`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eTgG+1Fnxkk41doVFRdnOsuUtU6Z8QFizpmi4XijTUdInvFMm6gzTNGwOr9dYurB
AvNs6I+nJdih1OLlo0EfAqLKZdhd0FyV0dqxjY/13JvMa0UcjSPUe2MHr/EjjAVz
Laj3qIhmggAqVWpQIbXUXPaIGvipeAq2e4owKdvzCZqoLzQpXeTYorUZ8dHBOlWd
omczEWI+GIxyEYKzxy6zjoNNex6wlWI6ZQaZReTLkILneZdwrkbe4MgCgDwjdzYw
qBDSdwmhixKeyqST1iZv+QPijQZCRUgv0oBHWYKpCC0A372C6hl7lYq9aLD+IFnp
2rV3GUoPDjy3gNeyAj8gLGVh9vzM+2+4O5cdRi6nCb8kxZ2wQJTpoamIoLlyywKk
H1zZwhKTRBVFCPBTYlKz+MG7F1ylSYwM+ikPaIwRSwLXgSwuhk4F4bCk/TjQMVpR
sDbp862mIGaDFEQ9LCci9RUwwgopCIwVCYBKsguH4xGUYwz87vPhlBz4XtWq9Yrs
ZtzKHnQMSTSR/+l/LwtpYhiG5dDepnHx6PgFmYk5pccp6L0IMHD2g/lHsfT03cwr
tYvOV10iyqpkv97PR+Tet1cGb1Mw8lQsGg0uGENoYxQA5BtT5g+EKHSnwam0lxQd
KBGXdotO4pLEV1KaEtld2A5MpK91h49Qc3dT9OyO9g1meMEMaocl1NaCrf51UJLF
D+h1+EL1I4mPP/fCQAXrRsi8QXv6bdO0E1kD8cJL5uipYAgkK2ms4yIqPeafRO74
+OFrl8CON4VtIei0AcamO9wl/s6LWc32wQ0uu1etdy7ymx+B0ByhFAatE+obD6hc
Lno0LQCjaPyEc9We9rB20aonU/rII4Qg+zf60D93mBEj7HAK/xS380zFQkttpYA3
T1Bk5X0+CnUk7K/MuLD2uADlD92cSdyvQcWZQu9KbnKR2EIodTd08EXlG1KH3FBn
DvPlckIT9jFV8cihX7u2jSHW6l+1njLLX6M7ec9jFg61BPLwBpfgfAGDE3CRYorB
/9R8dt+vRKjp2CUSxisP/CerNf3dnIy243uHib6moLqgTwvNrAB8xlaww0gHdev7
3JpzYI2PxwUY3eLps+3hN16SQf678QNcSW/8OF3Bn0Ud9TLw2P/Ip00Y4mpg6QO8
uku4qVGFMVAvrrJ3Ankm0Gh1xlqaQipywvW7FTCziODpzoDUmA1gqkxxUsAx01vs
5UjVd1mO73cqOa7yYvMAkO1vF5noLnonX3Svp4NmTZjFj5bTHYDZJz2hoemlgFQk
qZl/ispYUOvb3r1+ZOLYXQ6qbkXEc3pyOrjVJh0OXyVCsn//xEqHIwHAqWZakNGf
dJ6ssJLaoAjjpwkThUQD/BW2x4UtvxHsyDVpd7w/AE5bKItUrC1fChp4lP0hAEmE
Fa6r4LMbZFs3J3XEoJs9dDOsYQq8O53Ec8M9I99urGNfppgl8nSNGfSA07oEYNpy
qCRIsgbUWdJdH6p27QCxu9YSI2bQQN6pilBbakTHDUEJ1NfeWaIqRkp6HNk2K8tk
kV5E0IfzHImQL9aGJXC+JXQfIHN3zwsC4c8FahdDeFEpwHr6PVNlp8GBPe8vEsys
fTVF4IOUSCCMjSl9Px2cK/xFJsD6GJOn4TPeU24N8QttN16CUqaS6QCyCwneyZhq
RDBFYZ1ugAjVl+K4XGsSLX7q4w2uJK0uJqu2j8Y47NtmfuPR946Md4hWjueLSN9q
4yVAsfu+TxJOUnWAudZVT1maCtFbTTtGnopX8TZGcPjzcl5DDyB46+5dLe/sqZrh
Xrj4oNozJ5PZIwEFqmVIGw65rrBT2ry2jyJaIgZLyuqU4o+eOZsT6jgAaotKiKXz
EN0IvKhWXjDgU28X5PfFNk4EtKZ/588uS9Ijm+D4nI8ESyWwpAjD+v3UAuPPI+h7
KEzQfyWH4HePsALJcxQsMZiJm3Ha+YI0Hwaz7+EENcdEo/pIj1BzoCX+0fwmkPia
WVjDMZozWimyNJBrfwGxZcEhUWtgWyLOdfW/jWnc1UDY+TMxuJwugpO9h4C2cgJp
gQvfpGvdRSKfM0a9PlhK13D11RslfEevq2NuKhNRByA8b448P+OJlPhriyd/B4X7
0kdPyZ2tSqpOU9kxvGitAduQBfU1K6Z68SJ/tVEn3coI+TkoM1jpYP9Iv0mdVh+F
Mht7IvIGJrGK62bxAKvz99D35zG5veJAVYBLznEj43VfqMHKPnb0h3gJpX93GWjC
ARiRVryYBG+8BBN4wXnVnYF8vbBoSSb9PyNhFabFGE1AzwQQ9RwBtT3fbQviLv4d
hygfOA5wyA7ZYZkuxwNUQaodhlpAX70WdKKkRARcs3WwSWdy9ZjWg1vDgHESfXwZ
UKS3cXELu7hfc2jnv0WWd9BJ/hniAyQi+eahkn53YpIE7no62p+sIC6YyRuiJHMF
naqkzWX3OR5Ae0VWthpFBN3EhtA5I/uIJaNhH8TQKUQtrhBumDTkt3QnMa0uVCKk
ODECZ9YaQiMpb6sH0Jwp3rp42x81LmrC7YcIgTCPzV1t+/mS26sR5JYIcMIr3ZGn
9xviFOTpdtc7Y7YtKfwIWWe876PlaUPyyRhYnIJU8OTrFuAuNEz+EtKkfg6trlfY
HxFYLPWlZ6LOyjGvxP6oW/6R0o1XoPJP3jK3Qp7rbwkcgFheg0mRTbKhAqIanz2l
rDrr/Zl1sNT02DeZo7sqAAzII1cUnabtHjofcWIvTse5AU6A4iq1YASllam96lXN
r/tQ/t7j5iWvFGxyZtI0+bkbpjoSi5CNS+OSoVyC6pQLlm19L7fesBWreFAAYUrx
7LH0KH/HoYyXG4QrWwu6N9b+tmLhK8wa57K1XdsaWaksmo+VlAUbtDYUE+eg21ij
XkcyqghDtT4/AzIT7oO6Il34Gtg2K7nYtWoCGzyaTEOxNY537PpJ+G6ZElaY7CIe
xfvR5JaBuo1u0aDgvgxDpFFC3MnOO5yzFvBPPVk6cL5CxM+pBCT2XYWN5oeainox
PClu3H033KGieX6gMONgEY21q4lOe3T9Ig0eYZjewZqM//nSRNCQ5V6cYYTvG2Aj
nqiGaDvIQJ23yov9GqPeqzd7VJpnpGl0aleHzJKLldo/6IoQVriF83eWr0dMqeXn
g93QiX7IxlPF3ktwGXF076jS96rooxyxf7zyd5iPJm1J2zWDOEErdMrNUwAqrgxW
Nvfc7HRdLnKipvcs0xeEa1yw2WfhMCndD0hJ8BTXn0Dn0lcWQyONCKfGiwn5MBzH
G15OY3ZD3qDyo55hdHb9P2qkLmuU8zNXsGtAugFmu45XfgIcOafiea1kEfuXeKs/
l5J8DfIbUsS83PwPGqOs5GQInvu5nqTc3DfxWTTCPMNG12nKnWnrHVKJnKiGzlzz
RD/V4dzpaPUJk3J5VXNSvZfdbxe7C0tWUAXvqvqYTlDg9PsFmUQIL1Es/7o6VMCI
x6KIOUNuG3seUVEPXIyHZZKMO1h5/1tz9H8N/QHaXdMHKwNy6HLv2iaMEHfrlDJD
JrfrMa0OlQuLvAW9Ai9aU/JeslbNNmSTp+w1cOWLd6kZkrYikEY6MvPLzo8YcvDR
goHMTg9tMTwr0bhE6kEPcsjdSFhBFKDGkFX00Jz9sUe+n9UFeRgcGIBSXOi90DCS
+8/aPsWBKxeUmhKjeDQeTuaySvTstEQEs5l41hOz9uLFxz7oHwA3igTGlWQ3O2yf
cCJje8oMwgNNNy3ORBE7wkL4+mZCKFWNe3uU2k5kWDpp9lKzt9XtCPknAqxXeQIQ
tihpVS8l1VamqcWb9udz6XQMjG1bAuojxHeqsGM3rm66zmI9v8yLGqTSP9uou9zK
2ivPJB1Lg8/8Is82F3laJsjgDT1dr940MGi3/c3aRGY/rsqIpcMgeW7bscD1cJB6
Pa9srmmeFgqoxNwrsFKLMOH9bweGToz0t+DND9kIimghlPaJU7qrvlkbaM18OaFR
WJh8zQEKeiD2LA4dozIzfRPUVA+DKHBiV61sWs7pp/nmOxqfAygLw7/GC80iDEVi
k+AURFIrrG4dguget3YsQETWarxRrGn2vYsrOrmq/Hq0EoYe2CJLDwH6As6OmSey
YYLLPPrHhTKOrlF7hWKqPLFFu+xKUZ3nIKxY9m+yxJBLxCp3XqcX/BOM4wJfCg+L
DWe/pavxuXiT1fqH9OHPIXzYsuBQEDTObyLvLb6LMsIfJG3B8EdlVYvXm6QVhQwe
+YNJRQN+FEIAcwFuZtS5A7GALesSxqQrUb0u/9ujjloCdJg0/LGbroTfmN4yr8Sy
o+LJsGT9/3SeoryvWy/sfJE+ozO0qmKOvNbSytOI67AE+L/NrUVCFmzvFetKuxD5
8+LKhbp+1hBypQKHlRqNkF4Zz+PJkK4mPwKT+Ujw3zW0IOQYBq9Hj6beun+dmPpG
YLbK3dNuzC9vjXe0WrGs58aVXPgo661SUnrTQTzA0fmMHvdX6PVOQnt1uAxuzo2b
NaEEqmFXOsO2ZuIUFIOiCAnowtyRKWfVZ63t8p7pftx18tWt+9e6jMk1/bpuRwGs
2Ru9TdGvs9n+AV2GMoA0bvUOhkewfWcZsCU/8jmncuI0/LM5+RlcGBIAnbaRUC6e
3onGnqcOXjBqBPe1PypISY3AxXkJoEcVsHEQDQVv1R7nGXaiJsLKJMNzyj5aTVYt
JKTcERqFGjCsHVKBZIXK+ZMgMadDjzzxV1XvEm43tb0K7tWEz4XLlPDCuG5KiOSE
ZZmaBXKENlW7Yvf2Ejik2XAurAM3T//5DNVoiScnYz94ovWdYlOXs1DrbRzoT7jq
k6DIRQtiI9delXf+TLcsm+PKPdsiW0p5hsmHc+gWKLbZvv8479ZZngWuh4YCYdcb
KusG4FtHKMVIjtlballd7nu1VPYP3+AZzfjdLL9qJM2J4yOL9MqDN5HTjBtfwa7+
DS+YcmpOT7+y1gobJrPYl0SZzsTOPeRuY8+SIhyvnAwfRe86J2QR5jUfxGDuiApy
vyX17SMvoH5uu7iBCP+rju9En8LA47EKvyIemRsRYS5DSpJQ9Fs0HvFk37HshICv
X2umwxH6M2n71kKvhXTYvckwGrlxbJFxWZkTIpuqacumrmzJ6WJXkhbfb0fEvyY6
P2Qt0zxFdqCGB0oxnHuRSHfkmjWnlD4o3HfIjUpDVAOCoN+Aa4FNd+GhuFiGMYA+
vyqMBIRRc3DfSeJEhYfMD0rLguRUEF4bDAxwgy08xWJb0GGfi8dAcNn/8N7wSiFv
iI183ZbvZEGkZ+UWN2DWUXhAoa5I6sSjj1hD1LwSeqabxaAYT1pT0XOwMfEXPXqI
rZ1rSlpUcUMhxuYiOkt49DAEZunuP9ZMGNCD9do0Ic40LQO4Qd3jA1S7QCGP8Dmq
nIv2Pt7bi5IRmAhOLTChfoiectD+5qcJXZAm3ij0trXXe50JLmoxn088Dezaxo+K
6GVfz1j201agPjfj6ooeuf0lZXXqYC6pYeucsJuJCUEKeqtQSdkQ30FZpz1EYxi6
Ixe4zESjwx/n+HeuBVlZ/WpELWezAnqGtnJC+keKHtgLvKlsPezZHEj6ZbguM0hj
41z6qBHHLbwGaMf1LCGGa8+MRHsGY3LkY7sAiGQw2qzruXgaURyCRIOUmZ/B6byp
jPcrruEZP1aSGclAJjz10lUDq7JOtqD4yxJ0bYXfvKC6jHwGWy4Lc5HC8ZMUDGX0
1ROVwSLwYTTV0xjig4mMgNrfWohY9D9DZ1QOO85BbGrtQQ0dNUdoJ49bPQTMmYEQ
Mk+Nc90qFCUIdVJTJ2KTwBu4bcBTWbwjyZ9ypfDlV0DGnqjDj3LV04alDWOIwtJR
cAi0om6lyWSqaatyFxwa9NnBg5q06CJ9IcEMTKHSk6Ulre5acyy68qWtnVivOXR5
Lti8iAn/CEr74BDC9jXfqXqmTXQUueOhTRuqibFCM8wWAOniC0xRxyMNMMbTtPEH
ABH5KSYBvI+fYDwcuNFMnlU0aksflkCZc/FJBKRukUlW1gcb3Wa3xCbVqzXA+SG1
8ZWxErtGj27WaprEEeYWpG9oMhcNHAkK1zUWIqYCpAkhNTIQch2OmRkrxuMs9nfp
CqWPPEu7ZKrabfE7HE/dHZRpwv5CAZneLVhLw3p9o5vHQMKAfhlBjylaLvttezrH
FRcAm8JlXz0WFJXJD0+IV5vRzYpkkEPJ5P+Q1m+sA/9kP11yu8M/NoIYNFFLmNRt
47HWksnOB3d9hKWaRn4OSuOgeCQWqZxf+LwvWyK1shLQ9S/aGayrxBXCOdnBRHgs
RTSVtVhFLVvjcwCvslVAfdil1n2+NiM5HpKf9P26qNKA39e5jA1w12b3OTQKurXa
NEOwk0aGk6BIuArxIH4x4mX3FzkVBtQRExLmfVVxhxY9VGhqLDWqNTWJReWTZZKk
7gaZKq7ktFzGiF33xDFSlns2Y2e+7BnbXf/xRn7n31itmmwPPai471QzR6pn9Vb6
N9MIzb/xdT823/fZPFraROrORpX6pfokuUCe5VSAd6mRk+grJMp+quGFz55eUp/+
xYbkgtDgPIeeQ16nnQ71NFdVfp5fq+wr00MFWF4uO435jV0KeywiN9AXbHsSgbpo
iYse3hpMyuAOTLN43pNd9vt2AeJTzXB/sbXxI4JCpOStIcAijUXfmowIq6yqjaIr
znT0l/XlxZpb4/HYil6i1WbtJx4EyHrsmi8wycudR5TWXgSy21Gc4tYbxeZn/i6/
BVLwLEkNTIzqWFoSMvs2vX0cU8MTjcCzBpHSj2FBMT5VMTpNcZZcXf8MzuBsdNPj
t0vADdhNPpW6RUxm0B8YzwDQ9ajA5UvnkuyC5YSWe4Dv2zf+Nx992VLFpfbr3/be
alk3k7UdoDCY+QaenKZY/vRW38hYQ7OY59BFF5ayxNU5vkZHV0wyPXgCS0Adpm6J
WrCg8Ug38CWek8ZJS4GDP2lTWWErfCcLMi3GIrZbb+PSnaZrVnTMij3VwsW+8d4F
ozI4AFas2saludSXOC03jOUKp7HZFoSVMJVmYNcO0ZBsFMzo3tgZ8X4pat3IPNlO
SiQb+/hsBtczrt6pspfOrMRFsaokl2m8ziDS3FhHFbOMOMd6s5JQcGDbZ9R8Fo48
5RD5FpG/G2F61V8XB99zk6mZ3CPydZyzNEs6hD+G3Ike59wzJ3E9UEZCWjf6RJ1W
nejSHtrmL6Auwfbf8dPXbPcpmf+zkNotYjzvvuP0E0ik7RXGre2eaCIvMUPGqekd
Qcch8a++o+GqYeUixoyfD5wOQx5oPDUWynNao4eks3hvoHvVX+jcKGhiMsjemgOi
9i2n9NcRInPnZWXWrdo5cpWABLycFtDF98X0tjhsu+czZxWx9OAaXtJNHxrmwgoG
7YSYOr8ylkug0N7PJfDDf9vz26UWNc1wat9ZZ1mhDjLtTeDntbXMZlOxrOGfFHyK
5TQd9sGvf0TS8kKDkH1vlawhyd9DYPV5w6osW230yE2AgCr0aAScAb8RjRq05r75
MjeJg+ejxa+5yfE9Ish0+B8xjF9BQIp5TrLq6E6cpkS1foKjPFz252Cpqvu9o0MV
ITbA7PR53jYu796fw2xM8jUNNln/6PgJQ+xfFMVL9UpvXEchIWtpBXwhe3cc0nB6
QDlAEwCMcdCMQp1OsGWSq1tbm8V+sC4KGumQI6SQyzauXnvewUrq1gvxaHIHJv5g
yeqIpEY2ao9fBPVHrO4JBJbsxncbvta2b2T9g5cVJPO8/WK8FmIX6hbyWMB8Bwsx
NSzMZ6u5QE/ZT6KFTV1Y3LM9xugZ+KVQJq1K1XGhq1IE2PWA5cQA+d0C+f9NeKSE
zkGO5wDNvVNBZ9O8KwpzOmcFZtngoiCw/H0jd6fJVDVF11T4tXtk0tHWxBKhs18x
3131h4jXimx9rOtClLxnLTwbEiz3h8Jn7kqfp+eo+U91aK1XtW2pfsuBkBkx0mDt
RjqwejCVtAxW7jaDPrV0nu8d/rVIjEB5aRdYILekgTVM7pOPn80FHJb8u145ceiF
vzIw4KfuTIW1sOndZUsrko3QxdzBK3+4hoFfKdQrCjq467FrpIo1D9g7JZK9s/32
tiWyTeEOu74548kX6ZaD3FA3gfjja+MPc1xvP5517buw4naTP/1KwKjyS8yg1xVz
1K3T0+TFvzrfIPDa90DrxqPt4l/t6dzMxEPycxfXeMSrp0QC8e+xMRFYpfwCMERC
Z8bX4m2xaTKHaERsN7QEoeVnlsbAadTrPrejgRZ1OESO3X26MtEy+wdSP9IMS5on
V6P7zZji6R666FsF+jgRAHxXOcCmPUhsUxUkvtdeYBZRBJ5bjHoBVb3ajMtlHyXo
lUM/E+ccG7RV8lFNe6jYn8KGnZrxxTYlC9TSurmOYU8ZZca4j2SHD9B+pUc7/Oqs
JS3DkUbIMSzF3TGWMlcJSKI+oCQD4NRxT1eRwl4ONyvVX/PdoBYuc+DHOIIjwDpP
7mYMO5sL6+wlo0nelZIa61uPtEHu4w7DijfAOoZEjChHZDpxeA2XLkCayCi6wNFb
12k3/RAllaCNVw410v52wiW+fAlkg+J9Jzhrqg430wdIJaa0/iCarthBEfO++LnR
E/42f8gynP/Mg5hm9+fqXq0oqdQav417s058SYNgQbg1b0YfiUOocysLF8oohb8O
VxWi2dQjw4ksDwC3dK9dh0BnF5Ag8AojoAGSJQh5pmCv88r4SHPn3ACtSpz49gN4
ORsL2xRQ2RTNaMsb1zHZnr48KvComicbEeLq5Emdo/pYzAng84v81nOyVVPoPSK7
4PUX671XOnFHNdMiUI93uD6wDsgmA+uYSRlBRQmbatxhCIgdGVE1sFEVgrE0Az1O
DrhyT3a1M9bUUCC+z1IBJ+C6AT1Mr4/rns8FyFGN3G/q2552o/b1lMj4X6SsEhmX
plRZjsfL6qNpbckDU+R47XpT/F0IaVTkUWvPtliyeHoQrVUS6gLwVc8MIYrHZW5s
3f6uZr+VlnXWZyDk9i+JXp4o3rqSy9dn58ShT6saoSigu2EIrEuqILH1BxtL3Vs+
T8NjHkI8ROKGvM1ifD1jU6oRLO2HzCc8Mxb1GkbkdMA80G02Fgmi26ubwp6rxHPs
Kv/XplK/9WMUmMPPCXPj5CXRgkBfz79M7MmrextbRCucqVSXuszP+aWzXRIu6bYE
HqL57qbT1kW0d7XHpP2fsRw3GSHHME19wxqfU1YIkF4FDNom+IazZCNbAq9cAIMk
5VbR3vIWPgu/lh8cZkG/bxoDN3FuvZb4146GZxpZHnkVEzBiMEYQcnFm8MTsttR+
95lSi6Erk7n/LIdk/b5YVbfOEW7kWA0DnwllO8cEisBI/dMzRBs6MKo9esFRDaVO
SrrphsCCOBBJqdkPLxI8r9NFqco3DpcDeKRgXxIVMVrka3Z8cwwr9Ul6j7aeA2JZ
S6wBUglpWTNd2a51NSst98Ty+M3yXpAGnbD+vKHZYmJ13SbZypQVky0JUmjcVbLh
QkZ6f+NRDCYaZfFPd+4+MhCVXSAl0/SITwX0/aK7ciSsnFz4d1TL64/1ESBXL6gt
nJtiHts5y/lIB9WTDQBRoB9dnDOlTOphViIoTuWd99poh4n26oXbBhfoO+rGqkZ5
wmgd9rBf0oHDIE/tc8oRuSmnut+JjCkHwDfd0rCgmZQOJzxtwe+vi5joEb98vNrQ
zecQ5N34rCLPHmk+2FV7mizjI6YUJ/zwufJZdW+TvdpXRJ0xNDgkTce8wZP5jfHZ
3qquZ7FhYPWBEcgfVng8BnhhvdEX6TMERQKf7UkoK+sllWv+FUJ44YJcArxX0M6S
epo/RLR0VzwxwWQaG0Wbaf84hs8fEq8vWF/lJb99t7Dy2SIwgUYyq3w5sZARvQsR
dTSzL3g2JEiQIKRVPqKWVpLo7mWVuoYEw0SMQV+gnJ01Aw3d02TJt7P/dDJzAd2G
ShjwZxDFD6+9FRCkQ0GLXL8OSPx/uO4hXz8wl+9PQkQoJ33J3YJ/grIeZKKixo7B
hEjRmIvHsExqmF1FELpvTaooZleJy3QZZq/DjiqF24hJhys6hQTN32d8SmP5KyPm
SFEu1pghBR3hwPN0CvKHd3JaX1ObYemGYWhDpZoI6Tapvus890eQn7bqNU+AzbaA
Lg0dAgB8Dty1nW9tmY4Vc3f/cIIInUg4YCJKxffmEDNywtuuNQOQFdpNQHH8GFqC
PobbHBXcwGzURFvtSr1BZuNs+/BsG4TFDsfocF/QNK9gUOERosAZDQ9x/VYXiHA4
mFi4qOC1rCgrc2cLs7deN0/52nVAemBBRQXCCZYfT+94GfERYu5eIoRwdQ20vZt6
DMSbLJkw1mhNZTOFUA1v3bnnYo02wO+G14/yhXpHyETyTPGRwOzJNyfWDssEWHUW
wRPiYKtnEvjbvofwCfMPU9jXKNPU8pTTT2DNmF7XS5HP8YS7jb+XH+CwDqS/+ZtD
qp9loa1KzanvjUWx/aT0nje/rNEayU8QLhp1DdjWa1hInK0TCEhAyHMeJWTRXWwf
uX48eZ8vjQW4W/pWyOsoDmEqwOWK/1+TI8ZuHItE4fajjOH4jgoVKh/o84a85bn7
B7On4SUXrRRiMvyEID0KsVlDUTJ9f4ApiqalEIONb+dlHXqv0HWq015RvSE+1Rjd
uoalT5NnIkOHwvW9va3sLEmGdYeaS36BHp+zz32nAAgIcrcl62aOxZ4DhPFolR16
OZ3HaesMXUfrN/cbJL1JREGrw8mnLrRZJHSkvH0RsBXLaK2KBSmlF62VFPQ7UhFi
1rrByGFtNbgyj/E0GQ1nE6cUyYNeCtNtzvOxLkYT7Y8JjgUWHWLA2ePYY0UoOAQR
oSjPC2waJuvdLVMAlsKwIcpksVwez8ZFHdla7VJuyG0Qxb3rt7jHh6rWDM5VMQ2V
opV+VwAea1vZHa88b6CM+wW3Jga/rim4z3ViMvvZea8KSjnKn2+PwLgO4JC5DxnN
qpH1OqnI2ruAbK8xEIa7/CqV6uOQvXco9RbFSne9OK5qzFyr8uaG0C1zhdo19Syp
NwtJgp1k3Ld3oV9blnDGRvo3mGdJQJ01gZnqpgddkqhMz++MgaU1YKVc3q1x5Qef
+zCITRNJIT2SfDTxCp0YGnkW9S6LeNSXtcZ6VzI7JOEK7qplV7aIJHC1eHAu3ECs
RynenLrfLRFuprAspVKEpx7LRo0hJHrUOsjK1oI/zMrpot1ozjf8wOrUqjCCjHvn
d/cBVomulZuvADSTQE/Sq+1Qxj7QCQpaf7K9BrwMCQzsMSqh82DScD2/qpV9TRM/
ZHaDUKeXkpqwmKbvtL7ve8iv6cUkbMTHq7s+U3JfDQHuR+J9dB1Fc4G+8nwq7G3t
oN+q+Ix4PALRz+yJ1gr5n4VG/8A2vdLoVrJijFJDOo7aCx/Dd6XLbb77iykAaynG
kM/te4ogCvvb85V1UsrDfy4S7hp8LNNlB1vydVRsgEwACQIgfe7sciROcxacs37h
Wobj/TvkmmoWd92xmXwkteoTLn6jHhqsU/ZyofUGzBaVFrzgFnHlxlDhciUwF3Xt
/+7P3AYXDL/xWgyc1/n2oheoxgsLJVqTwRP5vxooSsQkRdIvX0sQRDmLouAtsCIX
/uAGbWBuU1d/RYm8wUbHUu0STzrabW7SEwW1oC2S65hGgI7VjhNvnh0PDShbBWDe
QmDX814KXYhGmIxjM9g4HsHD5V2sFUHjbAkc1RmdORdvhBSXGPr++33qgT1RpEfm
IiGDQzZUZk5fYmogmg7ORR2DMY9Q40XDPzacIK7iV1Z0a3os/xF6tr5BwhfS9utv
v1l9zCrywkjNHv2hhTQgMP6aGXaFIJKPJwdopUgrCWaJXpphWtjMBJklLkza0tBA
ckUk3xCS4hcJ41PB79UDdMkfYhhIs0BUJYMC7s6fNmI4CkbgzesHVaueWNsdEoLA
kkCoU0uaETn28dNU2LhSIzRhybtLJgzzV6jFU243w9uDQeWjktHOHZ92j+AxSey5
KioKouCJueY5AMYwDqUXhM2LIrDa1h3yOghc0h2ovx/RMC6SRxwR8+n7LW6Fot9A
qtEI3U5Ch8bFfqFm9JBu4dvlVlcOKv2cXh93y2zfDgTRQ03aeYEgsqIykosBnyno
BAKONJ8TuVY6yRFk++qOM7A2O8z9xTlXA3oReB2pNZhTLV130CpcBvGhp/unVJqu
JVQQmfWEVTJonf9aDsZ0PrLgduZdtHxuDINLe15ZCFh/lbIcbSvpJ3fO5iGamQdm
qaZ5ehduMngX86KIRz2ZakFB8BJI/WzvIBrnptbfVg9fhIadGXjDAC+BirQX2zgw
CoIdltB/P8PHwTX7KXpkbvJ+0mNpUKTDnhmVkME+lo8I20Df6SvD3lGMAYdjxaUM
gw+bdZR6RLbxAInvPMQ0ev4Gx6u31eSl97W9FW2NTsFcaWiYJoNtnr4s2XNw8CL/
u6Ya08p/A66PWKYR9bKOH42rkOQfy9ScxUDjgxK4irPZysDo5EEYYBlk3oZtDSHk
g37itmdRTuAJpU8X/rw7kuXVinTgioH/LmWRReEDwt38YJFoQkdR4JzLnncFtFlg
nPVpIL32Oc4wR3WwCEyNTPO9/vgPHL/WxP9jq/PMG62vUXKc/DEbFy3WVA+UglNf
Uho1ackGFniV71Sy5VwIwstlYmty0iLnqB8JOg9h2tLg9tCbtm4jSJyRzyLcbj3T
RLmyvHaAB+s2tQZgh4T+nM3iPe35MtqONNhOzxFy3qVOV7EbB9aawROsOWjaD8u7
hhbsdj6M3Exi1Oc4TpPFpTQYfMOER8nTbC5IafCbkFOFJw8+ewd5SmERfDxVaM8t
JL83GBTJMDx4L9c3Q+KsmnaUktGLm0IFKpo9La5xyXtS/c1VDXVFYST2PmxeU3Le
S0BbLq0Z2yekzs2KrpGSMZsLjMtQypxcHu5rKZC0QVi+eHbrarsxrzjhTkr0cai8
pQ0EqVxfC5RfI/nP+lJh2nUR/ZZy8kyTZ1ODMLOD3toSKTi5kvV1JxsImMJ7PDwQ
ZVQO/TkcRe+qAQgJO/dlRVjddqkpc7hni8DamNdHWSLb5d4OKTmaAGLBd42Rs5yQ
WUNVJMRuHrpG98D7NOYIoSKFsdUuBCoYyX27xF4kAbE2TQ82RP8emf19/7HHaBK+
w49iMSu3YsirFn/dhnVYELVBRGykfAQGk2MZk+plPpynNeoOdVYbQJYknVVOnf43
BXNtm0MWLRfT9OY25qbuS8st1k4/oXZuiMA416qPCOLFa5/DrbOOTCaVMJYKD89Y
IyAkBu6FTihjq6jBae7rJkyS7VaGIBIktFVQYLuiQutYzwf8EVmhNermc2DF+YAp
KqtdOXh3yYWLC6JLLxjGbQlVrwVJ1HHLynflA7TJnE+M5OtITA1DWXIED4sfk+zV
zUbIlGFKQaKoalQphJuNd87mRULrLCp1Ms65yQoBOv7X78DStHdIgxdPng/sEDxW
zFXLEwk6s5QViBcf/wmc/TwQY51Ia1ZFPg5/xxeyZIA6zT70Kxr51q0n8bynCoGL
zdSzExS/8tLr/yi38QrVTE/aur4VFSLNGOL+vmVoEa7JaTAIayik46locDGIPhim
xuc4tipCHSacvakc0bI1ewuXs0Y+Im4yDmZQmYjjSW2VRdhkmghJAjSOsVE2f1FZ
w9oIafc5UUW2FAPtYbq3hCEj++XNz80RFSLqXZjqgt/SjukvPATPaTqLPRIA8HPy
T3fMI9NZsop/fmpJ3Ez/sMpu3z2APwCRUzyWIGljLYMYbgNxN4gKp/D/ip5EEF83
O7i2P/pTc/WvxS7kcVFqh0tZ7LZKXpCU9nGTH2fzzDhPc7mqZ3fEoqbwbX+FBL/Y
/bOXAoRcesgPPzCK4gkKF0vXTSzgm+ThmYyQyHNZ2OUAu97pcVGaTo4DYDhiRGze
UvnrZbHh0rfn60Khn1ONCtsofAzisCx1FRTUJGXC+dB838t8kSsliDAxU6qSIqsS
i/LkEujwn53ad3rvzeKzpU2QZOuHNF1+xPBqCd2T+lt4sWkLFyek/aVaPiBZaQfw
rNJACNhdLfZIC0V6j2cnP5f2sBQDmqKlx2FLOzM024HK8yiu+aeEk37utMLlxFEW
qoYk5isYaDjCtuRUFMpGjNcAdQJEuKo+UxHfcS9Ah7c0RavDyeyZspeRGsZ80a/m
XEnHrveQutAM0HCkv20TktWyJ7LAlndBTGYQVjz6CxSSoVsbQSKINewrsqC0xFpZ
3kIFVb2lOPmTmxFtNoISZCRI8mcu8cGf6hsIQ/LnsuZmNcxNMEQZjtsNwgXkl+Vq
IGOqFt109ez81Kd9wira1HEPrV2OHdP24pZxW9Z1ACm214ayYSf37ruukhs/NPx/
0r+i1J0llAzIcWxQuUWCFqL1/lbAynm3LbRuBZmM3wwOUDnVyq00/n/3wVRI4sro
+Uqa4y/z1ZPA0a310akcGgQsaoyFGE+FNX/RqhQkx0XQq1ZONGtknjq5qIrKdOvA
56QECRWDdy0P1sJCzst0FDw1O4yuVABvgGnZiVs+tGHR4kk2NlVwPWzmb18PPqux
ULqRE9oFgddckXryq1xiSP8+QG9yWNgvVdKhOq5Up/QbnKq5n8lI0SD/XhoaUEna
wqhNTf4r9us7Vnuw+t3EHM4VL4AvziWoUUMlSq1owAFJTrYtc+IAm3qYdyxQBxX/
TusUKUrp0YxhkZrjv1Zsgv46z32t+xTF/CEVwIf6TMu20q8fgJZSXcShlCFh02fL
kNmXxz5d4orj7qJb1SQxQTwM6rSv0iIAZBSJfWT181GKOVc7zbsQvXQvjZdfYG1G
zzgF/dftgFkEXhHl3DEtffB6P9MJiwO23sksTTyypwMVtvGAfc+AdPW/enAqAB35
bl+On0Lh1Yrte1g/ybnADuozdN+pLfsahCTV44FeTxj5BLNa7fYD533PPePiFL1L
flDAPfchG4OpD3zuDjw1O7cI74jSRVqufzB80fR/LntldeNUFOnc23Tag//hX7wf
iWOo2l5OXBl4JuC+EwFD/shSXeXeSfMKWayXQcGWnquJdPeW6mCEZbL2YfcRipKd
h2EV+UqA0tLn2XiImd/Et9INyu0mBdNJrYv2K85uNPQ9+7GTAoEDKKd5opy3RxP8
HK6o/YE4ypJ2YyT/Kh+PcRQw/CpWM5875f2WOkGsVFV3611Emf3vO1URBepUVwx4
426v+rVl2bmcbycQrTnwsLgWqyzE1rKiNKJLCDSWffEgfKDQqJseXbGRS/vaL1NK
qLO8HjB10RPu43bmvf39oBK4qLhuK0IiF6iqpBAc2eJ3STB/rXrEkQyABxVOzGjW
tMzxgG7V6vArtPU1z/cU0KR5VPbWQaOJk2sq6vgLM498Pg06bUfEQ74x/np8ed7k
pfNsOZOafjv594ZolWhTbbnyn5oUfVtIHwybVFigR3guv9dM7S7UY2DQaXCagIyr
SbyyZ4y0bJmwP9AaGgeVPm2IwPQ2/ceXlee1m8kxObt2Nxbj7fLGU0FqbrS48YM6
dII1K+dA1UqgDQlpEpAVDlQvT9q6680T1Eq108IUpTq3l6lPDM29B3JnsekULrIs
/kKMUyksIb2xJU2+82xhir69W2BxrpN7vJK1aleMVvSqlosF3X9lp2cPqV6UW/xr
6KQ+qXhJR4XAkzZpMeXHy0iA/lwI/tvqqTFTxnzZ1DXGxCDb7Mz/lIWMzedqFNzs
nidO8VEISuSpujGc1RBHFztfZ0hRiaPn5tVosyWgGblJysV99LE37UNJe/R3UlBG
jbdnE1WW2OPoAx0iNxmgeTTCRGO1C40NQlmXms77iRk8dxYEso2eCNKM4eGGwNGJ
uaPst4pHDzBslR1nSA5+4qroh8S7cAWioxWjX00g/OEKofyuGWvvHreCuqWaOG4s
rNHseSZonDD1YMxWwVo3lvkvrKsmIgNLurM5OrICHFjrhmCuZidh2moamCg1kL4w
j8M9u9ysHhHMqpPXlcoJhhJ/ZlPGpfXPu7ROPqCkH5BEsPqzfpo7/4I2VYAw5kPH
q/Q0ZsmLLyrnPSEDFvngfEf8G5RJorFmR4fqLqFJwXxPAV837aNdCGlkNhdXMXej
xkaOBh7LJYts1T9y2DwM2xY+rgbDdHVBw5vbp+Uw+tHDH44ALjBWJrzPA1q8jpTk
vgKr3AGq/Tyc2V3onILMwHSwPQsrKIxat1rDiLT3WQyAfQHP9OpWH57XGUgUo5UF
2go6a7JovQP4RKnvesZBhdVv4XBGsTnaUaom1CC4VN1659UgSXxN3EIAHvqHxqvZ
GovK8uu8UiwtRYXCasfjYV1O6rYnrJYTgltCPHgwoGKFWEgUvDPxBG3GzQ2d7Rrt
BUOYhBXrs75+v1TvKNEK7x1Y/rOpwuQhgip4PM3OrmKYX3n1o8W4tVcfoXlpfuQA
e4yODpx2BPPW3DG/1k0qJqgpKofGaqHTOpeu/2QcRPUb0wySJT7YX0mbH4QSKk58
bm/6HSJ0J/4xGbjdq0iQrJiKbMuIvmnPV1lfAwtib46KIw6840Q4vx7JxQ2ZgHje
PBzU2AjYe/zJmr2m2/d5X3KSbURx3o7bAkzceCFA66aCV8VksMTgiOdc4H37w9yv
qGrIe2PGHHDKXrPr1INhZwkY5nuzEBmTx4L6X0Eybk1QELle9DPhZcLRYEhNZChh
MEACE/rK8LM7uHBjigDZS3uRX3dsQmxaiWKFHgCPmR7Qu7ynHgxfFyk8IvYTMIsO
vXGjh5jCRJWHPe13JR9iwoN/Bz9fVSqGNELfHtzOSvwMZhMSzV/mX1vu/pgbpFtT
Ma5H4t/Woef6tLn4bUJXMMN6mMDSvQ1WXu1gS9WHt21YSsaRjsUnG5m/yYu/yskP
wA3OexZIDylgACwGEdeWqVLgroaseCC9LSiZzhcLIWvVDLv+sD6mXS9MCybdETNr
r/20XhDI/+pa2ph6q4LqJp5OPXfTSJJbNLtDsI5MOCKzrnjz8wSghyZH8RHo4Cef
oixIafcwUXAguNlmWXDP2fPg06yIU82Huqn8rWHeEvjYZYO8XwKHoKVmUNpUhPzv
tOWx5sfvY8pBEH8z8xfFyS8kWjXUQIwIea5y6r9Xu/3m+aiMePqVN1e31x8sGcE3
vNmTZoZhdJtY2DI7ykkDespHcB+neNGlcW2mbpfLQdXP2vEM98jyNY4cY5/DvOK/
8rohCbt1HRxCdyKDQNRrxjsYN5fQOZUgPyjbd6dnZTWY4HOfMu8gvYGRNKYcjN4H
5dszQ8mrjSzTiMC+tMxkhltghq5HBk0Oa5bwvTFXS/oI8f5R11jGOuhD9pbQxkKP
W5RTtQ3cYnXGvjjFQsWIV17O44ME2hdDDjVMpYgYXuS1YmN0gwix3FBCWm7czsZZ
9m4xKGU2zM5VyW9lP/3ZlgrIpx1+iFhi59fG/mD8Fwdu47B4vRENF9OmqWXJ7+Mj
yZelPMDKheb99pjkxBaLOtMMp3ADBkFcmDCv+r8ZbMcnf1SSGCR4egCROgsggBXP
0mszQ1ftKrqEMGQ7dUqGSORh2OWP5CqHNqsCiWvgOyzRv3On0DzujDMo88a9ac3t
df3FsH/1jG1DCO5TUaKyl1bsvdjqc47jZvzaSenNjaMFizbNNXQ152WxSU9TxtFo
tC4linzYN5cNx8WGh/RaalrGDUrOr09y+skPzwBzETbf8H3XHTCKPNkav8nT00Pl
3JfMBNgm95kRm0s0xsk5oIzLx6+xRrI2si7UMsjFmBmC8t2nct+hmwsmErtHuwRe
OUGp2+k6pESM2Azt6kxTE+79AIoWnrg/HXRbXbASrkyxDdFhOIk+PyiBuchyl/hE
nYgCA/QbFLleN/eUWgiLVQ8klDHeHO6uwmztyG0J8zhBAC719RsRMOluIcSBgiYE
Rk+AN9fiKZHfJ1BMIMDAhsAihvHmH58qYG6StW+hB0mTzy3JF5ggnALNKRRiSZsY
ir39g9dgfLKnndsApYqon+rAWgyUQf0frdbWShw0P29X7HjlXikpYdgs/JcrsupY
dPbV59Eyg/BM51CuHN/5bVZhev+65LXcncIAORd/CwxY0Fk7mm3qP5ILLXgkzZnF
8ri+oY/TjDeAdo6ZhkHJphxjN8foAjHHQtoC+K46niVta51dNTHM1f1TV5FVpGb6
1qDDmWAzV2AyifiTiSWIYv/joEvhCbkja9mZj4Cx9Om2xtfC2K6ZpHM9WFlvKk6p
skkrB9/9hQ6iILtl4TsPGpjkWxi+H+8tQWHlGHCsBKPeLdN6uRrY1y3bXoQzQB85
GA/bO38ZTSi7ZEDiTux4jK0EpRR+RCkCIHw9/7cvgVFkKfXH8GvncjX88Ph0ev+/
BGh7cdpxNqzXXRMlBtBDg9BHlkcj7FwRPCeItvZob88SpRnYdMBc+LwPBljoT/wL
tuL4eERPjWCWfPa+AGeite0QzwqF6HJMXXj+PbhkBsQ+OdwOH5Eb5Lr5wwPhOujj
lEZ+CfERv00phbSqU2jMZ5qXTSj73SOTdkJPuoHPsg3wEsljbuTTIWjyt+762GC+
Xg0cwP7E6U5eoXM8sGSb6d9y5t6w3YJ08PPD2+h094DPPCfklDj/Gr2NXXJEFcxO
5IzK0sx/imeISdCaQqP4yL11kRFGRSjsccsz063GDIaScr21DCev8uYK8R/HTnuv
6HGV2uFntHaFWd/JrT9o6ohoUDiK5kKK+6QkP22NdoJgDHy91uhFoNVyhX2rhCkd
0NgoBCMtHvUa4RwWinmdEYFBnRsjYl031hZdoe4CNwGVXbprFego6cgrTqTcE0T6
t/R9CUAMN4wiReW2h/A8ewczybg18OQ+GXsUp+sYaVCcbHxsa4pLwserG7L0LYL3
byrsXNNex6KC+vrDzFVVnVCY2rA1Q/KAtrZhr0kMupn9b6B3GCLiISJI4rz7Qdcr
XjWO3wYqcpbQQqD5IP1EiguF+jMCmTC0a1gi8TmlRkazGcinK9BBuDLUqVTWIZxg
PoyXvXPg+WDTlrBeS12kZjet0M+0DWQJRBwM9Q2btUR2IGIlfEZmBiYEdDC0zkOd
Kr3HZoe7wpp3qFtwXmMm2cyPJwdWnkVyAQN46f7w/W0WUaVOCN1Ja08nZZbJ6su/
gUKzumUGJiXLGQJe154UGVtHQbTwWfOSmwN55Z6EZt3VSPwVpqBaU6deLQ0Qu3Ye
drKHI1UU8OjWT3zRSiFJwUs6tq1wSvthZveg9rirX4HQgsk/Gxf/C0FmuDjFfQmA
J7DCx3Ij408MOtVMiioz39UDooajiAqJx9irjH5BTERtVro4O89FeJxat8Of7Fgg
vw+vO4kIvce2ceBS0IElDMbhOGc+bk7SoXmvKeJUER9vW0xFmcEWU1wp9riSFks8
5RSA6OMH8hR7VxoElOSg4glAlecGEcfpbqkJ04XwMk4QWoW9XBRrKDAasAg3VmOe
e30kvrNNqHqFiuP3/Qou1H1NT+HET93BONl7povkpwzjqIoZf8F5asKu/cU+LZJE
1gvy4eTKhtW4s6n8POOsSArlvo/kA9xTbbp+QqSlJKuYEZDwiPDQ9ro6DaKY+fLo
dFE4YE6xAVxM2LHgDhR5HVeq8UNCai47cnjWEz0e0VDLhDLEoCOsBxY7tq/Mjkjf
qXNFvQuu34IrFAfONRbEUX6VExM3ThyQkpaU9LtXVmupYC9B0J7ChbTb1/gsW9or
4c0G0+nIKUC1O7ofB50YjSsX0oq7oB7mQpqXYexUmZSZ3RMedRl9XwvbD/xc2HVc
4O77TTRKj/BO/Jan3EJSw4+FNdZ3RYbD4U6BmFhobbyDNuMqBuYvQ/cW9TXfGCLZ
HoE+dNEKCY8LbePA7aTUjtDW8BpGNwenGfNg1FFi6rFyj2W75V4K4c+XpmnWOcbS
lHE/ENb8O2b1g6VrZ/h2jmawSEZFSZ6cQq9m/2WabC5d4LLIieSYPh+9jvGPmJqC
damq5SvnkiPyuI7wM8mEM4gJ/adRPZ1vjDsTJR8qLcXVgluFKrS8QLAdRuIyX8Q1
k8bFVWP8fHgxQw4rvGCs3/u7yNa1czIZFb5CpIcJIWYGt4IUp5tzCSDgcB9kyLKX
dILh4X30QuyPl2mgS6v/ZM3FDSaj5lKiH9IJPn1Nk9jRbRaAGq7++7UY7FUX3xWd
YV5GhM5wWI36VljaTJwliNLQTUw/VIUxluhDaAv682GNV6AWBbGhcDudaQFcp5IJ
RxKtkabJF7IAzQgNc2GbPrGbYBNvmqstgggdSDkbBUQsPqBKj1i6ZJKQ5l4IGW2g
FaRa4nYJIwBS5+m0s0J0HSufyBP4Vm/5obk65O1UdpmT7vOlSxWT7kemQNGDCoQD
PPrxSDSVH68q/d9A8zuWuitRBWvzDrs9BrQkJQp/vsFPWqYyqmth5Hfo/pEdRaIb
YmL/w6uavwa+/4r2LdGraCWbHpGf+OyIvht1jR/sYFjIrisfQxsNatD40WSkUfKq
vsKQteOzyDrWdqoWBDUTsoVo44twHonfIYVxwtsKzpbCB+usew9EDy/rG4bu/jyM
9DKO9asu/FOZo6ZhH7+x00Vwf3TtJrzoXFmxe5W5cmlNpi1VK1hLQL6JTbHmAsYs
ZafvsnmB2ts5WwbFzsZ7rPfIIY8Snhv3Ll65rS1nNdNMUxHCAjGc+cVsnBmEFhJb
zzcjBd+DkhiD4JduTn/TNZdExmv0KA1MWORqoNMfABZMVXgGG6t07n48YP+ayYb4
NAjna/sNKu5IXyrVGJfGw/Bu3KxG3iFi2OfhaBmA9beKoOKqC+bF6Cd0E4KZMYtJ
EIXwkKz5UexMrqjWyFbDnYggPBNbVrZL9ZNL9FkHzkvmJDeXd6u7th8hH/nVGCbf
Z6G6yzOp7OUx5B9EO22moZpm0Xf96+uTAe/znIaUJ8R0NuvsBJL4IQjLTvDipzFy
TympwAj9xl+XTayzTW3VvGi4fY45hCbigxjr4LMuvNd9e3pORm1KKGoxN0pNlkdv
fdKzRMoKZtJ9C840peh5FGMY8BrhNW3f5OLMSsAQuHvvwscBNxoT4yl3nupeb47Y
Vbi2zxBz3w6XkMe94AMs/sB2qFcTqNXwVyROzjyRfOqJCEvWGiMjkkv6WdVelrIj
ut77rCRfEpvZKDzKwNfJ5e5ulYFRcz1VB/Xms29o9AC9QsmMSLHGbNFaRl5EBRBH
f1dQ913V8VQM0JX6qB6FP79z7BL6RnSwRatHnlMmgSZNXsHNJpZMqE58oDgE2yBB
5708wQxl6prgyWI8+c2xIsMHHX4Eaq+1fV517Tevnchl2MgAPTeUlQsrA22lgP7C
1NMO4lESOrg/Odl5F4b4hnubrFoNj0+I0RcrxWriSo6AYrDBPyEtkanAi9BIpaaC
YgmttGPG/WfP5++BPfo4aUZCRDuUFafJqYLcr6WECfQhEEEqRGBjM0CmRMsEoG3G
0jA57yCo+k5MpccEho/Hn7gLK8pI39/LZAMUDmBRooVhI0qWqHuo2iUGcRiBJd7t
3X7RbQWcN+nbzHX5Nfz4i7ZDFPwaLOpAXGNVCUexxn08qorS20585+WfIqwtxGEt
PD4EIKpWXnGcA0lNe1Hs5h/vHNEq3EIOrUPHKXTpQtBS63Mch1yt98MaHKkhk6EF
N5ffjpdkRCiUed2eE7n5LskEq941oijpA1leOrB+yrYlXgsFzoPpa8VwM72s5HVZ
cr0pU7hQd0FfqQEgqTBbKa5lJp1d6+e5B8Mh8X4E50SC+MVqPc95qp//LkqsCqyF
YQ2Lcrtjbf187j9CYh5cLcxQEtkaPjhn0NVavW40PyXKeHLQTZt21eXVNoQJRQxx
snoXkD9k2uDEG1TbmlW71+77RG000aI+O0bnFpFeeln0Ox/GmItpJ34Oph/8TFAf
l0MgAat7/jch+EeSu6+QGtQLF3TtPMkVqoRIMXNYG1PTMc+jnEH5IlfDJHiyaCMD
ABSsZn5OvT/BCMY/eRCj6pYHVKDVNcDrlhEo0O9XfzI+oowmD+BWOCUZ7dNBPju6
lauP2rRBjeCfuYZrxBEXTI1THC4n5QfoaFDOKea1iBuAJ2g2XeexLnSRfERmTlNF
q4/5OQNDbWAdEONvwjQ2VzjIngQFC6jQSO8T6nb0SSoh8kc8Hur0/zXLU+Mz8HmR
8vF6Y+ZQVmO45dSvyKlapiYUu9HTC1altmKYZToRapbrvwmfWnDOr0vBjGmaAL9b
FA0pPmzy6JAw2dq4UPn0IZRt1Qm8ZQ24xDCQsz2nGuEiTQ2QYf48aAUDzUoRagf3
pIiIVi2SvXDhlE64fvmQhNQJrD0E8SIPQIVBpHs4Xw/IakDGKYBeqlLK1u3e8+Nl
ccnd8yyvjFlnTLNGHkudWsO6jf2aXPFrtZJXy9D+u378EoFyqnVcpuOGqiOP1X0M
nbn9I1pE5HkY1F+hYd6SUhSnz81T/lNy1yzsmZxfLx0Ezf2shktm4NuYUMgam/NQ
DOA3tpWOVAO5bsOlYqNE+/BjAyYrYxeRII353iaCIMW0IO5eHG4uKdeSeToYVgoO
FmjCy0FAMM69GJMQff1u9kkVAiR9lq/L67qO35/zu08kAe0PO01gBJYWvdJnCpNG
yw3tJtWLSOE/RikifXDy2z38NylM4Bhzt+vuPszOtUkZXrdnjJCldGso8YEfjZtP
urrz+c4XXpNmJUuCoCILM6lwbNfUG5igecN0Cza2gw00ZmsyA2fIHnQL/KmyU6/z
jXP3BY8+fUMeU5BEzj3AwULJr3GTGCPqUz9Lq56m/R/k4opaBn3ee/lGJqQ8za4k
CU37G3C0c6Vc+ps2T7WB0NBcUfoKG0ubKkvQn7hebqEtt9J6EHX7M+FEdBpKdzHe
FDCR3TH4O1AzsVYnqTwsCyjYfZt/DZrgsGsObX8oboXP4XvU6jHeNolOSHzgR8iq
ccape0bAZKGgGBIXQodsqvnzzGqTPDMdQJk34QXSJS2FpHG4OIxs/7iWaHNngiv0
A36gx7G/jqKgmjLEOsdaZBtHTsuV3Esbmdh2bgy2KgX04Q5cD96xpDCPDhctR92U
1IlGalisd/XJolEN4lmK27HZI15IEOd55vQ9AOucrY1IPi7dWD/hdOEt9e8dlS2Y
uRt/CrYU3y84da0zS/2QlG3Ux7ae6uvW5UkHnWgXpY1oxwPAkNJsBl6EmzMwAqNr
wZdilGiB/xv9b7493egcKhlzpxcqg9HfHqvJuhnqRMajodItO8LUa93Rw5DZh9qo
HptKFEgZueThWGG/XyM++1Qby6qdetWxFH7EjG0ObPeXYpQ7ItUBMr6Kh6PD49KD
jIwj94HvXNh+B/2LxrLpj4mUpo1v/R0gg3M9K/ozLxqYJ6Yh8kMZqzU4xnOygdpi
y6W2iSNit5rme/3ZucDcGk7r4T44d6cijLYqov2l+lbCWZJDIYFxIw+FdC5duEUa
d/zt4dBXSKMsiEahqKqlVEpu76ACGtlBrFR0flt31AE1uKAR7+66A3BVhNCtW9aN
G0QsX0Z9Ifar1EN3oY71WiPXGNrI4tUZcEtJ11SBUvvJbFPaxwC9Fc4LYb8vMO9t
gz5M7BGlrHLGLmBJBhZcnMH4uO5bLhvaljiom2iMgNXDJ0X5tl7Yv26D8EnxGVYr
ZxftAuS91px/JV/g5Ebt6+o8I3NYnA8zt3De+FnDzSOzaQvaClZoXyxrlxc6ToJy
yltv6BlyhsD8uMnR1/Sy848K/KJ6xea0PiNEwl+EpAe9ZV+70/sdziHhO2R77VWO
ufUtmmBKnT5zWk195GvixeLLxTLTDQGbWaA2A3FescIaRsXvojBQ4k2OQYbaL2No
thReLq5GaDaA73s0UIIA4n4lkaBqnXXB7wgMMc3BvO8Gm8L00QeecqDEgrMIkDhl
k5jQyHvOAXzbWr9F3ptNVaq1CP7sJtwfU7EoJq9S7QNeDzonWRwPZWzfztkGZIK/
hYv69224ENXSwNWIHH5peKsohyV2qb2/RLcq/0h20rFBY5UmFYEaTfxS2R6KXw4K
nB7wDlzWJ5a9YUEVIO9pKElItFtkCKj+7HLaRUA2LRINTJxlBAn/VlAEoqw+ZLK3
CuHysTv8t3NwgoQzLxSOrFFW22ywNl/+r488ly6IN1hQCZOG8YQdQ2cnA5l+ynDn
ZCzYq3iCLeS5MGp2Mn76RVEp1GKA0EiztQ9bhEaFXJx8Qf1cBQrz90hQNBS+b36/
3NVodj4wFedBElEKpuEUny68rGlplidLAWwyPz8apzMd9Doy3RC32mnFsQ7ceEIT
qUz9tTVRSNDmcZ2bfkishIlUPYoyN41xGFtFV1NTvBPBp4VLeamaiD1g+8XO5hDp
89smdRnC/270/g4JsBvTt2nqC4mxfKzWWlPKPDiFPN3c0rR/XqnJUQ234XNNC0DM
cEjOPi59s02tKI1w+ZPW+ENJvpYpaFqBeJGIV+xjoZgIr7L6lID8pYT5icnRiQT9
uAKZf60HJiRXpixyRroIS+QOQ65NCeCElHVCm2NuiAQvb71f71adh+YxC1h3eHh0
0mvdbYeD8ifONZrYw4mrI7Qpqqw5IgHDMI010n0KikalDfq9wqYDjSVukOGnrVJX
QrxdsDhT0d/4Hl9hzVR2YBLQzxtic4SX4i4PvHCV7quUSunYNcwUoc8EdUYOeqhA
5KrSRvjq2v3AdqEVxFmIKutX0mmcxwBlLhaDXaW2epuyBKvMLN0pr0nk1BzOgpCW
GYY1GQ8AHcHaT8LBVV891iOZ9HmPInj9Ykd1C10B+hAeevcYUb7NZyCi68q+Tec8
H3tsI+0H6ySbkcjbCp3v3nmCn1V8ihfd8kD60cAr/1xwQXehzN727WUih9qnIIVH
3rxLmRCfsDNPC3AKjmRRHgFV72odlb2siWbg8agRKWZfMIahf45zlGPjhOx1dapy
FAXR6BSOahBwthtC9Kgdb+dj+V3LBfFC/YPHvs5/kShOGxtto4p3hhXFCyhiDwsI
MbHq0UfGMwcGsYBRZl2a/ElKpzln8TcqDCP93PMk9UuhZ42MYccd2un/MAtVr7qy
rPOhrZlBMtWMBRkjB2pPVcKoB81uJtU6bV7GnQ1GltUOHOFFlnn2mRfDTt6Cyalt
0tOewEY0s1aTh7d77Jj6xEl5xMn00f3tq7OXL9xZQqJc7i3X/CFDO1GbG/TFamYq
vbHp7JmyHPwO+/G0DxDPzIXUyp5zgqLoXsxNS3dUhVUD/jh2j77YEMuyUI34gkF4
VjaFLD4n6mi6Sbw0vm7t61Patj9Dwfnd9AgSgEbRy10/TXIM/ry53kqTAbNYCJHT
6HcsnDbOdsu0AXUqABt8nQzn/rfplvKcXBq5bjhcGjLJEDmVJoxBc0nUh5YqlXAu
2sE4o8/3NNaqyxfHB8tvH4QUBDPLhXOI4uCFLSHGLrYCxB2a9Rf+2GWWuIXPIYdj
D7nPtnhmwsD0+tiTOyaTMtJUSZuYEQHdik9EQbTSPEd3PhB0idI25ihKDsxHGWcM
e7SCtxvdcBtwR67JjuKYBSj2IJPVCx88gai0SXdRAx0gYp50Z5sWtgSIgqz8ocha
Hdp4lhZU5RCjrwsZZ1k2BjvgBgwo4ag2z4SuRD5oOSBA3imwnXf5xO8XPtwOGhlo
wRDVCRo61evV5WnAnGK3TARb8zIupUYWKOmPlml2i45OJbvq+a97dYwZVgw29p21
G5u4UNJkU9IwK/QTmlxB1BnqwuFVCLdPyksF+ysKzd78U8OlTDQX9AnywK2s4wZK
xPXeh/zsJjNQit+bKclP6L0MsAuKT7uX90JnFmeSAln+1kH7pdNs/GwT9xYg+JaU
OemeBOSKCWkFjG9ZellfSsC7S6cxDUr/tqKWnUAKx75tYqQwvSiVPRE4pziPGU4a
B9gtuHAd/qLjkqWYMhraKgv0lYAnlPHLEKWAjWPSmS83At9H5YoxXAjKyWf2xI4k
40kW20FhpL+1zqgUB4yWUT8KPtyu8W6MbrpGWL/Rb4cbLtiM/BfKp2ZdbrMwokHy
sbYvynlGM5jsYBSRr8aHHqwzjtYFaCHD/d7HxjIxtc1/bbVxI8JaMb3ZFKFVssrL
v+UjsjfM5bS/ZzF0LcQ6JreEdx6p8um/kd1qTxn6UnbcgHZoQtkJEZihZ4+pqaqq
c5zI3CbKlfAB26Og+NqK4MeX3gOwiMCuFwjMLkjgm/a7HgE5c9xFxO2kcBnR6TKk
P6gLH/ztK7qoOmTb/yUfXUJFQk9K+l+RCSvLFWW6zEdLM3SyAGhCmk8i9XsBkjBJ
eNEVlMGxvLlgN0fLlc3y5AwnVKYCfosxZvNYPE3TYeB85E7S7B6xbe8M0ABTjG1L
ljlXBpOVrGPJPDd3inTRo9RKoyrkqVL6GyoRC9xZVBJra1R9FZh7jMEuS2BF0Kmi
VHW0Ner/lp36jgoeRUkrUSbl2UoL2xIEmeRjCPNotu2BBAlpnxCt5bU0NCueEVyB
zJb9JiIddwwnqC9hR6SQq0lbpKCSPZXKLsZFZzKj6qqFjfeqhK/NGUssSN43mQmn
6njQX1x5kW5xop2q9dyXEwkGn4vEqeOIDWCF1yDpsiglf1iu45EwJ/5OxuRBW4Hr
+mZo1xG3LnuEhQmllh81fFvVELqNuHAQz5JhN5s9bUb4XSQrSSCM3G0kV6Si458d
/EDFUuw741m8go+ueosIz8Q5aFw99b1nEaYvOIGdoZliH0kv5TciX7t6pe7VKh6L
dfWJH8oCmJ8iCgK24vxCFrCnhouqIlQTtrcDnhGqJ71gt7Vqh6V1YpkECc5hQpiD
c0rb1D4ZkJyjKQ5u6f4x1NcNzqvjzfCEASU2cX8bIGD1kV4r6jTtq0yMQL3kqFG+
KCdevP2kK+Mr2+0Mla6RWddt9eijL8Eh9HKGwb7zMWOvfQc8B/jzejbJae/yOoX3
SAyGMbVQ+6cwj2yJ1jleUIpmLk1MOUmfjUYbmVVMkiSjb2igTmWpU0nuKF96Ayad
yiVc7f9at7bqEqPVDjWaL7Sp7E+IeUqpHznv73iAv1T07mFexUM8EWawcERWsnTh
PQGDiHCvAPDDSP5xrMijTwJQe6d/QVRHVLbQA4LIk3r80uhThP1WWmidQKFD7MrQ
M6BtcXK5rqXm9kfRgNnK+VxyAnbl7tX7wEoDJfOifygXpXEczWEhmbuPG0p+pn3F
OVS5skwo6aS6nCXFrljCbVxhte2Q222/ROqgiYzugtH33EBKa84GbQj7el0zeBEM
XR1C/W1qpZuivYb2VCmtHrwVZqLt/G012RW9lH/aviqsD3vDa9QsWfflamP7l0XB
S5y5Fq7Fu4YRvg9oVv2tjb/BhVLCCb4aMmGVitO6XjHYjd8VZJ/mvLG1ac7As6pJ
Q7lnyytuPqPaM2ysDfHpcmA53vEJ0/poNrcq6oHepAOb1JhZ0C+5IIv+OnvE0oeh
x8365jKlOfn7XJGJ7wK5qjEfV/WIOyR+0swsAIsCvYsG1CaNmUYq3Nql/rOn9mkZ
63pJjd0TV1ZC0ou8sLZOG1hd2kz2KNdR5yeCabAAAPfWVohh7gYBcwvdTjU/Sb5g
a++YTev0Ia1pUUfttfoaugoe5Qw1xDjFImN1PerdOYJ4KmX7fyjpJAcOg3DsJ4Oe
5JHoub8yPScTCDnWX27QJFSC+RN0htaTRl1t01E/w75iA1KDEPLWwQSB3eyAebAe
OoTVyaBByYTuiAs8z3/tLeNVdr9RoxubEWoxBA1nNVUDzPZ0ipkIcQBe9yz9RMSF
7g9fnNkhc0J9wNMIjOaTMDxyw+8Cx4eWCc75qM2rG2Ct0MF/lZQ2ZgQTckk0mjZ4
Y/TpAUUx0aCYrrFWUfp8JuBbY6MtaoWRetCD3PzaxHIECKxC0fWLwZlsGdcbkOAF
v66fyZ9rCa1/X5jDBL0wLkLbh2sRNj14pTH6dCrifEpYXxsnkCEoiZb2cIxp6vSc
s2tZqqNGduUTc8btxjJhqra9GwUbmUefMlnCCkoV/X4YY2XW3LbDUMCNEpXygqJ9
WpxRUurlk+5wTL3ojhoslVVvHjJscfXgmrmxrkQ53aw1Fs1/mqWGUlLEppp1FzZU
OZqTn3HtCRR4BQ35u9sUzKFfsJm58I6mtwmHAnY1zkzH/Uc97fOl0pv15VwokU7X
ojL17JDEC+xjaUXe6AFZK7RNUoUZwnZvllA71JNVWr3mXI28qetmPBW3XMDREckB
mDGbEzX6MLen8SZtstTTEO8aOuj4PoB17EDyBd7X0PvU4YNU+6b7OB0EUMbSZjHB
neF+XYn6uBmMSu0wIClHVwzI/2kbjKoAV+fXSnUn3TKB9sjMd/UfHrR0m8tpbnyV
gbWFUo506Kxw3H/xojYmWmJ9HeTcuQe5RyEOj81nLCFHCILct7pDyy/goMsQQnch
E6ULNLecYYJnL+OZlmXTDUow/z4JQFVLaVc4jLnJZCSBEAsIroT9wmaz0gvX1jQ6
jAyzqXgZtnxMAoDIix4emY3WwE2YUcGsQvfSmNHgbhdU1BX6xKYHWkU14FiMMl4K
8yA9hgGEWpknoTiT2Dl/YXLpIehiBjErKpXNzevUQPRiLGxknjur2bmgTn2F8/qm
/fF+/EV2UKDU76sb1XmwEseGDcOQ5TmlCcvBcp7+IEpDLA6yqLZh5UoizV2vOJVd
ZzcUtu6KaSmB73oekisu2c1s24Aiz12BC8Eu+pL4z+yfhEyPERGIe8Zm+vX5Akuc
aDDbI25e92oiL0WFF4vhKj2XokdUYb8f7AZ+Oa3IhWt49oeua5avSDgc98EA6FWk
LfXdopk0rVeQ8Eu/flDRE+CAQddKlos7FvmY4uVqd+rlEQLxRB0SLNNRyJ/ahjLY
VB5jOKfXxZfnPYwNQnYtFjTtnEpMuo1ghVmzlT92jZMWjl2CMQCEuuS3elMTwzp2
sT/OwA//1cfyR6cxt84d0RikXzsHx8IBY2WWFFbK6nUbJRqvdltszyW5RY7nO/N4
xCZoZftWyxrykfAizvHJodoeqvEOTPKlqqNpBkYcqfJyKY4IRwvlh6/Dj4II8nOy
9Zb77o0utCxh4424IbmLNhx4qRsnv/pBBrviOj/gNm2xsad9DATXeF94r7bhmIE3
/q9WOgl3/wdTTTdTDY464MmwbHkP9U0/xfq3kqCEPsJI12hZp0X0asxgP8GeSOfV
XPwqbh3piczJb5F/S9/QTC+/B5N0KoF5+td+Af5lUOpVsEPnd9hvRFa6RXrgQ4d4
JDNviS5tTh77OmK7q7EEMGZeV7wiTALl0k99uKFCmYW/5VEMPhT9ChuKF+5FsSlN
tKybAp0PVnT50BiczaJxgSx9Zb6f/7cRUIEVXTVoFHxoHsgL02N3Epn2qTZRY8tZ
Q0slwhPKeXvrD85gtN+rA7bi0tcMbJm1QDEAYyNAgWw5SDG32WaUkmkBXOxq77Nq
UD7WEDM19k8FyRnnIDCKbP8doQ2YzP/BkBu3ga9lZjEzwzYAyNpFTldXyeXnNKgD
LwYuRZa2VGJPjrPG7RkpUHMXTl0b5jgaAirBRFiV4sUn2sDydeUZTJpzjVqyqWtD
nsnu+aUGCc8WShyFkm7VwjlGdwgAPrfSe3a6mRenXs6VTfbuQ+CtPreJiflvK0l7
UU3l4qQhKVnM7dk0AgRIPqNC0mlKG6jOT1e72IGEhD9SajS2iZgOWGfK9Q2AhQuD
6jKhprJddwTTRgu3yKJ8PJ9/BrmT3ioqV5dV3QZHtvWyNNlEMPzEENAsFl/FL/Ib
CfarxvtD1X0AZGOKIyy4JKKEomBsWpkv9miOWN2/lqg4uvX7tQDWXZfJvvnUu4LZ
oA0uR9p1ILXl63flwRwMxeDwYNmlwZ7j9vUQzm9SVWVApO1tmR4AGqusbsw6zk70
062Z8ot9sFiZV1Omi5k7y8tiztcNbRcc5ZnZRk45NVFPb+QIfJWXHfMmm7F+C+Y6
kH8O+MlKCX3gK7cRTm06AYMCj58FcDIabI6B1A1xzIutXyV66jwvWb82AiKSE2nC
6+Ma8SOUmIajvRwBkMBR43vBcpgwoyqMVDDLuObkg0r1Ouz2YMK3xmKlkL8NvGXx
ucuZSkw0OAiRBP8Y02OQFnrxg0c3xh8Wb8z39h4efaQnTaFcAhuzG9xtOTxxfp2d
BaUoeemgZ9Vcj4aX16iNIdygsDl1ao+9mqjfaoTq3XSokPNXqFQjdmY6d1HZJ83p
JAcbDreZOcKTyoYvwLYnPtON+HeSRnUUUkiJdSuJh8A5tnztZdinfnq2ZOolvNCc
aQRMXN9xITQ4Wx6Yte5KE7HXqDe/pTb6CNHkXIwh065et3/51CeiP3K9XpTRpCeM
FRj47kN2mrGQ6+5p3LKEIMLTRQGeT8IjNou8ZDy8M0w9prkf4/eFLHqo2EaOkKmY
3l+ylarJsin9WvaW3G0/lguQBQ6KGSQWhtrenKtf8FWjkjD+HofoKHG7UaWaDRpc
MTgHUkzCJ43MJd3l9VqK1GUCA/JxqRwNXzpn98P10aZv9g0T/q/7Ll1g4eqJdAfF
D7vNuXNjpK2DT7AwUVvSjRFiXfuGeffSJT9rL6mXsfdoCIVaSdt1O5/VIWGDgu+E
JonodcbQJUG6xzSXtc4o2g/VxyQXiCTWU6FmNjdyD/iMiHpGD09k+065ZTY6iw4t
gewfWzJA5KJQGvg2qPBADnumoRBmp35UZPOHeNDQLOecBmVwEkhG/dtSb6DJu8NX
sF8yNR7BwU+dS+lohRdmK/3fHSAuIeZ8EHRZlwMOplkHpx6eM6WbB2/paP6eMamA
Xs9fxhjulNk2YOhInBItYPk2QnEoAPbVUBtFvHi1MjX0RYOiDuFtYfCvuGZMXfRx
Y5Yu7907iI6g31IZchO5tCvz7T8wM9rdAUZ9+BMmfi1TMWpZb7UvdlO40fuX7vxf
Yfk2xkb1GwK6mymeW4Kdp/9zabJrdFGtN9oEkiEZKW4nJxsjlVoU/3wWlJ3wjnqq
6en5b7U9XWtUEGqhS2i5NwtWYmVAHPZjRFouBVJTbXW4O84a0QQXyvR+5aj22s6m
DkhC4Iw6TzRB+yZK0Za0ph6KxYSe0VSKAyDx+BrtZ09sqe23zFjJuqjfUiDpYj7M
l6z2xK1gX9X86WRqXUC8kyPJTA7I9u0vIRT+boe4vqNH76BKJXHmy8RAkS/HQBtW
io01mK5/qjdEaj+KjK+lhlLlIfvNhXMtu/nddNh5v64kVVTaESfu94KJMRSecrMv
B984ZObIYxP+PYGCNmb9mPw6ZMnXeGPlV2/NUF3CBDvFVBPhLEvCHN5ZBcr1uyI5
7zVrprAZ1kqtsyXACp5wfXVFqe8pafmhpE4boDtljhaMfnRrCmaw/yYBhVbypry5
M9XRNVRaSZzVZfKNjU4n98HxePb7tvmqzz2E1V8Rj+zG7HxkJtd2tA+GiS1mFP0i
KFLXwNEVfFs5FxEAaumkLridjgeSCw9cqsAzDoMvT/7kDAKt2O9NLnrkCFVxp+hw
Ocze3NovnrDwmRHBpt6LBE2E3OjpvSalcUuHzFgciB7GPazeGTUDeWSdU6B2nz6O
VbqTliIEwY/oftbWgYN/6PRZw/4/FKsz+KvzSGjhd7iyHNkFp67U41l0WT8X1kwk
a+/mBEwuQEVQvFbFLoPJvFMajhdDbGgbqUpdHtKeuYuLlz7jt+N5wiSqFrQD8upB
pztJe/YbBs1pzWSNOp/E92OVm7BmCdCI6KaNaSDL7XDk8hngt4flvDeKX4cpQ3SS
VZp7/YPEd8e2k9igxAGTh5fRCc9Is/Ivd461+FhWGaxp4qrF0ObJkt++29Fb06yD
u/LBUgMUG/SbWuzhdVaWWJKbiW2TA3sjicUUWBVp39pgQ0JxDl6pKwjNU8mevcPL
1s4Ego4pL7gi88HWk4iITYU2syolfyHVz4yJjWGvBKCEWvtrNT3XhR+9X/qNw8sH
bm1qqIzqybKwpJsAItK6dgHNPMLeMsbu8e09BvsLb4gF+MaVF1LoctThqR5AysUJ
ddgkAj4aoKgyJVc3VHmh0kd6VDTdqvzkv+fvd+yV+HPrJrwq0Vy1Udl1BLsEEJ5e
qurOt2f0BXivMqAxo8R0y+lD28Yce6NEwk7kt+O0qkuAGg2/k5c3+EYjhY3t5/fZ
Itxfk1otHb50Um6MAhOEZwo54HFht/ZoM2SwOHoXmzT470MuKijCqxeAi2YGogpI
KJ7PiQSWGkd2NBRiePKrw7fD45pyCNU0ZlLwPoEyHM+2SQgT3spUcUq+fxEdr7z0
EQo74D0Lkuve3lnCS9kD/fiFNGG5rL1+buAVWXZ/McdyH9k5X97pSYDQwu85ZSyY
iJVUY7rOlZZGFNY438zFS8KoQgFWnd4G8MA+ano2JK+YOQg/eEWhVGn6fR2wZOyi
qtLA8HggeVXQLkZk0JK7fFolwyoYaC7fbl2ofWwKA6Zq8m4C2h0Y33Xa8C05XFrH
9wGAaZ9I/6ezaoShHVmGpxilfA0+CQxyJelNWPQmMGOCHWfovDoIzxVPnj1J9U8X
1skrOxvkD4mGqatEY+/0aZCPxVBy+2iQIIm1gAQQBQvH42CqUaRb4NUt4n2Yk7qH
y2oscVfc1SOBjWKgnLDXDnH4F5TkN3VCA1D/gG5O7bALfSeUiOn0OLJLvFrb5d7R
FgCkfRBnL5ebwTA8NdXUVTP50V3JY2k1GT04OVSJXMXfLuoNnk2eL875nAC6Via0
B7M+lDN1AQQH0hFqqKwLSTAgBGCD/clfMDb4JSG8kkVLLbVj5SQZ9Bnyoov0bPMn
+pSKPv+7FEgVepuPqBEtATEXmj5dOlAIOJ02ji/V6prBfrz6hA4TncQt24IPkzOf
B+93ItpkgCdl0/LkjDqaxyelwtS5U5VwZRmHvRsmF2JRY5gTi/761LJfjxTuWTeH
Fi17La9yWof1bjoVK5eKOTcCdQpKxN+epHDO+tyWMVlxaM8CNNSRqEf8qDv2WDuU
t9AeH6TNxgTYnC+C1nCIRN1JcwG2zMx/198jS0I2ogZyTkR0eVKduRSusjfSidbS
Dbrw2kRR5H578L03EpvTjUFZTeGxZLNNKuLWsBdEU0pqWSJHU2HcICZhmRFfYHbV
0wmgFvrws5UxU01F/xuQC9Tlapf9dfAnLDQU9SWFalDqk9I2StXSaYVM9CxbhCou
FWM+uEHcP6jTE9aSXu0nfYc9GrqSq7YkibRY5l4hreR2nxpPhl2vQn/UvqmJmeJF
a2h4UAmNYl7D8FeZsHJ/RBtD+090PKalZIH71GofXiJwOzkFMMzUXf4KPQ+IGRdO
bwXigK65gyZxIg/rY8Kkg1ocXLoh34ebJfxrNSvZdh8mXivPJ2raRL0TuVe3PT1i
NY1vC1rOo+NWRnnb6HMoVIp4Q0AlvW67k+sX0H2TNi/t8nmXAL5OB1JlQW2TPwt1
eV642tLj2Ez1F1xSOGsehF0AmqZ0ikfHcobKq8Hl6tjgfm7m6phgNHog+L1SHUms
xnd8nB5GvRhImCzjzdfGa9X2aiRkorhamYqgFslm/KL1MJB6nUEJ+7gfqGxByDHv
fLaBboev6pFBSdcjWmvweezUkTdGJXMCf2ZP65ASFkTGtO6KX6hKluv+Z48cOfGx
BA3zTbVMNnCqv7FFvYotDn6D9tVBMTUVyFwn8+FXlWs2RjP6IRAdyac0j4ndwPnv
x+umEDlR56tPwcC90BIV/iE2k8G4pcxrcaZxuBQnh3TgspdcBqbBIQ9W+LdD0Jyd
2tttigTjaaa6V57Gl13E9/wIw+WYfNdg5i1rbHmr3PuOfSwhIIvqyXR0otlwk4PT
TOVN6gn9MrWbia3eC0KZX7/QiY4Y6wIADgUN6eZgjo8ihQAgKHhtvyzON+VrJoUS
eV4xBTwBfx9TfULion061vUck1CZ9UorUv9KobL3mJN5gZjfGCmi6tPRY1PVcx5u
dmKvEJ7lv6aczr5W+GDCL6jM+RN6b0zahKG9CypLSgvrXH656MOU5rJL4HjEANy0
w5z0mVuEe5pkHl0auUif4irFFVeDDKRIvdmElTymSBPkg984VGPNSwvQq50vbHpG
Yp3v+X0q86A6c1teBdtM2jDq3MvUTgtmhVA+PjytLkBflCZ+Vx92CAEFgRS74E2J
dH2fQfaa5BUe2QkmYxXz/mhhBlZnqzMOojNqOofNJoijNT8CouDoFYA7mUMjXLHN
SXeTonvy75a7KX7GZZSjUYAom9lknQnvu1IibNoAQ85ae5j6gAtrgWJ1/0V+P7hf
Pr5H+fntNen3BW7PvEvo18etWnzXFzqyUnSSJPPj2vy7J2BLSwBcma/M69w3RFjF
dg17BajITw+auN/9EHNAK/z5joBMUpVpTxLeIJzS5IsVYC9TnyUCW/Yax1o5uTh6
oM2GxSaooojqJx37av9pLD40sYIfXsVmLHpa+4pf427Fp3XWaXd2RyyxgZcrz6Hv
KbK+aIAXdMoFf6XJGxBaKM7xgS7f44EAyREIK0qfbXt3aY5dyytc5MQZI7LSz/vc
Eo22BkW8prM3DN4G8SXVwOIy5kQoACXEXe5MLEsqdyIYwBCVW0ZxsaBmuDdrE95K
huA7ve/JPOkXbB3qq94nuOFd92nPMIR7WEFUQQ9Vu7jJfekt0wOFWubyjYt9aw/6
ch1B664lO6ksxZSl+e8p1Vliv87RV0S+QGGWqlqdKbFQ7YxL0o7t7fdl274W7uhR
vCjDxAUhkXRFekCkmnwfWK9NpRofH3K1DbOg/+vIWzFTdyEsXc0iUeEk6eGTn3cz
+XRjRRAOOCUqkuf6e8pGR7TCukdeDjQrYyfNgIJh2fJimPYGobxYQgZgPezZoZX/
Anb5ungo6IMfheW3eT9S5+Ji851qNEV1v0ao0PqRH23M57lLFYl35nhiDnM8HxlC
WRJZhA2siJda9gA8+YgCURWx37bdaJ/5NL0K/a0nFly9hZPY2KGoe12EwRlhQC2R
VUHRW9ZJBrgd0y9lfUmYjH3heU0DPdPeYtsaoLr2wzsHiAs4fMNcCe8jHKaZiVhX
WNK1GalWmFtatKUNHRXK4PtRIGVmp3QSr5TClJzjrJWDSnYgsBOl4P6EVPnXbfiN
eAxL6XVm+hfDd+dC6/ZOvjddLbkpgywG5KDKvLclIATjD3mpOe/SYjPpzO+2Au6B
pwcXPMcnNZ2rDNd/c0Mv2G2f7OwafyOro8UAatfJqMlj5FdRv94/zC307d+1WPLa
Qc4BmZex4dIzViUj6bTgUiRjLPjbT8Fz2fuNI9/DVRaujDEKGx+75U+hUlH0Oa/0
gGUBHdC6qNH/02s8HC0Gx7zvyosrnZK8ElbdH+5RJ0eWwx9jkTVqXB47HNLzzxuY
nb0Nq7yDuyhd1N9OmKpZGyJccav2SRj5o5S4XxPKnKUXbnvtaX8PWYc7ZyTyJ6lH
o6ZPp/SRAFUUdIL/FqfOQB/k0IAKtzZ/K9N6NGPFleMDkWQXoAFeyim6lH80arvf
vvXzGz+EauTOOUCwhDFlINL062u7MzzGuIZDHb+RbAr0VVZ0NsYuEOaidt2KzEBi
EBt7qJgxUaVlsZtCrcHYNl7upq1Id79dRET6+yM399/D30W4G2gc8RQoXeur+5iW
K2dubUsTlYM84C+xhvOBQquESCrOfUnW4VnLid42VEDiAGNDqQaPq+7I30vNxcrX
OHyS/ZRRtqG+vuJT0bD2v2jy8HTGnkhfeyXzp2hkH/fRh599n95nXDdL9f1P3CGd
mjg94d3bQPoPHo+s6weYLm3efdOtGwhxOaguHAabXKs9C5024Hggy2mFDd3i6zYX
9Abw1gpPNXd6+DXKV6pbqaxI0xpFcjVipxbTrMrFjDgYkKo7inShdG+AnQfZAArI
GwlecMFLXdotp51XDnf5OftLCNJ2ioKDnu1ZTHU2K9WsDvJOgPfThIy9ikkk1HnC
2Qz35NQMzu4sHWbZSYPyx3DdmuNynMLgSs9WqYavbWarU0xGtomTocrl/AGOa0l8
FqRm6QLGASs0M2aiT6VjVvlZiTFEorl1GrDjVoRisA0mBdMBlh4/k5rssqSq/OsZ
8JJhqb4OmaWIGW9aAQA6Q8vvUCu3DNoZJBLgEHLMk/koeFDk5eOm0ggLkPYpyIfy
u42meiTznaEIA87Jm+2AsL3nI26i0/U+ECdgc8bAyUhSyvDT5NklYWEoszGDX5A+
2VquIM6s0PpA9XnYOz9U2A6z0W5oPwPYW6MBQP4nHHYDUD2RHc1IPQSV7PvLLb/3
GHMDA3lbQenoI+/X4RaheMICmIeSrdHDNJCrg9WYyA78PS3/vIRJwZ1+UPig2arW
n9syIz6bZkG9UuouIUbeCVEIslKuUt0/Cgo04KdkqAS7XN5mYskMc8Oz7GVoFmu6
nwZRPSG5V5EJ2oVnRJ9zlRchSAnAlCiVKZMKc2ma2XnsSXUIMUt7iKoubSgghgO8
ZIVDif38tGnqHDfxCEl5PKJNShMoU1y72UR3YuqVX/wn/CN8omOg8KLa+pUMcW9F
3zj18DC1r6cFbRCXm0AYa489fd2QdhsJN8u3dnDi+bPt7jCGZgKigcgBm8yxeOMk
qBCaRCIQP+D+Eb7sPHNMXsaoW8RrBrfks2omA5X9Pxq/pnOGDJFEZ5FE9AVad2fr
Yl9tNIfmATC/lpTh9prBcRh/Wkj0C6gHtyeJjGPcEAWohN8LN4ypuDQHfaYuGm4V
PEg3WlLCJ8P5bVifcCepTJ6/2egOuYMT2PIgycRluowDXew2s8KcAzyWk6dgz2/y
Wvx+MREAgj2isc3xD66XoPqHAZ5euuUpVxYXW31wIAfYjvoHwaEWIoE9FfKYjgqH
9UlAarOBVQFPXU3Tzq/8PY/EYwW6VkQSsjL9dG+PKd+TSuiNzWC0IoGOdKZrRO/l
s7auUiWP7fMYCWcNefwi/qvneJJQkMqmkeKHIERHdaLTCAAt0eYZ1WjTgltPc4n2
v2uv3xYO8gcyNm9s32//uIKQppzuYcq2uU9YiYCh5lYZfFZeA7JBv39ng0SNgkgx
7tCABaljEsxGid6COdwtijEooiidtV6NjmQz/LDpHIdXewVdhWSUABhLlL4iJ5Zv
ZHtpnRBwAnyAcaEqhyBbN5kHF4LrdqytEvau8oFD55CVaSZdtzmxJkCVLBgzuFAF
Thg/l0y2RsxbYpEOXPjocHftZPuUMbk01dEidDVvoY6selWpm5hi+TR1MfnDVFnl
M6x9wXIwEJaRBszBEcO9jEZDzD3Dw2SdJxg570+bRzjtzv7171GS1cncCkrXLOSq
dplx+RswwTogPC0MET7EArIMbyZJX5rsnAG75esKxDIuvyX8C8adiGMMJ4stShU5
St2pf1+fqvySpqcpranMamI1385Z4HaxyY0sYV6bPDJT+iuCEoXi/g5vUq/VR6PN
/92HcVlhJqVBCBE+iy6D5fXxj59oO6lElrRwAsBxtfO4pDB0EtCrTZl6XwENex8H
gkBsziZ+Fc886iPcrxOQKLOQVFPTbq63aCpso51ctxQB8/PIM07sh10je3HgHcvF
sn2ruXlCYqCXpNpiRCH95VvpvKrYzPy9/zIi+KKmANSUygyVyCmhmC/6yYntWkYc
mZq+A6wiq+MmgYwdnwD8WEj6aPt7/KQck3zQVxuDH7oIhZkKOpbEJmhN71JU2lkq
TOggpAWwuk2pspPT+AitQU/M9zeTlPw5h+6w2KzRkQWyIDV1i3NSWtZU3tNsZLn5
jJqd9ja2926yq4l2ocAoLSR5JtqUeb2F2L53MZJe/LvoxPxGC1jI6lTnjbtq4A51
HXWin/9UA4cls+LWQ2/l+2V6A5E6jmHcRsXAQEeAjokDm/HBn+UDMvgpjYp+ZNEw
zDxr5XbFvmmiP5uNdzSQkLDpOqWF2eUmZVBpzBhvFQn9cNjR1uhWp21n1DwU9y0M
eKhmOjaP3Zm2fOZIOk5WD+sI5w5zAETJkjAU5q3KWU8DLsE0EgB/b4umfHIzh2rz
5IXjyJrPEyzmHunFOSL8tGQQyglp93vVSXc+WsUy2YChaMU100muL2l1Z0+csyTh
jh/IWepN5y4xKZ6Jg4JbyFCdY0QHN5wjfgatDl9RU2oWZBDD3ocO5AMAgbw/7jj1
zrTKEmZJxzV15dRhrFgzP51WZ5jKnU4yIaxVqYpAT+MKSJSje3bkVm/aRZAUSd55
AuRsFRajCAPyKGi+Mo/OFcrOZr4eQf49hC5hTV641JXGzo+7p6gRMdTQ50agwPeM
lXZVPnN5IVRGthV3MXQCRTvUedVPo1Si44VE+M/bcBxD+hTxncLF6yJcfYb8HU7O
YZtZ1qs+x8zpF688LLb/TJ8Mb8REsHkSh82rSIPc57S0lQjwyN1FFCZbyIMCmQS0
E6cmGJJqnyM9pUDOPFc7eIuOa8ueFzUVbAeuIhsIJO1MczvC/KRE+j5PxG2CejHk
CGKxVZ/AZo48FRVUyPNi87BQfSbDFoRtiTFEuVcZOnLuqxdNNnKPMYtuyGCmImls
MJ1c1/h60Fp4XmwQrx03Bb31hucgooIvEKWH5ZvsZd5a0oQ+epX5uX+bBYBC9tCF
QvUi9wyw7hGXwcETtDAyNLZGuGJkaH3hg4kwc34inInY3u0j+55PES9BZr/pHCty
71bGOPVvxxrub9UkAPV5I8ose6SQS5KDJ54v8xJoxvax4/5aOvwNrpjqqwN3BmDh
TXEm3wn//ryMCjpnsRU7ouUYAkUUPz6K+sm2am8qczjNn3FkFQzg+a7W6uy6hv1n
wVdvWE37/hxjMWXj0Ao26RtZ06pl0yqDWE46M7UOtGjMGpZMSat9RDa99WEvDWKj
dkitGxjPURCb1weh8c1xon5NUuGVzmilM/bTmJpbAZjOc/0wfs9epyZKofZggZrk
JQCSHqfOoxDSw8G5WMw9ftUbOeXyZE7+RljBk9Ojr33KBLgk9x/iUsjvOff/443I
apCBnD//LK/AJ7Ml28VLa1laUO3E8KJ+9PdnHfJirdfrOqpMlErFIFNuFB4lRklY
prnuNQC90Xnz33dnzcUQZKXBFK9YGozsAtN0ZZpT0YaeKO6/4rHYbRhahwdqBdfP
ftmM5WkyLy8dSaz2/hdHou227RTsQuZuvW4W1nedf+LIvXQrT/n8TQgW+d0p6hZu
rPe3Df+soMDS7bDXrpKH2NY/OqDrVL6sFO3eW64jl+F29RlpCCtm7N5op4uFSl4I
lzaPPfT+KXnT56ggZcy1lYSYO2UUI4dE0qo7DlmQ/DhVLgqpUIx5wgUww9PHeXxo
tzSgUNvCdKffYE+RgUWFOu8pqcOWtP6Tk+dKdxx0HZzw3U3cUTE8Ua4dzZXgtyd3
RagxhOzSP7cBFUZan/lqBi9MrKp4SWvYY1DJwDn95zsb1mOyuXtfu3RPcsEs5Xj1
HcoPoGzoXVvAbroa+PQ7ZibesoHQ6Hy6oI5iEFtA8XGSV/Uyh62Sr8qoVnQwTVds
IIWvOvT0cP+dQQ5vSiX3aTPlU7fyifGZjpGWNaT1e75nopnmk12Dxsea4cI3lbmG
0LmGiGR7OmSTTCIUDi+pmuJxUhqgGTfab5BLfmfap6VfNc2A2VZCAwH47t2743g8
cGzlMYC2zfiRFWnTSVwIoWLMN8RSfD1PNP4EorX58tGGbVVC3hpKCKh3R8ZtRs/D
NdjvuCMNElx+8nKv9u/7dtToUPwG6a9O92LeuJtqQ7IEMH50tlVK24kb1RX+a6SF
8vd1zVC7+n9hLlGR2ezpniyb2w0xbPPJwo+WxlW/QR+tsK7K0se+bjwC1P1QnRX7
5GF8Tg26Yv51wi+On691YzyTOiGaJyDFBkebnq3mrPTOVToNsjJDg/x2HWGg/wSm
iafzPyxPv+0ALoCqf3Igfv/uM1Td2IGaDvtHSgKTWJCEvVYrg+sjE0mak8MEv5f6
YoQb4k4aQ/0V7h3D7QURmFoheYZlVjLqgZEsoT+lU0d59VpQe6IQL9ntoEk8/Swv
U2T4ZGqGphi0k1JM55QFQDQZg5xHF4LjFLEQhHsV0O/hRl+O/ER8QEQ8NShLjxCT
KsOuRhFjRUdKDTrcbZJbvVeE9WYM5GfFiBU+xPQPpuKIYrdmdINsf4JvDSVsS7rr
P9KTuFvVYH0zIMFb6T7Cjx/Ea/HjDezCt2LYjgIvvH5BdyAA2MZk+ADPHS8Qlbsf
Aq3rmwhXbQ3ClfPnj+/595Lkq5o+9hh+tr3sbm+B196Xm6s2dNtUEZWhlDzAkdNe
g6rTq8U0rYVwzc2SHMI4xqCoQFOkEd8WjKX7s9xSQ5RWDqAdAjjfWWNh3jVkrhzs
qT0/v2zDkC7LJsCrIlvH5KlbI+zB6B9aIdfe8dHPlNNiY9hXh2pAlq0JLYz9lggH
0Ha5XDWEvbvAaZ2O3si+l56rDp6WzgO0JRpg1uEqnpvPX7zJzvSwCOS5N6aFMrNA
7PqfA53CYLCVNHhcSP5ANpbPoO7x4m8AsQilT4wVpJ9kUuMSMqmuzAp5yH/ILPuJ
Zpw31ChXh4Xpnlpzi/XMO7xk3UoRzMNiJHqYVyx7u2okUAZ292Y7WkBF/8wz2XqT
ZT3GIOA3pghbQeIjAOVDDGEkYy/PV6mSNW1tOXYZOnGGNVdBmbkh4tW+cmcGf6G7
fh8fhyKfEz3nxwLfIgq6t4KwA046e2eWzsYcDKqKPOgecpm0/8ZDu979hGvRYmpp
sEa36vRME24I0M40pGIcdppH/lVEGYmnyZE1kP2tZarhJoNdreKogXuxfbSZhnWe
WWbDfURCzwtY/EzsEU8EaN5HWpW/nwEoQn5KkoXDw6mzmByNPve+CukKogv3ViFc
lBFLLhTYfutsZGQopkmVZSQgI2o+Y/biXG7pYdn2atzAU0IFXZLjzXL7xHnEC3xh
XB122mMw+Q03GkDmPaXX9/7uSsSfdPVDPyQnlQbxCmaayF8F8U/FuBOHcC2sIDmZ
9MbntZYc6k0Oy/Ew0gmr8Chi+suxqV1caMsFskyvFDMAPlqSl6LVfHl1Sits41bv
uP/W/CyTesIYPFe9VTHbp7PphiX+1Hgigb7CpLzLXJRoR1mmAo25flmUu2jpBDmv
o/KYDMY6y+V3Nr4QfdAcrlkwp+eDDDK7ecC75oJEEVSgcNGHJ/ip7iPJYWLteDcr
+Z52rwcT1lQXJxSHPCUQj5YnJBdQ8ky6G+Lh+Pd5rcrEGUB40Axxk8faaSFOojrr
a0m5qVCYFmg8Zx2LCQ0hG7sEFExPyyfD6CtDiVtUVWtM8IOY//T7KNYIYR0bc07o
Gk7IFBsaCCTnAEPdlpTnkVsAANec3MzbSbLIxBF+5iQnI4TRaJvooVLeWQjB3OAZ
0ktIxSQdahhrmvCwdP65i2EJbl2tqzuROR/taBmMlmNmXMO8HOs/LYIVQrtNw6dv
Jt62P1uVtMA0QjuszzMzcsohlR6jDARjOWRUyCJVK+809w/vb4APMkhFF1lMYsTX
aONfJWzdpxPggWw3m05L6xnHdaxmbB3Y6mrFlkKisNsQ0MbOtgsIf+MRd7ryadvl
97kKLLkYnig8UuNqYJVNuwkRbFzEUYZFpPmKiNckkrzbbJfD5K/T7gTcot8tixHa
1CXX0rgadtFI74sgPwih1/ksKi/7ERr0gO8xtR9O9btw7tijvEzrvJQYdDPeOAuf
DaeBX51YgFx164i4VyHV/M5/sYehy01pUO+2SJXjt4hxKKIw/G68IiBBl43gWwmi
g0ueZO6/oLs0/eAcBREuFfwvkYuVltusp8QfDG4tRhivA7iOEqZlYjsh2XJEpB9a
MjGuUOJxD2OIlYjfHih6VJMXB/MD/bgmrNK4F4d3AQMMJpjDyI+iK7aU4WaXLG36
8gKl2k+bObi2wndsD+YkWu0uuQud6mz6BLhvbiuKx+be5xdhrJ6W07j0HZdeQyLh
xNJr6oT0JAmvyIFXM2aSiPff9UgROtAakDLgQSwFz1qDlqQ3lmvdUsLFVAuSkGUr
8Rb8IJdtg0FJXS19RszLo1j505U/RNpt2RDt+q3d5vPjezAch5Wu+PwVKUInqfoJ
8y1FPtjI6/ODnzWq0vnqmcHxpGbpIoHIp6xZ1OpF1t1nIzDwmaRjnKqKuOXa5VgN
tveWcKeMcayQFsk5uAkmE5MzsrtwYVpTbo/Dc8g8TvGgO2ENG/Z/kmxiBZQF3IEx
6e7deW3ZI0uqIMLUZ5xAI3F3h4NaPHZnV5RjrUNfwpk9Cfpx/q6Y+e1FB2Gw8GfN
hPgC6hhcC+pc3SAc0+7So/LGUKKAA9vdV7pB9T9SNrCkQ2ua15o2HECQ0H3Zk9+G
1ADdy08wx/Z45Udw4zmnU1ZquQu2wDU44Bemo5q4IruSue+77ogeCdm3LDrQ3Z+o
W5/aNCXENJ/+TgKWQPf5oKkvoAzOi1r+S9+V8dWg3MgFR91tRj9en8OHmmxr4TKD
YYUPLMlg4uCJ4Ch8WZg4YAj8ooVEmQwl2vi2RkqdWViBi/iGmi6P/c0eCU43EeOj
o+9rNgPQGpvcrY8c4BXzOvTXF8DE5VsW0jXaT9PbDepvA1YuawZfwYfboGLLPYcR
5/r/G/9S6MdDBthrmgtw7F8DzbOeSjM13DgyGgOlaCPl4EN1O97fkUtv8vsH3fux
yvw0O8ngMhwyQxrORszpMJg05mwQXZOTo2mgCElNVh2Anc1zoZ0Ht0ZLDf6ahF2i
7t9oxgrVjBWhM2czffYVuw0oAzoOLVGpEDBjDhh0J6SRwed0XMHIfloHeRu0gsms
BdjT2n+vcZgeLbHR8Af+bG2ZEIAzYWl1ijWz1WneVYBDDpTVonC5ExwGtNESzhKv
XhepveE7q+AZFORhr6xs3zuEz5RhZ/eXJt7zPLbTeszgplcDsMXvI6s9BtOHX0Dr
Sp4AkTSqiDzdnbd8wGzNmsNJPqL1yiCnr9Lb9N6oLedct+Rb3ZCZAN3WPg+ikmNL
PK9VCoB5xczz4xflb96XJK7Cis2YLKkHpEz15YXSEDdqpI9dtvnmkMnhLBN+W1wA
2p4ckfYQ05RFHUoOlTWopEVjHVcjCfzp58qVPXwCNo0TIR1O1+rMyO7pRPqgoqIa
bpLToKnxp+pHIxow2bJ/s5LVnfCbM5alFr5vBj9/3JfnBak34VDK6ZE+dDTuS31c
GhqH9S3JC7dYo8rGAcJWErhd1qfCH15UAUgcKYkiN8SOwP0ShcdngrD3T0yz4ZCK
aoLECT38IwuMB/10z9U1swtuarwmoRwaX1hCjVgvtN84Y8MTDF0wGh9X/PuIet+Z
jHQwRt98bgJ+GNCK7wm3rpnmcajuMFn4tMrbX4k6znP9vZOw/hXzEl1HWzz4xHhC
onQwFGvKg5FiaAhdL0nI3hJXHC5TL51EoCh6ADERx/tuf84MkBizxbdLrl8qGmQc
JovdaEDBvp5HkDFhUQkEqwFOyABzuBAdWdTquF5sGqadCG2x0I/Y55/6O6pGPvVh
Q6Qgqm/d797jWaVkYUJvH6U6JvSk5jM0WAlddRHml6SxF9IZZZhmXKbLgPT0PztU
wPI6RymJ6y8bDfX16vLJjEarrBjWdQgFxe3Yd1YeH6R1htDg9bTDOq41yJB7LMvx
4M6lN6lZcWURG9x01zynWs5oAThW4ztWUmNExAsVNBbcIfSpQ2Oua1DmozZkczO0
tYeFyGucd9Urc4mFcU/ff1bVJ+mgmb0ntR4N92poWpXLLJzFZuMNGDCoWLmjK/Cx
1UElBDn/SrXulYVltTMkm+AfqZq831aZl3LKwAvYSGZoQmjpO+LhFN7XRcoR1ODo
U/gzU1i8YJIosSZSHDIsHL267XwO6HqDi78gyOJlwDzCDaBCwbb3FkdG3l5vQQt4
Ar9qOh1Q11N255kqpAI1gsH1vXfMXZw6kScIdziZrcHOMLqzASRS13+3Wff3VYwU
fmn8eKtVKgyRcgNqgOd1EcDrwRNfP91/Zt5dTrOjAugDfhxzXupUproBf13Vtxz4
4a6WjQkwSxhm8pikpmrJuGE52mdSZjqG6gAT9BvrfwVz2cc9x4WPxyMDLLQwtGZS
nschP9NQ02NVkt7sLxtIqMwi+zo/1c9A7VjF+EpSv8WXY5a0ubjiJdP3hxf3wduo
RFvj4RmY/laEaLxIHXli6JGpJkqCJ0O5spd0y6g6LGoHJjuXtxR4ajwkrVg/mVDU
kVQBv1ARwrgJSVp01JSUc4LRFcJH8K9phKPm7EY37mCs84YLUh/ZbOb+W8UypNqx
e5UdkAPu8xyg/yXq7+XTrwqIgH0vxT0849wq3SSFb/wEntYQdVUmfxqZdhu0qOK2
MSVK2lBzu7OGVbeT+tr1YhFYWQSHm7tocwx/VmN3JMOcIeVSxA6QTJbq1Hi+n+lp
Xqt3bYiDxPoRg9xFGdJwTU16QpXHaNgcgoGjOiDnbPL0gl6ENUh/hL/89gletNKN
0eZDSHYwNBLp2nuGp7+e1zCiXzWkN3oxB5wrHxhVkyBl0otDprMqskKzoDxc2tjm
GppzewWTjJhxSivRPhhaxSRmiRp+78hjgUsodK+kcGuDH65RkFdDEFOAqXAn+gVg
G4U6zv5k7Ph1KZRdoLXLLp0wSy9VmrElIZ+fEJS0HgL8BE8XC4FvEgZBQdFIrXdG
CgGhecyh8okldGJEJUs2EcpTHmbMkjz0lAO/UnM9cd1NbBy4XT6aaTbiMjAdrdB4
nY5S6cs6+ZHmGotuJyPNoVtcnCsOs6C/SsY3Pc3Mve52SSk/vTVPMl59/8nyU60M
7sIKIdrvlZ+FDUyOewlJaEW9RwVr8aI9IY39TeKKUsOKK4pnLpnAiM2eqjLhutsi
lf/1r0fqku43MCIHGqW/yKnP0zh7XT6Owb6+WEBZKMQCxp2T2dTMUBCCsuk7B2O2
ktg/XyXtDSjUlBEVNo6yc4835EAXor7FhVUYcfhLWXU1AMxHkZYkLfHBxbyDFL15
ZXhElTGhNfb+cUlsCJnwCr1LH9rh8qfylGCWHgcqb0Bn77YiWHPrBxNGNWpJ6hov
Man0GVfv6MZqV0Z2Kvj3wXM1Q/S2HNmPcwbRrGWFzXSHz4tDFO8hLEKyoghQLyaA
8sYZh5AJKFoEeIgJl3gQAGz2gsQk0KUhyr+SQkP+TLnv8wycFP+7wgwVgLKsokkF
enTLvGKkTka84kmhcuFmunommkVxpMz0OYHfLbNcI00+jw7DcS8YGd50C9ynUDJP
mKKYAYUfkYxiRizfW8C1FSGcRLW7/eELxBOqXnsAaEV6bL7aPyJb7D67u5kp0og1
Nfy5qWIE4prf7JeOJgss2MyQl5CvJNNb6Ya+g1sR23B557fjb7eJSl4E2XPTTtQk
nRj0AWiTSmIVHV6rZCmVPU9aB0Ah1HEr5YakJAt5Dk2mGitS47fO5E07Zd5O6FNZ
y3+iDtPPX3bxlbk4MLpkNSXM8N6FSEUxMofZ+KwfltM2snM58Suh4WWHbeM9O5+l
57Ib2Wy/nSrQbY3ksrAeYZuvEiQZki3vSCLIhalrzywQtjoHtwHj3XgdZn5ljBAZ
6lDEMbEjOwTNhzbxq8+lXLB0n7e3Lab/BYPzaCBKV2eyD4v56n/06Z60A2bjFmH8
oFnxoOoBuehOc6E0VQV5lOJvVBhFlOf30Iw2BLi6v98f2++rq8BtJNBsFgvK/ogk
HPqYSNIWs2HNhI/As3rTOHpH0bpD+C0ikNVpNxCYrY/u/h58MiAuvQuID5AsQ/Q8
OfFAESDb284eLoqKawlh68KSuIfehvsRuUrLXmGKwSTwgUN6pWbmwUSyPq1zuz66
AinV7xBLKmbryAbUD5C4gHMwEsXopbXJQxpUulNjgHV9CqRWMmuiOJbw/nopj/qa
oVkMvvRMpD6l5cQQW3kie6/ROzN5vtt3xK+o7VcEMe6TKBm6nAuWPOEzaW2BSKb7
mGyOR8rEmyvdYk5q+AtGv/ou8ap3XHNztuncD9QGTG+k0eJWB67IkU43RexWSNtE
DNhCC0SRZl+62aszP7AJ2GF8qKobuMNrsvm8ooFLAsCjwTWl5d5hV/L76J1umhGS
bxYTayUKc1V4V37AZQzNLu44MYbzOCvVx3uqe5siTA4jLsKfLdE/uFMkstwUbX+F
+GbZXg+XFGhOPbaxBCUyFz4E+CRW+iiMbiLGxftGcm8PhwAHyN5eStoiqCl8Uvq9
Qglo99YBdDJwQGu/WOnZ0i11u3Th153knMcjwe/Akx9ycufKynJ//jpODLBDYnvT
L48o0cqiYvWhiHs67X2ZnwcXY8qCh8vtzvokNTXJEY79ciOnAE2HvXaxlzUV2pqb
UMR494l44cgzFmLdDDtu8dZ9qbliSUm32SMybfgUknizBlxDhG2C2LI8yeKqHg34
SlN8BI+KMNvoZVryvm/HMiRBs5rEBOPqwOCHsUIDdSwRYTnqk9lPn0dnHe8dLDeu
60nsDiW8Uap95ljaED455X2ze7Hx2wTl4SkmX+9OdOYnIk/XlIEFL8xW7dC06btI
Gdz+8WAv6IigcJMnBbVrPp05Szi8uSFP0LpFcQC5uCu84WiYSOw89C5fe2ZyjZrE
tActkPS5R+L+gt552hmZQNElR3lfgUjM5XCbykCrw0O/xDqKFFAtCQSSmXEK/8sq
FUggEw/ilfMS2W0dsMiou5vbw/SleuW4oeQPo/tCJKoPjUdoSb0yk35hMmTM5UeA
Jdpmm9smYVVtum3HLL7CH4zRanQklKLUDgm14yDgk71/JqIQ85zpYZuAJVVM7Eib
fTtmJSnYbPKTRyBstSm2DssWKJwuPuVU3dB2B1zlpiFZaJmbbfAY5mK/p4+BXQmc
RTrY8D0u1Nv8C2PyElXOW/qv8RDQsIuIl0qBHYUSKmUakq9E8OFsqL18jbytUgYu
eAinkJ9ehIPAOy4ymY16aQUQRP+fORdOxWn9rHjK2dyF0jT7anPMwZ2u4yExQuD4
sSVEMkThANG+uKbCOfCX/rc1uOcox8dWPCD62o13eKQ1Sjb5enNTUSREGn7m2P1o
WVYtZj5STzy/Q0kOJt3rrE4sVUB/XvDETh8Ewrfde+ekB5o2sRaI9negJDyy8jwo
0MxbcAqcAix09Xwlvcbf2u6XpMiiKLfwJ1jBLcxuJzn/w3dtAYtS44Q+BA7cVIEb
DFPDptmy43f3gmV+zGqlJwVoEry5GTqFSlOo5wPuZsNuBAINB5oBlCb2CuHoecNE
Zuo1zqBgAdKzJRGkjNJQQXCkOoubt2tXdg2Smj7YjDJHCBLIo+AlS5fcRjEvBdVm
ty5Byfutu8uI49XiBbqxkw3P6OP1BhJHKhsVdn4pnvCyFDXBcGIV5OL3msa+JAyb
TD7BT8j9U4r++5NcaoCZx9nz+C593w7pCrz2vgWhnmLY8lGarVUF8t2aiMq2vW9P
GIiJMytCGG9JDWKMCVpDGI/FfclAy9qHr+5d5IhrNHg4jpJ/KxDC6VDtersroJXQ
/nmQ2BAdxZaPSVD+V01DqcrDUyzKpVJK2u1nSGKwCh6PXy9PrPb4yUKKby9Jcweu
Tn/v5ey87vAXd/2ueoaXW126eAzv5YyTMOaWV2eChqNcd9aRbdAVIW9t6yh68a38
yYrizcezJfxhX832A8cigu0qNxoASSZghda6RP7J2jruUTkOHaBrcs9NMWICA5f1
JykjfqfbRCmRdu+FWAGVfxcR52A1MsBEATXUddiArzXfwJxZOu8Ka7kQf14FyUGc
0VORWWAu/OemkqHil7fYgfou/RLICvskv5mpSU2hgFZSPEwX739RZi0RL/aa+jmF
rXkfOy4K1eYq8E4ZZjhHMQpbql5EWHu4baV6SFF/sCYOWbFIg4FTIS56GxjcZhLo
9UXfSvHkk6vLYbKHLvA/ZoSgAm8pWwRGpwM3zr8E4BKLizavujIda4GDMJJJcNWc
1dYTbEj1sZI/Q9jIDFhVMt8LZvChbrRsNm8q/C0s3tousv9jf93OKt2eyvD7BSXX
fUYELZ7YGIYSrtvITFGnCq/Ju1Ec3i5jDzIGK0lLu7v1IYdueuzIN6vzXpYn91bB
l4fdlYOwYt6QMbBysi35pK+hdNdm036K17WrcSpd9fYgtafPctIG2fSZeMGlAKZj
GdLzWy7uCrjv4lz40f6DqwvIBg1orrmYpVtO5eS9rn+roeoGTx6XoSS0K0I3T0dF
JqnHi6EFq4Csx5ScCNSdebQdz+9OS4rWKe1Jx5lZpbYwoFfwWDbkMAKiPu8PLQro
0EcLnpfJlGxWHSs/I1XOAyRZ9Oteef4N58+ZZ1HSr6BkTEicV45Nzl3q8AfnRogP
6SBLKpsBsdmlwqHmAp9JI76B/JGoA8aEsWrPGIUBhYALNGIGh0qGFwzCUAI79WYq
PPjMR7wIhREF+gY2S6W+FVbNnbZnooPqZLAroYLuHOGu5jxKRCPtFtTw7/kDPc2K
Np//+4EJoO2C1A1AX4MMiTwdJt//NTF/vtxHjdx5i0OP0A8jVcTOmMo63teHtXFG
M0NSXLvpnHqI9nFzzJ2kgnc3v3JnJqTcl54ez9WUYapY7viIervoJMRrbTjR0ZEu
eaXcY6pEgY7nSxzDG34OIxEFda7rSsig3hrL+QExRP+g4UXPIa9lgXrkQVHofaGD
O6uTvMEGWmkxgXn5OFTx7mXdX3x3wCDaOf2Daq6MVon2D38SdUd2qpyHAeq3TCwe
cN0FZ8oezoK2MomN2Q+SoWIbkupDR7iWXaaeVUrWQwqfw2i6srUxWVpa0NRoqV77
bJHhqecD7j8sIPryyaxwRn7bLD7kfpFM+n9twSbof1qJKuPbdgg/46eVi9BWCbvT
yv/NKFvTFjNXlZDnDYTbyvS8BHgrLjkxMReZ57CRO1PpjuTT5qAM7WdVWauF+zoH
NFYaFTyq7a0A3DawsTszEy3o0WicxlNiFKMp3Vkr3zC1JdAZ1GsWXn4Wisjm/ncR
j2v3gVpdACI7vs/zq957oI0AfYfBx+iZGTx1orfxzcoKIKPolohS1e2Sq0ZmTCmH
T/tcJ32ZrUooafRS2v2DZiDzBuYGRIWzuQp8Rk+U0M22wyqmqMm/3rRp5S6rM4qv
JTjZc0SZ91WrgwPJeClKDZQKnsc+flShoizhnDttamKBUsJBJIrBieUfKUt9Y0N3
rnh2UlS+7xya5SX2lM/M1Ok5Jo5ct5aaUfTzBC04tVISXsT0vj/AXRlV99Hzje29
EiHYRKwnmFSDkD7cZwnZZEkhvyX2SXlFuTcLbylNjI3tZdNgUadgAa8PqXWoM57d
2Gs/AtvNl63pRqXMWoidvalG1wkE5NCJG1KIHE36t0yCEHp5Mr0gPnO+H8rypuV3
AaEEBiGFWpBXIL7JnWMLz1LLMqhcHM816HLK16AZwnaSvJATbOH5fDLOuyNM6H7g
UaKSK4yHgJoVYsS82xBGkFneWG/Zxxheifm/PRNB9C/uXBU0ZGoSn+a823B0El8n
wDc+S5g7Q1l8w5/fYfVLz13kkFiCSmTU5peiHbUpC/wDgqr2FYH3/fmAm3WHHvki
MKXcW2dnJnfd0ysV/HalqNkM8/fvY8Str74GH+gtL1gxBCgRKckXu83Xpt9z1pkN
dm1OF0nLj3aQon3uk1DHu50P5iyzgiHe24xXldfQTXGBWjogWHnEEQP7g3+ba+V7
iESBl3uQFucbCr/UeaU7vQV+yBSRf6G6c9kpHeyPwZWFBbVIEpc8TeIPeG9q9llv
qeJdX37r0S5KFN36eFpZ2H9oSuQqPgH2MT1OSVhcFnBCfG7CIGFXkpHWgC8zXOMN
wc99ApDS4QJVCaWlBqf8EEcNDE3Zc19Kilg+h8+0CGA7luWpEVKervcbx7ReJddV
l7/5eEM3bUqEkVIe/bb8hdUk85KdSg1De6zzDIq96pRwbhhviWuPK8ZmJDY94iyG
4GXz1nugkhoqs/F9E8iX2yB2t4fkV6x45Ao/+ui6k1Qga/b0IEb/L7V4nyp8C+i6
t1qQNaXdXHOqCmIh6iKvMQnBl6dpkgfrDn+kCnd2SJGP6iUi1bgeHCTYW/WtuOPL
41rUg05i2H+lvIZmeM+N79DosALaamSvpe02NBynUaMt+AnLcffyABNXWzopkjDG
ErhOYGVw/Se9ovN1RIJe9xibwQYkYS7nkdRyVLfOUZHERqvV6qkVfRQg2iKp+t4N
vBV972pgTnTscwJFU8DRiMGxErQSe0NUJW3eVMBtdy1D4NtSMzKh1anFWqY99njT
DkxdpXs8UATlxfLRAj2p4gKGNUDG0exaHOZ7XOplfDSEPJjjiK+9CQD/M67KvkMc
pUdl9SlI1UiTIPDdZ/37PnsjRYDg4ZMocHsgMjjZdxGDlA0nTw5LkzhsAYyAPQWX
hcuu2rQNiDXLjT66B+ynGkKACFPUVc/OcF7gndXw/csV8pFYORikDKL5+6t/ZPhL
b/fMJBwxyroINLbLOUmYJEs0jHWhVoS5+NO+7/mEdBMHJ1jUCuJ4IyoUce2FOs5J
j7WxdLOOOzlotcsnoncycjjiI/vSVGdG63+11Yl/nw5kd77+XQLstAll9L/Url95
r2RErcMXi92+1JXowD9O13C2a5DQ7ZpEiJOJXyoY2vIVfUhlUqzQq0urRr+bzzzn
sP/aF1IMQc5XwucoRMWAAlm4p5U1UJEdaoOnfGHk48EvNiWqFuwzyvYranDYig0N
BwKrhqeWmvXW+/jaLE5BcPym0cpQTijEktWpg92YbuAKJR/Z4ecPh8YsAmIBXOWf
NqAi9Vy/VoNGIt6QR+EaY83u2lvHYlo0ogkTv4Do4ZVNXv4nHZ3xNVpyHtzSSPWh
QpMYaVzGKxF58lMkgtyrDDsshrkgJ1NBaGLQhjriAFWfcLCVi04hdph/9uJRtGnP
jpOX9bDsljZ8o0NRkn/kdqHamkxLVXMiJVd7B2yaK19NuQM3NlJf7tNJv1nCun12
haIjogakltuj9muumHpm/KP7jFW7X0Hlmm/TWjd42jmaIgEcGM2bvzyNVCndYHjZ
rPc2e3kBq4Xe1+fNOiDLJ7xWRUARGjpOnqU2CyeHJRuN8zd3dlq2VDPCAQ9UJKdT
yeuGGETrHow9iG5FGpea4LbRvPsNvqyk76CnDG3D1d+mn8ihYHqDMffVeIHqG7Un
Scf4VVmR5HyAkfhI1YlQSLw3H8frpfMaPHOlSGGnjszk1kdlz2cVXaQXCbjaQ9cd
MhmJKBS1NqTuBHIwX1qwydEQ6ToY4LAa+OCHbdZyGZgzPAzADMg1cbA0b0vVKsLP
3BGCvieEg565ZaaJpt+IrWoSzzq4pk7EXI0dU3EfQWppesvefpNhwNs3huu+00SX
DBlFtDQGu8KjPo8toUbHpnvPhqOYhbr+B7jxUsTSO5cMEWVulIUHbwoGFhAj9JK8
Mhum22dd81D5A536NyWnV5PMpwztNX0C66prD/aSg1oM51IAFw4bKkdmhk/cU2U+
86o6ChtbhiJdT184DEjx1HzN5EFCSWcYEL+TlzdJP/22gGk7kq8iMOy9gy+RxsW7
s9AtGBC5nwbzLjZ9XpeKFhOzKLqMlDGId2Y9xoS2uil2voc9uu22+GeMYNKqY8Q5
mAwLPfx8e84RChMORD7QK5EutHFpU+q6l0igBcIV3tLJ4HOe9zwcWfzxHjrZ8agw
wkhWcbjkkyaJrwFRFsxvgPy4AikuMPICBTDBogwPgE3FUPJXFMnj7rC6+R5zRts/
didpY5UFH0tHv+NRZXo7yRpXTgiGiG3cNKVz3gnnWBPcpbCWpu9DOz2kJA5/abr1
8kIv0somBtYjFUchefL8PJERG5RuAi0Kiza2lhf0xc6qD+1edCKi7t6IzkjbM3S7
/Q1+Moc5Dzz/CnEwRYW4K0NWGUm4Ex4lqpuyY/kKk4t5jtRrtqD6dBJAPVdfbW48
WaCQmrVwCrBHHYXHH4DVG93zBdRd2Rz1PMr08jKP4PODH8iBoXBXJmIAuZav1nED
0hiBC0+iLLc+9aU06U1hR/p0HCnFyuYrqtin5QSjQkH2Cc70T5Mif2hkfJVum8tj
rEkNj4F2FYZpxkQxDagf1DC9oIMc3wB6yQ5CHve57WNjpcOetUhLfpbapTwox0U9
F5Z37vvHcnUHSjTuhlDxt11bpUDnNamsm7zJJ14GohOhvifu81+SFxU/ZBxoaYaC
3wjGf6HYwJkuPQnDTD8CJstP5FXKMVCYXt26jTrEzxp/i4jH4iHue0usHOKokR9A
ItVQyF3Pc6ExE7XjVCGFshw5CCvcKbUxCA+n1q+4APxdA4rfKSoWx2+h7xH3cpQ9
o9I1hjHiHiA68CgcsJnRGU+3R88ELZdBXhhSbWy8nca/gmEwoETmx8cobXkxsM+I
H9/mTy0gFCa0BEOsZnBpDfw9mVRPlvv2jQ5xmBpHcS9NvQ0zNl1boeu4jYShXq+U
wHs3sXMJY6DMMMXQFpu0zqSKkkGtYEHPk9hA1qvWb/rJ9GZ5VrIr+SUDUppo9GaY
j7sWxlsWe6mz4zyIBC5tVM+fGs8ldYG76TMUfpsriBLtCUPTneuGYeKzk0yIwK2R
/u4Rv2Wi+3leVPufQlkfWIqUNiSD1+AOmG1Txt7oCyFNUJ4FaCxFkwleGIC3IwYz
rBikD/7xUP64vVk1Bo0kyuRoa8buBRW3AD8t8wayQ1YQ4Nn+ZnQN1Ge64nSdeBml
YuQBlJT1awyRB/BDvccJw0xBV08XpPIaAY7S317Gvowd1cVeY9x/t7tas2VoJt80
HQdWDPQb+26NrAcGKleW8dN3dcRCyA2qzW1VoEWaNRHzsan+RctSSo/K7upSNN7F
wn5CsIbuzO00L+kSpdw522H+ubCKyfV0s0c+FepxDE+DAmcEQedDepgQxqzpJdq7
1uwTyzr3xWsduj+hyVveglsbgdTx6+oFg2DQWVvbtjwSeo6taHUiO63GRHCeC4Wb
RXyLmmrl0WRxFjId8Smg/Yke8nARgkLGMhgd8lTRheQ+Y4qHyPsyossKfjpkPyW8
B5L5Nffp0ojqX/VEXc/4RsLyZAxzE1cLeiZex6pc7aKu+TzhEtRedyV3Gl67V2M1
y3EnmkRsnEEcTPSxXewfQLYaVyGUGVrir6oPOhlXc8ThMnBIS4CKvkKPXBzigphX
/1+VjtWDC77SJdkpbwQHi2V/fK5fexX/YJCh0ggF//JiYjBLEQ69A9pVZf4s/Ujo
2rGdnKzJ1rI3tyXEq5BpggjnyQH/XXAI7UvJeUBKur/cNMB21RB2xWgLkgll3cdp
VG14QbGvR5V/nEgZMrFc2OtKmLx6wUdE1btcf2zlyWMig1pOrpeqP979iZiGAL8g
j88mqQoGIhF9PSFCFQ0DE+UDSdrVZ+Jj2z1vNokO0d5zJf5CwRiA5punbW2cb9rI
/+GjtGdAWBjWSYkiJjBcqfPPMbVgN/kI4cQRL/blrR7UxIcqG36ZaWOtNSQBojnd
cWLBp4qF9qrwvCg/aAu5QaBIHCSbI8yPJA2drUjXjTr1mbkrPCiylnWsU3NFKUr+
qV/O1ioq78+ApqVxMdp6O4wCafQdVOBteMlVspzs2OOUNO5AQlHCvTpzxTR5bdcJ
Kha9uVpFu4aOXLW2Sy2Kh7RA7yJLKeW+BLXn7OgWWhuRN/6HIKtYw8896EPu/9T3
uVArZkYsmP55rw+weSD5JoW2/NGv99arH5QsRnyNFQ8qMNvEu7K4BjUhiD196AaL
mzE40ysdNMbgRVT26Vbvae12SppIPn/g1/g4vtfPP7EEOEeuTwTadQBqecbAo1kj
V0RXJg/YQ9TufA0smMK1FDyiO7quKMDouH0BCb+f41XBjxBjWbp4GIO89YpbfDGy
IwF5yRyPCq4h7+QQPXsiMmLrUzcaxfuV/mLFbw/fJZS5EKnBEHLOIuUL0JHN3sqs
XK3eyAP9kuD57kRm8ioGc7gk4E26u9qb61Jmn0Znx67NeqOeVwg+HakJaKvAkgXU
3Dbk4dWd4rOqOwxeYlv/AkGpcoA3D6gaK6usdof4rOvdQQwu0XnleM2ugHtsqJtd
Rsbs2+N8IqGSFe7ZnbABraqqE0/9FWbNeOfnXrJF9IbbHcanmRStpP6EMMa1l6Bi
T4JMEURqzqC3Gqx4HHOeSZTt1KioisRwtpoz6wSjNDCOwl3+uAyZnvIytwHQzaDY
yEpgjABwzjeH0UaV9csKvAWOCmUAUVzWL5URjULUszCsOUzOSoOyO+u+5IGnCfm6
ZjuZuhSMFdIfgU3b91Jc/jJio0Sl0emKFexrfL8Xm9WImvKHTmeNpEP8UR8wrPnH
qkztpEZMvbA2bQR1DSICHUGNIDuWNOuqt93V0ymG2tVIvoXN0+Svf6MUqamOdXWi
yhe1/q47z22+Nd/BRNS2aU6pyVLxtuAABVoUE2BOXXFjWj1zf1EvUBJDHZlBbSoA
z2FqrekYjyQGYHsYQxBbNwtaqR6CRt1QIUYwuepB7MQGaCAXjTzCCE/p78a66i7v
HqrNczGG89x/Rr+Xusbst+9BaDXGcSkTGUNTL8BXYLJooZqSMfag8KHznGO2PAPV
ZIAwzEBrRPOUkc/kIPtq1fIFgLQMtowhDjGn4Ca/UlFG8MQ5MoXqhJuaRV+BRoqs
baOwJCMFSAhLmKA/C4FeJt0kpmXoaljF4iZp6EQhHMbNFPXcLE3WdtmfGssAhRQW
oTs/I4iu3EChIBjdadTdHoz0Zuv7h39QlIhRJZeA7WFUF1QLFrxZK6y/lXIF3nkc
lX5zpMwn+/boHjmIMPHO+HcutqaSdA2L7ZQB1PB6k4f8FdniBe6DIuIZ5QIP2cT1
UFrtBzjL4e0QLEGdWZzkSF17ZdxcTQwt/wuWyinDXFFcawRx7cO3es6hcBT4CHGJ
PxxQTlUKHtx1MXYLosI72kn0qIN57gvKorMAWexU3Tpk9UDepe5Zu7TSxt6F68U3
wtL09C9Wipj0MYYaRDe8nmDcRC1YqrS1uyw8DVND6MOm2NbfkVTlFOWaW47HJYGc
6pV8SbriLXuW/qrMChMtCU4JJsG7cd1RWs161m9MYq7KmvwA2C+agac3sCwlc2UL
HG6UFxGwEBl1TfYKCveDm2iUOyVjDsRVKE2kESDNFQ8UX0cqHPL0Y/2kY0DEQyLC
g2HN16RIAMLTe5DJSLlBejRDpueCzDJbitFDrE5RhRi50Wffv9OAo+WLU4E7l7YZ
Ngru/b1STd1lzxVmVpz8RPQhIUw9C1OEpb2mohEZ8KLsBCyzcl7lhfFPHStL/G0K
ujCiTtikiPrOcWYtaILC8NaAw+piN7RQZUjAXtmXK/dj+e08HpRN6bY1ImpDZftT
fgITqbmnVPUpL5JA8X+hG6v63z7HpEkNfOTFvU/fH+TG9+EfbmdUryyYUk1l+syg
kdrwlmtp5nEHMnulEWq7oYUnikbrwPJ0j6KCB29NomHE2TDXEp1SXma4Xn+aA0MM
8412i+bZsozW1C9LPEghWWexuoaGaXM226ohMJlREX7ZsuEdNbN015i0TaBA3CLy
4XQMFRmj79YLgK7UKSszUTYYX7BPKsEi9y7TRAtRjeAotCnKbW2CMGb5schCG7MO
dqTVNUyTuhu4xKNci/Oxu52SsnjhUcPIpPB8nSP2tsVaXR4oSEx2JMZW9714YfPs
jy+07RGawFacp2cT/Gh4lVo42da6zoON0eCfRS8PEDI0B3knvpfLDO47ge5/sImP
RgNYDt/dcOFZoRmHHgqgXokuq1jJPuiKFLG7zXejuwJyIg9/yVxFHn/UJl6zrJLQ
eTtbr8Lpo7jRzzovpMb/JRfmyIsNBHKDIgDEkgxo8UA2vKy9OOSzL9xWsagYux9v
MWtViAYQNAtovwMfL9NaXEjL+PWyDDvo2t+fxlBWknee+EmLg4gzymBnwiRMq8gj
ZqqkzwTdL6VPVh5Wx/72FeAC/V98Ze7ulcjRpaBGc5fNf5FJI53VlUT6X+7qfTEu
y8nlzSRWY8/xE6lBSkhLl25wZTtlh7rl6luDi9n5W0Cm5fS/APtWcfdi0Z5TwaXX
4Rg6ZjxKcuO5uEt7Ey3ynrs6G2YlYQQF6pZw3mh1H5fxfwqiOX2mrNzvw7pxYGPn
Aq6aRAMQYKHj7LEBWX2edSDWNUppObWMwjOtS/6YtLE1h7D/yURvTYXCywYHuaRt
Ng9y41GGd/OwcmfX/NcmoJoa+15IuCN/vltQCScG1Cyp66DBDlbFrR3XcPPcQIMT
sN+jf4WyI50HZQ4pomx2PCbDpgzWd+Q8bV0jatQqWIxApKRDw9WO6v72ioLW5i2Z
3oAMT3Io7sP6EOi1zsxDjaSvzbWOmPHl+v9rxTfV5gU0MgH0Qci9V4BXwwDifX1w
EFfQ3eID8mkzsuOnzK4oIXe1KozfDaDjfl8tbF0gQiWJpXvssh7OgkQwwFrNBg19
YshjoJUVNUcW12SsRrvjGwTWH9eoI6cT2K8bwoy80YUhqv0Q8dpbb9gwiRFiTnMV
RbInzWnYI3yBubRHiJutf/kscD7xwA3CVwkZVYfS009Uzi2NV88kxAIEdXJd154z
G39Jo//e96wgxi+RhjFH9lDoZI0UVlP+6Uj+4T9gzMzIcazVxEAcv7FfPpnebV0+
9HUGuX1q/ucX/Ob9M7ssIEaL9N1DCP+qb4N8Aywk3srSfOA7LO2FbmETtADNJbCk
dACT/HHR8bcyUWZC68yxe2fyWFP6AVNE2uuBXeX9n4obhiT9z9c3lKzNNWDqj6Km
+1eUjusjaOuH8mvQ+rWVVIyNncFEPjCDS8vdYTxWAKEmyORCwqGhPYIjk5U2WrCs
HAomYtCgl4xIyI8+dtGuc2KnGUjCl4LifEc+TYSxhdwPO+AbQmLJldoY8id1cc7P
d2SID4uOqqJnu0bFvAacI6VlWlJ1G78/562nd+n2r6R4uOpR3sIO8igHZi1tXUN+
RGuh4DM46phl+3o6AxKAog4BwZrUOXi1ZrcJBO3Za9XW0xcIbxwf6WiWwpg6w8Ya
S4NiCPTijRRfr+R/KVXXX3XAOVdYoSgf28iBo29ZN/UOhSX9tEaS2kizFEVN5A8Z
WX2cBxb2fenxNvJRPxkWYjWPHSXC8yBIkiJw9tra+hwVgt6AdrDK6EkVCMyA6q6H
nPtJJmIf558ndVolM/ejXa6jH2H1DgxqDI0HbpRIQ6y21LdDw+R+BEz3As58tzo2
OP8zlMSqK5SFoaxwMhgjX4gUC6R+I0tyItLSuU2mhvHmlXjbbZ1qQoClCtA9CmYT
XswCiRW/aseUgjn6zZ0lFvCIpx7jGRga4B9/2T8NYPFNH4SU6+QavFx00Ky9JYW0
EUAR/UbDaB+2tOZgTfoJ558O+b5u6dwpMQjdCSDgO+n2WoxkbGx152Mw27gvoWRM
orDQy85CtcRIN/sVmEWjTH72WCoLrvaHI6RY8zCfFyNuBmFsjtOoR5LeaQe5vkFw
5i6r1p/a5cUJyE3CeszlCysIirKthsDaOAFmQEG4hpMwOd3O0ldowpWDnMrAHTgy
pc9b+7cFIPNHvFBieah451r2585yjfhfDTXtbXCTzxoMMquCXlwgu1rvbH8LLVUN
Q6emqFAk7bGsndBi/jCQRiJdsDBbFHpVRNhiujDPLp7wJJj1V5aqQEeA9mA+dt7p
w3iaqDP4CsFWhitwDSmOvqKWp8eBNDXX7dIChenMno9GcB8weQ0LgWEttQfHvceO
Ch2zMYlU4KomHcx6X6b6uP9P9ZOkUn0/RPr7YwbOq6ulV6u6NIG5UWo1OSU8FH+n
Tv/faJpwin96eXylyfVk1KnmvjfeJFICI0kvbwQUCL/T/QeiT2dsAWfBLscx8aua
pYVnbGeDQKadAfjK6fl+Y5G/jOUL/R9pv0yLTuXUlLIXpRVvtOPsK9fQ6an1Ixql
VwLMwoIJznCp3xbxX5z1mgbQQ1Rw2x8i3FP8NVaRSq/lcK91sNcwSlULBCjdwAYf
VMzkyuONUDNf3CNmik43sE8DbbghyaBdDYqd7lvgT0WGQTHngfZh1Xr/CagmiOQ5
EyGTDuUN4L00Y21szc0ImUTo8DbqW9MOOwFC5BR9MJqRRL7AJI+CeK7awcYrqTzW
vTAcJIRWWbwxuYtjoogRhMA/tmBkI2/ummFc22cBHPMF6gkIGQG/KaXIDBvBe4Fp
4N9duUdlSmgfWpnoIo23qhTTPQulk32yhQHSGq0hjXO1GM8h1gKNPLpu6KBO+B0l
yl1bwkmOMUqDpC3ZIai3m2u9WGJ5Ct17Kml6MjGC4s5J6KfN9zAKuTlfXkFnXIVl
4lQQM85hLtbsJ8dfYdfRPAuS58AUqFXQtNEjotgrpqnteN6ERJKcfr+uZTrCxesN
qZPiGjaS6IHEZPCAPPLIdAYw+WfZOWRNR274GGA3ixQU0FKgxtfZCG5xKCPgdXHj
WCpQX3tlO4RMCRTiwKMksLmt3edEE5MXUTnKx8FfHm1BVQAXquiB1sYRraGKrvWP
/qJZaW7PzLKX1zqZGUHoX+PKHl4z+ZaN0PQ4M4auU13d83qWxiig7uYS0AtO5FUj
+Q6eGVSEJLj6QmF0qc4ga5mgjqwpC3+lR9DLaHoZL2QPX04itvFrmIt+JiK84qgY
9y0j1Sbp92n5epe82u2SGfN9uAhGtUo1t7fet4ItHcn7H5NG6GYvlHmau9+LAnX4
5Y2b2znkk1P5Nl2fz2DInB+Cbuk/F9XmLLwp2apxK5MjPNSAYYDruIJH9YGZ2pQp
TOWz9SFM6NaHt4bHzulmIlblpdl8cs1PgZ56QMabLGeMWeRyhoYvFrnk9NkevEH6
drdkkgFKop9w7cBoOkPOwgUHXTaAlB5JZvBn2SqW72ApixJlfnWHtctxqg+XBG15
qQ2CANHru1qxBJMODY5T13ADBDupZJE74ZWSIqzMiyNgIpLrYQgWv+WlbEtaRyLM
JYsYoujTTpTH+k7BcVOww8lwtoCpwTnn0UGAJLZmpFLJ9f8nNAWWyB/R/+7EDrWI
sKvnMfM2lGDL2fDbW0PjW0coCE5BZzSo2JpDKDQJhW1AYkqh+QznZDD5FI/C9zqZ
mYZpHzpGNpNcpIKXlAXgScbwr7g6DqhzZzjbWEKPb0Bsd9pJ/YiKgXC01xIXGESP
wcGkZuuLdlC5h8VmXO3bkEKsEEq4X3Wmgt0zX7Rc1hrwyRVpQfFVXOWWnUcCR+vb
hLcZbKSLp5G/7lEB+9p/wIpYyetRgNWMX2TjpN23UE/nF4km2JvKkw+X3xoTIw9A
dCgyWHdRM/Z5WglvCXVVIMjCp50ymnv6zMUpyshjXGdG6t0uNnbwxWJ3d28O5HIE
mB+aV1tSiYRGZJymRQayuBFEZmqyKlANLsQ2Mu4UdIMfX2hU5PZDK2z4MyOGXwp7
4GsZyEUcFBFy6BQ1rhxvLfE8qACKYMri4QWQ1uhdastbpIQTJuOrrced+BxrQac5
QN9gxZcXTVFMxPdQ3bRbrJRk6VY+y0KB/C0sAZe3dpNsdMdEJkDDSJEKyxUiaXgF
01KpGqvWHrL6Bp0OmHBbtzbh3eXix1cOm8zNrMUOgp2JJYAnWG6tmRk2ukZ4BwJ0
BW/Lqfg6w+pWwjqwJ2JJP7bZm8bKCI9D8Z27CwNRrQMR890cRRj9SpzdvCdOR4fx
oDUaxax8joRimnmIFk3D0TgGnT7+WvMypHx9gi4B47h8mq7q6lj0zk7cbeO93hA8
+howVCoejbJeuQrjRZPkXoZ8RVyy2MA/NqPf9CAaIW+Cd03FAi8HpGCaXAJSYKWK
zG0M/JwoXN3QAFxHfNLEV1hhPUzMg0lfcKjPc0//LWpfF0GbR1oV3BUukqkuw7Ui
uyUqDlFDBLmZrltPV5PisHUaq94q3gi0xXYFIudOpsmirkOGKZ9uHSCWFPAebpas
wXBTyi04zfKaegLjcXY+ZSS/6k8X970HTPnooJrBMHBVfC8QH/eMRxFYeL+MHqI0
/4PFniM/7Vub0I+99GN9VJOUhIYlZiXqQJSb/NvYIQ5Sy4yuQXC60zJSAqzl1s02
f5w5XDaMRIe00sKN1rhbpxw89Vcg/WqjN6ph4YxN4jIFhxoVu2AFLU/LBvRq1uQW
7uJ7OR6ZyuehWz5uiB9rcaZHRKCAZmvYLOeUaGAPZMOE93IoFzn0mj6C/uDG4l84
0uJ44B4yTo+H5oVnpLrKiaBe8eNqOeuU3DOHjJoqWc/T4DhKDeY6HMDrid33n8LA
y3PTpOPT6xW/mbn+NXmDysx7LjOOs8CkHneUtGCxiNbmAuBaSt3fMnRIygCn3hBA
xX8UaKzF8VSZKfYn/B1CeUsaxa7FGtRIH51+qflJBwfpM39fdNlu9e6yzsyLobWa
aDTszLoJFes3K8TGtSCWiXPHtCylZBFQCDIACHG7seGW4loj0sXAN7rJUwN0Bt6a
4bOfWpUPcpcrKATDh8/xxYCmz0LeIiKey/J47XQmgB9lVX4TEfWlSmvoM4Kwupl2
5siRAgktNJtPH71zypgj1hO+3JsKrWfYgBJDkjU3Kr5uABSan4It6n7IktsLPysd
YIiXro2pQZ4Q3pLqFwzkvwVTPqv+glpVaLCeOVO8E7DmYLNRR18O4Nw2A0cg5ZgC
37QrVx3cmhjeA3fdVjYTVGQYynOUrQRJWbfKzbWl/LX2Xxu7upoqjucL/ctWCWXB
4UT2yomMJa9LQIhRxWXJmq+MzjcHuFevjaUbFBZ5M2poMbP3xKsrgvCMDe6smG7q
FUk2hbcpI2x54Mh2i/KN0JvD1VUM6KJvPF0gTUtgnzhu6SxXfM/IQjDdRa+XNZG/
WFaJr0mWB/nAnhDEYQWWlZczXBL/ASEQ4LCxGbB2qdQFgoPNy13H6w4TzLDsCd2+
jlR1Ax0JcZNX6OSOmQMqkcIXxe5YOgb17pEEbzYQfkR8jgPjnfvvCNhJz07dWtgI
rpHO4r3WrCx6W4RPqTNENZ4Fu2EYnjAm2bDp59KwBEe55J0A5fyOY9C+UxcGYkE8
kTsQTxNfO6U6fCW/mbgnfPBkqnPSZiM96Vh1Ct0JmYdNITzZPbCfC7BaRh2RHQI/
mVE6fiF/yX4BmRUyFWrjpW7hxm+ZBDHQe2/Vg8dz7gwOSg1Y9Z1fmOJElBAzaAKD
/MqK1WO/qIRHI4DPl+5HNQpmETfYg8b6Sstwiz1+fsWdluAE0tef3KZfDYcjCfy4
CKWFa+MNZsXabrtRsMa7Y38JVoZuxeOFN5xyRAEcjkoaNShw4vXKEznG7sZF3qer
O7+sOURyM9XJpu8aAY49ez94yPie2sPrB9wmH4u7uQ/oPip2/xDodGEobf6lK9cW
YsW/EUdrgHvgdR4/Cy5LeRL2CS1j21XuEkKCn7ofRD312U5Q5kXeR5e4Bk9L/+oH
yWGudWIfpIBC5hmfZRUnY+8waigc7/DcNHz7FEwKvoqoQUdy9KadkYFhW+1UCe7G
vTzvmulIy9OtJP5bZQqVpGXup8Pul9DL//vcQA3pMdcPhUS4PX62eT2RtLZRCEks
Rn33kGmogrJgYF3ugH2gu/vdK+jwapPgVVBz2acCO78GS6QRTxDyXTxHxj+8KhGb
2/FX1P6+SZHgvSgIwpiXeM0gmCt5cj17AOa2rw3gpRRjdAlxqGHtE3M7b13KmCU5
bB1dvQzzEAufbY2RbuOpvAIxZnSg88KkyvfIgffXyg3F3AzvitI3eyvwBQ6KWvPV
BK6uLRO4iUtgmODCP3XjTubiH/lO/JPjtWVF98glpkWV/8rr1nrosz/z+lAgGLTm
o026fZOUoqR7A9OHPhDxAHUaMDkXR3PgPEohQ18uG4MzGGjXxOD9tlws5vRVtn9S
WWqte5LhXMgkmFk3oJ/NH94rwl07M7MqZoVAWeg86e5vS1YIpb+eYUSHHrB/F49Y
FvAiM5ZjpOsQvYs79PyvqmuyasvbOTxB1tPs3BNJ9vqBYme2F7f89WPway3IhaJl
0cW4+ZB6UANvwi9ZfnVLB5Crza84GVQgHq1wI3iCUABJZi/O4mkeBRjb811NuIZM
bpo0RYlf3ntncHDkqLbJ2Z9Ut5XWJId6SCZwvkoFS3ixoPtuaZI8HnVKWpr+0Yyd
MnHsXzRXbusewVqbyEbYUoHEj6wDQTcoRK64JNdtgAhaqus1bmIhDuC8yoJ9zGEu
GV8Q7a4sAIudIFu2AwgRhgr3L9WtlEeTcBBoA69L8hi19nF/02UeZm/dG8FdRwVt
DcUX2jFVO/5HyFxVCepyU5SMGvxBMim//zro2tdKFPWlUhyBfRMgLUp5R0qGXTjI
cLab9blwOyk8OnA0hUUrLQatY0zgCb3TWYx3NoOvXQCeyHgt/Zr7DZ5d4Lg6M6n3
w05TjxCs6I5PYiVXNYV8AvqFGjqkZo5iB2T3HCGuSYm2eUrJSEnB5+3rmKXcH49p
0Bvi64XrY+Di7G3xDFm5OvdBxiZjfikgguI834KZKI5o8bjgc1V4XjEdg7QsaxZ/
0rrFKWkR7vAvifvqmC0JUJeRP9hvjXM+alfTHAuGtKugCR7Z5VBKtrBi7sn4qgBP
tziYnqeNljNuBv/TmNZPltEJ2KbDcHAg9C9wYZYZbebIQttO76sY6yIBmJBZ7LYX
JVwbfEAUxCGoNDlu1r3JUFw4G7/63qC3d4pCT/JnHuZjsLqbPzXLOH+Z0SSc/p4K
vmQI4kmhJJ6rNtU+9CCF6UOmtaLnsUOb+ts9cML1PLNhZvNThqRXKY2eAgza+nX8
upM/Q4ikjLJl4AMIS3t32Z1BvCk1OaU+leVIZqdACFjVXB5suSopxU/BUicXWbws
LH0M9OWcHaPXmCeLOekXGYjMuZ5jDJSfq3TSRr8ybB7XoYsRDZ/9fHrVwmKpd/NV
4ygR3AOJWJ1QFAvbzGL2/9/lsyTTAtYsT8g8OZE6klP6gvOBMJHeoNYOiymRFYc+
6EX4nIxO2Cxk/4MZCdzls6ZCYHldL4tQqoxKkkU+Yc0vqWWPDpnxAkyzAX9K5Ab9
sxHNeVu6zDuM9CXcENvldnLAzPscUvHbhXNqRi7erbBgL6KFgvqAaOL9f9ZwTclO
PEXghJhYuBHuLI3GEKoNnNgybK+4950w5BVfVrLbAyE+/eG48kKhzxot4+sEf4Aj
f7j13m1v1ol+EZfpNs8Zf652YssChi6Pc+OY+Td8G9J+MQiVnwW5gK4hYsCdYH65
ELCWn3RqqLgX1tvNvHpenozjl+ZwuPAHb3289HLXtFQFLNGNJlB4l/TENIs+hAjO
bfP16B1kD3gNz1b0vNdW0m11pecpHKUoaef34nic4zIvS9KlQ+SpbLvbuyMwCVOy
hy6o2CB7a7kxLUvrQ5y0kUHROz7u8hLURL4qe/rbZSCqAQiB69/hzopEaQKyBA1B
/ABpRPvRcz6wkWePPB5K+lgvnAoKYMBqARg/DfVczMjQ3bfACQX8sCqIbLuIVzLL
f1sd90T/MZvJ7Q4+7ZSlIj7EjT3O8LXaiLGz5IhhsQ9163SWFLOFzLY8zixPwr4w
agy5SK9/b3wAS7OgVgAFPWYIfDARlklpqUELU0HEHOCO9zf54OxE4LPW35qi8PrL
9S4A5VaoW2UNzlm9WRkL8HCboz1cyyv+aQJW0hoxweG1xa1xiGsHTv6mR6GXbdCI
+s6mleV1tFODMu8PdsHzkO3161e5TGM78wlh5KVpXmM8IqE1+ZFAwk9ylvqigmxF
yJ818XyuVbu+Dl2eidjb9UxOCy/LkrBUscakp3UhVLZMSQ2N6ZcsX3Gr0/saoLh6
Oh9rVh6RQY+GgrXxEFXmT3XZ6tFLDi9XgBXvtOBRt4WMlqz7IuyisAa7qNYgLbbr
iP9kwAfzA8VbhdGDDo5QfCcVZ8u/+fvao2fV2GpuSHP3tit/Ouf19mxwqe0GvIGU
iS+pSl3QYgGuiC7saU6ik9MuCqb7wEdwkCa3v5eathUOm2/51FQvJNbHg/yo9q2H
uH+T/EytLqhgsVw9eD69RaCszkav2/qYsFSgetvGUqA5F1EqbKuPhOqnj9xqTkpU
dvg/D9IAPAWmR0RdYQHeuoHF/FPB3ef6GHPLJgexYeZHvbVAvS0AxRQaPqyqM7eJ
1JnfmpfZWsVHwVGT1jsB9XFyK20twIVPTd2m3XHEtopeWmx3k7+t8bbQtk+2ZHoG
qEsCZ8Rp5sSJWflgqHhwITs5AwLIjsohL01mJ6taCqFEZcxs24nkyLUgCfDQqhjJ
dvKszeGnzgtO3CMWFZ7KiHfaP1TyWl3xb1JuD9WibkQBl+FB9QogNPqGCsWFwSeZ
n08DokU8Y6R/rjN5X97n3ptDHAlkYS5atuTpBcxOMd0p8vM5fHfBDmSZEdzZp/Mm
p+Ac2xURF8+v/3121HRUnNa37BwaFrPokGWrOcLcpflP+kjpU+yZ/5JyTuYkR1Xy
4c5FmGN1h28cPqIDDDhanc4HvZ4Wwy7INnBrwEUKTov+V5E3g6U7moUF9o9f+LYG
WK7cRBqJ5J7p76vzgwBFpL0iX8grYWoV1/NgcU8PV444nsTF3GNnzTRlpgSo7Uy3
kB7FWuUCrrb+qQUapn98qwkrXOZWNSvqhZYFdgbppLBCZ4I2nG4sBpslX/thMOlw
6Z/R/+tHUXp5T72ZGlbguDMKLCAM/2aq8hBAf0AcZWNjcr0jfXj7tDrtFCqEKH2a
puPsg6YyBcSfkmAwCW/Lhouql/dWx3hfPPaJ6Ractg4eBcZJLFUjnrEdTQvaDS2u
eytkjn03YaqT+lvROWxoPz6s95k+a8m2daQCDWnXC9f+05j08K1l0sX28l/niETJ
dxLP/E8b3PdoV0oNG8lNlpDta1/cPuXPLIbUdlXvZexaS6MnAHBZCqydkqtyLdUH
mJtWiS5mtuiM1ikFy3tnsRsTWQYM1fGsSN3wLiTNtUvTPWNvzge21YVKI+b+1bPv
CPEbd1brgtROrIpV4XnLO0MRckc3zJAWRCSlmS1pjPj4KheI3OPrzbgyDpjBJ3Gy
Pf+OPbHi06u40n0I9AGGW+3wdU8ysryrwSRiBzVGvsipGbfCBDO8r/N3gxjOEFNC
fYA7Ske21GWP+VU/SKfUlbl/TrxBeGwnh+UdwTVijr8yyr7c9h2rLTlZkZUzFr8L
jcgoSh+zpOFctC0CJwDQlb5u6JaSHfVH5//5rMd8ZJXboZ/j4punS0cpchw5jS14
ziExJbJQZzajU23GqFKNssUzad7hVPzh/6WbGen+777kVZfEVWNhTty9vqghDy6l
C4YUNlpMrJLkhY02xvlLsG1Q6G5VHS6uny24LPA8FTHoJnMam0dv4JP3560bZVWk
VFWbfJXql1tzxy4RfN3ZrSJYP2r9jdEjKCrbWnr51aAfNwsJBYgVYX25LBakHDZU
6ak0tCOMnZBLfVi6aVHgirIZKeuUFRmR7miOQrGT/T7jwBKkFAP9IeBFDswy3T1v
8jKTaAonuhXDCHUOMKN9rQ3pTBR79fnkwMrt2pjR/lmSjG8p51beUHnSKC1vbkRA
wp3V/iC0c5zIWWFGb18T/9fTYWeap526rHOU9Soq9R5BWev1uXCMVicU2CaecyLD
Yrah22cwGMNdDJDpi46YMmzUEE5epvhp3AiEUYMupzaLZwpE5m6NRookZsF2mG8M
zQqUO2mA4CK1iwwDztRtrS4asQ1TIaBm2NTT+HeHzLKRGSWKMuH9++x9ys0R4819
lVv8Qs/MHXvq0PgOYDPRO7YEHUHfZ5+jvVttwflENnjD4cWFBqqu2GqlMnAFBqRZ
p0SyNedwMbGszd9YJSVWwS1jRNPJKx7RgypKjgU5Bj5PQ9SyDACHbKdO9KnH1vI/
2q3xMjJ+jaG/bWxDK0L4ePlGJegqm4rad/Dqj1X1QCUntuiLl9WBwNMoJqRURgkX
4uwu+VpjQHouCWFac7QYQMu2v4npxv2EPbkYdC1J+2wFOWHvG4JcgN4/eGD+3rdk
u7HaBBNbvNx7HA6YIE6uN6CZ7vr9eDEldrjtHfh/3KhW2Na/BWy5jCAkCuDyB+vb
5VTiAlsLiZK+cgKRIlsw3VMbSHw5oIRHr1wcijLVcTfDqvSYBpQsxLpHoaWAaxpE
SDUwilve1oeFLN3QqztQ5UEfXUYXgIc9NH3vM9V54DwOuPCbGYKfapgcge19zpw0
JlyvUO5nePeE1O0MQDFNa9rXuQXpyiYyQzZQIAgVY+AuT5ljl+1HXhrLp+NPbyxi
Tp63OmZortvlIPpO5/DLY2dndARoNhJpoUxGefgACMwYrAcYETO7kCY/uVBBw17Y
SnK1fJNjKkFt+paFaV7HJzNp5KmGxQNVpA0oZ52elPRVwcg6rn7ukXRH0vMSinR8
qjJcJd2WEh2UZcsWXwMg9pUD3/uCd6qfpyzB6r/vJUjZLkihazg8kqSiG7ShjVyv
2yYIRWabD2fbTIHwRGCuJ09sjFxrqXS11y+Tc+m50hZ6JX3XMlYceUuMQUx7snB+
BP+PyCkRbM/z6g9eUDyzpzR86uqId12v4o+Oz6ofifR/MOAVvDh7w3nrwsubDkWS
FMQNn27oKTbNkRI+qUsmXonzAvq9hu5NuSO3stvJ9drV2IEwjbJBIWMv4x8eLV2i
h9SNU0qI6fd1VT+wfPgbFy2Rkunt2br4IE6XHzne0OefnDZ0Z6nFayYIoBL80t6V
f5Z53u5TlZb8zFyN7iOQcAvJLHIBC9GMuHnRR/Iu6x6JcCQCiqhar1SpPeXMH0II
eM8ipEzutJ2KU6gxzgbdpcHgOX1nNQen2FvdPsEFcroYbjY0k6iZZwAvgkX+IQWm
NvVg+OgWL3eCzE1Fmz+3EiobyHY0VXkF2ohTx/ND3l3Z4ewEaZ7LaJqA5a7wc/IU
OU27omvRBSszGJpnMX+IYCRJeDplqDk8THPPg18b2kDbQnElYoz03bf8X1qD/yAd
VEo6Mf/0a63kpglTX92gLomzMAnG8btIapmq+iFZt1JBIlzTnRcqlumad9ia5P5A
6+Qu4T+8rlxLH9OGMJfRPyDQmmvGTmza4YC9FuEpE+5wXfgWYb1ceHY7PPumd0uL
6ag5jUmrGKuZU+E910bluBSbF2xW+quxaEmmXbRFucxvMAdg4Is7VFw3qC2+8lB9
uVaAJU0cI+90N8oli/Zc3nT56z+WMPFLTu90uOH68zkCaiGwhKzxrEE0NRMHtcE2
3ou02CEELWRkqzwxeX3BiiF771Rw2vj/loVxyigPwcYo9azxu56hc5VA22JV33PK
7dSBhAFFGfWFr5G1nih6Mdk3iOaSXI1NQi1AX7a4v3HY8owJTHvNB0X2N++1eo2h
Sabxh51acXwOGKluThTCtBPfLo/O6ywGsaemaQlrMLyvbeUFgkrkb6mpNi/xUYIh
SEvoVOKETLaFzxraT9NheV+oojicULM7+u1QVFlJuL4jWG259ghSMr9g6pXbns21
toREgGTzQWXZeoRAagXxjf4+Je6MLz4W8ZxaSe14cRawYEdILgduEZhiCI4Rt8jl
d0578+V5zoTUJf24X9uAERmCFoC+ZP16HYBsFrmREAVQymYxO87ShCKlEjJMr2ZR
cmbRLO5EeG8y00Y9Qs9J8zZskN1s87huzm6NMW8HKBuLZWCqJX8A0QlAxHA3+5cw
zedrfYttROQRqt4RPJIW0Lg6BTo/RqE0PDGcH6Q9Ysq3oXg3z5F1FtUMoLkTurTz
9NOnBbK8E+eAQaLOI4sLR/k/2kTZ6HCHZvdvZvJDYRjEkAMkmsr9L5IDIJQ3YB1p
wH313sdgo80NqkhAaSKLn8+2z3/rng/H5HmsuOp/K3MqB5dXKmWnz7DiwIbhm1Fp
Itk6Bv+pn7R3u3ZaI4xSqoxCcEAaj+O2zPycpsjzm83wuL2/xfPXoly2R4SgSsI/
WGxGWQrL+0oDXu3KiHZecTPz/sEJZ/N6Z8B9YRgSV0XgAz3IScltI17xcY5rGn7t
l+cr7hz3pIDd/UQiuSExdyFSXD5DLXu6ebzi5rn01QNqiWxFAczA8kbo1wCiYZxL
AIr1+Nry6W4YSkBiRCV8PTp73pqnhPmOQ+hhV2+9XlDmyTq9Xicm4VB7lH9EW96H
5CRRQq4vYuEjlngBxnwa8y/gQQdgg839oJGo3ukkfQGpHDX/U0SivDvQ9NrSmE50
NJA7PHTEPemlFbqQOSr5dqH0N1aUOUCfgiwdH6u4eaTfySivxVM3ro4ovMexjhys
7dgLyfBCIr2ALSjRCMpCQTGHoR8584PXNFMXzVHrUbGMkYhVAz8AXVgKX4r/YdtH
ULStG95CO/zCeXIYFuPMcKaOmuVnOdt68vVrT05qhsXPT9bsb0Pt3aX8FXyJCtH3
ONIrsOaBnwq3lClnAbfGnBfi4MDXUORswWwJYpsQedbNCMZo5N2t9e77QezC5GpT
v9xV6hD2f5SPE+xmlfJzfmBfjbZQqqymNyrm7rsGdAUIYaPfjkWy9T3DUZrZ5uRG
/mjJASF0rEou4ir8+U2oxgY6Jo0K+YldYiiEdttIEJtAv1QRkNZsvWiipT+TvKrE
p8x4FworIdgVaSBSgxPVxuR4fsRSWF5T0KRgbu8F8b34ZuH3UTT1+Nbbq+vB3O+4
FymB9GPjZMeHmkfnqiAQ+lXSRvqs9jsVhBeXMFS6sFJg0i/5cNfjtWXhVq68CWE+
A6RFvMeUSZ3w9BaWuBHnP50SsY7Pq2gOmvERRlK39wc4PK8fSqC5PIpJgV7I/3zN
0+BwOJsvUcb40JN1dhmrfZ7yqXLhoHmovbeRUG1BhP7CorwAOJ3cPUideKkirV7n
/CqCTwxmnDQLSHthLYicom90r7tAQcpaszoHeXLfIVdqtQIVv1RKCXqmGz2LmFDu
ROS7Vjyc23duQbLWHvclpRtcWBZDmHgA03ki8ZGczDtAjBu+olkJNuKN0AOv6A/3
8BPp1qNbMOxjaAPCQ7h7XiNYDWxQ8hL49NTf1v03A+g2D7bnxXQEHdMaFEnqEm1g
Q/i+BZtQIyw730dTfnPCFOu6NE3rOMR+B+BZAQSj4kEsoOm28WAlPbO5wKnd3dVM
o0Ho4iXlH7zleMMgSNbvTF4B6lFvp1VggzP3tBb4vhL3wKuRfLe0z7UR2MR4PlY0
aMgiD2M98tIoo5pZky0Iy1cBDN0ETUpyQVRP9a1HpiDiETHfX6nAE7F4YtT8WJbt
+LU10h8MWsRyCkcnbLj40AH4o5o9hi3WbaUFCqmpasiWqymSbluEzN4iCFdLr2Y0
pyrzrrpM58CwJAwv7CU02Px619d2vOmhs+ZuAT1xfgCQ2ZsSFniwdq3Xh8s74c1X
Y6GSRj4RDOomzFzPi5CfoV39B5g0ZAt738FYG42y5HL+aT5CYm+J3w8iuBNxxjn6
9u1KuoZKij/L4PSuZfrEorlpquWd/UKPlFwkSVzrBb+updX9tMRMZ+Vieo/BY8iu
dZLNktS2Ij8lIDmE5w4iPeTLTtlyH6p0O2GGRxdS/ap782WgRw4yfQqWn1R4HgQx
8Ib1PuVW7ZIDwJbACyv6K1kdVLPeY0arO6Sa8o0O/xUYLLcaobbQ77XEEirq9GCV
fOy6+UR0B5D3CxKWtDOKhZ8pKBjIQFLSpslUqJcxmMLhgNXKMjORf5dC20flrnMR
Ng3vJ3g/hQrogJx6wnSkwpw/ZQ+D7dHvldPZMdL3Qqe6lcZniTJnYaMhOt7/VIQ4
d1uXZA3X0X6d3GC8jzUYskOWPH59OwuQQhL0Y0mAF2/1co5SoIZb5hlEIBaW9Wk3
9A11of8F79sm+WXkjXk/B7guRnbwaQySeyiEJIW0QMBVOYJEzXqcNtVWBGCTr2gz
Yu9pGl+FbvyJubZktyT6hx/CaNdfuSwdmbLbJWEoBvr8J1Dn+3ueMBWM8iHPOJMY
Cpz/GVb6EE7KenZKDTrMJSYwfZXn3m2YKPDmY+/X1DTDlAo7oj9Bv3QCJU1cuRXV
C8gyY4EfLINk/TYb1ZywGXDEcKhEZTEGhOd7T5/+w0vFkx46EJAH69bLzb/nZeWI
4NOkLXduEC0VWq1cuziDezJWIDBscs6VYY5yAa5sqV91Q/RStRHk1FkRTbi3ypAb
JaO3JBvslHHgGYjmO2vG6//YXCG5hyEDSImLakDr1/O86p0OKtni2N4ZVxi9CVsd
qcuefkt04JfeaRllD6zGEynUZoSrzW5VOULgROt4drP2atlSSxq2suc3RKlGeTaN
i9ONYG5zrRxNEhxJ31K9maRjAVSilv5dXJXRsfmWCJsqYWM6vo3SEk8oBYNpfGSY
EIi30SWGrR84J1TD2ZPMlGuqdVx/6wJR6wBWsZZt97Q8986pwN3g9jR2N70s2qeH
J7CyUkGWI76dVV1nMogFKmH7LjckWMPU01iSgRfHmMYt6vk+r/M+YUbiHWAwMPk0
RRE90W1rYsBPgZs1aK+40ZpvNF6UsnODu87goqpLzusopSbjM7k8J/fyH9LxrgtX
MJLadLfi+szsG0MLmk7/ysmP60H+COQQzK8GgQ6sOMg/wZ3Wz+CCV3t/jq3V+aDO
a1S5/Ibg4aNPCvEJjtjTcSuVUXh2Qw/t0snIb3KfWjfaTC0WZaTdhS1U5qN2bpwm
AtcMRINnEfEt62wy81aHSQ86ww2raRuMoUm2DQ8i3QqJzXy/vEBP+OgxreANNirb
/GsLVKWuZwN0bL//9jc1g0LjIbVJ4Q7nWZA8ephzE9joCFC+7xW1ZqlZtpEN/DU2
1eCURScrZWxf77gCQ0KxGednMlSOTn51g/0FMbEGSyBp7zVeEcKeio01EFuZ9imL
42GNgc7q/S9J7L44t68sY8dw7th7AHVNMRqjeNyr5rngzTKAT30jTAJbZIRtL8SY
jZ45Ru3AFC0xdNa+ASc+B7nWdfBUGxddw73DbCC1PSQ3mHOt+PTyXZtFj5Iqrc2D
LWfUjK3YnFQ0HjQ22djnOCteib8S619IpOzltNBadQO1OGfo2FgMEDrcOySbzhuk
R7T5GHilKxCbgvaZytQp08M8pBTlTrtUkerORx+HYvpGDKnoqA3NgpjFUueIpgMb
buREdBvgS6mJI51miU8kFQAKNcykQFiHwqj0saXahUoLdPLUm3gzEl1ixMAevppg
PA/zcSPnITcvh6O5+us/76UyhuJWkRqfTZ5UFHlEGf+Zj/dUsELCH755ifp7TFsw
WGLV3lTGkL/0C2c9EyCCfic0K7C5YHWLKmuTzaDl/qKexyeFsj98JwKTrcDVFPqY
rsb4KGveGt/0uXMeKX5C740/MK8x8Rm93ROOLTH7+ElPy3uPdE+YjF8NfJlZsidw
Plf4qTLq/Oks0L0LlHsQIgWpITSuKUd9uAlJjcRg4/QnPyUfqqmdVHZ4xzLY4nIp
VMSzU1VwtkrgDge3ZF2cZG0nLYSdQr6KoEM7HOh5bam1/rcOtG3GVpMWgeFsTCyc
VLxf+RhQRt+nxDFcvkSxkDwlCFbLNotdSsMAnUCT/P9T7ZzaaA5zOKsMOwG0Uh7N
mtXVnw3276qstnwfQWvelSLTupRX39CLCegNEcpVMC15xvwWyo74AlzUlbqOfrqZ
JqeLEPq9Gku8c2hXxzE+fISHMeAjSKTWXzRDkGglGG6d3fejT7yGClJf3qH8vPr1
vbtmOiYpowd7zks/uoH/MXp8jCO3S+qIOaE48YziXCIAcHBmU7dyvJZ25ODa9Hwo
qlS/5y99NqeopaVleD+aTSJv1rbbmNZOTOztr/VHNIIe+xsneOTR8HWyQzfZezrJ
oFwyY01A11sFeP6tqPZzBWgh6TvFIjIgk4Vg2fguqtmDAZ/BynjSUacaAwaKFXcF
MIpzO4eCMneoR9Bp9RKXLf9bKzeU252UXiXfgPQybCcxddLIG6mjT8f5+27iiBQe
ugxVAwGkXCJubygC9A2cCyEZQrDJLhVHYUftAjc9htI1s29DpG56T9zM5qso7Im2
TEnYRH8DcwvMBJpmGYZSwxr+NbfwzWcjZ9imzva+aZAUx0xYr+BEcB0oa75Wt7Px
20CbYcf28gECaFIfk3IX8D3FP9lS0xswZZHq+LGEP8jmGBZecoObEGsbQ5Ig3PRq
Fwk5bKnpRXVrSwvq1LRWjaZcU3oZkrb6BOL5O5umsxjVjWKvlPvJzgJKiyNPQxru
fXYKqbCqoWfnfeH8Zks4lxuYINwCs39qBEdb1L6LynQj1myshz+DefuadTQvBtKW
ou/WIGelDp7ue2lvm4cmke0dRubu6840PVwsQdYP8UBl4H1arlbAlaCKVbccBzpy
tpDSpezU8MD0WSXW1akuLs6topfGxwdYHcDiv4w63gbHaHh8S8ytvxG8z92SqNmA
PKZbfYideVMQZ7a08n8aLzZZq01Fs8rVF5ny2yX55MQZwzuBcHvp2J5/9gLT5xbS
9UP+oINxXlJWO+QplLhK6qE5BJ43LyedHamj/K+RXEXWYF8X36Khpuj6Kee0zd9O
35/C1ajIkQ3Hpmg/3ZoOeDII44+hXXFIwoIhWjFQ4yJJLqwYk2H5DoYiAweCDAPF
FcEg8O4kr+hJgPnBy4mj4LEUqTZ2e0X8GP/c9BG4ZjTsLFNU3aGiNUvXWMVQjxKa
WU3d8rLMfxQ/XBXzzXgGsFYgOmtKeXQ+Uy2NZuH2/VOmDAHqeBaKntaH1Pbhckux
tw6DuooNl6pBk9sduPVl+e/tNmUBJkMgxMVskYB7DLFy/q+f3XMX2vipbYGHsZDH
mqaplfEkfuvjH+L313es2dLPr20Q39Ki8MzOzPwRy3GR7RUMF9xuun0THkZtrQYS
jlH6iPWFprvbCYFwOFe+GuwZd5VmzgqmD79nPmk+F8WyjWsR9V9P/f5kSAiQcsZM
X0Vr98XiDHf5eUz8fexWPjY6KYIxoVriGQo86vHJtfY21yqMQ2vnlntxVhZnnUeg
KlVi23exRVqxMqNs8AT3+jgeDnsX/3BlkmQ2A/3A3KZlD2uT+NUON3OlnFQGKugk
sCxZifZhJjIclMONSc48vqub0Zh4KF1rMfxdOvnVRR6juZpO/miubI3wQAaoL9hy
vcks1bfvP1rcOMnmGLCxX2bW3D4HRu27cHu9Ll8LWsg63uNfqT2hyjHJ1/M+Yfge
cHP8s9PRh9SYdlSmCKtdgz6dZqcuoqqw1E/9fDp4REPRS3jS98fDxv1S4tBK1SKP
Cu0X/vkBRB0OeR6W5XonEgJjX9Qv6py9ngm51arTLqtq+zvl6m7e/sihu3yI48AH
9CiINdcnKVovC4vZzYUCmZ9Q1b3rzccbhL4azny8tw4xJrNxGiBr0Y0LcykZEMkd
ogZofL39belZ8LQSGKYPNoKykDu1c2c/lt1P4AAT4nrFFaqrNxfO8KDRgZclQN5A
UMnqnAG7CvVps7RKnl0PzTRGaPSey1534CDCfGqVqNAEC0TflcH+GKIGYaTZn6/G
XjckOMG6bHrEGA0lJcDbe+IPGjZQ/afunYI5C+mQ/XfTRD2B4N9VSIpJvsiEaKFx
qOM8aWMht56ZXA8AErLuvj5nvgPBjUe0M2ltHxvwrEh1luGEmaPqRylID6tDc035
mqkqf24pPtCwDsUCA4lNQYjidLA3YrjRtMcnprCBl+L3887aV0u3/ckqhWV51u1m
HmHbowGJ6iGGYkDaSGmE+IBI1brIcj0lIrb/TkFgzJaJ7Wj6PsDvfrt8K4q8hAd6
//tzcE5UACWWxQrGTpLJ7h4DxDclc83nQexBp8TFSj0yuwrT2gUblr9Gb1C3LM6C
Mr1aDKp4gzZhegpXEQvZ5Dm7GvG11cMHse1NR3M2SVh/txkz33pFL5eDBlgrZAWP
1/rMHKYc6jlgcpeoa25cLXGOtDVMrpymjVpj8Nf1fa8GIrykS/vKmKmeSkDveKAO
IgBY43XIx5b6REhTOn/5wACpfxz9OPreKz0SmWJtcQkyH8waIC+XRxWmANkRCnYz
zU+pZm+LNKx642fbNdWYh4Q0n5ebUtDOtAN2WLCcOLFV79lvwgr/PhUjKl1hd/o3
/21WCEzW2ZYruxzKLZ/Pb9pAVs0G4N5xMihrAI7ZLQpgH0lofn0ubtkJhQ4eNbjZ
NEqjK+8JuNGXwXQ3NeMZ3KVdwlGQpAYpAiuWsNgFLVoyr7RDA0+NfFvqkG7fNnD7
U9LQcVW5AwEmXmpea2gREjbtgacYVUuurCqwQLo2CMl9VzbJHLgAikJMyXp6jEGq
YdMYeVslUkvJGnsq1hQjSdB4K6abMm0OC9TXMH3plTQW3WM6Mpv5Z1c5KRlra2b+
ydIBfQ5gljhN9SjrxOiQ6jmJUNm2D6Ccqiy97w6Knb4znpXODR5SuvJ2jIgUMRKa
wKKfIva3W2kLjAxTbC0mjlTwFljaHY6XY7U1//G0+bfpm6NtOBYwQ6Ak66pmZKs5
DPR3l9JyWW6syrzWI+ac8FayJ9DSoIDHJZ8azp4ZScNnmXL6Jwf6jGSmAa9cdKug
Mkvn2iGQOcYJgvaF31kMTAURux9UtDTFN2o0LE4VSWxy+7L+UuCo/r74LO3sRw8E
FBpjmeXVq8gBa6KxPaFjr2v1YB7IxX8RmIfni3wdlFuYAWQZrGu09Crz1WWeJSrE
QiC+i6RJgDJC1tMMXOaB3HQSu4uF49xkWutILkXdEnjDagRS5Wp+aiXGY8ttYGX/
NUZTijh3kCvB2gcKSbMRj1qQQvZR+YzaicjqUor1UlrBZtr/zFLTeyS8ydOc+rot
k5eLJwNqdthFZ7bSUshTzt/GmWIJ52r9FWmBO688qLXO91Mb1xtF7Q2Cc357tGiB
nQecpDHWbUgyCQ3xwVcF+LLg/1ASTT2dF5VY+Dnke88oof1SvyYK3SRRmcbQPVGT
QKMBQbuO/5SNkengltxgi5UwPasIXlWrdXT47EsL+0Pq/9FyE1Nj3kgJXUfbgC5X
uHsUhgZa40fyjVYsnpd5fpJKj4+z1POtiWvrQMBw6FgmEHE1/Ab9JrHtfDxkyyw+
gJ3Sbjw3beW4405qmfeTbQSD1u1oU7BfSo66E69KBi24Cw+ZZVZH6zs2Whi1+8D+
81ugobX7ioeJznoBzG9e54aimx36UCGEQL249R68Exn27+EAJuSzobCeoRLSQrhf
3L4tAVzkieRTzxyHDFuv8WPT73/SxVChEo+MIrL2C2VWh0zwftyXHg7myqcsvaN7
0JZFuSizmsiMqMBb7WwuB3PXLSZdWGk2hbSoYy50CkwriMlv0plIwYQ6Igw+ZonR
pJGXsUcONbEEUmCdlNYI20CFrZErnHAdBUKLnaQiUp84796uC1LdBWaBS5H2pqY5
4vc8Cw+lACdM6pOUAvXk641P+6NkWEqr0oj1TDltF+1c1zyGQ/YyYLxWF8c/Z/0e
QJ5bejL/83kKD+R0Nz0AaeI+s15+zCgtr65+EFXjepJmbTbrwKwqfvcHFmq8xymc
HSG4YSjgGR+wZUq/Fx2WoTld9vFXGxYNFwH2EsuMFknywtaXd3b/AXRG7tYfxy2f
HVrIWqVry+zU8X1jE8BZ/X3uDUn4jXzvJ5n0+6M0L1YS2yFZVNv7QR3VA6vlixUe
wyemmqWsiMg9aBop4GIBEJXOxbkL5oRK8HuXD4hgk5LcfRF/PjyepjAfCLBF/Oax
P5a4L2pWPAnBLyu2ImWiNGq0d9XaCuxHVeajhLAXKhbvANqu166TmRq3P7VyzJGP
48K9uJjWudgrsodm0T561ANZdldYttcDeZWglYb42yc8qpsCuZqIECuNbfu/eN7+
0MnKF7yiLAKB83lO5KfPbIB2pgOPz8um+qQjzgjtOOqVwV17H7s3oxiN6K3P/Pjg
w+Er2uINCe1bmXEnXLcZ3O/TJHmR9iaBoDoUgaOeGG8ZaCSdupBFueDnOApoQqCK
t8byzY8X2AirDbQkIu5bBYNcIieTIKjSJxhNHcP2L2ZJbsggbPKVGGL7GsIA8Guz
RvBMl4QowDRZrcUY+y9C7vy1ZsqelBLBY5htSaBYIlc3E6ed0/NYuA6HLt77xcQy
9fDbxoiCuRNfPabS8UkAO18MkMRazWcQQitv3FxzevCi4JRpcf2fcND6Lgu6N6ud
9kWsxUM32qAUx81M+ePQfpTWULAjMdi2hglKKiKU0iuHEj6DxZpqkR+bA37G5MJu
NjZpVl9/sIxnk3I5Rx65n9SCEkK+BrpxdIWi/O0pg//0hJiX+xACJWWvWFzl7XBq
yUF6AR85nIWxGhOR0Nx60jEqMY9BB+8K0sqFsOO8eZT79/r8te5dvgNUlANaW4Ww
zwxgnENwMbW1bm1N7eXGXDWkK4u1VVw4WhGrSy/MI/9LjiCL8NT6w6Nt76gp+6NT
EqmHKBJyt9uqVwtzBfGFtQZjrtL5QVoFnKL0s4iUMl/O3N/kw5SIEkmgzFUB8rvT
yoTVigJ7FxX0V37BK+87DzdCTfbWhvpg7ZrNH4u9jnC6LqN1mOYos/y9tbqY3Abv
Onp1fWDzxIVcvrNHO0IJa9mpFrkyFgml1irY667lgs4xAWwHSFvFuwipbAzJsVUU
qmcus77ChQOdAuNzwK6YLs/a+EHuzgKkg5fGNsuDne/VtmGr7uo9ebmMxOpZUW81
i+Xx5npg+qXaRvbVC5kXHWLfCujAjcFVXDRq3GpGkcSlQcm3YPu3DRWZzNjQjC6A
Mnanha8G/9vWKQxYZtEOqDMXb4ReyuUo88eEQiSm2A+P2je2S+6KId7rZzNgeVO7
tjl/Fq0GEWGqP+2Lm/U19fScQ5eDPrkovtGygnVJjkmb00yn9NcPFNuxATJ48R6H
R6ITjqfC70eb8Fx/TQJD7m5xRhAs1Hgt3nDhzWKu9xx9tvmh7SlOKsFaiQvErzpQ
o7M8td46btEQQKfZIg/5UJG2MHkXpLLGqd0Imlz+aoxfpd64gYexi08dpPV4jjMz
XsVfVJj8NEkzVlwOxhoV/7zsmKw2RLoluNkNWalCIJbSk0fDhI+ywiXUHFJ8+4CY
MI2yCIkISA3qHrxshO9uK0/wBObjwdfcBizVFDu5HjokLOgHHRMx9JdDaBwdlot0
dg4Z+MrhVwOu5kigzxUIDBhsryHQNObhsFcxgFW4nYK+WzlbnsvepsYOuAv5o/F+
w/q6WNPgksM7ih24ntspecnq7ZHQGscVnDFtqRIwR7yXjlon1bZznv4rfjVwYeLR
DEZA6cHWuIWGWYJHlpNIq0pDuLQ+Vm/MHCyy1mmunp2utZeDAFVzIwiNaxeqkX7N
w94SHS6Q0CZHBOIcIdO+PrNYwvsiRlw8Vu2Y7bNmB2orE2h1muOLkN9xQitu+JIk
U/J01Nf/I6PfVvJvzPfF6zYqvfO3XzzghE5/VGYF/dTDhebIKOjYDUNAjQ9Q+yTO
86w7Q7QQTcbEW4UOWW6Sm7rjN3t6i5l8y3fE5hojMr6CX+HWx3lMJvHRUHoNx1Mb
EOaxryA0qOC2JPxae0itF1Y95SGSIc53HFidPjTNFdjHSLTFnonk/dq4oQXo2t7i
am6lKWioJono1Z6nLpcVKKXcHPQZb0denVqLI/StSTB9dONAKEjYOpBo9o+prnLk
ANJiKlakrMxymMKVoVgRCJ7Grjd+rs6rTm+TvhWDXoXPwlJokxdLeepYV1ggQii6
XvI3n5iiu4XD/T8LmysJKDchYAbxJTCxpc2kGpEDNpXEj4Z9auob5OWZ0IdvLxM8
vRM08LJ+q3bIXfefbFNt+Z5r6CVdFsolFzb0M+pyBgPxExEr4jFIVfnVgzJCsDZL
lxownvTmDxuUzRzXxHjILK9qW8OjNxqSsjmxK8R6/gRdWvmTKcR9fHK3srUljmi1
2mziO7osc7FogHdOTDFRwoFTxi+fQfGPynld5+Z60T/Wk5RahEaTKRoPuN8+VPZe
aLmgUrG32fyNEWGoEzFAtyIj3lPwaNaxII4wCvidlTK+v5zruCeyyFMT8SWTDIWr
M7+Zh8GfVKdZLDl7FOJLbRbt+z6H7FUyINUc2qwuLMJmn4mfuM/CsQZ+aUImIyIO
v2jUOyvlEPk8LF3EhcNWcgnqk9DFsKS4u+DYjRhMavv0U8jrO2kQjkaY3DoMBu67
oXODOGSrqMOvIJ6EXxPZy1y6mHNvcbIw1RQPODsU+6VOJEpvcFLNwIKLiKn9uvVw
kWI4ekSCJWTBjXpommGETduEfIwjyWCrFLx6wgGdCPXHbrKpn34+J6laHz3QjanG
qgBN6OZhpptH9xrofs4QZP8XOPuFtboKpVDEJyWtwXKkig9uYkJSX9xwazJRv2hK
1O9zp/qKFmD4GKscRvY3PezH7xUHnO/vCwTUYoe+BCYPYWfN89ESZm4zCDpSJBY4
cXlw1sWRMA7P9yMseRF87huZGgVHadLTXjmsYANcgt2y4LdDLAQrvY9qQXwDywFz
C7rNJ5sUXiZ0xWfCceSQ2jouK70ipw0G+hIIrkWagumAelQKjxMNUq04w7xt9Gt9
mseHqkp5rv+uNoTK298sAX4XxQ43/CbSO19p0FlTVrPCafIq0xRWeK9stsN/kswx
MoLSfnM1K7h+50r0x0tzCpLtCqWX5/7lJMqzyK7BcXP6JEetHH9ob3gukSfKYUNJ
qNj1U3FFek3156LYSsaEMhqWcmwMsTDCQMLtoTF7saRgmEcYWIr9wFWXpeSYzI5/
qQLZI1NV2rnDktjWP5GytDLHX5ZXQpv5cqyj2sIL58d76DcSnclVKsgZyPfr3Yb8
Ct5dJTdTSmNKWyqmpaKMZPKpD1IQ0Xts2qe/03I90mS7k8ICDwOCgD8OkYJHPHQP
ZVNvFuJC0VrrnarmfE7NeK7uORQX3jBgwiX8v8EapQh0eng4crov3Yb39Qamtkto
M8RnoKgaI5TBXGP/1L7QgRg8kstL2O/11MNDO6eAfh6igEnHUrEX3zFfTXuMGOHA
tLnrgT0vv6Q3RKXIqMBDteGCp6cA0xV2GKM+pVR6qz5OFDEfdIZarg2Et7oQmzOJ
jEItI+KylALCemsjD9PFVZWNd6Jf8pnGDL+weylosE6MWXkM1AoJZNTMyeiXDgYw
IOPXzQOuw+9uLi0JRjs8mtoPzDxU5UcxQM3kkt8TCTIJ0oSaIRsTFDTR4Vi9YAjt
5MKU3pGCMsO2OM4KKe059i6Ay/IaCCMnzWPJ5wOpzJqWYJKiQ/F5KV14nFNyjXjl
OnTjzxY1OESpRMlUc+1FUYOSIgFYWG5mAONF32o29L+SQskKNBjv7izP6Vu11aeg
sBFy55xv9cmNrvn4AhyYfahKLPObakh4Qj4zE2dFCfSNmB95hr9+9dui5w2bX3N9
rLy5um9HdsbLI4zNMgN9IcatiowjyjnjxGNyGDcIWMWQW2E48IyXzfyVsr64yIFe
xbCiIxXWGkt4lgGJ1XXK6PAn1U5SU9gpTKMIPyIM0nJIPCRL+YKrctR41vbFG6Go
pbaxvEw3aF58h47wDWHEU3vzHbEE0JA+HZTkCPx6geC02AckzYWyFU65f5FrmVK/
xjTup7CM8FHEoJI8uqU2ZhsXorMbZ1VMrj7RWUzbqagDvSpLpT3czWNXj/nt/lkF
sQTBoSrqsc9FN48qpy/AzmvUmLeaxhJbX1PUss5/jOTV3s4wdS9hpQfDc2w/Liw/
I+1M+4LM0F0AzoBdDVOOKia6d/jvSkv2yqcqZktMkFEuAFcPGIp5EF17EWnwSwSv
EjKF+6VgknmgXBP2FlvtC7J+GHZRTUKTttfeitMOoIvjWJmqOlr2aMRuvu4o9OQR
8ueRQIAbM1laXOrGh6s8nnJwfC4VjmV1rkDzpy2Pq8C88C8bOQxH4nwWbfgBK/TZ
mWDkuVo3Ias6MTYs2FGEHh3JNVvTOVr5SJo5pqO70Qx3Psr1qAk14lmUtVKdrZvO
2f6y8sxVpXJkKaWwF2qWJ+yiKgkoWSqlQjK+fHIZwpZbbP+/+v9dWKemFrIJgPp5
85SJGwdZ66BDfDbWKGroBU4tvVIJKCxDEp0/ow5N4MB/FEHb7f+qGgp/XexhaXrz
tB9k6AkBWWMvisaZRVViWd+4+inGgmEYr3xR/WyAtpAEtfa4HOHbr7+64aMEjO37
w9+I53yawxRjGWe1JoytYMNX062eEHoJn9sn+IITXKNaHF69M8iMPoqXUt4OP81F
TNohdu/YjEUlwTf15jcX2f26F/B8Gk5scReHHUWlgVyUYwnjZ222wuRXGRm+5U/d
8bf7osnc1Bv7WlXvuAelDuolJ8hrdxFkGQdc9hufWR62qGfL29m1evSD3cOut3Fi
a93GThpJHzwoGpawIfzs6KANOISnGwgexwLSd0TzZByuPIdAlfZjEs8V3yPS7E4b
jv3HTyABzjpSsjyEHbvcIbYBjpIuq9rkmbrOtIn9hD7oc4Te5k8mQRDdkjx8uGk/
w9ZdeIG7TH4ioLCfMKR12vcdreqPN9s2Zm/3i1A6T4WziMtExHLeuR4nItkTIlUe
cWPjMs+k1/+uDlMbBA9x/rXUeRc7flaEBJn9RWLgFCXYFvRRrjDzG6OyOwxUrpP+
Siw4DjJZYhMJdI6QoNeFZXrENICGOFJN/sE//L+gbdhP6muebqM7NrFV80bzUhRB
EIFPJZmcKhXf8YQL2p7eLcs/R/JPiFc8DSYuk7kND5gs+PDMOZGJJAhFLtuo0h/v
9t5hEg4R/yvEg2jiCrx2FghSDjS/SBVdcjXRw0StNiRIidDtdVf8Z8J+mcDiqpeZ
E0uUBf1gXoLBFCMMppTFKwy1/f0jMKFKM8uZ0HZFRD1oAbr9i4jwXfNq4WnI8+OB
0mkMFVG0tmops1CFj/CjxOBFN0deUWjTEeQ0prcaMYNVgHj0EgqUR2n3UGTfgtZ9
sNgxynYlMakUOHR7Iyq8hAj0LAI+JeZFcjcZzbUyhhMF5TTuXh9dAezeB4+Dd7ak
xShZtWWX5XnLKueix2Tg8L+oh8s5O1fuRap2mC3BxNApGlbykH6ubgUDKm5q9DU1
1VNInKfb21OXqB9v369XmOLGrvHRtCifqI8v6ZxYOP/1OqZI+3kEA9KTQuHm6aPa
Ggr6bn95PUD70GZLjmNginVWOLY41sZ+94tHa5Ojl+/xyXK4kRsWPJvXSYkjWVNm
JE7N/deon8839XffCq2OvXuaKA7ft0b+9scYHzdBfo0tNefCLjH7MmJ8Llyo5t5w
RGXa4j1b6QR47Usbnxzw38AB1y8VrEp0TpBQJZ2MnFc4xQ/tTk8Xj+XgW99h1z6D
Q2fm/aDF3USahj5Nvx73hfpDOwWsh1EA2rkkKeVDavwkzHSgHlzX1s6nXXdY9C5I
RSuO7M5azEdwifTbEiVXFyG9gNg1ax7HToEcYqwtRdeJq0tvh7J02L7VIwSlX32S
O4FeHVstoHj+v1qj/9037sjrWIN+g86VgY+jmh+ms95dZr15aodhPYXK465VPB2P
WSQ+v+0GNawYDKxvRv13DLClkFxzV/OHiW3QAdfSONy+Xvl2sBjc+xdSZzcYYJiP
skvA0jEo0GvXY1M/cBsb0djwNs/Saf3mJskfJGXo5km9p8KMv76wAnywgjLZh61+
sgjxIBFHbvfG/mSoyamp6YgBgwW+Np30mw5aBF8T8yt07ss4O9l+zvy3LIWuWiZ3
DCdmoaJhO32nq6CawTlzskwB8KLh/DpY/TiHbc3QiU8GHJ1TachgoPmk4LXXwQF6
O7QIx6nW8IsUmfORTFMg005JPmRSovgXNU6TlHAvZ4i2If5iIRM5LYzrI324H+LM
cYJYjehyEtwuW++eUL1XDsrt00YFTuqQuJ9c1GMyA0V9KXCw7mXNodfVy/RX17Jb
VoOADLnSiL64df4UpBG05qwpU9iJG/rkoLe5luROl6ihVDCqOCvPJb10QWsf+RBN
QxGdjPbRFCKPVKDSBVqvrfMoBrV3YTjLEyaznCluMxlf5CW0vacu05NkRS4ss4uW
8TUoDNPfP79sJnscYGfyULEJpBHjG7AslC6s6UhYuC0NDSRviUkIwc2Z/8pXykIc
YQiAPZilSCt+25tbtDY3MBsJFxnskKKe0dX/HBF0/25MJtOJENMSAY8qHipIVe0r
hJ/hKWJqHa6gjZAMlnWyagMmCurbhk+nXdClgvI9rzjTxFvehxr2kgGVxI7T/vDN
x7p9Ot1m8AcANc1jb+xjsJ7B28iUCGFwUPWofkq0veeqfuHmbkxDrHuXivEhKuXf
9dy3ZghW0Dryebu6VJl3cVoFJrqLgSRS+YVs7ehiH2Kjl9xrlv+AfeFmkKOeCwGu
yUCDj49faioa/rSeqmv2h3a/f86+OToWpH2tuXGrDpnybDSVvRzxqwJa8+YDnD5Y
Bscs7c6+S9/VY6jPaZfcwyswJxduucJRZhbZSqqmwduT+Wi9s6TWBCBV+kUMDOzc
IhPcr4V4dIgdRYVMseffP7iMdzEuSUgmMvP6JMpIYFo2S4tMn3YrwNjhJ+8yZGuS
3ELz34mo4HcS/HFCIC8PWZuo9dLYf0XJlT/x81V++9yryo5uUdtTdUnvunOPztqp
mc+ChLmbTCMkBV0SbneU4DdajIhxbHFD/JPFtFupm9Q6MFujJPGINMW5abrGgUgi
0mfBcdqpTqGynDzXaQac3DeImCO/72tC5ciboWfmzwyr8cUk61PVecjGDjq6NMZn
aJ9GAybmBIqXqdvrORzCmqMuoRJlLZPhjg2VD312yu4BUprnOoTme+npZqkVuIL2
m6o6j+SB3tC2pfBOTfTlu/oFJUvkcdN+KJ7I//UIRge5ssCnVZrP6eeFIZFNcpzb
hpn1mWULWyJRj6BK4ovZBHcsjaALTTM3QZliHEUmWgAOpKxWGw1otPiNKnwqTgOz
u7s22Adbt7MPjiZKV1kkxF53JDH9Kp1tGhMeVu7FX5B19/avD5VaGdiaqNWtAcvp
3p5i6KxdSRPZENfZKlTDcC/31qRzwmCZh97D24sc6yaLTT1/0OleirqVLMPeInhL
r+3O+nGZH4NGSptbpLICjobT1Xls5aWhoijqxCITgx2kjKOGsEdi8TUJaq7cg77y
coZrYEkr/HLtR1F7c1k6jXkMilhb2/YP7fikTleEVvzgA+icNxOkhusSDv3gL6uR
x2n+rBV4hrF/307wdpW6Gw9MbaMTglU8KeRT54+ePc3IXepAfMvYEc4Tl8eWUksA
jY17WbD01kjZML05F56MP5lYaectavqxrEtZM3VCK6LpH2L758rybE8v6d73t1Yl
/pAClGrdfSORtu9rmxJzfrHUxOkFY+O3J+VKuJLHwXrD1G/4wyZMmfDXmKsAu0Wk
b5WgdKJDXnp/OoVchIlogbGEpPSKlj+6KprtLh0ajYk8dn3mI7ywhd+SNiReOtdi
TMvIjCO2KiNCzpWtuDxiuq3oXPwZJnvbFXikbRaLY4kN9bp62vlDrDxTQkS2uVxk
sopxTTK9Um0F7xWlDkMjA/Augg91tsdGTOVMuZhJ1YBVQ6McVPewPjpbuxnMFneo
zBMe187iaqEQrPubc9QTO6D4t9O8cKcxWFnqTwM1rDQVu9TUux0zY21FOykmEEiG
lgJeRw3O1wClmAtqufqy23A00XPiamV6xSj2eFhslX0WDKMb6p13qsp5AKHE5RAD
eDu+tLiX/tWbHgr6sLq1XtjbwuZx24SaIdWZFqBUkdwN1YATMajcJMiHw7KASLrb
ASyEGmuOnhwRGt7D+K5PgcMOf/7E4Fe+CiyX0+QziuhbjHrzUJHvLrwzSixbnp1U
6ERlxUSxXw6bWCcSia9wVS0WiJPI/QRavgollSjrizUeZA1qb5DNqZWLF8Qn2egb
UyRRe9j2QtrMNvzG0H24pZv5+HUx0J5fDd7Wnrm+GukauxOIazCJLoyyVPNkkSJY
FLT6ME3ufZ5uX53jQApBejH9nggt7tF98M9yb1Bg4fTB1Cb7gTJ8rbKi7CzODppo
py1dMD3021ni8hmbGvvzKCH+4E3VN5124giHGcguAgBQKDomvKSCsg5ky3DJyu4y
s4AqBYv8GnI46aumiWJ69yUQneUlf1pGTB4AxXfa+EnOd89wY2qLv15XusN4KK2e
mTYid3+jK0RyliDXWf102dXxMBfkjWvrEqunFYR8SEEHXe8XKCMKgCNHcb+8nPlJ
u34bpjv3JPnkaL3SC5KfXrBm539J5FRjO1ZeVZxJ432gX2Kr2PUUYq6cm2dach+y
F17lMV/JpU/tY676ZHhJkwATga3d/yxYe/hV9BAoyMxRR1G7yAWCQSr0Ei5t9BQy
zUASyjqdmPgqFU+6D/qWsg9ryeagj9OKKCF4QMBcnBi8irPcB+i/tfkTdObdNPqc
1oI4ZrERPq5/wFHdADRxAWBOgHFAHzwxAAZlU1021dko3QHctW3EbLEnbVD5UB4/
r5Z/SdMobmOi383R7LivvDy4HOxitXF3B5wiOjXDTa+EdssKc+bp6OtN6wvlG5Iy
HcAA612r8prb8G7EWqmrEcLKPFieSJSyvk7yfmaJtnfHY2LfIo+QWziYeJ0+tFcy
hc05g7qODVDNeUHU+LenZikUWDetMyVfoIdJvldy+O0/NztDOy9AB5gA2XuLjLpn
BUBybL62BDr+7aFN6LxQYUWiD0R5oKvvl/ih3FhGENg7CSyTNQiPMobd+OZlDL5+
2D+Tm6VBKnx/cVEmZmYSxAmWgMFm8BDQbZrA2z/KsiqBIrL5TZq7U0fVqHX+nD/A
pl0KMvy9mx14SVUAL8Mtb6Plj3GRyUrvD7UO9+K7kUtoT3KtKlR2Yq9O2bnMh0i0
xbJKmNfuhUHoA8EGgnS6BdJE25bE8xVS7LRLQpO5zpt5BZETE0D1wnqo3nIPUukx
5S7waZES9zt9bCXlRRmH9n4Iuj/sc8Exk2ixC9TkLrIQoyzsVo9WpADsxg6ja0o4
/GwAoKAzknFR55H7G1V78BOL9WGm44PmU7I0LTJqGL6J/GYg/4gg4RmfSCB57i3Y
v4P93msZLRrQ7EZ5sIMfVIw6pYMwBn1Bqc8i5LIcWCwDE6RXypu6gzj//iPjEPCP
sU2dP4x9EyLjXnpXtB/GkvDhRvAt9KdR6o3xwOJdYTEi7RsAEOPMQvmicCGDykWc
/JLbsYKD+I1yxd1886ZlV9iThOsGqDDOETP+nS1BojC5xmZYxsOqQdfzZJFufsHm
EtLv+J1425WQ+UVAFxJ9qvXfm19vObmhIGUqhZaeKB9z7ah5+1/o9TbiZwA0YfEf
l6ucVlpjeS/FPni1+lZGccdyAN4xRfa0D4Qw4HV39lIB24LCaiNu5ztHjIilgYIf
37YWehp7pwLKzZeIdEPlM8xFoEb84kBFUJ+Cu2XXcvA1rPPxf/Pogj/MrU0++Dai
TWoo2FBJukWQVIGRPD2GhSEAuNUdWfBzilxWMC2ponTg4mRTYfP7ZudIoAs+zwBX
6EX9fQchdJDkAt26I+TjuAxhIXK2znGDevSx5P/4BPOMBgKBO5ohuZQ4YOa89mWV
LVr2a7vANV0b5icNNQCPsyOQUWa+oWiTz/D0uG0GRA/XLHQvn9p+Iz5ZI2DqlY7o
QW73stEqYACnfkRVidS+fXktGwBu6s14L3AFMgD4XlUcb5Y5sjidRrDs7jxat7QM
8bhdXKqwI60OeoWVK+3ajrmkB1WMT3hM8u3onQjze1JmErF9exhAYb2q4tvB57aM
cQVrRwzvsJtW2llRrD5ChF0RcaclymEiUj4ZUMJrcv4i4dopNAIJUhq+t01hPTgn
MLCcyIg0PxpuZ0P3wWnC+daBLIjL8nUUNyU5D13gMXmogG3j9G5EqB4dKUKzRFEC
IfVl2Gd84Jn738K0FHTgpVnRC+rEyVKWBFnE7IJbGpYjumyP9JyxXvDPc2ysuoIr
49/y30dqUoEcitGqOV29uEjMaK9R+8jDK3+ileiar++Y4duYkZyJMLt1n6pghhFr
qZzxrw6sKnPLvAXLz8Sh76FYXmtSmHbBCWjsqoNBMBImbwXDAmRmjZ8zQzVi354a
zXFjhV4jszJxQxB9frxzB5IZtccE7+f+aQnDzSmjB8xNraxjMirxk9fPs+GjyHaf
UR70nB1dWJd7w6HODeyOQPvutzKhDfgUJKp5Xm3B1foNXztejBOD1DBWj9mnUN3u
wNOAZCwOubdoKH+tMCvk7wYOHH4XsC23CHoAQPI43U5cf06gocu+Si7J+zNlc7Qi
S3IXYOdglVYHuJauaOgazIV0H20tIQ6+bu4RlsJPU01XjzhihAwnedyxY0QPpvO2
I7Xtbj/bg1Rj1Y5HpUuZHcxpwL4QbTm8VR/ZexnMUWz7lMxgDYhv6B40jczOJ4xx
yIMVhyPqmN3SsF1PB2hZ4/cxzESsyACVlGD+rB0ifvZiWFjfB2LA0Q/lHEQuY93x
IzGUCMCdj0YTPtZh6Qro60Et0JxhgtZKdyT6VXfgwmopiwJtFOyp5hjgllzOSi70
2G9ObDcvGNINh2ybRq6/syKfn4G7xR4JrkmjrClVGhQ292uQ9sVf9dypdIV89Qbn
tHj6/BM/1EbVUKvclUMngcNovHutzQd4nYr+rMr5fHTuuakVAbHF/CzH/QbgPAsb
+tfgkMYh9swuseoqbyQVDgEOtcJhenv/0pG8bQ8xb3BmvonPUUM+1+e2a5lBI0YF
gCHH4WgMBc+80Kvb7ybo6QS6u+cUnwGM31ZqYipZtApe5FA5vv/+1dkgypxQCh5Q
f1eAcuLB0zCPN3kyJ3J4sPsDu5lz7fHXMbLo29giUuCZQ4z8O/zupY/AR2Yt5pHj
VUlfjI8mzKbIJPxecrYa9Yqw/bwn3EgzNGYE30KNCszcDj1FhLtD3CP4M55RjIxK
Hu++CsP+Q0jMSHGGNcv3Wpm7glAm/NrXdgnII7+2a/+WGWwoxgoJEv9x8BzL26qf
UuDuzLUWgIDWPMXJ+0utyaDuBZ1bMWsO63rZbv1XhW63xSR5OhMMS0yKzvUTx8cW
QkneVvpsa28ZQnARDCyinsID0ZegZiWgmCrdlKzSiBkh2MaDpbS79ShNMOAJjB4E
GZcbtNfo8JDOIvi6//QejnluzXzit4xnqVXLaJhpZWwZWC/TeQVjLNqLiPAQmHXC
khBQCA9TfLASIKHIH50wnATZMavmhqfv83xlCd5caLo6ljjkOIypjcjdeNZJDwPt
oStAhDkj7G+24WCEoOnwwgpihNgSvnzEtJk4on8j/5HacxnOAb/Y+a+Mi+RXy9mv
lMlU9Kic+3rada27wzojvcG5f4t/SCUc1lhiJxsofwsdTHAhALPwy+RMOb/H0Ou1
2/ME/YchWtuyx5NNZWILLuWiGhf7jf1TXJv3H7D+eS7abMCL0JAW3CqBH5Qi+xgD
icNATbiEKOEyFQsD48qCAfoT6g12E/4+lvYPIjiBsXc/tW/e9d4iOvAtlrWohqKO
PcMrHaYryrS7575FxTsRCTIaxUomGAM0rEAUKi5TgT0Kd1a759tzn6SkZTZkvDUf
jg7d+dHrFHn+mSulbU2elFibPSD8NaoVLX+A5QoEHmODwqhZZ4N9xPkaHjXJ55+j
pMe+7Luzp9u9ghWnerr6YRM9i3s/+74X9veGrNyJluUWzaUATvtSq26ZBneniQ0p
t1/wLpCzawpN0CIj5mf/PzNGKq0QbIVelxgg+CwImfTvQiYo8sjbnogbPTqf66dP
AavKKCPcojqUwRwHBHOcwhGuFToFOrhuppYeEzREs071O9COby0jmpaeMXcAEyPb
l2YM+P7UPKYaMIk89mEMGuE1mXzrkP5XBdUw1xkWeOH9w5wEx+vVvOFE0hdSi0Bk
3dEuHzrrC7ugypmqIVY9g4Hr1RtfK+MwEJi2KSIA+G5P3T/6Or4J/vlKJJ/fIlFM
tRJLNbrJ5cX+8QJvGcSF4Nx5becKS8XHBPDUcOuNpn/WCiaNDkeZnAJ9kTevS0Ar
klGRhyh/sHzVe8rfEVmes8ypnRIg0UAB7J1U7zqtiTcz/vfC/hgbNP0+BrKVph+5
zbt3EfMMIYfZGO/aM6gjZOUxa8WekctIjl8pN3UUnkon8N/vDhI7bcGZjeuoBvdF
M1eBsHr86z9oS+3dWgOK7w+2/vFAjoyKcS61qSjjQqsoRyhKfZdhRqD1uaSA9bH7
za7uMlgZHUB5fOjCX3CY5BqJy82Ug/AgzNz5Gd+zjjw9C9LJ4/yg3icPszZr8koO
/4S72X4VEPFUMfdTmutCYtwZf4duiq3ICt5V3vaO7HrsA08ubq9FGvIHYw55/3TS
f+uW9+nCYAVpuZbrO1FLrmEVIZCJFEfMs7ZqPS5x0Hxbz1fGxldZUBRoZSf7Arz7
1UbGX0X7Zoful5kfNbOOV2n2vHRYlmjfXqplWpwiRLSP1Q6pRWKT4lzOa8adcV7e
laeAm4RbBMRZDx8PHzb1HJpwZXD6iKP/Ot4MUihgZhrIggVyAhfDwp0LqAbGN0Ss
dQ0vmphJ/eLg0C62lLQ3awdVGZMJfadiqsoFAeKumrQG3TT1jziESxmvVnnZW5yt
IfZmHibvYDiE7VYzxWaLZz4+XHpFjjDCG+KlQur81GqDQSaJn4y9db1p9NKQUM/s
Ik2ehKUDo/0VztmNSIsgSiPqAxMJRS8YGVRjLnPHITJ3Nh5SOj8eJJF6fqusWqyw
/yMI463iWFSyj9WWL2Wc0fuMhpldxgY4thOn2SOifKSiUdoiuvC/koju4yyDwG4f
AE0Kix/nqQsq5+X257yocSzcqcx9nrqSaPMipmPaRHO0ksI2ZebUPB13PXzWGrnC
yimYn4/MkNqCxndd1h6OPAWZdgxam77uCeoBCvdCKbPuvduWv9lEhFlGuWMaLN5y
ZFCgZ8UeHWHvaIrDCvDiKnVSrOW6r/W0UJRhAAOOq349dohwvArIs9l8gRm7m4fa
oIjOxm3TxSPjkm0dt597QorHEksaWmGYjP77A9ibtTRWGbml0jnUOPkUqgPPXuGp
3+4VkQ+3+6hjLsYbSiZ4laz70NNcoOHOM6cObVVDYFGSkLi6zYyjzOVMSyTP7Nf6
4LSIdi1C6hyGMj6p1ls1JfG7ALcOmdbI/eaLr4/wFXjhsrqLC/e6NGx4msaC78Zm
W83wMZF7ToiwqLgtTmg3WWYrL3mZtH5qA9ODr/ijh2MP2jHhS7r9VNvZGnPxVuvJ
TTHTJ9BTwbQlIgfX1S2nr7so32Zpsffx2yFLXWf4JYD7BgD1ifNcCQi6JX4ZJzUD
vd7sR1aLrW3yW40cF38AwW+t2Pz1IDeuO+jX28Qgkf7STWcPuuVZnjCy0R23tLlw
yZjixU9tEUn2VbkTZ2CAN06R4kPa5yAskX7+Q2GSMi4xC9TVdFU0MeOdAkPcnMYF
vFxGUX/Y5C3k5BPviiqDHJGLv2zBsPoWy0fEvHMrg0kbTtC8yFUygD44Q2YkgTUR
HsnmMugvuzyeiAwNeP4VU40xfGmZBGt5zhCBc5eBkIYJH9DHnzQvfp3VtdpjcAV6
G/RW534xEBQQsdekl3KIAJzQGA3FSGspLWhV+4UiAAaqu1ASmNeDI19baGwiS/zi
Pc1gM1DgjlGxsv0pRs2/Y8TR8wAoK3SDqeUm7wnVnDPTkJEGQasrLJshDgTYLq7y
jBBV75yIsK2xzbTpQtjdUrW/j2cjYNZH5+cnh5Lt4OIxsX+9tizGTBu3SruvQLtm
vJoKxFoWeSeKWaxhtne0Alei3/EEg2WaH61PApUiExbRSOd7BmNeqouj5yO8d7PQ
LOcxbRTOFUyoWyuxFrLJ1nMAlQW5syTAS7R+xIaHJ8KAfqbMTmKkq/vsZwuw4FL6
fczcKLFKF6Q+deRx7FkUC2K30hm1xS+HkmFyJOiGQ0hI52sDmEJLEVOYnC8JoRAG
iJAvCreN9gRlMyB50NQ+xJdt86ueU9O1gQyTU1yDjUDHXiAz63mn9dTY6XX2KGNs
vB3Y6rb2W6maORBF1tQMIMOLJntrGIwtRvnn+o3EpwHcJkkPnWy8UaDdD5egRB9D
22kiCnJG1S4IR3z6LqO4wUFmOZ/vZDq3DX70Qf8Cd/VpoCcfddwTzbW5rh7gu4gC
S7A5AhCQz/OvAukncVii8NIq5NCo1kXSSOyhAU7hNLH+vVAbuae81ptSJc5qqLLU
5jN63bNFt3lR7dP8FABVYZ/VThJTkq/9Bi9UYUscrTAudwDyYtWDOaMjjaapD8Ib
P8Ahnk4W6PqMiuDWZnq3sQGRsG7GhOr5crEKLrxYPTR2QTECvb4JsIDfXUsH8/H9
FfNURUKuW2KOGQaMtQxGJRYEofHFAsd95mjKgIBp/kqy05vDGyHoVvHF935GfkVB
SSdc2T/3yKt2pMOzBftpV3ZNY9lvbEl4B3waz2ZUaGhG2s3pzn7Ym72fd/XPE63H
W82EtKwhr+b5XMrF1fhTB3oufHtmn3aTIYy/kWN/796oRw7NrOlfmLyz7y/cKbwl
3BrjSY7Q7++JdlTvx34bDcvSVxsFZuTDFeAVaAUVaZ8zb85jdLlLTv1CoLbmbdlo
EFtTgRJi0ooxvWgHZCtdOFiHI2sZt6kEhUsBxDYp+1xBrYhrnJA5Xz7KJMVAzBKY
iRhei3MRljaTh2lQ1c9hHwF31/eorkScFcOA4WDkacv9uaWmIS6fFlKt776KQ5FZ
EKOqIUctI7Xg9h9KHWGk6i3b6KHCk/uGDBcg9xmwpfNOA1B3Bj9JfxaQQgxtLb8K
KxOGMgTAXARLL2eSBv1GW9xO31JXR2gacX/imhFBnPcY2h6vzxiHna6wkfDK7AR/
XzJCsWmDDd+jKiU2j/DRV0GJLvpe2bg6MHEyqD7BfenltCJoVpaPDHuHlyahx2bq
KE5j1ga5Sv6/IQ/JpBdWLf3zs/hruHESDHe7gsmM2zkEJUYIBh5vu5BMhU8kuLwM
Sd7CY7vnLXyzAJEH7c6Oiwh+owHGwhko2yLG35Y1f8VqEpidWSub7gkdyVNi7emB
uFroHMwub1ad65tQoS2xU219/O5nbFJb/DW3kfCtXv7jRwwKcShZP6iD96itPcmS
ZlZFbji++h5sGhDu0VY01UHSoXwEZ86RtZQZxK0/yVHs2pvAQKzFH+zPDw5WXm/v
EmJLwq3MzDwaqwjdxvQp07CGGJ1HYVFYfWZ3DLljA0tjWsTual00uPZP8Za4foYr
lw9j+6q77vtaC/0S+POx3fm7qcKya/3nWCzk8fm+zuO4uOpo5ngiI6sfoBZ9Mlpa
+s9YsOy+3IeI+19xldEZg/17FjWXM4yJ5pDmdImHM9tVlSKYkzzvFRW+Sr7TLuD4
P7FAfmtyT7H26J7JAW05jdH/AethAGnj7cqn86b/KR1uSYsSXbeagNLBLx7DgiR1
84L5WQqwnpothloPwt92wCHoMFf2jZSuXrmdw7A8Gve9NDpC9+mvw8ZhqRNw+2di
SzD24R01MWrZ+irMMzJv/Ukih4eOAE2kUlkjnCW46KFR4lhpRxiBmcKRm0zgopPK
Zpa4RZHxv5dcUpzpvQX11YQVspkY7WOU80++MCkQlP1VUqzhq2d6rxf+fLETSWQ8
mMyQ4UZk6HIVHztB4xtY8Zu5G5gUDHGo153uZcH1aisvypjdEt/yOQEZ5kvxPRPV
gJrya4IXyPYBTIzNax4n9DdsZiCvKBfJDEAstUo5bRN2Qxdc4gHxcP8lrlmjw35g
H0Xw4h2QRPRHXGMbfZTiL3ckl0rZlLGx2w4TFyUfog0hXnZA98OvnXL9wxBYxYry
A5sqvxyMxXtdQMcDu8h+fJk2/XiWu39gj3eTTIZj8AcFRMu0xWRkeQsQ3QvGTBBV
MS7JJns1n9KnsmqAlvbS7VeJggnq5r0qaUQ/7jomwm98tnk9uXCnGFV7uyIqbBMk
PV3UDus8KDjizh0DDn1E9dEN/JvmhU1nyCQgF5bbCryCGH1CYizyaRs9RYvaqBpD
sht4Mcf9Pr6zcNUUZk4zFX9hLSbWayRhxV8rK396SJ+9V0U0bmfWxDORazFX0SgP
r6jrGyZG1eLBxMGlOfgrtpabkOqqLEy/ZCwuHa1J6Sm3kF4Qhsm3Nzv56QZ8/cDk
qBePJwjMyGJDNvTAa4xHfNa/yNgjamFH92WJyRoFZvlTUuQNTMqxJRpwY9p01OQl
M7mlW8nGl1LHX1bhJykTDyyIHyIUtlG2MjCsM0dBlhzJsKU06vuXYclgDJBlegHy
HJsIYk0hJMHMpyTKqBjNpIBhKkpAtPQ9xCJ96QwnLcTxMQZ1lPsxPQ1gzaN3xnIU
CeDDYbF6YSpKs8yJVAtHeQzY04jD4lIaKxdG0YQm5qXqb9aHqy8ZZzAar+tf7FJO
4jp0C9rp2iNaK5V5CWUYhyGQ3zeSe8kfVI9qzSH8XGBo3ocPpePLDfJcwMdocs02
xIj5Bldd7eCKevOd3qlHJ4T2YLNO4skKbetKAXZ+slHl/hBVQRwiuOMayrX4gNnu
bLddQpS3Se0ERcl46Mycfj4hNxCfCHgXBe1MNoaOW8BM5aGoy7w7aOdOy7yRs5ob
dEGn6RCzo6MulkvJDWZBYD56+Y8GqiyCvTf8hDQ82NQOVMfNJitjeMcu2W0OHU9j
FYAbVxZam9hS4vfagBFJVrTScSJ2dvTGrbkGccNbJADwmM+CbuugQ+wo02FNEzts
3lcdtmBGBxdplIid66YC+40JHGdZBmT4ZCKa+JKu/QGma+YCUgumrk2FHWcfHA+R
ZrCueRGAurQtKTortlxQb5I+jhqpnsZjXASlfFA+cgPm+sNA5881BM/b7i4smvj2
iuc0T5aB0AYqHmaoM0PagKuK/MTk9Co4jMIB+vG5xW6XJcX9f7LLBcgEe+X3I4cY
fRmRw4oaxrE3Exs44sDoGTN5xjVo553W9qDuTkb50liUle7Ha0UYzqpiTcUuKKoj
Q+HXqdMx/5w9xIalAym498z7aeX2LVVk1nYUOYTT5au5O1vybd+o91/ZYhY7f340
X5QCZ4bECHdfiOgei908XBRI4Nz5bl7A6Vmt8pWy660hW3RDytyonpP5iVZooC46
cZ4QtKoM+MiGTBoMDxpc1YZoQ3Sg9I1OGYRtCiHiJqX7gxRXyd55BeBZzbtUHvEh
HMEV7LjDuQfIlpGfKuRLv/ah/s0x3m1Y8lMPNTZpxkgcFjcfLTrgwLDL81hgTu1N
wF9ucn6xf9AQuWcdBoqouUdSInx8PnEWSelXyyTP1cau39nccDTF/IQFx3q/o3V7
u3/hkekSotk0FnE0UVIob8dkSy/DPEyUJp9S1WvJ1HlbpzcFltlmJ7yAE0LBI78Z
LcEdqrPGhnlxKt87SMeXDKpU6qBN/3qZ5g25IFoYAJBSt2KS2lKO2Bld/vLPqX71
0MJIZWFbY2I3vEXjRi8xSkpgj//+dAncssf5QowBhoM9roBpdvSzJYLneWOF3cUs
DRK83H0VImY6g40zgZQZgtr+k2AZ4+imd9Bj1HZ7d09ECz/p9q3Q2jq/z3hVKgDx
F289r1hoevTL7Yq+VFOr0SlBpl4LwmHywFzE1FVDoUWW/bFn3lAsImFcC5BSW3Ht
K8XTaNiuWvLUWxtEgJLhMKnKPoh9/7GBhoYkpaRMh8eF4C86ktjby7R96Ba/v0SL
oyu1ynOuMJpc5EZTswNsUghcVYUsTlQDvoBm+maL7U6PtaeLWzoc6x/B8E9u4mGE
ODT9DuNlDW17EJC4vOC8VgTEc6ZnURohacwOveeQ50Ph7bNfTumvMw4AlELlrmox
nqKUzMtMVjJQTuWGxv1iPDGSZn+/Fc9ApQ+zskdGi4gC28L+Rpf9vuAcpG+RzKa8
llm0sp/EsDjJ7rOAwZwVcBmP1bSzQVwHCpm2NPPL3alH2dL0FWjqaudQkcMHYltR
wGL0CPxPsvfx2TIKLGF3VT0DnIHuURvfL5cEJdELOlikHLfqt/ARFOwL/h44Mv/Y
hCKoYHUg0qq7cjaZatrDZnS3+bdsIlpNcah9HZwhfvOOFAf+ZGmkB8L2PrtLY8uj
suhh0FkJYO+f1RUj/J41f+MwKkiEN0Clb/KSl5ZbdeR06dh4TR8viI3p0BtZ2crm
Q9n+DZliLVYPPVXjseuphB62zPBoshYjzEweoTKyNXbBWS88RphUR2+Pvh3EIEGx
rZaGoqLSQX30KFuFX5qJtLIWdCvtfDCAoz7TELnSC6G6BzyANcNjejz6p0krfGPY
qNbDds6xCP0L//UwIgr0mM20sYIyeKe5O4senIzwmODzTiZBShlE3aHXGphHPpdr
Csu9bB3nCOO7UvcnPvDPEYNCS4Mpf8/uXMCH8FfQuBa8rtdjCieS/vgXCLL9F1+A
U1WMd1U/nnT3zcocYFsD0yBjGSJM6VP1ksdWXSsHM6vNRdsxVpKrr61n4fIt20of
36JHBY7AnY9bdIoo+KAK5rzEWYwcEn2HYJldfOjMRt8KTMnLC7eSfFVp8REYWsdW
yNbUQJqK+VD/RtZi+c9GSx97GsaCHs41JFK6dSMSsLxltZ1MT1xwdjz7buFAnBUz
CAEM0+qtRWufR/k8hbLLku4P4UhilIdd6TyNGyt0A2JJyUzQh83lp3uJCIqnEcbW
VkpAPRSSsaPH18jynHkbGxOiu2ThJEWFRA7MOUBRFfvXgHETJnP/jO1XpTWYz2XD
0d8S+cQRFzQGDx0BzV4+bKXpxXh4Mo+1ezrs/2cjqF3WGDVeyFxXcphqjvCNsAAa
UEdFXqgpqXeDmAG/xMTREm05jd/ri93oILy89T5WqS3AC5nE5k6/Te7Y9YSbm42t
1O/SLR1tB00s2d8hFSnlEGxkYJ8rJvcTsBh05wx2Z6Cl++1PfAxNtSn8Z/r/SdTr
l48vIk9Z4d/yVntqgNliWsQPO0vQ3Kex+kq4Ibe+miIXwaKn7TQGaxBxc6aCXfen
/dcxM8koTD7ivdbHR7QJbxbj/DFtxwK/NCcA9+nPOL5QxZ2vPF8wSI5AIG75Nb5w
4cjFBMAC9QGyzoxoHEL8GDQc4koCIduH48JEZscoZG4oCFShJwllscKo/QkMEMPB
D0i/Q/InK60vgU5RaPwCuSM5i2ELSJtZ07KXU2G8iut1tuBmsfnonzDYBC8W4G8K
gXVOszRoWh6CSmOW1tKD57FHOHUVHqq6KpoQ4qlRNPMkSlPZ13VJWG3pOk60Amid
LPs/6L+DxIajgds/xhHdABov/f0rgCs8TVQo63ocLIvIwufFqEBMXuE3KzHJnnWa
OTBHa66Jo+9rOhyKsBoZZRpniEGwt0V7hMZTICzqMT8QQOYnKCQ2LTxGGWwrReSl
VQvDWChZmHtuUwa00fJwLIm8Pe+GXWnIGf4RbtT5Xd8rQAWzAdJaR37x8MCt6ksZ
I4hkEbvqNd/rh+nOGhfGGNial51I0mxBZzOi6dwdHJwmjmk3YndDgU3U/y5kvM1b
EklV+884XH1tIzqI7c6qLcRP/mn6UNF+UNfAdPa98V2MdVsgKtbHMDmE5hPw+Tuq
S1x7UTXigv3Z+yK2SFleatpq2bJFExCZ5ArPszEwhdoMgHK0vnQw4yelP6acN6qb
HiZxT03yyAb14GuqeAWoy20h7a+PI1PYNnf+sk8gFm2qRT/S4QnOF6ceL387UAEs
wkf+Zg+P0+TSo1v4vr1lsZyJIOQCVsLhSGyhQTSFWCfJYjNeFAezNhd4Y+TgYBuC
Z54jbgFUNyw3s0sAq0OmIz7xSgE3l4WhxIyq7DgrD0lZcBNULdYXl//xc4Kl75d+
C2Cyv8lHT2gq3JBfgBjzxFGrUsmgRYvUO/C5EvaNQ6582ZuGRGPZn1dvw2NaanlX
nhUwDzJlxW34fbS89iyF/TM/L4fhyI1sUHkem+6TK9S4A63DPrbiKvS6IB2HcFSe
rtWtrbLWSbCDNUflZ71/CONj9jhvuQ4wC7rTBhRsnL8Uu4TUrVVrfUgAIyDgLbfE
O0NQRgQQ1gXaKgtN+gFUBh4Y/fsV23tf8qk9Y0NxV3jlV5Fmg/Mzz1nXISvF0GFO
WHni51upof7bhBMSq06p/ljk8fpOQvT0Uldm+ANGKqkV5vEpdYoOVt39ac+NbxWE
d/pnixRIhfBz6B1P6HMurw0NitHnl597oG+T7ybOcf3K0ednM6872S5a4lUH3xyY
wjYYg+FVK5xmJAV4flgpaaDLqJhYt1qL6LG6TgRWjhNmYZVc5U3BfMU4LhiPWoI/
EcevIdd3ht//PY2LVoE/4tNaN7bzOxFUXZ+18x+h0u7wLVh8FmH7AgzoHRvIhSQG
GE53/WdA4dSCK+c/R0uYZn0pe14e32jPU/IUUm8bhjXypl10GqFGKYs2kCzv+lqj
Ai4MhP5mm1ZARuHU1yYqUDm0mCntwLpP2JIcOAlh0MY324KWlyHitbrRDr4EpWzl
XC5D43vJyuV5tAAzASvUmTLDtCwyJ6JascNBiZnEcjAjua8+R9ho50v3X6DBK1B9
sx9EVD2iv1bDDCak64kykjt8D+SuHffR6NmwgF08I4YhrezGSVFWfDXYIiPP+/2C
zPwLqrScIwQuEWOX6VoYYs+rZ1wHUf+sF6SoyjhlNiuJQibTNf4X4+nI6kDmJJVy
zMQj2KM4xsT57rguZV5BTUUmSPqFGnvsXcVehZqYN8xGm9U19OAmxPMMFioA5NrR
CyQT9J7zM6x+weTccHWjyJ6/UqSUEgSDpm9ko8Ni7RhMpBtF1n4CbmL0Icx+h/4k
TVrAnMqBJZ988hV3N6ycmx0a0R8Lm6wf614uP/PKO97GPRtJcmDFO5AApqWaY4Af
kqOt6RohJVDskYU713ITV8phCAOzqp1Rrt3riehUaAopBOXz8qdfvKgkYd8aRSVW
va5YGd7lPYk/X1SLGzbgQYeWq9zxrKUH8FlBqhEzt1irUEuTDssGE1gbEYTy/aie
YWxcS+jWJ7q/jPaJ/SCvDzu1Tt3eR8c8cLz7Z27HsJCmc5asJRkJxP0l50+LSc6R
8rJqlJJlQuBEKKQDio9/ql7KnDXkPLUo/UEipVAadQBvDZufiC/AM7LW6Urc94dR
C1A8qmB+vVE3C4CSIcG5faJnXOoL3f2vKIqR5xpdQzsmBbh7FNKLpOGagHzyrwM9
f4Z1hxFdeJCUC3VECiE55l1PsRnUetnZFcsB5jvPjD71wajNIxyQFo+ckORsj9tT
LtmlSSM/6FY64VXrIFeooxch0kIehCFjdLeCreIySMtarqLpmcQ4PW86EiGsRd5l
Pv87DcQId4ntMyJogw3b1dmBkcfAd1D4ybbBOA19CsSgfb2JGEuZo2tA4rKYoL1G
YHDsB/qhWXNwKX3BLnA11VbQN2DK5PN3YgaMIq9VRk1w7jKwVIqbneJOjbcFWGg4
nTg7DJ0iTk6ODdupQpQ0RwsTqCMeoRwGQykidj8TrXADa6WM33va2lsYlZjpfnOP
sZyvYfUan3y7uK0JiWXl201GeFfQ//BjSnjiyVY1mMk/W062AmodCipniPGIL4/V
ql3Fe+8y9jxeFUWh+CknIo81ry+sDo2XMtVFoMOmU444XxIlmymlg1quY1H8Jaav
7IjbxrkugcUPAagEyxGSUBLuuyIviGDbhLt9rFhV6Do7cUBYgX2ULcYdEkSw7RIY
rA2u7evRT9TIjW0G8yIhZl1pXheFtTookvlast/eRQ3aGJVFHvpgplJ9QT15RuPc
tkL1dqfs1kLhA/6bhrxEij+PXMvQvCH1/K7+sflul0GUeSucjo9595/+l9qgc8Xr
g7VckDulYbmRdArRjFzocbBBjY1OZR08ti/ANKqcwOOXphxaKKnUVbk8lOQ/Akzz
CeUXvrYl4hnAasO7E4BrvmqgXtpllBQHYrZnInBmSrhfgYGeySFcN2yvprUW7sft
AnP6wVs4P88lRolK+Z8/OpgmPzyR1R4prq6/6nwzVWwUycmNxmODykZ7nYbIcu46
Vmw6ci2DVgSRcFJFyzKYu+YAjVlfr+wXx3lYjaisAF1wSOdy5Lqd4Q375DLBj5Xy
Xagfclytc02N76UCKJoo8jgs520bXMWC/3Uqh4SHZ0SD4/sj7/gOQJNj60kTEmyD
M4PUdZ7TLGRYy4pfYFZe/tQ1U23sUQW5t2leBYoNYbsN6NM73rRJy+PDRWTmyJ4w
fHI/cXNcYpCbIDAdH7ILUygKZwXmlG94NZm0LgwIQx3kdZgH2ih7rUaywS7RnuVy
aDZVibak+0G5Iv7W1ahwJ/qtB0iJ3dN9iLcru7Jxvo9ojHH29UDEkErgewdy54Mw
FqpXa+MNtEkIay4374GhcxVg1ryeBBqdD/QWdvfZfzj67gzuawsmv41FuFJFbpjr
xZDPrC7BB0Cz7Hr8SLqdGCAJMOke/m8WRTi7La1Ap/N8liktSO70YiEpH8fpUNJo
g2rlLm9wGTe9ABzvqW7yxtwJbezVIfMUFGVTtGLXhNyrMA6B95SpRkoigcDfSPqy
R7tSTywmtXAFzbF5GfYev/sdHVbsiC17Yf+I/H2ZZiGO6aP8ZLQA56I9hYMqtyLs
5J1iMIkd1MrQzr31rVQSmb+HTRyLld9F/kmCeFq457trk1G4P53WRptQJu1eWiYi
sgr35BbTfmFwa76EfPevW7g7qU9F16pKai0RzHRSluea6eoWzjf7+1qB1ht1xmWj
+tK6FUjyDdLAJUHFfgjTnpYC1XuPg392rkjTMOxn9jYSSPxfbms0d2yHF2D13VD5
5/TqWz225A7ny2HRXAKvMOSUbPG7U9o5B7kjlrk8IPRhy7UUDvrFfcBA/J3GZABL
QVOrhtg5O/pHb0yO01+UJmT3OqKNUoU9Bjvvws3Yugxh9qOupLMITgWJlsf6paNi
fzYSntTR6nQy7xTaVkg8rbZnyrZ+3Ccf6lxHdAf5ZZ1R2Xf1GO8sFsvhF3FW5s8B
KLeU+Js3pFJCcZfMuAd884cwinVr93i4k1ync6YO+JTQowCm3wTcTFx+OxJNXIgi
H+vcXpxg7qQolonQGELlNZ/jicfb9ODVoM6B+3+u8U/IAcf63NbrrnKyOcbI9neZ
EuzgxAKtoZSk+DgV+Z6p+gAouArrKoUme9vnWE+rw5FzjoHMR7yfE0jBpmpmL9+N
bHGtf1Cpwl6VketyZxCE5KlFwKEthwp8eByQJIlC8U+YemBx9MoU3hgodM85gw5u
Rx7wHkRGYGXSN2n9gup902y2wPUpCnS+cFCfyEjsnuBPPl+AtjomUEAumc/uVTvg
5hEHO0ymoTE2XWdRNlBdy2CkgGEAnKRVnlF+6uxARUWp94+WGtIT/1ROnUMh/f98
t1DOZs0xdiS8kSE3KazKOtj+qVoGY7XaQPMx7HUIM8zrVfRdvuqg4VQ5hjQ0CPtX
V1sgptAXBjyrkx7ZUnxtAaC0Zd1vXLQ7LiUP7oqtPhctKsotal2g2BSV381EnI8M
oYKll727NTuDSWkb9NZljvZf35OP4w9mqMqRMtfYZitGVtd7/LH7PyKoeqktDduc
IFXAqrNKKrKW/0nkWzsi0LPGJ+18JQqWj6Kg6fnC70kB0lrT465SZX8rO8m+5L9x
HIuryp1g16nsyrqEhPDuPlU0SUnEg3S742P+jqmCfYnf6hwTZeUn0nuqlJ7kApwV
xgtA0tNbQlgCJ6XwOckfKe+YTJ90AgTRTn3FJt4Aa82W5xLKvLytbuxCLqM7oG3Z
EH9ax6BOmQTYMUCLBMlZjcV6Zedc3S13B7eU2AbP5uIN2S5GjhqPsCqHbip11ftm
izV4DDTMZe8213YpbFTDk7VffAE0mTet6zg6Ltgir0nomSH6d/qPg5rkt9KeVIMi
LHcWYDpP7ki/nUj5ktJCwSCwhgzXfJlQ4xDuSLzeRcXFNuPdFz0woJyjXuVPMNAE
xd7CTFyrV182jZnTfVc0aeUvbFTvC5FeB6t9tRlT2WcNbqNndT4iWKRnq6/GaEef
UN1/oSqfyYCfipmTseobCLhRnofBCVju+hp0H6xTPELcOfELlsTWAZtSVD4FzonV
sR8lWrGxQVeqEvZOH95+BRiW876KZ3fhaF7kcgV/yTgr10pu9ESlm5G4KNbyAW62
EFjVhI2ZvNrKnsmWclCYAQkLLvtlB/KUf6yX5G2QcZ3pHR5Ao+/bi++G9XguPZXA
h8e7KPeR0wDCa3mBg5HiIsMJhkhi8HewBim4CgAY74J1wi/zbQZBUP5BkSYlWhEq
P50uoNz8yg8m4Sw9OLK2Es9pAgMZpFOs8qqUfGrRFHAu9HhVVM/FKJCPqcfLpgf3
ZxRpDQVn5SxdP91NGc2CAfXBYbynyx8sEogcRWxUxH+fbD27p9R3+dZuOJs1wTQD
68BOuNoqARoFikBAIn6yrC0qhct1MEh1tqbKD6TlCMOreSuM4GlTQVMvRP2RL1VO
z5dds9RArJ8KdY6EQjcxpEcNkdlKJI/qZ9Leb/Ruu6Od2vau9+ka5dA9yYnsulU6
rnomeIOq83In9uf/WhvfzrFn7QSVmdV6ujd8G7re1yvTXOKFeeEFuXn3TLsR5CYR
FMUl9ZbVsnP/7Ig/02LYypLtX5akXUCq8Sk8VSBoUfodbGcbP1JP49arCbqCXPMI
Jf79pjox05IXgs4wm/TUE8/nk+N3JffNom55ZQWOth8jnBtzgOjVAV30BLjbWDtb
ZSZJavRCVpy1KtkVuDy4t5gIRuxF6qeSBUSybIu4kPeyPPU+5HGCHedxTButl4zV
2qKb9qmGUwF1p9R9oenObiJ1tqMPGzUz4GzcZwnvUeh0d1N7ypgBGIyqQ5l+myIt
Tbxs2LptckzjJO5YnUc2ZXOy9F5ybC8yLUZvude54g37b80ILnliD2EhSubz0M7M
yuoFxBqZh7PpLXbMK8xcLC1O33GthERoA+mNUCczjjqiao7SUEhRo7wkk0Jg0tnE
imbk6q2+69/tmZbk89i4V0I+92sNy6fMwoeH5O0c1iUURjm3DsaqpLGbKZSO6zRL
l9jG0XViyLiJYbIMtNj+rcxM354XtgTZQGTEqTgtW8+Hlq6jJoAMJhxmiUErZYXL
iKdaLbZcyieNZOZDgPI1CyknynP9/+Q7s9qYJkYVO/vkHfQG+KakX1iRzpWpjTzn
DWRFhkBLmuaM6r47/IEe5dppbnf1PDCZ8AGWiZiQffM+6tBe4CTAty2hJbVDAY9A
fmEfVuYCBJ+859KjXx80AXWX2j8FuVIzGgcTxNv+E5u1hnf9xdIrXGvGAUVS4K4l
hqM7pjk/y5Pdc6SPtaYQjYQKIEjCcfcZNK+nwkeROKJGvUIF+lJU4nNn79EB6Fke
3BAixijBDFKnd0ny5+AYZLrx7geJWGRFVOZ+MyHzbqpgy8RIfbUK4JG1Mc8r2dPq
6cSrKSHk0EP5I3YZeXh9UuRnypijW/0mVuX2XxQ3jEaXOp1U797Ou+iYrZ/EHq7A
jOCoAj+AEpDXavC57mj+gUdYDTOJPH18L5qQMkLuDekL6dqhJMlQjRrD6THIleUV
YCGhm9h4NbUAQ3Jgette8qPoXsWE79j00Tom7gvXY3IuHs29HZfb9eJBIlpGHKu5
CRT81ovVWEV9UxRPkYmiHKVUgG71Rrhv9zzC5V30iOngnNr9799wwXdIT1S9XHr1
fSTczI8eTU/Te1DclYDsuGV5qFNDeN1g0FhHseqMxmB3l0b3htqReJm6WwSJVWV1
wxJTBhGw3Joc2iCFc+jGn+0NhJhCqWarvtAnouEn1rzUPFsCNbVtC3K1gag4Sxp+
Mnh6iQJGggtUIa92I6QTqeIvm3C0xKdQ6PXa0N9e0GK4TvkiGs16ttZGYJt2nMJF
nEfjiADlZGVkXElQn8j41p36vzLflX7u8QP+J4owgTCt1HtEhyHiR8p2YUyRHoam
JLGDG50Jq5bj5oVm6uo2mQjAZm18shGUpJx8Y60NhfV/L9RLsJdw7O/s4u5SdDjq
J4PhinwQy9oNL8P74vF2NiuNZ6hEQAU76/7P5WiG7LhvZrNu3vJEqO/GD6W2cxIb
EDLborG3USYpiL2XrjOUgjyB6trcf3xrwRB2p3l0k3TWrpNh2GYwcFWFALUarD3D
HNBS2D3m2Bvqy/wXxDk9WPX/kRQxRTqr5hhUGqwvvcQ81S4de3IwKTdee3GVsN+V
dm7pqElozU9c8OZ510sscZ9H+DQhrfDOS/g1FO29qGTLn9gLau8wOiFgIpXvYNOc
0BRptFK4N9AaTH2iqJYvlDXBawsyM7MGPCNzHmoZ3t+X/H/xhnzbZZhcWLFqIRKT
wHVAVqbE7r8rE4dHZaZjg7FWMvDO0lqok8EoSbxqFAjcx4TBD1fr7SxGeZIE822t
E+fuHOS2Lht+svPA2diPWt9dzBv04ccYEvJ/s+Le5APFErcsxNrnlfKROZw4U9EM
23+AZ19FWl1MOgZ6h3pBo/7hyR0au3uU4pE/bMAvPlWlKievm9GgT4cZSsAkQT3J
W30g0SFkXyeiT48CZ+ewFVUB6vMhh7TiZOYWF3ZNXK6PvcB5ZV4wNQViiV+tNkq4
8xALef5jTDcfV05R13f8IEsJmrrAZcuQ+R8WJMbI3zOQJr8SguwfsSiU/xFsKg4U
JFNV/5H070iD9s56LmGLzOFhQ/IHd88CbVi269/C+oDsRZ3gaQqTNzysOULSqmWX
mGdNsgL5MGbdvK8XgRefDsUuANupcGkljK+u1s0s4KBOQyFlku8IntpGPcHwtfar
KD4Yg5GvS7cF14kr+Q6c7r0oCKpHd3UM7GBNkkh6NnaR7RjkIkF+cIgXPsw7L/zT
IUnPy+LB/zoFCi8oEbkkiaxwTcYwuGasaAf1q+VHLYta/w9AGKSIGzSQ2dy66QFX
gzEEDkJdHFFWLSF/vZPKqkVXD5zoIuGiSl3lAsoznbdzzVdOCdy1tbofgofaZPza
0obRfWKoGyWM+HGOndPho1oY6wBHuCee2suYhUohpVg3c+jYqubb/cMmKakyTOGH
/aubv7IfkEVhEpOC2pJH0Mp7rjEZ3fsmsbm6MqpWCKnBX9gQfOU8E4sCiIXkuQZ/
i9mgo9RvfYvbT2AhBAR5ibPt/Ce051cImefBHKnK1wXUZZUrT1dEDhFyyfPJCziQ
VzVxUk8sXKiQ486piNuxz9aV7pbYL4S5bv7x8mbrJcGPSDFxtkD0UVDiwUbkvapo
AQIlmCFFqBMQE7ODHERPJtX0CwCG6JVG1qTbwmSCvUh8I1SGT6eg+HumEWtp2HRB
x5U2OpC0ZqB3qBaj6TvxC9WN1cF9/c6y6EfHpoP1coVoMDe/YuTt7O6GN5zgxuzE
hIw6WQoBsd29c803oFkTS67tRHlzmi72p8cwBHiGB91+9iOOQUsYB41F5FEmve8r
DChf2hZr3Irb70TYIBTTVF2QlKVI6AUzf24hgeurVIUG76ncnl81ShlFXNxk83Em
RREGkg8RR/5hmfnIs8FPfxuoIHACYP5I7oPzRr+SVTRBBfdfvIvTZ1HjSrH8EbJY
+t+dxZUiB0tD6dhRQTkribM5HIbkhcqN+Cb2cgfAbA9qj3iW495LrhR5h0OrkzpU
kpeHRuAKceYOr/j1RE3CkFUog7xouFwyo1dw1DWBf+o6YHySp562L9aTUF2GN5sI
dEwehw3bxRvEDGj7XTh2ns9O/Uo8HmggGa/z8I28qOEemI7/0USh8hdyCBuYVpzR
pBsSUJrSS1tYGFRGmOmf+jx2TJpdCqmbxvfJU3L6ph97RxoBw1X1RblRhDTeeIBM
tFN1scJsFDUPQnYm6xrFWAj3zde0bx8rlBaI5hZ1E92B0uUbCnUJr0y1G+QIZMjK
6cOcsYnRAT1AHWgzhrOtXEHxyokoPcDgalp+8pnYKCTagl7V0tjtCspR/mL5XMaQ
/OIKuEdHmQDBjsJvHpD+Kjcv4m7jqFamOLFkeOb95+3lXRhZsBSyKIkiJhU/iyrv
eJqCbzotR1IYi8pNExGmDCrXpv/i+fqdvziF2T18miy6BkhhHao4tedHe6upVmiz
/W+lkQS9DtjNOwkmnuf7FF10aIyqkGd8gvNLMH5T0QpE4ONF6KQosoH4/TzAprXO
MnVVntwaVXRb9c9VXcPu/GV0V2P12uvhoYYjot+YnPniV5cd/ci+AAPdPFQcpzI2
JA0nkC1IbgKIAg2cjOfIUSLOi1DfqJBK9h3rwGlUcmuB97KBARBF+ZgxRP8EGfzv
I+8+X77WB2U1FegmYM41ez3Ys6MGcPvHvom+me9JfcFQtWqSf/ppG3Xb1eTpt8Wm
LanBzicnMwlePlFytPUSALllx5iWrIrjXQvNU1FBvl4hGnXQKEJrboDkVzmqZ5vh
W72/4jbz9PJBKijD4hujySJf4hyJP4USCLNlgFr0NCTK7Mq50CsJvHIYLmR8oJf6
Yo0G+wIQZXHdd3V4YPJ+knfq8R3se6vZHWH8f1ThJlh8vJDEXIbw8xilLh1DUlKz
8+PNjAGV5s5AzWWYOOiQ0ml96Wl9HwEGmvivWMaEqXVXMtoOHrlXVJsuB1gmXFi+
o155lClpUXFYOkuMgtA/BwrhwvuVM30q+xzRtCtpQcq8OexX6SFY1kubnYiL2Y+4
peVbvI/uZyps9HbzS3ndeQXubNKJUGNPc8oo9dPZPm4oG0XhQVrAhfxiDHyw8Vii
Nk3Vik8SAam5UuUsQuFvv2K3Q76IkTN7uHeNsSJDsX2VOmq+T3oFyNghgT5uBXDR
EGjE/Q6QHdL7P53RtX8r/8gmgHAHy45T5uYlEUHrUIKCxNhRhcbpf6I1qG3WnuMj
zimAjizhL19udGvMuvEf0CactA04ICrN9gtza0JBVgMpmB3TuTY+AGDb2eAZaM1t
P2k2mHNNp+Sfo+DXj8g1BCM89h90LJ8Z/isEbzqLpGVgRH0iSe2LhURkGC6I1psT
jF0hAh4Oc1Vn6yFCk2NAniaDiugvJ4GAYhtvpIsV1qX2ipXOGRQ+Hko3Mt+ciPkL
pVvwBKltmOXxSlyTnkny+nRq1fRj2T7NdkH35+3/i8BUcubuQcVGMsgDVpOKxyUF
7dffpPOUu+lw8DXVVVDt9tyRGCn1XZlwYV5fpsi3JL5fsbd/CDeTh7F50CqmbQ+5
pMQuH5gCPIv4LpvyEYQVawEYp27HO4ye3W1n/n56NiPVc0IA6GBJ3LgkpP7zCNk4
8k2lgffWL1EhIviR50jza7PThFn4m/EyA3NMIOTaxw09Nkcx+7DIoSO4ohootDzt
yuMBNgkg/2IOsNEUkF1z5CYFuY97dYYOtoqT96mJxrBIFY7uoXIyy/DGA4ghXbkw
gY0f4ToFrDIIVu44V3A2rtcF6Hw/g/raogSah91O50hNkY/OX6CVw0UmSaAAcOHU
KeVAy65Iopb52EahnvTOavRiybC1b/9thIo+gGYidibjqhCsHQR78oByQ5Ng3l63
4K3cxjWCdsA5MMlD8cc8wIXXU2ZbvVSAK18qewyZddQC+kRh7RkKizfIXytsI8lV
HO+LKu+J6BTp4ltoH+JE9FfBXOtirhonzITfPeXXYSFRdHRo8/Gd8pbaPeftMC2N
pYU1P7GW4EOXZR4M4wvnbHaNys8nsmy1+tAT/Ads0IzWWfBatmYghj6eHYfYNfFN
K0NJzJDTB/X7W+sV/7HtREaLLslYcEJ5SoJbjrVwxMK+0ho7baej15GQZY5GRUwL
PZL4sczZLs1ojU+Di+X0uHmU/GElAvGn97xTEV3qXU2M+E2OC3I+oRPJ49WKzqnV
sgDyPCpMRGyxxBvzCEKBqT7jGq2vCNVizBbK2eM+01ZS4z2gti5xpk3NIkBwD3sw
+rb6hTTq2tQUpaDAvuG/2lavObf6zGPsiq/iAEO+vL7mNuHLur5x9NCFohQldUIM
+UNgy+DG7S/CQVRSmDuQCau4/WIX8bTeSUTbDqOALO8uHxsEiV4IwS2xEe5n0U7+
ECd2wtueMk3HyzX0wL6yhzEGgw+aNqyAARmN1FXmnffIb+J/b3pcwjkau9oVR4/P
bhNApe9QDoA/Krf/sNKxqfdNY0AlyG4Ue01ugui7IdZW47k4UsQqYiC+YTi9s1kf
tH9PubwAr6aIoAaKd7YOuK1KTcvhKbW2BJKj44E3AJRJEGinOfJ9Wm5IJ9c3pAKn
U7DDdm9LfjR3zicmL7y6G2orH6z3jFjFgI7CyIiGNk6v+xr0kOXSUhYQ2jKSJlCu
Dv7Bka9b5mixnocb3tGuT4DLk1MWwL1aWflQPqta3j1QJvUi4QqHPAkfPnegQY1+
tdPdjhyBaxCdRShHwUMw9Kpxc1jNJX8SM2z1A1TAqfEy0cbA0lMx7Y39I8NsfzYX
ORSk466XZaBlXs6Kkx+WHw+4X9a/187mnFFuLWj3+z+b5uycTUB4coEimY0lUJru
YvZ2F3OAal4OK4yam10pTevCX/aqrchzvW6TBaACd4B4M7svZobKgU6XsbhX2BDP
BRjKDpjNdlWL63kSUfM7b1+79//iCyfSAGpKB8oe4VKnqOKY/zuC6bp6UW/mxjF1
4av0khjwhNLFDZe05jyUNP8A1pqqebZFvJdtl+XdhQ8jg4MSIHKfpEjwrQDszCYY
wcteLbKeOEgx5QEgnCh6LQDQzzHESYb/JIbRsnrZYoarq+6Q1+CLrWXNfq/mDeQr
J4Gcl7fC6jsNTPsmoyIvKAFRVLx2f+2Z0WiJgl9fbgSEGZ29rb/z+g4ZNc/DwQuf
ECKM+M2zEkQz9JdVe/BhA/yUc42Tnd3as/JNriBBn2yhhvzqJFs1FbSyGhYBo7+A
I5ZJWTgVwqJ+aSqipqiAcuKiNNSsbUdblQBAZH2Dhp8nnxMXYPavLSk+Xy3MIe23
wZYwdT2nAJiHP4UEp1W+fBGh/4mAXkHJB0bbN8Zrgs3kjWOmoIGHvK8jvpmeT2gg
8fLEEL9q8xMLcHsy+1E9Wo9MI5/vdsHUIozaOVGY5cu7etrpUdW02pz8+YBiQfOX
fHzjSKaBIQAiZmDMD0x+H4WRtd5ScZs/XpTjFxEk5zmc9HaYfCFsnjeuHSXL8poX
JYbhqHbDnfd4aQnSuXdVYz8j7t1OhaBArgV7Oo7Vtb5V9A03v/S1m+GI80izB528
4Q7iyE8g6Uc9ubTfnPihlh2lmEIAc8Hy2WRNUTDcJZuPWBFxPubHRE7m6ogNhUX4
f0ZptnYi6W/jZZ5AGtUMKPjEmBDD7Wr+A93V0jiPv6UIZuMn9IsDsztNOhWQ7Dqm
khf2AqnNxzG9W3u1+qds/Wyv/cuGjyzQTjjoJMJbaxfCBa3Rrx9tityCXPBLUOPC
VybMOxAxCQzmssYz8IS0VNG/00E2locToGzx10jusp2pIcHClXTIqI1tv8n3lCjn
/0xGMDj21za/59G0P+wUQR036rm7PRRyWHic2rfL0RhHhcznV6fQxBIGxV5d2W2o
T22nILaNYO3RBN+ex4rk6VESmHN/q5gjHUH7apLxrGGcjIW9CaTJoNk/hLKOmGvL
L6N2gBKUzZHZrgA/2Oh91Nh9cflm7aiQjbEmOsl1/+8Nd6ckeYBGr7at44ppUHdX
eTlrUAKMo81PHDhlEqIfvP61S0fIbejlCKR7Y0rla9TT4dp4BgQGOgxAaEqRjKiS
CBkj+w74Iff/m1CbprtLRt73Ijlyx4LVhd3Nt3NuxBT5bBry+jbI4vkx1GJAu6GG
/wYIfuwRFZzY8UP0nwrl5prypIurbs1as5yjcw9+Iv/dO50ATZEFMz/X9RfAXT5g
fZGAcqLqFEgUkd0f3FvXUIlCfel1pgvS42GKfS7JDGvEVt41BQcz6itg8T/djOBS
zNhvDM0TKEMgIWFdDmUhH5xGy/mLp/URp/pCc6hrMVOw3eCVljfCnmB47Yu6ZBOr
sAHXssI6ciXd9KSXrOoafTXiQ85T0Yxsh4VYcz1+xnPYvkcyqj9vC/KTft6g5zXD
QKlIS5urpYvEDjEev/FHsxRNm3MJae3n6DC3eAuKbMi7XahkOSNSylZrqMCkW3EB
RdIEJp70YN49J33/8RKNCihld9iQLOjlrNycvfdj3ParCnVmTFmXTS+5+aJt18L9
H07GPe/KP6t+1d6dLew9LuNdoPUlnfHEpKO1Xifr9y4AoNRvrTyeT97pyepgFFbQ
OaPOWcn5KGFIgEmpGAcUTzdiAf8Dnj6TEVDtDwBQ8DR3fUJTU9blll0sFgRYWAJ1
eRropkh4LMapKkgQdCtSfJpVvs5NHxQ4NcO6H+oAcft1MFpdavr+R/TxzTFOPb69
s5mHMriNPjHYXiQH+mJXCLhNlwgO1crSNMZvumHaLO9V+th17+YX5wLW29fraSHY
K/GitSG+Rj2ObTWu69qUO/nJh07D7p4WcJWkplfOhWaEbRFz/8fYamA03zyBW9QS
K8H6xpYnbPBowXFEVfAvEMRY3IgjnKoKLm8vv1Yi3H6lKNL8bRjl8ksCLUv9xw/R
+JUUbGiWIMzquDlr5Cl8XIboEO4ctPB4NMYXQ7pPbc82D/yLi6Tkg82NQIWVWNfq
6zWup1iaxMHnF1zIOPsyy6R0bdbItw8mbjZ2RfwFrww3KElD16D7XPhSYu9PDJ8e
piDYrbdXtuadSthzvMJPSYRGJzF1Pf8QFlbwLqXK79IRhUdlcsEIHAXGu5ywguRk
zifl8iyEJVGjt+ZFSIJx76buk27Hl5WH1vbl3XcrZIuBsrBsTNePDp2OyA6QGBKL
6mvwiIRh9Yij7N90vICKLGb6eB0xGTgqlKVj5DvQwq6kJkeKffnwkZMfzhOYxP+T
TC+qBVZfKMueC4Hrim1IgLoLHp/8h9SgnsxUoLtZU0TZlz8xugx9VJrFs1nViLgN
0L9knXOrK2Jht2JYEBZl3vwQkrdGK5LZlPNRxtr7ZkkFd5Lc2xo1gHzzGVEpPk+I
AaIe7KIEp5lxsAPa3Avxao8VLIoK+blhFd7tQaosyYSvB3ZnqrXAV8wm/+rJAbG6
7al/GoxOqAcKX+CxTRTc3/JKKb1CzR6D2Wr7r5oS/BS4E5p3rr0zam4OzJi914Mg
LapPJQK02NAvsvbBI7IZfvxTstI5LuVUhrgZ4Ps1Tl9UfwXzdQ3KSrFSHUIedPar
ABUreeMEZcf0HLx4uB6ubTTc5FAMLm6xavTyQOOlgq7FytKVkyTjk2brop9uP4qi
EJ0EpNRkbsQ1Qg0erL8ki9KnZdLkFR14BfaZA99v4Vs/k135nSkeR4kvZKuRICkT
Rsn+92Bb+TW7UcKYyOLSL7cZHyt0TSdzAWOSP71kJg38pO89BFyayLMB0SN45u1k
W+5FkSKPcbugqPHBHTkgDWenqqmc0tRNy/tcCVCDPr2O5wkrpz6JEe9YCq7+FEna
z/bTkFE8HIeTTYsOH3hnMBPuOUGWZCkr+DA0WZGvWbXOJbsZzRgWulRGv4ZtwZoJ
f01ZDkjyf1+R68uw/q2/l4N7HDZSjbnEqv4X9UNY/2ct6p+UnpgEYDO50fEcJt6o
w0dmmnPRvacEsrkdTekFlkxHJX2noPk4FsVRuoMy9/xTnPMKxZOs6vWFH/Yl1IJf
XDzoALrG+iAqg/E5/JN0emwKZEdtChozyoKd94VJOqMKGRdx46DaMZ8Qfgf2kU64
BUuuBCNQD+56E2Hsd4yqwRX/YUFoy+DcwNNWhpid9yoVqo41PfTakTlbooxVMKb3
4uM1sEgYhz2MrapgNXYac4oqCX8PsIsEunKW6gRKYbl6IlapSNHqJDP7LOyTi6BF
kTZGFR5K445l94cCP209dCmzMcRhwBFWrbx0AFw+l3kY4O8ILN4pEUIYwyoOylS4
r5TLgE7fDBzlM+iCgvov2vYQsdauXaD7UZs2fbOXyKL4oHArrHNv9gsk20TSzMBi
axDSvq8N+jqrpcPChd78+31OsLVnYxYhH34oQI1ftW9Tb87ZNLfA59WBiWBMHdXG
o9cNAoJnf0uQ3AegQjkIwnIbfUCbpt/CjpjsDrfnbKjvbfG43AVB/ypgcG9mx/cG
8Bg7UCHFVgaO+bVDOWOQ97HQ2MWtkP6roWOr0U+2mtVbb/Ow9RBv/gsIJKCGsSq6
krLrdlDhJxijo8iSlXWWtXotLitJXQX0sJZCf3hyUDgbkq4cdHw3SszGJOE38mE9
aMhL4lUU3786Fv8yyhKrVN8/btEYXXwbI5bizQG1Fka7LuCf9xM/+VCnselH3u5o
yzLg5ihLNwGa6qRzMcDIjboa14R8jKMi4jJkqlkccFx6AEPSke2WeL7uS63sMprL
kZfcNGMk8wlfQhz+JURV2FnECS1q47GgDnT9UmONheW0uQrc8/da2XoPxZzVf6cH
O9rMbqd08/PKWx81a9p2nnqGeQgmLxtUdUtDIObfodKrS5YvcKZhzPgbKVVC6cnn
1kywHa9ZKXbnRovY9rzKcVqAcZadUeoT3nLyk/T9trI1cNShvwsP/vAb7ShhD1Qi
CVchNxdgZ+w5iwIpqazzddHjN+3k1Sa9U9JvUxydkxGwdqqHG6E0eXkv/6EYNyz7
l52gbeobBFAEPJ2FFtnWGvbQZ+9BZ5fWJtvl9dX+6Q07IsSmBQYB6e00MIfhQPhd
5FEeF3sAlGGd0X6d0iIdl8DBtaXTXRdIPqcVzCRiDuaNEEfpmvq81c3EHeW3CpiJ
Sed5/UvSPbFOioZI1MtEz6eN9+6StEVcBwTtTGjj6S+MD2WxJKvNUVQ53SkUEdPA
I410Bkolw8ddvVZWetUlPPyc3IT1bXbY16gE9KZQiIz8/+oaG55X5KNkg5Xz20We
ZMIUABXuJzny+Yt6w9Y38Mwl604Psi3/IrZIUd7ZHESugpL6QISKSpgFJZE+GWC/
d2fSC+9wcKCmChjN7c+nZ8gLoZirNBa8D5txQPKAVUywnWU/py0RDwOhfimV3VHC
MN9WGq5ExWSUInSU7U1L8R08BoLjzpxKKb3EHlsKy/bE6AWzZPiEbV9E5TEIzC6o
WsniMqeJjnBuBA5wVE++P7CBf4Hg0g5Dx/6chvjAV9KkalAZCSRfDCPTBYCtAjxj
NklkIdQr3mFnTW/xn25eR4LfQ2ShbxJupdUEqzIyFmX3LHCJpvNc9u0mwT7Bc/s0
VGn5/JeQloRhbdSQtdhKFDZ9s+P6JQIjvyjTdkpLaAUzYst3/9dWVR4MdWF9TB1s
yzVRr68zUn+VLDYABctTAya1KqIjsPauCVb4UkKGECSvIRqO6A9OwlOVFFJogstK
B7RY//uB4GsA1HP4zmmlZVikpqSox7qeha08y4FUcz7LxgSxaXKnFlqrpzoY0RQZ
e2NThPC2XTVfFo4wM0WxPTr+kDbEq5U3O3DRDf2HeScb/QRtVIksh/PwxLRA9i13
4FkD7VSepBgJQ01nPqB6afSG9MynRzIJHqKAWEP9xLYdSbpINPRwyKUKaQNqDQo6
7IKGd/3V88HfivU8cy6AFbmAanTdLXHTMa+TL0pYkZ6AwibZzrj8zJRwUfNMRMNk
np0x7i4oaI9jeI/Hr40rHYTtYGvYakxMu6DSBGirOlcDIGQxbRT8+JNGdH861jnL
Ap2QNLuBF+P874UvNgFnADQrEKjkVs3gJLr0+wYHpu19Iy537RTVb3tS7VKEfhmt
Vwl8zQCQpmty212YmN2i0czQqv0/RT3KisEApGte3oUaqrz/vAO3eKfOC6qsvBXf
NtJq9+YdShsrYGup3eYuSqRcse6fetk3ykBR3CLXLCYb9MjYZuGNC6lQuUhMD1gd
M+2Fmdq4xd/RV8gIWA46g0cMWQYQPh/eJx68AHucFLMnqWcR+4on0utLPMNJLy2d
vURrXfcKk96ZHoF/A49mCqzzuNj5GMFddfAJ0CksuB71hUdpk9U2BgtrIB7bQvrg
EiYtz7sRSOsufj8yim051xfFtWc4mo7vGYbl9VkKJcMN+ARUqFnKf0wwYZ2vDDKu
xRgws3tZ6U8CFMHjrgqJ0j7VIkUWJgXoA89LxoK+wzJ34bGB2Sv6ZToWH6mFWSF+
yTrdLfsl9gQHGNtBMlXKTRcXud6/LTq0xRAes+aURUXBnisQIn2UK3mw7cUVmRb3
XVzMzWi6IGL/BP5M+xuX1MfAfKYPxJ8IFKda4HHv+7gt+V8doBY8SOoZf0j61V89
iRK6S1Y36t0E2pl2mAxs8Lr0GAJLJp/B85eHhW+CmQNyPHDHfwFjoP/fgqDleQAT
MtMYI4p2qBecEI7tOgRrmqRBKLfo7pKPhfFjRDrzvoCJGRHy8/1ku1MC3QuWZ8cS
TymDob2tg+S4Gl8DhKPtsEWYPP2VnL5hmzhARwg2rmePROSzf45+s6hFTYIO/+pP
ABth7mg1567STysgPWGYcwBJD8kXA3JtONwbz9VLWTS9NWlfPyohk+8uiIcIfI7Y
Bmgb1wAexWso0o4zlgnb5cjoO8m6lpzlLWjgRZse2+NJFYJ1KxrQoMjf8RRjiWHK
B1VleO8vr7GdsCs6Vv+mpNDIVY+9RD+YBLziWKdvqBdhIaogEt1LguJ2y0K6sjHs
gzTL0ZNrg6/qismfOFkGNYJ4HxpB0xNCq+iaC+mlfxNooSO28RdHtTSsrgsQKDPE
qjRlzLhYf/FjnHEbGr+rUX2mzS/qFK0+0Be2EiMQx/P5ogEGDWrqrpRsoFShB+YE
alTmAVr/MeHCsGHxTQRmTpHEqUGL293kEWZLXlMEJNKutUIajexhqVbmfgmBXVs5
QfeJf5dGJ4uhhZrV6rBPWs4odCNCMC+IDWSakTdPyOYM4N+YvquYwgA+7tiv0cwt
wrYi5raT/CEVkIvbaco6jyQCJBbE1JNMKXiKs3Ew0butH+8t3QruumuAo5odhXmu
2a+1/WFGp1eAVQ2NXUgb7QZH2fRYTqYDpbOpYfK2IkGfQfqXDtE5Svxd5I13N3W3
moyThy4ADlAW43yPEePp9kko/Ps1DiBJQON4x3FrJA6GSprmViRsS6XGl2MkEyB5
Gv0f1j06yuiKNmCXAC/3fobcINwSyaLWwx6PRvCLZdBheyN41ZpEG8c8lm+Kcblk
MZrMwAB5Tbld1ATem6ESVri80+UI5HOkMsVkXdqj+PRv/iEj7WjXPza9DOEIKn+e
z/Y5CWbeZSRBDYoYtiaKkdfmdneJ0JqFF3JHakhTYZZD9xxWEVpE5R23iPE7QxR8
eFUnQPaMfo5pqp3izTu99UM6ffYZL6EoHRahFwqHBQ7qHub/CvaFNAqjG5/j4eCI
BWAd274a5G7PSRTAfzb2Z5nptlPkiW6UrrCxUZmJIDLL4+fbf8v1I/5CnO0QW7f4
GuIetm+hNPT+RPrOrG8srkT0kJZUlAF4kmH87vQrbPHG35dCdlQ3YL/dTAKgnZ74
OYoKlorQtIQLBfcaBVT+COjDOhKxR9HcIoXi+62hpHvVLBdvH4lEycYiZOJ1OzGJ
TwbAuc4Ky/cAQ72rJq/iNN9uX5QO7Q0v7ij6T9QDN+Zb8ZpDTtVhFtpKqZCn1VcF
s+gXS+EGW3Xjt+UpCXUBD+is9oTXvKqy2kdUN/bM4l6PPpCVea9YkJsy802p9lMV
Hrl4lAsLDjZfJ8HPnUTUe5RicMQ5YfyBne7Xbq6+8xFY6o+9+EBrmQ0AyTFEPD8J
VZ40jhYBPKhC2OoAKPlRlO6sBE6RLBurRZLHPzLOlpF5i/i11bqvPf93wPvlsvmJ
UQv5vFecdsds835sO+dVbDNE6pWvCvvOe4GkarGMikMlkQ21JAWKiukOLw9iAdrP
l9GLiQEaNQvQrqvHi4yiZIJ+2Gmoza8aUgyZ97OKmMGCiTEMOc1KrgPEfV7SuvPn
aLAwqUU4jiDXSy/OvutBFHO1uBJOqeED4t4LDfyqVfOeBSslB8c3s/V0c/8M01Lo
60isG6n4l7qfcOjKpQ9rbNoitxUZGVJhRZT+yCXv1dhxLkXE2Td94BHsx6v7QSOs
GNmDoP7aEbvhy2nVnfuJVmvHDlkz2It1JiP4CZO9AYtOFSHNOOWrwX9rFDFNRJRy
YDz9Zp18fgvJ/VmRZarp3Jg2PE/NMuF2L7bEDoLVRUOL9q7QPjCz9/6JVZTT2MFP
3Y4n81TN8bdSSUKrb/jlynsfvHESAHb6/qzBNbhoRCAqsmyNebjBmVfzHL/3SB/4
8622Y5iEK9k/R7y6w1qO1hl8q5nJ3hBOf5vJOkiyxHW6683sWUcuj77V85TrQFEn
Zv44hwetLoppwLJTt6ZCkhzxKSPjVu72e44GlQ8XoSgfECkwDRn5Q2Q/hn9evkL5
kxdaQHw4X70lnlqBCMB8BYOYfwoAiqrBaS1a2YtL094tsERkkUyefwo5+MHsKOw9
BXGmKA2WD8YyapgL5BIHfCBkcEMGIBRNRU+5GmBpLaT+2/VtN7hWinl4SwAeCVWv
t5RQSR7A/KVwJ1jXmvZy/wF9D8ozEqJKliB9PbNdjmsk5nKFSVJ/XKHGcxfeex2K
pQK8Kh2lMY583zuwUbO3SUtPB83IBSxEulVvIb1gWkfe8Z5us3qcHnpDAjUGaoh9
0gJTPKOpLMShCxfYiUSPlhooLwjDlDg3MUUZ+7Sy1TF3BXfsRc71VS9pHOFb598U
w7CwJZXkSidyQY/gh7FtbgmW504r92qgyn2ZkeC6nbMvuD54JvXjlI5h5u7IRZzG
bNcpp3s026q81DLHJxdnJ4B3BSYBapifz1j2TEH95Vr8kHWIhb4nYEGG90pYdRtI
gA1pm1sylY4GsxfW4PrOYvZDvainW5NKsgrwffu9eSxk39sCkhHOSFjwO2srKwGj
Gx+IouhwZFAQbQvvsr1ogpFpasQvn5kTvndVVrscQ3yPRG0yt9K/GehyX+iSflGI
OhrmpXslMTmrqnjc3proEEHICcUijqbunXvUD6Y+fibwCJ+npt2bGEGd/OyVsxlb
YwHGKU0R8eyNwF7LrMxHFW5kERK55Vfniov11nwnGGbUXttGpPl607OFBuH83hpU
/R3jH+3RmhcD6RoCegkGzZa7pVQ8vfwD5p7+JVkZjKUUBGXht3lwyviWBqVJyTK5
17NnY/5Z1xpRzJm9/1rRVFKYjWrOFpo9mEV10g+H5cWhjXXKYKXvfuD5MrbM3nfn
ZGmntRzthAyj0155Q87Q9adfYXkDJGc4hgvzsB5UHKS06I+b9lFS6CXKvAkeWGhV
SzfZfnT2xTGvYKc4jxDubML55TLUwARKAx7RkkHG+euJS52LQCpTqJwIb8VxzSw8
agnHGG9evl0XwcrdomMAaPxhL75WHvh4OXJpkH1m4Xd7FnG5jLT3TTSVyqR7Xy5/
gm/WYhi006yflPiANHAPwPo0Rp3Gc5rI+oN5+xk18PbJcFyn2U7prJBpS7Tb7DxK
imXZgUGoTKI5/VfGhs1aSUHf/vQEV651vRzCIfBmxVJG5soU64ZaTol6tBh709VK
i1jFiMQUAVW6lI2TAefzyYFPMJgt5+ZqoY8+NMpTS7HDDLC8cke4SiNL1be5yOig
vOfOr2Au27A9X3gy0O5gQMuScgORvcSqpoIkEHMXI1Deq3yKLPkF3zZJ0+MrIOFN
YHBly2hL82zbFa4S/pj4U6bld+VGYnD2106nBp0pom/Rjfz3VQIpQL9JlUMRMM5L
13PrzV1+dgdY1h1EtjlHhLQIhxxjqIxhsLvkPbSOTZiTGHXWAQlkXTtKjYCfWWTC
Hv7wznsRCsufxLsK/JcmmCnbJyF0fQy1xBsxaBt14w3Xb62CDs4CVX8adEUaX1lK
kwOb7qptJ2J2uUPJ228qCkEUfI/XvWZu6zgXoOZH4PLqE1sSoSCL3hxIfIrOh3Ev
rwJblEomSNkqTu6MmJF95dtidCi7NDeP0sDRwCaes7RlaRWHW1iAzrWXOBgJBTSZ
8/AGJx3hn+f+8mMn/4b54agJfYwD69EJfbQBwAZD506wm2hFYAnZ4PHsS80vTrof
CE13T1jRF1x8B0bpsgY/zZrn0qEUZPukR2fRxExRdL5AJV1jaXKgMYY74D4pLdjP
F5Rpw1mNBLWs//fl3xN+s5of3ZAmfVbnsU6FC8BMQKiOyA0w4+k7QlGfbXi1epAP
EvV3zhu9tSH8HpwKFxd8ynjNJpg0eAcrqhpuLrI65nk8QGQvZ65VM5eq9rQxK05r
1iZDFpgvse7mXc5t1aSaAlJqwBq8paEgANLUSIkHLEgKLbfNrms27lwpg2PwA7TK
fOrtntrooUmvjUEcNUNmbW3lYnzr0uypp/+igEGLkPK6ikjS6YBNZ0l5zZUHLD2K
26+3FwkNUZwKa5DsE0OxLlri/ERF2A3oMuqrJgmCzrDs2lrLRdX/uybf+8GI+7T1
xckqTA1njJuCg13wrUANPNKHc1FgzR3pcPBmshCH5jkDVVbLPMMZpxnvOqUqpHo/
AqG0PlUftT2s179NWEVoB624ADgzbAfDlPm5AaUKnoR/2wa9ZyDfh6xacGT6/b82
5GpBw0RKHNA/O0Ixr1BJDw7jSqG0SeI0tBrTP1VTv6lEPQ0IAgw8BEadA6St3ZVQ
66K8jWSMy1QdkW/V0OrSBMM72j67fQ4Z7YDuyJrVKuItkIllCrlPP2nIPcooHru/
ivhiWlfKIM/42tsILfrGypcsh3LkhZ7bq2hyooIf/TvH53BFqtMzgWeZCujQZlOJ
XnFAdkia6MdKiTQOJ5zi6+UV51BXX5vXgGKL1olEnaAo0pG9OljaWHwSrJQAggay
K8/XfIB/cd6SeEzVukIf5v0jeS2fteE/m2OFcpb/yq2R3TcGWDEplmomGX2yRxMe
4jBSjHkeIntbvcL6g7ROEIjIjSQB4w3kw4HsJbiVCZlcpuGWAX3nlYT4y/ePtyEU
w0bW9IsOSGIxKuTXVCp2b6762bhS+wAxH9VzbVvgIdJkDt9k77StcgWdHXJlhJOQ
nCGMtZlI52ftF2dGHL8lDlG8W+yDxlCxbSHfIQcH6XwQ/8ryz3NQ/jLmAB16fZD9
oeniIexBOzseNx0CWLUQfZsDNhYYnSQbXmIXdi7toSjuigdOdBbGuPId9uOoH3RW
vU4dVBENIPzh3t1VckMy5p5fnBUHDlf27N9fRJ1HqgplnhsrYaanUTsdMxJufB1I
QQobZ8nEimm9+ZAvnev+5V0SZyV5jrx5BIty5kppQ1/zMN5GfP32ujMZ5QHplxQq
zSm/lk7N3KEqN3PrxAsTEAhl7idKEWxUoZcmvgKlWcIF+VCVdPoXNeBR6rdaoHP5
4HSyNm+7IzYKBjChwc4byp3mW+87Bs0ThsLBpz+rDvYKSnbxhty+zCALFxAiExpF
JFttlI60YNxxmMh9f/J/Di1EBiBU8R/7PD6xfjFoIvmhQZm9Oa0Qd/Sjk6hDCQ+v
4d6REzWyOU4vCTObYRRijU2Ro6GwE1qK3e83E4J4nBOZ13i4arYRVHBaSSAog0xe
QEo+yQ46FgV1lZdF0wA+VnitxWwxxF0bcniei4O1mzUDc1wAeJDT+hrWwMP/doQY
MzkeUAdMCDyHIlJyo4OS0osrPp0I4gm4BbtstAfFVo5EqPKIcRM+2tEj1mqisOWs
UKp8gvsJXzfna8rf+AIX0J40m2PktMPL0Es6Wu67hjtlac9Cpg7DXhqVRGvVnms2
jVJr+1w3UEG662Xmx7Ba+gTgSkw8oUDX8NsRuPNU79Er7/1UHPbw6DFrSPHI3Ei4
AiEVJeWBd0AU/uIM8RbnW9B+otNgjIVFdX1luKxzL4yFoePUDqdIjPoCzYbPvHpE
ZTYpAwXkPDJOFEIXI/m0+/skCGC86Cn+5RbiC1x0Hrw86Ieu9w1fzIJ4zgGaHEXP
6kTd5LN/EtdUT0SyIHPn2wp12oLQusE33v+RyYEKkywxt3xuYjXyX+4QsPx2H80r
+SxV4Kpw3b6wUsg/6mcXhwsfLf1E90Ddlyr2C9IH/oKefLioxAUoa1Wu+qnktk3n
v3dZJwSiQCzqT0pQ8CAzCnkBPtp6UxdAvj9MszV6G2f9+joVGnKZ5W369th4/KH5
VgKXXFLaY/GzPT6flKS8FwK2sBHr1lLLR5ha8whACHn6i1/xqXHfBOLzRU6iH7CD
q0/OEVYLtDtGy1JT/a/K663riCl0/VRBFvG+aotxWXaVDmgX1djQgzhfQSYMoIlC
0Sp36fBV0h5UOeFhGT+qql5aOrYnax1wutlXviPJL7bLrwyCLB+aHT8zz7DPXMVe
5EGSAcuNq7VqaLqNP7FxN1LgYi1Rtvi2/sLqo4yuPn8KuVjJXkQgVaLFlciuBoz2
luzcbsMiiIytHwKrCzWTGDLe0qC/VlV0AEKZn/pGGoM+0gpDdtyBGWgq0J4yU7q/
D0cqm2jTWpobiwNKpZPXWBJyMv2X0XnrDmGQOkVk936NERsA2Ki7SqO5uDz9aiv0
EdkYEetN1Etd1xIh0/yih0uzzljHEDlEaLj12WCmW+WY6tgiwYhUlgaca7XO8OGK
tuFxYoBkj++iLlL/W5tv2M2x0dVCkWiFxe48+hFOXDdkS0PVHvI2cLwoRrNfXBci
RJrx6lQCnPdxT0olQ1t35k6Vaai29DaoQVJa2VXHFGpOgRgI2lPgOH0OKEVNXEUX
XQ1DXn0GrsxAbbVPXBfboH8GhvrqAfVaRJsOcnRyk76l3fmWOBnPmNHjzhUxXKDP
rJF/mWCmrJg2PJVwi3rha6pxJy99g6Qg6hvzMF6nnIpm+f+WcSgwIPinh/H6iDEu
8Ksk9jT0+cAzD66YezGWWhrJmqQPsrFvJqRDd5aTJqlITbLTXPY0VrIkNRvB4Dcs
z40mKdsNK8mePkWukYk4X4ybhSuTpHYoVDiDJDnQWCJIwje97yfmXB29tolKl4gk
AgcCLZxgXhPePVpbJE1mfBk+oAoiCyObU4DBi/LaIXmGVjOiKXG+BtHaW1Naubz/
FBTWGBpfzeN62WqleEn8Fovt4MAEzhYob57rKdFtSEBDl6IxaQg9qOxtsyq1hm5M
iySdMG+uv1vZePf5kModAvKCII3nKWkpzXJoaSpVBlfxlXSNBUawhw2XuOpuQ8vh
+k+j9xmUd4dQHRQFSy+Q6FRMw/0huzjxgYZ0cX1w2WTmiD7CQLLdnhLKUXDBqO8A
av6F9kCUZk4AZ7WCL8UGvE6RFXW+BvMWZi4sOwSvxhmbfUIDzFycIugaXgmIaREm
BePKZb8KqFI7aCfH+f9mLE0PQDeWCLdCrNnbIy9bCFuqUE/Oa/8WHja75+RZE8HK
vDr8sdu1UMkdEPt7tG5dQGoC2I6gfFxq4B3+2vYJi/ptGHfQ5HWVXBdWacaZw/gg
LMqL7zmFdMdxBIfdt5uCvH4BbbaWpt2MzNMv5UXIILgCSMJX9vs/0EIgfKoIw/A/
V+8PnITvoG7YqHHtPLHiUBi7U9axqnvNdd1FSjwX9gHGaQu7LdBQraSUBe/hlHBH
eXzwLVxE0zrA07nyDQNHUt7U7hXjxd/m8khzZ0ONoNV2QBxp428gbdKP9ZN93HrA
RUrFOxW7JEMYIiLbe6pzqpCQmnTEd3gRawLCLPc+rizmmzkRm1DTO4SFLS3dcWa1
CfeOMjxgf9i6Vnak76yEID+QXtz9zA8lpNG4EeZsy3ulF23FKwZsePp6TDtTKvdy
cvmR7UvWkQLbvaQqzEBTcsH7I8GegBV94ZtFxfF2FW9O9phcatD4ANKecCRScUPU
ifiyV5gYZ8cFAQMW2NmFPC6dPWjxeJdee7vKy7IT/55PKSR+kKmpI2OaVPXCXOQM
GaYhNaTljvMd0Nkhy3SI3UAWwyTTk3grSi+qlpMoZIjzwVPmcRejCvd6G7qIBsjW
N9qjrj1NwVhpRCeIH4MyPtVQB7bx31qcLSXl7ja2JhgzeyLisPz1l+f/9VOw1nPK
5njUuuzAFD3JmErTX1Q9xBmlipbo+GBUPndpjICZyTOIPfW+oh3otjobZlVlbLLD
ZFj4KsJgxBwV4DWbKOq7Ay4x5+eqWcGrkjGDCxCokly9JRK/xwx199ee4s/8NnDe
rI1MTN7ep1lkYiIxSqXRAv0Af1LuAcChKH5lC8NvaJxGASL8NykrgTsoRm/pcmf9
uhgUlMsnfbLIw4O/F7C+c+S8F9v3vAStwOkeAzk/AatonWGrff7Gh24E79eYv7Ea
MX0YJ3zKPbHVkWBcgmxM/jkwh8bmR+UaVl4twNhV5kADPlyLnObI6KeJXdH+1ijD
e2JsFr8Vg/gQqLSXORb7GQAVAaqfsfwFxiZD67vUaGbGF4xp7e5KjluT8gdf6JS5
HQlDmpDlNtIuXAFgH1J0ZJ3ox3KO8wjwDXzlOE6WQA33wMXxVGaGcDQE98Hiqp9H
ptMELdpX1JAgoCqz5D9WP2Gh3b+uw9e12zhzvpXTSn6eT63+5sCcGJDyIEElIOnj
TWGMboPMkWOnvXJsHNON83UNSVYJ4WsGmzq/P09vORY8xC8XheG7ZJ1Q80SF77G1
UZYLhFISQlA2v6rs36AF0aDyJCeveMMLygQ8DYt4tLBxEzUfTCMb+ox3SAOXUEYQ
McrurHyUXUWfgICSpvbYyZ51UiDqD3pKot8vH9S8OjaXPHKzLnyAlRJao+JFABTq
fZYxqkYfeOCXLXpf6ByFeH6MjGAvgnTQTFxSwEqUonKdztznggIOFIcuQl1YsOmz
0yXZv/BGHA1ORRie5u6D6osZSfe1OfSRTuSzqOojPUJLCP7WCRjQkkcwNdCWCp1u
24OQdh3/euG/whtEsgoK+xqfQfYBA3vjZ2wF9NYEwpHw+Xa2K9fXFpFKANBukRTx
R0GLmcHwjQKHF6ZJljErz3wAG0hVbK4pIqPD02/Ibt9ywyZNvD1jRxPX4A09jqzl
oZyiqzfbZr3VINjqs2yF0uR+7dluJmldJF53VjioLzZ8ySJpVPNsea8VOjyY5azP
JEnMa3BmTR9b03Hcg794jRdq2y8uGi3HP3z51raVK+rJv1M7C0/UhEUiRfYrY3jQ
otu2VIM/01qIk7PE4SJ2quGnKi1JEkGqq+CWapLmTE1Ui2AuRR8KPL8c7u7HdSY2
Cd4CfDlJXlYjS2z/RK4jULuBQv2ywowfdnSKuq81l0gpIoXuJ7jKLkP8r/vFe9PI
asqTXshuwg0oDxM+BObhbenoiD+DxuAI5OI9190iEs/ryJ9f1bL7jLkwdjmmMV67
uKtgYKmJO9hlP+YVzwXDquYAf4qOIl8pNuOMp9vyOthe6sRbGqhdxfh+ITH/uZB3
RN+Uom/th8koXKZKiz7Z60WyS4oVRM6SDp+quYCewI/KP0jjLZwOD44vEg9OKCjm
KotcoNouWsWt/6/C3V5vRdMDB1OCkaDZQmTinQxCHJiz9Zm/JnHCI8+CR65Z8ESI
xC9/nuqjxgPsT/QPBrNJk+TOciIXMgZCvB1bJJcMQFTYTkE1M9ChW5K4C2ABcWBA
TzMwlLNzCR6T/cTVk4ZGlZQfLW7VAkbUFVpIvYHwXPvZd4wsT9/W6o29EY/ttB12
S9U32M9MVnCwmUprMiO/yFBdpWHecer3B3iZgr5AayyRDudMMmRsPaseycDwCm0I
pOsBDFzur5CAUZPvKp+QSc6GRoX8mHkJSE0hXmjLOy7ZDOv+G9aFHItxmwfJVmEG
eSP2B9tDEu9f786t2p7isU8R/bsAqddobl7DqiyXu660fc6ppy7dZwYXSHCElYer
MSGKWXE83dcAgZOk+p4PoNz+Xauro1dnHYN64zzFmru3p9B/BQ5cIX6Qvhf0DUtf
xbJvyJ5P/06JK+a/joG7sCH15RDzEwXNiRRHuVg0rTXbbvD8HOyqAZns0An5S3zQ
kKPIsysQL+cgN6WTGhGpAIityabuXwOIgpAQxXK0GrmHX/bZ4wKq+/tEMP2wprNG
eL/0CQzneAz3gSF/xX8tDXvPxCMVkD43umbt/B8T9yeo8TsV5F66IKhnpX0jSo/T
y40csJPwMxlMD1XmcyP9zrKXYiKuBp7gqi53+AZsmdz8ufiVd+si8wIC74nbaGiT
nvMhaGS6P9ZeFSr9HYFoLhz971Ku5ZR9EIdUUHZoEMKvz+iM9AoBZVPo77jgxRL4
wV/81fAwjh7rZDdXj4STjZYzeYTWaQrRQ5fXOV7XnxyQanMfzjpdb6yqodZmKS05
mWpnwXMPDntfO4ITTiWmNDGXHD9iqoEiwjBvrAbOTwd2O+U7qChqscQZX5ZFxRSR
FF3k7XWn+0CBJrBD6RAf2waetmrV+TdXF+zH2i4rOoGB9ji06spXJxCbAaXdviN2
xEoU4qiEFkz1JwxR37nAAJ7mFnQlmqJHYiv4nVx0ojhYbl/i8IZouUBf90umOmdT
eo/XilboRAe4zTU3ALAQ2XC/nCkKk3vE2W9aBrlgBRhkJBE2sg5g3ipsvU0G6neF
ap7h5uToySOsmxsx588HeJGEO649hdu2q/3Go/Ohc9oQ3trlmgBQY+g+mpZUWQpp
Y5yYSdEK661AvAfjhBoCdB3e2aXKLkkXdghb3zT7WDH7dNI7nTAqmf3Se6qyw0r1
r30auZ1ZFBE/zoh7B5X+FSSEraiYmDsEO1f730KsuhHtB6Pb9PACRAehmM7MsHbQ
RGsQcsBEjKyGT5bpHwZq/C5NDQoDnnqUNmHabEF6KDe8diWBrj2vEghpOlc9AiK+
EpBjRGzMCGdKBtQseqgwnAx/+TQ94+ilxlJxcqJ7bkx8XhxKDIf3NXEX9Y5VKwzn
17ISBmRl6hWC9x+iTnba6bisOrge8hjNwUuGMcjUHtSJtjEpTIFcbfpKKUD/mmyY
04G1QaqW3fAYcLpAFSYtk0rAiTzbinf2mSmL03nKOty+WzBlgRFPsrX7o/6R33uJ
T0F9oAuX2GGtBF0AUUbd5Zsz0HdmKDRkz1/knkRk8bmFUJ8I5U2XQ9w/ONtiLWLn
4YdeWQbSddonN/OlTLw/KPavEdJu3jrP+38sBhYLSZUBbRxM6tPskX7vM2CgM4yM
sUkhTCvYUDg1jWl8zJkluc3lu4DnFweCiNVbovSLfPjJzciav/IOcJOODhv2M0SH
shG7TmPpWXtTZxxbPPduOI3J051jAg/uwp8v3zP7t2/GaIT6Xzq3hdIejbgrVEq7
IdOM3lKQiMRbdNolTsKp2AFtSWY297WYeVVZe7ub3iq4qH1fm6Bp9RNYM/3e8e/C
HUd11rnzX4hjmqCpmgC37zpFVIYPQbcT3Eu14Ewk6QAdkDsYEoacES1Y7Jb032yl
tm/vjYaZG7MzruvdbJKg+lDSMq8kmF0ylIqVuwOrKSTHqYZaC98R2WkM0GnfzvLo
DBxqYB5qxO1Wnj8fJ5HPUMR67U4+SDpo946z0+LrEh/fAXb35g9PBBMfL6jWltFZ
V0xcJB4QdtteFIdkBLyRp6WZd2SjnyDurXLLNVlnOgsGGwqeJ2dZ7AYTX1zwD/RK
bR0uKqpimamLjIT7mQYXlL2gSu5O0JOAVVXa61eejHORbwfdMuwCrqGPagipBCAY
Tar+4A+NdR/Ht9EoFF1pl3/oRgT+77mbwzaXW6bG7DvUP0UQwEZRrMt9A68OWRzx
bbOSSnpwBI1Jxrg4dNG/gJnOR1kd8PjoCRXipQnf/LkDgTGxb6QS3zSF1paTwvuw
HILs24jsDhL5Ofwl0onvkrnrfe69cUUJYS5T4ew09qjsM9DqsUyvLTFRi3RSumS1
AgEL4DsGpubemPKSfMZW4VNRCnEwtKdafRX63M8+qos/pGLbq8uOgJ6mChhruWDp
+6CAj2vW/TYBYgx9ozJUy+GKEXnVKSqzftsTC0F03t4xnoLyoOJMZdeRTucmNP81
k+yE+QMRDgmjelsrBrpK8/rG1s63gRbhKZpdzr6IwxP9OiyTCqitqzpZJU8s5VKH
PvsFvmcRNwiKrtfG9UZhHDIAvMWigXSIJGLRRe/Ft/o9G1oHhdFbqWQA3Qd2R8eA
tUzWGuYX01CJcuoZCNsQ5zWTfJ/Y/KZlzopEdJTPnMFVWHI5GNv4i562yslQaZQ1
S1/8w3mTI0CCa0bgeN3S1uooWVwVqIlb31GZCFSBtV9ns2k3vqN5m4W3+IGa6RsP
gXfTXBv9qt7U+E6UpZ4CQQ6Ubg/aPnh5iHCRI6bNAdrITVNjyU0yoani+Hox03xy
EWudiHyAJTyOewRFqCozObSpSqgQgBz9hsTsrjbf3QWSMI0uQ7Q0DZg4K4zybdd8
9H7GmHaJL8u0+puhRPwWd2B8w0Lm3lgzkmO5cZMOK9/Ij7KBD36odflhsU1bjvvT
lSf7O1+6F6BtEU2M9K+NHOtnLTMsz+PcXBVeoi8y2+E26Uj2VttCw7d9b8QAZvj7
WlZz784iE0kltO/fyOjVTJqz+vd9zyoUSXtnW9+2cKmuChZy/lhGxS8WY7nwNPVa
eFhJAc2k6slmNjz8SCcP1f/fm1qbfxkHvXMGwXNos4MAGL2KSzK10og9ObGaxDui
1NnFK5MVizGimw9U8ZSZzX0ogYfHY9AFG380PoLhwSd+JMhHH5WkogGbiLUtE6UN
azEtSOPP+waQo7m8uEOszReftDVGQP0qv7YpgYjKVdMBQgIZYtAirGoAA6Jv9qvJ
Sstb+RHH7tgF2m+SUqtwnYFMNd7GfQwixWl+O/2yqiEATg3FrgpPA3UN/eTSm0Cj
PdVYP6Ka6RGE3sbtNS5m3qCEv+mwADNof4MlqdjB75mKf0swMMcWY+HROXc67bpu
6CRG5mSeW083tVlyY53SA/bahz1fM4LIp0hH33ClMagd+Wb1TNCJXm0le7c1uhNh
LwHpqfyiff3GhGjHdNUww0JjUDUiqEcGQiZT9xzMiLU/BNctWTwXhphQ+9MzxqYb
ueLQbNcETLnsMaTAQ0qdaID+cqbaHxivO2FB1cWV6olVozdHgKj97k8kM1OVPLiW
kSHn7kzBhB9ptPgfwhKs5DG9L2XRmk1oAzOdI+ZJDhm8WAAX4ySc5sNhVAXM82nw
nwq5ULP6kIposro3i3JxHtVvrKp7xrSKydJISQJOohaJZgfBdDTb/0KNGSukj4o7
ZvoQ4o7ZiKVbVPQXU9889CNTiLykzzWGo98kj9qYrx4OKwmx8maUG4JS7CHEnPUx
I93uHrCIYuC+pDYMBKKagyJsvbZSpcNXthVRJUZxtgAe97/2udsnyp5EXt+iHhJ3
TPJVg+xMmLABvihYQ1lsiY68KiP/TJXqchIHdV/Ebi798kGeoUrJIMOvtMp0RlyO
STBMA35Tk/kAkiA0UrAvkQfw2lvkJgf0SsKM8m47kaXH/Jend+HS4TNOVir9rI5l
RtDA6ilhYhUNJe7WSSOiFddkEAUYpILu6HdxEmUKkCXkxS7Dn+JCn2/+3VSzTlnV
kNosqvWOIgct8/P+olGXEVEnAlPmAiBRlm8qoejApy1qGU6NHr1KxebCUVSzh/IF
EjWKfedxtmJywIAwJKeg0qEDdibUvLTGcbbJ5QWRYGJGGWdHFMgJo702UCk+67yi
OVjyB5SApjTlCZwlnw/9dnfnKm5HKkZwmvoMRyhQRF5gVMgr12Q0R5xLYLeTtiut
AaYDjOHOCRE0utQ9CaNHZbj5kipTd2RpnjwSIUk0BlofbtoyTdOTAG1pdcSgpTLN
1Yp13srNtW5Zm7VLpHuDtHDXzVAMwxoNyP7D4s8SJZHVcteNP5rJzTh7gUOsKxIG
cGCkno1bIyEvqhxt9uqOh9i5NxZkZ0/0ftCws9BXJiwvmLpwXZeN55kkCjg7x41C
+GtA3LM5rg8l7Ar5WW8N+HzLXtfrJGjLRyv1K3INpYzSV7RDSX+NFMW9+IXtYL71
APE74jBbEQ/YGbH1vk2sPeF6QQk7vWYQ9eQqnocn8082UhREd8bOwP9DzPYIlEKM
4C7CgH7Fqm+NbQwtfXEbbRjOEhOa0lQRpac1cxTtV98E6Zwzhe/A5Wt+Nj+tIBIm
UvAL9mFGLTxdELa421YaM4wn8Jm5F0uw2KeTpX+J9toCAsBRRMZ6smRqaZXfAcde
6Wt1u266tCf8qxGN8Gq+Ko5dANOaTFVhdECyuk0Dn0vhoDjdNydkXCNmIZHoo7md
/YJw8IbPWMJVJRHtcDzK5WbGBi64Opa7M5pdq0dsFrJe5QOkVA8tAkjEDLZKO0yZ
hDRaLjx4xUFYDcjWFByx1kZUqa0eHIw5ksoftR9NAH/RhVLIkMdbdO2FGRWuFG6c
oJ1zw313M/g8JUEg2PpR8TLhU1BZxdu1gsS399TaiyjEh88FaqGTASS0hwenUhYX
zedfKVPsBliICQv2w1NFl/3J/942XqEfp8mvNz+eg3uNX/foCxh9u9kOMxeKk2ls
Znb1Jhg62BvwL2f5uyrU1fFBlYRhjN9+KQV79ZV3M5tY2oz6yI8GZe3CZMXZVwhY
7BBF0PBFKFSmXR5O3obBgXBmaagpIcvCQGWmxnZPOR0Ex4fkPhgR5PMvmCIkkhaS
50iScQCmd+IPugx690GM6RlfXZ3ir6JwnbxolhvJOVjeVJvcXvwRlSj+BLHFPDdx
t0mbthb+miP4ygTwx5AChyXtSsf1DVAAIC+fkVuiYQkojprRK59gzL+R+ZJOCfax
Ezmh3xls3NX/XsWm0Q9YAOtcvGY5bOV9XeJsvjeQBOQhvU0JKdOvZPrVMOPX8nLq
RZZc8pPvtj7JNmJ84Z+NvWRH8Et/a1zjQFU/6EviQ4/Sd37G5e0A7CBDjOUjq610
OFp7sSpOYk8hWkaP2O+GfS0jt5j/NhEpHV0oCoskyNFhNXJkuDO8TzfQxKOPzEMP
WE/KVOmsTAllZdx0MTdygsWs2LmJcGPhaAACyeKon410sgnTVwVjOhsLSxr6C63i
KedkPbJLymF1KDUQmLqpyas+4eBYfGXlUQNiMRfbfDCTrOMXa/F5GxJHg72nfX7y
Ay4WYmWqQek1GcUcf9qn8V82xVyneNHGFJduhoimX2UFyvfVx7AuYanK4SkIV9GF
Ldu6we7xcRitUHcvA4VOlR+qE/VpPRjhIrtyItvW4jWVBAH7ydx+npixn6bZXaJ+
E1E8Qt+JFbe41n6M/3kAbacxZWMZ5+RRVTu3OjrD1HQe3PYpllnkg+ojAgZlCbzp
fWB+gDfYfYna2WjblCQzgytT92+HPoJnb3K6W2yKPV40qp4AigTLgygoyFcjBm3y
CkHjZL/cUSyxhdZDZS+jUbGmSH+5DAlxbkzJoJ1iz9BP0RSnBdWngaARo5ODKEjw
ZU4m4si9cf+HSLCCM78br8w849b9/Mv6YuDpHAtwiTa7+6DFcA2QkMSlDJz+Jkan
9ee2cjjmsSR8b8QdSf3KqXZFVVUy7ZeaceupYJ3+T/BkxzUdL3Y3PLJtWR3zWkWH
sMvCtW/YaeKWpdkhOX3N/H9Aa0i428bo3bBIZ4cqrfz2IVNoX42ZZgR+iZxV+Glv
ccmDAQtMmzn7eV5gq7nSbkJIpL+GG6vxCihtJBTKJssYUanDxu3CAtYYF7dFnr04
vTxFSoouAU/IZHOwRjRqSbZGq1pdlj/owUEn+W2/nfM6UYDiUoxnBNPet/QIiBAj
D96iehEd404nPXecaSdRGaV2m2Ge6ty6JdYbrGGcyJ1Oy/gML36eUdrGWQYlZHi/
TlIH2/y3HH+/pUWKdbzrulFHXxjAle6y7Vwx0JvHN7nruuU6ll+ZP0qn+PrcncfV
yKpsedRzlvJPlGrjspf33MAaLSRm4LW15ke8AzIEWxv/jBmJFseh6EHeDe+ltlOG
dU9xk1UDdd++jOyZhS7vld8S9/BM3r8DuB5Vbq64IrM7TC57tXUTsQoBBJKfbxkS
u8n5J1fXXT8Se+xbmow3hL8K7Q+RA3JbAjXII1wuKfZn5Wff+jY2dx8yyA5wGlIO
mdx++a5T9I45oGh9JglEVWPUJPwEgRkdxmSCWPw4XvAw1CTghpy4OXxSnzsn5vr4
A7IymIrfFiu12wgDXEs9Keu1gD9NU0Q16Dwxfq41bT4DReiIJzJmAiATVdA8l8tE
JEkDsvmWObLm04zrjvhYdbJcGNca1zlYpQnQpYWhxoelMptkf6vCxPdIxBuZgrH/
A9pKf3cjXvCi3WYQLcn/kRCIrAI2c7Bz5omrpG8fKFzFQts4lqKTQZMBovS0Nrv5
LVeaHZ4x/Jp0d9DZWeFXFcgd0W6+CvPZlY57fA5rlZUrINRHR2YZrYlGbVgbHC2W
BHtgz4UtQi1Q7yTergv/ouEcucbHlJyyEd+qoXIMXgi0tFTP25VmEEcEL2jGBwrS
An5wccJo6MCqheJ31nQWlzaOpBjT3QPKCX3V2kRbDN0HQz4FAHc7wToQDEvZ3/H7
sToxQHQd+hS/1Dz5FR+mAxUAYVjBVmnLlxG2hNQ+yV9a/aizi4mDaEAkUxCyU10s
U3p0/viyGK7UeNbIR0xa31ZB50qIbOIwNm1JiFa+jp/dLYvv9pPSYOpqB1CQ/J6e
jfHV1nFIs2q2dAgOvot3Se9ofMvHjFPlcJx0yJQkJjejc2mriJrdQjezi4avy+GK
1jSAnlhk2De7kjc74YmNQ0ERNZJfgfA9KIqSOE65ddb1lzzzzb+UKNpYC73LDkUP
9dq7nyQRTeq0ns1KFT81iHEg8ts+GhxIpdqOi66VuxT1+Tl65seyToKAnEtNqC9a
5+9JM0NbYmX+FkJdQr76T3O/8viOCzaVgQQs5taToQHjqXaaC+dd/WFniAbVQ+Zs
13Blou910QGPuA04eV1tRHtpCkwgfVP6mEH1cGzadt7MVrfMC2Dk5p4cHj5wtL3X
JFeqrDZ/weleb18iMITksDdIue6lav4i/PKoAycMElJ2W0ucX65Ba2lw2druTeSJ
r8xVvkWqUxYRSDGZZIYDaKh17PolwjcosWCv1lnaJUGl/MwfMv85+dK0vGWEWV0s
CIQoRVLv6zSYXvtOpIYEJceqW5b8MTlgFhsq2GjrS0d7xqLB6ZhQah4uZ9IbuvVQ
mWP26hTitzhFXooBm0c+5zqu8gU9j2Z+fEUbp2mThfemR/Z6RLo/hVyxPMde6ywB
YgaDyPEH/xJFl/NObwivq+uWBRE5pS4x128Y0dmEK8BI7qB89BWUDCkqcMaY3fvP
BpkB8PBn28wRyGv3e+PxPSXy7V3lYhICHzlr2u4VpHaJ4aI8O3OeSUKZylxaEsAg
9xuaFttfjUoBpzGFD2XC+2FSnmB2d1bIYgYkZZQgb9B2ptHMCCCw8ufAqtfI/x4B
KIoNRYOvVwv1oEzpXs87uiRRYJVVr3mN/il5BSpDvrT6hAZslZMRBgov4bcNGFDv
TLl3H+2f/35yzSOQDnyRYYI8LADvBU1P2gbQzkHDpF6GGmYjjPZo45269zTAy24J
ZrXjGuOdD1sbB4Jo7EejoZItfuLh5LPvC5T/ZjzhE57iCD9IS42C4vGb6urXTx6F
mSoA/qtUsM8FNb7JsC9Dt3IQwyi8Ddmq65cr9s2hOVjnSHr+3v7IotaX0aMxuWj5
uM22EqUHeG1uKu3pbe/E7pMOCwfDBrpZOTjQQTWpZmk07Nl/q4O2Gd7AGeXjBGb7
y/K14aVbf9X0NnWbD8Ytecmx/L7IVcMjpSor0Sn5SOmBUqgUI+ORLHJWrXM3aOGJ
2P8NXT8WZi5G2vzhcjt5gtfQAbcDUSRpp/Mv5jymu4BRHuUoFUrFsEISlk/MvdMx
h1MMMLjkyG1uHCcUlJO1Yfw2tb/yEQAu1sufD9nyODDmaz2PAxcYOm/dvuJnlBG0
jHQ5ud0qMFyBIvJ8qVZraZPKhK61jyCPzPTXWTTjW2PduGRxOdJzGvLSZzleMI32
spgNKc0QztP2BerPm1y8h3ZBm8+2uQfjStjLEs91ZbV/SMVwTq1cM1+1M/S8ejH/
WDDRBgiBeZwzve+8GJKLit1vGop9BcuQdqN2gnNQBw6vI1I8zvh7sryF+K7mCKIp
t80JB64+ANHd2Trz86Oq49VWcDJjenZykZkYrGXMPOcM3CqOZu+9ul0nAQ7Yec4b
OM309A8EYwsujZzqsl+gXXm0Vnt98g8q9lUv7dDGANcoHI18H3+4qAj0a3UbUHnY
hANZNweKR/uQpFxr1HCGhkUryBSMqDzOf87HTi+4eLizErCJydSg8Z9C8zaA7Zn1
lATpEeVRN1hblQzm+wXisvKRfUE3U8YxIzNiGjQFz4M/9KiuIcVsEBfiVH38v4Kt
/INGOXqgTmqlvl7JyMCCp50AYrRal9+in7wjk16Ma+7ZDxFz/22T1SpMvrmpoRCu
MTJMWBWbpCXNKu5kv1k5AUmxZj50pfXOQpzSmdovbq4ptZei8AScbEZjQ0CMSZRJ
TxNkVPA2VXWp5OtNkUj/Ex8x9+vNPqPzW9ogYTCquCAl0yAs9kEQ2aawh9WsSFQH
PD8xv7Zp2cJZXHHHi4Yj8Fu4GJnCcrs6Mrv7euKE+OuRf3V289OlAHgJW4qZrTkf
HRIpqxAJi4atyeWkmOPNufXnyqFt9L/mR5h5St73w1LgVJCNCAgUaSp9DJIouOa8
Rspc0um0Ewrv6sYg5vmKetd6qiaVaD85WQ/vq2ycWA6SFOIpnS7Mk+xU8Q8ytTVQ
443KC9QFghd4XWNCB/GtNekxHnm8wlaQ2m8fa99pQ/T7iTjheHInUSM+Aja5oREj
PgFkp5SAyhWSOXVYIswq3XjQkS7tKRHX+27IA8xDGZu1Y/ZohU7bg2wUlqh4yhYj
C5HAGOjtsUSuIxIR3TvND/V69G6QobkfGv0/RjkckEawalLyDcicK2xq2jU4S1k8
kSOp0A2e+Yber5xcIrCNMld0aDnW26XhHjZLc+qVaHqqXPi1429ennHxlt1tANeW
9o82yCC5pucldlEDUm8Y4D3gbqZmewziu0NPMWq2h3CwztCvhvbUzyTbpRcTAiXA
Ar00HYAhjlgUli/5vrYFINorc8gMLBJ2Evf7LcE0wac7G5MsubU3ZpglWBgqT9y3
KdnUu8qFYSRZrk3CJiaFdmFBGEmSjvhAY5XfbYZ7R5TPrQkfsZ1oyL89PIq7+jqA
oT1shSYJGEdfsE4oDQd2/KT8RDYoCATLQUvQrkmUffusLogkbbKYNuAOvd39smJ9
2vz2dvFF893sHPwezxifS8qyOum3/7l3A0T2VG32Yd5pafYnbmZS4jcDADQ/NtLL
5ONhVwpYoU9l3yy6otnZdlR8+mDFPrF058PALmu0OGOpjN5wbdSRX8JXY1VuBZvi
Jsq0EOytAN/XXRzmSXGbj6Jvapf1gnthVwuvh/jCvTVSMy0GZo/c8j8Gfjw9l81e
lqwYTrTMLOEP0bilSyKE1z9V4zBWsh+fK5So18S84qBuP4O50wfb2yfxQkUy8KHz
f3FHoUFFOxjKuvH37kBVgZgagPNqwe5OfPrMl3TG9s9rjmWNvOdmaEO8pX23vIeE
FX0NGUcDrU/teiXD+EErEhfU7RclRsCnJv2Xj3Tw4BUtROu7nsFuwguv4GN8n7hZ
AzaYeS7ysEyrCbTeUyhlXjJVU6H7TFmZRhhvpelR6Wk8QOUQJax0dDJBXtnFFPaE
JH1qtAv2o90S5FKvzYJmmXgmeHyWpeXCRWAGD6MBrZrGYKrRsJFcxfyd71ovRW7U
WGJI9T5zt2cIZIkGb485hsGwEStF3AHDzxoMdisFWqGCVWDXFndWpxyBC94Z1TeZ
jzmvndKJhxXMdCgbbnzzpEA2j7NAApYAutV2+FhlYdYWLt67hy7j9dC6LRhOF9Rq
Y9d463ty9OxGhzwTOH4/f7AtBrjl1OlHPYs+rZjiVgdqVrZts8YomsG5Rv1u7tPC
ZwdllpX35D87PwHynpCH3L9zeuIoFwjnOhmpgQTg/UHlDRA8Ev1TijwHEVkipHF9
QnvCMQMY3eLdpdw1EnIDv/34YOLT/Mv7i/Va0pPsiVG12vQBEH32xcmjq40K2SCw
YThFWqapC65ijX6Vx1+8IshciN6gZL9CME9z6Yha3qO+R+N7gDBmuU1mhSXH2KvY
zoCFzpRORpkDKMUzBkvCXBpIDWL7r619Tr1dCIIgTeu4J5+Etq7VWefzbp3yE0rx
kBG6PvUbRj2APIT9pzsOIRiK25/VVJYIILb+Xlh1+/Kt9/mAE/b/PJQHPfGo7OpI
MFXInpUNTSJKgub3RodjbNpqSjGWrXKoDw2BWPv67xwdkzbku2E5I+0oMB1Hxs2h
RhBQruvg3ZGBHhCLmJDaRvO5RkEOcYP7p3fXA6jMCik4lH5+dpdXS/8lY7xyZ96X
0T2VJToqt0OW7AlZkgfm+aVzQoW7tHzBFQ7qEeBdUlAhxSHXrzyvM0q/MOh5MJjE
5+0DkMu3jOhYxXSCtlEp6YrP0FdfvLOSBXhGip8iv0FUwq3S5z2O68tofnNqUMAu
95ZEHMaJtOA3EwXlUk/csp2Hmdao8tZxnTrEg24vTvSiIurL3OyFiQpEr+YVzQIl
bWAqhB2WrJyN5HjnUO+i3YS6r+k13pCv73fWkGsA/4AkRCF+VkGUtdbZJisxiePq
WxBx/o1XTjBnBYQ6Ugb3u/blbZfZIM15NNJgxDdwDwP+YbA4UWMe1b+IlJzpsjQs
G4v4fsIcNFDNLmWQeZS9fcASgLOUKKPQu7jUsdW1wMREMDI/7CIftd2XSuElK5bl
HQrj5FU+5QSGa3wkOaeAK/AVPRe0EFqC1haWEEU48jVX16LazNCOEYH6vF9Fwn0j
Tw76fJXVNzKe+e1ToJOqYipFlTsx2URxB0AsJk+kd4o0LAmWyGYeiOPc5Mdx6tIe
nWmn173UJjXjEY6ub5j4aj/06tDESh5mCGZ/QvTIAPVT8/IHrl7amQwaf/nHS752
dyqFYQNRS4atTeEON5NcV6e7tfNNv3bdY5IZPu8PCdO9m0ltgBQevUY2DDMCzAIe
TOQ4+a+0I091X0dRpZei/GHPeO80GDLFw6895vLsuxCUNIx3PXeHtl/oXEe3wao9
c1e1e+5QGpYl6+UwuzB/2iCOm8Qmck21KB8VbFsL6bSpQlb1LyTM4gzD35gtG0l3
aurCBbAqzth/Q/mAlsEHuk1YHEwXLK7sK+f9ZEl5eQcPpL1uDfFDfF9uVQvSgto0
0cPeqAwGRyuyEJM/6llfcNIbqabDRA/E/9dgkzksVp/5+F/DI/lUNyzMKI7aT8SY
GJrzv6/rgNP38Ve+t+K0C7+SYmtjVn55FVy8SKFlR3hhesWYvcfuPmpEfDHGH0q/
Jk9WCnPe//ApVbHbczttAMLygElnwXTrzJqVSWGKjBWyVE21PzCOPWg4OkB/EmS4
Y85u9iyoIOnSQbAt9OCNDakBKzhs6xtYx3fVSOKkA3cOAfIeA/rEMxviS/H/h8jm
CfZNaNfyRSZiYSzxHLIEgmtYZM35f96kgQRNB3wv0Evzfg2uEHwQrYZkwO/ed1hm
YAEJUS/jC5Zun2WzkYCzmVXKY/kPng0J3ArrSS+dzPcaSjSkO+PfCis3Y21wQFuo
0BYpTkZA00CYEpLXvuv4GKNlVxGw3LEZY2Zt9wdae4L8qaQaGoe9Yz5Lj9YPo8Gw
7IcEjrsJAh9OYCQVYYi3jNE8hHMSwt+SxFwRry3q35ALEu9lil5z0fjtaBkZe46H
MZO9rZ9I7gvX9kAlpj+hPR4Nwd++flaefROnVEx2xvvkVRcOz7RmSvx9QKm1A+s5
uDsB2JRVu4S8vDx8khffDEfKdn2MausC8E72GkBGGms9Zd2LhMtNDJnrdKLd19au
PqEfNwDBo64X5QhyOhIA8x4q5Ja5ZH/z+9TLNp/ClTRJQ9vxJP1rMxRGuANd4BeG
eTYw+7I9NLf1izJrPQt1Vdsh553KnkN201ayGnyIpu/PxoRBbASNnmwGry7Wxx3O
PoqbLo0tzhRyTPhp9sGAhIBhwfx1XiiSgyYc8G3IOWUIkG8ekQqZuKwIB07A2flh
Zs+NdWyiz0b3XVkR4K0n3jX1DfethCqfOpMfaD5jTiaXv3rLHSk0jpkHsDnihZ6C
dVmtOOY/w/UkYV5GMnQPpmkzb9JR61vQNZIUz8FbcUCVtpS0ny34gQsYzUWF7R+Q
ORHGZptHDdyaU/dW4u41DOLxGkCDfqeDXzFso1qIjys+kvh60iCDdDeb3tCdn+s2
6sf4fM00Xb9jc84BIo7qUBWentLF34ZvjNjyxXJaeDxWp13C7oThhUCHLRRP9/+C
8OLvgSdzdQeAQan25m6+yjyKFL5ym7LBQ3JvY9ntcGGJXu3M37DDoub+m2zS+71I
gJO0EGKZfwqcM5lfWGwTKn3aq/ChQ51mzFt+BQNrN/ImCvLdfFfP2SIwWfmjmyrp
tMYW0CXq225EzRzAnvAc479DD2GcX2ALQarU5XZWTicNMlCuIZLfFvLHHYK7Ufb1
yitV+b1XCiFT9AQp8DSa4TLChUbUqCSHrXPqC3gBkCd1pWlSvEI9PX5gtB/hvr4u
mklbg7guGX7zBmaic4zRXLUL8Um4sbIIVJ+AsI4g/XGnr916N/fAcbredrvUuAt+
Zas9waqdxLLODepUIOBsHx/h1X7IaYPe1JmcmnfhSVtvgUSVnWAYIv5GRwa+uFhr
KVKQmrH6jTXRfqpB1rl8uaYaxd07H5q214uQODBvUspt7yzOIw0DvIkR7dcs/Spq
9BGd2O/qOd7qpZC7i/8gvu8GJ52RzGT23lvynBgo0hVRGpKRt4s11WOMYPqiozx+
KEPq0gZFz7TvHwau5PUq8nMzCnqFH1gfVIhukOSSt4rSare49GsM/HmIZqeWk3nI
WrS3ikyBAgSfjqkhVOWDgKv8ID0n2SFjnl2AloU+5arxEekakvfQoHihDq7graJ8
Q/+6CuQ4leKC7fvbHAN5sBVdSvXLS6OKgXUgzmsGQfEn2LtKmcWpTcqXpYgkzmZA
yIwZscbxp3ZUb/Ax6tUVeogz0nnrN3YhtYxWlWU9muW33G/EhVXn304gbXshPBKP
9DO8jOzPtFdLHinIKhKdbQfpk2UJc6DxkVQ4BMKLJwsWVhNzKdGB4d6PYZs6CDZj
jt/w+OhJ8hDsqx5vdA83tCbF5c2pwAk+zud29Mw54OQxFQzwz2ErpJyqiKXRZelN
vAblelx9pFnh0mBQbpA7f4CXVEoYrrDp0D7PCffZXegBMgh/jjm+r55ZSOzfgbE8
hB3RObochoPovfsZEu5Qyi5vuIZPn7IWa3fLj4nCCjeb3BNqh7MZIjy67qrNocQR
Z8jkyt3PBLwhT+dJE5oVC+e6lIlt5mRzqfDuyODx2XM+XcmxizpkLK4BwVSZ9UE5
RFpsrAsElsH1ulpzDxYGLqTDzKtSQ3no9qziQ3bQ1+7ZPuAIfWkaW949tdHZ2hQs
wBm1UCCBmQZc4RG2VI5VAvqJbO8WPk1p/cGI68PAac/SXs2z7GkttQpSbPwNdMwx
lFzR1BCmOa3CVcn8rXQN2GUwNaNqrov0GFQXNy822lKFqhHsrHK2vC5ynOgFjntx
Fsg5HhZIKYZZcO3sBRlD8Xfd4bsd283Uw6kEONM6LClrhScIxVc081EK3ofX8f3I
nCismMSFT7zwBmt0d3OEoAyrjRbwIBHKyf+Rf+UoYqFUqHq1rbLaqp5cFAb28Hum
cQmalFj7kTgryD2ojhnpB0LwjFfji7MdU5Xc69fOBPL3EKjFuI56xJv6/uY2m4rv
W/KzMNodgkK5Gf5jVwh4eta3kENWGx9yaSeNqHcwQfelpbHC0rsIJnMEWCy0lBxJ
6omUAfI7oZWln24WcfrIScaoPJslYEtucMB9dX8wo6HyOb1Deg/qxixcoi/F3S63
sIORDCg8zRzvIj3YKjq0vzKQh10TXBzlbKtY/6qECfhu3DZD/LFBrz8C1SokuzJ1
Ot1YUG6wLggu4PAoGh4WQGAGuJgXhfoRj+KIiRKU2dsdd4wNJIsLhSyXAZwknpKB
DrHmYuN3Dn6w1hAUgXII/nv4rjSVRN28DMX72XwHY1uubSMimsUrURkKkYWwnGub
J8c/euYUE4/OaqUWi5pSmVrCYdWXSMxJzMr5c+XmT5dYGosK+KNDeS2zYLiROPMF
EQRFOq6QZxL89btuuh/lvNFDD9Vz+6n+t76j0HO1SClnsOUxzPeucQdbRIRAvczv
eh1u1ZKs7wdS45QjeFFr88MLY4SlNDe2kBjFpglGe6s2qx2X80kMvJUSVLWHFwtU
RM91q3Zyh/h1nVW2qp8cqlaVHt2vvPv0Cv7mZqstVxELfBgACWoahN3GiSHf1APG
2/BN7N37DEfKUeQmQ6cwAEYrcUqmR3/QpRfNW3e19/tlnkKYL1OUE+ZkDgmZZOhe
qqmP9A/OVanvEgwYs7JQ9A8RwhvY7wX1/epAtJDbpYtIk+3IFxAlFiIMDZWdinFd
OcunWFlXFVjmts9+5hF2xrwD+PwGIthI5AaGUiLpBdmY2rHaF335D67kZrUK0xAk
MTwz7YM8dCHJJIyUQyiKzZ2GwaanP2PFBVtABznjtbC3djfGTpr8QfF/FiFfbuV9
5FFmHEwL48Y1CHrUNZtvJx/niZ5pctKX5yotency+frVdJjOO+J2555tENumTuvC
U0RJipKNXnzV2h/S4Id5oYGwaPM4sQ2NQ3WMsalopSaRsvuPFeL5wTaqbPKo436H
jwM7hJau7KWuAW/bRbULCRDomKwmIjl22IFLZREbG8miFnydBUrwlUBAo/JDdtX1
fgSNzJz17QoQRgnTKMMo1YOIhbF7f0UaA8AiitFHdircBsl63g/Sv8PNjthVIfwR
lc6zC2POhq71JZzU5lrruHDWAk2GUfTeHXjNwC+bRnVEDSrLlcD2TcC3vvEGGczY
Zk90cwKJOr5UuIwqGFw6OgFTAViACf0yKJAEvpPCe0rdgUoK+cdVP70TgOMeov/7
vifH59gm5XHdRBR/Mwe9gO///g03r542eRozgewnpXJLX/cOsA0TBmrWdMlUNEDr
ZWnOdcP9Mq3l++7hMwaoDaz1PaALB6FI3WeEYnmrJtwHdLP/+jgKgwPPoVW1DQHR
vNVHN9lXldlQgWIQjeLBHkBPvfdikSzT4e6sS3QkbddZuJsDNMaOOpyhbDghCvbd
EKTeixOn/dIn97HSKHr7U8oMHc+HU3b23Sd7ktHniHmOVxUIbg6epB4J4iBwTwA/
3r+w8gMn+soZTLy/6/2LIrjqMnJqFslkT2OqVf3k5DQ9H7MuXE4CLw+NtgS+zh2Z
M6S3y9CYr0pCBuw4S7E2uzcb+Z3+IgP5Qs7cIzseHxCm63oYiWVyO7nzv4Ld1oor
O5K2aTc+6JFD12pa/DOSWfBHHHsuT9ovbT5DPRTRUlsra1jB1bohmoeayAqlqH99
npSnH1iJrUAckqf6epbWr1hGyXdqLmQwTSYk5ESDvioyEu3YzkxxrVSyTR5oto1T
gLVOos16A+QvWU0xAru8/xvY8zL0EvA+2mbkHhG4HC72ddUaOTqX0KHAUHjsxG3R
ktCRX5GV1HWL/ZY4Eir3KZtT0lz3PTY6wzlpopqgC1thhPoejxOk1I+tp5YhI0dT
PBuBJ3LOIj0rTn+6xo1QhQXNHuF3sCXvzMYo3Nbt2nUJldHzZ7h+YTtDnym9+a5i
+n5cb64nKxe0rB0tPf8lgMSNOFN6aJjUAzeMCgbq4S5Lixo849yb09HjFM3aEVoB
Tyld22yr25Qz9NWPCVERMGZlBmABl+m7ovc6yOQ6rHCPsHWVhdMpMt69XyfYMgsx
oi1+5+hqK4f0IsIsyvp4I6SCrjs+4v17dlEhTUaL494N1SyAvUlyXgiYy7tme1Nl
YLt2tjo/IzGp9QCUOt+18Hl4Y9ikwiwgu0jRvnUbDOFBid6lLhXnIlxyIoxxSRM8
KzquxmEIQzxDNICkd53JkNolNm+UkBGSFi9tFrO0FjhnnctFBpYDRX9rx6t50tqT
2DXHoyceX/YRwYhYBGjWZxKuthqY49y9u+400BQebhNDRFUA1wjnho8LPKC5oAo9
vPY1OSnH3vekUbuPiBMM85YskykXW14Cs+fb5rdfdRxiw2HlsJcX/BoYkAYaX5Hs
1zIzC1sUwyvFhwVDvvnrsfDm88un8jUk5i980+2Xq2sMingP+Q2ELKOz6x9uHh7V
MVZok5wCyERUytcN9KQfQlLkkkFBtLUTLaV/f5zIMR6lsBIQbH7fBwLqCbOEmIEa
sp2V5VJA/GBxKZwoVcpuiBBZfBu0FT65Ogfp8hULwB3Lx8z0nB0inrEfrG4zTHky
6IpcrN2u6W5Duyqf3m4/7s6AZj/qUjhunoAS0ImUUkexthmzudt9H+EvbfmDXVoF
HsJ7cW69evuwXIHi176u1JinDgrRDKfaQLm3y9r9buklxCA54CHK7xGIfksAapEN
WmC0m0RGvGNjKlFX4h/ocBomJcBVxCugrdySqbWfc4FwfFFwjteXCbvO9VVHz+B6
kweEoF1uxXm+g9iYr9MzAVjVN+9byBiZu3ild9xyoWyGJS3etCjIXY7tW/kGPfhX
mmUyuVwdHYhtN1aH7Ox3jwlANhqKYBBPAR5gjwbRc5n8PdAlebpuOhLnylUwfeP3
yi4TrohXSFHlgNe92fUYL7aB/IrrtL8PZQsk6TuKBNLemA2a7nVBLIgzTM8WWmpX
ndPQoA52EJkFuaBfU1aEKBE1lQy2SbB9XQZMsx2aGlVBMCUK0vR+XIMbhl5D3gXT
vwk2eTFDkJL+DO+oGgVsxJWOPSIQo+e0F6hyGx1ATVlaC1FxXhpMTIaE4u45xGyw
krdx+4TX3oRpgygZUpCgVGHzRPAVP4E78unbi59vu+qhdToxuslyRulu15AnKOCk
ebLUczhCArP+M1OIhLMLfkq6f/rxn+DRz6P/SGsPevqyvaz9UhQn/zeLcDDyGfAm
bJYpc8OcKzjmVfAMshDByzjS1vpRwpA2abQzGAmeCyn3ECOfAQPPJG86/wklwSQ6
wUleXqIt/NfiZFDRq/IPZiaygy1T8sdHBJMiJ2DkKnKle7rhixQd5KCWcQovg5Zg
OYRVKytMGXWP92no10cmFdI0cJktpscYO0n7iSExoKPke2FbrBsTnnBZnwnQ6CHM
zcck5fQ579QeVDCnDGqkGJSCArc3fBvTgD1j5cPdI5E8NhFWpsEkK/0UhPtnneuu
Th4hrOTD0NbimceH5CPs0XfXIFul3M/4Ia1PMl7KOojf1p6llfo3YHBwcG/Jid7l
j1CklJRPwYrb1f7M9o9GPwsNxZzX+4O5MM7nNY9ZjPP/Cj1l2SuHiUFFJwfT/iOA
ZSbJBZ//MOj317hJYhBEONpv1WWEfKfK4C5ACd/WN07K9WKNPOiqG/iK9FNOhpEU
6pJ92nT/h/tX1g1M+BXFOHdHvwwmzlBGMT6aGwEMxaq1F3XLpzhUNQTun+71zrFC
DtkRrb3GTR0R/qynro3Sap2GZejLKC2Gx86NnoeMAXAhlpAkKCrNolJ9UDUaA0GA
hnjoH4619LaUMk4j/z3//eUwQCZpEMIUYadD9Q539tzdQX3BMXUXOZIvSJYUgved
Y40E/+zjfiY/3FpA5YaXD3XaOMdkv7rh01p2Ehu/P6Tn3cIf6Ut+mKdt1bTnq6eO
vNMf0BNpzfNBtddgmpI/nc7jTLTVbDNof3kLXRIhK7WEDcykEuWK9Q5uyJuofjG8
qJ5Ill8BP6Nryo+HRxKb0jcmei4Id6FJTJ1BBSm1++oRAyO+i4Z7VIinjpL4vbY0
0Pb8CLL6wCrdYydI7dYQLizx1OZUZnvflOylaoSo2wEU5mZhCGB32ZQ0kiJNFFZq
ceePHepb+g/PXbeSN6ePDzOPiRpVBgAO2lmg348m9XTba/xv5tB3tnY0slKsNvgA
RIbtmRGou+/qw8twKFskr9Qx2ikctLuP3NiLquz4lOYy9QFOg34h87JloNKxFUFx
ccb6y4KwnH8xo/DIRtA+eYQPlhI7yKpDp07C5dapAscCvh3xKR/hYXxA/ST7zWH0
9NdXFTaXn6xOe8bJv0UHFG0qt14AVWcF/ucMyvmqyYNyVpIhjuNbhFNdH117C4HT
oah1hg9cMzw6ib7oGZrrZr42k0zRj28tvre5Iw9gM/qSgJotJ6KUxwrK/J71Xa0Y
9otQjC61YiWmUv0MfzdURU7DwDur+QL1tqbXR9LffAq/Cp+WUCh8hlcOkWo9ddx9
pf/XtBCmkIzko+MtJtQt39cB97HMyW7nB6i+xsYwUrcIYjDiAs73wMAWuToq6HxY
v6JNdWu0tAhH4YhvXGZ2hcW4xMT1+aKj0zB/KJf6LiF5Br9UjCnWyxTX6VznEmPB
/qgohz6TYgCdMAqEWv599lcfO59X1ORROZhElUveIsF6hGCPdepxNoPnFBiMHIym
JPOBplMJN4xBaz3gfGXH0C9K1Du8y9j587H3vjKkTrIU+/qmxdKsLRyrC7hxT/0s
14Us50zp3lYUPyqtC06VtNXPd2Lc6C/fFCI7qUVCcQYMXQpd3VrflNB0cqjEPAsj
fM+m52IB6FSrPOs+7uRaUJX4/cXg4HBZq7NjLlTDDzykguXEIaNoe5Ua1Q0MmFi4
ygVaJ1QQTPRrF+LnPYE/tq8iywC6LPn8FJYyStQQUKONxFC/Wi8XBKcxfgbNsQkU
lhZPrKdZhI3/FbzHeiB8eeS3dPfUZdlfp0UrBfU+r7OR57enkdLli/X03pWaK0o2
LrHYdsyrpX69zNZxcmJEXazwq2PqHtHGtaiZ86hINBMWQNkRWf9dNl8ExqFXgL+i
C7fW+CFWPgNrd+bik0T2OSTF3p0Lq/d45zPdOhTav3nPPSwYMbVYeZwEpwbyjLH3
aspft/YUMTQsgDCJzutshqnVeL6EQVtgCEcFLJhxhYo5Q0RRpd3Zh3nfi94onCKb
0BsiV7Am/KEpDX1fz11JZECNWJQPLQzhodfdY1nf6cQ8sdR6m33+CASGwDn97S0Y
PhH7KF6UNftSL276bdNy7FHIFJw5937F6yN1Dcx/v0tl8WSjYvPnV5Q53pwHbFvN
drdtfymdySfzQQ8iUovgkoM1D40u/1Sid3TURQEL8Wn7uIyonGqJAIYZcZrHOaDP
BnQc11cWtb7vwm7DA9yDJ8Lz0ZHTKlwOzk0w4o5EH3UsY2JYLqjd74kuRdgJRrke
BFC7y8bbrUmD13TLE6/VreuA8e+XZFruqoX+uxCyq634QyVKHfr2VKWVQj6YTTK/
FkbIIQEpiLsBm0pM/86FFrcZbgbmnTq2pwPYQQvhaVVtzQJsnxAL96sncPr3pCTO
5NzE32PnGQnBwuJrSMRk42HXrrGMFpH5zgl+3EKr5udAOWi8Wm/PwM37CBDkfJXc
xdUlIuneMlykqNxTAEqxnCYZxULfyoF+hPdM1VSiOgRmJpP6I/1JJgqmpz5oAtuP
z9cNjyuu6qCrn4m8krJ0PbOPUrB4P+6yv8q/OAzYLokZetgBV5ub3y0IPcjeteJa
R278noS6qdfIkrfwIOig/2xnOS+n2AG1jP8aChuKijaGymvHH11fu5CgUnNX+r40
g7rgjpeFsQLtkdWOg+pIybDk810KYsBk6sy4uWGqVXpdWUSkm3QFwYzYHo50nYtv
WEfhDl85o/8e6tu2qLOAHzBUq4oRaZ0B/OCpBK/NY+IxotkIky9Y2iX/yZM3+NKj
Fm81FKY2VePZCkzOMGil/YknbXhHoJDuhpmY7GTVJARDyoDblz8S4NVN97krkvUh
U2HFx4dRrsrq72iEenBLmVRULuqXILr3xzdQS1WDha8m7Wm4qTElgK6oVTwhwLXv
fNvzWW1NlaaiPFgMhuNZIbyFVRn3i2uUETeNQUGJFUeLxB97ZPiitWXukIYgmkUk
XdUpT8FMlYgBZDw8zc538wBjEE/1i6tPP7DXh1FHQyfrhMOCU8bgCQmJUCnQJtSw
Z+VxUbUoYSyFXy0EKbDlN+y88V778UEJvSw+UFQ7o2obQ3D18eNlGaFoEV8uqLC0
lXDxJFvJ8zrqw0lAT+jZsT4QcU/WdgN3HPA6YPlp2DI4OhLrAfmu0VgdgeDbZCes
5zg7mbuTuIcnMOpitnnUmdQhTP+Xui/5qFZjA6yDo98f2aJPLwZ6/7B/VatKzniH
OrMae/Ixt2et2kj+KUmpRRuvSFBKUq8OufA8KS3DhXQckJDTZAbTDuR/0l008FGP
4BSIZCGeLD/edAqBO175v+SLW20PHGaN/aor0+IUw4jSohl6CvS0c0CUHV1Et03A
wE8a5CG32bLcC8HKpiiOJopbHT88kyUIaIKLOjoubQ2f0XkVaaM5w7QGds/E6p31
GzfZ1BcW/g9ScpDm8HR6o/rO5EB9vbZetMfoWkUWOD83OrXIxoq4HIlo4IQUWJNN
z+y1CZf/RxW3TYNrNgj1yehkCUX0ZoVpIMhxi5v+K20onFqR9CAxsZFPTNainStn
Tjgu9VxY+L527UsdcSU8J//5YJwpoL9hw6+LTvWy2ZalwjsYtxHzvzjCz/qq79kY
QG5ioqKT6h4tYAjTvRVuQjMbef1R1+xAvlpBXhtsg7HA2WnXvowDKDHvYLeB+aMl
+jZ9aCS9CEoeawdpSSL/28HwDdBWzSttNOAKV8vkJ+LOFumOFa6AN3gwmThYcpdh
+8hstpzEvY+P81lwZsBdHh+2lpXrJPABqS1nsU0h8Y8+nbgjSL6l/gR/uSngKOiP
09kILUB3nSUhUK+w9koPgzzJv34tJKPrU8T3BO8cnLxlEa++Wm73UkIge2hjXR0k
HIMGGtnaAypo9E5i1ah3xc/Rlie7ob9uVNwtS/dJWW02VV2s8IJ1KYQf8LvPmH9m
E2zQi1SrQKDyreJRLpt7qHbadOskq8sYWpb0kfkfNxgzcWWt39t06b6eeYsY/hLE
uHJ5f3xIkABOtGUZXTwU73J0vu7uginMTEE8sbJTE+5pVOcyGky+kETv21nIl4zx
lZak4fKlunWao/tcK01OAoeJjXZPoRbZSUn0YL9QPdt60HVRBwyOIHiH6oK6yG+F
uqAjXh10brjlKN0b1j3LW6fZnA9VvFjXnpgummWOqBcfQSyTMrkBCfIgUXXJTmf/
iktXvRrgjs9E+dNR1AdEDkUIKRjwd+7InBo+7p0LMd5/pSlkLwKSyxy+OPytJX8W
/yMd60UYg5x7tktyXihoDtu4M8z5/ejtXAzLd6qN4tMhphMTLQjUXdbNdFLxnVBg
tuHB7nM4Td4qSGKj1wjsfznjOX6ObjnL1WMtcbRzxqjj9b/sIjv1Vptn9WnkSuo3
cxKP7jmUXQDObwdyideiivvrSF8cfM0g7Z8G1+f+rcf01UTYoljIg05Uy6qeQgKX
Ogoz8Y8ER4l7XSbglWoPCnlqmWulAu92mhdtaZ0hnkMUZhBzKCpBCt3i1GyEOxWL
SVQo6PpVHkmjalkppCh/kngZ3Hrav9jjQ+FUaAv1ooJW/FTLSrwi2etPBX93i5MA
XBk3U4aivEeQUe4gilhBacUVTyVvonFce1EGcFUb9u/trJKesGeAxCpjy+9L8n8L
IJVGXzua6XXbmjzUjE5HgUOAUOoy0mqRv4F6+1j9b+uIAWEWq65gq8cqxl9MBXEf
27KcE2p4mysQ9PTuSjlT8fMoZ0lsdc3sO+AXiotAcsnCZPhM9+AhLj9won4+h6zB
CcPy81EZRLwVXsKs0LSx1BYhsMptvXaVIcWLy8E3SxW3jvE7jr0TGIlqhp0trVJc
Q7jCYtPCvuCuBt4H/KlFomgN8vgHfWlW9xX5ZDvbGGr5N0ISRQ1spAbfFkpv2aiq
gem9+XvSEtVTZbtWFXdIa/9fWREw+z5HZGA5Dy8MAUKezDO/JQ50iZvk3TEggc9t
IzAt6vPUlAVehySEOA/OiWbsl1ktoUEuHnNIsP/DORpPKuqvAZhawCOPZPNXGFh3
D6jRa3vmFhHWCpjYgIYmTb9hQevvYFoYhk/kdBiz4Xqo1xE+wkvsx/qPuREQbwJV
7mszifFeDto/08+6Zci35ia6d1mh7kcmiAd9Ui9qgfiO6QnPZ2+KKmqmL3x/JM/v
7pQDvsYMI0bpmr2euC5rmGlYirmxy6cfDPUu3tDgkJGhwWgnxfeotQ4W/ekYNxcJ
9I8BoLHrA2ZAc+kNXY4IPdN/xZSjz9uuh2P0Bmv4UJ6VccC4jZHuRcxnnfZLpicB
iujDKgNqvlXVsF6wvVL0DafbJAOoPeegrHHugYp7bAuzZI099lgMaf/OLGxcjkY2
27snoTeZ7WGLm8/DiZGhlihxwt5RXBNxUlTaoyc058X2kwtOhHjxfXqQiNf9q8GH
MVBOFkt7nTLuqgtR+OwAmFHyTrliOvnId1e3o5uyLQOencP/KgyVDaJsMVXG8nZO
5X3lhlHsOAuxeeZoX7miAqScEAs83rMUOm7qzFAbZnHP06sjwHvfLu4FIixMbA9v
WD1CYyCLG6qtQ7JUL36K9y/4z8RkXl5v1jGQn+wlwinVmm3orfvREmLu5xrcsHEx
ee4A7mBcS4kwqzZLirYy6rAzlotXLx+5z4qlR+AeiSynd/R12d1/TVREofHKoC7G
FD22w3TBpx/zIidvHdflQEazGdG6Ufd7cLTvoCtHs+FWKa8v7YFoOS6LsmoGMV7j
pz9j3gqMTY16mSmgg/MDIaplbAbOhIroS+ulVi98C+37SVi1IxTbsuP0+qUOgnvU
mLDjginfdw8KHZ2rcGq8HAlUmrmvJ9y6iLlx1KCERzPsym22Va9GDDdyc3mMjgo/
NaP/AwpZP6vx9pm12lsbi0WKo+HpCfw2wK3DNtXk8RXNeK+ivoSMqfHlXOvjD4mc
zHIrTdH3GJ81QkPfBY0L/vaTplf/IzzeAxHOykZQ8OqSGCqOEXT9xrZs0NTWI1Jg
djLRzKdVME5JhngIPq82PAbeyP+/w8nal5ie2j/4eS3Vl0Ik5D3fU5GnufbcCO/2
0PLLEFvEW/0GWSl4L7jBX+xq6BvsndLRbKf5U02zZXoyFB+9cLlrYol4XCqCzfQo
SeYB1GXSYh6aKOIgiCeVNm2qDev2Ynq3/zXQiCv2LABVclRCAaeZUF5t6dDV7WkK
8NG4nHj1ncdrmrwWsZDKqFEJXnVC/huUnOq+S53IYA48RV9O8X2dp1aXWiGrrAlN
ioNH6M+d2dEOXLjWOr/ZMYFfxAIN7kCF6zS3CaffABR/JhRouDFRDW7jX0eaBf/L
tIqDgT2THyYM7yJ+N8yKTakWaTyN3fP7yqmMfKEgsGRnAjshmmlZYmDF3oWGTcKt
55oudoLfIMIgG1KawFMwD7hQmvhjA9Bgz77CdwiHyA4t8l/oFSPviqIKJkOB0Sgu
TuYu/r2021P6P7uXnKOjhxCa5IzMRcvSlg3J3OhURLVnKE1ysJ6xiHiGh8zSWp6v
/CORY3ozXb97qGb4R6g8vKkFGASJAgyC6C3CLB10yWl+d2hZfqmQ8LxLxaPxm5yh
mm11K81RU1b4ZwXwkGY7yoikq9dKEpxXW3gTof0K0jw77dt1F4V794D37Uk3bWgW
TUO8pCs1zgQyGBvSaiI6zEedM2I6z4m9is7YyYqTr+0oLQkWp+wS3d1vHVEx+q5u
BlAzXNBWiz0rCIBb98uDW4Q8+3j6qpQd/TV1QIMUXGqFESKSpovCsawbKo1FRF8y
jpN6sBGkkLnYHGYuCqR4NHkd6nlDUeecuLLhFrFDdC9VaVGFqfBc3HC6dgHUL/dA
vjWOJXnTLhWKOnUJ13/Ku3etVojqCYba6dgByU8xeD10gWDU+QrHqEtXmeJ1w9Fd
uauyZP06liKCnO5tBVtfIXoeGRMhxKos427bb+cynP180det7947GTKaDT2FAe8c
T8ZXVXvxdoWP9NSBcbwiNv8O7sVsXgponciseqKznCvMQd69PMoNUYljjqe8tIsp
o0ehsTiRt7SjZM//CV73XkV5P9fOwUhyzXKewroIhnkYofWlvsUerh+nqyj0CFqK
m8Gdnx6h6y4OmmGo6f/+hiNhQirG3q8RdRppuGLsdJIXTq+ZLmfqzReaSnWJlLm8
sQgIONIqzKmu1b1bHh9JxpHjpI5STrjlRhSAvpKvljM3ZhEva1gCQm8usFi4L7zt
5ZTqbV0+uXqyKUmQvAjq0Ma21nJdLIQaxuYMBIpR+o9na88FgFBqrKZPfC7Awh0k
TE7K93DDX5sV1UAnHvT55ccRcmSOf3IghyNX+QMOhSuJyfxua0T3HauC77CV+IpD
6rXz5B0PRzAjG2KfgyLI39o3a+CoGxZabjXXwpPB1Nwfhb6UOZvrQ46RKz9mhhmP
nlwzYLeKUAYkdYE3KSqMg334zFhzM0/YudrutMZIDJEI6OA2iq+jfVv9VwxHyuRd
W4vucvd3y6jyKydE6opJDKU9QWY6cehp65ozO+xcmmKUe20xjCdmEwfDGOOB1XBI
/rvBPUAbVSnJyTkNJsu40ywy94v1ho7Qpu32rsI8aIizTqxanXapRuMcEQ91mFNG
uoCnqBdC8IhO/282ki4iaPBgsTPYpdiyWPXm+QeLcqSXoor7+Xx0ydMAnIi+BnFf
LOwMI7Uoce/YNTJdiACUGtsf6K3c2aY0qyve2WSbnYPN9JRlXSFqJL1MTKmoQlkh
RLH6xddg0JZCKgI+yyQ2faGz4csw8GNpGyqHVZXCkbs5LRnUFaGJhRm95/8Nwtgi
Azlul3NtjhQuug4kE1GO/sPiGRT2OzyL3U3Mtf6f98z8NCA4wp0FsbxbilBsEpra
gK6vRlxD+w10OLDUEXOvJHMfH/qacBP6vyQYeSJFpK+ibwo9PrCXRQs0c0xaSUW/
l1zx1FmXN0w29ywVpdacPD/XPU66X1dAm/b3/e/Rzy8GM9V/vp6gnErqf/J5x9Su
ilnryQlICCLsdEkF/+VRz6tB4xTN39Oj0ZBdLB/uCBnjzK9Bw9nN2+faje6OEOpM
Q0oRZLa5n6gTOTz1I0g2ciCfXDoAmmNdzltvTZv535j/bMijZpwP44CgkygiECKr
igmNEXqe8mv2CY11wd3I/qhi7s6Jm8ybykuomPbxCaJ+1mav6upd6VMF7XwsPvT2
KAunMk+go8exI/dES8mD+UgcPchP6aTY6U0GjNEgcsAFHF88Q/X43p9NTD1YR7nz
Uy77RD0lcWnd7OLfbZR6jBM2f9iCGRtUy0YU7w3KwkTLKFvcIs5Z3P5gpl+NI3fo
4m2fFGZ+o8C1T9NSgFAjO9uJ2xnAQBYmduwDK1Xu+a2TEqGdhyWchJrS+o9ln6Yr
AYT5tEmokPbYgiV5T5m5BMFSqetMXT+lPBt0igSjN5fdAY88B+BnZz7AfRuRFnix
gO3Vd2WujLkIxy6JPbW2dV7wuzLLUpK2jW0lURqgK9wAvlUyBIY9V/g4VJY5SOwn
5qpzGKO7lxAk0kft9dZVjzLFYM95/7WqiKEECdE1yoZCwW4wEIRv1C503OrNdS3p
3w9Lg2Ggad/Am0EtHXSpqJtmfoGsJMeJJd2zG/FCEgL4uDd7oco59Ofuez8qOBah
jx8xetTwW9YmxBLBBCqcVaa9z+7ighefrnEhyTMGrOLA6lKfggKLQXZC4pnOecQ0
bcHcGtJVnfZRuBlj3KY/EmAdr9p7OM+TZoDrHHJlQMgG1EM9uxvNNjfe5pQ80vMA
NkZL1UU/NL3Cqmq7uOaiuXt6NkEtw2IJA0d7CHOwxWXiQh1bc8OPciDa4eo2u+SC
VMZKiQyPnKBU5javmhAjthtLv70Iy31oKnZGtmNG8lYy/9IGqzwPmenkqKFQbe30
lXSVfsRA0dUSczSjS62eHqFXdxDX3USeGIJPa7CSzxtYc2fjD2goEPZE6VWVGrIM
L1yRijN3wW2pMNcLAsI8UC3MtZO0B6W10IeylfM9o+cV6Ah5vJVL2qQOza3xxD9s
eicMEWNjgbd+E0zYOVPYDM3Ai593XM8a9cL9FR7h+5l9+vjBIdsbJQTcVrCorUg7
vNwudORx7oA90Kg1I/Vb2JWQ7HWchZH7h4xJvyq1jRB9iTJ/0W0gjUWIclgz3a44
E3U4+YxUD1uqhNYSJNqTAGB7oAAY0Y0U5JgC1d+Bxvfu3WG6MnCf1jqoCc2MitYE
uO7r5CNqYRuWfO7hIFofCsm3ZmO3mAbKrPggNJflDnw4TfVAdsE651GcZt9rt/aF
Ery48e/t6Yc3asHxQSLdMgMbs4ufdw+/oeeUrRt08jdxFXKN06bfqe2p29nywC8G
wwDO6FacigQwBWz39keiix+uiyUhcwgkiLWNiINiyyqIq4PvfSb3+RckM30vnWmQ
vtgfCkri1StIR83CbZkG0QU3kbs3AhcWwsygMphdLyHG6pnjgjP7PupR+pf56zVV
ZC2xU7c3GZHw7iLbeJ4xGDBnaBoTR5357WkblXzf49YjnkfO560fMgkpR+oATv+R
+dTVoM0bZL+ZcDMOmm3VecLEzCRZXebwlqt6e+ohJ8sThXmgEpAVu988LwFKyMUS
pRtlJ6xPQ3Kq9f5s3UJq0IOMFNM6+Q3xGtQ2T+IlRrCu8fkiMjfklrPE1k+8JDLP
rRhrzq5Idg4iEJbxSsOrV8tnEUMqNB5xr/6oHU3ij0/Hu5VZ6jgT551H2GHqL14R
QfGO0OcRb7QcYwKgVkSwBrw8lR5uuPFXMqB5oSZnd0XRLXAD42JowFtPOV0hVqYm
9XidPunDhqHZ2PcPi4hdqe1CPIDWM3+f4cslwSJ7OKDwXeHRM/xlxQ3awc/1005z
PKI5kWxt1YJBQiLv6zmgf3LZiCF4wQo4lr0s4KzlEJbf/yr2//+5Q0YBsrqzPZH7
mb44ZS2z0dMEle709POXiW8/40X/krIKLp27Lq/BSLDVf9NixFWt7rLBoVRuQbz6
11LTHQ2qeuXJQsN4WkSsLcFmCR/lGCHz1ensj8UHi6ts52QhXOHJA/mo7t29Ug1V
ZEBneh09NJMjk1D0LA4B2MGMURJ6F6zWjXoRtq00Nq8uw5R7t97xNCpXzPrmFkAY
LuPpM2w1GOiv3h5ygzOc1H9v0UyLqXwzjcKIsGOPBcpIaWn7rpnF1ckM9gu+l33X
HEFS08XECUCv3TZJJ99jeryaoKIT8jPZtadFZ2G/m8VtyHUfzgkl11IUGtzgZ01U
dQOzuWJ9iRKp37h8QWcKH8KJupSZfy4LvaGqS61hrPFrkR03lufwJgNlfjKRH29X
ZupUFIAOuXjoM1JaKyZgtDzTWWYpK4vGPPS/nkbF1ILYvCkxG5l8L29+iWrsSoZr
WL3GltQy82kfY/RH2NXS3MOrg6GrXq1stg+xtrZD92PFg1RWySUtht5BXHCDMYD3
cC13z+L2byC/ibOu+lF0PuUYAUBIsTE8HZE+n5/D4nr4IvAN01eXZHAbWSTHyd+t
cUmLn77flgiCD8x6rLdhMRPL9QR9TGLbCJL8CJ3k29VCF9upR2O/TYY2fAZOCXPo
OzDB+nCmKvQxulPzMC0GkpXTmj+GX0TrKYg1kcIne9GhlmLz/O4ugYflC8e22FdQ
kSCNmN/R8eXI4JEkr7Y7e3uy9c08Kk9Lv3ga+Th2rhutR5C/UfAyh9hrWBaiEzby
hIkOoTgPlPIL0+NhLXdYaVoDfksZhApuNX/yYb5mxUndCcs5DvVp5HDVOGAT+iRL
sTeqsc899G8+F8CS1jUDSZtZjjmeMJy5/7feJGCinpeKvCKolW5xJuxP7ppuW+3Q
u7mA8DDsrFlKiXt2hGFh7KVlD05ymbnASd+q34And6tH33ItCFIK+o3mK/eZwnkK
g9hCuX6oyk9hvpBpZeUZMea/4SvD0IeFyUW8bMZD8+GE4GqqAc61JyryHDWxvrOg
3nzwcMcyncNj9NiE5qFJjMJwvKusLxy7CgInqRJlnNEOhKa5nLrWHaItB0x+s4nH
uwK1SFBOGKlTV2zC5W9Q18sJVg5kzwoDkwh77FzfEY4O5EmOeSZ9tLQL9+FDddoz
RxQIn9myNjcBzBumm3L24mX0lbIlNNtV3x9FotbQBe6IfJd8nNHxakrUi5arBcQT
kgJIsUYsuGP3yfk7O1ofCVG1Q40OxKgUg6sQ2sPoqy3nWFWmOGIYkxUwk6/kUH22
HwhCkwyfZwm46JVc5DTJxT2rz08WGyr4iIIrZss3BNZQOJQr9qxPB987Um5Jgslc
IW1DmC+6oqOtTJc3F78+qIZBi1guySxAO5tllfasE1LJfNQC0NgmPyEPoab5xfv0
SmzavmjDK75XbpK3dksRGZ6RK4HR8hHhBtVK72PguYYITFJd6OTdge8lRv+HyON3
aUQqeigQ8r0qs10uiFh29iVjmVrLeaHDysSF3yrwGZZRAyhS5t/f11dauaM1XGue
4u4VvilpfuMTvfYET3O+7Pk+VFgDMKN4sNBRwk29fxqpNewO4jZNGmMVWuf2Ntxp
WGgeasLLNMGhyoW2frvIfiYBHO73BemiABh5zdcwxxRNdiWKh7MHyfgEempasaxQ
+7vKEJ3OkOXyErbb6Lu1Lwjfv6KUfPxbsuj3iKTn0AypXXuQTXXqvSEISxirGCsL
V290mFO47yMuIX2Gqy6XE8jJaNhUzqbnpk2PrLr+cgMru6yo99ScS7SKXRh/m7BR
8BWAxkf7J2TqAMFurFx9ztIUX+gJCQwC9u0nEuCZ32hwbkjAZN/IbsInHiDGupcw
Dt1Idfyl+2RZVdyakOK+7giODNFM/walQogyyxoP2sntIhE3P38U+aAncHd42eq/
YecUd72yRiaW0MWKDYLs9HksPI2foxQivIqWvDl7XLC+fWmcF2GxikF4I/nV6wRm
t/hYf249fmMuM6U23B3jD7VYhZoMEuwhOkSC8+p7dEHFAU8MmQpCLxLD7ea/lDBL
gieh3K+vmiFMCAg556YHlIiGuEjxQMe14Voc1BsWLlq0yYk+kHVKjSjaR6yRBksY
1uHiQI/Kj1jOF/zFFzoNR+3Mpz5fvOS0OO7j6deKyLmytVlTNKUQ5WfLJIR8EQA8
MJ2D6zELHnBu7f0iHV5o8y8QkU2U1vsjmRloXLXg9+VEPqmypLmOtv9H27JBp0CE
KIQwF7kKruBl5enKiZAJq5GIvjBvSC52lYje9lN5eLrs5nfF2FqCy2BDP51vgFNd
DgBcDHGPxFl9paeUqp9Yq7V9hJ113Iv9H5XiuWEu1QylLJgINFXsy4J7srsAnobC
vYInFeniH3zgZwt9XsUc+zbfvQqTxgf+hL9ptICzp+8uhpdCl/M8iZKC0p6UNtvu
sLgQaq5A7CensD0ggPszTvjXbCvMLEnCtW+WR+ETJm7Qozpzqa+Ow/12VYwgmits
+TWJ0/flyF9Ev4KcCFwZRdmJHfGD4kOSsGkvc+QJt8N4GMicxOz3i/hoeLuD5Cmk
WyhyJKhokQR0l8W8gSl04SBEuyeuzXhEekj1nLjgAXWn/C9n/OqpqRwb/eEzbCs8
n02P2pGq5XV+JrGBICEN7b8naNjVufM064rnvGPpK8dl7OxGJfvhbjOURWfGY/KN
eykrGjRFPZCxYtMSNFda6Nlcp3692XmpXNcRwzmTSmJrOTSbolCl8yC7NE5PppzS
H31n/0jSo2BETxfPtU1a3lBHwu3tES7WB8DNKZudjoJFZHbUg88hd/vKlVAC9q6G
PP3Jhv+1GFIhKDBF3XGFH8Iwd7tOv+SBTMJiAoxCH0pHiUX+L0cZl9cc/acBO4rC
5n28xkQd7e3gXT1QZ5n0Cg3cMlqGsIVrsLExVVz6LOyZJTTDgB4LQuY9p2TF7qXa
YAVlAAT4dw1tqJdu1tK9PoRtcjHahi806uFfMw8cu8Ekojt0tqnXPRSuRAX/i32/
4igoltpZUufQMTSxVc3LLhOfHuuQj6mvhE776WoFOa2R5xOAts07VeHxFdPCktg+
ledXbnhcnPHtgHwe5KfWc7YhBHV1SUiVn4CT+COmQA9/WatNOWAcr/2TBUfkDPmy
NDeYLbslWikqSVWTNXWxmL2qnZzfj4ipDynP3abG2JegIYpDyIZPDc855ZHoje1O
2TJYUG5ZCgME50UVOs3y6Ebnzz642UUTMFGxkq0lk4CDAlSCde2+FZ00GqKueFEG
ge93BcBypGZsNbS5nKSxRG2DKegtN4RdpI3JVnG4ANsr1xuZlXzq7WWf2H3xM50X
XIGy5q6SuwVczvuMU8RHqy/xMyA/iG/8Vvh/iUAI63HCPQand4JSVEMJm7cp+8vO
8koU17Pha1aZXPxPvuhQqHCkPDv/2YBg1OPftWuuH1tyMGA8lnrWC5g6yBejlAb8
LE1i2/VMY5wunNWD29q2GoaRv5ptTtLV38i+2ZO4y+dqxS32Uc2zGwW7BU7CVL3R
3QTwCWk42yN7TDu9qKDJRM38mAza2eLOO7Doch4Iiu3WuBn2Ud6tMk8zEB6oaS8j
nW6LhU1BX3NpL7sDE4PcMj2IY/LV+xjhJBaC1VbQfV20aM0g+58f8j3pZd5HVdch
PzGZ/ohHN1DUEg23Ngh9Zd4CcWl+oKIf/ovoG9HFBWQM6Izx8XGe+GMyTSmZM7Of
1Y3Oj8Ofl/Au+rxTq1AmPH4vALRoTn72rKvyODmcip9QoP1Sc2qbhBN8SwtZJPkt
dLDdTo6SO1xoMGEWO64f6hy9o1NSl1E0Joq/yvZzYkupz6lNgWaPJH+072OB3cWh
Z79+L5miuasuCSozHCl4flsYpeQALAoAdfGHvxdXHyn29FE5mh3a7zw7BBbZmalp
qFAViJxGmTpSu72mgpcbGLR3FSZN9xPXzVZUEeHG8RNaNh/I/gZGiVJQS7LHt97/
xs6qWSb99cl419vhxO42mOPHh3phTWDoI3Q50cf9lQR6Y6fRIMLazsxwKpzBTz9P
bETr+Xe6HYBED5oJ5sZxuhZ5XNYvLv2RA8s5wlo6MzpRPTxpxQBPgvEsjfmxZqXX
bl/RB3EXjLrXdNQfbfCW+KnHblziIJ/i1VDK+pgQzzBrVU+Z+lTG0v2fUnT6mwth
kMTO2hCMUPIfy0zxcvsaPZSRnOfo4IovZUwxyrris4QILdzpydsriA2nVoC44isf
zmWcJ+ijt5+1lr4iJkFxhISzuNyVot9CCX6hmcgPiA0KPHvMf+8K2YVFiAIKqWG7
YkzSIOkmFx3czh9ueLzz7WiNtwKNL0fA80qUt5bd5VZKMGub31cDSYKsdWl7d/pg
kTAJDopqPVLxzbMl6Q9SSsMeEkcDlRhPF2iBXpGLdhJ6IU9DcWzruEcPBaKV+MBt
UwVw9yQmVrsy8SZy/VcgkySGWdJdoxi8UmGJC/lYeXtSg4cjvccn8zU1sqCqbTCd
DA2LUK3QgkXmQzNWKinrZ2PmY8J4r0y+hoEwJL1rQUTQlzFua/NfhwX9uagG+L/H
QxIlSmU6DaXFzPtBbLHVrem0KtVYjXErRu50c2SwsBwEiKb4lloPNO89y5UgL8fi
+yXS5bPXMt1zxO8D8hgYu3wddCafhE76/X3ZZOuKy127YVzABdfHgcJq7uK6jyz+
ZDpIr9HRBtANw918MeufTaYJ1ht5nTxVyKqT1boYNBWz2dj3dtZxEq6PV2xJuVyS
kULoQLwnrF5NLKeGde6egDaPgw166JJitG0CV9s1GIVGctgUGAnEHG5VXy2hVjMl
MEwYlycJCpAkJDkn6nbFoshlcV7X0cKta7YPPTgb2QnaXuqrDuevSuE+OyFvBhv1
X9OVFgWMWJIRvJktLGMARh6iSTpe+E+ysGL9/fDBclNFNtr7YlpMhxU3s621s+wD
4RqB6FB+NJunrhfT0For6FIQr5VvZf6Rs5BH21JzlG2XIhb1UfJgcfed+yxSKC1b
6zp/q6WYLwZUu9DWeBV8pm8sLpeBmRbOnUZrRipx0Pjwgp1LNElI/UO6splFKAwT
cWGQvgeRBz1ykU0t+NmEQOoVF1lsJ96gRwZPeLdc6D4t9uRYdQ8ETsB8VP4gjbwC
JQlA7/nfE8PfJPKzLyR+EUCDnC/p8txntbJDNIa4cyX03hV86Y5kCPL9OVVFeM+b
WlZ/N/74PPHsmG3WooRxhaYxHei1PndI7nLiqslW3Fj4GF5GyHBQCznPagaO5Rxw
PTkmoJsONl/f3qJ3R9VEtlZRpnUUsLTYndkthR9jEcA1uh8AmC+h0gTg4xaqq9To
xQoak+TzjY+RYsuHPaF1ziXZ3wID10OE6IxBweyYmJOC54xBrGdLOZRgteJSCpXw
H/S4HPyfDhQhyPVltpEWAq8oEsFZ9ZgtrVWTvMbqM3So1lVyvb7nrh9c88dYKhF9
okvhbiZ8rqSH0R8vA3tIOT6BFxiOmTs991V9np6EBfFNZjB6raPwpBMfFAcmRFwT
fKMkKJcUSlr1qopOPs0tMl0YRjPlOLiZDGpKSj5i8B9od+5IEWtMdmeqIQRAKtHq
MruyLjpKjG9Sy6yDISTRSJGNf/K37FKIrHhj3/I0mDYpupzrQgox4BnNAqi/O8Ut
a+dYMtp463NSu4HExk/g8IT3dKDvagy84nXpWVR7dnvkoJ/WmvwzWIiugvteYmhA
LpZvfkN/KvVRXjLAHsnYyp5bATgtH36D1ubl2VT33vT/L/usNgwWn+8x1lVMJQjx
G8O9evRGfdmwHyoCQgT9yRD/T8m1so/PV4wdJ79AC9Purq0FPgPN6qrgigV21e6j
NnvA6Fy2ldp6HiV/8EB1KaRIPUfU/0a1y3F0p6KBcQRlXgMDVAe307iWv8vIPSyc
TOojPASfDfsTmPORSTMWTJNBXpbKfbZvv3klOLewzyL4xKtZuJDcy1S4J5rdb8iu
FaHKe3X5cFX+V8WWtPX/Tp18PY0gw+TcnvwW2zXjREOmoT9bfPb02MU7C6mBF1gL
rprNlHv/I7PKp2aI4MGNDaXT3oQpxxI/NdRm5+Xuf1fVOiDRhlWf/jOWFpONf0f/
4fO/u+aLIHHOjEZSTyQp7q1Lo2tEEOL2tRPxucJQlgVYMPUXZlirR2/ERm8UpR8m
8L3lAD7Fw7POyoSWepD54KLznSRm+Wu/jZNJaQEsTNDZBqvi+gTt6rEjuMW+ld5i
MTz1PRyB1pyngN7Ny1HbTOtu8kYiEdxwfoM6Jl0C1rcAuhHPBduGwdqHF2n9Sgdf
12TMYhRqiFyxBAEnBp75zp0gxUEZg9hA4Jjye4ba9DLQy9nvz5uXsc8rBPKORCYI
3RoWJeYqVJZO7BiV5860JnT5NvmEnUwFEiHATp+em1G2QzDAQag6Fjl5AbCjbQp3
ScCdwCMz//ErlhenUxg0PGLC1JbSyP4JifOkciLFJ6ah5ZLHTgyhVsl0lZ0PZpcD
ZwBribV8iXJIz928h6hjk5IP6Md1TeDBdmDT+YC+2fUDwwH/J97EIFUGH7MwsT1c
QQQjSfQh1fFTKEWYP3+wRrLLSUjOO3DLUiFRa9pOMnCUzp7ebmlaGHLoGi2oEutI
MgmFyHhtLRm1shO3+pNPAirikdzMOY2YkmbbbAXPdB9WWHgTU3LOoJ6OMHTwtuwF
7h30jBymLBuEy6VBTiK04bQ8ETBAt0WwRqj6eb7nFOW36eFANTpARbVF79XrRTHT
ALysFVscEnzeFoKlPGXq9Pzflw5P7cmWWeYZ3OngOJclF0D0ItfVMYLQMF8kkQwi
1ahULEtjdijzj7TbcRRnKdQtJWTriMYP2QSJS+J6lLRPaof5R1hIvmBXaB5cP+rf
gH7KIjtN1cnvoqHH+9eTMkyyMn2BDaEmW4hUUrIUClZmvkxfRNHkZytqnOalYdop
hltv81X3o2zs+pFAbXjkEkX/xgdci5CpzJQBx95dGTqC1ErLYnoFjC9/NkS7tbqU
pRZ9QVCuzoF/B32rlNV5C1CGgBRjMPKCh3WMpeqLM4Enf2F+EZ2iPDpLriMSqp/W
BuHjAtmx1AHOitL7zCPbI5kINSmkA2HjXDIh8HSZyL1l5H725g9MLi+ZoLJz6Ohg
fa/WiDlfv03mxabMPSDUDlwRx20pD0oMyNMYJLvEtk/kllW21BF8LrTtsURVoU78
/n6Cu2TlvpyUf+vfdMlbnV2uNRpt+9TAOiXDUFiYLHVzQujaZwFhhrjFcqgIqD9X
pUzlPvXllTt/hgpgepThGGn954pmqWjNr+cEjT3TSRVaRXxMNE2d9kHk029DuXnx
GMNCD5PwycKLIhMx9ASgFfoqP0os3VhE7i1VN0mnoXmiNI0Va3pw21APkkEdEeOY
E98C4Yv7sp0eGf6eVQWjaTUW5MEAT3E68YDcbQPtrTjP5+5mfI1fy3I7d1ilHUFG
HnvYg93U3zdqWUQYffKcHxb2ocs77fDs6VJFwytB4aE0hMe1IShsIVGS06PS607A
qgCWkcQAuCjqTEbyCvunfvmy/QGct+fSjXU771ckExHq+NjrzhbzjuhedpUltuOR
pTTy+3cErgC8dbNjtEKgZgxFucZF8c42aZyA2dwSdIOIXUz7VEhKfg86e+yLTfn9
ESXzFmszYSfIGV3V2j2tQb6PdSZBwKb4jyUY356zDVbnQ92hVqCSHeOd3sBzXbd8
FiQLWdG4/NfcLsmnzC+6f8JH3bsFFDTHT/iAL/HWvJjmL4ruR9GNrrZpyP4rAvj9
KqXNPgNMOGdivRkeA4/zQ2594mQENz5WVTVRe7plSfXi94x8+v8Ikx2TrKLIy281
VkFfj9YO9o/VT/ZZQJzM//RsO+347NI8XK75PCVo/HTTxNoGHP/5gJeRW2iQEYrA
ZezsyFKaEy5AyhE9vkyz8cTt/jcac8n7MOeG0CvCFqp9onY05OfgpCGiAllmKNwj
i0qEd4FavJYnQv6siJVKnGrL+9Z4c5W5+T7KtS84voUn/1yK1zpnkU/zdufMAb7+
0sb0sRd2gvAs01Wrd5x9S/XwpPjFOHZpT5BBQD91mg99bNu9l1YxVCTfr3qdYHhJ
dzAq+mLJUJAZ2OBEvE54CQhGDYdXmaj/Uw9Gqi6CwVltOM/60MjI7eox5q92xG89
l3w348oN3eQ4ddtb3QHKkbznF9LXMsza1gfyjOOC2l1tpCGKIKd2ulVw+ENpc05q
W1oqSljBiEhLLOUvGvyqsu/aKR17xNK2c1G3AuHoKH1aan+4bXxENyQaK0whzt0z
fZeyUfzuBFSdYK+SSDlW/4AYuwHv9L38PDJiM7uSTf8l6dLN/dlXmlL5l2CUSQYs
+bwNKjkEExsCwLYOtWyuFHltIIrER2M4QRaSvMGWzxIJ/sRK05gp8Fl2lXM7eEwV
dv9084m26EmET4kxpWEtvyjVkdo2hsFn8YCHj5kLaFn2OM+dU0BhT1AMNejiUvNP
phmAlD33hwHig4Dohv7YhPs9ts4/Vb5MdndA4HDECxp8u3z1spFy43JvCRrMktvF
nUtsmUoHqarMPKSd5MJTIxepmwXRTyFNm04EQST3qGHlL7abw2j+oOnfky7Jra55
cP9TtQTOdFSx2B1c4q2KLsAvDz9DWFd2bLJf4s+F1smhJbW7GPjsNtreS3HsjR7J
4JlxDnJLpbIop4x8RuiGqCKCITd/fCtf6zoe8pO+qY50lXjS+Jlnja474ld+++59
tcnkrDqldwxaolyebtHf2qb004S+Fqqqsn3OkzCJsuQBmaZPexynOVIDY3vPAuKy
jDRyH5LxjfcGBir6MHaSBxqKLaRkc1pYoCcLfTKuJ0TN++8QNu6X+/Nt37/VDoQG
ZKB/8KGLT2XyrQ3nXwxY3WXKLSZupaImRaaYgLU21aTW/rgBHVXYrlI56V4c5Xvs
JJIm1Xx7X6Ch/HCxIIAfU0eRBRGW6RnX9owjE+IvwA8dncHaKRPYnPUCtfkM8x5I
OZKpguVo6DuZCZbbpmnndcB52uwLHWUxFtZV9kk/9m0MhP0KiomcWy3xS1TI6N+d
3wlNlumbIz3H7iDDVApAXX/36na1ll4/lDCYhmiH16AS0SQf4j4Gg79ILn60JrFb
hPfBfiQYUncEAhDn1CgJTlKBrIawBxVHxbEq7GKjwUdWCGQ1CF/wcC+QPJesGZ8K
v815tZ/rJF0WmVC7TcJJyDy4NYZcbL2JkdVZZFDs+XNTnSMXLn6xclU5ZbJ/Mxnh
xfYmraS0wldOx6kogE7UcueAZJh6HwJqOgIGMCBTlv27ULTW00uOfhfnL6jZr3Ke
+zg9RX4ejl+UMEYJz6PP9BRAVvqO3T4h9IMh5BJ6euCGl5n9SlZ3kkvRvS+w6a3y
PDjK+vOsEJkgrcKH1Z4e8xcSwkic71YHnRwT0AtKI2sOa+NGA3S/aOfZfWkvYsAb
l+K6dPGpdN0joY4Y2gHIWtPAI1qNbLDwdvYLIB2MFtCbDS16Q96YGn8ukiHALUI0
eYs66d0dytMY4e72znSvffDJ99opznItWGnQR9t+oPz/dEqqs1yWFngM3UnD5CBG
bebFJZBezLdxvN5HMwzBjoECjRMjRrrJOd+5AKCBvyKHbsBkGVpQX1X/VgRPyTC1
uE/0zNEjCybUnj69NViofCpslHJOTVVHwbdX0CQtMj+zRP/U4cS2QLjXBWnHAW7P
bthX82qO+EdCn2OsR56NigKmJfPaoIOi5nWw937YOJ+PWD7DH6st/u7LUkZeKyYS
3/2RP5q/GsGMciZGLJmVmQDKs1hW8n7aZHZWgBMGeovdMFqjJvYgE80x7+dyjN0x
jg+So4gyNFZKqaot+71bxSCj3kEa0lTpPrLDA8ZXwQTU2gsYaE4ed5dIIdPHqiYJ
RMsWKrvYT/BM8ZrnJRNIrIR7ld2qavQFafuRWQpNclTFFGkWRdzvnC48p5lcpg3d
xM1AiwIk16jp5v3L7fGdmjgz/kl+gbhYXWAcMkpgvVeNGm1sEPxUQaNcbKln//n9
+gE6rg1jLtOUO3/+H/yEMvljSrXuzmxbdntL5GPK5EyTHjit7lR58f8So+EraK7r
qw3cD95WLaipiDxvOU4sNwHn+jOgQliq4Rf07gFP42BOeApTBlZgjPvX/zoliqOH
PmN+6XPHT044WM25n8aJ+cbZYoC2pZHs/9jVQNaM8+SKhM7vojVQz1vxiOlRVa/O
YBXmfcLkArke8Y7fsEDh89RTnoxu+1OcOVfFY6Be6whTAe1U2pcPwv5oz00Tkr+l
B/nnUi6K8/kY//eQUlT7e1xQH9lI00+DzArbHq3c/mMZ/liHKdq3N8o0hJrhWY5s
N63rj+kEW/jfexpIqscjNoUJlAZNWoKLdC9IDKtZZlzxfJX7oP3k3I8w0DYs8ULX
c3+vyRSEQ3U4IrZyejbZb+y73rx0F8vDLwvKHtIOoAbJYWH9QbDCXtB6QwjSQaGp
yIAFFI46gQ3TaIxUtkCPUfWcwUiqekTut1mQObdrwCgI6/pymHBfmcU5VHbPXgVi
LXSbWJ6/NqTRhHOuhuOuGNTk2WjnZ4JTzqLzM7IdoQy4dzyLxFINJDVmg12HKIPX
W1zhrBtyP/sEitcRhtDNJke3rgpfJb4TyHP9N9UbXVeF/cjWhfXPwVmDjXQTjUIk
ZorpLRTLZXHxSnKSwkrf1mV8HgKrz46FEn7slbBzlC4EeToH0uuw8ZoYbm1V9KDs
NS8+dchQg25LstDppZS/pyadPTNlGr73Q4meuEdmCUvSnn6ItK62p9j2Hps9we2B
NtwjJlIFZ+b1fTrVfRuoRzicx+v2IpWipTz+QmCUpUH0bZIX0kZq4ynJzc9WX5pi
9nPo6AZ2Ll2LbcF3ef3T4z9lStTQ5cMR93fUGJoIQtYWgbGRF0kzrDy4Zgjsqr6X
tdU89Ps13lYRIJkrnlNQEicFfj75NyBTmmb2TRgZPNT7j+3nXjwAy0fPU6ibU7IF
iwtVzhR1WxmEIT6XmXHR+Pe3CemzlKGGBEaCK93sbF9HgL+9q9v/4ObY770vtRkZ
QjBecW4JAWTImpXJelZ8UgTci5125czjBKmPkFl+j7OwpellU+kTHS4RwDw7C+v3
I02m4H/Dp37YiesPUqabJ+DbmiekTqbeDtxULkp4FtbESZ8uLbP4u3HnKK6I9Y7W
gEaZHanb3yL1/uBTOAJ2vbySt8Z/lnp4K6Axsmbx/7gtO0jrAk+bRVsK1zhrp4O+
3gUHeENhxTECtiFLMkwZLDDGyQTN4mt4PgovFAjGBgqbiTAp3k0EE9B7Tvh1KZsu
7LMFK4YbQpQUHy5DxXbarhBeT9TgHeLtiRxgflo4oqO5OToLWaFM+Bhy4Z6llzSm
NRIqTIBqDCwk5NZlXXYI/LveFIF3OQSTUJGcDQIM5Dfl8LbbP+qRUkpoYk+ss49D
/JebjIPFlK/xQZCX05xZv0eUjji1QUOFJT9FIFWudjzHyZn6VxCT/dWe6wkFFjdY
WRllZtbbtcb56y/RZJOpqX0hTUeuH2lPj/z35pLF0qKzJ7yORi20qjWcW2KSY6xy
HWZqkFfE1X4EhNRKmIa5DvDrXRsBfrW9mPLEPykCgHA1vZ15JuSJXrpJcaxd6uAw
sQCFs8UQkRrUkWZS01FRqnNEZtXrYPyT4GAGD31y3C5XH5NMNpChBnRpsP3hHbdo
6dp6IgCCksqoKo+N/1HREvzQnadET2O1wjvCbcKNz17KUORxlY1GEx+sXBNtImem
hTj9qiXJUQT8z4dSwgYjBupEF+chDXBq9oIkSXzLjWmZYxCAC7KyvBhru72zecOh
leHaOpNWw6iqxi3BDVegmlgiSmjByAq0xTpTem+WTl+6+/uLFGhdqhHrql/PfTIQ
dToDT7cfWrNciPRSQPuWGU4pXM0IWa5vp/9pIfPorX5id8x8ZhTeDD870G33ftHW
7jR7HDS4HHc3ABw4E/ulCpFrw2ERiI8cG3xhW8iAeKoN+HxPOMkxAMkw8jB4KoMg
x6RcWjN7b4gc7pz0sKOknZfPdeykufpm9sE1ELNHE/KegXGcVP7eQ4cKEinDZ+WC
cP5xuRVEuV3QaXtRZeYhu3wfW+5iN5/FVPKSWK6ml9yv14ytC+mN55C+J8iKQ2sZ
AcnDrgPpZ96WQPlNlHWFtC1tPfgKNkKmewZr013OJlsoZhidUh2io4f1fVjxhQwC
fziRpcjXJTY8CQRAkPATI6c91OvirK3y+nFU4uExtXLEUrgdWPQJZDjwpKiAdu7X
zetqfVoVjeA6fOctZinuce+l4UGQ3NV0R7fqrsx8z5OSQ3Gl+jkYiHIEj/HYNSrm
ErTIJGjvyWuRVqbjpmhML8+IZHkSkkPDMsQhVGpS+x5A6SlOVtdMMBD/4Vihb065
x7wo1tz/X9+aFBPw8w9aV+q2hJ95kUY5Pq2AtG9Ere2/1an57rtHfZtIHxSwr0ql
2l0v+Jp8EGgfh4HAl+R0ulE6KmlCNhcBX5GNFXMQPFFjmWiUcAyQGGo2/fl8AAYu
QkDR5Jl6umFKqt+RTkVKT/fDrn68ZinhWBDEB8iscvOjTemOoWwnJAANDSgKRCnx
Dqs9gVwKl7c875RS6s1nEXrM0jdUNkwW5YfdtLaRjFzcj7fyRALS8dE857gauOzf
jXjYHqmr961lQkbA/wJjjCyF58w3Uj5LDYg33VjyNZ76dBKUjZF1bzdCg1lnSlO5
7oaQN9j+JGtwh/Mh7FzZzCMm0VnNlK1hbWy3yh19tPGqnG8OVU16YJv0E2DWiPbb
RdCoSMev6cjXezf/7ohWLZy46GWjJq6evWsBTtWOlfme0xGW4GLkkkUMDFpf8kQv
NSS0WFrVAuVKmX/Tg4Jc10UXj8y4NFLmb+CixE0B0k3XR2E5IvJ3tOaBIf1i3GmL
r5n3oW8YrzLE4jqqLNYf1cA74xN3g8saKyYMD306wizo0BUnJd+wdZCrbCj8jtOw
XVJLwDFhPMTjE2wnXhc8efy7w4HNVCLyexWrnuRQz/XhJmHMmWd8bFkzO6ulpl7M
jrf5bhbfnEwwsPGJh6eLXPRWsWJ7lEpcfKKYpXiA71czt3KqRTFR06ycsfZaEHVy
5eDDGJ2KIpeaMBkHDWL13tQ8JSEvZ8ITN6KjG5NVNYLBrklotcfqY0DCLzokuTzH
rcixJMsX+4esvU8YTVYoOPmEA2eM+JMwfVZOV7a062f1+R4O/CvKiKLSXnlgdFwY
ta4hcJwbUyWlg2M6RzriU8JfmXuS6vPRVAiEtOUwWZON7K9P8Air4HE37l5lmLLc
HzJVBp57eHEAAiaMsvF7jDSY8fWmJdrwEvRjxUFNRww3VPRAjAYMYocgamQ6tGsZ
N/GnP6hmIWP7zL+VWzMVYf9GlJAa2T5U21jGcMJvaAL5PwBR6U9KOiS7Xdph0V2R
+JpKWkx//hQ+Nnc5l5ODOnlA+RV0KpEv2ai8luuwBmV7B614iSpX+d9Tbu59E7P8
9Eby0Dd3CR5VdvW6vl1fR6nXiw4ayo0C3tWRQiyF+FB2I8sjZbX2c2Yxwd1hj/vH
Tjj2zcUbutTku5aVtDCHrsAC/Kv5MS53IqQxhdsYSSbKiM14EGOr4TH/8PDqfTxG
UW4X1JjRm4w2YtdDwC6xyA7MDy6//kOKNUauFh+grOQAVBaIZG72vifP0Y7X0Uun
xtfmvokDpowRVX62F/mdv+8NcdMMPm7kCoqlmLbzvNin9AWMS8E9jfd57gCWze/C
yDKL/d5xd0yX0vgu7eX0Xo3eY7eMeFqLcAZEvd++G9JYWdcjOWL49qnc8g8LmwFm
UE6zVZcZtpZBUdkYyWQntF2/JenrJbFfUm8Oj7ZDIRAAswe/+QuEdft7kffbVEbq
ihlYbu8GIybdFAZKd13F9hlVIYjE9+ZOYaEeF2pVbWWpI4ZFMNVzibRaHhleOG+C
V2pH69uMhJT+tLrMUmgxHFXIRw7MnEwS7PSVgG1LClsYsEqJ0i6eUnhuuDK6qjBY
paNVquvATab7uI4Dx9sJrHtk4CCGgMeMfeGZ3EcRGPBZVDlhw5d6vyi6a9kszJVI
l0Ocz/deI2fhFxXWyRKtlxMD1kfjjMyQoFTyQsT+XkfvRJIxKD5yAyP6cyBSmlkN
tjDIfhyUIdP0h8pd6UyNLEZUb/969ZLJbrZvEzgEjZ37uxDRGUBVwHZ5hncF05n1
9ejQjYLGDSEQASi9+TVpRMKcSpJ8vj8vToK4/PHtATfQGFY1bqaHCG5wMYlnGWJr
eZdix8s9FkbrUo4ys9+B2vUUZBMWCrUTh58MTstFvKc5qyJo8rj4CP/eatPlAUw6
jcACQh6BpocUKqGTQgkohE3uDf3rN7tXLiYOPQ9pp2kieODfX4xl/64rgKozAJr0
o6moBoXk2WePR7c8FX3ppY5YdwZDCBJNChUSVrL7PRPyykHdugs2shkl/aNbKFt2
+tRdHNJBBARsy3HvKxOvOJitFbFGnqaa79MF+IoVZSv3PvOcG1NpbAaP63GNIAiV
9u8H5tT/Y8XsIPvR/OPBa65hIibqIPTCnV0NeAOrXVMHMQUI+suqpHddkP+K+4LM
srIabfbIeWxOGjTwXwDqyFgrMcTo63CG/4O/ZEriCKTof9SpgsPN6NffGo93oEjX
LPyqDUEOj36KmBkgbnzlvDJ4Jrc4nw9Gy6EvhRvJOULgXB9pHJ9F8pz9c4h0GBoM
dnFgQAA1MuUOerg/66scgsbNV22M9dUuRnFw6Znq9MhQwZ+emfyHdSM2YOnzNzpP
BAPydtuSaTIjdW9yJMSTX1mD2wrPhdTNYl0z7+d/8w7BIddblBcbZ535QbZvTamm
0S9IMxiAh02KhQ4dHooKokx+Op1PIXmJA7RB+UUFK31NbNMr47ouNlXdQteQA+Lh
q23NSA8TciRrXLe3RHit3EsmMRwFTMEE8Wbn75CvHk1jy2kKH4qbyrIL5C1c+1E4
lSNFaKtPAIwGr5wSMORZmbPbkW0Jy0emz9CpTXxbfxlS7Owbb3tp65g6t7AD9/j+
XTbK9n1F5sW/L9dFDTOxcP1AoCELLczV15Tc2bU86njdU4OF2VlKl7iTWpNhwN9B
qDoI5yM0Upmc/SG7TS//tK6mrPze1KoFU2EbcmmnhsZ7NwDDETzNNhns3JjSyBFY
VNYKZFvCZSnhCsjRgWWlfOAaDri/gWxHDq5BkuhAw1M9HLU46zhJbHFdtyRDBd9h
J1J2WKrUSXEtOi6ELXC0NUqXLiHL2z+dKygogt0RkHWCKXB3jki6Diu5Knz2CHA6
IufnPL0GSGQy1CWp5MQ043XX9Xox64odNn9y8pVGCxcW7Ojp4qLETAtjLn+HtE3Q
d1k4fiLh6BC4rjcp2U++tC4D5T/T7j5nOaeUNAQ62kMcBfrgRVjrsLUTy0wXXLcg
5V8v3/QSFlRmwuNDT9uwnjQDZWH2ZvIpP7gK89wgin8pLQ3sevu887u8caOSoY+F
poICxtbdOyoOxRLmRcepNelwSt/3djc7wZH0yoVOmWX+CAcXDyeomNZwE41746jz
mutiZirxg0efXyoUC/XJ9XGAZVtSRGE06CQlAFBpnF0SibbOQqNWxiGuirvX3u7O
A92w+5neq3VJ+m+bHJY+ecU2hyNtiBWn6npdv3s1Kmm7fv1vviUQ0dGjKDTXnKFm
Q5PQdYK+QrO32qaPVGdjEbH/X60sP0IL5OOLlaIN1DG6bZfA9yVuRQKhWPj+4GNW
jI8l2olz7oL9oYdJYOnd11GUiyBaOhOCFVIJzFScYIZhX3Ek92vyn7v/K1Qd+4bF
I8ZTbMu+v1mwy/vUkLapynIiwVyh8HWcQ8tHUn0MCObQ8l3HfWp5i/51qKItaCfG
ECAZdz6zefI/xWGosFE/8o7VQCCSYmF6n0zzmHbDDfZ/bfeXkj3QHQ85Jr2OuyT+
dDTBkpaMNjxkYCvJN14Z2nc69Pq4OcVll4Fb4ViKJZMK1bGWoFbP9CcjvKA/1dxz
Bf750V/e7nbR2GBajeGKWvnohsWUBdTc4CylRb5CSbu+h5NXYRDRj3jUicyJX/Kw
SLCg56gVRyD+/7fzkKCbgLLIK743qU7+KpUbzp6uxPCY992wzA4sDHPfxz320wjR
53KA6vKYiTyFuy7TYHTBgSB7HyWV3zRnPKBv7T5P8kCHgDa6ELVzfiWxxOj8yxaF
fFu0qrzMsa/gOTggMQCSZNFv5finvA4a2SPOeSaq2V13Y50gxI7hMyfc95tFIN4p
h8/ZpW6MAjPC/Oa8N9M66xZ0nCL0+3DPIKRS7XUhaSdHkDQqJc5mGSTRBHTwwxsu
BTjN9LdtVdXk5HEejLtD+Nj8EPVxn+lGre27EDbVwFmLAR1ErV9mE/Bf3SedrTTn
2ONpuK15e0ff8Wqmc1QYRgk7MmrqwxidjnVmJfU56yEpFSyuRuqPFs26r9hnVFQl
U1D7HNV/pXjRsd6O0HLvIFrIHHhypp5z4B0Bg9HEe8Nh8zHf3ReLCL/fA4uu5CI/
TLbAsbfTtJmt751ZM5EZwWe5bChZ8G/W7YDjDeVVR9Y0jRC+mVxWcswQfh/ku+9w
18MsiotziM+b3m4ckG3hPBBjoYCer4BibxH1nUB/orRUwgrpeV9DPE9RtYS6V7rw
h+0wsu00jQgEB8Ho/3ukNAI4xc3v3mT/kJMA3VsPGPYpBOO6ZZOcFia4xwRZeqjP
o7Dfpj8cgFw2LStS/jW+OsUTtkebx5qjrBB8ZhHEh84rdBPSDM/GVI4C6g4XmHRs
OCnwl8Ac5Cf0tz5FOpi4qEGbCzQoNiBiCfzxGm6dO7r78S7VOYOUNhjASO/+qFAG
hubFZgJKgVacufyoK/jYmpNhYUzZrdKCDUX8Gg+BizVwi+rk8AUV3BDQ6DPlnTJl
N9snD36i/J9hlq8JYWxl3eycbZPT95tHvFbexDazRT1CH/nBHi5eS0D1MSKVypqA
JL2xtQ16XbjZgrWOjSVnUCnz2QsquBX6lN4Hk5x6gw/mhnJSaeIA0fjnAiyLtIq3
QeZ54lpyghPnxJswz39VpaAXWVXnEtZwD6dfLQbGmOF98FXmNo96n8+rj+VjLt+q
aus65+JR3xDcUrU/QyvbJ9Nux1bTWDyCEsmPM9pKpQ8TzYJ96q5EbTqDWkBB7sSA
/GTNGY14NmG583mU+z/Y3RKy9olK2IYr5k3DL1Sbs4bIQPKLu5Am/ITg/UZfe6AW
24/V8o3dCZFeDFcjRwjHOMDnYjb/bhZpmRr+2PdZNQVvDOI9QcO9ZfTqraA3UcIT
vflpymw+EWbwFLnOMSLbVFpUE7kzKfedJX0HHaG3wxyDjXakF9rWyxuDexIn/7cT
8MLJ8jOZss55qkI4JLQ5nHz3UWtuJfGElGS8/GCTfqU3q63gs/ZPsfzkhzHuPEuF
s0zT9wNvUg8Jykpjxanpqfal+OxVRb4CmBXyy2GmJ0JmF/z9AEHSj4j50dDy/0cn
aUVA4HwvPY+nHgsURB30AQ8vJIgTpNF7hHemNhkdgp8VVGOkvStQPY6/2YG32bJk
xWLmVd/IX49Zid3jYBwRpv0iAwlmIS0quHlp7PDW39TwBfGbQQQt1dciWpNXijqx
QH5+BhCbJH6XqAzv2L5WBdKfmzDTKGKfZIsnG/k3vgh9S21S917PSC2Lobg6/lVa
xN6AZK60MfA3CRxZR5r0n2BCk3lJEFpuASwhvyzjPETvdCP9v+ZyvBwR+9eZIpRh
+x/y/RJk2lK7hl2ysMYnbMwdStp3jlkrFidSrDPA21JAPtbq+mbb1ym4ZyFxtnJD
SpobhGujeztT1SV69+CF9y5lSr2ZvSRxa2hitUzAGHYyReZKPpLR4+vMOhp9eyzu
/QwS4LkaZwTmEcMv6is7ATuy6mE8tHiXs4jJVm3TVOBub4d8HIYlY9j9qtH28RBk
uqsrUW5xHPot//PLXNDrbB+VAvvTfqAqA/c/THDJTvd9VGaBIkFsXPZ9IARm5PFG
xuXticT2noni1Aw5utzckFyEQBWsoPMiH912rs/VMbLafMDlM7UMkVRAUKJB+kj+
9oXC66jKMjoY9zyMR2GTvkgEjg09xdQhZjlIuao6qWB4UqVwO8oPRa9l4Qemvrje
xDwL+8aJO1RCqWPWZuC5niy8GaxZnmacu/Y2q7D+mBJmerpPAX4QJu/8DUko4Nyg
7uf5Q5zxCWc0r0uDOHLuNdDZjb1qifrL6Qd1pXLxE3/ZTltw42CV9d5rde+lLUPj
wXWc4lWyZ9YaSV0OexMRZwKKM2yUp4rd8Lha9FqzjVj/f81dKCAPtkdG/aA1prB8
0x/O+WwQYQTLorSXJN1q05j0cpYb3YD2iILV0ESmEL+MgcpLvmNH+Hl90qTC5kXd
Pt+fGz3mqaLuWdV+hVbdrDeQzp5TlSnZUnzaSmSrEIZTnf1LKPTJceGFrD1zPpZx
pWQEcRFoQoTC3wfR+5nsddzxPYfeHXdgEGgg/DPVXjZrpyzmlb6u5OtJNcdS/QNK
qcZ3EdU4Ae9VEMCaNYseS73OtXRg/YJk3exEq0Xaq3d7410k6eVo4s9+vCCehnHM
xSAR0FLHEW+tovIS96ttK7qhCSm6Me+2CF930eEdplWxcjzLNhmr3+iRJ7YirhhJ
MDjJgRs+i4CTp/qNqoyjkzm6l497W6pOPwpEajWS+dGszI9W3zpTNrT5aeB3JpAa
L6pXJtggQKu6lWiI7yiPehayJodKRJYK8GxGl2HGKt/gHMiFR/eGKp63tjLUwy2N
3zlhCwOPWQ7yzK8XbOhybp0npk0fN9khPMXNjwcVnXSkd0zkm8Z7RjINg6vDd8Pv
JF6TM1avNHJ1POteV/6Nq2HQWSF5MaqxBpT6AF0Ibjtt+qJzq9lqeTHYvS7M7jHD
MQ+2y4bS1+lyC7qcwo3eUaBUg3VqoR90EMUbEH+pzJxeDFETPMpf0Y9v1QktR1+1
OqeBHmPJ+j3Q+a4Fz6nRfiBjkC/eAvc+NJxUnWU3J3lSo6tXhCGcc4GK+GMQBgyX
YXVUuow1Rg/IV8nUD6N24Yu71jFGAS6nNrqzddHtUe9LvUMRh6OHohlRH0OM0fil
vM9I69JG4jBLqF1TNxAGlJldppZ9/b3aqMsVa+XqVovUA4qqtw5wk9uzFngf1Ioc
fB//8+hU8nxbD9tMcXq4KSeJov/vw82LMh8YtFe1bo9ExdvDxxm9ArCGqt0XRY8q
CudtbSViM1N3gBQZgUJix06hn9v/Ail+S2+aipz3/YBLcg4RkiUlvVbUOR+/79X3
mnaXjqezp+PT4qLERCNi/HDj0O5TmrRQyVsUyebMy2C5SgwXmQIGwffftZMGfL2t
oPFQHZ198q7zTPgxJVkgboZaDeF8BHaS+PGG+D8tpnGr49CNAOGkdHXKfXQVJ6BM
3XfdSgyRX7u+HpOjV7K1w7PlQdsus+/9fHiJdi5obAY0AslTY75iGHB0Dd4AVVDl
gBKqc3uN727eQ8oriHZfImMjl8A+uR9vjDsgo+nQ8qxeUEcRvWQ4SfLtOwF60v/s
gObOCE7xypp33FTOp8pMUaYFHJse+28v5m94H0gGYzjAUAv1QMKkhaIe3OJJbtq9
5FeSLrJJ7SukDopRkMwwyeTEwjYmEbY/vGZlubmP0urSquKRnEsDlQ8sCSVAl0W2
K/MDiK8X4vzXsyb0aZk8GaHW3PZyacI+WpTxQLrcQqwGe3xYpWUZVxQ4IztIxZuJ
ogNB0glOIHLQ1bBS7syzujtOGj9lgg/FXopwwo8PbqQ7PGIO8SkwrolIS+1vXoQ9
7uz7sD89BOQUFyJm+barmdPlIvWjlUVsCBD+dnWFIHVYPbmfcVxGQr86lAjYoC6m
UhlM/sqqiMxBBYdm/EFnX/YI+CfyZ6TjfnItNYenchIZ73Swa0bOjg4m7xCY/ue/
E5lXClpJ1rdIsnCXly9QadnM0/2R6YuX15NzEZBnO9youyF6kWst7DDcKkgRQFZG
omeQ8SKCvKiNtUsdZJSPuVncTe3oW31LlGsGunankzn94nmjTvmE1/JUuRWs5yjW
Zh9RHVXzhN+5jOz1+d7TBzrHfq1y8yIKWb1IiSJjw3A4JdaLV1UBFyleZHazKNYr
vU9HC+ZiYTkZITir7d9KdLelo8IG2gl+VikTkMtMQzKD/F8Ir88EhhsT0PxTCHYl
1FgFRHai60mg1u9YFfh1pw+/0qPVVWL+xS0079YPPa9D9JYUBIYH2p+3aHw34eV/
rjyINemJvfD1Qm/G53VWN7eBvQOW0K+CybdYBil7j9Js8KE354L+bvtFEWhqjJZi
iZzrOTmCJ4El8n64nMz4TJpO5itM9Rq3nlVoIaxSjBOcoQ03SWEFkuXXFU6rFrJy
pug1pXixsfMwxVgA3TYlsK8lCD3qii+6erBEu+Dx/eSwszxMlereIZGQ6BVYyBak
Igra+zAl3Vf15+AyyGb83Yk3jfmXzu0d0M/+E6y6yLvdmNy8WcqjWUuzjPQNl5OK
FXkL5nky0v7c5CLPd20iwO5/nap8yZxgdiDMQuSp5QSuqZ6y3QT8VQouo4UHzjiq
1tbFd4XXEZrwQ+UCO7A/KOdXy2dyjHI+Emhij+gr98PoOT4SCQU2PM2f41c/ojII
YEjmW+Usv71bF7sDoHd2/+qXIDbwAYlj8F2czc35h1hx3/XJpHDzbpoJoySNGjxt
j4hlIboAy7RL9RqnX0KmHlWJLlIlAQPlT3/nDBVlEKeMvCLEcBcSo++D3ZBO3eNP
yQCOIhjV8x3WbAn7E6XeQOrL06APhCribJmXTEkpcmz1WVdv/ePAsVhH0q2yO/ke
JuQNopvS0+7PnPs5p6fFGrgkjVjaBvmRhG9aT+Poyb+nucHcmeD4qqMYF8NYuL8V
9KRtxtI5NI+jt9xJPsTuXw66Jv+VoevT7nUGyknpyt4kMn71w0dqclRQoXGSyGYZ
Z3kdGVe6pw1P5xh0kPhFRtmc4lTUUZUDO/BVQUBNFRjMlQVCYG/OfjIt8sXq+xMX
x3SDsWKpusf24rYAUoTO2DNAsj+PZL3ROOESTXl57GW9ZIVKho+/LUY/dsQz8+L+
jvdb6VzUVMqSTin1DN4FwEWfp6z8pOXUe0XxSarp5EEM7rsZOhc+jZHQtmC/wQ3U
9epmui5VrvFinlzDyVexFm3EAjazrLKT6cYuc7lEd1VXmOgpjlVEcL/BwypfRVhv
rw36LB/f2PKLKAgHINLMIqSdWoq87TbxZZgURibO54C6G4jBMnY2liJWGzBYt28x
HpcIriQuVKg2RJtn4x/cya0MMHxkswiANFCJKvYD2gmfgiV0zxTxlB1tIgRBvT/B
glqQJIjlWRwrt5eJgXM/0lYmTHjuK63il8KrIcaaIpbfnLsXF/32Cu45K/qTwGBZ
BMpOB0qJ++ZUQBBN+2mybjFzDzWBYSb6jy3IwjJWfVS3wA6JK4BT1JtcCEAlvihv
YNWn4OTXVdaVPYB40IJpBgsyXIecUBDDGQGkzK3/FEZDWEEj2VTuNuxKEzx6T1df
Dc0t/NJnrX75ZPJ0luNdPWInypMXqiPTAfonbKg5oeeYTvErVVH09jWcMyMXivs5
qSQOxWymOlAZBRUyT7aMptiH7f8jW1qt1qRgaImcthWA+suXeyW4OUlFakWK6dL/
+To7e2bqhowtkTy6P3wUznfVuy7n9znIMi1qBR7ucOhWUyqAACGLSX0/hhsBVm2V
M9glkf9TmKFn3rFi3q7EMIiWCkg5oENvcEIUnLLEyZCuqHdM7GJEJMgQlgQtHjvH
fcv5aQOT0wh5LnTWxqMk7qDh/j0bHejStoX+VcalsauvoEt1HMDL4t39s7cF7Agg
9iljL8p1fTsyJZ3gWwwrZ6Q5tbmRt06QHn9iji0AHAvNyDwI45uQp5uFxYfqmno1
LHYNk9HCGndyY4Zjz+2CsHMGeA54EA7HiuX65STLvQPUkTlSZFr+2sBeWeqk9bYr
5Gl/uw+wi+sKN5JTriE7pbuoMs/FVjyqUuAxZOTLWytvw9/boO0OIgl+BW7v7L/C
8v2czuBkFYbHifBJtEYL0vih3/YCBBc4YAbeSeKC+WMOEg3md+A+RmEy8sk1HxkI
GMUXYghWzTku+BMSxueLFTeeyiVhUsjRw/i7JcQbRqTqZth2WMC7ZtmINLBkkSv7
7+ksLaZfwyioubFb2eJB5TWb6cDaEkY8Nblis6K2GIMaWRlSYPGiZevm4N4f+Hon
W12taiJZrWbVw3KDjFAoFHSlYya0Gwh8DXnG033v5CsoM7B8hRbJRvM/JiizMgMS
K3GOIlw6+T77aLZopMjgo0BYGX6GlPPoqEDb6Po8f7D7h7ncMnJIsSLX2APLeYPc
xxrpgxqV1Ll+lIucfeB6FLuSk520D3RcLLoQAj5Pa3nsdUWELAs2PJ05rC+/UmW6
hhHrRmdMKtLg25Zhi4lXXekeQNSofEKTYI/3mYfDnM3Z83p+PMmR/JPP3D/mc+VA
H+01PGqimUXyCbI2l1Rz24C0XPpgKidh/N/QS7EajO5I2ORoTqRochzyufXtAYeM
GfeGD32R106c5Dca6/xr3s1PvSmoCbjmLKOQf0VpHpf8HJWzHtC1DhwYjv0P5nUh
DtV3Wfzgzc+8JGNpBjDrttrmWxFeEXiitJyYqxWQEUw/Drfhdj3/wDG80xJGzJe+
gYR1/uB66Tmz4wmQwl7EQnKg1i+eHHsbwKmq1CsWyCL0wD9jNM8OCdCwN9YrpUfh
GytASld6H/3KSvxyjV04oSheVWFxKv26n/DBAXbuvqc6z2F6Ya+dmv7I/jx7eSIv
JJWIOrflG4rfI2qRpcYxbFcM03/My800qG69HuEpb3libdv2XzYXdAS0LvTF9fF3
t6Rl3uehiGYLY+HO0EPPorSKhmNXFqJVfdaLHyGhZ9NcPabOS2SW1f/jUcaxPM42
Tzln4FmwIcpaEszlcP42kKWpETi54TeDhTJoaekejmYjZ9orx4cww6FfCApkBUb6
+SH5ZwJmyKLr9efFSjkF17CzWt1Ujl3TkvnRK+zpJU/ZRVEceuLoSG0+kPEDEArF
9tOm37qS404sywyehxpRr9/07UpImFeSvYTgtLXzPzOVspehVgnHWab2Gxp+AkcW
48Oz8iqS7zBfSlGviiVUJb7N9guR8pTAI6XdAXYnSjRWj8kf/Tohhxa4rVyCDqOo
0xHCS6v3k/xThJGuOZBbrNXCzhUdnc/enUuwPjP3JWEYeah12VMuAvRIUZV9VqG/
XVSnXeWEOugPGUxQOsXFWMERgsAlrI0bc4CrWuU1O/U/zpdDabTtATpbUGUDeXaf
0YskG2kfM7s8UBOHlTCHMMURmk7Z8At/fP/abgYq5wS1Ye0cRwpY01rl/VyRqZfw
ckOGph8F9kWvAnscgGR/Yw9FYU/397zlCk/L+ZRZTNsfmaE42/+wqWJp+Ild8PZs
/HBVukoVqclIQXk7I8eoBT0BBBr44nNQm2zYVyy5qqS7GmN9kPCwaS1ON+fNysiE
UuWYjqqrDev424mOLKlfk6En/PtwjiVyReMvquvWU372Pm+yJVFvspg9jgPuTirW
bn93WbXMr3Kzw8Xp443jHPij+NjLpM+BKWfgFGzTYrE+5f5DEc2fhPSG8lFnEIWZ
RG3vDcMNFj9cwlreoCRQCuzu03yTXw+h3Y1WJVOd5t3t9PmYilB4GlQZ2dX0Ltk6
Axu6hck+RF78gpByBeLa/rcbqliYsOdnwUtldlsGMYktL/WsBfadMUQ+5bIscc61
Cen/kSVr97BOXIo+P3IjwKPj5RqsmGU1tBEHNtNoMsoNlt0c8NmdDe0j2WpdSzHq
ibRZ2qLqpIiCpS6uVwgqNEUEQ2qK3pAcw30LoLBgtB45Cc7ULUGNfYWx+ELrDAAK
npgcIR5SiJpodin+uSbm7VSrSgn1+MlWDlIKpO4uYa2L9ZpMegc9LNN+7QqmDjQ8
tA+OEtCcHg1lO/fJl76O+jFgNBqJsSpp2lWlTAc5fBVyWjym7Mq2wEQ96HovahYJ
lJkHsbHguqvkVmS2oTtRRJv1EY+FzNsLBzBf+nt94OF82mVYVqRu0Tx0KuWEsgk0
sEYPLLm1JFLAe1lsEe3VWQ7KDQMIBDSIDNH+2ZT3w0KZMyQyqnGbhnZCe0qsS0gh
IuDalbLfestBzvTXcHGztd0Wq+ZMAq/sBwWmBI+CLvUsDKBJXP/83hYdEp//2RdO
JFGmFweBHWyTFCqj+74SnKrLQCuH8CnTZTy8iWEqi+VEMEFrYXaXUXGMnzlsK53F
jxhi+BIj22m5BttPSCcU2nJzcFEm6ZGI+AXO09YqbjROcf9J/n5x7hJIlgOk4NLt
BfrxLGBrHgs/nJ1FQxhRLkv2E40qWdglD/cS3cgiLK2r5e4c8bUj530gabl05WN9
GW4RzEl3uzjcXXKOovhGIGlxISkoVviwrSIk5HOI3z6Qqev1AizuECtmqmYrx36t
getXiiG8BAUuixxKUxbtDpNirYAl/SEjJ4jwFPe50EWswqzzb7P6iAJWEmBr7JRu
jYkDkjQZXAloMSytKP9bm5fJSoa9PeOxaNnxYiqv1OUukyQNGdb8C1nmqR/2IegT
KCgITbEK4BqVnu8/TTP386wdT+r8sPhqYKy2u94h2FJPSTyihi0SgZ9H1vykb1Uf
upsxq07FaqsaZMEs+pscxw96gAMWCz0bM0FwnQy42+w/zkcGiAq61evsQVfUvwHv
LMO51dkrMvpavQkiVTqOldGxyq0Ofgr/Vstfibmh45/GBbRQ49+oXiITLWSqlZgO
DUIz1DdkvVs1AU+T2zwEuFGfe6xQWYEoJF61UC5nOqr81qj6Wa8bEL9MRrSRvMkx
Kh4PTcEpR9Y/w8Abo3I6lnjTgsGx7dyn6Nj4TT76Nd27cd+ItUm1ymvYpayrvQ8u
IxmmaGIOClWm3DF3ZU0AY26iTujK6agB3GobsUntZ8p8jrWOCkgmfsj+YXVU/ag9
kNDQToA2h50lLEXOxCBeBnF9HT/XejQ3PKvh3mH4+GWo5GyUiSFTBGuJxizhWNFM
hSV1AUwivgREBNGq7PmVg9CmzWVFKGUTxi2vdsSxmpp1y0XUSe0HFL/ou5wWdAl+
o7mfGGPF0N7UBAvpXll4u27TVBZBAZaq8uxD/OAYlPfE4elVb/SI5MNAQvIEGmb6
bQLnz0gMBZnvAGgHxpeC3w9w3pDmTHEo+8AHcF9VmyisERe1GqfBusqcGDrqcJ55
0lcKUHlaVwlBIrFwvZ3EIFYgy0ifyHA9kV1XnGDkWtxL8ZpOMbzOjZ+fihuSjdHU
L2hdC1ZYOc5nBYTjS7F2pa+C+gfpc0VVvJD9EbgbdDtArmMR1YdHrHf7WUqNPAZh
0dwSbbxO1E0xVMCA/LiVPEDkqUZNSnH4hSmSBszifF23NSN1jpGB0sHOMz7YAfGA
8FRGzfLwFxK1tD5rRb85DGl0etlzOCo+1mg+vPNSqdWUw8QqWjgV+jDyP/gmViYD
wE8R2lUeiqti8woFtSC9C7ybbFMR6ZUDBRxxRiMHKcZmr60EufBzzIGDraNZRFId
DTa6Qmi6jscVpAjAn5Au/uu9H6F7IEcrhq0zzESeuYAWlkAZ/p76e+KLdLQ3L3X/
XVla7Gk7IcbNKCyyMu/7aQP+CtAinMNFQYglGZqWjrUQ3BzEamiyypdpOZzs3UmN
XAiJkT0552vEHCAXSeNQOcelij+tyiIAXk81mZPRLthgo6Y7/R5sIpZx8L9eT+5A
JBkU2oFrdeqVOm1oglTUn7FElztvltkpjJ9HttyZVKyCFWRb9XfZchrU6pfXG39d
pAUSwk1bz38dWnghzfqnYbiKq9OIm6Rz4RCKeHWOTMVbls/jB5gUDdGiPzkAmxdj
bbPzJUc7AIAMz13gxv+YPYId5ePy3ERN92C1CqhBtdi/a7388Q0fcGiePFD1ZSyl
PGf8P2fqkGV0nmKoT6QvcrPH6VB721KDinoxCz5HCCK4S/F6UqU6uGqnjVCnHD5z
LIiZXh0s2xQE1zDB1YfONd+OI2VD90pEpZgCkYJZOxl8Mdo1N3jkOMCx/Qa+buAH
KegsDMoH9hkl0naoQXzqsYFIufGEYqJNmBYrVY40A4J3X9GBPSLlCa+mWFU9H06S
o8ZFd5trpNtQM1/UloKvL/yLO/oUFYeoeP2BfQMoTvL7td9xLj4TA3IvDkKw5+PJ
hcRGJKtizjMnOpAhXqWs3IDIKTZVhuPMEBLFs5EnzCKQPArICxwAHBgXBPdFMOyf
R67x6FhyQojbNNGVIhUstCOzPrQXo1uYpZ1dhaNlQ8++7rXpfcyxN7K1xx7Hk29A
zPQz9+An9AKctwfmV1WBwQJFgbZD7U2y1EV9ws7ej5KGTe0sA3nhBAMOQSV8XOaO
/x1famcyi3sow2cOBYAPh/6Dse78WIldd7O9YdZHMcSemeiPMrjzHjfuO6axClYk
TamrrN/Qu8rUJORXR0lzT7olcJI//WEIFGfD1f9gw3DrtueDeA4Bb+Lgu5kN3PJQ
uqGUEkgNdFtEpMnTi/oVOJtZJyzhcbIaIXEb/vkjaht8bcKb6TRV4oqfdp4tEgF3
eCsKEvPd28jvqejhmLCVB5MywfhQ9Jzd2dFL0ydg4lVILbY5s6Q5l58H90ZwswCn
ebmDvf1odMTAPJ/9Q5O3odZ14dd3rp2mrBgnS2nYxLmy+0dwB1dWWoYiDgxt8GpP
s0tZ8HF+ZX9vDsUunIIuw0e0Q+jP9Wu5IbA3Rzb6Z5Qw4rfnslk1wp5lci1iThEE
siXSaI/On1/1VdBf0SnwLZS8v3JocRuoJQFiBx8YC9su9e6KcPtA4tW8lEV2ctOW
tGA66su2Ej3hCvmpQAGgYestxsTjoKeU4IYh3h3B6OMHFsZSqCHWUWJ6iReqTVVR
3EOgKhiw0fM8Dt+jhx8iIiV879kwUkESWeVbZFr4EeTd+5iBLYzkWNmc4bfb0aLg
4P+oH+EsoezkaUdIMK8g7XTvshnlCx6vmpjaB3esb276WauL3trFhFMQ/c/w07qv
yH68rfbxGgUl4gPmlswHtQjgDqu/uCLVzXoaEdVoluv4cF7NBNprZ9UX5Mr4fm5B
wwB1bolT8JMLN4IKJEq7pb/FNh3nNe57pmCnhM9BdLn0/dMiMDg8eCgjBkYHphdc
CnXCQzcWs2YvqfVZWOzcciBUqn3k7fugxjsagtTk6pvclo9P/Ecq4cEgR82Hj1EG
ZW9hN/OPnRK/ws3DK1fFWe4vGw78F0t+ZslbMRBEWM2Jv1Kmu9LrQrFU1H3SckMy
Ru83L2GjEQ2fAsBDGBveyOwgtvjK36ne1LY3SLefaHXLGRB7qQ/tQTq2dTWNaaOv
rSi9/WRKSjpw1m8StdTkcCgwV77S3XZtKmpej94mctxBCD+aXUtcfmq2lM/zEn/T
3+j3t0Jnx5qabf4YNIfMA2rCEwRF3gSA2hx8NXxXMt1MtZvhshhsAfTxDsn1yLmZ
Jb32A7YRs7gcAQaHhov7fYhb8W5k87KgPOjaIUMDgnby+7fMElacsZPDDhUR+EOJ
Btsi0zrKt4d6eMwssH5mRw88dtGAn+JinNULmUXgR9pXbVKwfNjLjI0oCBequ5IC
PadqJIjDSM7kGN7xw2dhqafRM7c/T0NSPDRmN+qJaDUxZKqbY4OcXCdIpXPd34OE
sWhOjvCyqlXkQKNVMoUxeh2dcdcQFunnIv0oxHZxkdofyxeHQrNf7sioj5EcWCHp
Tj7zYr2gvrtJYET/vTn02jzX3YBBOHfI/Ky0HGl071HoRXfxH9xD9CAj6UCnj/YY
7acGuUhsuRXcykuI9BMcow6YJHHgBcc9WWnP332tAl3XY5/r2kGcM5M0MG4itK3q
TF4gVYwLfgI5i1d/S/bAGF76MoJT9OeboAK5iUu17+/Vi3bEeDDvNP1wWLRoMU2R
z8YW3oSLD8uwpmbJ7W+T9Yyrdg3uXmVneS9itM/UiqzYf/M2G8xsD4Spz0+z25sU
x2Sb7hNXj5eem8vfqsztFsQoYjHWVcugiqmp6/9c2qeyP2BR29PCySpLPcwUKfdO
QejSjdp/nkXR6aARtvSf3NrKY/UHIboIRgmCElNb5Yi9+wYUYqBgdm2l9ddCf4HN
cUCCNTpPAzarAwrwxtC96IPiWt9Uu9pn0Q4s8LMe0CgJrrcHHd/SNCjr99X9hq9T
cWy6T1tu/DqlL/D6XNdE7u7VSULvuMQ8crCHdDbUKBEoOFCSH+FwouIIxNehr1ve
kUIJLneCb66RYvNTpl/4/cYxTZGN7RYbZnSjrlMwRPO5jQPsMSZsWnKEhFMJCbxW
HcIFJPbAhQu+iBZLs1mWJMrbTAIaJtEfIqLi7E17Hfoljvvo2Ze+yWo1930wRj0F
vSnWYLfFsKqD3BsrFJs08IVCWunEf1IWA9Yg6gQpYEg0/FBHgcyA2xKhC5ITMCh4
st21btQSYYo7cRx8u/4bGuHHwRoVWMgGEw2nLyxnzm2nKiclWH+ufaNxE2LGqnnc
ireyCoM4/mTs5NpVviVjlk7s/RJ85LHeM29UDUGZbMkTBaIt42kscJNCIu0McOGB
z38hZiJB/65i6NcRFIPP0RJCw8quchgpGpx//x5ZZZDqLywp6/sw4TQBL0iz9KH6
0pUgGYpHnOMMzkMzm7ug2eP9mJr1k4wQSrEGKn3wAqXFmmM4fOy74AKdzzrceJ9j
aGMNHHkIs6W0Po4WGOvpzyiVJeLJqDc+oTxWZsWqEm//QY63CKjIvHs8z6Ys7ID0
ocjM3dMi2bZnwnAhSUEPHhbD8vzs0I9wzJ0mLaJvnq6G5Pg8/XWPQlMk14xiQe9Y
wLZqkteSKvHnw/CrAtn/ya5EGJVrsKAtEJvXgx3zOprnHiiRglFZ1+w9+793CYzW
Qg2VhNiy7eMAexETZZayMvuxbibyw6iPrTIERNoV/93k/GMZYpzg3uSevH3rWFol
enHgAWp+pLZuKsEvOg78H/ukspiU85NDNzKLIguKLpt899da2a7lUvW62H+nLDN8
FPzKneiVtcXl5SMQSSZfgXrc/RZe7xwBBnPt/JayhEuGo1PUvgExnALpgL1CJn+L
pmKlBcYXsn9DemTf9yKj1sEExhK4apkfFmvUOyC3kVZ7DGbzbzbRdpLAQP1sC4X5
huWUaB0YUCa8rxf1jy6oljFb7tD4jE0OEdjSWXcVxO5S/8nRFGUp2iNQGRC6Mv1U
DvxMGNyNCi2U4aErKIN/8WRgRs/c5oiUKcM2fO5SnnMQk7Ex5q7+7wa9SzWb0MvL
oEkJn5eclC/uoGdjN90a2POl6CFnTLhQSPrkjRX3Vk+MgjS1iDwAz+IS5ymaNeYV
9+zWIu0E6F7v/Qmg9+VeYS3CgmSEaMEDnb0ARNyfV2d7xnjH99TL1SWNk2gIT7Bm
CBkwetoBs32Sbaj1mwUsOGEniQ0uDwJZTxDOZQA9ZwfWwSbtBXSOd8ZbgevI6cQf
q64caHRB0FBUXeap3b7XmtYpJSpsiHIquWlnI+4silavQaZFhoZ1qIj2Bi45+Fkw
J1HVa0ibwR2Y1qbg5gcdPotWTbkmatiWmekg4Ch7M9bsxZfht/LXhuHK8e/SAeZH
ZnCjwFsFoLubCqAnSdEu9T1AgRdBx6W0xVTXOvePBfYAodUoOoM41sD9NyxadYls
8O/PakHdchzE3fSe30G0kb4kAZRUXuMYUZz0U7t9fTFnuQNKTqoqoUt/WGYBfJ0R
dRIwYcmYpuiIoORZJBzXzre4V0v4AteRBTGka4htrIAW4mujz4GU0rdyYzA3KjrW
lZtwapWkuXutG9in24l+nWuNQ4UNxcPIpY/A+bhoZNBjCsurbfqALlLVPqq4DWEM
ywJPLhgsCIrwLubS8eHAZz0FP9pj5FZuoZdVBdKhzLNbUJ2f18XZsNtGzbIt1bzb
HevLmW21+DDdnQECpK74obYnqoJVitk0z+KOe8wkXoo88VFeYjA8RoDjtQub0RaH
sVrJzBSu7sPLGWSjGWTBr52uCyGtf1vmaw7oA9X84poHW6m2S8abORCwsyjNJIUF
s1twrHOrG+7ugFnTOybVV6Glua1RMez8qyKbzOMVF1jxg42jsDmkgqli4asESq3S
JrxjczDcZ8fpgH9Pj016lcyTurXRodqMflxlyHz+0Ifk6PV6ZbzN9MisDY2H1tZB
p13fMf+7TBkSYWkNJwoSNY2INtbR6JXlFlxt7h8oscslsMeNIgZWFhso0+OAJA5z
AQk1sDyvM1dJhaJ2rzB3AE7gUcSYwP4RBEdyRxSFbicKVdn3qdEA3ULgD5fTVOVM
dO58nn7mEPkVO/q3m7Xn1P1OKw2TgRPp/Zsrx97fWBVz8W4xHeF6gKNhg5Lq+R38
nN97aP19jmk4nWD51Pnd9hFno7vGpfXVq4BMxXIeLdiOBNzVQnj+FWvd135mx5Xx
d+2K7MPF0yL1VQLT6FiCfToXxo1EoC09Jxug+3EGX05NftUU4qAm2YBQ8fPs97t/
Ke9WtiHjec3OmPCAh44YdOf0Lh9yuj+TsE9Ylmt64HYAoKhVCPtECeOhDOWfr8VI
NrjGXZoxnwL/Zysz0tCZkZxZN5mAKtrLhYp6JzsCeuxD4MAa4lZwjKD03jw+KSJ4
Nz0LXrdqFNqRcNt3Olhic4e89YtrpIWLpYJvA+nji1nnyp47NcE8641IEX9oOJl4
nz59U3ac+dhZYyFseXpV1jXjeH8ZRF/MJIvJmts45O5ayAbID8QJMJEX+RFhCU6o
a9idXIIB74V0ukVuQcVF/+YHKd7uzSzhvvKDejAYOHIlF8V1c0uWtEWuY50DVFhx
PRaa2+BEOcslb019Wx6pO35ozIe4+KJCC4IbCovSMX/J9rwOy324LDP8sGkMwUjV
qm5ExYT9CvDuAc28smpipVL4rZy7qGa+P1DbKxb1BCgloLe1YjRDbgER1nKhXwnv
Yz2/iWXBKjZVsduiyTjwe42bUBEQ1wITeyxp7oo8WOjHjoxVYfVqtpbUmZCX9dM1
w+0JKQENVgUdWAOj/SSplcXNxo5DnGLB8hv9dVU5r5u5AptDkNepiPCDQb8PSgTx
rFzpil+sYxHc+bUubFdB88M8KtdzABfvKYH/UHdS+oBwqBSSKBhP1TsWEoQQ4Bfq
KEdEdkwliERsm7rinREWiaRcnmPw4OV2O9uvw6UZxM1lCmSgjQpII9sPNfHs2aZ2
spDdnSCbRa1lazWdf9zgKztsA3A7CZrKZWoURSviZwcIEfasEJqIhZV4g4dX+zve
9mim1EzdxCDc/ZotUNLMQPTRIhm+D03Zss7estL8UQxg/hdTSvzf04DoYnGod49O
3A7LLNT4hiH+vEbXorKwrWDShz8XUdpGrQFNcrU/NhyIbPHFCALftZGyGxNDia5o
lJqR8kp9GK427QOVUl24qgZNR2ROS/TnYOZtkS/slH5OTW5d6H4q4RWHSuW6wOiA
xoU2RpiQ802NsUVf+l/hhkku+HmqfxKgmDiGITsOaqqDb3CQQ24yYgFpL4suxBUN
w+on3t73jux3hE6sTtFvQoKGyYkKxxeX3CTROpK8qJVqA+nsGPO2NDzbHwpQhy5S
lPr9AMbnQ96It6S/wmrumki+nXj/gKoPD5zyf8LXJMXLBmkMRdTftqGuJBmvJLl+
k0PrCE3iqXvriUymduwiKNmGQDcMEFD9mNn+0giTDs90kNUsZIk0P13A4i80n7aK
ieVZ7HKcNwvEOoUyhrTgIPRlMC+/VDE5BpKioKLMdeuJ4KtFOVaKpkt0cc7G0lhX
q91kknll0Re0FVKVXUXDSx9mY7Q/ynxOG5Hk5yvRxXANCZpZmhJzI+gdxPbHiMc8
kaiE5YwODNmy7XQwvGExwYOO775gfYLzt/hWpw4gkScpCtMcYCkKDJbCotl/MH2f
dzlplzU/LzlHsv8dNz3eyJoaUQe1rB4/ccmSFcBlBUHtOpiO1/fu1ydDLYI3koTf
pI0CSGUDS/KCl0iwiGBdeBcsP5BRDLVqslIMcPKt911bevYx1fel2XGJeZhC5xpg
V2ZpL91vucq4Wyv5psPpdf/cfaT10OTT857RlJZPDJGi/5O/PBgYhylAIiqC/r0V
LYbVPPtawWUdpvUNgkO94oahSH4QEnwE7t/Jzztcw7ZlRa6Y/aUy6UO7RwWj2Lj3
lN9Ivk3+JJy0RobkofIQJCiQuugJPkEyFwXbYANZNSJV9OrdruyO6iuctELxxOGl
WrxTxNEB2ls72iM/dMVkpGxERCMJvXUx98NyH/AmKZAglCmbRY9XTtl5KMagYkqr
MyVAvKFiM+DAfZpx//izpdc99xjB8cXfHF7WOPdH5Zyf8oQRdx5eSEfi9AyiKTjn
Q2ObvsWQ3r1fTmOD/1TjR9errqNeRB5Cn6GyQPY36HA9LK+ccsoDKDYMtSNAu9vR
4BAFvYH8zkh9qX2O+4o1P7yl4vW5bh0/RwSe1xgisZCEOglfazQey4D2o1BFmYeW
MA2XdNQERdJPM96CvzfvNtOdV5pM9sUDlB2UD2jaGOB/OisB7RUB5Yn+tT25Iwrb
Kxby6hUA1ElZ3xeiGghqAP2eWOOXn/4H4JkAZsx2x7ykYlSWabETLuYJnDwt6+9e
WHymsFG07WZoqKdg2QJ6vykGTGLb/4WsfykkileKz0qM2yJkCEJfrb3g6IHTbU2G
9fIt2Iz8zrBOrnVLuHHdtlNDpTRQ0RdzlewWrTFBT249VmGbJAn/pvlTRmDo9cs6
YuBzaLAP2KEnTftcUZH9ipBCBvoEny10pcjqsCfiDXafKdCc50s+hr5+669wrMGN
rneq92Ih1DVD8cyFKAfaPsLmFp/Wv4v/2ly3f0Zww5gp39ClnufLdVuxzVi9oAId
TcMprqaqdexRThvTmDLsNDfQ9UUszEOy3e+tH7yrj01PPKxsEW+G0JZi+KnaIv0E
7DfoUl9C9iUneVBKFsQTgY9wqGA8dr2lrlwpP94Cd4ly77vk3Ap0pAgaQM0YVTSA
drrxtSZoDHuQeTOcqaySKAqBfacD0vlt2LcG5PEp5Q7rRUFcPVqocj738yRPE79V
GwLVY/0wn6I2pM+VEgoZAr72qglhiGdTkUcWUN3VAgD+UsFFJmuEeiXCxUWrq3Ye
e8XklEpfdPfSV1KDkBU6pLjXjkrq1fSaykFOazsC6z9B9ZAPmq1ousm3Jvxmqrfu
c7Q3xMP7STBpt4BBGQoWvTZOQ3zbbmLK31Zo5Gw5ZqUoYhzFTxb4Aj34+mFlPZI8
eU0eV7bpLCDYP+D8XvzBWhtY6BukDEY3jHnJFfET2DbVqlFSPVrI40gTYvEUbSWo
an+At/76hdbmt78YJ459xmADZ2t510q3EMoLIEYcBj9TsUb5tSfAoEKlStY55ngI
cv99grXHQbp9nNdrH4FX73bzuoQn15eCcuTT0UhDOZPVMFE8QRPNS7r538Td8F4p
JokBAhaXP71KXvJIcpIrllEljicj77iIvG0obbofO9WeoYYqfiq6QxtXLRujTtMs
qLXsBNONcYO/RqQlUKYMe26qNFY6nX8wlAVyHHnt5ACbMbYpHQq9lkRnXj4umu2c
6xVHVLW+XiwwwKE4D21zINqIk/0H2Vs3LhuwSydSJV8bvuk/B1WTmWOpMgPUA7N9
JE88sQDj5o5r1ZK/2Bvs83/lLUhfE/cAYsCwm4mGI4da2o7pSWOAK978UkhpZJ9I
ba7jU9F8GWgH/uNw9rIl6lC/O4TRo58GhzelNvejNyFfimY9IhWtV3q86ShxRB7w
nMECTLR3iuskHz28pxkoGd6p9/OFc/fDmMtgBZFLlg2yPVgQpB6a4GjfbDExDJ+L
sU+bILDM5d2qod0yOXsB+tjS0fuEXLCky84wB1UGAtaSxHcKj969pmsgxSRttmAS
/yShuSF1KvDa6sWvuHIqiuCAxgRqDGLnifYcVlkvct5gNnfo9CheNmROmA0iZqYC
fHGCwg2FcXYYqptmUC4E1dWhmIDsyEm5m5xN8xJtPKerSLHM7q9xN4uhSwbY7NRu
Iu4HbyAQN2r41L0wmRgl7Lf14qfwQawQrlaW3mggF/+nKHSg/Pcsmbau2dknJ2lc
cX164iIOiAaxHQ7OFGqE4IxhP80/bru8+pUnQT4AYviaB7gCu7CtXYMP+NdjfPS5
Jw0BWheEkiAhcBteQg3zZES/I2O6MXJli0ti7XXvF03toVqGx3D5jy8uLm7mRa/c
qAMXAYEpE39Y4FqPR47Pnm1xjLdblSJm97jeIF0Z9mWFsqoXr56ExuCWQkg/Q6Gc
0MMDBhKVOe3PW3RX2QPmEEMobl6LWyf7hvLH8EdEkvPuqUxKN5oJn0P9t+rDZeX+
S+GwdKh+JrhrmvKpFD5ROKR647M0ikMaaKQMcQZrmU5ZL+34ZFRg0syyGHzYTZxg
mpB6tMCKsCG/ef07AWfOtuAESU4I0ED6fIzvlOjKFugDKGx13PAoM3HzEmZQQXcf
7kktzQCkzurvrAmWCxsFJdYk8sqr+pQ2qERsEwoMq2oEaWtPoKAaWBwyaybLYN4x
gxP2xdOiv292T1LO17yTS3vS86B1a0c2vj/3PsCn7JnG4ObwkWQc3b33WzW3Ec6S
oonsa7fVtblxmdji/00qkNuFX/ofVNj9JIJdAQupa1dOoHS7O+UmMqpnkiIXkKog
GptiJ0paw5FHhJfIrt2Gyufp4km6vXUZNvLQFzMnzeS/XJ4QVaMxBA1LbGrK+Bjn
qUOZGyHOaOkCcNPeoJb0TBVx8S6pNlNg0/z3pGl+QmpmW3vt+K+eRBAtXsw6GROy
3XnQJQKTnblIysDbTN7d1hz3q+Rysq/ZMbre03sSe1h0cmgjbRcAhm36jAGWpdnA
UnBlVNJu+Ig85wAJQFb42D0fPr3pIGbskG4BalXs4YeuCz2tmcD5eYI8LqZ5vbxx
sEgCAhHfSzLY8DCZ+w7+txYI5yZW1Lx/lwDaFQnfkzlacrImMrN5vgqrsN9ZW0+f
dHmlgV8GcRmFZoyOzvKvsvZBDXqnzSUppMesbQPl9BPGoRYKghwcwY49/6Tx3wbr
2mz2aEnUSAxT5MXg9FoarEx+H5R3T6Jj8pr1mHDvUxi+m52T13r2uKwpW5JXA/do
sk48F5KjAstssHc1sb70y14MzIJsoboPSFCq/43+OoTYGE4ocx/JlmwK8P0S27zm
Bar6ZBOK6LWk73/vHkCVRS5YMQQbXmUc/5RE1p2/qZP9YQnzgUu3i4ZgPf3L5qC1
RicY50NoC6FEZ0Lo06YY9mwOZxirq6abetsBpbtiw/zmpcNN4AOscDwDeGIH6nqF
OAV3d/TiFJMd9K9CKGpbluDducFkIB07jSak6Sl/HBLky3xFSVmPRvlDNgwqDpkB
qXtG3bYsa1jpsIP8XG9W2PsPHf9bwC6ru3pvYGjk/QhD9esPnr0BWJ59YnlsnOKu
jN37y3b2JkU8jYueDLXWJ2LpCz05hcjq1lIEoB8nlWAF/B3j9KdrGq9YuE1knlZE
XDUrespm9AMNpV4GJwGLSldteEJQUVs84zMSumJnRPD5k6gy8EQEjkgbPmu/6CU7
e1yUoxKtjFLDtCJpxv7/vB4saOYdLKWVd3bFw0+y3oux/3pwpFyyo743fhIhHRcp
ZfuTsFZ38QrH+dcui/5TrskMwDpbdA4JfU5Je14sDUHGWNaf0zcS53XRNGpUOq9C
NNs5Xnc9ff3lr1buA7Dw0XZ8MW+r6TmXkqzf2hMiT2Q/m07dZrScRn9V4LMgEHqq
4z0GO7R6pCEtC3/tq65sknk6qsVWfGLtMd0AOUfjOn0rTwmDat6TjOPpQvPeYaJj
yFcRsMnu4MkTNuSynXDh7SvXsr+oqfvyL5paClLm4fKaZ9gmCrK/BA/UQP54Y+9y
mJzi4ISuW6B7AjXlnzwhYDAhQj7WKRI7iWHJl5wVsnn6A1lpJ3deluEWaXvuGvxJ
aWu6rhepe+iZ+nYw5IBS+xfCpVkOhxXRK1avK22P+luCnRzIW7QS76u+i0+0TCUs
+dFv8di9dxzyrbDjJQmTrwNPTJ1U7wfxbNSCa6mSdiB8w3nwVXiX0jOhT05c8af5
qUU8ZOBJq9pBhLGndt6X+g+lLkJ7TkicvUgGQBBxKUEbkAUWBiwUiiWMVa4rC8vT
hLdSridabgCFz5CeVkB+DrAELXz59c3A3eJCURWhcIJ6PWsyCipMjYYp73J8k4RO
lSCl2vp8XP/IToELD9M+Z/kVmT8eiJA1EjCth7GWPYoZUHJq3l0bXUeCDJ9QgM7p
zyaHsHPC+urrbv18M29LbHLZnLFv+B6scmtbnLG4CqYPjXuEmoXEWnk6Sfvi70Ik
IeObRBYSIAj6OtOwdR4hZoPZH0bhATO4AsQtAGuQI26AI13DF/ddT2R4m8T/rJCk
RbyGp3Y49pXKH9qhpCcGXP3s8RWiC2niFTGGH22314UU/qjDSwbub3VLllCU6nKm
ocCwx987ljnFoiJDAOdoRRuhmH3yGqHyIiqYJs0Q3ce5tMd+QvSnLpIhYj0r/CTo
90rqr0vtUyZf0tgxssSiBhm3DnqkuRliTx5aYL3aOAa2QPLTD2C544eFRQF9V9ni
nvLPTBOQaTuc5mjmzoFPzuDj5Y30MSh2NF5j2x4RR1RZ2IcglfoNf8JBpH7VdcWa
doN5ecLOakZEx8moTWbZgx10I2v89n3rOxdZFujp0nhKULQfG9fQ8srSWSGHipVw
nOdek0Re2gWpuIEm3LZjaI6WhM8Uv/uOoYo1JI3VqWt0SsuAtK+MgLvO1bLQL7k8
/hOSBNI5MGZOZnIsB3/yOYDYKrFGBueIh+vUTwmsCBb/cNkAVSGmU/94XZ4vZh6t
nDLFaxbFI12GTMO/aCpfTlMhub0uIiJCrXXr2dMpg3gZWAmmEVFfWNlCvFSz9ibN
/xJxjA9Ajq8qDviO2cI9mltlBwOFKzQW6APbBkRLxNof9RP3sXUs8VicFAOYulpV
IBpj4UOfnNZvUeE/LsfKokgHE9ybWs7Sa+06wtYDLmnuiyW1jeTBanRNpaVLHsPl
Zm/8LCso5RTGl8R0PjjTIPnfVKJLKjdFHx+XpmAA9Rl8Ju0NPP9bSG3LsULRl91D
WRPRfGrGUgUed/7D0S9WO/yE6FNFZ8PGxGDe4Hvfru0k+XQ0LU9AyY3mbjTQD+3L
0UzRuAtbBIcj1yfTrAgIpsAPf5ZeFW4Xyz40cczf2PN4l4lQzmh80Tl50MQGsgjV
flc4kmtZ/qSFQx1m6ZZlyeR2tu5t2T2WSIa+mPQClvEjxhE2XLVGyu6IXCtbnPBR
P1nqruaJkk0EICrmvWhDnmYeTu4yGiXvrXUOEVAw6G01ragi87JFNGlb9jmM2qgh
7pDuk46zLtkwd8C+wNl0f3sVkMmmBm0qOqw/odShJ0/uDQBLbzNOFCx19A/p0Ea8
TeVyHngwz+pLHNtX7QujJI9B1AfCZQ0Bi9KlqbZX99hvCuZ7R8Oqv9gJQDiUJFD/
XmGZVYbSsQwHmd+MuIlRWKdiJY6zKsiyyUFfXXYTww/TB2vV/A1uM7GlRjk8tbOZ
9k/rPytzzu2f7Tu//uz/obCZ/cXDlXOeQ+VtEWtNjoIQGqiMOEzKYUdTNXPjH6cV
QuiB5SlhkdtBIfMi6kSfUZ+O0XsVw2AlJz9Iai0xIcUnT82c8S68zQml3jlXBChd
jM9tZEC8YQ0bSzbAxgLZyLpwI7FovsasIm8CVo5sYQRDMl/jieYhxQ/Za4O+mib1
tAWEeu1PUN2pJd7jWtSmRp95HeiYaiMz6fhzo9Vxwx+75UZGDtCQNHvF4TAFAI3S
+NfF3s/QHIrlxfvOafj6qzaXLwEvqHAlQAw3JlD3lELksDshRSG3NuU20iZbUoJN
/K23yWhreYB5dLlolTG2qEK+s8+nxMRsm7Quk0KRVqiSHXYetiaZ0e/vcO9jPXiK
t4h8xhLyE2kN5+k30OOj3gxh201PcdCYpJ3VTEFH3xRo+G9GDVWCUlT+mSOe5+KP
YSxsQqhzfbK7TYbXBx+sN4xWXjBwbLD7nEX5BwhVg71uMwbPXGddIlEtWmgLiNWm
RMJZcRz8eQqd/WUjT6VAdnmKPRW+0GYiakEjK2Kic8r32HWIit7KTFKUAj7hnVus
MqJplb1NmssRpIUGM+0M8jNKHMBnnE4PgzyI2no0yvwHiyz0P+ZrTR5Sbkw24XcR
Diz9LkLkrNKkfK9rvaM6OwwBUWqYkZVqWGQU4lSz4Wtk1/Fiov0K7qHrhlXsJ/q2
KNaVDFURIdCy1lTyK2e/jUpbww2Lv0ufIAx3G5b56Iw+EurKR1+wIsNxY42grd5n
WQGou1IFLaBPOgsEXVnxGhxP1Asn9BiNEMQFTBnjYMtGv7kLxjF9vyEqsHa/NT05
hwJ7panfn9msvBPmRcLyyW3bU3C02k+F387mYNoL4X5I3nSQHNkqblySR/euMY0T
HLm5omcb48yiG5Y0jF/2DcVPLxJOBPORBzp6vQT9FNq2ywesA6bye6PGd2cUAT8B
GBPT/T0bdcOKBqXvvStnDd0SJnF/17qipICp6pocLfuIBracDQzZjdqh8jl9wHNN
+kmynsGoCPeEYfGc4L+agR5fwOhf+sAYzkVyvmQP9I8d+OQGs9cdwkSWz/Y7B0WZ
QeEGCi8IyOWV6w8lz8G1wvvUkvY764qjWC+PD+vB9kkJ1txDIii1QflUts9Izigp
XiaiSlDfSCPerRunk2Z3OC3dAhJ2rVYzsIlteH1JkXhSdPXU7YqyHCzOjr8jmj9c
0TDzXI85IhlfNdL9Vt1++rlXRmZ9nHFbv5w0Btg689qT6IMgCWDxP15oIslELP6p
AhiF6akfyx0W3hrKPOPZQinZuS97ee47uq9tLO7dzOOBAM7bkVNKVtJd5ezz3Kpf
hgwiYawwXF8gIlUzsPMxcHx0jQ9g2e2WumCVm294aDypo7yKF2IBT9glB39Crhir
t38C46TUggoarnJF1TRCtkbGW3WTPEv8z6PWm2wGFOMetPj/aGjZAGPrAroxPa15
rBsKOyjuC8cKCgwqt1E9ZyzyKP/LSJHvvr+XcjIjDIDA7P4QbQJkhSYaVRLkt30K
W6yY2kvd4WQz0rAt2tA21/0A89keALAYqZVfFY5kwwAZdV8Nr+AxZlg/HvOdw19s
mmaJ2Pt7QiGbJfs+4HXoLYarUeYUXYACOXRSLkJaWEIKWwp12GFgasl+dmH3ejFx
ypbONku5NkZ9qBKPY9SAo6dg2BQUJrdaxfBs/MrPM4JSzsS8dedB/5fEgscD4Ft8
3Ea56Egdd1Cngw8p/a+6LyVYGXk6aOuglKV5TA2w8w5jlDbOvp17bI2HTKuQ2932
tdzB2REvcIT0YWxiIP8XPTLxYzyoW7yITw2xTxW4W1VnBivVHnELBm43f9h90+c7
+a/RWP3kx11s02px2XbWIYMi7J+Tk9VcKRFqWO+QgeSxFcfQctDkJ9XvK590xRTw
bLHIfy7rHbb2NsW7xasoJAXsUdSGDQJrFC9SH9tF0gdXd+PP587XehaRCv2uZXgc
DmQB1D5i5aYiZz+lSfNTpTFGpkp5wCmj9c/Ks9FizuzDwHx3yT+Hrlp9WCw9kVeC
YpKnKAOXCzwT3wmJlELzxb+0SsDJBDSCYHLjogUnQpqecXPAqJuIjmzs0N8vJlhD
gqaanWWB41U505JKn4neniiibjTqSlkIHPfsQFKg/0XzvJXonj3H/bfTsUnTNDHc
5Wsm+PnAsMDwN0M7AVadHG2OiB3JA5m5A2vtFayhLz3NZVqNT+cB0FWmB1XvPLPR
QAGerK5oDC58HWvK0HPKqyXNL65M/sy8kcb0ANYRVJkJgYere3sX1RNvwceV438N
YG1kulljFhaWdosRL+3sLg/PGoDS/3RlGFpNlBZNBz1HAVjG9sAgmmzQB0lHAviG
Sp15i3j06mkmfe1r42djQavHTx9w0u7c4G4Hp9DDUle7t4fzk9GM+5auSyljgHQ2
4pmOMeMETSjt4M0M9GVGkz4mCuXXfI1c9xi7T3OH8n+KfEwIzaGtT9KEWy0nEipA
C1qoGLbeVP3l7kKqq0Nvsh3ST5qBj/b2xmHQd0EMQpete9rvQTMskD90HXgivUao
MM6FsBNQhy766U0A2CDWiqP4wc6iB8DPFbCRsWn7Vrk/kRgZsGREVUIfW0T+0xHN
1Jns6sbuHXYaJ/8hCVhM7lO5xfdUSSIIhEjBCNQbYj5+OXq9+3GMvX6pGEfkNr55
2Y0rAm2zYMocM4KqU/hKV19dV/n/yEv+G6JKEbD3aKCVpvPaXz0lYw2d81TdNIra
tzbSMgyq8FXyZd0oxyg14KS60NMz+yrxgFJxqmhvfT1ZGQyCQK6B+Z9YFRVSAO5/
XSntFqLPb7ZKiw37VX3L+Jh4eUR1TNz0SvEkTStLIKI69flb5rs22UwaHGCvX0fN
hbRhgU1Ol6eGGzf8vjD9DTKymCUbPn17Jdtym1c/x3oAbxyLlv1L/BX+TvZOEIeh
VM9X1bH2anNZqvW9w17j2aGlqVOhY75I/dbm9rWXmNJbB9znqWGhUcLU7SThlhL5
+4rh323hvDowjmHhVb8qgofqv1Va51mAh0fxyZKAJ5hHkX6uW+7TEwfp0txTGLHC
9kcOWKh9KO+eCvy+aunR+Uza/adKwULWc5HVGD/o00Iq61tKloKlvZIxbvCQOdtY
faoM7twgioKbt+XEBwSzkR6ZhfLiHBkrI1Um1o7UmockiWT3lpY8eTX59mM67rzV
m78FraT6iIX6ENVzf7h4jwKUGMGNj5g9yixpOV2YsR6n+CLBvBTHl9rXYNN9m+XR
jqtSg5gtUD1ppGvHlSoE9Pakn0TnTWLhwCLKv+9t6BbCCe5zTfnt3016hsaZb5HM
sbH6Y2Whw73oaHbTKg5sKraWJ5HHTiX4ov6Midzp5nxCDoKtAL9eGi3kHeAn7RtL
CpiNXgVdybywqqCim8Si9u0EgK/ho2oVP6j8fHRRo9WNXJmgD44gx3AgefuLZ8hq
v8m6IQ9UNNfIdUqj9U+lGRdcAuM+Qi3Qzll2z773pfYcvxKwmE/FpSMMZr1Ciogr
tR+908cGnk+rrfwguPNN6Wsma9Af2Rgt0jn9uTaLxkxrSruyzTBPVSL+Tqcxyrcy
F+3kSIEJkqKXL0bnnvWbaURv37c032wsDm3abblpU99AR0fhJN3KzSFTR3K8AuQp
rEbmJ8wuM0RUoOecX8ETHWHLxTBKVcYzm1LYXG5tObgU7R3U0hu4LgOOOMy/3By2
fmS/v02Euhl0NexTFQM4gGSATcKnbE7+lphPv/byGIAQ5YyHw/7J2B7IOYv/VR5A
P0FWLT3vWzKq0DskGhkeuYlCJRhytIwjqI1jWmhzAjoUhlp94Juf46zH02yy1kmZ
7rXx9bmxUO31Kb47n0h+q8xh8ZNUPIyl47m5z7pcD8VYB0vyk3uB5ex2MMljzWa0
6ww9YLy0lLmzYPgyLgz7Spi9wSTDyRSArxCXSX7+KhKEVg1nE9HGopLgwy8s5Lfn
fpEdPqEwvtrew7eB6TH0WolN4YseBCLY1SsjPabJZl9iOwAIMJ0xQUmmwUaKXh8L
Gy6qUK/6f+lzkq5omXqnXKSx2bDy0/M4TDqrOhOHaTQxeZWhsmg8qjSwpdscIArs
c2euv4T5vRlPwR49Nv3LBZUKyqhc2HTlDKN9pJZi6JUS6iRC4+Dgd5sPpSlzW/f6
Wg1QZCE1MlSW2QYZUap1w7d9QDnWBKwPC5og4K83pr8+ZHMj65O2YY92WnZE9K+h
bzZ+XP0Kl7omDRTgrMeW65CGPIgKq+sNN547xnRaWXqJCLXKl4waARawGcLxgqaU
jEzfBfjB+GT0UjQ5VxHmmZKhgEE9WU+pQK8f1qVeKVRvC7YSRnzlhG+VSn3Tdm6q
IigxAvqyANBZkj0HrdlMclKyEZJhXL9KeUjuLVkeyCmVzAnzRgIx0juRMUqOXxdh
IsJzn3Ves5G5pGflr/4slPV6d/XuY7J8Ij5RydIddD6tmRGP9kyhPvlRs3hTwGI2
0azMsJNbf7hTO2pJ1RcgNxdgXmdSu60+dLPMhDBWamTg7byJyn47NFyf9KReb5wv
xDx5f1cpUcsGaFcE/0nM9aI1BRbl/BySEXnPDJ+xNWt0m3CG/8t5QIYnNh8IgV5b
uGw5shdmUKWF29j+HMG+wnlftkC4AJpdAcJ1FbqhUHjy7a6skmPZY1Kz/0+WMr6u
fMUlUbpKRFl3o4P4oMX8HIIL4LcNKWi07O7gq4tHKvi7EBIr2nYtOT9Ze9xspYfh
pchT/Mq1jM9ihlO9HaZ9FpyZ2RumZhLe785B7TD00w28aqC/tzlYr0laAyv1NTHt
jbM+g+U0A6LKNVcShsUJtjTFbMSa7pUUBqU72IyHcGm2v6NmDD7XPgyG0FgNk2ff
0gpKJnKCskQ2Hx8gr6351NCk4ywdJ5JBsGBDD3AF/zOm9YIAcPX+1QxVqJlnej/P
MPl6BOhncQw9jGEhI4Hqsw9PKPahGoC0OXiwA6Spg2RFpyOq0sq3LYxMRpGFojXz
1hwE+UBC9/Qnq7ILM+tQNIkVsDbc+EXcKb6G9xMyRnWpoWZSYdSTraj/c2vi+HqW
HmyT/fcuZd3GMlfU3fHIsrV3mnv6+FMkCcesII49UBgX6902Hp2xBWWARE6GOrCK
zzsH6G/8v7ycv+ltoG8pMK2Fx1RV7mWq5Y1uOqc3rvHKp9Ujp+ilUucY48T0Fsch
F4IgacZhfnZ8i78rs6XM7q9qNA5Rs7wHLYI85EPly/nDj/EnUPh/sX1HhFF2LdUX
vmYkThGXanQXphwfPRuBjLrCm9+LjIA868rsRZ6blMSvWCXBWHdene/pcpwOvIMk
dZkaiwSAIoskMYFs32clUaiXEu/reSIce7KXwsE6042XEfYHPJIH8j7kr5LCZbF6
8JPvLWWcdPLy/GxHWCMgIJZw9Vunosi04n0imls9kJm9aYKsGnSrHXYIHRx37S5B
I/GueQFRGEJoA93uDz8rAWVFYtgodn0kxmCoon+c1gq5Yz3unsIcaG3vDHKN2/sU
GHSOpCBfppCIxA+WBD3IL+Kz/2a3PiK9Ey6P3KC0r/tfvPdOL5rebO3nq/LdiP6v
2GeMUcMtvPvvTXhdymrFeZT9wH/Av8mC43ADpP5P5qX12v7cpVlC0KfNJZnr35nc
q/pjhoSG2tnHgJAW9WN9sJgtKiEJZphsdq+d5c2jaaud8SlescGmPSfGCDO4dp2b
UBy/Y0nYcZjmzmDNu0bYvTR2NGrWvGGN33fMU69d3+cjzSyQ0cxStWv7WKgM8+l0
VqKME1l+F/lvFu21gg0VybDINCbVRKffw1Vy2LXQ7IhYOdnHa4bQO2ygZlOSzoJW
vEgS2VivfcRSjNLLZI3H+xMKVwCd5Z1Y/yNa9jgeRCxPiUjq9hrHq9lV5Fr/nfsF
zw2qBzNdaaiYpGbflejSA2ZoKOmzZxMCS6EfNP5/Sz5Zf+U/lpSuhGn3umxxeTQb
KuyDoEhcbPdg+LUSALgxPJ/kjfu5hsC3U35Mo5hndXZYGXNn/d8Fc9Q77G1lN66s
k6DqtytkguHtflXiFRJ045v57tbKYd6eCGn1jiIkeOWuSfcHBUfQ9cbhm3XwavLy
EzAkjN+0/M1AeaXYKpLf1FRVZt7F0fF9BDPypnSJwzC0a+Z2VugkS8XQ6mrqReQz
ZO0MY5W0b7MmPfxJKnePH/XZRC0G4vS+N4QmEEGPDKSoROTLPdhzOLv/pyjVMMJh
AOhbSjpCsZXYUCkukb7d21ZrIpmwqqTb5P3X0daBbZ4hg+tToF6+Av8M9zvDcQL9
DiB0uQMPM+OOUBUbHnzq8+YO2Ilo8/YF85ggng90u8CukiO1esVll4T9/sFsJQrg
Ndoc6cHcPB20N37c9kqRFYzqeSCAPgw1WHmGg9Oq5+vW3QTG6fJ5/mkPAIPJ82do
edO/AXldut7UefkBUrnHJnveyEzNb4s8lbdEQTWim5nuyfoQI6iI/U67WYkxIRca
f7DUXzcUSsYbymy247hzq0RuKOQ7X4Lh3sZg1fzIUqV/ZK3ZeW6TRh8UhjOUXViJ
4P6xwS9tKweXZ0map0NbFUSgv3P2frr34fPM4Y7lgC0ewQC0+mSz9VaQgCmK981J
PZaeGiw+RxRCv4iw5bCrBrVNxj9kxFfSxKQmB/2f2b2pW7IF5nx5Ihvqc0koXHm0
AroDrQK9Z1YruU2SvfvYoGNtOU80ecwnaSd9fjl51+gsz8AoKAuUajbJ4pgdGMl6
sEh7T6qTFZNvdGKY8p/Xnc/D9I/tRkwe1PAPR9O9RZ1tB9Ue8gE1b44IdWg2oq1p
n2qlmdcXZL+zhDXDm+EdBgXrMcfH362TEK7oUJBKusf6cS7nq8lpiHAdpn3+swF1
QIB0CqWASPKGUt9Phplkcl3GraVwapb9B2cQ7Hzaul2P/DzK06L+q3xscWpNdD9P
uSgsYsVFN3OJSxiJxdTcvGrF+qalKI/lsaqsMIFqAJIe960J7aaxbttTm/CavODE
aOEMFTTm3BimayXhuAA/SX1dc5JoBfjld5FzNAzlFxa3z/Q2SJYUAjv7UOtKT7vb
PnrX0srrJIbw/q36QbIooRBEpInMWtBD0TNNn2ChdQ83x1d+iz5uS61/4V8jmO0B
tr3j/OxbyBuEWSUEDz8r5IgJK1qG3poNIvOIYccoWMYgJbRdnidAHPYb20BSbwcv
+TtxirsHex79VY+3o9PJYDRKYA3EJ2t0yZgBwF78P8LVpCgjKbLjONsshCw0uNm0
Kpos2g843MnzGuJTgy0Zt1ir9tQJo8zAcUCWtx4XuySvYvqXTNfyuNeKxZBWycJe
ab5K/lQ8tj6F5zqYfipwQGeQF6xavoLiLvcytHrYSWtWk5YBl11AXbyIyqVtQg81
xa6EMRPU4lQjFrCiEPA6Qzt+q68oNr9gNYUgNxaH7pxjoVBlokOWOyWa7TIgOFBc
eamH8xDrCEfOCma4ARFgurFcifAmylC0/Q8lGJ18tfO+9ClOLmQ6qoVOXlgUjfb0
2SAw/f5h7mnI2btRQd8vTz8PnG+PqJs4oz8VT0PaYM2GcEnTKYwz0O23zBtAU3Gp
ijIURHJ3f3W0wpGp3R9l+IKHpidedUzXrB2ID29dqlzqgrPeNVSI7HhkbqYArbD+
aZHonhuFY2GeQ7g7aunbV4drD+wYVsRk8bnfIYiUkThMXh4oq/QX34HeD99uZJCS
p8A4hkHLsZWhdIsxy6/MINm6jjLv+W3CCbmpXiwIx5XrlieAQd/NRW/zYuv9Q/yL
wKJEfoX186hvhXtYcmKHBxhGZviMjoekGgsYamqJ2IDDFEIJ1xA5lXOZ9a9lIlYJ
ef54Ts5myXWAAXffzy+VYiyrGHFR4xGpU3njCreEzd0K5dLiBloU7kAIyAHLPL0D
/U+57U9x0xRwo9+o+iyKsa+B+wqUAEVZQHn/s5W35Iz3OB9pXeP0sZVsnGQlTRgk
BEjA1PxtqmvodFvM6dfh6YrxjC90zegRocLnjasXW2K475mYrf7pqkvm9NbA83J2
BiU1UCJnGhzmTJFChCtm7PQS5vN/fQOcuWiG7yaQWn8nbVTR/iAdE3UkqGTJMD5N
T0nTHmo9xLKwqOdIqssPJC90SkL8/pW9o5KV/7tWjDdw0b9vzUtXeXr+e5XVAhG4
ptcer84qzj1jMxIzKE2aXcGTdF0IZNHIvW6j5Txqhc164nKm3Hfhd2mlsGM+/nzN
rgtHy1v2vAWATGZTRDztJNwWL63PcGsVRTdfYMkuPHCtPr76M+Zb19ALxSe3d6kh
abBYgoDVHl4AEkRJ1oR5heAKmPcAGGSshMn1Io4oOChPPT8q8OioUgpKytdW/ain
NX1/dCx2Rvuj+39jvX7LmvdSd8M8qUxw7n3BpiAQWbQiPejscEmsvV0j7MDtUz1U
g5Z+M2CAz3j68elJjKFNWjpqOHIreW62lG0P6+stFSP36MoNvdWGdZel43BRbV0N
vrtcdpiCRF/wiCrzRZD0uIC7T0Na/9fCmkNO+kUobpgZaGAZZR3PELCHOOhF0TLo
lBEUODIeGlwN6zkK/EejC0A6ZqAi2AcqKcKZFB/qbZijEgmJ+twMtOaER6JXuXuy
HHpVPIRx7v6tHEK0GOpfTzoEmb179RiO9cTHjvaeW29Jbj2WMe9T0rj+ZiGBMRL3
UWtstMbhjZBVZBnDWTW9ItYD3GQOfXr7WA8EFXLr2tQdmYElpvcGwW28J/VIQZqP
X+M+bH6GuPBeTaBYiUnOSLuCMI2MGbz8FvxpITPmZ3tRhXyfB6NAtuhqzws9ScjK
/LP39z+94UlDk63YISs1PUqrrV4RYMCm3wumPv5tsLTzMXsxzCbp5BSfrGJInE42
UR6FOTF3ojKMTCRUckSEu3JTgOmbJXQ7d/gM1oqzZ8tK8LJtylrYOVQjdvRxDUqG
RxSg+ePv9suVNRg8OPyqzfHqvh5A5jF31ZTlhfznB5c6AvYVq9lWYJLzJVuUULC3
kUpHx7Qq7pvrtirJEPG596DilVUyiUNkovtudKI6L7QvoAnM1RRLGfBUxGJpkCzT
XPafUvoTtBmioV0XAm7DrQHaOqgB3+h/nLMbH1I2mKuydUl188z3QRMByi0ZjMYH
szZ/Lnv9/ZgmXbjCWpBoiu2ABu057V5N67FExMFsJ96vGznnJnF6pF28gLTliWF/
ODGfcjt4pFj6N95XPvsfBNae0krmS0J7AN4bUpzBaZqOWChHbFdN4H5lPF2o0XEh
zpuy6Ca5TTDvWyx0hPEAoMjDGhtxMGPa1RnbDbraLXGL1MF4M1WWaGJ7a4nUm512
XbDXC63VoVffVDt6vwUcraIG8HQ2ATemCDkg6mBD5qOBs+nTQm161ZAMR1SO6PfK
vw8zP+0xibo8G1mqzx/5tJXum65yLpmfLfQdp4ljX8kI3n8sxPlGHdhBZUZ5MCJ1
zIX3d+YSQghuOR6GiNrISMHbKtET2wlvI66ABWjIiLegXvj4LmALH2m5wZLjUxkO
nkcl6wTTeQdKL+xMbHWu33KRW+nPrU7SxgvourBQ9kqDZ3nWbIDqDNEZ1Pkk1iR4
dxO/Sxew+j9eErXcDC09r5C5nsc7NMHxsvpZt4kENGYqlsendS2BmnYc/VYvnJJb
toaNTfM9GNthYPNnu3rQJRoRyf2qD1lCXhFSGJfbiKt3gMqH0stVr9Sy2OlHcxh2
t4dK567zJXY0GRiJWt7R3mQdmsR3zzroKsXxw8pHRA8KhdU5FQf3dFmvEK3rKA9b
SMm4bPfSIZ7WOnki8YNWtKZrH/A5OQPNvPDjIx5UCsI2z2bbinfbbxg+1Es8UdDz
GcFOorWyou3XOGfNdC0WRTeVFxa69qmN63eL6mVGi2igIqPRfbI3yKvEs0KIJGil
4bRocEJN6MHR8j7iNRDG6Wlj2QpL1N/AMNqQO9Cf2LSUcmNgvK/aD2kFjrr7/4DF
AHs9KEtz2/tdaXq6POVSqbF33Ufm3Zc+A7MZxvBRG7jdpgv+h3pbMYVpozkMKWrZ
Hh2P73pinwIpmSbUMSzUC4sEt6SD9VzxtIMWE6PIamSwRZ/h41SI8FJyz53PkT1O
+G+OB3tmO/A5whix/5AX9qsRGiGUpLHOhX13AT0RcIQwGUivKnV/pMsodLK7bOLw
qWsWam7E9yJFyk1YAzkdGYJjdV0nW3PiyyLQUAcC6EB4OSw2mS2vZ5Eqn1gpfm8N
EA7dBU8tOOPj9pV8RCUu1Xxse2nYrOjMrGHX/ZhRPh/ROqSTMg++eWpQaazqHL1M
jp4e0rQCe9p0lKP2MMohcUqb4hMUaxTZk+Akbcqefp7AnrqE/VrHHqtOgmjEKGjX
LtKp42kedXfprMe+azTlsQbCEFDc3aqNMmLHa2ClUfZkAErbIDZk4X7CKrpuQkm8
kNac3/O8B9MDExUtg9+ZmmuXjHGG5RgqNvQOHfosJFfTQqpaaZSc6d/ZYr3LpTk1
yf0BW0L7iTNqpHdYglf7JyKH1J4cKF0kM2erFvFoFHElZq/SGhrHc1DMHLQs7lHb
9SODd39Fy0P4DeMPDVgp4Vo4Ev84rEB/PfbuFQMPfLEacsf9+Ry4zDlBjqag5ddb
uLbqxxD5wEQ5Q1IIYQDNYT2oaq92zWhJVvBUlkJFY6bF9GhlBlvszYbqKCI4fDAR
AVivCT//cDgpnOjtxrDadWDVYGQ6qE2Kb1+wCt/hRT5QQ6bKMRsMIVs1wARYvYYm
Fy/paXj0D+bplqXRcj//jD7+pTmZJwR/Jbo64sp49VYNeCe4LwHvq8u8Gasplxyj
P8OmAtRaGZnjZsQxPYFfneHXL8/WIaytnDvHu4Sr9VglWtWh6ToGvwPM20aHI29v
VuMYQZHZaYhAtWwWQp0L0DiCBJYDJFtbT08IqjvFeS3ossos92ZXIcUVKPKqPTD4
/GJxE/UaPs+D5nB0bGkXr8bfFHr7lLMTfYFdHyKkmnFYGiTjyuEpYpr5fT0g2r7I
M1uPe+ML5ZFooHfoxfkuUoLKaqtTPA+2UVnUJufNPq0A7ftYWs3w7Btsxe4FdCy4
aCTd77oSeZVoAX4RLCCpNJ1C6FXA0r7zj9j24apaNwvbUEC2VJBIxf+RlTfYSEmU
vDGGiOAMo08/+ithRvIBkq1uk/wFwKj+xS65hNhpZTiLqLhTjEISl3SQj8iFPAx2
VfKCql+Hv+RVJhlsikBvg0VZlZeh3jdZ/W7kPYNZ+9QiPs255GxaO6cHGBADgkdS
TH5F1bbxYtAwhdW5ywQgBug49+gokt/F8Ot+O8od5AVd241Gl5v3MMZ9CQXSeyF9
JQ7LmrnRqPHa2zWM01ClF12z7moZW6tqzE746leoUtmqbxYj7bdHRr7k2iXXUJg/
RhjqPyJB+ngWiphWsuZE+4VJI+PnuUli8rvpQedet/det4VmvR8JTOwBDzxH3uVL
7NVRUbhvbSzT4VcdGzx5ehBvjHBj1+2t5lmGFLegilSGU78sSBhnOnJJRjvQZC0M
VyKpuZXYob9RyBrLPHv7iUlj/260vl1skCD5uRhjdrGbKHnAm/b8oq1PIQx6usvh
aTwkrl2VKJNe6YVBxeGIkxA/XcWjc3JuOu2IUZlbcu7OKJ6TaJnVoaDn+l2UYVFV
JtwUdyU+J8n+EUyFy5X2qjU3jQNlScz6/T0JGwY96HWE/92L8cdGyYDcEc/QkYL9
dvDiNa38Q9/XKeht3Awg+ckpGl/pS746Q4SpXExrnKcsQF+Ryp1LC5AU4YLBHVeN
FVNy2fk7t1e+MSckOtyTT9NCMCBxc9JbTgAPeEE0qLnmvSkqn0iyNEwCjisMq7Kn
8hr9MBBndrBoN4ZP3pWrc1IlBGbewupEmeru51sOthtBrHZcN6mOqPkMvFNF/HsF
XUE6C3/DEOOIEiFJkf0w+vBLz97JRXFvT/NCjBMR4e3J95KN1hW4O7aNQ3nGM7V8
S9A23ZMpuKg3HslkVGwL13MNUpIqChGxM1HL2FmtzD8yHv8FGMUY/3rokmGfGuTs
aWbb+O8SAUCWo1H2Dh9Z8JunvScTNjQevht7uSiDQKy7ZAqc8A7mWLnsw6t0LO7X
ZxwC0xDCIy0JSHrVOioBvsf9xvkFY6+ykP36vjL+yfe7iARrWgLaG122lthihIWB
Q+OB6aAyJcJQJ3v2ffHZIPEIYq4ur1/Jfd0JrtjMFVCslInZqTYEn33p/2Rb+4gU
1tcS05UUFElUik6+X3i6SH9krmofENJh0ZnzZBR2qE5x+HI8LaZO1syLUUIeyJC6
NsrgwzLk+qF6l9I2PFF+iMYqpYhdnm7ieF9PC5mZSIdUF0onvUC6kaMhnHQHmeEs
nDw5Xxzj+chSnVf4rNnBD/2Dmn2wqkVm0lumIO0LeARHxHHq5TFNSMoUsMxC1ZXR
XBuMCazpO7mh624ca6JIJ3ZmZGg/fHVfcBDSyZVy0OyolGCpjXJsxO5KXqwBqCzf
62tge7I39fShoEbxVPqLBys/2wTseGbJ9cAwBXHvsS1dwHfQsXGYcpzAUHv3GyWN
Q1+bGyZ+KeWpULFM3R4qNRNNATXfAOOtRbx0vOHqaKr+esmHExBPOmD+k0FnbumN
/PQRw9ZRJlpAQ3abE7ed3f54LNZZ1Fhv8c5aBxHt1scon2BJvt8HTamb3ZJkkiYG
3FIQpwpxE7QwsMtLuvmagKhzPOrZilhWS4kCQixPecbBh2rrslMUFyAqx5ECW04L
Uc4wLAI7XMWpKP7h6h9z8f/83J36nH93ZYE0tnpI+qZAs03i87bYz20o+YMhnZke
pJYwoJLOh52zVZcsu077ZSMMTdJz9UNDmBiIHBex9ixVGSRsiIUhADU5hSLfl/y+
+2moRmYfAcKkFkpcWotM0yzhW0XN9XMgy6IOzU0aAdcrzVsisJYGYBOqdM3UsADF
SansfIzkFNsEUiq5futhcjBIfpSVlzPz+YvLy3p/c/vAejXxcYCxi0zFwbi2g+22
QYuyv7H0Mz3tUXW7Zc8Ota9TTWSLrGjpTeD933EMJ0DcyrA24KGVZLItSDp+7KFg
nb4XJESSQZvaaUQYeWxkVqv96rw4Ze5Fmgv1BPgcHjti0tzxmeKPayrr8FxktN9X
RPtjGJbab9UPE126PbdWCXs2SiAWictmAbHb5Rqi75u9nstWjSiwwGutjD+8cvBA
zC7iU6W0JAXJT9yI/Fp/0l0uN4Dxx6mbZAPRuABv5RUoQQldd2crucS1T5ZoZurX
ofShqzonfyX9ZH+PJpapIoDYl90wcJB269PE728BMCpTrV/ph57HDIYkYB1gDXD6
20Lq/zQrGDLu/j+MoB+ruN9NkN5C0vIrPM2q6YIkErFuJi0lM/mqo/tEmEgvoxW2
kjcv8ecqSNmVZHijv/VnCJ35oof2Ixi9vqGdJx9Sw4aouZ0XGl3fp59lWe20uXge
T+0HRWKGGTNPX9ZwdlCvYqhbp140oP/5opodrtXW7d3g+W8lkn3QdFyp/SaVCU5p
YrQckfWmqBXbHDG0htbDkmTY08dBo4kAXuEtN+sEAlFFubZ9eDi+JEl+Hu8JRhCV
TAjUmvt0CkhyXDFsGPD+X8ftZzeWYnpnev441VUnVHnt6CK6k1ATgaGQyIgH1DHa
P05qkw7gVpRc+WZB0IAZPcEGMbinussAkfYLY9QhF2goJS88GmjA1kacEYFMBuRq
ITZ0ziWaso0u59Rj0/GW0mNIeE90GGI2TNvSY6zB5ggMIB7ytTFizm1wwF/yUrcp
g90kNr0qlME47SOjny6o8qwT0H77p6eozNKPFr6EfyZ7OydJqDvbKKC1Sgs5+ClI
mr150bePFzajAJDFKGGklrXueuy7x1VwBmD6CjBzi1uogayjb8xo/oBtzSJ6DIU3
DUOcy7GzWxR3qlp/zaJZySrL9Fth2JLBzSG6wMbRTWjKoFck4tHxYxVkTy3Gwlk2
RG+Q/tPyu82ywhsEm1/H2rJQrVLkMNne7tyJzyCiL4ovvqmNgIY5AVKCG2whY9Uu
x+xZM3uEfb5K1PLjtcpKIAp9N1zQ/Xqp2WGX6FnVj6ZP3RDzJbvFHW7Sps38uoFP
SGCIS/7mwTHhGnBWgbJmxDSk06Oh+vsEk+PAnKYFJzddEPGyKI0+pCORBhey1mqJ
mJyreZPL0v3r+c8jdflE6AP0+D/JHBRAzFYprgtylEDAuua/jAPgfe8inDnls42T
F01Kng4yHmzB4sarcK+LtecF39B+x35MGhlKRXcg6sKSKsfhN3m5I+fQFJ0f3LH1
9FkMZPxBJoMvFXTzYUUqz+xUFk874EG5cmsiJCYA8hzrNkNU7sufniQ/pa6FHHdb
MKRKkSbyJ3l80YbPqVQHbLjxYD6HU33mHMYnXXG5Thum2wr/HFKGO0B2LCVfDIRN
NMOKBo39Lpnb076v53LX8Xitgvyw7XNEBYHjr3VdmanRVq0JEwkq1jkjRSwBQ1IM
qjrvxQ8VyWTEhw5jDqPCX20EWIIaIDXQ7CDULqVSqyJdItdV6YaqQW+NI1slHNQs
jc6N2A5jwKpEZCcNqyfMcmpU6oVgJW+o5AgSB44JtIoAbZqxkE9ZC0XZwxdqPwbP
zmdeCL08noAKpiyVcztm7eJSftgOL/C2tjWhDliaaV0Fran8eDk4aOzGehzqigYX
59I7w2bgDDp7IHiShsA4IOxzLOuU/vjYCP9fPS9A40qBU1PyCMfi+Ov3GVm7cfa6
UHHU8GHWCKpciFxCZmQPkAulmESP7vbGap8zgM10pg/WkhwqeR5NSLxwpLBS/sML
y34BiPdczlxaAv5+bWEQY77oGqrNrh28zkqgXVjFMx0eqv2v8N3MRJhHoisnoogw
mfl9jfNyOPDY5rmzcSx9JZgVZ7l1ef/aLH1elEalrEKhkhInImyz3pJCvA0sl8me
mVVDHZjT8QlfX8nI4BGEa9k+WFMO0myL22vkaX2patYb3vDDBSMN2IzK7GUndjqZ
kfv/jwMnmBFZlsqWBS3X+8aUrOxe2AQT0vxLYAuXrDbnDki8PyCRLz7Yi4qSicud
TkfcsETk3U8lanyRjztvsjIErdzoKle1jD97bhwAifMvo1TxYiwdZHfYy1v6q1Fx
kveQ82C19tmtalBAWH2zSfa7eJhAskqLNQtGTMpH8+sSiVzrmXwJOJ7QuFn2I1sz
EEAW3Bv04xMUv9lV9ulfHjNfSsSFdM3dui2sY7TT6qNtKtPScy9DE3tPfI5z/6LY
QbcGGmSJy7ZyaFynHdQzSkead64dnvQ+LKg+OQftV0ktAm2wUP9IOcZ07i2w6JAs
oCw5GJ1OY5oGthMLE73sNq5ObvGH1C1lQtOogPyQvBYTlpLSKvzh+fY3LDkihH2y
A7ciXKHUlzjFNM3dCG2QZQKW0DFMqvTmRJnEElWnAvCukTLC/4XPrpmUxLquk62W
Dhj/MnYT+R9XNLr5nkaaXznRE4s2L8Wq4JrjunHxHYmQEvZAnry8xwZTMCcZHqAo
RaW8tL2ayd5hGdr2rftSaqZeKQqvRAjBc/kr1G70tM23eWNFBnpUt3eLuZ4lE/mB
NiaILO9t/Kck6KL3t102W0T2wfBmkR1v3mxwFk7aJ8IsfBZEBvBHM++n1eXl69JQ
kP99eyFE+9I3XhSOTGs05Cu9RYNKjv9YmLCi/8WgwiiwPhoVeBG34RB8LKXWr+F6
wyCHoiVE8yMjiJ4l7+lR/O0C+V9dE3oC1JykibzNAnzP1hkkAIxPS6gS61ONw+/h
LzdLF1URtmRnePvwR6Ky6w8048sZYa9oHWm3jGx2AP2DiZitth2PoqUzbWE611ww
vXoSrHeYNW9tjH/QxuvmkoxAUOAIYHEhwbdJilJ1FzS+40eU2VdX6m2nUe9LlzoF
HLBrRRPc2cxoHNPUHa4hTLZUfIcw8wKb9f3oBqCuBt7PFTF481fcR8Yb3OGRcFWN
is2bdooAZBsRJJg/7InGeZ8XMYtE4jlc8ti49vcgJ/hpN4ASODPCOyAZjraY1fvD
sTH89AUG7QBhuCkJWYU4zGa8thoBxCBvPyYm3TXLiEeETgLyo4yC0mpbiLAZyTtd
qgdGQ/liYeZ9RH8sOsuroZ6qHkLGcrb15LuA54+l90HnKraRAGXR3JJEoM6nxDSK
GWfzibhYdjHJAFcAlMpHL0qeYQm5SmlsVrpDcb0lYIYroY0i+I4zHmgb6gYY6axI
4KEmurk2qAH0Gcf2F7AHeW+dyLrfFg7IsrFmoTZLJsErC33MGqpSECoehRf53PP2
e9CJjnYzPi8aDJiL3YJqw/Wtqr1235PCXbyvJVN8MsTDU+rKVGjH78o/EAMm0zjA
K7SBBMnPwqcwSNzh6A8P0QMgVvMhSN1wokInMhEhGAFiKg1c02/2Bh7C/4Y5jpDM
wgN1LmvRgbiGv/sGh9IQqg0WiHEQtqyz8OWRnbJnlZG/hIWLSoxZE2cVtm8yf66W
BHsgp6HGpTgdUm64b8Xm5zAGx5Tyg1Ppxcj7EfHvZ71E9Pk/TDCmXngueFP3jzH7
zgzbL3YhiyB3ti8fYGISzGXKbbNdPsKEt4MJBMF6tgDdGIXJ1c15AbVUGZ/ok3pQ
6qXTF3uK/ivqTl+tk+OleWWZOanIEOjXVBVX8BAaBo8N2aXirnqQUIktIDHwhcUf
E7rIsjVnm63Ym8P3ZTPBp3ggsdcIopJFPAvtGtvArD5dOqeZNlfvM1+beJPdtcRQ
m1D/xoz8br1aiL1duduA8OJmZ0M5ujwwzWBJKb4ThrQDIHc+z01due+2hYgCUXtY
neamovgAHQP8gRJ0grB3sGYIP2xzWx8H94jrgV7PyVQwCI71O3m7CxDlH9OqAioM
+AkIEZA45Y4Z7iqye3wQAgiJFmPOgEJYpYyHXI4VJ7kAw1pSx2LqzMjVQBWrGdMt
OwN+SG8wiWs2EI/qhOP+UG8M4dJCJSVNYTYVpvUZERVbJQirsAXGgRRKDFNoEkuS
IFd7PnRQPGxhyeEoRULRtZ9zbze7ow1N0wGVSkzT1bHrczl4KCwLfO4kEvoHT2yR
ulD6ACNFEOv+R2BMwuKStS+1ztOCk/Z8YEB6g/Vc7LVtkzlKCTzzYLWc9ScULRrk
tX9KnmQRBVDcIB3PD7u8mQgvv58s0/s7RfkTYEZGVGuB8e5TJZLnAq/eYGlAxlS0
rNKTdjOPiiXMkIOfzBkYpFT6MhNFZMOyb4AXE6bN2dzZAlK2egIiODTTtQTC+fZB
O4R2pLPA/VIVrTPF1W1YMes0Xkd6RRfgo8V+2K7RBDoLQXWwwi0NVsB+QWedSpdB
iw5joHtKeDlnKTDXrqHUUmCcTmQtztDDoqiSjzHo8Gi8gKcNIyUEoCqCczjwcjD1
wqnMbWUrJe9e8Ja22W26AVhlgxbFZs+k+yuw0IflCnUDcO7wN/CfkGoeOcTl3CwT
MYZqxB61scWDcwjQHhy7YSKShNuImcu6qutPvMvUraiRJ74vNyONfsPt2n0hrO4Y
fn0wFOJRafLWYP2D+eRltvt86APin7Sk+9iYfoeumsIEKNdztUbT+YIfcv7rLk0C
Zlt6t+0BF2sXj2WWe7HWsQRllQ94VdW+xXEQD3FpUVOWbEPjqi7rW8jRdYm46xsZ
ik9G/muLysHuZSpLoGni0w+7Nnm4LLKI9YSrVCvAZXK2wYhj3ejiN4rNarpsxoFu
jsVSBm0J/JXcIAIIV5wdNyQe/6jtACeEkUTPejqwy8jhKOlhtDNu03xnbaMD80c1
OYoOPmNLtlpLbaISWukVpkITX5jF/pxUasVRg6U89SrUrBT1JkKZAQestjrdvPZn
2NgTbB/Skxeb6jXEdMX2qskZc3cGP+7QUlQzIgI8zy0/u5MhcRxeDIf+WrGKa1y/
AYUgt/SOU+iFxz3tDeYWI7LxzvrQO/PP2U6T3x0CDIETGnQbEDzj35CBvgkWjbEA
xDHVZps8SbnrW9Qk+Cq7VQ+udbG3tCfqRaW87qdX3GwWpdVpg/phCm8vRexl5s1J
V8+s5cO+TpNzbbXDpFq+ZUylvOx0oZXgpXR8dqorBjeT/1O5axytUoYRIjCuXOAx
52FV2k4StWV+qg8UoXR36RkvvksyDXAbBNb3TFS8BvdfwsARs/0AUq/QSQpbziIV
oIf1up9uL+ShgHrJl+K8JvQ9k5AA3VKjrkzCyq4nfwX9HyUoV2QXPK3Omj3tE734
Z+hMJpLsICOluZ1zXTvpWdY1oQnE6DFvgZl88BGSyLSgayLiRNNn033cJlUNWLx+
QQTvwjGhBG67J0cVZGr+joTzrYYBKd8EJO5BJyZVj7npU9EXddSljxR1/MTHS/Q1
F0eHfiYpQJRrQeyUdF4IcqnS/AUqqe8XMztgtJ+gyYCFFP5iF8QnnxwEdpvjdzVa
NEPum7PrIwUdsfVRfOv/i667r0P0v9BFn4wGQwpmdgjH75E4eJrAiLnp48cmHfwE
49eVABBMCfwzx1v/G+ifkBKqbL+RqgPOFbrFO1xoWZFCPZslJ5gbVlR5FuPxrEhi
IO+SPPmWnmONW62ejEfdqtSfPBNmcoaYt6lxEnDHkNutM720FxaRaUv6hPF1a3e2
MaD93ZujsjoFRP/RiJQFbPHBjhfWO0NbaP2Bco2JAtP9T9kEUKauH7C/DFAudSia
lh5fsWkQ1/dZwgyi1ddMG3VKyoeH+7qORJNqtbCSjpYg7ZxOrkYXdRjEH2MmjsIs
19yOFKHFyoK8ZyMOAUDSwqYFNZ4h29a8bhp+lZ9we7VxoEnW4yS3b+Yabv8u/7kA
5n2ebxui/349+rSvsuHEfpnZ42AcyF0hS9vrgzZU7x54669raNPXr8BiIqoI/1JE
ORYgDEo07uADP1w6H9gsjnihMH70H3VwcH+UkDsIQvxGny0wGusgpWhD9aWAngCa
qkfv2w0MjmPKaXdlH5ydjhPdDUTKprzo3He5lVKU6FHj6YSw9+huoPPvBH7N8DX7
t1x0OhwsG2QFhp+L5zxrkzEsD1wfB0OmYsEuzf2OntEOnNFFtaO63BZ+vvRQxj97
Kv4IvA1CxsD/pjMpusAKoyIutrMz3Y1X7MUvHGi2P7z++PIkYtzXunlQlPkA8c1v
qjYAiewsta6/vxH7F8xpZGm4vIW+/NvUFZebYZ6zXrv8UcqpdpP11dTBfPQY+T6u
6QBXSB3yCpXbih3zOr4rvCjqDsspgZT2joH4ZzpIWol8mGewFSpXqTvkTd4M6bR9
kyZBL176XfldhNV8KCWM1GKw+i9S3DsPs/Qa3/86jnaVEOeajdvAB8JYWEvTIpGi
uTsYkMMMrR4TZpill3zAjbLqq2eYZK/zXhA7zI9LcDElgLuN9ywGcX37W9fs7NnF
le+yg2jV5oyvJwAQ8cPJZA9gNWJH62ZO6p4qUPHi1HnLpRBmEXJxIenBOeUt7UkE
S9bYyvv6/DXqLnk7/fjalTik6cQ5EV0sIACCXmv8M63ZpqEAJHb9sikzCy3XlLhv
Ty6QBoAOEZaAJen8cx1ywL+FZarDP0rv3kji2uITTXmGAjb0umIabX5QfXhlc2n2
ECwRzhZFqdl4wkm9zAlAiQXYx/TG+tI4gsa6wATb2KG/VbeBF+ugYY6Cg5wwlksV
fQVAtf1+S+neRUC3iqHisbuhiEGHNyDDrYa95C/tTw0qwndG6/qUP2nNFVoimdrh
uaP+68XpGRDT/kwGzbxG6SwPHaw3dE1PntVnNH4pDngpSSYLBpQA+EvDN5q7bX7t
SoYkJ63Znc1nA7isfMNZfFnWcWnNJKUSSQzuS5VzpKaolNxcLe+w0+69yif6mtAA
F8GN8HuwrewvVrRj5++jQ58fTVk2XTiadWE1g4yhPMMNDC9hohVuUsB719g+UohU
UazHNh4Sgj/dUF8z9TrJNQzWGZzY+s+2XcHyuCz+oT/88aZaQtZ7/5mtKDd5f4bT
cx2pMFkzh9HYm0GvD8GVWUVZUNWpShx7WdvBVbaPcxIqhoBRVQMrbrW/sFfZlcHw
FUg1oMEWu65by+rBq050j0hN/voEX3o4NmC2gsjmXM/MqQStb3Rg9Th4Kgz8is0s
rFSKow7w13xWsnyNsgKw9JNz/jtmchVbxPhxbXSt8CfkBYkyKyykUcognD7TOhUC
YT/cBvajkpN/gzKjBdM+NkODZvkXDtxpqavxkt78NGK9YdHvfzcB1c6puqobLrfJ
5zot1nMT212wEptAbYhPVHUd2qSLlURFM7zNOUuIWS/8QDLQdZhPMoKgu8hBdA1l
FC8uuxlYtkXAqCLg+hHUFtQotq8bVKcA6uLZ6hYc4E3VVQV2T2iNyOFEfhBcUYqf
D39WUEc2nnxApZJp+6krSTksHDOCBwsY5xuolDlzpMAjLNJGWPPPJjDo887Tnzfx
OTN5JIwZf4gM69f65Q69FzzrI9Fm/pExtV4UsH6vYsrEVj1tr09OsmE7zRZNMhTV
AJNGFdh49TTO9RA0GhbbtDz86h6/IaY1jhIwxp+muOJngdfU3mNh/ScLH2plaBTV
w5l3CtqD1QacOzJs8DhFtWmnqefihvAVrt+CDjReuhVTdLAYA+ZBxWMDQUfUBYck
6TkPScvTnE0vouolJ2gzYS0CfWXEWDBBxmBmPsmLyI1jwF7Uk4eVxJxm4XlTbe6E
Jq2c1nEgHWkKgFfrVpFVLVhM7M3s13r6ew3hVwQrv9Ol5UWgXY6eHdpmH6PQjZwn
PJRW38Ylijiq+QL5fD0PUIpOBYLnSVOWb4w6li1HF0Ii/II91UE/j3aIJIwu0ndK
XblS/g1ihxz6/jVG+TcA2KstkWMxH4tq/cYKUhsdTzirxEKLgnXlb7HTejb2d2Hu
0v08odGu85DkZFcXtBLJIDwvcUP4E9vhoB4nRr74q8PfWlAbKv1ca/fhxmzQSyAa
XDo9O+Em7/ZMK3kmFykFGBe2yDtJvNCvTh0Hd7bB/bbqzAPIsiVd1kekcBBHJOGr
IVD4Fi6z0K5lBYR96zVKB0yRz4gbNcut/oANHtlo2C0lYP5vO6o3EhYVVoCPTDoZ
qdo+HkOHi/5X3FCoHcpBZvUy/kFhtxLjSRQGvBLqVUWPA8xY+Di3Bxd8Os70l5WE
PLSOkmiSCys7t5d7t8H5S33I8oZ68A1+21yTywX4JEe9JBqNCoRDVqp/7MOUsGYw
p2LLhoxMIC2/PidcMHgZnHeob5ibr070z1yLHIv/Y+8nIrhnI+149tKe0ibSdQup
Q56PfQM7o1WMhSxyWOU/wxdLQ0LVGNnhI81v6cD+mN9zOsX0RLQ6tnT8CAMPOTUa
V55W5U/jsjMZPNiuGyHWt/i3ezVPd/xtTgziadb13KzTzUg+IfQYy/kTqrwqUsU1
0STXP5/+QWFQY7HaSrBaNWZq0mayjjmMRFfJy64VGFk0lt7Ds3pDhPzPeRUMf6Al
Tcdp7465rIYes0P09jkFpYoLbmDWjRSDg3n91f1v1FMch8fShZdrIfjU8eHGdfRK
uSX1UUEHCXSLUSKtHQpGdq/n9vNMNrwf7ke0D8hhijLgDzYx3bEUda3Mr8S/7rWq
TZsJ/nFwvPr/5/kaZgSKYEb+Kv/jWptjZkN3YOSgnmfBexWk7TXmHirOly3Qf/bo
/gdYPxza2GEHLGjcwKxxbKpqVBXMRVh8cyXkU/e+Cm9IVfQsxxgY0J+w9EIkapOq
woWKKmF+ZEj2opWCXUzlM+caATN2XvykeIXOlQevxFPxYacILpvovoxWoeqBOhZj
YNN5DD19KL4t+tyMXF/ZKM++IylVaCDh/m5LHaxEZBbQfaYfv8P0vJeJJlmzW4zz
1MbCRk4uluqxzFya0SeK/CUmHKdDq4pLKFBDlnDogaZAFnlVP8uvTu6ERPh68s//
53zgs8FDN7szVKdzWKlVmbh3aTx0WXU8rFJhisK9aLB4JOaRs72trG6x7ERgtlUe
sl8ivgwJN59YMyYw+e6/kVm5GsWmpbxnryoDrw2zMkG6/AJpjbVzlaij1CyQEFMb
Nygpn9YFR0C+Bo7XA+I9jHE89GvYSTKOdHPWiQASxj9x0LUisHYtnVbFIas4Tm1t
4+7z3q2b/5uE1BIVqDiM5eIIbDExhxhB75umkjalcYuxU19riFnpU9pAHEibFy16
QS95cxcYS2u2VV1SWJPtdRTcp619zNHCwyaxP8EAn/4xA566U/aFgC+iptRlbVVB
M3wIQSDrAjA1vJSRMpy7Z16DzYTDuRUwMVSzm6IxpIngzIlYWX7+TlTvmHQsGFhS
no1Cs6Z+/wG7CSP0jtJEX3E0mdqFGSgs6DoAGMrdMUkV4CTF+Nus7Vo2cFvDwDaq
JsdEyQl3RcZylXV6QEdCX4zeiIQNM2iB8MNRThp/ynmy4fC4MEV5y5nihVa8qDLf
/qO8j1rc9zopz3L1FqpVOYJSP/p1wG8nKiGz1fyxWPKogmIQ3wpKWLZjd3X9+Nf/
xhuR2Cvy8OUepcQ7k3ah9XwW4ivxXkH9SigqKkUGOqvsmlIU5z7SPtgXVsGKgaU0
kBkofuq052PWwgbQSBcvPrcbhHWQno3h3Vjc6C8KZbvPI5Zx+lw/BokS7JYI1Ld+
cqQDAh57c2L8OIUYGV4LJcvdsEf0OUx96BEDqqJ/PLkzqb3yLYx7pbAsVLgIoVcw
J3sxcZNLStFhFwUBP3mTHJk9Psx51/LvCq5mzyD9eRg4nKMcGuKm2jy0whHogxPd
czhbhle2qX5Lb+sQaNA/9TqHmq5MkRq5X/v7XolkbWcE5K5xPAyt9fH6Xog/yRLq
w4wijZAr+A9Hsme2NyOZTekeVUPoKFHdrGye/YZClYgjGlRrrDk3KjU3sT+loOsv
87EV+Nsr9z81vydTpN0mijrptlONrbKIPbw0dGy1Pn9E+/hf+dLGaJvolaJCF9vO
8ENgAN51MwqXQt9JmkWmYocB/kpD0HOfrDlemb2Ir0uBN5tg52OE8+859hyfZDxU
cW9qHsB7mQcWCd9BsjOWHXd3S81Gq7/Fk1ka9IhlbdNozMoxZv6Qd6kM0Ah8JNPM
GhfYw9In3C/IqgfhRP+ltPePg+aUDamKKaaDwJ2OaiTgndQUkG985sGFm1BYUgt8
c0K8eBHWmIXzN/T+l4gTCbGTlv1MGlh+xTnmjlJFZ/UlokCkikbzGhUWwvglmaui
VIEIHYFUckVLQjrya/HVJGfVQtmZf7XBf91mtRAazXmtoH3cVmNmYKDS6EF8TY3R
MRaKSSWnHbcj82k4uoC4EskXP22xy3ooq6aL4JVrWQlGMwXxq7fSXmGjAqM6O/U9
75iUjIUF90iNxPgviofna/XE5rKsGTdVZJldm+qxvZzBXb0TkGMen2vyTuWF2DEy
JKq0NbRL95u/I+zBgrHZFaOoseHXj/yq67jTTrzsMz/HTcs7GNH/kDqQRScnwyJc
kgUzvIoSYq67a8k5lQ7AC44rnGma3iEdgiI6DUAriv/Fv36LClNmZI/yyGvOVEFr
s0lluhTsGstTZP5cnG0h4qLrIOKLOKSPyCnM6NjYgTI0PxLl/UzbXAL7v8zlwvCd
1fV86Idv2aapy3JX0LccBUylNOeJtlgpjsTz6iJlbEsbJjLp0P7bJFMsq8UeLApv
EsB3znL9m0qDeZM/XhOcBheuAmJduZ2g42ZvslMJxPnNrCU5ltLFTTs82aT8bGNH
2ZWP0Vs43DNUmpbs4YFuXurCyEijplcITg2G4q/G0/rOUWBFXnG+diHwiSWMCgR9
QRmYCsQmKWI+gDkYrhFd55aeuJzi8MGHETaFn8oevX4nVwHqxJ+CSBHNuPfzDQi0
18vWwV2GzBpfHHZwGrQPtXAg2Kt3YV1S2JvTo5D0FiDYPxnW21FiiPuY4/5gkf+k
k1nOeyQRnKU0XnX/FU6iS7eMtpiz4+Xb+mFUxhbUlvGgP++xE5WGEnRHYxp+vA4N
7oBX1k6o4rKy8Gx/Q4Spnyd6bCqUlB9LQE4q70v5fr4Cz+PCFxFpH9iVzEvJQVX7
5uesgdUvXBboBsN7qXkrmV4tc3CtDo75EDrgiu5M1dVR3CNMsXKKtc9m0Z1OUGox
5K3V++5lFALcnuA3FAItxM7cbyDLmBaN1POz9X0VIcXyqAyMk/bE8+nusSha8SKc
24U7QhgOUdUoP18RonFfQXqkxE2PqCVvoSnfduaoRvtbJlgn5FFcshjuXn6R1K/l
8ZMvP4AnApy02u4vbqoCloLE3lhE4yfZq9w1N+OP5vO4hBstDwnEE0v9Z7hmT6zX
F2l5qF+O705ImPtzATOYX3SvGEWxqp6BojiFErW9JeICD/Kw4J+b8Lj/X5zidQqi
CFFsXJyBHOuVmMIPwaf1pdZavi7Di40BZZeXNZuGvlbGfZegkXVNLoYJnya/ufYV
0vMizdBQNakMwyA+L+1vdpEcD13DiLwJqq3W/7wd0pww/QrockPiM68/Z2iY+e+6
vroPtbVdQA0zY75q+oUu7yN8CcyRhfRsRGtvj0L7dSBBe8LUheyXHCoDvI/EHgU6
ugJta7WI43A6YRBnQBGSLZJz9oS+OBPENN5m0G6IHb8ZaV+cQRy+fbHovtxNPZvi
nc6vXFc+sZBNvIGkk2dbLeLtYfi15adWhJyirEDgP5WWE9mDftcHtoKEGja+gR5z
l1fd+0ugllv9vMd2TavZAsymH41aAc/wCmHvaiQNSL0+Bl4mZuirjyIQLTK3MbWi
dQklt5zA0rokExc4Uod2XI4AxEDKqhFhmiGPGdVb0ToQjzKEo5g2RIbhu97sOYUb
IypQRWspPP9QXpXOGTG4hfY0qisYSrrXipK2A8sXyW7UkD1kvY3O/K9F/UZxlNQt
yJmfR0x221yz2hcA0YCAqiDKPnM/9JIW05YAlCfonqw0YPjdY/PuqdXHiLwrDgdu
d71yEkKdznCz2yt6cIDP0/0dK25MghtigQFBuj8pfHIhM/IrxLFYm/wEhIucMuVo
NjtU+RlvcnFfbdvKbMNDFc/7pUuqKFb/jUWDRq58tPb7s8zWlYhZ4HcJpLd/jj9X
K5aliioixQUTDrGIkowVT2AFJe8wkcfQ3X2T2iTw6mOYxno4orJQEK1AcMrLkAh6
WDFiawsIM4RWaR3E4OBVAVCYdhfewIHvlKd/QbwGcmPtYmirsSxjVn5RUhf/xDOZ
IpxVjpXF5K9XzfnBERu+3ueq7FizbQyE2dXuw7eFbcsL7f4qnm/Q6eQWTh0X7FCK
FPQjZ9uXeny6nsN4NrEgtT/HwQ/P/u1qyg3J/fYtU41ZjZW71IdR56eYYcKUrtu2
DQWDZChrgROKiuuKp+Fs+4aWL17enU6sZtRLalO8D+jigqv7bvH3czYzSZKYmWNy
qCyEEQcboqR/eR8mrLpQrj0pj8nOTzicTbP+ZjZSH7wMdSX7YWOToYnfZ2C7SAmy
pPqMWDQEuIjvI1Q1P+ZZsmYy3ousNw53mlPyqB89X2k2EzozbewKjPtYZ9aOioeW
aTpSR43E57NA+QxwK7MJENRZ8jDcyPLr7WIRfuPKZmLHgBRjqbuHMKZx5dav2SvN
ZL6UEwZMtDDcQCRyIWapxmSvt0r/y7+id35RZMe2mps7sFv/rHrzPtu3kAfH3KwC
SgYpFJ0OnB3joGe5GWO+EOR3WNJMkxQLKBYm9rbUAFlC8sQ5YOGnG+84WufhhttC
86fET67uWR/dEQvsivlg2icG6JYr4epPGnj/EVklBsnNe9k/4V94XWAnfIVxevoK
bdPlo+8R2W7cP6VuE38cXw5NfBQ6Ep9tahbMJqXI5yzwZ+TZNqP3FLCJnVtASTjN
w2YTPHAQ47g48A9aJXY31OuhsGBoIvp2QVqKbZMnggzB0ghqfaDwX6+E06WzzLlN
TPCNPBN6+byZ4I8lhk0girk4xsAiRqWUYvQZYgib0Gx3zAGbuS3d/292opq5rJz5
/HVtcWavm39l6Fp4Gc23uXioJaQ+6BdVOXU4s6JdluI4xYfD+InTsnnNctNh18Z/
wpSoblj9l9nQK0xK8JMCKa7is7yE+KdCLFm8AZjpxWMFS1SOPHi44/1lYNriPcpd
BcvBLlJCJsfbRQzLRZoNZsLYH9HsgsvemYfp4tfBoqme6v3V8VmMduWKmXqk5ul+
c8SIe6fKsxHI18KkMbtKYivikLXYOHgDJ+wuwQYnXkspRN9dk7BUv0umdxVbRJpL
emfOTw1R9Gvawmy8POeDlShZ0Nv8dtWzTvy4F1R1afQk7E9tfG8IdLvq3B+U41rK
XWcTC2JnhUcV5pRNC10xjTjWuRf1CLg1QGNCejFdYV7qRFnHBry5CMMLzzhnTLEV
6qIfnzuL8NomC4X15UF9YvNc9z/rz2Jqho7rjxaSzyPjhapSljGp6qG6BpxK32SZ
uECbTT4amP3BSeHMkhwnRLRJqYYDRNrLcwgYAHlvHLZ/5d8k67Uu2mAs0uJYKi0l
ZZ2DHypB2MveDnGx+DZaFx6tkM70BIsfuzyiFcHINH8frZVCwBzpJHMDthJ+djit
t3dHoiJDd+ytNVcXtDcXceB6Wmeq/OiRMYB6nPQBs2AF2Doa28/aF6QdUIxZZZK7
Hsi4LygcE8XitlbuNpsW00vvWDxVGXmeTLLMS227/TxRptKCF6vJycvyGt6IbhqW
7joO1509mu4e/da94yD+M0CCydMAQwEvo69zaKK0+Ivvg7CH0MTTkmDDR0ZrgyFm
Mc9QwD8dZyVfKQs7/tbuez/OTQCJYQm5YifYj2PIWUSmGyol2wasHKs1rh1vkEt5
+ebvq6kpkuspiIhnOlZ0L+OYrYF4MfaZrpNN3vf6JRNoADKZfB76QP3p/BDco5MB
bqcBfRolvOQxhK5K9uoVFGNLUs2Je3QbWM0DfFz4PiQ4v/h8cRItGJL7W47FQRXe
/b8nuat1NOifuRErV8qN/WYAJZzfiiVRHbzIiNqujdnVO2v71bfZ02TXGDZMnkub
UTHKb1jAnasanH1XVMjjFdAMmWCRLD9CqTfy3x/AIlWO3ZFZp2ow7OYL6MlFxM5j
dsMw38WW64xergAv0dHl6DRadThBVUp4wTrS+SJQPTeqI/vAcLvkwRoymo9rnZHi
V9Sn1gLPELXApV0oaFp8csI3yyB6Lalu1NdlKZ/EauLE4ekIHXkiyz5OcgXGNqdc
u+fnPeXLzE5fIqxry21JGVMfll1rfv6h5WMZJE7eodhgJ8EAz4SrpxXZ8fzHo4M/
QpcdeVVM2D/MmqLzbRCXLTB5rk5hcWqJDw1nmUVWqj7FG0nCr91bqSTeONKAB1Lj
R9WsVmWxLcZ+GnKlE6v8A8qHTEoKpGBpAkc+LSbyodeZGjV7DlTd8JMnz5Pc/+gg
gvUN6x/jElOY2UjUgQLulfRhGWoN+o2VX4aKHafsehdA7nT5r1p4TkIn+L4UOFLO
83Nh2qz/vxmWxOYRfk0lkdu9quzN+jyASMVK7AVrd8998jjxMp94T3hUiN6nWTl+
i2tmN9cRsQreAZno8titk2Q9PwCezA1SAvzALZOrfM79WuhERMGEZgPYQH5Po1jk
WGNNEA/XQFLPzaQdz9XqRFnuz6fHFJJQRIlt88Bodi8wnzx0/PrxDIKj+jGSDd8w
AZaVzGr7hqWKs77XFY11N5u2x+294i8L8kzFrAWJ9gFtbBsh+sL3wUoF3C2MNHhF
Hhm5u0fZOdiwMWnjGwpfBnMn1nrUXH96Y7933uNHZV4Xn4ps4oX4Qf+w24uGeDiN
1eA6DZkztC+kYa+j16yVxU7be6X6vL3X1sG0wGZon58fnaPmSuElYfEiq3w/kW8J
M0+Mq1E5F0w/Hg6QYm3dk5Ze1ebNYgQQEBXI2wn6IGdUbpdDEIMHLDEbq9f4ztKF
6y5pgKo29M+gXF35B2IoXSJviC1J2GUFCsV1o3ImHkqcB07oeSA7zntpie8uGpIK
iuB7+IgSxiWEDf+z5gq4ykuzL286epsVdXkekQer0xStGPfMU+XFToNBJgRn8RG4
kjcqWyF0XK1qVxI+bNwwkoE+y3DkD6p/hVhkMi4jt7iXZ+R9T1E1Bo8MiDiFOJHt
/5Abx2N40C0DFTt2DoyWDQr0rSfg/vsuVL3zlmu0iEbqJmv6L5XJFztjBL/awJJr
+N8MiF0q6CGOB4bZsy0dpN4/F/fmwmByfr4owTydMrHQGnJwantACYUmzMWHhV9z
7q3knfconqKf5CUNfcHA9gchDMqLXCN7rDfgEHGwHh6BMc5bsqKNE5dClzPyVdzB
la2Hq77vAwAqZzWK3nRXrLgnr5mmWIrnjJa3x11w4gYsqw/NAN5rC6TD59cbcH/c
1syQ9hJ+au14T3Zz0ROdzLdBu/pq1lgFzyCiP78rgEw41YKQ6Ytt7OXVA+FPR4yT
QqSr1iKI/7d8Hf3fZIhuz/GCeeoebu82yduyQEN4YQVdHoIcri6CYWQD7WpKewlg
c8IqiUX2NqhwNE2mQJy03gndSUFg1nH9MWcdAZ8nT2J5xOjUxL2EFPXFJml47fsb
3ZXK6fAgToWTPRKlXUKsbrId5XZ1THhnRiiw+lyM+1AhSmAAgKlRscYgo0XmDPyr
KuyL12l2v2DruleO2zoXX2YfaGhLMeg4PsYNVldAVdDPyJsnsimvjgsyQugQ9ehk
GO/IzA6xchgb50A4zvxVYLGdVK6FEeF7CCUyagdr5HAcELmKMeIr2lEz5Lwl5Dg1
HS81FbzJT4c9EHHYZYRu6IYUPHpus/efq2jxEVZQh2DmX+BARyHKYe6iwxXIowxW
alJYKc7uUDCJ+DF0LbPU0ygpt5s8q21LRPq5kFH8NNCPNZuSLN76rH6D8yj7SpMy
ta3+5Zxo2/LzwFY6ycokGakjzjiHKqdQoceQyWi6GqpHo9T4RkKQG6w66W7s2XXM
61mOtjQ7HIdseyMpe9uHQISIWNQ/J8ITvwDtlXmzrpTGgUXEP6qYOUFCGkEj1jGV
2Fd7lLgjw4fncoifP6P3VJI362EbTzmYJ0jm0VZktRy9vIesyLCQlOKGXpVZ1MpD
/aHYqi2y/lp7G8uOE2SongWPYchY/aqdLI1UFdAW3suGNk1nWe0T89sHDQZDYtRS
qOsVXYczoGGOoAfQBGU98dAxaScC+QLvh/V2WI+mjiSUVIwIw93OqchpzCRqX7h4
UzcdAMut7OSfrSGUPa4EiJWlywjmDNuxmtJMl1cB0h5GJ3mQTqHhLWXBR9QAHFlK
2ttgneBA979pGKdhIAaFionr9KRJ4v3UayfSZo4dyJTczQxW5Jk6gwmTHM5fRlLf
UrmtFbcF1AwSIEdUYr6XRPfJRKjBD/vJv0eSqhGyt31Yzv3gIybzH17iHXTmCekp
++UgjH2ADjMYlpOs2bollu7QhbJRTMy/MyLqN19WmkQqOaeaPgkG/dim+NpeErcI
L8dpWWBDzFVM2ap/1d94692Qv7fwkj72mHYGNPP4MJQun1OFF7z+YxnYkBN0MqxW
JDWmGk56RxBKQxfpXITcBVnE587lZrIJCqKr5kWMocf6IpCziCZj0hOyWvYOb7Pv
ZLn5D7cQI1IHbe4IkKz6/veWoBZQRru78kSrtYElplsm7HQWEECHqdrlTwYyyapO
ZlDGNKPT5z8yEj6nAaXD0KbBpEtrzY7svcxeBI3QuDu+9CBWX1cRBAU4yIt42r43
ZTMnesDYxdkCq3JDdz7df2tyrSy/nxL1YrXSKws9JDioQYF/Wee/0dh3QDsy/7Se
vFnH/TfOKUqKq3P3fGh5jx835rSwu/Ms+2QaUjcq/QLv+Hrgs+kSRfWgs6QcBphv
yfd2hpofI5ATMtFBRwfOOuydxC6BClsKaJNBnDuEhx+TZktkQmRUKaE1l2g9eFJo
gjEKGPJcd9g1J2AA/QZtWWzpTphwxMPvnvQzdGKPOenCvS4qxhk1FiBAu6bV31fc
3DU6nR9twDjRMIMEWRikiGmn86bTNlU3dpUtvWejqgSHQyiJA0Dm87P6oD8nTfWn
DHA9MsFKWUrsadL5TnueNZQZM+MUzBO1hfoM7NOgfZKeeZlwFYODi2FGNSjWAw3D
0WBvR7XX2UpEOI8MMWkse9wQLA2jCfLLvCzgrSmcmIz0YufstbiGb0gFr83ICScp
Fb7S+kRSjjHBKkQRpdzTCGJPB1909gNomPDaeO+yJqAs/0hzfFI9rza/ztmqNTFX
JFwCwZNCO9fohNy9H8Ejq1OomUbP4V2UAO/nyrVhkkqe67uqZi3S2g2KFikTc2v0
U0vfSKxEYGNwCbwFDLczHkl+isMtECwT9wD+hojrMkSa9/4AFeAep413twkeHJ+S
LE+Jv8loUsLk8VtvU7qmqUspR5/2vz0rdNK0vsyhxH8jGeWGBFZ1ECKzkWXWLIda
ujc/7KDWe1vcU5TyfG0n9b1rNmRkLi3yZ7DkdTOpFEL0gbeKWQpW0MA9006HLxgf
6DN7OChKKqiNzU8/ZUL7K8j03jWfK8U6SavpofrrTMBZ7OGDbtrJq8Bc1hB6W7qX
oi6sq6ke66HHJgbuxG+6pusfxz1NRW7/HwWFZp9QdvWSV2dLFsLtdx+UP8djMxeT
vXd6UzjTen1m/WFCPe6zdoe2uNyX4dMpzU8atbx++ZkcoGPVJBbBHVhO7EQRv4ph
jqnGGEimO2PecNB/qLExngzc74xjw+9+TCR1Hx2yMvyqcwrEy1H4Nuuf/ZW/XIh1
iR/dUpBFwYt2nfaNIUCSh7p6+yRNVt7SVjHw/z8P3xbrhoGACsrYxOXkyWimI912
WvJRkOSjZSpyPErjGXnEtgcF7Gn6yPF9QSzyntQOMUHKjJM054r3O/ZpHrCxARD7
240VwOY1HTMWFofq08BoVoY780vTGkkHoqquBY6CTCATfm6bXOwCGLbamOB1KZ+4
MERDJj0elfbWYn/h2BO8Q2VCq4yw4rXh/X0ENTkZSf/eUhg7xRhlZSOYVMxj8wHL
hPUWo+ij7MzClY9sFUdsJEEmItbETYP+DIDUOeUOc/LVtKzaXXEDmODB4ITW0CjS
ue7tzdvgYKvr/y+Ugvfz/kejqftfRTzuTIJniZ/QmP7CyhUXy1ZU5Fuju2GhEq7K
z9HWKWgT3r1hWC5uGZjdmsk0+cbgbVAvp2eKMnZLA4XtUqvJ2TSOUdNw0m4odfoQ
g9xgOpEe55HUHeX3Q66nSBgK/BtrQiMygSZLMdwm++/kRasXLiZzr02zp4cfHUK1
S+w1S460A7rui2c0UfEwY9cI7gjPop/Abyt1/GWbdD2GdzUbIv0DElxSQbfJJLjf
375xiudhCSMPLJZl3zZSbOaCxSbxZ5KkB+KJS5zaOSXMKGWyR4iq5ayFQE/ARNP6
0HUNXt4M8F8F9gNEwtHbC1OTBgAgPuULEaM4F7+YUbYM0TT7Mb3XGikTYUCI7dWt
zWg77PVUB7QGld5V42vf6YokC0FDpL7bRpuLogFip5F4vsfrqNZkDndI4JlLngN8
+HIYYl+HZpxxqwMedCQgDIsjkrGLy9cqGv633GjmknBC6nn4J/o+cduhwSDmBRH8
Y3HcsfCpLkCjTpSpZ9TRES+qlC+YEKKKpPBAkHI5EbuS3UeTr2N2hvy1x2wp5G4v
xj7vQkr71FL5ru7bOzeZ7MivTVXQCOeQhOt3eur6w8B69ufX0YMtSBi2mvFHW3Qh
7CQnqxGAy2HsR4wVDo/nnc05D97aNOorBe+bIHsY/i05o46xIs5dQQKambJg9sGt
c3lwLn1w7gb2v+wlr/XWL2+uhWaiFaxTijNRMr3sTHXCHM1p/KyWBgIkgHlp7eK0
TnOWqpwg2Muqlxs+Zve00IKcP3phKwhNYU/eUpAHy0jIi3W3WwzvYQ2Ck5+IEnBW
REsDnV42fGvYBYgEFgnxdGU+w6U6YQq+70dt6BPS7hikNS7Z7eRmEDNs8ZlCPt8C
rhA9e1v2aOtjWos5Wxrjc5Xij4qGFyTE2yN0H1aTQAnosLw+Vs0e+Gb2wG4mCG4d
TEFS+Ln0QB53TGKyGEpHV869le9g0Iy49oyPH2VZYBSpjIrHT48Ug+Z2lNEoYovy
00p68dkDlyLycuwM0CoME+CprJSA9reoKWgVqyI5gsUh3pw/nB5J3FxxZXHDVrnN
xzJxcAN+jB3k4WcmWaQcb0QEAkI8WMzkvWjj8mvV4j5FBg60wtRRBnKFMfmrZXYl
XrjsxXWLHp3tCW1DvbOmeP8G0YJhyAmv9L5b1sqZ9r+WdknrJ9SCcwt6rq6nYzzp
/mXbEWextrwfIr0+GL2wBAEWMs04rnUkoEmlXQg5DK+E7BAeqxM9S+cwziD11W5p
CG3VAZNoO/aoltfQHkPKCNSLuhFIHAE5mscnzuW3ttMduCmAwkNyOogYjc40UfCn
APL7NlbI0cbczLdJJnNzlCLSaXfvBi79wdTRUzNaHHn2NxBG2YxWYRtdGfjsl8qV
wveg137maAxBgY+mdUXi07utPbd5z0CDFWWaubNnJdyt11Tj+N0JBR4AGFnujdRF
ZYN6uYP++OblDh96r0RZEtqfJZ87a4yAdR1+0bdzFI7anMoh74lLiLeO3J4tOzBW
dJjw9WAVgJNU8SzY4GGO+HeAGiPGd/BCPGaxBTJGSyFOTAsODQc6SlT54QeqWACN
iC7W4+5LLZ2VSOjbdJWHkTH8j9KsksLcVevnURVS72WUl8L1+ShCUmdjypPXyKft
YxtJKL+E7FjKUl1nIe7ekVke2FSMSLydrB51DWFrDtJ6J6f2B/JGmzl4q3ZLHGCe
XtErqI7wt8ymYR/zGnZ9roP1gq89xu/M9XMN+r9mqhVp4JU4zI2uh/hv2hgZa3H1
/QjQPG6EORMnmQs1D2k9afN2Tm2KjCfpfWCdW6AXeYqwqJ8RFhD+psgHQW/nUSjn
Pm20ot2t1qJpBke1reIHsyJjfrYtsxjYLjD4wtIiJ8MYYXz+7BunqUDml3WjtZqu
HH3JXZf6kzIQFW9p9mTNWuSvJss8vpyZmz9AVPWNreSrZ8wlmZTeUkTAIBexQm90
tR1ODRH4eskcABiCEQlKwXZrnpUQBcufzRKZ98dMtF7kVimmrLaqtQPqUjfCuHPt
Bu3MNZNhCgECxz5EjiHqjZqTccyJUF1P6Pl7EqJU9kEHTPFrhVbW43HnVQ7u/KZ3
VeByQJt5VHtR3+AtqCDd5NKtTJWx/cO0CgPGa2EukvCLEeCOdiTOihFBv9F+MCL6
HRHwraO3HUI8e8zCct8nkqApIRsmL7PrrMJECoTxFWEOTLOC0Agq1+hKjrE+Uga8
oegACOizekQl3Cl+Ez1NYKMHl4etZ1uLD/t+/HnfnPKcdBAMIYaVZ2Vwuixzj5Cq
Zy95C3oFB4rZ5Fs3+kTGwq4sJtKaJAA8dLpdWPZqXijADdfwLVMVhhmmM5YKAV0D
o4Vb6N7uYSbbS4+sEi7jkHbyHDQzaKSeW3W2hy4LyBbT1Php2xfx1ChrCTWjoiQd
lVhPaychR+YULQT8T43kIRfJeRXb55tsknc0BorOZP77ZNzJfuFeH/A1TSb9hrKw
ENdSeEh59arBxfnDGkvyzyw4d4ASEzhRbKLaBpnqhdlOSy4dGwmsQokuUx8tMJif
EcrT5XLXLiYReMvpyfuhvbglkKU1qAXmyKKwGvLZw9+/NnoHTo/Df+WQwphGKfK0
0HFNDA8Bvz5/CPGbkUSi0Fhzvt4sO2KZLEKlCYWbcOKAsLyz8ihh8o54FgmkubiR
Le4NPDcCBKGOcjJpg3OnlkJILUmPrOwTbGPQDsWxvsxLQtGxJbXEskbMCHgSbn2n
O5a4MDd4ypmHkgf+nNewVVouefo/GRkr69WnCmKJ9LW4OVir9ZtCQxra3JrORrj0
9vWSm80+xt+r5oSvyItJpgowNFE+TWE/84TqPxMxhjqpgO62l0K8Qum8yemXvo2h
WMBxnIq+G4vWbX8N4KBBcDwq8WzVhwKJuYZNvKG0Si7l2nPOMqBsBigvaMyOBnQP
tM84sueMYjd0+GglH8A4Z6gdxxo9SPiqzeNLSQuJH1924tpc0xvs8HUbznFBjLJu
K97aqPxWfNgF7ZEEmQTQbRHLI/EEiR6VYDbHPFbxv+20DrD7unxN5RIyTVv79XNg
bFi6+j5OBD2S9mPqS9AdksUSMsdnG731XLPl4EK73FkIKbaRIYenkNav9yIckqSq
Z2UPsdcZ8e5VG0I3IErPyXcKhM4oE/HJ35lR6SVg/20GtEMwByba+08gcRQd1Og2
0jDXABqiGBAgksIM9vm3xfEjZS+ytIJ3dH6r8viUkzIDRhV+GvIrbHoFeWz3tQMf
ntvLyGm29xzbsnCYbQ3J3/Nr5HWDU6f5oNWXD9tA3YBUT5vnJRiiuXiW8DMCNUbP
R4M0paVSn2YGUrJGF79jVtSM/YMSM+TSVIF1OkI8FWcn/Wu0WMoZnf17Ggq95EIQ
mKW42EivUJH/WadWxNri5knDhggrAFmNl20mz0T2RW9/fClJIlAv8tZiJ6fsopOW
lPB8x8yVNBPm3ASzCSkYYE9aq0XieHUzVc1KhwEDeOLuWs09OxLErJYjniUZPjLE
6b0oP6As+e+71tik50xpAuY1w6A38fsRAH9c8tZH726oRT4/qU+ikUad9i6ItLT9
YDUnZ0ZwhiIB2Al6mQix4MRZ76tnL2SF29vJv6AWxu9usg+LzCKUoxoBh/WoAxtZ
qeEoOWGT68IicaybGGyDXXStT2RGlEXH/C1GQo6FhjWOtwyZHzFI64rJP9xsGRS1
DxCIJc/lbDWFnzv9cDFZT5phgCgW+sU5Y1RgvmVIqPeOVpSArTW2Ja5HS8GdetQR
8/HvohvzOohlU5Z49C5Dy1cton0SaFYB19AUl+4pSTEJFdgctXXyyL7BnLaVCNeI
nYngrjyL5DW/nVjM5/JssXVbp3Z9pZMiUEbu8Ab7WfsD/cN4qKmpEUWFDymkc8eX
SBhtam+zkRL6g0isN24Y0o1agAUxe3cBhOAgbZO24KCH4tDnJXNlsChlV+ng5zmj
2pIRivNM8LG6oUsuO4CNyfenDistjWmEU+yRorDLkyyLUShJsRo9kPAexPDfEo8V
WrWMsJ6VcnN51LGeowFrvwv/BM+rLpf9f1dxXk+x0Xi/JsWdCyK/feug6U1ZTTA1
Z9tF1vFw5XXNMhzgvRGYAtalGtqd2RDzWZd72BvJPeEEvRWczwQOeCFEJQYpIddk
EIbCbrpllOyYMizDdPbulRVQylBXhUWiKyq7V7tjK9k/vgYt4xfOqZBzEB+3Fpd0
UBfZdwxc7EtIyQZLcjUxWG1YqRdziApMvrzoBidBkevEZ2hnER1kIEiw1LZsafdc
MnIgXJps/q2jSzO28e25rERp8BFWZqYkri0Q5gmsA/7fNnCUd8RWSs7NM8/eMIGO
JP+KabAXS8berN8U/Biag+4czpOT8hDrdGa59wftOan/nBYhATtjOTfNzYc6cmL9
51fidWmi+cKTqIPH4iDGEtNeNzeaqP5eAKQikWV3DmaGahkxzBKLqah/958WJqn7
CfZwrIPCejncbf8gLdy+wbtj7HyOVcPZuePNMpW4cmwtC32Gk1Oav7VYa4N+P3Tm
OI9mGlzEQXszdSt/CkPWiQ0v8kbshhISfG/uS1VZ7Xsyd4aTkvXYJ6AxZIpNMIM9
rgzs2VXSUP2n93EkcGvY5UP4D44TJWifhswUJ+iu3DjguWtta0YBnRXUcIv3QzfH
Ek3uiy55zDT7JT906qHkU4HdNfEdAQMHCz0IfsyTVzOmcsBGap09/NXFum3Ck/oE
pV7uctRDssDiTT5XutT8CQ7ZTf0TX6MoCNWJjmJeZVjgaC4L9Pt0xthv8JTdq/rJ
qXsTHYW6cZzRzMbwOIBwKqmIsyJbZ8yqIjjN/4DSNxEqhQzSgsnPMwGJMf7/lIP0
LbPTu9Ql/CUH1MuY/LuPWn0KKlFuT/dDt9eSInXbYZY9pvq2ndtg5Ja4ZamMuBDa
MVY3k1FnUhJiZrsgnHpidm4+DfhLXzOQF6tAF959TufLzw5HsffO9Y5pSTzMl6Vo
ZW8nP3NEy+uyCAuBxB8I5Y8/gTAipFpFa/h1RWd5sgVII/oDOcqPgPccr8IaIwc5
+Ix0BI8JbUdfyu3Ox4aNMrqtrMmvQFCWpvfxP89t5acsSvuCionsqF+Qtd+BKfSs
/bz/jdP4TOdpMdFd5z3q+GNPGqazpa48dToUyD4n6Dw5dw+GQoTaCgH74fj4ilnS
85lhG7hs35ck/4cf/ICH7/Oyw//JGKsDQWbsrSBIR3ZCG+h+LXCkvPlrLWgMizFt
v+ZgGExPke48kBeYohygRjpS/rPE2rhwI+fYDlcpPhe83r3mlCXKQKKUcCtNr5sb
loUTsUFprwu5CJfGoDBLTJJZI2S1UvjoQHNDXd2lHjUO6pBWZLv4jUINHBloJBP4
KE0qZKzwX4s/0i8s6PyIhPZIQWKE9tSD7uNGhQI6DUo5tFxBxhQwB07ZdlT6qvt6
5JgCOqG+QzTYKN+Es2jbWSpMa0GUKwGhYYwMcHZp0XcMliGpCYU4wGP22fFWki6r
cnAjc1yCLaI+f+hk6QcpqKIqRifS1wgEWAwfekJXJYyWNnAfFgJySvhxOhB8nR8a
VCa0luss0aKFpiZva+a2GQ2LL00Lorh5TElpiyQslGtNAObAcfP11LABCE1KvbSl
CiFNoyygczC2NonQaFMMAR3Iz8sgS9vASmDG3YaofNJ2x2zlzc7uN7b8VW4ubIa4
fjRJVpnPLaEjHVMzzY8V1M2Fov8PTZzI1oXsqr76PUkNq4Y0R14jC74ItuGOcG43
YWFOvobyVpnOCxUZsGOkj0wckwPeaR7Beijp3ImVEdDc+zlsPxn5HvVhJjCmrrGf
0Ct+x2BYJJSRMkIwWydi/1L9Icnq5T++IHr5/wGqt5aBnJ61Tol10NOat12hBQek
N/skAtpPBAFZgluvsx2SY5SD2gsr32OVCSYWRMu3HfJFN8PjKSOSJA1oMh90+3EO
hVV0ZTHicwE5JDr2cOaZRm5mIh/ocuBPotQRD1q4N5xe/Bjhqs/T0ALNSSp9Hj2p
h5QbxSKhA4G7noNlVg9N2+oz9t/sPmyEB5DRL5XCoFOSZmqMoXTjFUsYTX2AGAzD
NKGLo7luKXbiuTVMRCivbI01WNTxE0UzSCmDPrXvZyqcqY2hbSzgPihbENJ6ngut
gjToNWi73oX/NJMJehJBl5i0NtYErYliyGMfOduXwQYUGtUQnBjkyAY3px8LF31M
tdvNT3pz1a55ITW02Mjyfku9ov2qtPQEHJvnxV/7p/hfumBTj6+iCnjXfvev1qT4
9wd5rRiEvCODFUcCHyyfTvV5gRTiDC42NqsxG32UTuV1ubSOgJW2dN3/izAcQhpG
iwpwSVs44hsYojyaIdYJ8OR5rRFrlwg+gwZVAnh2b9wv8ZmwnpNgyp0cMetId+k8
oplA8CfEbQ5RpVPmP6mvW3XvsFEtZ4sQXmWI2dLlqZZOoppuSKkP7vTy1sIcGEuF
axEcnG1Wmh6LlqBX5EYNJ7NPvyM96pSjoX9mJ4nEVbTM82o4U55hUtvaeWoYco5T
oVPY48EAR55DY88j2YAuHuXiDorbEmhBI3KEgybR2EG0Oc//soFJ/tePkZVlznYA
wTRwq9cLgQ3tv4NdI17iK6kbAQS+YhNCVPPY+aaWWwDRbVxH2UAV6MT5RQv+o20s
EIYmyGDMGfU8lCEh/jBZmJZRw+bFARBHA2rHQZssuXykw1wMvP2nlKIgC+tPd5Do
rBV30sj6BRu8+MOMO4bQdY/+zCVT9PhJa2t5rSy87hFv5h/z50cbjbyhZL1o08Rz
WLPpX7C1eQRSPFWE4ochFb1KhseLHvcEwO1z26aVsZ2xjwmM3c81TkeXzsoFQOQc
A1uV3tqk0gd9vghNxWG4nw7pteWY0ArLVsmfD71WGxyKl+t91H3TfHJrl+ul5DCK
FfiYCn3+vH+9MAiYlAh7FXjIMXI/dNVk2ypoyEKkFgynkHbV5a5QqyTxoCm69SMN
p7X3zvZPsz0Gfw7Al9/MhjjLkogiUmW9y925odzzT0JZKHQsvk8YQC8dBr/BseTz
HBTBoRMIi+QLflr2xclpRqflYkPmrASphW6tOBiGtgv9M1DlKVXF05zpXK3DgL8G
CyoHd5vZsgdI7E4yY4IpxjFNzYQHSJ/EHWQEIuTUDUyfnOAh5BHT0xTF+NwPOSBS
HtIOY9W292HGO1bN0xRNYOWO0Vr91HrfMzCYRZVuppCYaAW43k/LBaO7RRnMDUIC
vuf64ZAc8PMASrsDJaVKLzu6iK8nxGgUYxPWodKLZ/WLojaqyFdPv0srO0O2lckB
MwrZTivNANVn4xsphJVRbErafLHkpByMJx80OL5RvDr5Du+amcV4smSKcz97GTao
LKmMWnruK9o34SpFY3crC/wPkqHwzr5sigfJpxxqN87nJCj8rcovMF/dTx3QnDuX
LAUHZ9vs5Of7uzVaO6D8eVvoxfeUQiBwE6oetsSGymuT7XuM3RGdGKfHx9nIqz1o
436IlT3D7MebF6V8OKJbtibg42sPfsdrj3cU05VBSuPuZqpxforCslc/kt5oGj2K
buzRugcq+QF0jPu5mECjAZtusssgzPPd2K/Yj4lCCflEGHlbEjADl5d5QIj9txwM
ejO8/avhAeW7FHdCwX+5A3YJukUzVtS+POLU+ndvR/cXggdWPkS6/qD27F64AUE2
CDiHie6SWAtnLdxoNvB8zRyWZgaQJkoFS5N+t/pEDuGg34axMjjODOCol7jerifA
FwTbUMxsm5G+K1j6c5GwX4lnKgQlClkgAWrVD97qizmKQKRT8w/2zm5wndWFQaEa
JZPx8ppk8sHd9Vk1oL6MdKNxtJtGUtrENCtYMxSekGyJVTx1xXClrWdg3fuAcd3h
XxT94VXZBpJeurw1nt0WOSVYeYgR1g5aY+9CbYslPQIbrBOhMnqboJNrsSZGVFNY
kphfGO9kIe6pKsOMpXSg6S+DvFjJZMb48jcnwnhCClfYxU6fZC9Xh+ZLQAlZW5Ek
UiKPszMuFS7yh0MRUfObfAqZqFsnVolflds7DlR7mW7Ih9KRm96Qx5ljMsZn4plM
AXqbDKf1sBXY5ipLtZfoF4I3yKYSjeaYDPm4TW5qSKYIgMgQYkA9fazvCiIbB6j2
TSNwdbkjG0Lq63c7U5h06AscbemFXSFmGrvw3hnzydtKEj7df1+VWkeCtLQHkmTW
aZTlBlotteoeEUxpBotcPnbnm7wCDJ3PASMKxIwAIYmG3ti1JZsPycDCVnLKx2Jt
KwhjR55Ascw7KJFIKhw3Wd9Av7gQ4IhGY9WWuofDBVhY8hpSv+Ge5GNVgzRr8lgf
DrJSae9Z3yWppUCxHLSvFvcFKpmbGUt/pWMe1qzqt/9pFkYtFqkAFZ0h8rroYWqW
F8scm5c2CkRK9ZHenfr0uhdTxLK//452nwxYnPJsGsC1tx21N5nzvc8KhtpF+Bkv
ZNAEX5eL9qqYadmF1A3rjy5vQ2Pp0IBGol5EJ/lvNMQv2BxXTX+Ovns+mml2pPkX
L5zwXKZP4pmjs9/o1Wy+X5XcpKENnSMai5FZXSS5//uxf9wMLhGOZtFJDfp9rlTQ
wXS2FMB58Uwv7/qWv+usPvV1ii5W0Zgio7VACUxyyQgTH+i3X5GK9MuZWHrcfhDi
FrlWnyyZ0JMBJAZfhoK0ssajs15S8VFuOFm2cJGML3Tp3Um8xcKkuLd3QQZwykbO
O4vn0YR9yKN2zq7DZNBhCmvqzwXD3ODXBLKJbFFAlZWi1XJwngA04N/07YT+UdWd
nPRvMfe2esxkLSGNWr5eqaraMROIqR0UiBUaJNELI0wfSDzv3VDIAUkhBdoBTcPw
KHLHAnxPyfL5IgGcmBygRKBQAj8qAQuhbfKHh645sGc9UVRh5IZZaJBCiVdiKroW
oADC4T4zpfz6bl0Kz5QiPIBWAyjCYasdVMD8LJe6wRFVa9b/8yW4b2GWphihLbg7
4cZBiFtwopuCNwtFnVXXrfnLpAsYvN0v9Qs+gmSf10qY/mjnYOL4y7onjrG0U69y
keFc5y3sxkgBVd/BPrDTMS8UqfFoNnVnHprBQ16yGS7LFa0uqf8A+caeIJGSFwxR
xs4t70u74QJRuMMcG0SqvPEDPsQhtsrDqBTMGW1E9+tPCsYnpFR/M2K3EZk03s5m
ofFgnB90v7bD2OHIiGe/oiM3yPdPGYoSYmA/jkSXvrOeigxvOWHENoQHSiSXheQ7
Hubg1gxYOga10dOE1ZFKJ0ZEx849eGW9mLX2Cn1C0kp+ZppTwcOy8bWa+vdzKpu8
oaAOFBEysvOHpllXcgDHpGIm6IeiMsduCsSeReb47Jq6dhLZ5xWWZn3FI7TF3HOT
HKq+y9CHHOQTtP8okl05wM27VmLza40Hwwleeo4o4+dl0yNM4+Hx4p3xyKT4KD5J
JnARZ7xphsdyifpYUopNjZ07azmnLafZ23jhX3e+49K9unfbTb8CcqHZxcFlGx3C
PagSYq8/IURnUH53lAKcsgZ6G4oX3Ws/ISdwQuRXKXesbWHlrLJwJNp9RBYOzHsT
6qo3AVrXVHm45fwLi5m6ODJfpFzof8d7mB8zNi6h7yYuN1jg9u8AlwYhTK00JjIn
84HZj1kV7KvPM8TXf+dSCLXRouF8CUkwRm9votaNg1+/4jhFnmIft9cWUgA4TN5q
1iz/fSAnduyccYjjKdtTs9ibttGsIpz22aUUqt3xXOdWu6aQARoa/gv0A1F5/0Ck
gfcl1bpR6L/WXMwNVN4TUwu1mhzvX5WpmKqMz2MlETuUXhgfrMLZRwPiRE8yqXHb
Y+OGMleVU2bYUpDW7aO28l3R414xi3oW7Dt96UMOebGBVFj9GXZoOdm/r05x2uKB
PfAUDUUcTcMsFxXUerRRFtvnRX+v6Va/RuOVS02S1K/VBYPZKS/XOQ7lIW4ki+qL
eAHpqta2fzwy8lBMM2P9i6atEkcm6dklIiWghWKVQv8yC0s8a3S+OaFFmO5Emn34
KiHhS6LJDSO7dkSekaRJPyS5/dVf1avCo3cPst1g78DjGwqY63NHHpvYD4e0NPl8
TfbkVRFxFNxTfVr0cb/UM4FehnpeNTQPNKSIYI5Tog1iz/O0/ogPvo7B/9eTAbit
Sv0oIpc+j69TOWKkuy1jK7XwR9BLJvlD8vYpjTX6a4lnrHimmL0NxYQst7QcIjeH
JgQuawUA6srj7F0UzqWxluvRAImruYfYwVaSJU6dH1fkFjMHtrM1Rw8dCxekQMiE
NrMj7qdFAA6w5WgeTb8jLRdwM7xE8T10jqufRldhwe7PJrt9N4skfWBKT2yrBTPR
P4B+hl4pkUVU3GqWPjxsPI6ftDlyCywmyYdMRuN6VaRuZuNAg5h14nyKQ0WefGf5
Yw8UGphIwGTn1CTwRw7jmadzYZ36MxxxVT1HOTWGMG2IL8MacjjOrR4CmOJDk448
qhSwKdasPByZO40UspEB2Ua4le07fsnhAPrNcWIvDgCq3Vivh0JByQd7t11NV0DJ
kmbzMIMolmRDVN3Bpy4t01PVlvgtwLs22AwyjfZ7Lp+hi0vAlBmqtqpHL3RB29TW
oM9GeKQZ3sDnN0PvCALX6wNlLas9LcKwvkH29X9pMsi0uh+UZ8lsNp4veVt+ktSI
CxaWVaTMvW590BEor8bo3FEBR3DQGCoeMF4zpuHAlsMykq2xIkLyLIXLwfYvw3Mo
48Mhe9Liwd7/JkqxdquWPD6jWIijmLmlXO3JOmHjppvPH0Gs9DiXQEcqugv7bxKX
QlcvQPtBXondAGOO+mCyR9tC7lOZFdIR7QWvSqaekJf/d9nWFt7+bjpfyJP8sTI9
ExpvLpTOHEc4GcBSGbOUE9XhSblxIwSEsbKI1FoWJ9OIG444/4ilXJKVoKsTUH/m
xlv9F22DpR7K/QGzJIEz441Za1AaRwbDOqmex+ad/2TnG7npj4PaQxdTkUXpTKOG
a2rkOzy1lgFbjCvzDFRx3UMKf8nJVMJKNCLe1U/xpzYBTjGdtvUZdp4tAISLrdt8
4IqURlWnJ9pN/XhMPjdHQw/fD28N1xZIJn0Yn7QUSgk+a5Ylc3DwmDQAIHl9bsLA
d8eJQ/GQVD/Uv9ZnytB1mTMKQV+J9WdLHxl+Xa0lHjnX9flHgvkpIRjbvCbcRtW/
B8CYRnuLpFnmrQkSgmy8r8rr/H7Er3ykYsA20/15KQ5MKhacq53V89yoidA7SGvq
VlJuKNK7TOb1/6SqLikoIltygiBxEzWUKJ47Mx7ZBd5KzQq21ichnvEx4XSdv+xL
8FgXbHJ5oCPpgrbtzz2x0JmFlaxJ/W42cvGwagDL0zlVEU5pNVZCxTIoDi+G7Jby
m3nngQbqyTmytqxtMqV2FWrMMH/rjAxxXpxjrJwnT9Xg8xNeek5ZIEsY6P/VEJwY
nq7jb8BwvdGjAu5/JwpbVhJyO/a3rsj489oAXlOGoI6FbEWm/ZGWBNJ0Hf8kU8vX
yhy6ogecToqHxp99LfJHDWyj+T1Ols8/VlVUzaoFLTjd9GwMVaqPJYcPdgk3sW7M
D6bNbbbGGQuOPsIY10XSWMMP0LxYxM7COrJmrduYxCage9milSGVEc6lKOBR76M7
wjqAozahdjc2MhLBDG7B6S6nbKYGWPXD6Z+lAFU64THq30IU7QJzonfxauTWdPe7
0zgtHZZ7h43E0bTKRRpxtYvtqFKidWabOjRuReqGmp94poHHwR2eB2WyHQHuZdJI
TWROg9b8BfnOiy/tkBIsjDcb79kJ4SUYoXDC/VL6O/pTAdHo2JGVdfhtZwisyPJi
DxTuGvsTHQYfjuxwM4EOsIFKieYJX7ZT8eTScQLfBN3fE+r446ywttVqgsXfkfi3
hP1SOuobs/KPTb47zgiBsxIN07NRDYiM3tpyDasYjfne9psp/NXX4hrIKXalOSfT
nHEJ1jf5u5/OlzHCzd03wyMqgyK5/cWaDQChYGmV5d99JP/YOcK6+67MWiusgmc1
LqMFmhmXkM6YsZXDLkhi6zYmcHxRU0UyGbtASq5E0XD+Wvk7pdJyuBsCI9zzOZBb
LmJXrSK2ZzmHI9JH8vk/bACE4ZLQpgCviTka8m7Xvw9vHEo2uzNHIS6s5DRJjfGV
+wDvQJSaeJJ+Z57u+/fawRSbt8IJGIYnDxw95c4u5ASbn1GBl6PIfgjV+G4V0VHZ
DdlzAcP2enTsc1Ik5V5c8JEZQYc4o010tk3sm0+F/R8tKqAAsYzI7EDu3JwCmpRT
W3yUjNAe9cSKTY/Oz9dw/TcUTeShy3YPnyw2Fe2q4FsTiHsBdmAVN7mNo3hSB0yQ
yuV5IEat314YIgYNB6DeGixuYzP/xYIX+2HSTZr8cleG83MVxz4k38hW3qARbBLE
iijV27Qb4XV8YuZoWRse+TBKroU3fdSkUxwa3Q0Z79UCBewHhFswiW3Z2YfsoTr9
I3+exNdwX7TFXCVf9q5cAXcP7q2oLMvQzsV8KQsD1VlXOO+isbLFK7HQ1XELJ0rx
5G5uzhj+rX+Dp3AFiRBpiUQ4zNJGF3kgnOSoe8CwqFssQSFf+ElkVUzhiv2ELltx
FTEsxN6BPDlhQc63T6tsHBP+ExUYgTzR/eYAmBYh329wGJTTUsMhW7iL6ytiF6lv
QyOETHgY28lPL0kNS3/9SjPIVgppAQfUkMVH9taebVcoZEzmfA5P6ZUKsmrpsI8P
l62AUM7MyOBG7Xns0abp/hVvEO2VK1Xu464P8iin+kJruZe4pjN64fvM5EbmrI44
JkSUTeMcpvFnBGoyH+u+zUDJLURbSqBz644Qp4tDKJfgeYahLRnOlheudduhlIZy
BWYc6HQCjh3BU4cHGtnYGzT7nzE9eW9RRfrWt06QSUbUvuPqtgO5P5MPbOsfgk0m
ol9Lr5sZGq1ZI7sfuXymqJqvCddQglm25AP6Hc5R+R2SVsRgNoYTAgRrvtV7rkWJ
yLW3SxuVgiFvft0/zJ50uoG21QZc1awCAksjoB9Woc+q5zZwuDLQQ7+ZfYz7G/Pm
IPw8JLj+GfFM2mNtrpalIO0KqO/MXeTM7yFL6yUQhpjDRqF6/RJgDiPKFFGOUIAR
yjq5aSzXBxJxklTUWv8cDGGeAM6fsjp9r/gFJkaI8ZWOU1JVeuWvc+LpG8CiuvnN
ngIvHabs74LhQZOWedv+sBl4yWTQdAxAcrAsubCA2xlv9vDmASkju9mGFfKW9XfB
4gxTxHpiX64v51NE7kJ2GK0deDT49COFTZ/WqGEjPDpSOM3ojHtZq3xFCx3nBH2m
WrJBKU+ff2LKWvqzLZc2ovTP+rzlalrSnBw+15X/C1XzCloA9P/DzDBc1q6rXgwC
oe72gwlpfO40jrdojWPOzdLHIAKiOdHFwkWRdMW2H564ZfPdh0Sh73tSCzvS+wWX
tzWB83+big9kJiSc1kJpXMGqvM1724wUCMf4xmhkfSmIaVXawoI+MPPJSYg+9hLf
X5ckxXo3R8sjFhL//YH/VlN4Db06VlZeu+GqYf8MWgRDBkluQ+r5kFsm1t6J4QsP
XozMSriCb5an3f4gTSY5ByqSisfXVzERlKoGQKZZbbuXIH3r3mj2S5AMsZQ+sh0w
1QcfKaTC8mVWlqHTnwzhi4OOwyiT2rlVGSVWxOOW0FjVGhSyZNll3qQTo0Lg5Nqh
4f54WL3UuyiRI2zA0yUIl3sJMiuqZxuerh0Q/0NPsm03UQ3uFKIfb/HzOzHtrt7e
EYIPpth8hfUI1RLnU5NX7Qghdk3loRsqcd2pg32uB/YkZvUbE2yalH2TMmPc6zTj
LV9RTPtqlgXzLc/9vicSyhshEZKu1d9tTiLZBbZSAOy8o+Nl5V159hgy+1kFuiGm
8ZxlFeoNBqC4iO6KvTTp2B2LvxnMm95sguBziLPClA/OQf3UVRZMoSVZwFFpEulF
Lolg8Nnd9czxq91/lNtytl5pXOkmkm4vQrCrNnX2uA9eIeqGpxVv9nTEh/u8SqWa
BwZdIkh7BVI4briwxZxwcWce7o4G5r3sd3tDoR/vHTnvZjNT1vGcB1ScinfwC7R3
Cwg0Bosixhs7maHdMpCpvGMngQpKVNv08o8vAV6gYRQaQexGe9jpjoQ0AMZYIWAT
OJF+huo6bSjEqcGQn7A27CK3A54byH3nBJcYsXM+kH4uJo8q6NziTpbFwM61SjAQ
8wws49FKMsTYkEeFlk1UV8nGnENfOgvsKWdzR4shjDgKDy3AX3pmkC+4RxXsiGiQ
UTWXZpYhPR+4zGDh34g94+Z3SSq8CVlL8nR05Hwf/+44VdB6WOMi8/c4sSrBOauF
rc65fzEN4MiA360/KKvg4X02lYN2kkutATxciwFvkvpUQ061CuZhFgm10OKnTVA+
bif3Q+GDu8Crp76Ec82bL6i0yd6+2Dm6S6bl33q68RDCLihwnm8r8ZY/nMs9WdcD
f5xdT3P9qWN7xuhAHZZD67NWftkZhS6Mh1sj/qavSRvZqUv3+3ecDywPWHgE+mEg
PFf53hpeh7ErlvMzaZgtCtFjeOGcUvL8z3HmwsE3xvAcWEPiq5l8Wjqdle0t0RKA
HQj10dg899l6qVgW9eFpksxem+JsKg4EwF0lFV7BcfTvX5HZF8lmoLeqVdnp3Uks
P1nLNNIl4kI2AsFhfBOIv7fkZDdYAfpXAXNq5AG8TKFN54K3TUt8BckwHz843N36
2Nox5TVjp/Q9lED9JmyoMHklYvLMro4rXb00Ey6BtGIxKOzAgpU0CLZP51H9zWl/
7LN15pyYmZ/s7ORRZ0x9wDtfwRSmmPO/idlQ/8uuT0lOMyJmJisChcvIh/k5FDCO
672V1AUT2lsefDSw6G+InGhLlpgD3EutM6fZhTS4M5HEQ/zGemgmr00IevQbxV55
S5aMb1aDhg7C41eUXvzmYivwgwbR9QBufP+Fe9baptL25OT/QDy4Ah602JdzuWXs
N4+RdkMylbrBbx3ntl9IMi/GjEPK/hi7izgAttC33Ahd6QztnMn9zmblTArtItmF
tvYQseUcF6OGflpmElsce1stEBWwvwhOZ3hTPeFr/NeccLvwYzb8p4gHt8R20wKJ
/IUImtMP6ScHwQdoGpcUX4WU7+dlVy1RXBFDvCNg8LV3/uEfX5DraIe0RVCvcDgt
TZ+5VAsR7na3VEb+uhkpEOn128Q0lNOuVchiI+E9ZHoPKT9YE5ApFRgupQVm1RkJ
MsV0gtTwMT/4ze68kkrcunTZPpe9FuWX75V8rGl0POHvK0vhTferaLiTFYxw6zwp
VH7knXzkgnZfw5YXL1oYN+EqMEHjApUbyWfK+CIAmwlM/HAOfNWShHIyARK2yVqI
bkscs9yu21YESWx75t1h9gwOYPA0EcRCYj+6WRO939EJilOUJeaatavzZytKOzYY
Isq7ZCsKyj1ppwgC56SLSq8ptLv8/azP8Ye0qesZdwyPUJ08mdFe+fTFq4utEaeN
HPwqomyu+9OGlGURJkvf3NNqXnj55KPk2tIWp9MacUnqgz2R2AAqeGqNCP1IZOhN
vhfmbg8yjVcnqWnU3SwioCFkV6kwBOc8/+2fiqqsoaZjuey0t+mgkOSJIuNXUjXP
NLwJZl+xfbVyREXSxtz9BnIr9TkDRJc1ZAITpOzlLFBVbWVadmx2uIGf3L874ZHA
jNjTlJKjibSldHRvcfKoi8g/7vGzi+R3RvjySLkPwtZxaKjo3q8HH4IKSlPo63fb
oKjNoUVNwpEZpsaHdKjohOKFefYOP4IHJEDfgKk+IuJOrXB2OFgdoh8zXcoEnA5B
8cCDLZQqh4z1sug8eo+XpUcM5XqHQJ+d7PX3DcGPzPPt2moLjWzAeFRUfRyFqyCN
bhmEUMFbcwJ6rCo0YvOqU13zfO2FSEog2dZggya9HsdjIsSOPoK1HadYiCHDrhBj
5IEZrucLmQR69ybxTwqsYRDUONjxZ6flYBhS9F6tGTiqqKftIHdSlXZcOaxo/8EI
kA7ReNcJUBdEmHzp9/qwhVnwm2yMUf8j51qXSeYmZ5cP+quaBxcAJIrLP0qGwD0N
3fR6V/lW871Hbv5lk++ET9MvV/gcDgc8V3c8nErV/iMDuMIqjJvdRBpSz5EUZ3bG
Bg7QCPYSNuC2UoBRNWtOHP3waatIvYn+dkXMxxWxCWnAg2lfAn8qv/9cMKIrWpXA
cbuAZhr7jTlUQYsiOdVrGsmn00eYmFv5mfq5KPpjRIcYoIjH8E1vmheIsQ5ynsxp
TNo8GAKrlBVizVR9/X7SmuXmZj2oTedsXbUhsS6Nls+7O2SWWOR76jA51ThMyI5+
rmd3e2AcocqQU9qRz5zDLLxX7Xp/mSMUGCJAV+2hlgfyO9K8USI+s/VJt0gChEuX
Wo033XnwWnsLWDnbkpUUKhkPuFW7pr5Sn3wwGOfJsFYPwKsH/3gcB92HpgzPdHQz
GKidw5wd8cB8Ray3cFBfKDJQFpAOR5lVA0Uee8zuiZutrjJoOU/Vv3A1rxfHO+iR
hNZBRUdVVz43j/j8WhVMCE8BbHB5WpTdGIHArwU+p7/pCAKEnFLrSZjYXoNI60By
sxGnF2RY+nzAtHmAVujoYA/x5ulYNqxQsdXZknrdjIMeNI52979PomKhXMgCtlP9
kMaKbvSfX/zttTAtdZDzef0s9qPmTvvqzv+xXes73IJcZUEtpLH+oq+KJBguKCYQ
jG54vyd3SLfh+d4LMve5zf41R6T3LsjfBziQUYRvjfiwXoj1WbVj5jPvveM+5d3H
2EBHxariucsAHGZBXQABoORogIIKqBJM75kBj6sMYnl7zYnuhDLojPdcs5x8T2Jm
35GpbyVCGoJZsaFKeyiZX0sgYVSm1J7Rem8sRQ/8VqLMxjFSuDHpsZMWhbiiERer
9Y5MGWH/71YwymPTNpsCjGbuIDJU864y4WW+AZ5xZkz6tQYzMHiDiJAihPPk325A
ZeBOeRLD7oPMUgXkxsp5X5tkzm+4uWYZzpg616LwKPW5Lj7WBD524B5c3thtZorp
n+VMN89RMljlIUrn0Ms3CDYTwgAeOYMs+BldtiUO7zLx6SQvOuH/KX1raAOW+f8k
7AkxtKIcuQapyHHzl+jE0yDqpCasaCkj2s4DqA3yQqRIVc/f4phH93bLhCfvlOH+
KAf9yzrQ8iXLcmE6bjryGybw+YgJ0kAsVVi68SdRfCnBd7tPSTbCbsY3fC6X35f9
bGJCJh02y/L3BqliJmuoey79feKfmwEH+GG9KyA8EIcG5tsvhHDKbuxDUN3q1l2l
NvZQXHa5DcrVXNO6fkthj4pvDePS6Fr1+87IDv+x7VNc4p84Vwadodfkb1m8ku8I
fFxr0NBzsgQ5GVSg1YYqqGR8FlQqW174Z01stqCedadZA5hSiH8qHitM+mTT6CAK
3dCdSOe5aFRXwor1Gt7tKmS62H2MksIsXnsUFYIrTwlxDp8lYzfSh3proRvxrbsl
xrxAZUkN7j5HoCxDoov79EOd2pCwclSOUT2ILZ2oy3SsOwcGqElNEhKMvDQXqtlB
YZGuu5Q1Rqy8EnP2ZU9JRa7vM+ZWGZJKISDKeS1j8TosLVNDO9xOS6clsZ9cp8ZC
a7zOY8idhw4Mdr5dUP3pMcBycsGY+bq1Ql77sZGT1nB6OVFEp03HdQ71gjxtXPHu
Da5BUp5eqS8unZbwAxmK+PHr5u8wHJJrvD2aOmceRONknx63zXUGEhNNWobqPHwb
zB4Stf4zLCE8ND/532LJ5m239LANMfrQYOsWTWM6/MyrSxeV6ipz424GKVTJSYK1
3ZBeAwg8ntPs4I0J6RzHw5FKJPNeFOmNSOSzUeWNw6aEQn4HhVHfJNNE2CwAUPSR
SrtsGsWsQSJZApA/NHgmp8z643YCFUQX/7i26ktM+nEmfAMSoanIDwe/o/j80m22
qro816tNnoKB9UlA+VtbjLtwkoNyTbaJVk/gByqL6WSqSeft9N19UjensqsSBbnX
x5BXLtzcKuLDVYKMmJoi19K6AKPDy70UkitZeYHi2YDPTRi2T5wVXnx2Co1ZMfxf
ovUDMiN5g3Bsjuk8Q+cpWiB/Z5Us9NMShaK2Q2Az+bE2tJQGhmExTxcNLYbok3lg
XZvyclrTSnotERz/rJIeFkJXX+wwFpLN+Bp6iZKcDzA9+Q7OVWv4cpzOvcYtsrRD
P02kd8rOtNUN3DeOmpxT1JBP0jPVuoztLa0REQviIaKnKBcFMnFufnx36bITQfc/
cQJwunuW/+Mp5WTzrEnHaTEL0Dx0QdIFrwUyayU8D4tAhlhfhIRR59mABBHk16hq
83zbovXm/hEOf/gZtPKrGNOSahM41aCxac6K9nNtk/t/zwLs5mGqry8Xy1QNHVdA
aeN4P2rKZ04p4yY6NBej1y3bYDfAgfeGiIEJQfChdt8Mu0dkUA6+CcI62+czLXDG
i39i9DfoUwsRHP2sUuZZvfpoNtVwttxEfeg5uZN04JtIZqPBL+NJaMc8yad/6kOs
NUGQrPo6wdtQktNRfv1FLZemxIpog8ckX3m/+YuYI3Dxn6mKCIqqtLYB5lHib64T
L0HCRmuc6sljUW1Wn3aa1MOovuUTfWwtySwEulAO8vuJg5vinJV4/+IVtOgN3S7S
gwVBrTFM0ejG+F4j7huZatnud1Wif0tMcRX8odm4EjKDD66ApLxoC2xL62OUMGtg
Ls0Cvs8ExRqcyCXePZy/xfqZDlWdERD2Xs4YlHa+GEQbmB1NTisJ2gzGzj/wRwr6
0uYm70XF5FcyWmWKqstQik7HXki5SoPV6cvd2UWYdWZuMMhlDv7DTml4piJuTVbP
DsvLe/B3oVVkLUISRjSi7cfse3BDz+rOv01OjOm/ufSdXVGoJtMaFQakHfNCj3v6
S1CmyW+MSwd0LWJsdQBC3pNxdFiSOXV3hpQqoqF9snT5NcNPGQ+tkOCEXAZYyKrR
4sPyk56apYOytf4vBU9b4ZN/bDOa4BoKjtZqonAcR/nwzmo1gbPwT6MQk49L4/ip
Csf/cHfWm6SsUckwiNuVbSQiP7xdt5r39lfhOYl4XrvF+GPnAjoJxcMpBPY403AZ
4WZZra77l7OZltvzTdsoJAgNA/IlGH7QUMBfomAFUYmapOt9azw4mupyvcLrJN0h
cuETooSzZF8pvyzNcPnWDC/Tk95BUsv7mSSHLZaafirVzqfWeeiJSW7F/vI/0v/y
8dtmOX4eCrFxRxbyvtsI1eov5SB1vyxYzu9WEBrniK+DbrAjBMC1sk3MdCH0RIyl
/JuVJHY73pqkY3h3xNuqvnnc2FaCgrgvnktadqvrKzONBjTqb5Yst4LEKDla8fID
5+BjKE15Gl0DtQfmIIINsyj/TyVC6kb+Co/58urY7p6KaItbhVML03FU+AEH4Fvu
D7e19DFxnCXwfB3Ro93FdGu9Uy4uiZLph7VX+ltUJfMik5dhbjca8lfcPIrp1oJv
0UAJlvAWEJbqcgs2fJBLaLIURRwlGbUmChaRY6agUpVDZxZwTVJX94WTw2iqVj3Y
BdvtIGITej5vOpTm07T+aUnJTs4PNciRBuW3MbPaMzJMvzjF4/gGSrbFO6gXj2XX
6561fpB926/I8hTPWMGRUk2aHYJMWBW50UF7wwXff510oo6efpHvJftTJqtDLndF
8vAY1naO5lZtCgn6FHgV5rBmrLzdc65Ymcu5WqrZVZyD9wwVpbUgyPJfleDGBoLs
X8Ge6HbthEL8j5sueBzPEBFGNiW9km+oQnc65eD7womGp+UcI42eQMgDr3cJA1dd
CWGPC4opiqTB1HwkfY6dutSvf/AFeevUSbwJ13H9WWSrhCTWV6TiqTCau7JsLQza
RVt2k1BEFzv18iRcWI5RZVzzw7XClDL6MEwkrD/GMrrCjrMYWz6ROFIEgM9X8hh4
J5LSsWkKjvFx8hyL8mt4CUzMRq3PGp67DzlNfkFTVvHM03a6f91BchlyH3HA+q5n
kp6biJCdXbW/okAHQND0ZVa5BJn2mvBiXTzc1EF7BQQwiyfQA9lnxEywh1ghMeGK
DT2eCGTmR3HJtSrOsieODhYqicDazxTxvEP6yCz8O5Fw6oWiFAK6xD/ICIkFNseb
FRL0LxuFpvCGaQcE3DKS1oaJdwJvoFPErun2pvkUq9rIirfhuMJZpB9cLvrpp0Nz
5O9ZONvqwVJO9zm6FahTXtmzrOuPSEP3hKTVxgnaVTA4GJ9yFS8lPoDgj6ZjeAyX
Oe26HVxaRhKTsnnOipDgpk9etaFIxTky5avDpYJJEJSNboPUw7aTPURbgLHgVbnu
THdp82UjKXT0uSBFCWhQ4Ku/wJ3w6zlvZxdGltojNJsbLqRkzR1VqZHLoaRcdCXs
2OL2o0rVbGWhTDL8l3luIDJOgERvXkkdyEPL83ZPrRL612F0QDPiIn8XyhWkBIoV
48l+OGkbwsVN5Swmhei7CHwunzmy3PCAaO6hrMT05qS/WQYXfX4CskDL8cPXAYFN
4qu7I+mvKTovNqBTXM8F25fHf+/AkPAeDmFjaMK1uHALcsDQI7HNsOxu0J/VUUvI
BPdqdjBdlOJcIHKRs0BfMae/NPWTVrVQmi85HkikJiBIhgFo+RAt9PZFutXED+KF
SljPNub+gpni1RBfEaFTZ7riCR6jVvGNLtQhpC+rFrEx6DF5XYyy/LrLlSjgSIiZ
0nQsokdc4rSWnKjSx4WaU2Zp3howNkdaLEY4rPJMQetIB+CDkVUlUB5ARQYmVx5z
M+gdsjSUDeufcCyx6e1s428FYKj+h9sQZrUiBKJLhwidfFdzHS/aY7ooAEU3qvFw
nm4vI5G9NR6UEJ6W1ofTFd/1nnkSVunMDJDDzjjh/oOOnk9bSeOgD5ExW1zTYZbz
ATiqw41ckQmxFkkrA8zXhmGQH0SE36yec8TwhvictNPERH+JkGd7D0i8/h7tESdC
pKmXQ6Sfwj7bpqGjd5akTExitqnT1bGVZsRKeqtlLjxwXsCx6wmGRCIIrlawsI3h
p83qpmkAyCv4UevkJXgXJsyUkgCuqF43CTqx0qAxhkuIJ4g9y4BiKNImeCpgaR+B
mTVg5MG/AEPA/b3zJ8wToaJ3sB68dhasFoYVKglsCtWzp6cSTSpCAbqbOUGF6q/q
3FkH6ZJoa0bJIhzYW7fXe7yEo4M0lYpCHQdhvADHxdap+S7xxgSyGB2gTswv3jvH
SXrsJGhlv19drDUXi7q+EmQnPMMUwdqSt0sUZKM+DVgW3jJBDxDj3wLoDYe0AdtA
g9bbd+1RxyMNT8IjLD+GIny/yF//EhugPqeSx7baaIqwy/1f+O5zzZ5TmFyl/QqO
PS311k+mM8pCGHQMLeefLSgHlzbakxT6QV0QqcVdAnZ5tcdIZ7Ngwa9UiP1eXOfv
YmJWOt3LMN/YvXXhrlCm8zwXPrnoNR729APiKxMN8XmMt5PJgtx2nO4QKbsdinqP
r9nraqsVx8mGLA8/xQjJz1+ZrjGxy4Yr79iB7T6lZoi6JhxWO688tGYdXAn31aMT
sjEnHH7LSUsPFjQ0JhoyhdcIqCYvdp8vgjm2zLrM15At3I4UHhOHAo76YBqkRDbj
LpzHOspqGqoMb0MYH5s5pQ4oRqXatldpo9KgJhXaYz+WOnAC7lctlom1RdRpCclh
qTjqwUCrbVgcZfMcsnyHxVH8p13/1pTbIRAp0PU8WIh7viCbDH3XjZKwOJla8ybS
7WdGtJ2isp/HKAotkj9d8e8RrP7u6l9phpRlYK00FcaKL+5CIzdgCs3Cd6mHF95q
Sb7cC3z4uByaez8nrICTkFLwygdRrFlo0fMSWwBeDuH9iZfsAnoWHj/9iGZEkRYz
aArylrnhnnp5CLUV/d1BtMIj8NnDjQF+snEyOTy7NcgciYKj/xpxbffg/0i0V1bu
NgyHty9aniTuLl0GRYgUGf0vNnhMYH6MShZ65lbchso+uDeMFYs8TPFqiJAUhaT0
X/iaobOTulH4sMqyHr0AtvoOVh9V8ibPU0o6nbQnSaVIqlvlcHM9qIpRUD5Y1brs
kVIU5FpzwlDK56ILzl9E2XuUv8bupWzQnL5DiFNCdMs0ahfDAROEMiIvzBQ3sAQo
aRBkhR6+fCjoBEkdPq4q1xylB7/vd0UlCZZPJhr6i/FPlxnpYUY3DqJzCNtHRsTj
7xHFov+D9Bg9zJ2aXTIPLvcp4+wbXVIdVE8r7v3m9SeAss8eHq3Qdy40yMoUz6oM
yjbwc5FikUHbHE2UwzgThGP+nFLQWVwcfpgJxkuT3hjuYbG1sTd6QUsSx8d9sStP
Jp0bdFWkG5oWZKx3sJCG5UA3SRTnUsBRWbZ3amq6TnOcQ4p7WNtRgo28M8Pn2n4D
Lz+4wVVygcDP2CUL4pEnVjIz5yffFT5jjoQhEB+dyo5e/4/QeZzs4eEFxt5TU8sB
XNTeq7492qzECVq6ZQ6grlpA3qFxdZuzYEN7d0outbarypysiCdxDZf4DfUKdHI7
+DR25hKrB7ESeeIyde0iJpLUybrh/aWsSAb5Jcnhcv9xWCTZ5HGYnJO5uCqzc1Wx
Xv5eXUljvQVSxekd3cWcNcz1f17NyWUzBkLWKi9pzVl/nhPNOGtpA2XsPx4tbtu8
vjlaXuN7qnj9UE7GZyo77TzfN3ozlFbyodhkTCT94CtPMlUTtgfgAtBWSesMLk1v
Qx4sWqZrKmGbK9caKBaa6NDwA5+O/lwCaOsZUINyjGvojawdavhJBeyCkCXEgj/r
6/WQy2urhWFgdDvBNXcGZhskbm5ZuDYVTjnFwHTprGmfMjm+DFDafvHCvlIa4bBB
HSL7LxVTHSiZjvaX5pXBbQUW0j9/oRP5hS/VTNxZf9jpqn+zyIfJmqkWzZomHpnn
sNnYsJHLFJkunZuwufj3RITyWJQZbDbqJZ5RuBSrfgELd2LUUZ6wh/VH0hUdN4J4
K7zQihe8R8+qmepbksOCf55+7YkC9GTMfaHImhmxUJaxDjD6iTgBUxUx2HR00zUX
U/WFhp10bAxv2eWaONp1owAeM6hLhCR/oTF0Ws90NW6VQ/0HW5yJTAth7uoL1ZwS
jtX/cqMCWo+Q4HknSSPAAF8sGp7zUPvBWiSReh0wF2LP/pUp+nPftFvw5vQhyiO7
M8Zn0fVJSiyNxcIfxmX5Dc4qgjgG0ZZDGpLKMMLUmJ62iHKOimJBoncreWkRpotm
6Z5HW0ji2ZxMWfOuNhQ67BSOwbT+gTASIJLxB8ppAtwW1QGx6JvqN41JzVV8AH1L
GwFhDADg2up+90eDXxbd7z5WB3C2tDWZ3b8+1tWkrMQKurMIE0dRRyvC9tjYn9qd
JvCEdCyfOhSLwEPblFO0EeRXlJxGEuXA6GTeF6/lEHSzVW8u+nKLvkRHVfio9vB5
3zpFN2R2qN3mK487zEzsiP1Fu3PXT28blOC0Uo+CzszXOn/V0e09qRTcT1OsiWdx
8s47+9gG7j9246u9GsrIRdEzRr3LeAudWEI7XicmJQt+R8x9v4GrfpG2Dla7Nxam
TD3NmA5V2lfDluOTVlo59yUgK/V/DEay9pod1zYtdSyoiLhxjenuScYlWWnrDZT2
06MQJOzwLP3m15B8dSN6UixGj3osBrEyqy+Xtvf7lmtTSX7FOo0iKNmVgWQV92P/
ggLzBF/Fl9/f/ERXLYoLMDknl93zdmtoDlqU/JscXQDcNcI94jRCe7uq9eHBfAQH
bKP1dlVlU3tfvCXx+AQ9ZhrBNXQ+yeQDmw/ccjg0r+IZUqIxcZm/fiomAomBbI7I
mVhqbhFZY/iqcvIRlgSWm+lkFS/nfzuSC5+WuP2LH8ULHAukjkXKP0kmtQh5Iiib
Cb/KbJJpmtTqVcTPLTC3YFud/R+f24CzP5YQjLz546LQTDzSgJSJICNccRfaBaWe
sK26eWCrbhgCPk6LpdLnmh6wkv4DhvECQHNjsCsM9tEARKoM9Zn93EesQXOmEB1I
t2jTsiRQM6mWvUAhlwjKmeRTzJRPIDCSJoM3aho+JzqP86H+IHlv78ZE27E1ryI+
VkjxsjTMbKkt+VzkF3zQG9KdW+qh5jKWqoTcgqTl+WQIezbSK3QleGeODKMjhii4
y4/7eAdmfcZqfQCptP2i+qG2Mm37dEuKMZP48BM6IKrjhVhKNQ5qrx0TNiZ45rve
odyxmOC7wHrKA+uagMSAyhRq4TKEZRENYLY6daqAU/XQEFzMVgF7uBDnWBrVcudS
ccB2O/N1ff/465gzCIU0O2LQ9Rvy6rgMhHBMBhs0Q8SIdQ9anVDn0Yvl5chcGgQZ
k0Jrz6qExzWeoD/ve792bL6eYe1c0bT5AhZnEjnedvm6ZCsXLSLxauTjpIXRmW4y
eidfCjDYM3WY2jxH1qmM0vOEFfW8+3ev4xXED2VSdztSRiA1Z3OUZbw6CCjFLCbH
vPnMBdpfEb9N27vahia2BfJUZW3+rq8cJ+fHQPrtlph2p6SM4PzGMg/xjdpW0udJ
HQBpFxHjcmWEmziAo1K+W5JZcNa9fBRlnJEYGnNu9ptMSsvV01RfntGQQ1XASfY7
I4lCsih5eqa13p/JbTFKk9KicbjRSIdA1NCOBebjECHA5DvTxS1ZRJj5ktW8L/xE
TVuc6imraQfa5I27rFWWcnzRvFDg8EsXH5Hs9adNdzoEl/IR4dF68x+ifDpZ+Klt
uDwOMVGitbKBKQ3tRi+GBHZXvSAk+4ONxuV8cYejnYp2NfnnZK1twPqXbmjZn08R
6HTdqcqgnQUjGuHbZKwGjPXnb0QxOosqJuQwMQlIe7xPqay2TcwsaTZM5STh8B+a
aSdSlYtVBOXi83EiR4f5OivgvMn3V++nBM+UIPd+yOLdy6MXfV/YVwDkKJUEn7dc
1z0imNd0BTuNCGLu3vVgJRrYvAbfrwRRUg89NftYn0Aq6JeV4gMehqBp0JqgrpDs
fAto3+hqsPp6PS4SfX2YpVckkYOlzjPaxbXF8C6IrD6fsL13w8lprNFsf41XGKbi
Cmr21Kmsnv94AY+bLlnGbKEaZAH44BOIsEfah1V1gakrPFBh6ByXMMrB71BCK/M3
uIWGOEmFcU5KZl0qpkzAwhmFgxsaPEu2uYd5jnOObn89Vfk0v89FefpGMFv/W+aX
C/N2En0lKYH7mqvmbW9hYiVhhcJOUByOKEDvFkXoLQww7cFsFTcCX+Mw3lSAhBu1
iOtC7yqZIzrmIAFuWb70mRjTooXNybNURoaBeJWhc1u66MJFETzTilQphUqmeLh2
Id4WqysOksDKlwN21E+oLH17mh4fyOIV7yAApM+U9UOCDTDwRbT6rpFqY/cGLaEf
WVKiHZqXyfEennZssLLcTf87AX11fg805O2abiiMzWg737cR4CDyAQ39uuo/5sjO
3x4kY1Iowj3WnRmABdp2QHmoi6V8sfWdSeMxLxB33AoynXcjl4NEViuCmofb1A//
nYatVrk5xGxZ/oLJV7w9qgP2pnN76mrTrgSHuh3O3RT3ZUHUJNvj+o3Z0XAj6Pg9
UOH0MPwhuQaEOBuSSPu0oL83/uBy9Lt7LG2ss6R/QkAMxPdjZkn1i77tAjxoFBXT
nwrFnhOBNZZXFJzOXS3ZOt+cLzwmzSAN89d8cugd5mcZu2yDkz2HAHAoDDrYjscj
8YV1O9q5YF4MmiogIv815KN/3lFCwJ87dL4LVZcqH3PeMvYhH+WvZ0gMDEi3cZea
Yormi/axMyVInDPo8nRV4KL8PY1uJeGqpX1N1NHutsFjt7ng4Gfqn03Xa79o0UdC
2pi3Qo8lNzujpVjtHnyDH0KPIYsHURDhdcOyxbtsyqYctnPm8ZuACnCrXNDJdiDb
oOrKyj4PioBjzmc/15JMkSeXfM9E/HV9E8ZQhujIMpYSlV8Dud/7e9QA9yutClac
egpPxSoN8acLZONXFUQ7F2kD/MwBvUlLp0qDryb0OBRkSUIn/G/4rSlXUInWouVV
5SedpwXbaVmG/ciGp15Pfp+Q2tOB4FzE5WlUoVAOVgJ5als4QZCrTAoCWl3bXlxK
oTM6ynygc9RmUpBb6o1A/kSRF0Vyk0l559jeZT3aYJGyLQmnUcqVgWqbYfgLkz3s
r6EbaovFqWqoirkkkL2PZ03D9RHR6bDzaGFkWGRouU/0lbF3zIN+zv5TuCGILyCW
4n5SQkAfoEq884n6qHNlKMeuxMlQAnqAIubPH9uvPZWjSSK8T2Hfi8uf6aSDTnR9
VB0Qsn5dWidhqYeKB4cPAKcDtvAEZ+rL8Z8nXvuL5dHjSCtHFgTmNTFeQh+CQq/e
d5TwkWpLapSH8z9mpfThKMS31sV+BdS5cPffjcDA+XBEmU0NEy4+tJq4b1gVoBRT
O+YR5QyYZ1Z2dVw9Yvk05itGUZ9CkAJBOgDfL5LxGK0mFPT3DehkOLXzulU14Gxt
umZTPKjDPzOvBSgVKUMPNKlHmhnklrkYz2eHOA33IaAhM106C4CDOEBDgElGCAn7
B8rOUJIyXem4vThD1UVGzfOJurWyqheF3cPhx2L532zs2JrdTyf32p/xSgro/DG8
DFsZL+QezM+87guGj44jqeP3dEklyWkkQZNxo+0JKaajkeF+s5gzKNFCXowTNa6Z
p7qm0mFiab3DdwcTnQKyaCRLNymgBfX8lT0vOEJkqfiZxM/Gm6q8XpOwdb27K1/2
/mLWOy4snRJ1LkN/uolBYLcoqPe/n8mLBLTKeCZrH5P7/vLhgTQchS1bbkft95HE
yeaMjRjEhK4JYQy2cta9gSzxVbAuLJTdDoH3Kn71QkfZK8TFiMq+iOzKyghwPasC
/f9T4ycJu+YtSALYAwFlOllTvCvjexLEDdUIRha12TKvYxUnROrESSoNkTIy3uH6
JK/Nked8ShuPVaL7KGz2Kp/+xzkUl7X0EA9r+yNgOIfmxdsgyIwkDGIiwAxjT1mD
SsaW3UKiJ46fr5i0ShL5T7VTRlNn155AlPZ4pBJgkqFDg9i81dl3c73ob3q71ndN
dPU7urSVx2175fsc9U9irIk+kk0EugoTgTCa2ceZQyAXpFbtN0ilWD50VWTubufY
Cq77W7IJuoy60sjLEIhfOh1A7sYr+m+zfFdFLCieU5h8OsJnEgBv9GqecYsFmegV
ufZQeaij/7xUWNHBCa9hHKNEVZUyDElfiwptZF87n4twXiZ9Pjk5FE0qYAgf0Djw
bjQQ2sIl6rx/qgRa8IRQ/XFbPFd9DJCWXnJ9pbP5AKoSKGRvcHS+Js4avr7P4uaT
IwunlKr8SySGXHVM4tDJY2NtqxGrjGc+A8LLBZpShQGidOlMhOAzZ/XPCyuJXkRu
tfrBwiNtSKaR5FQk5r4hzZRFqKXjD6n5FSVYjHVcwdO+teE5skKce5Cy8Rd36tgk
5rhnyV3/n8faRRNsleC4+yC+DNswT6jY1hc2yAw1gzJWHAsVLv7na3sRWUJNFvAJ
itZnnCYNvR7d8N9VlmB+7AoVjtSiv5arSZXnuJqAblE0N5EmTYyax0Oi1/oeozwq
I231fV+j+C3qyMYPnq2tlfrYmsnkRPHZZ9bqt1XXdZswb/mBR85ZgUovYSmDHv34
QuxK0cytS3zd+vSAX3pbWZyaeLkNtL/AcARGigQ1ANK1JUh1wR4M4CwKkA0P0w88
GfoaDFbV+jUmwEVT3dJccX6VGy1tHM9SC7btsXDAiFI4y9/mvmAoXXarno0QkmcO
6VIvW3hIPGKz88oiTGNBAF8WP3WX3EJXNincV5LI8XzE3bX5aCi3CvCU+4moGMlK
9dj4WasRnPBmGw0fg8hl48pbovBC4sejERO5jIt8dw3fl/FH0OjzAY0PtEEN0ApR
Tu/NmTZRWX3OQnzKHg4VVmHv1PefF7SLSk5AboeNlBuloO95mF1Iev4NRyNPQin/
TXNlE7djl+peg56mOJox04RBRDDXGVdpxmnp+xMfjRtOuc+wIozzsTWJtMgJSGjn
dZKM1zwCYSTFh62rImKBs0kDtC57z3hMcYJWr4C/IIoYcl4l+9zETlU4bMTJ3yhm
CIe251b8STpfjC/3s1R0ZO/pZF2UQCn5egPvevkAGiePDx7Clx0OxOj9wTsygV62
cLRp2TqAJVxBZWMENVrUa01HtoNTfUB1b3iROTqSVda7+pN0BUSclWhiqPARSsVJ
yakcJ0RlgsO3+hoZ1qHObPJ4hgEQO2/NMvrk3rtDfrfkigD1DrlnPPpoIh10Eku9
lCcHBRI+6nrf0CNImKx4BOJkU08xgeGz+7bCB1PF9WQOdpIE//vW48Hp/QzWk0RG
796bzs10B1O7e+HCd4+9IhDlWRfl0r2sR/NqliQdQup4ixbsb7wI9TwMNPRsHGOR
q01VzDRdGMFdLoTkHH/SOw2nBWbcgzELLgnjeiUi8Aof7JatBZ6WlVV+pIqaO83k
CBZbBior6Nz1w1VNdPWAUeimAth5xjp+eMYutSNozVdSuhfz+qbKr87CN9wEO+FF
wAY3SDsVr8UDUWPufMWdfXKV5BDhrS0ZTpQWUUP35Kjr3z5CXqRonDB3j1248V9F
pIFRe29cWn8O6dSxQoZyv909Hotm93nfA4zA/WN2pz1zVy15PMUVmqPp9g2Z0W3X
T6uKnE+QIv1LnvXwawRLbE5gYdoKbQsE7E9bhXnvtKnuZRtmCU+xPBDv5K9u9m6G
uWE99YUPiTh9mr/keo8+3ZRND01LFvR5Sg72CLTIc5s2OoKTpxcB0aLm8UjQbSUs
MTATR9JKtgnxV0IQvE5UowXBFsqgZrgbuN4qDTBRwF2WyRKCmWrsVGZxLnmCZQ6Z
2/mn60gFbecFkwC9OykhBEk0d3BqWPbaCaq99ZroeoJgs3GYW0gEn90cQzrvYFui
MD380My+UMLfpvsbC/p9gAtg7UfnD0hTVokRdXNk7+/CGoTZeZKAq2R/mCeRTrFU
TT/1TInIA/0ib79CCnWBqJW2sEsDr/ea3rHGITN05LTAWATCySvEEV2pJgqTJc7N
z5dDdypKym44bZdKVZrr5N5psmIB4M6I+0hKPW36aB5JwldaIZRNA/22I4DUtXHs
RRTnF/eGaGceCYFFDgRnwjOFFqaQSxtszOjUzVyr9+dHmVeq3V9AiRb6gOd3Jg8Y
lggmBlFQFYAY36tAQcEvrsFjY5M3EfB+0OvxY0lBK3ChUM71H4IAKANjSpSTcHaZ
Li1XFZjeyjvXrq5e9BTs9NJSQq39vdKnArVZxfVoK071u5Z5dyJAzqJv0q/vjzDC
eO6ucTkTwOTuQEzWpXlxP6Cd6HiV2U6wOFx/35Fe4Ugta8WUQP/pGj61AiSuqwZW
5pT6dwWFgYYPA+QDGmun/dSX6zTZ24yLvccB5G7PzBOF6GtK4QsadjCn/a6bIy8b
M5MZPu4rPhcn/rQ3pRqtBonlyZh4gUV+2lPlTKSuJOf81ry5r5GaNDuKRJL686rG
pyme7sGbbltse0raKVG7nFveQwhwzpXxES6UUsWvCkiXSFwD6gVtxFF5zNwi0RsN
LNTJ1xG6xdY14oBOrIk4vIVqXaQ0028uTJWV1iu4TxbO1ifCpWoLOfHjn0THasEq
wjzOZCoN1qPEBMvegNLnds6l6PmLOoVVWCIqXToQ+gst6P736DEmgTLZWhghiWrP
KixeBvM5BVzrrN4z/oVTeFFUoKoezDdoBHkp3IsBPpLGbnK52PmieXJPPzGZJWBG
pqT8dMjIE3fg6k0R/eVF4Iy1Q9jOoIp4qVri4aUd2WC+yhRHK95vyVirvf30bj2m
RhOxmpXefgAZ3S99fMOZDAJeWVnW865KPHrVwdblmjtS/+17YSqln7l9ERl7cmX+
4Jv12K8GakAZeNttC8VXy4XqbjE/xPfZ+9g5kLvYsV5boS4iOAMfUhYLzRyZrM7X
DXOw2OpEzk/jB9aPY/GzkjN0jvlz7ULc9YLnzz3HQ0kkDWFKG1qSEAlXug8SyqhP
FzcWnckiZU3DAvhfwRDPMPvEn09b93clamsBXkT+R46vs137zEQSXiJ6PmvIKRtI
yk403vacyVrFZlIqChUoHCTsyuChXAUt5FL83zoAx8Zg2dDUAt2LKh8JrWh3TBAU
Y569UaMeO/Da8ELU5FmfQqbsb/6k4RqUPJXdlpjI0NzPC4jCQB0zI+OBYPP4dgpd
n/Jhz8kAmyFYPsHv0yJ75PGV8x88myW7G0Wn5K3KS9CW7dHqG045WExIT25BN7nP
+1LZS5EV6ZJf5s7HDTOqnSZYSU/U771Voo/ffCLTaSPlVJJlZzlEvFT4gl+jue4w
E+mhezY8JIILIJ38km5/M0gpHGFuLWmSH53JwDf5XLFDG2OWn6t+HsHw7NAgMtok
UKY/RRlFUIGsq8Y+vP8hc3AD4Y3DkpHYnvQcVvnM0w+ADPpAtdqj8H9A7higZm7L
UzSDtgVx81c88IMzFt8JNUbdcljHhE6d7/GTwScujVunf03UcIRDhPZXxGzTqGVC
sw/zjUceslMOjCjAFV7RLqzK1wPLtBmaejXw9fYyhaXyAk5B6sBaAC2UBisvPZ01
jY377oxc3FLJN9E5Sjm1lX/3r/M7OvQEGzZDsgIntuJqPHeTGH2v75y+lhbi/T8H
LCksHkzyrHXIlVVE5uRZ3Nt9X6epImjJzwySc0l+CkSCXJu4tqOhbxq5jTr5886g
PMeOP/fTbfczNz1woOSaFY6aKNN090g6WlJeI1Z6WwjY3EmwxeRusyvsFTEvNBAp
oFzX8vkl7rts3R0K2Lo71ltSrDjKthfsO8Tdg/7dYduCJpM3L6wdETyQxQjq3mOw
hokzq4BxogeqQM4p7/IVnl/aU+TyA0OOxvmldWm1RAlms1kmIu+vmrOMUaKXOKwT
Qfn6d9ypcvsFroMDj9nTot91A7xYsXYCNRGGOpfa4s89T1baNNw3GNHw3DkLmaWJ
QXyAnwpD8Zwju4eQfPcDtuTny0gtfwQx0cF/71xoGxoAvZBpsQgxwbRZzwdJ/Wci
CRjFbaJ/BrtT8tBdsKqIt81kguXWkO4QK9UckI0/3AQ9LYGI3w/86pY7l9Bw2Eax
ze/MPwkXGWBQVWfTQnuwiH8QVDqIY/yT4WdBcUNEO86peAGMUsKz8ZAIOPrDB45j
rwy6n8F/X6nsg6qyfaAELmXyFIwrbEJYPsETUlAlXGZmhY1jLsXjskEkJ9nIJmV6
GJpjGF2KGMebL+fzCiftiTXIgtgDdqwzgvcocM2Gc3Iow4PA3ix4Npuu9b2W8pEN
h+sx5TkK7STqLOIk9XMTufw7SCzlriKG6KKYE0icyZTjxouC9Cynk09chjchjNuQ
9qsYe17OtYn/VeGUdLIrALYUKUB6usZSu4Jogkn2VeMEh0+JngxszTePt8VBj5cz
nO5O7N6R9Usjs57JowHz1FEJ9Ih2GEH5p/by/8Hxwo3DAM6MlwLw3hAXGlAHZm2b
Dn32jRDAdr6f7Siqignar6BzTuyr5jHL1021hZBApHoECb7Q1jvuz7MqCQAvMW9g
FQHA3Z4MPhfpqwn/yoTfI2A+h+FRdzVNZH1NDTHRwB5s5ShoctY6HdQ1fuN/c8p4
0bhj8IwNJdn2pSJSZqMF1oD1cYX7gF9mKw6pKl0DFIXFeWcbDsKSJHb+EKlYbQvQ
i6nxtlWeSroOqXSit4XBseTq6umvRrp6PtqwRxqVBKgKZhWZ+wQCPGVoB4d8hfg/
kFHjxu4o37qsmzTe7vzFflsp3RQM3E7zcSxqMAVUwuzKc1zfDPT8Fxaexh9xB0VE
+WRvT+NQ00GFdXss5immUvOZ2BLR7AoIeAibQpSqXQvxbbCzpW4T3fIeRuexFptt
684vPz4fVQs0tUEtmGamO7BqEMpiPK8/eY45HXMhaVuvEiiABFwkPwe8ex77Km6U
U4RUA0EK5hY4ILhSqUI9urlTwFyv1tVqHX6cxoUAyL/Osvg95Bq9dLnptDusC7Wc
TuZ1CG9S8BEUAsRbZBcUDiBYZ3TUvzNDlIYY0FivKi/1ppNpfHEWfQ9kN4Rr6mz4
uWCoyky1bjzyOgpyt6P3mJpRR2Nm9xyMjf0wm1ZlTP+5/3/C2FxbyA2ZxrfqwOwo
JO/AuTXyvcxa8Hp0Ea6mwQ8f5NDivTXv73FkF0a6MW2A/QhWBjVwgVbJCTkzifv8
kfHz7BDjmlJajp6u/QAw9/4jsArsIJVhGYaSluy++tNgppnOxeWXX9xuS1CrzME5
bQSN7P9wN3nXTUEi4gxB7EFPxpr07s8hotqItvOJRVUcaItFWhvnlvbeYRc04deZ
jAr3vFsNB4sYN7hw5Bxic0osBAgxDfOHnJShwblFqtDna/JDqp7hAOmgmNq5YHBe
IMqiR6YPhRJuYsn2AId6j6edk0oW0EwqGgyUXYJjZ2sYz4jizH92D6tZNMnst3TT
34nGKXYfnYShowuXfK68vQkFqzAmBp0iY2bpIMWxoMWIw7wIbWUM4hHgayLkT5IY
oRJ4yLPkwMAR56LJYYMMCMoQeVNa9FQz/YXq7CVkL2RsuAB2I6QBVcYYDavEs7df
u87jPEN+HXVIZm+z2wVvQSHbEwlU03AMFrY6E8jQHYzJIyXgkqczNtDI2f/Hsoov
DsnqhaFNpW/NTV57/aOa47hZO8ieVApSC2Juj9GOTNs8UQOsUwSKUXL5MPWrjEq3
8PiN0A4vxb9iSGy0m8HX0NocULvW1b+P7XDfRvFCVJ7IVqggjY0gJVB8h8233e4N
sQEU+D1lhixq8CbdXFqE77Bg5Trh9Ll2hFqA0MfrcToDPUKnQDTwnnubGc25+1SL
wy1UOfzw+PB7aVc6+x7A+qDqGI2dnKirL4p3XZV0ibhoEaYNAnYu0JNUy9N5gXAx
4ff1wRMhh2D1zn0/W7xkKdLl+NZAuF6uVHdCw6VpTz0NEplJvf1jfs1gmm5fTCfq
kP5PQZhP2EOm2RMiQaHOVKRVyWldeGZjS62bCLYSvxqEKQNnG4W5iaHzWd1eyg8Q
vazAy5t+37TjjqeTijYpCwrNSz43/inilPALNzTfVcz8DUhxSBrZjIY8QEmdmeV2
CG5EL/D0H5hbB8PmNonhEz8tuDCzQFsR61uBsuA5cbsP6znhKpKWS5fCgUOwJPZ6
XPsL2GD3pBvs8XwRKY7fV3r3RkFaBoOqtnjliJsCaa1W/Quep/2D4PevhVmL1oeS
+VFvB5iK6dYa0GcspgF+xCApnNRB6KvBPkSW79Hy0gXrEUj5EdqvAkZg2QSGtt0E
6qOeF3vWAS0nqZ93ntlHE0Ga77wka2n70AWYM3eAI8qT219eqck3996UE/4mv4yY
p5ZX2gH4gV2pBPASbJ8pGDIlz0bWClLHE5HyRQnCFeFaMTx6h+xS8DeCr8y3AaD9
IN3jXMiIik6aS3hy+tL2m8QNyplTri8Q4ZJny3n2XSXIRzJJNZ8vlTX+fzhTepca
qAeuWV19Ky7N30ajHzzdHP/RXa4fifDkmiY/1MJzqbGSz2cDRhWBbOPkqtN/UngB
6uwK99cSvZ43Msm/R4hnmRkueP9/38H5oaSVcQ4sHaztJ3kcpRPIDR+jP6Y5P0mW
GeQbSH5MmpwUIvrFn60hNwxCiPWXO394JZmDTUQvBmrfDa5GgFbZbsAzGtOl/L8A
YfrL3kytZLgrVi73KYuUlEH1kHPOxna8HUT6gQlyKdO9IoihXRG3tPhsnyiM9/f9
+ivl77bmCWZ6lSoJMEL6C2tbU62paBLYVg2UAFwDSjKCMXswkvobpf9VTb+sL/o4
5rWHCIM8TX9FDeEOoQLK31aH3pNRhSInA/41O5bgLSL272RN5185j2jwT02REP1D
LFfMvQUyKpLbCiRW6U0EcbfQpxUa0VHAE1WpifkUw5Rz0gr4zEgtTqTgJxX1FZDH
RCTXZm4DI3Oyzkd86+5MZ0BjaVBUHlHU4GlskYG3QMO6BerdZRd13G5veQwUAcG4
vH/buzFWQbJ5sKqAzmlbVLn04Lpg8q0Df9QDhWfir1yCGu4jcp6EBR68ylz172MM
Ll4uLy1+ACOsYtvoffsdLF3PAuSoJ8d1q6FwF60LOnwlC0RwTByiZ68ifML/cj59
Sk3Q06D+9HK7y1jQygXdNlZ7RAXEZ/1hpj6AdBXyRfv0LF6yLqnhuoWXfW4OLkWK
dqc8LWVGonZzgKtFfuPSMy7oksD5LZWXce0hdgO9ItbNP1qcGXZffXlkIZRLLe1F
6H19J087hTaS6wpJLYY4bm8j/3eTkNFeAad58UPyUmIZKSWkfoPaux+GOl4JR7Iw
QHVB03+RcRBCx4/Bzltc8d2VwP7wPjbcr5cC3sqoMRUkL/wd9HNhJ2+S/Kn/orUf
V4/sOHSVff59hnwJn9XHuZA1/b4v2ELh7WFgBo4O7cuDSy1M8LZrp8wFFFbcMJ66
lVS7vmfMZt6/G57S7OJ3GWiL75FOQU0y04qBn8B6RscqCAxJtZAG6LOc9dzZHsek
pnPwuVLt2gnoXlw5rvAkmD5cvuJpO1LZMz/okRrrjNOAkPhKVm4AQK12rGigTwOZ
kpQw/DkxtP3gPS0pAWcPBxZdw3HTAzZsmTXj2xn1lDotNvtvMcZTByT6Q+m2asNh
fP//rsA8o6+KXNAcKTgdhXFzdwHNGa3aYNkMLdnRZpqK5e0mbLoHRMKAhSXBqqyW
MKARssgwutoC/jazmdxaX7+iStKiE+FmwQsp6qCqLOIP58OhWUOMQndlsWQEjiss
tFhHqjRD9RR7EUr7g1HZubTv15GrAMdhYkY9YMkkYZaJbWQeXFMbFcvFvKuammzt
1nMOsn9tWdWbMCj7gXAQKnO9O8b8D7iq+3AyDDvW/aYPQd7087dnNnVgG4LDDc4G
H7HWpsZIHQFTRnfyO+PpWstO1QtV6jXm7vPXxcuuqdMSjHHbyXEYijXbZxjpBr8v
eplTzIR5ygfm93qFWFbpUhFs2m3FIkCWY98Fhm/04XCuBUfOAlrGULY3TV3DtJcO
9Gu/oqpvjOSWmDahxaWUg11a0U1aSg4/IQg7k7dZUFGO/je/onf4xfElLY2v9KQy
EzrSvE4xeweDmkiKb2Y1l5DJOnQ+lWSWfRNvaLrmn5ViY+60M8BQVKIzIHIQhVQD
BAvBelVLziIZ3hH6exXQY+pVWCiCEa7++Sr4/sD6Wcqc3vpHqbDksweiONhjh3Ny
WmJPeTloPQRqB9rC3GIpitLfCowtfLPiz/wt6ldNXHIJBTUeFv7Q4RmaggixHfSu
jmbKuWffuahVHy1H7DCj87JnJzY7OK0VSkZHEcDxXMoict5iYSHJ34Q08bZVFt0I
2I2DdM8UVcBUuB2e8cdOmOIwzFLzpS10kNd3aaObgNcwkjgBiMm1jPWiKRKl3RPY
w3P5NfyNGIelSml5+3QYMeofyjq/XV4fFBTWJ3DYRC6GhHxbf/Lpec4Ai2RrTiTo
oji+hJsMfCnGV/7ztSt8vY2XxnKN9OR2nFfyQGia2V4gktvpD4fF/o9A+81abKs7
9OOjEzv83yigaRssrhgGi2vd6Rt64Vx07MKJYEOFQ+cr8hqwhUuGji4vjQ7ja4P5
k6N8wA/6/JAEyNqY546/6EO/x2NoPQdSlwsab4ECNCvwbatkqM2ZhmFkunqwFxY1
yctKYJpzSWxjQKk1EEaR8yt1GjCdcshzLfpV9znNvR/LiF1wXsodGKhInCnsNm3R
US4dCotOaxUQvQuQJZJ6qRkB/ZK8+F+4mf2UjGV3CluDmLx2KhIm8qGBbzNWTUwK
oi/YieWoN+c2xJtq3pdvzCjEePJtgu7YwV8ohoJ48UsMwv98/tRHADGr/Gwf3yIU
g6HSSnNSmHh+IQs3Wg8eHMg+n1/qYatITBlMg4JZHIJdTn5MdN+2lvOVzk6ieSpT
mNLPYdwHsBignJlGQTS7KQu63fGoyU/mIjiM+sEv6Gsw5EyiYUixlyiwOuHgehDX
Kf1UASTgzxpVVNXRSqhZ+Ls44G4BWM2iverHn/FiuNtvtY0P1ahbYVmUbdC+u6b7
zXjnmGa/DuiMDXlK5IDGUH+ODbiB4QnUZwcdm/od/0e70QNE+D6w6ZA3wZu4+jPM
XDDgUz7apn6p8ZTO+eBcHRW3Q9C/lk2BGlFCpQrmCN00r9HWDP3WJh6yzzpUvPxZ
7G8kpxxnIxsXPYk3OadAoTm3wv9ZsehenDqybGf45/F3HgnoHfJeRoxxGvtkSPZU
ET0JzYyNcxud87GDAYAZ8uGqdJTuQ/6cK8OynwXU3giRAl5A8QnK/zqSSB28gGZC
Ap9xTNvY9QkRSkqkjofWjkgfafrQc+/bs55cvZ8XictPpTdC7of+O7Lo5DdcOgu2
plMK4sdvShYzU55S+ikntfzwFwLwbpRg09Ote/ga+9CUJOLxP9uh1ZMxll6T8O+9
AYdMAI/qDDYgTNq51fZ+Cm8CVuQbs5Uz3tzgQOUwyJgBdG+QAikiC9sKfnDuSEAK
Nb9C8AQZ15rwBFA6LEDbWytxl/ISkS00K7a0Q0jImt+HXciMlmq16oja30D0t581
XRbaQZRwys+rz/tnVp71Y7vHsPzZHeUV5hirEhlGcHRQ6ajw+3UWVvn9RTfkZ4xc
Ga+OpntW2IK2sANCZ/sAssW74zBbDG1WyNN2GW0a1N4zjb7QG16uOAe4L1aEE0/z
LioHtaNu+d3RvmROr5h/3/1m0urpXvmbCrt0om/NI++No6Y33kqhMj6sdoCyygfi
Epk2CIkGAJUtCj2b35Vcm3HD4b5A2DP1XYYTHV3dsSquv+mWE5bKalsBs25UWoBR
oxS3y2YG9NgvWR0zbn9QHEPfaDPJDiyfzb01mqJyUHK9ewM4RasMMSYcjRuoOSti
nOzYmI0gUQdJr0ywCHy1Pm766c4J62cNuqKyIEIyw1dMn39cJ5MwoxVxAhT7S56T
/0zlDW0AgBJIFoWLQQwq8VAoDNyAcJ5IJNNN6ZjSAVOgSLyqkpc+pdBz8akpweMY
Ly+Eu6cObtqq7Owhf3+ik/jMq2KtS0U7YCeuj/KxWA53eyiQYqV0y4KyRhK6ij5E
5CSq0kUlxONeaSswswk8odbk7SGaaYeHkwj7CFhF/k+i1c+FVNEKFxGSsVXC7qW8
EAGpxS82oWsp0iGBFG2r1Wdxnh3LxFJlpwtIu9WXEf01RUonISRM93YlFv20DhWH
bXiTr8bjB9Fs4PeYETpBP4hF4c3oPPqgepwmwLcoh0fT+ejgDcHaOs9K4z+X0ug3
Z9bME0jqjRfmsATXaXaqW7huxSiseo2tLqLOQ4hay63Uo0DzdLqN+TvnFdY9c2gi
g4XHx+YSEb0m3D2ep/G4jWYp36/cR77SI1B6vUYEUrEtF5BvuvOGe0qso+ngNo8H
wsIj028KWWTXHSK6jfzEo8XcKSp2LpIDgOp7JLX3y+Q1hqc3x6Y5A5hqv9rDhKSY
t50wmTj4wDpFbCJceVtFOHz3saujuKXF3xCKl2COoxeyXsd7CcHqxRprxTD/00uD
Za+V604PzlRJhyV3g9d6V7bPfkZl0NFLLd8+54GtO2Xd53nHQ+jrxBrDoR7Q7gjG
7h8KfQ/k1DZkj78o0ChGn+GJXmeOkuXz31nL9hlJPZMaSxlFCZ/2IY7GhdtP7jfN
CfTO8zCpTlpLyaNAklPXU94tRhAQZ7AMVX06ob3RaWmRkPNQB6HIJXpxtVoNRB96
IwIgqQDitAxs9OTn6LBq1/ygFyGMY5SiSKVVrMFks6RPKt0Z1Xt6nGZ2D1DWc+RP
caMUbXBsDZMubvDDt5ZBwqyTHzYPSc8jO+JQ6o8x/Bdenl2GqVT1ADSkp+18V/6n
cfJc/qc23nJtFgB6lYr/1XOrYpTO+u4JI5Z6cN40B2YHw+AKFZgxdJZZp2sgA+wX
D3WUqUypQ4JqP/SM3LSW8dV3tBtWZ99WKRE55CLaL4EuGaD9xVrZXytHQuT5EYmt
n4EYEpaKRgA1P6tcQYUi0TEIGQTBaFaYURIPctaw1kNp+qQY49nhAQDR1k+cvKVp
OYnk7cO0MRPePCcRYQHNmPUOTnC/yXJ789kRdNwkSzC0arjaHkST2RebTCxlPMKl
9MRtkUWdqc5VxQT0A2A3CIs1R49LhH3DVcODeiameaM9MJlgGfuRXcCEU4daE5d1
sVFvaXJqKqOuMc+GVtqY66Q1lH7ClVfm5NtjsbgeL29k25H7CzbKZRRmDRW8g+zx
bjNHWFMn4BfqnSrZ+EOrHDUMI8HxJim276wN2PsSrbFDXXQ2w4aRQ78Tw3JYHmeg
sUbbKAWYsJZsewpQEQhmJah4GMiuQQjKAszQcC5T+a6vw9O7rf6z4E1EWihQQg7H
DZnhF8QItds7YUpLSAQLJYnXdmg1sYqUljqqeQJLH/Jx4GPMSq7GIaRJY+7S1kmf
QdOEfeJkuzr6NRyfHrH5DNGTC+C9j9tmTtpn0HmWoeD1dzGQB2fCBxIvWMUmBkC1
l8bn9lQTKXhAsSUsXVIwoPdncQT0zjN9sZX8DjXBxUns9Fzkvoc8xORrZSzeD8Tw
VyHV5yjroAyf+rg5ZZSlczWI2gc/0U7c1RJvukk+GM8nsKV7hJ9XmLUlZoYwPI6i
DkYi+kZrDrkSIrdMevcxVMPBVX9SAooEo7536tDEWwtrm8FpMfcFDo8w7i+pVFVL
HYdLvj/BxUWT4ScEhSIaRTDH5tGwrX4NfmJHerR/sksT6Sb3YpaeKGSuk7uXsy+b
/YGjZuA8L8jvr1AQ1ptkv9eMun3QBAxBeQWAApmFAG5tzx+YaGcDhHmbcBVTVIoE
0asiVj6DbLn8X7w6qLfvRyA1XC/llOzHJyBkVrzbiDqRU2WiHsBD0Z35DEIPTvpv
9oUC86V5aeeO44vZOB7TnjxHhU6iC8FCBj2F2e4HiMQB8f0p1yiivlAqEGgoI9hb
+EHY/3qbrgAanVINnm0x0fZmwUEd7TsIOO9c6UyM2yqoY7OChadQB/APMdaSzlNr
1roosR2fT5TH8xposMQriQOZeyAOS38zAfy/Vx89l5FfPTXrqumgibaLFlL30/A+
4+yyvklmA91QONcMcEjxJc3gK5Lmd59J/R3miKtZqHPKrbst6c9PA5OqfdpHivs/
xlFSKms0Tb6A9nMP10KxM+4vZP0eU0kIK8MF0q0mmwkMn1+g4DQQkPKlDz8L52vv
J7sOUmjRONpijC6smbOii2fKLJt2zPOr5HXnZMNkQEhLN/qcIxyGsxDHEaLwh/Bw
xNa4OeNBgOblx0YJnp27DyU0q7eQ2UBsZkuIv85BtFx5F3pxqEAbd+TponCANIpJ
c1fuZin+RVvNRYvU0d3zxsD0ugSojHhlQmnJ4ClqGb3e1LaIxGG0S82UtRHZACVB
qJM/pfYBkq963AIj4WTjt9+jarGbz+V/DjUR8q+t4nqlfEWz0crEnd+yJy/4d2Hv
A88NvLQVA4iPDJEJ7BiNV7HqZdJVsM8ewZoTwhBTAFcMgyiJwOxKHYic2RpAuP0+
mLc293Rk4A31d16i98fKQnhZHBn1psEmXZwWAbgKUrZjOpO4by3KdpXxD394UwF1
Dn8IeiECrDjkUwuVVNL3YQkS5jDUn0EmfpFf/CmQNeDytH6tkMe2OzbcgNOmPcIN
gXrfZHv18FLXLAh7tVTqTM7gSwm1HJ20zojkQURhzlp+c7rsmxW4oCEkbvysJG8m
gQIuuDfIUzIi7ltc67OKbiBUp8/5GQZK9R+l2g+7NOEai0wPlfesPAdk63zZCD91
21PGksjk985N4Ju6zzlkpUxFpzm2yyqPi0/raoUCPCyxUhpDaWcb6tCTeBK1KYnQ
CLPAn1Ofs0KQtKA4UCbcb49LpxTe+jn3tmUD8skU3qobqLjKW8pbOYQwv1I0cMSD
LDCNNGq3ojZuU7l97h3GX0PVquWca7+pBvqEnf3R6XzygUXK0HCf3jmTIfF6qn6h
vWBjuRSNdh5jUqu5oL8hmPEnGPpiG0JeMxwSUtP5n3I1R2Sv4DDeq7cM5mdAOoWC
dDMGcoL1Kt6X3SYmkiugQGYvIvldxOM/BxMksyM85bTPGl09W676CA03Wu8hoRsG
+bcayTQy35y+6iMA53x9uGQ+4u6f8Usu3OKnAtEhiA92IU7spdU7kfpn/GyjVUlO
fVgK4umUz4KeYX2J+6FmWGbNyo9EYqNRgjSSRmZOneb5rdmK1RxwtW+9BK7nXo0z
Qm2ieTWfx01/9ypuzMsl0GMfeSdQ+1yezploy+JiUX4Sv94p7SJ2Y3c3bSzaom9T
IZ+SCbM3mN3Bn34x9znANnWr5GE2Q+2tR/qSaeUUIyWEWpndLkiA0hxini2n5eqv
+QJmlB4kfvnyqqDf9PoAUWeLtGVXHC+5N5nZq5BjvvWtZA/Ht9Ef7PZM7fHz+C7/
tj3eQms298FIv/fV2PA5OooGlqSmK/wGkFmfBx/kMUcyeyuwH2lYIArAF+LW95I0
dUgYkLB6mYR7D1Kt2YNYRg71ev/kNYDBKUHyVnK+AcOnCoMcuYja6OfFoXM4Ose2
JVg59vkoLbFkAZ8w2RFkQ0VJ2ukQWpwuSbSiz9w2D+W4X/QoVjq1tyJ7DsxfSjY7
y9t7wx3nNQxKt2e9e3YV7NOItZR3zfVvzNCr84CwjGl61Z236kr1UcKyaCwRfun3
VJVLfmH+GbcAu5JHqeqMXD8JFVf+5jliR91wENX8p0c/jn+9VY2DXmb8A/CRkaHu
xvvYLjg0B/fNGTrzO3eod5uQMoAgQMFSOO/Wv0ebdHpFBQ4ZlBO0EQXzO6Z/dmOl
dDQhE9zHiWY7OQtbWWcw8CX+stY5cBRHzCeJcgoolLdXOP5asXW5HFGqiVNGkl9N
ScfonAChvjJBCKQgi5EuvEkCxiZ0eGBwT7NVWxkUzKSkShSFDxuRuAKHH5PBOkUK
uRavpX4oXGzhUl5spe9xasA5BKtT/9SeN/BOG52ZQKY4EDFtgoNj53Ri/xhtQlv3
dMrUIj764KkvRfHY3jqyfAZIRgv1cyLfbE//9tNZClY9/lCGtMIq8vuSxsmBr2B9
j2l9t2y7VbbJTmuEVSaDaRPkZitkLAKjRHqxKpwEZKg7mmm/9JuzCn5GEa5NF5EN
Txa3sxQpjOz0kfIM4pgk+AkyzsfW3HEEComLurXYlv5HKYHpZJytov2HYduBhJui
/hqPVfwg8XfegJA6s5XFJkS3AqbFI/buRTNAqtxmyOtxUmzfbkfJYIXKPSSnDSfp
i7pi3sV7KpRKsd+8JWtUyhkf4tpoM4EXwSXELuST1AZKWBVbe1T/K9FeX5Bowr5W
JlrJEAUvdYqQm3kZCZuGJXam5ms5JwVCLDirkj+DZKNHWuOACvZDjC4xt/BdBCTD
SEoT1VMsOseZBX7euEtcVDvppvjVo5I0lJx/d1d3JWTSazSIoQcQe/xW9A+GQpe3
RsQ2XZImFylXBmmRwAAUopygSYSaORuqLls3AaRQGt7wWO7rVLxuqu8j4r2Cciv7
xtusDLQ83tbXNoNt5eKAKoXm0D5IzdeHTqRNXIKYgyDZCMji2x5IzLOa2elVNWw/
EIA5jFh/vp+crCU68Pbalkege8cshyRAunj7k75n83GHjDjs+Z6aQF+4pd0x+AMh
M6hUp1MpQNPCTZ5FzglSs/bKPPQeP94GbD3vCLGXsZ3q7+ZgfhDJAxTiGjwBPuGW
zZrHatdnlcuwjqryqccxYtcAQuBIRpUcRIs7pNJhTlL2LTVd1YxRm/Z2rzgZ6VID
+A2tVVRMw3GYk2ZcWDt3gcPtif4QaPo0x1TJEm94oos1apSXQDW+z6KRZRPkdJpJ
qa+uZa2RplJjvDK+kkd7QY01H79NU6ljz10+Ixpn8sLPq5dMOMtsuYXJ8t28xIpy
JAkUMhuDldsPOarrWGq3CVPZOnCxYn8Ona6VLeZFduRN6ZRXqAzn+kHe63Op7CqE
kqQp4ob7pKtmj1rkbL2jl0snZtDT8LTyMokSeUtm4sOHroo3SOs+h3Tt4MgrBec2
VWNC7VivCm/OAoVZNbLzaJE9C4fFoKTLGtOhT5gsOnfjGEM49IKE+sLJmAoRXHpJ
VPDwspzHacM+XZ9qQgRfmf7blE0bMOk+Qcx1/42cuCS6ccSw9iCitmsAJ2/EfVk8
44S0QuzIcfNTVywKddOLgjrfpYIXFdpi71LJvVfU22brThk1nHqocXReMxS7zkxm
eQx8paim8sOJi4hB3aMweoZ1I0MoZkmdkK5DXB2fS02SthIopHfz7aWtCJDHNb3D
dROIX0XPDfZbNE8f40G/KNiJ7Kda3pP/wPpCaQ3v42HL5AMHqkOYHAG7R2LoAjZ3
TuhdBCmxzU7A5qCaT/eMfsJeYwZL71icwSRCtudWeXME+sqFTqRTY0aIK2QeGK/0
bxz7P9qQmIW2MQRTCOFiS+k212iZK87U6fG8OONVUo5p9hZ8bxWfAsJkj4iJ/GiZ
z0jg6paxcDuyJeqo24WLrOHQ1G0bxvW1WD5U18jY5NHHLG6vJEEK4o6eP6WHPMwL
Kr09lwZe/v4anD3HmLeq9FN00BK0uPbfeaf2Ccge5n+zrfq+cGiLaV9COoOSaJaV
pAIg7rVEVEEdBPY3sg5qs7bKx8vSStD0MTF8PXBimDepiDHNS+V0iNqAnb+ZseWf
25TsaIbtURwH/BLMV23cdhGx5Fs01p9HNw7kFO5rPAWM1Aa7LOySiU79LEUiSAJ6
CSY7dIC7Q4X14mBjVu6kmXkj5J7ryR8uCXQ1KCX8ekldnPccufL/jllnq/js7ZsT
DFZEN/bXnubnCQ4zaugzaa2Hq9Slf8sPoQEz+1ni+mTmLis2SsN+YbUsPL1N/kku
07SNxYKdmjJHkjYXX8us11naZZpwtkU9ZuJCWdii3z2Od9Ze9ZZgzQkpPfNJ9ivO
xGM+YSuxm8baGzofRrln5skgl2hG2RM70HD7bj/SSJv0emcqR5tIm/TgGl59VfxI
7x26YnPLxsasI+uw6ZR0ITruYp0yYJWD7XY4ZXNnhk64+e9hKuf1VxCReTH16dd+
m3Hvy7yQe1/9zkTaCJkpXFwJ5xTkrzARk4fR2zc3ARBj7dKKU/Mz4okx1OJ7pQe9
RxBWuScNLMaMn899C/w9aE7r2V1X/Vz6xZ05b2ReA9/T416LqpbWN4KwMsxJ4rEo
TuiIPKJiAvndRDyEC2XWpVYFupv6K5H/gNL27zCJVVKJdHgIEeKJv0sICM+ODRKW
6UGNLo8HXn3rmp28EjL/ehHb0WUjIYea4Qcxwmk2vtK2t+9WzKRXmJFusd9z3Ixt
A5OXm1Uig6p3WcP66yPG1J5Aha7Vgu9ZvuyR9OF7fES4piHtT5qJsxwIky9rKGP+
JYIQnnW3vbWtxNljOs4J0rZzCEARt6oyMWRK9ARmUEOlr19o0xhugncZmotv+kcp
OYLF0d9A0Ajj9pMTzMRscpLPQlOH4ae21DCb+/AR0HajAMjT3uxWjDWNrzkvrDMp
FYTWC/qEEAY6q7FJW5aXez/f7JzPG1GS+IfrCZYwG7pCSQ0mpWq/roWGEYyvBpUX
jHN9cdOXkiDKuNKVTwZa02os4KgVB/mFrbDGP5BXraxGGpfngedIkWecGkzFJ819
TaTkdmP66b8Ke0UrukIiXVl2agjD8x7eNpY6w6ClCPgRL55gN65YuMUO4LScPq95
cr++ZIfhoqiOHIHPXz41G2D8RxTZcNXBn8FHtVTMevSEfH5tSgopGT+5UgA8b9n6
6ArPZsquznmk1AdFYIW8BUbqr8KYu3LKmrZ6iJLmAtwMYYLBE71aDkmlbqU9rj+3
o+kRjHl7AuzauPz23sCnvqS8EpoCLFUiBUiJrJXJsk2LCrxLdZCQnTOkX/hyFLTt
73iDxlRVxm0sqBlXkipBIAsLvqiMXpjEI+on01YTcMcdz0qfZdc6QynPVR+H4t31
Y/aHsSm+QUPCO1x1c9wm/zMPEhbCyUjsqi9ajjCq58g1Gg7LpXODt+LBvrkzmVvm
qFa05c2EviJQBS/MZti300ydqEjsb82l6426rSaOUDGExpvv/SJF/T0Nuaavfn2j
HimIvgI/aSy2W6zWo7E3MGRK72sX+Yy4miDbVM++OTA+eqVbEqwjIgA2yd9Kh2sv
t3WreWgWAnRbIPMuuUB7b575EVeDeIF8LN6RVcVBPDIURodbXiIgWiastMYIS/Ux
WaykwvQvYHT1Q4Es43v0PA67Ulqj4RDHQ0tznzhED8HdnhduO3QjuYZdn0jJfmyK
zacfNSD0UmY9ORaqJ6ldLxZx5p7MxJBpLDKNzpSn8I8DTuedFz1Z1CyWZAbZSIvW
L2XfHFMD3I5HH/2LF0nDISdaRvgwtmI3fRE4qHIRfZa42TYs45B9FwmsCX5hvor7
XhVNOo2RdwspxpBoahheDVch1MftAMutlTE/AL8UvcIp9bEjEJsKxkwCHh2eMhSg
VwrrKw1OSYnxIsBAPjYiVV++dFKfjt+2RVeedZs6aekFWrSuIY7jZ+iEzKl6IG3l
hdE7YmHiEyOcwAlT4jOitOXdF8AMXc77cy6cs222SIhtM+agqlRZaUYZIZm3pdrS
8ON8jOFk+FHMQCWiPRxs+KL2MR/XAaCZtqBp9L2IN6ipS6AA45VI+LE7+GMQQccR
rV13mW1I+tFasD4AFtf3Le7soPk/fafPwMnjCRYFLssplWmntlyjD46tbRo99tIc
9kZoz/J1DEjR+XH8e/mLE4DNl93/K+BLTLhVTaWuKEOH/CjpyYcmxnJgIXNWFCNp
PB4nwv4hk25/i+cw8Lbrh1oUC3VHCGw/Vu5hVMGTPBtZ2idxv0+0cn5Vm24u/Whe
X736G0/TtluFoXHQtrOtfS5kVZn5962+t3BZubM0eaYuqRlO76PPiBZkj4pgBD4N
z68hdctGPWBDvXGL3CLBfwHR7Fk0EisIbg9LDUaJSgGY0vzmkV6+5MS2L5zESZf/
hPrn2Q0Qt3oYILPZm0/4J2EktEUSLuS9Cf4RompupS+DcTeJS+JPZULsZxevzxpf
ogDvMIj/RUxtq0OzdbDNkL33VELg827PuTo2XqOFXhZ9tPJU6WNVhhEXd5aTBlN+
eKoPC0C6aOWMB/YsdtYf5J02HBnA7JkwP6WMD4H/uIviw3/fK7ETOb3PNEnQeNG6
fDuzSEHMG8ZPrb+RDq9RUH7txQ7/6gF9Sli3iqgywqbPri+86Awtsu075bbHQdDm
ajl38PsKGt+N9mqgbkbA6UvvDaixhos7dy65ZDPHkYyZUE4sgqf4gW7oA4eXUt01
cMgXSFSAxYYtYpWkb5sYMwQlwlm5I6bGEg16Uywj8L2lpQTwRtCWJMxSq/DU/Dds
rmlGHygCxkX0YtN+6zJctK+SJMRrQzakfdyUF7EMZDCsHaMcDxyPMPDLRTvVDiex
1KH+eyLpWVUluDEXGCtbQ7z4YSjMp+q53z341UI+XELf9ud2KBihSAEH2vpHmQhK
eSZSrlrjrtfB6+cwCyXkIBhGTSfQxCusZbLATHAgiWfsPlD4QOp56Q3NOJmGIR2p
uR/C+0iw934Z5PBH2EVeD1qWMt8Q/noiBok6Ogp+87UGe9To1WRsMiQBsDiGwoOt
Hu+e6XhAqujJZxEJjdmPYeO9XEnrSg3NHmfSkA3BCH9utENL2rH9g9prnBks5Wb8
oNWTP/9VLLJy6t2Hbjpp047g30gekTSHifJTJ1lp444FMoMf6I3VG9XiXMQZ6Opr
hLnaD3vs78xtly1nWlebLb32KmhqaUrFAEz/MfDVzOLgjRld3vvQhs3aEPQx63uJ
jzX18HHvWHYu7+/P7+NBB+fjpCBMsRKOnezJD59Os6fdeCOt1agCoW2Ir68uV9Vy
zjTIofbQOn/TMZNmXzPYmNx/PCiu1AuKP9qCWV7d8gg561s/KDZn5weGApKrzbB1
Pg7IIVbA7gl/7NNbKW+YRMpZUay7ltq/+EvQ08RUhyC6918tz90Tak6859A3oSis
5LOVRP7KzmYD83UuCNatmhFc/mdo9WvYhcJe+o0w4c04TAQ7OTiHh23teHmgUbPD
Opy2Zvp1quKK3YKy5SA0J2Z6ad91YQI6Iu+QRja9cGbsZt4jeqnHoo2HfuaJ+Jw2
vrECKd9wvHS41ZtvjVHbcUz2J6nIM/KBDSuO2A8ojFib6PJDnjgu9qpDuSGTMdrT
Ytjh5q8zTevy4OibwRQe1d1MmUz9ia6m72dwJp/dL2PW38EtpybvCnfXNgPd5s2m
qC2hZ/7QSN+/oRy9li+lKa5XpLYglF1mmewp2t0wAxlH4zTQr9kYdBWNMZghv8Ur
cgcW/K2rX4LvUH7BHkJ4bFjTUGmvmcyqq4t51y9CD354QSHSrugYMF01CMp5LWSv
bo2MPH0nB+7tDbrrP2suUpHVZbaIg3LEyQYbmvHDV4SXvnQfzDifMAK8KMc8blKR
p2JsPoRhxcHKQF9d3EgUjjPESfVo7tr3YPk2LagSEBpcmLKfxMuVXG504hNOy8Uc
vWZw3KVmnIj5Sv9dosv+KqFIWG0cPWz111P8sS38nnxfEzhFczzV+Q9Hbo8SWXhN
oVNjJowsvfWfhdgmZ+Je4udY64webUQBuvWOo7pct7O9uN+u7Y2Fx0i8wHBwcMMC
/+upgA3iSziHa0n225FwN3BkaYF5L76Ig+bxqecReOaE37Wp2c+k+1BWYPvzdtBk
mD9cVyskGtcEfGxTW+NyGUc2LV4+nWvrq0xlLCWeYHvfsGaoxRb+QDz4fnhGa9X7
YT3490ty+AJGzbwNAosdi5/7Pr/vU3kdiaGBIy0tzej/YmsUlPg1Ppj1BpFaMtpk
TY/9V9S/sO0X9RIu2hO4SIsDu+VI3n4Rf7LisB3uB//y5av/Qp7baMwpe3l2b0aq
62Mj/B2hGmqHpISRjAA5aX+ssL7IyPxhClZy4Ls4lnCKkEfbYVYrKzOj3WSAABqE
vmpZxYIs7lm/mDZf4JtjqAhvfFECw831FnztK9vfGY7x2XR7BfCo0W9ZrkSzFAhF
ytXE/zrTraT15ADhj8tbe+Hd1dqKSEyEHTBZDRPkdJYrTiKoZSHGQngL11O5eYcb
8hAiB16Ah3N5vGsc/9hegSwokDUUnx6s/4wl+I7EuL8tDt2MzmRaQnoAqpBSE3QE
LP0CAoZAqnTw3P4vc3rAvQSMGjdnnlOTsebFOPOKtfssRuYQzN4zPzp0YSFCzgif
UDIxhcCbSwlNyLmOAFe5ri5afHkL/2fYSiNaSVrXqxkVWmOOrb8fM4GLS38h6FHQ
27mYh9kSFFeAzkNAfeW5XbkKVVOQiGMPS0lpkvTNesn7j9irl3TbIl7mDBxj/Npb
eKPYFiXR6LyLtjEdc9U/kepLWXq/jl7YRdJCzmBL2JW/AO21c18xRcwByb3aeG68
GxgSmDYDgloHMvAsyWtA4FIriLwRgxSh8vJlRNahJqCsF4BCza3scK/deWuQpO3y
/JcG1xgcBy/bcPBa01X0ESmiMbTV2jY1hWYrUYe8L8enB0sY+39xFA5zD+j2f7/T
lb+cDle8cDaLL6fmpucv/IaXslhvsHR5ju52WrJzoDJ9rNkNVrKR3ikW9RIz+ZOf
XWWqicLM/GloYqcTE4fmVqSfTMOLg56BXCq1OO8g9mcT5F4TDhnq309N0TURBcEZ
6IxZOJc8SSk3sHGIbz4jTMLapgXlbs1vvE0BvolCr4rm4HXQN4qZHRG9f/70fdoR
Ynzu4dn3DLwWf1kesJHQI5TH/lhLriHD2h4TpByr2KS9keHIyxR0Fv4LkYARJCrH
6BjmrJERzLtD+oUzxEOtnP48D7DEvoB/2O4zbY4exg7Ud8cG19HrZnddoroDZCBS
dljXKzAMBN/HpWEwbE9tS1PSBNunxJ9JJxfy+4B331APRRlH1Ir0DhD0ZEzWbOyY
5Bv72cAJBqmNcRqVBJwopPg3eFZjfmWhbOcOAGUCEsPWV+eSmpptS1F1tNYwDqEn
0VgGXaxMfGXhK8D7hURKlkTuUXdf5jhbMJ+yWgQ4T+4ZDmPLFVUs2CRnBKR5+GOP
tpeMjK4safV4cHjGjZG17oUVVaTQDMKAfWErmhEMA4ujpN6vVF746mTFykpf/nCT
wBIf/frspYq9j6oLh4sZwQpKYfzwvM/QjHeo6YxynUFLgFv74sOSV9DFM3II/6wZ
mcgnApAKskNNoZrwbaKfYxhXdu27+CX9Ip1prq8ojoL6fMp+Zg8eB6sMuaE6Qu7V
axXdb0jCr2V2iTQNlz7rpfurG6UyVw3i9k+wRCXVPKrDz/tfQhrYMid+akD0y3kD
IGOr92AEj9whWJM2qReQg7GiR5+KsjZjN9tgFw4pX+w6+MSfDTk8/qVLkv3nuJoW
B38MnH6FKLtvLL2bJo6rr4l2p2/ZopT98HsjD6NZSTRaq3e1NbfBpd9gCaS1jUVi
NMk95+tQjOtgE2FmxAKwqwq6rS7nDItNT+Z9DztxO4QWGFeJTYbFu36yDJnmmQFf
prTNUycjvprVSSYWmrVCXEDTofz1qn/kMlsxZLfn1HGDq0vrH1UaQqp8a2IAxcle
Fcf6vDlj9hQ4718o9Rv6WPwZ4PJYall1Z06PiKFKfNxzoJVbNw2aEJBG+GAol596
Yo00HMeINgcppeNatZEuPVaHlW7SFH5ptEWHm/fpqN8cEdC5AhfuH6mdcoBjsU1s
EvwCeSwVunCQm5aAMhU7AWYn7441FnMJoFkforBa6bGTQ9PhzDhV9UdO+X0Q/aiA
vAEJ6Qqt/o5+oW0jshYvAYriynNF4r/yHR3hDqBpV3uVm5AxptOmAnH75qO0gJ6y
py1i872RYTAgztgHbg7PN36wH4gRJf7A9Rwh7fNDDJBOBzYcezNhxKd6y/br4uPm
PyEMDPkjWwL7ORWXjXMxMYi/hneY+UKEfSWl9Xdri+O39clUrEtPk4CDrm986sVS
E+jVD/abKsaocpbEb06TG/pOUwzWwL4m0edCaUR9SFu1NfbbitO+nbIBI5KZ627q
hUy1uNs0ZH96MHEotuL5ff7oPXbfO9oDEomocfhpYdd+4qfFx5xTyxpkHQ8iUJwr
Pg5N6MZUqLlFOj/z2D8nn3PmTsLZf8x4gkTkYQ0OVO94Vkm+U6IpExAN88ZL9Czt
JKWlVGTLJMEeXn7Zb9p0VUuZuHKg5Ja59DOWTo0EADWarlSEXXEtB1mUFiihLGNb
WR1PhztKPP46MDB5StLt93lxfgJaRERiQVSt/wtBEPekdNZqxxpimI9oeuqgBT2x
8jnb9iGG+Az6fGilQatzwoFY6G61PPBjKQ1qkP7BkcZT7qoOFwjuHJKvF43+SSoR
/EsEb0Eh2Y9PW+hcCZS9jmRwe8nRxJjhpV0lsGJgrtsGtwGQCl9G7M+uDdfN83nN
XyR8k3KXf7T/B4pgFRQOMcvjr5g4rty7bkNpuoefk/ZGNcImS2DJNvh9gG/SvYed
vb7Ry2uXJTpmEzn6PaQ//kckiThA3TWpSnHeRO86W6VX/+cgSYGiBXpERCS4vzmE
nSbezFBEBOoKlnNLztd4N6AbA/xM+eAb4eng7d1vMWS9J0kFmDpbwU2WUEVeJEJm
0sY5dlFnuN2e3B/v8Kk1Ft465ZzSU9BS8K5JmzoebOQWS1oHttO7GTu62NSwBiZn
4mrTBWAGwlCckCK9otKivp5ZVRzIfSVIRRqEhC3zVmSa8gW0Ev5IelbIUTSqTMF0
vWkjrJQIB7K6L17Gh8FmwA70zY/OtaSCZGmE8JBaM45tBERnbMJfGqyNf8Ekgwcn
bQm4Sv1KFY6xPc3qS3xnmWkZK4K9RCyqzgPubZidPrlV+IFRbYjc4iO77dxxvB5D
UmyJ3sjSG6t9T/w6XqbR1Wly4A6XNSW8yPG82S6LFnCeD7KZdRyO35B+ZCGQPykG
epXtIgAbBOFGH+fRQ0k3ELgxcRjjTI1DOsCPCAo4KKLFZDkc84uOrkGNHYNy7RU7
oZWjPSB3TZPwXjGFtHp545WJyFCdRDhfJt10Iwrg0B3sQnIj5fcGyC/0q1zt12bx
WIRmYz/Jz/nW2jdev3h9BBxAZBpWldembCcTHdRF5zRZ7WA6szmM+YFewOhzg1Y8
Rrfpvl5NJaZbWBr+1g7a/lcAM5MfqJ87+cXtIMEWWRzZLsNl5CfEWWWTL3yZdLsJ
eUV2U1y4GHmBgRPh7IcNRsJXL9pLNYGhKHkPW//T+lXpSPz777xBahKAsPws2b3f
8eSFW4g//kciOTAOPDmDhbClLiFTDneRBYswlOChuiqLuZDGDoHrx/ymbZTdQizy
jHLg/n+vWmvUuulY6DgWUR/dV8hdh+lPsYrHdNIssnIv7L6Rr/L/XntssEDJT+bF
UvtIRKxBofyyv8+AsjyENtXFkyhsn3IwBxgrlNftg/vDcAA7sM7HmCY22IN1YQye
3cRqF9LdHT4kCZaQy1LLgcnLRm3jb6rMWbLGnXlHKOD0bMQ8tozeW6+i/zIDWXHp
0wIWV7IeaMsdrWjJ/Rbh56HEYTbr8oLmoHMvu+lw5376GZYpWAVCL3nqQ5Pck61d
z0700C7dF6gRUjGajlKHkFejeBHMBjOAaBYayhUfL2gXATBb0H71uV8/QIEO1A9C
qhzL5pR3ny5S1a1TSsJOkJppXM+X/RqAb+YAZ4sXM9XOdst/xvb5+TWK8luv1hyt
oOjkkYQDSO4gfZqdf2FkVZLZbB7W6h/jhhXBbiVGjOS5e0VpzhY0bHmcZXKJLUd/
+V/nfNCsG+cPocvUttUtZzvDIL2+s5K7RT3TQIEBYiey0XsiFzZQ3fOSr+aHkVEK
3lEIXIUXohWCMUySvBVcdTXU5FI6Vvw80LgH22QiioVISDLfzRBFWNercpGy6RsJ
wqSGons3uDBhnd0wjU5VwadE6cDFpOxPNPHD8oK+dg7FnuHpWmXkk6EqVr9lVyrB
Gj6Ep4/eVXlBrm37Ts1Wq1MjcjmQDvQ6QmvQHCbBYiMp2/ccOuO1f1iqf4lR4Tc4
8WpamjYq5fgR8BRZhZhY7Dfzye6Amdrb0CXDelPcSHaNwjWAjoxrKX45dMcHvoKs
OtDQELstkPDnTHDSKXfgvKBNhOueWsZcki/ZB0bxRVMOROsqOGPg9t7X7oP5uMNM
gIajkG9oQb5Tup+Tmq/hbwj4wsw83BweiWLZ7Lz3pbiW7HIsGLl4oismW1XuleIV
pNteDTJQhs05Q0YTyuvmjMhO7xh1eAiIcEvn5Gpvk8eq5XRVRhmardfTB7NmHB4u
bWYCF5RjBW4yCkoNTej06/XkqjFmNQMx31ukb0q8hx0LsH9vBx6CG6Tk2HVK9Sd3
5l6oQLOU3yjKuHLQMqdM8v/4/1b6jBT1WyqJZwsQKx/AC+ozw7ODF9vLxdQvcGPC
EYRDw1mT75e7MY9/Cfgh4psY1+eM3XZ3cwhlovf3fbx9DjDHG+bLNym9e8om8ZU9
k4JjH9wRio6cBeu0AEbQjTNMvpXJRsyQNBb45R5zGLS5ZlsrqYSy1+FEH/pg91sI
PLlJx13cQScQhmXARZO/WguSpjWG5LtncYMCQOGANTLLOcbYYEyyDE4MxfC/HQV6
byKtOb2nDSO+MZN2Y4VHBIaPH7lmompGSV6+7JY2HT45PB2YwEDmpN+yA+0meqzo
EWDLbRdYSZEx9xQqCSnUVXCo0sUEmMYIl16MqKnYmqfkHzi9ncmtV2bbukNZ2vK9
t6VRvAO+d9NUwaD1Tc0g3qBEIWm1Axrs1jd/2fQsjoUvnQ+kLy+TuRgYJh5dSSW0
h0Z6ozUGuZtxpV2u6QvmMeOC9Xh7SHIEwVmpPxcw5t+e6dDGpR/JpZwEihNZfDlB
xh2yE1eUuB6T9dyl05hCJJ1YqO/gA8yWKiVifIywZ6EnwK7d/8VumCHtv+FE7VF+
erUg7jyQ5Kxm3PZHrH5sZHvV5NAQJ/xyPV4Tf7apVLIcISSHBTOntYkQV3vrNM3w
iEo2bMiCzMIGdiPeZFCYJbKBfSzhGPuA5vSqCGBVdHBJ23IxJF8i66qKE4IBL2fO
f1BysCqctsF5udgFIO/AMpEy1d8q7nfv64ROsfUDnUXb6unJlUcmJl6HFXpkBUbl
Lz8Fqxby6I3zWnxYLyvBO+J8ejsDIrs0iTfRnFHXNp0zpA3zwpC9cVIJ1NHnfcFX
Hsk0Td40nZAT8M7SJezRnNN5ls+w1+aYONL3Ga/wpcehuq7eObuY8BFkvQ34IrPJ
w5K9YbrQxTdgC9h1cRg3XxTjM9JKQtqSie8wKLPXO2st/uRnCUsIw5j4DoflBQzo
C6JIUOLd3w9IcarW0N7lGR43JTNdkKB2irfOY/xuj/eplz0FLGkhg9mOON2QKVOH
qNp/2DeGIY2oOhL6Cg/Qk8isBM7FSFGfQtC3+eZ+TW3Gg6nilynsWAo8XcfC3XWJ
+GFxX9edcCEVM6a4xAXspw1vILnKBSy7wEixlxerud6X8QiHPAO1PY1iYCdR9/hM
omj62SlkuopMcDaWFU+XZgSid1YCt620Utpo6GYlefiTUAd4PUDLujtENDPiFSgL
wnbaKqk4w5G1tuSD75WfInta/qdfrpLuoRZPrBOeAD9rmnnqY5SMKnsVAvdfbNkg
dALC+bQP7UeAmlarEHiMMRtnyo7juswLwmW7X8OvaDKKRb5ApFmh769CK88w6Dmn
zkTod9nYom1t/meOjvbu1gJg+9iZF/lI6BtYk4pKKffdm7fBZcWRk6+uzFbBijFQ
zdg4mi0KH1kjXEd3WUhmsV79740XOuucGNb3iRBL0ayTZwziiiep9KIz6j+hZirM
FS3Zd3HAOKy03PhDxsqx7FlwryVd5uMxTpsdgt7rryIvk/aIP2dAa03I03Eq9OVM
XzqWH401AELRdGL9P9Hb1mIPoDGpQ3sUWRy7UJiYB7N1Ho/gs1yt6fNbVTTsQQsK
jsQYuEN5heNNypDWV2DmQ5WJ5NzB7yDfW+y95v/n0wwnPBR53+dgG2wnLMoQj0xN
8dd3KUNmwWbhDzeymYeiMzezLcdWRvjE/e5hgD236cCyoINrvAtKowb9PCtkSv/O
c6crpPa4k8UhwNvOlOVUwq3D11cPEitjjc5ylLboxc2kRZJwaIEBC4Q/xSExSqoO
mRnX5OZj81AOutAU4e/vufJD+ozEP3dK+48LiXVxz1XgkMCalrj5nLvF6yBn1VzA
mo3x5T2mXQMLJJ8B8t4WTkHd0hNxRbhRfBBaprC6BK8yVpSXGwnW4QRBs5MXWmCG
famn7owZg7UJC1ANd+aTiH3+1hoiloLgxKNcG8dKQQ35CPFCtBiMGPNwvBwoyhYD
7DHh+DtV9RTov/ig67dTXIRADUplp4HULMy4ze1U1ZMMeYtmGyadfr2vMbh3BOtb
qyAWo2zfpSnorTxZqmh4KEAeubuSqBLdvk9IKlEPwrb8NsBARYiy1sCOChapTMSm
97yHILP0kHzAo3PKxCFxyv1bvC+AstCqi1GJSR6e0va9aqBDG/5JuvFgPRuAa5Fq
DKohSgFlyOHywUE2DR7Y+A9OX8BPUKiKQbyT03jikpsr9Y0dlpOorWpBWsGaoNbv
KzX+TuE6Kd08xI+AegYBq+O+XgHc3KU88B9YYk6rOhdBP87G0jrzTNDqKAPlQoA7
TcqhvfG6nM4kpTcec6fJOkskxlIhM3OylplOIy4bTohzrlwCPh50R8Lrt8oN98AO
XXCCAEyJM6Etezhnd4Gh+rvgYYthDanjiXsEBq01jYoyExxCE9k+NNFIC164KWRX
p0+DJARm8t2QsXKPyrAHJEjm1e1KEc9x93jzp2Vkgj/uRsMyMRU3rkixznqgLVw6
6QqoY1HwIHNPu0wjiGn+4KU64QPQEzLYhx4KMFq/t+sGIM69Pt0zyLuQ4+04Xq7K
tmog5ousxlIgbV2B1ahkeEyRSU4Yh5SdCYdjxloQYX1s8Ljti9dBxY5iPJfIAU4t
OZBjJP7bxhyY75XIaJsuP23PnCYENGgpwHtK+n942QHx5W4n9wg9rMhWnJXATTNK
/L4uXEVyKJo0NmbSI+COH3DgGRjvyIEVWJzL+xed13E8ZX4/SORilERyLBkgGDrr
uFxTadLLHBEfBWOkHAsQKmtUiagvU1wBQYtHMaT/bVOPztVWCUcYrbvzbszvi1zr
3mJFEda/5QXyVouU9t8BLSmiHpwLGX8pQPoAKD+0J+c8EUs5yjTdZBv4dISpPAWF
TFgY2ISxN0a5rGcxSM667XATreScYLXhz+OCAwf7Nd8rFHQb7Qbwsn9AQRyXyre5
vqflmkuIB0850KeXc888nY57A7hZPHC7rI2WLAo7Hqr4SOHEXGWG2Iy1OX8w6iOY
X2Gg2xwh8OSTc57aXS1111vbCREkuO/iLOx9SSz+H2nR0ixAjb3/Us/TWP7wfE6+
bPbnSLbjHmbHLEP6Qgpv/ufcbzhOaB8Tb7aX3K10+tUck9YFwG04u/asCb45xGIS
7VrUWYbxe7d8zctlJ8PKdeA9GOwodn05+dvROniVIJnKObq5gpPQNIK+3aBW4u52
FPqJw8FEnw+53+vxtZNYSRTp8XwhK6CPQ7AkQP9n1ZGCYP+lcoV3d9G6hcheuXXt
aFYADQadOv4bb0z0IEGO1oRETmfuq5hsof5YUL0s2lL9ad84aZduwLqGBClrk4qx
FvyxXTdIkFs87f+fq4K9cS6cDHnkR6DhJaHXztY6gzGzC4NwtF3obLb7yF6zuq7Z
vvy2uAY5pDgETyaS/6WmBgOKijPgoxXyQbHxLJYaHqYCFglY0BoaQYXPy9zQtpa4
5n8rScvfKwnCrCSSnCwYReI4p3zdZM4Ar7WM0SZzDENH4vFSfzEtpIxq0Cl9neov
QGk4pH3spiRoYKD0QsQattb4KJO1Q6y88sIJ9S7CR9vp1QNJnY3VxRe2xqmywLba
GoHfpEht4/fYZncrCn7sXU+1uHPYaLjUHlnKltH43SNZaudjxaxBU/silGxyFBnV
J7poYB+2ar+uI691DHf9wPCoesq/MI/2I5e4Tp2MVkFkFzPkUULXK6VomLK0RZwm
0svMBz0+jvzHLP7ponqgcqpV+ZLZyEdlkNtCSmaMNYY/kmsINP/1r9ow+vuj06bi
sTWdYOTx2I+o8nf7qxT29eN+6OvPcRud2ZF1taP4RE77/QGtp3JBHpRUMZq2mJ3/
/c/7gNDtZk5AjEb9/E6Occ/G4GJRuNs5uXnau+mB77oM7cjlF2HsW8toQDaMZa+R
Cf1GzE9SZy5qHqlpCEWSjICli99B7/69QqjqByvQ+0k2orgL+cvUIiaSbDnztR8D
GVdbMuhWiT/Kvm4eLLqJUJ2BwHIB+jo5ZCqVg7KUHAGEyhPQbvOm4C5fE8KvceZp
ckFk1AaA5vzlqxbVXsKXhyg8DR0RJQOQr0fCI39F6YiUnjvZRs6BE+qXAm9Hwl1D
qxx/a8IeopSlDaa3vGC1pxvAIsC2XWdVBhQdy9y2yZZyLEjF4hkSLBcU6ybQCSUh
3tiL33oD9qjuvDkgTVSJeNCT2YYJH64jXbDRXyFcRLNp47PYNhenBt8ReLQoS5wa
Tf4sNdnF+wSNGzAGym+T2mIz8dBp64/CCPhld4900CBYivzNMUXxLWoiLhqiRmY+
KpeyKaSfmDwrmLgL+MgP0cnl5wA6CN74kGGqSddhrYAo55in801kTj3ro7fXcYIE
uvC4k9W8qlUr0HeTfePDtoh9eDuAxVWxx/NZaGS8/bmAmQHfsuxm2KoRE9Oy5Zy8
turdKBjBEIbmT6EooyyGtDHqh8VK9sPmGYEENYtoCu/6Fd7OPMwa3MqWdUn3pdFe
hdfHBr1bssxMOzSiKdxBZskAS76jBAHWSqKC1etdYnzjOPzVZRVC0FuaUBSC40wC
qX8jOmJE1tpxw4NKFGVAHt6VDXsSCMv8910G4HW2TzqKFKgx3/W0uTV3DMIOshEH
HAYZ/RE5ASoV0wnCWB9kjXLLCINTklKDP3PJX3pioi6mibKcM9UztcMTUZ71wewt
G60R+k3nR6KewnFR2QmvvsFMF9rBSAoQrYUd3KqtR4m96n6rMV8NVmEgrZ/gpnsw
xg+9hCBBtHDujty/Agy2yXvUC+IlBNhi2EfxFbHs8ImNgTUAhuAtmsOuH8atH7sk
4Z/J/dJfzvoU7AuVZmR9yQrMVmogQLEI4qQkbWPTmwHNa8fYMuG/wMsDDepdmXLq
exFXo7OKs5CdBZCxzTjs5RB6UuqeQDohc4gUof6QsfRVPwHkGS7Z3XgEmRWqg4YX
4VaXFDVOwHvl/Ol9wlixKtPr7p0UIYzMtD0vG++1VN91JC8T0MtgQ7ED/CLHK/jx
UdsHpx7iZ9DnvOd9ua3ii5+1Y7epor4D+IdmhJnl/743ZMhWwK36d5iRp5GST6ny
GVEPJjkiitH9ExjIpJx40pG6gUHRuhtRAr5FpFu3mzcJwEJIIAcnplmIe4bLSQ6M
W/UzGXDUwNTSqJQlVLliX7jt5hVsNaKxFfazdDh21Ka3gFyQig4UOxy1ny1AhYRk
gYAchduRQ05HErLNu60cWQkLEaPymhEnEnDDHgYzXNAYYGoQr3LDBJRBNXNQq1E6
jNV3ISAVOvFj8OPgejULAaVUUEB8zgciH9h1MUw8lO67+Ms5D0CuGahgE8WWb27S
zuL2WjjfMb3rMTz83G06ZYofWBL84aA3zVHrqmS/YgbJt7fg24xNkBeM+KMY5zc+
nSdVcK7ZNO+61BIGaqrgwFmVTyElaoKGZr5APNEDb9yDMEqnNnzxbYCl567YJpQ6
dnsh57Y/sP4oN4Cbsmvr8a/ty3T/zqT+ZcPPY9L29QAh3uKoQZxn05mQBROvA9Wt
EzAgRLr1fgkuGIiqHEvAfuUHjeA4FhpURW2Q6FHQhtjrlsYCBscCA1o1ON+LAjtZ
QuiQceL2vafmMlTYHuM1GdXu3DPq7dsNeN+0sJtiydmAQGdS3ECQSOOzPkXf/dq7
edXAyLBEXZuKA6j19nZrBxTYJw/pBlQAoZYz6KavBYBW/O7q+RYGxZmKT7N26/U/
MI6uaLheYvEgIAFVH4cAxRJJ4pEGt6ev9FuQ8+J+ROE4l7XDQinn+cSq2KkL3D+u
1d7dfAqz0woIHmkyLYRYUbkmtR/RoXqbOyPBibIb6fdR27OZqYJi/4lxcXWU1RL1
MzggP9p84mOERpTVie2pZ9rBg9da3cBxW1q/TWPTqC6HFZY1V4cXrX+8GL6hfc66
yljDk4bmtydBAex46pxUbSARbgrAtYrnBBYg6vBV6N57x2BRLD00HjeNZSQPiCer
zoAU6OE6iRemlmQoQq0F2B5nt0SCx7V3MChX+Qozdb2hA0hCzxBCT39mbknaCUKv
K779hzaB0HfT9WjR9nCw9u87YENSX5iNU+3jl+Cc8LucM+CYxQlE4SSyZR1RQxgw
7kDFhNIQpWF9XywGFWefB0QL5I/0D2exa03E2OR9EhlHrjaN77oCY41+LYIbV+MQ
fvdgvq4yhMczJQaReWhoXGS2coA6qvpZP5oYV1d3lcDLOvgVE5XRYHXVzasqWRwK
GjXUsE6ZiSDphSAOpqiVP5hwrt5lhlmGRPKDbIyS4Pdo2/6CrdR12f3j2FL5EZyZ
wPaJImO9ZIwXNbkPoArZechWNtgRLSxjaIDVD9oFhamd2EjDt8sq8cioIgyLh6yG
i4GbNJkDZGe7xYHvv2ON+Eop4BLuxkvAzgaEgWZX4EA2fXpIKGmuTpcsd+FCaV9+
ywVVYNHCBrVvwL/uZX1P/D1X2WWR+9iQ43OtkC4ACHd/BJj9erDUb9EL7KizAdxt
cNI8pzQSTLJxoMlK6P5sK3O1B9Govmrxem4hSwE1tK5tQZZa5IQRsaYlfMA5+77w
53U5AtjnucM/OcKahewEdY/x+oSkb0ckpdeX2nZtlZQR8qAx1gx+pjGeQJzqI5bo
88xveRvH+L7wSH8ihkvgro33C806zWzQ/ZPyAsFEdqRJgQoeaiOfjaKmLZiMAl6X
ix3M7fEZZSk3VO5w0CNGQqCzGrJTTzplkwBHtY0Nql7D5tYLhxi5nhjitBfHDBvZ
9Pfyidrw9zDY5UWUERBA9MbMWVHtKlVJGhFQpToMX2ihi8V8gFUK2ZtVmyJHtvNL
LWpI/9HRfS8H6PitOWyls3jZtXLlOW63glikDqYdoWZb67eaUU8MrPwqW0XYSv93
GnueXa1uDSTpa0d/s91SxojNBq5FaY2Fo7Fl+GAlYsOdKcmIXTq3hwTNooxrIKgl
iYWJAkQKsg9/Y4ahG8YhPe4kbHx5QgzNtzbQxfcniLMlgwER5nQiYPCXIP8M58Ht
T6KsPU+Z7w/lXcE+SpOq4AYLf5UT5wQIUL7tzfEt3D0pUcSC+XWLo3FtvKXmL3Vt
LMlXZVnXEouA91A9OIZIzzOxSbPM+mt2aQMgZiZHG3S/5J/LLBXCH+XFEGSWV87W
qBaIpMIv4jK7GATP2jgKoDKMU/CX+6d0aIssKImPh8UIpQ0ptwmsL7fkDGxGLzzV
C/I9iUZch6a5G5Wm6MgNSdkwROfkE9Y8MhqQh7H64v7kQpyPS6xQ5cZEd/MWaQqg
/wNFMCBiUO+LJKhEoh/26B+z/yslfyPGcsPNnJDETrwpo+S/1grROEsEttodztnC
tViXnxumO0fR3N9Fsiaop1bwrYlOb5NravYkA17c1fzKjGfAxWTtYOi4UkzFDUYI
gQNt8VJ7aXH8aiGR6lCNRr5KZmu6dl+cg8TSDEczddc/Dwimh3K/PN71d2v2RJ5H
fXiUobm+XwgEKNl7ylF7XTsebseG0z3I5bhzk95YzsTOyhx5EOcm0PT2U3jlTEZ4
LvDfTzdagosA7KzPzeWEGNtBzqq98kFuVVFz3WXIcTi0nphI+9EQ+ZzoUGPc3Fdm
iWf8oq0zz24/edGWh2KJipyClLW0EFU5qWeTUFFOmRVJFo78nSZIhDN/RKtcRyE/
cRzH1cLevVMUySEKKt4Ot4wuIauFzYmpW2JDD9E0PhfZbZm0oaoYmJBwLCduzWLJ
Ks9esuPSB5BLQx6VCa87ekv5ySZRHavB+24x4z1w7imk1eKNIxAGVUopjpmv3tHu
F7FvDYEljIuL6nlc/ZerdcNaUqThuzNwVeiub1GuTAym37iD6lHCAvS+i8oSAaBx
Rts4/tED4Gs358e1WfjLjqGgBWQHEfcd+wh1RTYZYRlK98oze6OT3FKGOwJTMoZK
xWeHlieD6aZqNy9+F5IU7yshLbn4PwEHcSKhL37hxocKurJTggJsGKDlH2fJWOCA
PYKGe+akM58W5drMrjgpbY3VSj4Q5j24YneDeLvfcjZQY58DqzPOT0/geS6mH+ZL
T14X2rvac7gfcttdasPs7CFfsRyy2ajlVaoCdsWLDnGYVckvaSl3otduZRcaEJoT
N9DNGA/rxmnbz5swi+BS4sV0+znhmncLtBWxJDJR8XAvc1pREQwFaaA1+1JYCL+n
eTAhDSxiFNnpIhj2w7k2PVg+ZKt+WX40Uo/qtU/dSR0TQjfPHNgCm2WT7x0qx/v/
wqBjFiSx/P1fJZux087+63MvlSz8nWOAAEIDhhtq/CJxLxuxmaivJXN73yINIS8I
wzW/61yWIZyFmbnD2Ob2NEIjnz2Q/XhRLTQA7/MW9VSw8TCquK0e0HQT9ZXZ9sEI
kWZaV6zLIyWMh/BCiSKi3ZtM6ptFCylN8B+oWzTA16X0ua9hYeDymCw4nzTQyEVC
1mDYnyoSRK1WLIaoPuf84lsrxNXuvL9VOzszAoz5Gpw7xi27XjRdIDsUZ1LiKYYA
jCP6r0Rg/i72IydVf6AyXqH5kp2kJa9i/AL30mwxUWYBcqwZi29CEOgp/LPCtGdk
PQeX8fEhcww3ntCo0dum9Z57PxDhM/o84DmrPHDLtPBW8zUeyhGhxayfoq+bCesx
o6gfeSeO1ohxAQ2EBRZLr/U/7BmmJ8guPP90d3tf/yxO74/kP3INcmhy260UDppz
M5O77TQVFig2azghiFRpg8LZ8Ynn3M8wSwqtZVX54/r96ZmrrShfJI2GFRTBOt8C
txLEyjNvfwjJlVuR/Pu2fJ3z5+fzkkr20VXPyRhQFf2CSCpVLlgojvwN/NdWdztw
3KS8ssw/A6Uh+RDE6mdgIgNucSH3/bQP+WxmT2UldldeScO2lJGGjeSWCg+zUhZe
HeYDHjta42w0OSTHLzcO+/sDHwOBgzSHPB3pybndFKokttmhhAarWST3xh7WaBVF
sB0suFp3ptfc87rz/NFiXDuYI3HK81lJ9YGajHTx+1iJSyyfA3NwO1y2PSHisXgw
NLh4xoPaWd3XEK65SxH7VO5GzIG3XWG3Jae0ChIqbxBZ7U6zvPxxExsUzPzv0hSK
aoxDAMsPGp8zGIW1/pui8UHnqm82KzzvUXKhX/7/Wh2+pRYRHDeXrVPnczdg6CZp
2q26B/E7cTp7MRd+lJuwoFpFiG/kdhs/tthoHr+q+RSj6BxqY155y52MxazkX921
lRepSMBIojUUKZDxnvaTi/xUyORPCqqg2u12rJvmHIr91dbVG6pTys3foLiiUQ1I
pOPrCnaNyt+alXB/fYQVRvFckKTuka0qBlPm/zJLXEYtEdDYGOoid8Ub+eRXA9L8
aDcEH+a7IfVvl7hrbajkf62vl+RAXJgTIancqfPDy6QtyRYT01vk421bbsgAKlTE
d9ugMiKM8PKhR+HhDLoBLCWbXHyyGauQ5RA1lXwiyos8DLXHWV2j99fPfb6TuJmk
DCfB7xqbjIdoDwksgypCn8G4kZVdZ8NJ1QFHmpx8tlSwSmcafK38Dh1l//L8DTGr
xoKAYdL7N8wCFdofsbbW2AKQLu5eBp+GBclu96D7HizOBM4+ZyQQS1TJC7a58/00
jK0cmb+20kPLh7dORyCXC6VKZxcsxuapkmPTDPN1MSkR8UyrtOcl/srEK24jQTGF
nHXgExRsXHL34m9v7Cs/0oQ4zYUyS3Yy/Su0ucPG16mYOyf/nPHSsQVONlVvvLDo
5Py0Ip4tZ0VDXTE89fnOV4TKXPoN1/QqK4Me0puQkwDA+krHgucG0JyigH2I+9Sy
btSnrvvsbCafBdahuaUfwI/bs3BU2bMz3LmtHR/Pv5yeTWnF43WpVU84R+thraCL
vvMs4ECWV1wPqPs68uUhjSIKicaRSPKiEm4ZAE2CG7M+lLQyTbpZJgPVmqOdyeVc
kwOKElggTaWfL9PjEaCHN0XNdPj9Zo77ejF/3wFuoxs4obRhMfUinLrvck7ad6nC
iI7VOw56YeqxMjmMZf62w8B9n03t8hTRwNHYmBlOWykHwcqeyEckV72f285Fbv5/
TgjlSXQrXECNzIH+OeqMqbK/JvplB2vz2HSjXkSux6XR5nQi+Z8tfPZ+CqV9ecaY
We/Rd4+/8PsplYLhvlkM1ofZ2VIBscV1CCpA1XnuyzPvNCMBqMTsNJjEA1Lqt2P/
8N2JuEs+f8lXChizzjuKI5nZhYTPsqs0juWNiAy/Ah8ZyJOAugxW1t56kHshA5QK
PfTqhawF5h4A8W7T9KDE2ddHfPdoXgsP36z6poDc+JLxLfpDPh2qq+uUeE8UKr+e
pVF6f+enPGN+Bn15L429YYC57lds4kKfEO7SoFN1gnGq135ViNR7OeVDYePMQGVT
yzVJ6y0LUcKN7iXsVvYRiiNDTee8V6xzc0vhFVCwPlBLMSRkXZdjwUFvStbdYPWk
/SWfgk6lUA0wpu9OTwZPsxmcGfdoUk2YJxmQtBK28qja+s7KmIrUmyJR9dSkx6/y
rP1rd4bdwV/8kdAYiVNFc1vAvW7tSmwtfpjCNiPmGrgrBDMGk2ZcES1XiAY8lk4a
7CQjjm+3iQAvErI+mMt28ZCPeDSJvwPFt2avkKnTBx8+ud83UpOeRTE6qEg0k6tb
cWI9mTBIbuDC3pDxPaVXwpAPWroKQxz+eeOL6DRsP9m2ePQOeczYky+rU7ys+6rl
euv4zOhDtUXDu49UNPCyaHlafJ4g2EIl8pY3/yNIMKGfpvE4ue4CBdMc40GPU5iV
lcs5PcxyTk/gRZHr1FwK5w3dm/H9TPl0JCF95vrbx3QsSYguKA240vRbK+Nxx9sq
O+kjY1qHDezm5zsDdMgONcwR78aAMHpUsOqZhHvSnU8IkuF0S5udSRK7AVwbnqgB
b4S647lRdTdL5PlRnoqmEr/D2ccPp4c7vK/n3EJ/ZiPTK5xn8tSQqXNo76cbSQoE
qj80/f8hU7Kq0WP/2CDyQvZiN+YpuVN1ublPpahxDOmxf7A6aPvta0bxtCz6gfc3
J9tnJqgSlYdOqJKwOlADWyeJhu2KgwmIXg9Y8wTIJiiG1wuOBzK4Ntm4jOoYuzAN
9hK6PV9VIZKm++9harOYeL0tM/dnHsNuUVOiYPLrochOfC/aTUQgkTxX8xJSkZKZ
5D2hHMyOmnpSDR16Xy8fAV4+8L6S1tTvuQXmtID1N2eUo2GJPVvl5IbHYfJnTht1
JP+CCGFP8kraH7rYPpeDji/GCZHMOU8UFsCsCC7YAugxPkL3sElt1g2xKVaFqEE/
dg3Fm+9hEO3IAThb0LK3z5c8AuVqjpzvXCsOZNZ1pHGEnLpc7gh6i78Z+BT2bcog
NMdoL5qx6qu1TjzEbLtm6L1TuDwGENHcbdkfBidguSgdX0Rgtme28As8jiotWMI2
ClXxeV5dPHqwHFd963tPIWyPabAcfOCvF0EI7Ff4NM9mqzALLnCBRH8x5hUX2fHI
hBSPFl88MN6Sm3Fvf4aryy+7GcRjm2rJekY3Pc45XU8zd6ExdLsc/RjnL4Agcvbc
a9bT/EddAof6vzL56Tnpz4Vc9zLBioWan/h3fMGylCtLLFheGRDkXAy3qfG152tS
ZbVcyoGDFs63x3YXPFylZ0HWX+gWzthzAsiujM3PL9Nv0fugM1HzZ2dXfYtikVAc
i5dNGjDvbMpG/uKBTa3QGL9HcUUjc9EQtL+ynD08bGT7mppge14+pVM/CTR6Bkss
Y0igtTFB0808TdnnSSCY4xp17NgZq0lhJwNMstch92GS5JowHVyaeYAlBePj9ZWx
GYN4EiVUnWAhH2tjreVLYyF7JyL/p9Da3xZTpVrSp4+UlVHglAMIb/x1GqwNMRgj
Jp9lnZ0RU4p/3iFKdW/FLGL/izciRpA5p25xGW0Y0mAMeiDAemCm/kGl/L/cd0KA
CKJko/I90M3RLw5/GJCUrOzHCw2FyE/uakIj40Bc1W2Fg0GooNFinNbIYB+CD3LA
Vo6ocsc8C2RA3AxQ0BD6et1uyhWLTWFSz9z+uBL7SSKKOu5Lt4ZS3JyQ7HYldVlY
k5KPnIwOlLH2Rlw6DazOh2NSFYUQsR6ImONClYZOtmir0CHkqG4lvYRaDFVaJo8h
OLLfGtGa2ddvTYx6QSs7P2zRgzZG9gClkGruK4QQ42JmzcALYwreBSOzscm9im1S
K+SZrArhRxZU4KkrssxlDwn4gTng7a6taAkRWTPkdveQL47Gz+zBJDURVHBVlBZ6
k7ZdyGIX0T0sSwjB0Nh/FRGZ05EdTM85mvt7AOD7JgUI7Kv9cMr6LQKOFsSje7AT
sccEXEr6qgwf68kKOgctX0bf62x8qceuszVKMycqHSN5Y1xMlbVsPB7imKL5lE/q
dUVbsdOukect9zVfYG5BI0WEobnbXDquhbCTF1rqq/2X6lgrtAFaG6bZOUseRTEU
6cMMhKvCiRj5CE2E9yCxpE1a/v+12lg8c2b/mOrX4mjlX/Ue23kGVSXKhe00T7hU
sJeUuD/iuiYuap75ny7LKtNG299KesxVUlaRAI4rHRV//qJjAMGYVJpWS/iCBgU7
9SwilsibdVprpYg+uqiiquYQw4NE8jQIlos9XkeT+V7uqMJN9ZR5r9VPryzCsoK6
st7jPDGnb2OquwJtQ3qc9fY11CjkN66KFWNgYlGSbjjeGx7NdiInh3iV8vJAob+H
zFdJue+f6cjnc2Yn0QVNlDFKPES2Rjsp387guCdsVwgcT0T67tJQJefNfh/VL+tx
jBnB4/rvVCmhLlc1tw3tpp1CpqENINvC4hN8vxQnPnHdtMlfPXi27ymLAd8nQ/sz
4TYG2zFPWtzhFSz5sI9NL9Q94dijBTBmUB7xi33HgSfYoDNmNvltd9XXX3cfCl0X
yxb6aCWcGDuiafsT3KhQZPs4AaD3CwAsD+pdAjJgiN6wbuqDKzjk+C9rRXklGiis
ymh9p63RZ3Mbx95nnBgppsKANLtfC4xoSdSLfS9P8DbgubsMZg4zY47ZfgOhsqZE
Nx318zXb0LO8DOiQ8he/s6IwFSRDXvQbcHxk+U4MX0yo6ibPDi5OiA4xNzIqZeCN
gYNAQMbpZLrpjCceSMrU6yKmsdngPFzawwpIlj/OrBf5tzL6SVhI9g4St7gX8ZnW
xggWykYTJAlkfAyVZNfur/VqCyYvazcr9UsEe6q+rH6HThJTqRE1QOWht0zNdR4t
ZFtVXr8G/uStbaJS239ZZC/Rlqk2MYlJ9UhtuQVz8ISRATKbrQHiWHwhHbRcNABa
1YAFkzhhx/voNmJa1OlsyhD4V097kJhuluLDG/vCXTQfXQ3QI0LqmpFRbhXN/6q1
JS0chrafQ6SdNS6emPlDCZ2YSgT8j+grYtMwSzQ0jjD+7j3wnqMQwajfVeV1D2Kt
AOvsiwRi5mLfIkKk8SFAUXaveZa2f7d5ZVGBQPKbe05OBX1Xb5r1GnIr7KUBQbKw
mlohtBmPPlg5qdgg02pGFEhgtbLCyzZEXeh6z1XYs1YtkWPh0eQlDkCri/74ldlA
51cMN4P5v3vgy+8aHaUk1gvgfqETNIGHdWhIR7pHea+bRBXRPRK939dPKDdYeBjH
lzEZfHpL775M80kmTno3qNPdyhTeHOdx0KkdzvtE6KUFqt45/e5qmvHeMw6vmHLK
SRp0AvSFrnGtGaLrnJt70Vc6P4wmPUVpr84dXHVgmOXWXip97m6qfpHIkyXwH/Vv
UmFXJi59/QcB+qErqFsLWkKRNzTqk2pjXT6021rr+vq810rqt5V2GEWFp/17cyg2
fpXzmkYVh7bLbMZIXgUOf0f1sY0lcUKBYxgpaFdE1sUgL6mxqv7rDSklvi893I1W
9KBGwUau7nguiX9doNC0m4gRHuieQ3TFFeeSw8JFv8j8+mPvqwFiXXHT9jv2uKLO
1VQ4+wsEC6kj1dZQjXc6icr7cbjQGTfIjKMKHruiv2PjHH+VZZViLUYyO7cAs+Yk
UByyP/zU/UQ9eGKhGEP7r0SAYDyxNaWFAKfIE4QWpzYay6AIEYvN1/cRXAqHRejn
YC8nBBz/M9HMLt6IVHhGBKLK7jNIUWfEwXpj6YNG4sDwpUXMVHTNXjdIXXP0g4xY
D2Wf3eZaI88CEztWq7EcgGVYxKNBT2D40eiIOjObYupsZeGUtKdtCPMI+bMzotSf
vsQ5hPbCWPBI3wg0TtJxr8x3UYLbePnskdeZ6fKKXoMNmg8V9aUlzQ7/rUXqS3A0
KSucaRunAZq/7twnisb19EiUE1zCQQF5v9jDjk/aCE84uM0sWhXzR0orIVcV2Gmw
JoK44iqi7bDowqCvLyfKba+Nzklf5udVWPr5LQUxWblRUECU0axE2TxnregDd5yd
ueNRy6EZWDxfZUsLrVlfUk8QZdq4cbAQxuO2cAjrGN/LAo2jp0oO20uQ7WEGm89b
xmfBSWjL7nccw74M20zrleflLC0hxaNVtPFqQP0WthpSbx1stoLdg6xWG46D1gIl
5LjF+VYQPKCajtCLStqPXkYStrVZGwZovYmZFVL6Bs+T/qtpgeEp4LIS90FPajbc
aSYozCih/iPpDVYb48BMBCEdshT7m8PJrA8dD7LTMqJsTEbbva89zOOYTo7yorGA
ekHcSsq6WDEO5PrQZEY36C7E0wtHgK0dsCRj81c7DDvouoZCSjGbxdNZ0T8A+dop
uD3qHy0H73oijDtN72qE5VwNxQ7AqW3D5pYc6Sd+95BvvN3Af0cZkW75zVi9I8Mt
ujZX71q0tEtkdURDQDXMS9niJIz8GMKL1pvrgDImhaF8kHDta58O38a2FHyuk16u
uU+VYF5aP9h2KKBy9G+it2fluZmXfGzWuxV6D87Xb2V4a5vFHcO5TMqG+ngfBVcK
vGvwxK1i6KRxhEfnlpULpWS5k1pHus0FgSnBIOrnNbhlyHpktmvZ0OtXc01cuJoO
2ezX0Qkv04NxpQGzwXB/qN+n9YZAlxLVz2p4C++pB6gmAJBDbnAmax1AXdVpdQXS
W9ncn1+y0/2umxJSiKXP9E/b9v16x2vYtTIVqzSjylpNKhN3mfgU7i9RrtqCM8I/
iin59ahghZ4l2rfECFCEzizW5tglnxSn3xuc8b/uGmHsOKp5xb6ULuM9wDJ4RI5g
p21YW9Vp4SMlDQZKpF8rsAn3uJ8gqYfWWBSMCgGrFlNGd/FZeIYgaXmG4dHXCbS0
XEq9V3/aQOahxZTUEY0bsn41NNfXoUQJ/z/CsyzSlQeUVKwjwBp71tHpEcwgHbmr
qY4ZDzGhnrz7tjFzn7DgrEhovWhjHUClDicEwJ+qi8C3Ja/Ok8bU2gmjJSwnMYnU
75BixHlcaSr95LuJfEB8RfSSVe2Sa8r3M+odTG01Icqg4rywQwVMJuGBpHTxfKK8
hG9PyoOJc6MzuPU06CSDUrR9nAXwPnP5WUgIQefWwZ5UosgZSGvOycAZ1pir7pSX
H25jzvMSnrUM0b2VmYqcDsseF8rhpT1zSBqb5cDRLN/9EMWwa3+k7DeqiXEues7S
KaFVk4NHl+AG74rLR3dFT0CdW6Hmd9PYazpYclaamtUQ7Yi1DNM4tXG1xmE8DAN5
GJUhhOX3t2Kn2bkRhW95yPwnn/+NBD7ZALdaZ/1XRzo8R+vwdIoEC8IgXQlFgS1N
MJTxoDXeRzViLvqgtWYYrGfWo/GRmu7dGGEqssxYfcrJzoPvAoVR+jFk4Po3ZETI
/4deA/zfYxedArHfqNi270VjgPRW7pGY6IMWE5vO1s7yO24xbmvpnk9d+mhRL1dn
dDLZ8hbFa3eMy27FQUfd9lUHiePLJLq+azJbxCuouLHTQDcEZQQDM+rJdr2gi4sP
tk61rb4BJj0Pr/n2WlQPUz6tZm0cfpbhZVHVslTPw9mlQmwb7b+5uiJrv1Q40or8
1X2ipFLCi/p5LxbHygMdA/48Vj1GcOMDY8kP+z0l4J0hDyhwvfTqh+jxULDML1gV
tf2C9PwayzbHQalM8ziaz6G2V+GwA+GilwPlgEj/etWsk22mXmVX0Z2mZwNUjTZ9
Sc+fXLxzpPNTFT0xRGnUAg4qXC0EJDjxP32klFYcNvFSa5C+FEtec4/MDV5Yfbk6
iUCeCTnFGe1a8517w0OjMLjMKPa4ehaOAz412xpJJsAdAJDM0S6WZthEOjd8xu0N
SLmNKoRnqSgt1nkQoGT3vHG8YGwP6RJ8XA8g25h7+8iKMZX0Bxc+CYoCOUgQbV2E
tnVqLIKbwO5RL9jzk08hzN7KikOypYLGBRuZnRPjvm1DaChwxYUSFk89a4Po7weS
O3Xw3psdhsBpWM1ePAInidRWRpoXrgnNSK01PDiwkwkob2TbCL6nke1/J6Z3gTB0
gQbth7oWcDb6daUOjRzAKXCuskJEH9NvHntNItAJMnTLMM7tUbbU/tTH2Wmm3OVR
tMzqPWHEXUGgJ2jwEF8pZ+Mbcj8xC42hvRBzi2uqsJmUjMGn/h++j0tz6BZoYxz9
Vdg/QDbrG2KrB/CYixX2g8kHMatIeVid4APou9HB7by+Gb8JCG9QI+xBJBGj5171
fl7uiWZd0BHNj+REblYRpuqtweLOg7yjQ7q8o7T+I1cqqUfZBrDFejIEQgUzJbsi
Ke+dz/BxDgzFAOP1f8rhNamfuqj+eyZSEGA2tt4FpyWxAbjRaAyKmMccpEfJX8WL
A/7UNt6SwXrgvc+LYEjgB1ywsgyi2KyYmpCP8GxKzFLtH5kaVSq6uDynJn14Wjbh
hSArkiLbfZvPh5i6ithVBuohwsxXtXAURNj0+ixYdZOWtqLcStNYskPu+A7Uuvcy
zeOFJvzZFbm6mIDlF2vxZ4TkdlvFS2/T/U/0dVPvcJw2yHG6wVeupKFZ6xUW5H8O
snj+9VaLfe7jfm9x9swNrEc1o6JAKvhDiWpYHRMSEmoOY6mFtp2HL0MASjSn0g7F
U7hJRKz5W1GpGAmV8JixIwuiLCQuqemxQUXjGdsGAPwyOg8qR++2Ffp19sSfpvvI
YNCdTHk8A4+RSjg83UkKY9M+q8uy6VxKNjvSATkaR8AEssqGgloABkuHhkPZWDVT
3MS69GGuPo/1xvBA3fVABIujGjw7fzdoFAuZ310keVZwGtCubK0GdGSUWRJ+YLGP
r3bpqUW4dHT5qZeE/53PWTT/LA4ZJ+XBb29ot7rm4UBHutm3OELJvRCJZ+0jVO3n
cRYCr1leOv1mLUtdWC65sR/IoEB6SVdriPvqF/ZBoe1LyDT2uMdXLVtkWm8BRUFj
4A1Nlq+soi7OjXaL6aCTs8FyZgZYTJXV3u7nCUD34ZHP9R3bff8FQY3sxOGwTMM7
dYyFFO0imcyTn4g2qVuo2rS0e6xZlcG9GwXQfpdb8I7KDIdXqrE7nvWaTYyLTs6I
Yar4yCCG2no0KeUXag85QOUzOqfpj9cOu6hjOAdxWXRJ8cXKQTTYyYk0HQoKL6oD
FqjG7eBc4CFOPYh4w6M+PZWxIuWG5jxjEbksHKAIdK64XFoseJ+3WblegssjBva/
xp7C30iLp6sFsrEpVuVBHQh0hh2VbNhiYeadgx5O6c4HtKcaRWJRJgkr1ztRTuVp
Z9I/YwXuDtFNSmL8D4N7IQ1JaFT1wbj73GUWpO/9SOLVVQRiISx8C2vLrYX3Zduk
sQKvWHo79YQfKsHrQhzWapdZPQPPs/M7MZ2mbUp0QiFVsNhEsBzYXwfvUwi5RP7O
e7RM7SURQaxNQGcGFlPV00KPBC1GvBPn8GNC+O5rKPuOhGWIwnQvwxz6etp6pjtV
WF8tx7n8eBrdq1PKpjb5Jz2txC10g02DVvfcXQs6E4hvA7O0clTYQbrp2/i2WU2G
M30OrYUiUpmYvN0i0RqskyMgVK4e2kCTWjX+lZ9e0UTsuaN1QUri+p5CXPbe1J+Z
oTb3GyMoCFpjH5P6+vlnxprCp0YVPfxd3BBGxmW/qn8u5dhLY1sj5nTGNZOJb42G
1nI6LjXJS5A+IY8QLQZZkxoZ0621GJCe0P8DQQPewPJLKAY8p43z6sGQ7NtjH6ec
NE/uLxqkQTugI4h6EQOFZM0vauR/FM+ApFId2Hgl81nbDYsJoAgeHw1deKc4xIve
5hcZCC9dv4qVrItSk4gpl4VSoJa3oyNIHW+sLi/crSd9xfmiIRYckRAcuHf0eY/X
zF8sA80n87IfSQoViKUtXkVYnMxjSLntDPSvmm6VffC54SMJIg4ruXkNNZGkOok9
Oee1D9dLa9o38FKl+bCBccyOg5c2SMAfM02BllqfoHKAGfVh5h1ycywQziFUpUMe
m7Bkc/y4JYbSNCXkblq+xG4io6nYIq/TAag3BQY6nESAHyLyR2YoWX5DXiPzvpvR
ELS5QgUqWxgrG3FGZk24bsPxm1JHofHTMVSt+wpx0qRfRhlwAAodpbCQwEQ/OpiZ
M7FNJMxL7InHmfQ8QX7arIIRQ+5fXQeUFMk23vvc26zpEKRWQajE6rd5PV2zU2rI
5hnMfTPa91eeE3TqYd216NngyJvxwMGILl1Trt+hOqmtduZdho8NShX/Laz2/+KB
guV9Dm/Q8u7UOjB5wjiGowxBWeRea1xjQ6Wv0JqLClEQiT+jYYkealST1arM0BGo
FkBS9flLCn7CPVr5X263OVxkyccVPFHoXuH9ukT+hPI2j8cOTGQ/efhxG0qJ9BkF
ayRvmBkQhxn4AEweuEWCL8mgyKoN78pOG0wSgGwEn75GASg1stDrOWnFSXZtDcWO
wJSIAUj/z+VNzh29Q2MTdtVRt6fWlE/Pa5agADSFFqkTJzbHOf2sV9wsfRgQP08X
o9jdoVUN3XBIl0q0yiccYOqlVaEuAPU0O4VhkqLCbCSyVb0TQfUAWBXnAxhv2bD3
25BBK23P/GHqmnrxB/3djYP6rq88HPuHh1Xw7DhoTH8knk5z0LutMC8se9579AsM
XbIsehYAV87fqayc8GMQH1aUVpWuzKkaZnQE0xZmxdjjhuVaMutgoaYOfxshoLzX
0JBaDXWP8qa6okLlfUZX0bxyWJH7/jQiwo7Qo5pBLUUqsAhCsejf8FBoRXPZF9VJ
/5PcldFyPb7F5MOiMU/vUxTcFdbrGBmPpKXoXMSalMNABzDVwZHTGPMPY8ga7aTG
i8cIpw4TVYXl1xcsN9IlsIRD45f4h6FIlEqsWx+EjHHXdQnfnoguAnIug/oT0Lw8
wn4c3OV5pgRIp7kADffRN3sovLuBs7FJxs8PR+Mq02O6UEd05o1NJEAtu/BVXPLB
o/KFpkj+zunWJH3V2Af9h8TA8AeMXZOeDvtE0V5S3GGkF5jfGmH4ZMDOHt8MrxZv
EtYOyZCNdeG0fIAD5Q7kOjHbMPWcmDRmc7OSzgvmwPO/qMow/v48k/Du49VmNkOO
sk1s9TEhD2vrFgZ2eZl76arp7V19KhEz7ZaK+ieUn5B9MN8IAKvyxWIy+wjH3Dt2
H/plboxp8lkQWy5diOaBDcpf18p3d2ABiFQwfTGbiwstyHfqOoFQubrCN5V0XtZR
RM71/Tk+OMfBsXoZyrnZCnge8L8OFJCELOwpdtFukivPbR1m0u0N/vkiYmGfpuMh
CLFdgbKaUjFI0f9/WgeDfgGOctAgJZMq6dszn9A4kHK1koH0iqV0J40PWaBsWHWj
y5Ti8KH9BFYZ/gOeOy4cGGEmjigWbdt9PkJGlBcpMLPqBmvGh7UA0l3f3dEx7TVL
Q2n7hE9rObqea45tJteXqa3YZX5Wd3BICzCCTZfd9nWG83AEz5Rzv+Y0scledGqs
DcDh93UKq0kztYoTrCKN3OdhiOZVSHLTgPIpKVu/Wf1DA8rNVs35rAezetOx8Pxk
3XF8f6PQzpy/CNJWAeiPPoEnovXTHGX/OYNVpsLeQGzqIeJpwRkzdXOa04NYBQ++
SFHbEASaVmvLwE5bcnCaT9HBqJZfvk2yHzJsVn35rkmjDn9DRuM8gWBmEgKJXg9O
lPHG/bKT7dOuYgUH4EJ4wPRZeI8FuK5tvuFd/C/R2ffUQCF2adqDAH+3JaAXiB2Q
cWPBS7JcoYXQijQk9oAE2rIdjhf6Oh1Ge3UfL/A89YmFPkvS6lCHmuC1A3w+9SYa
qsQMi1AQf7JT/gBOAYUTuCtdpoeLpKBkRWXVniYofyZJ/66x/kW3PXAysZWKxxsI
UZgKGDY+8ZSgNGD7xixPkvGM6GWS96psxHUKw5eFxUwXXdvtyndlf4gUR6cbv/5i
wVIjxD6/QU/BX//9q71PiqK+li+JTCaCKHY6mPmamD+G6u15mXx6PK6HjYnV2pUo
Tjuj0nHFbx8SJURaiyh7cxtom/aIvEhUYNsga4xO6Yvk72iDvDR4F+FvANv2hUtx
CoGM6t0SvJLjsEGX52zgpx3vSi8rrb6TjKMIgZEdrmfdBEnh46pfQhkORF9Ox5N8
wTaUPk4+bK8MFIvD0DBZVZIcNMGR6VdNif/CbaMf3DeNhlGar2q56lHAs2wi+UnY
/jSJQPtkcB8aGuOh5kcE5fREmH1PBLIukQT12DGwWLDbtkU5PnXOeFgvHApOmiwD
RdRBA5l3xI+xFAgsmRASov0PnBNZ4MLqKXMWWur4e42bqKtn1S/eBoh6OEv08jfD
DoXFJigIBBAEtr2VwZ+aUZqwFe3Bm/hTIuceMM6pumGVwzd+kKkzIrrMeF3WF57A
1u8/He02xjUKYJA0I1pTKTHqcE5yBeAN5UO1mKhhkXyOIY0js0HGpEpdErPm1BsD
HsnPLm9chXHmLybddCoAx05YhcqIA2kBoq7ABKYjkWCJid3VebTerxzxLvoCCW8M
RSvc8icyEW+EOcrCCw1Qc+3TRNsI9EPnn7q8U3xlmLV0cmAyHi/m/MKUxY6VIAO7
/116cMSIECj4o3uGWmEHY93rweE7+iDujp+4CFWKQfks1hojAkorodpnK674bLA4
ureQJ3IP6thmIwqpntnKtvYGZh6H8SRUq8aTIUqEy3JqVqPADqoQZVA7hvZkRQgm
H/J3raYqzBVlead4Or5DEnL3vUeV9mmSi7y9qEuJaPSBdCkvDyfMjQG9LtTS+fBW
VpiGH7BzOvNlKXur1HuXSz8A/Vhp391x7Hct2QTVvKgDpBTBU7QRDz5p/u1h4Jkz
fhnCACmG7z7o6bGdscG6akjXSZo2ty4fyEzPT2UvwDtRG2zSCWulJmYSo3EIjUye
S7nOdbbea22GGFaHcbty4AjflW3Yoy1zHOdlzHbW/ayInnLH7u23v//VCdhqDsF9
B4Tb3hzcsOW9VNwql0nhKLamvSedK79MyDxwj+qlk6/F1LI9nQ+jf2L1LGp/Rdz5
GlFOfaIavzi1qr/5mfAGRIllFyWfFBHzjIU7rsA8EBVNfQBzj1zp+DdeSuSYGiOv
o3vOt77HC6AZujjjj1NlgVvOS4gewz1qonPINpHBz+hPFppzubiITmJX9cAiMg/I
xdxx70eUhqNfo5Z3WRuVZ9lwaUSB+Jz4YEIiKdFtVb0ZWzWUpGkhhVJsmYAvaA2f
DBCRKr2YzDhf3mMKiO07aWtgsyPJ4zvoH++Dk+Vo0FXe/E20bMkkdmBj909E/4QR
lbuqO5ukEZ2/fvPjfXG6f4/CwIsFh/AKdxMjjTeB+Q1RAQPcj5+oVGK4RhCxYAQQ
PZ7zORqFgp9uiSMXJ3Zem04agKrHu98TdtoLX6wTY2bAC09kL+9KeckuD7J2dpbJ
Qwf+UDm2gKo47P97JLfnergPTTFGyGXOzPzYCrF9zzkA0vhPAvkDnkE42OnwxVW/
QYi1kf45dIs2i9UOeO3HjO8asZGWWyHDF5s3pjYdbiPVX+i0cERR24rIDW2ysaEh
6ONjPq34lE0EZvNw31bKEh3B+myJq0p9cCy4nYco65xXOl4QK7P4Y+qebfcnhVfP
47HnfNj6pT5CHwwl2tKZz9bvYG+DiROpop0DKRIopft/rP65syxfArse+hnpi3kv
i4syBlUUJQSFBkQckv9U9S/+jyjirG2iPIoilzxtgPO7ELg/ZZ2E/5CV482fGRnJ
2N9xqL6057pGjX4acUJAQ2I+2sxM75b7TCgtGGmaHHEqZSgVKlNTNqfPemTZrfMq
QDhD4oZ9aba3id2gr4TWGoI2roQUlHyCIv2fxjSKumIPDcR1O60lQEaaRvvNBVNB
VnJQusEhZ7/Lv7UeaqBFfXFT7Yk7eo8DY3bZbP+6h9MbUz11BIYuUBqlTQOsv75g
xFvkFU1pe4IZBwXoV1epR2gF6zs8H1gts0NHSpC8J6tNqbaIDWzwETqFGyX3cVo/
HyXDdYlAaV6ZGnYNW8xPM/0JkvZ+mcMzwoN/SCQnDc87RUms5oVvMA4ZbMOC6Hfp
3JQf8xxcq1wHtz7U4TrBQaaYTFzT+hGMt+v0mwbw3jefIDpVdOUS+9uAxXOe9+ws
b8Iy9i8Ny+8oqWv52zl9THWT4QKdvL3cAMnx+JhEMV5/zTrshQ9SJoZSKajyyeAy
Wl7l8UTo2tKm0L6h/bMtDbELGZiXed5RWkt1eDtIj1F5CPFDFjH257XXoFjksrUu
6S9S0aw9MJcWSz+sOf3DUq2+qRzeQ1Jk4u0CWhr5WxT4N1MiEsO5TxjCVyBjGTXU
Mim/7wMvjw8P+zX9L+VJ9HZBK9sVFLEM4xF0LeTkgmI07qsptRI9vtnoK1sViE1i
09+fmSAXRsJdC/VXli83OfZmhfr2ktpVeXKJ39FCnpRRKPzUSU9W65S4A+ZK9/K7
rKkyOO2sFLz496oMeB7k+85X9KBTJEavomRkGdV2EQH5xKWhjGXRIjwMj+7pJ/KU
CxUj24tvzcmYjqJbtCEpoPYP04pJ4kvp5ZMhsJGswQx1ksprzjjsje3IpnAbpaXp
NqC/90RWCk4bzobk1GDlq/I+290rYoXFsFyL8InzIUN5Behrai1/T2hjroaQ2cwU
9dOX5tBQ2cyvv1BrwIuFpmbPUaClHlmaeQ9Js1bq2LASClA+nEe2+RHIeasXdxlh
ayp3qa+0lffIqErcpFR/dTYDnYytG+WNsS276uECKqOVYbP+qa2Y3rk8KlNOLQiL
BJm9yoyT/EF5epZgbi5nL7QGArHQVnCD5BoSB94qjEcr3bqt/Mg/vyeiIOgCXMMj
QO0paR3k2SyFTFRCyRW9YLumLDyk10HhJvZmZlFNiraow8s8FZ0WJjxIZXuFQnzZ
VYRYTJIC2w8z7cBWLyWo5PMvTQ/n5Xdt9t0073PPnyT7vj+jiFGDiGSPySG6XDY9
1mtyAIqqnlxdY47uoA/yhC+Vo0suZhwrxK/oxM5GGcgjvLVuseP92POmkqx8HmeA
JtwTMwJaA1nbGhp/BCpPLlTFpVXES7FnytukbFfV4keVA4g4QnO0/p/ycn3x61Zq
y5i/urHAFSd1xhPvpA7cLhC4EK485Vv6P9A4lBqnE4ci13DHQ+Ug2IDFmuxCtkVM
0lXjcb3Sru8FbpNpbEkpOQLDWg0JRsFAAGhYbQxWBRBw+MS9UQBbcS0w2mczcMcs
VbdZGyvZnikkF9F3d0GlQ6PINM7bCqiITyAEAHV8HqsIRodMheNb1SYV+jU0KAsU
LpC5QZ5WzAjnEwFl8Vl7lxwaPiItbi+ZBCOq790Str1qFMtAfm12lzi2JsRc2qbx
R460S3FzgUivNx5gNcHtpwJTI3OjlJ0P9flNhlilPz1hmhtGLMZZlORYWxZrSsGa
7k7nreM5Q7l4i6cyX/kHoY7SNyrfmJQZmNM7+9VkBWaewvhXmlGjgw/DJQvnaavH
k1sGHKalbPEam8T2//KKuBIXWHclg7GWYvij3ppM0s2g+2w7LgxsVhOtyfryfKYR
srtg47P25Gpis1dqMvPEFldcBAUaAmKgH9zswQxIeV8+d1kGmKlBHZut6tzBIgTb
hryeOEqkbBJBxIn7CsMny0rWUPfyhSz4oP9X68BucQ5bifVFuxL9FFQm+HMY9zbL
DWiEknRV6pbBHT71dEV02COSGWRj2x4J+soCWwWEaOfHD0JXkOZPx1l1VJTvn4F8
RSHlrWL6XAt/iAk14tISRhtf7+8EZLqvOs5uptHiydcOfUDYHxd26Wopeu9CUlRu
hhF17Oisbyi2Tan8Oc3DjAzSwwAFm7Ya/T4g+RIHxxSMXdh11ZIA1D/wUSpnKWjR
PImTuH6EM0EYmKfrkMkLgP1KWqNdBZmlMMO5uLHE4w11jv+g+jHoTpg78FRFOjvH
ire27cJm0KXw4Z8ShEWOHYj9QH4gwK+z6rRhZMqHqsl9IJII2MiuQT5Eqk8RtXZG
h3HznUZj79aXT6VhB2WjJj6BVtUJNzx4FYNqqQl9ZyK22ab3J4F3HBZq64h7paaR
YT60ut2guqh5qeqgcx2xdFYcLTQtJ6k69sHY1EB9hk15MrXrZZkxedBnPEjoQz8f
kApuu/NfeF2a0KPHa7/hWQComRDuoOzooT9ux1Qi7C8PbJZzDzBdOHN4b0b9jz20
SB64Fbqrx/P6hiGysop2TJiHo/RLBZDbPPCPMSMuAaHil03HuCOY9dmUyENokYMJ
xHPcrZMzAQemekhbBOtR57UI5yVrqst0xYljmUxpLKD3gBqrzXw7Q23mN5mAF79y
RFWqbaW9OhnNAXIEmjZwX/N5IfFRi3AgkIqUeF4WLI7RErRJS8fgkOt/XhRJyUpq
vRadqQ2om7SDgFhXBqhSqLrecYOcra+C6Zq9A6R64wZDsghfla5dLBRApEzloNiG
TdsaQVd2SjByGB1pC+C3dEbqdfbdfJp+hu9uebW8VRhDCtLcBmsmlUTBbIT+eiNG
1UfFMAM36+TWJjzJvZKT3WXWUeTFkmlBDfvkkePt/eVEzEUjta0MMgn9xiulAvMN
t7iSI4oIs5uQ31j5o0QwVBT1eZUZMWJAGxVbjwjluuvG7DHQuy6g2YyYKDoHQcGJ
ZMVJpUDY/IFTENwON0ZxBG0UZ5E724f+vnVAXEHobfc++krwijH7WlG8C1XwwSb0
1FgcRDrmUnrWguKIe1zJ1++LJy01t7+YkNXMHk7pBH4KXxSQmltHWNTQUB01Mit9
TK6GCLZrf2RjGGy7xcNI/IG934kcoh6svoVfkjussRPWPMnuM/QP2OxBo5UYszq+
kklVfYDh5zD4p3h5Wp6maVvRBHQQHlnUSnV+HPaGNW4zFWhNPwXM2qJvSOQJN3jS
k66G1i8uUdlbZJtDMiQLcfrjMue8hKCZw+/+cO7LTRSdWdRXlgMSxMwSNJ61dGB9
zsDcQwWyO9Exnz0Y4qyqXweM2AWjpjTEU22LBcFmSEXtWrzzmvJvNoSRmLS9kV7L
8QBxRjfKzMzjE3wizV0NT8lzAt96jV7vfn0KU4vT+PrTm/pMZ+cKZqu83gb0JNBp
kDnPy49T4u98zTDREFppD5lL2btAaKKN4rqycjb0t5wcANSw2+rqth/+KdemMxmT
/ZWlbds1EhyNCiTKeLHTmBpo0VTAJmdYndlFXvvefDGhYrHjUdKhfY7APbwG5leV
gtKTAD21szCmqg+woMZDBdXJE0DpTxd2yH/HFzDIWGHHKlBaZW5uMipyVqXHvTeB
H5kiqmhBfJXkJDvDjamJtdGGGE0Bfs7k6JAqnodrOuEhryt9pzcEzwB9W+aEXi0A
0ObXN5xT0h2F7mPL+Xtc/TiNKjf4myqn5o27e/YehFTn16vOj3k33bEPOL+ELJEv
i1RPvb9xsYJrQ+IxiWXZANFbiwadXxKeo3dHLpAi0YgpQ2AovCVWYw6IorFG2Y//
0ZZjyKyDz2D7BP8SaO/fEnpT66hKXrmGvxRY1Uj2OZ+wjz+3xElwM/HMrK/4UJ3d
2drAvGj7IQBywiolwybiXh1Lnph2sSV9XaAqzAteNE5K1IasLTD4fVRT36RRwnsZ
s2r4IoFVvGkm4Ty0A35w39zoAjk19P9nxFLFNF/iQpMM68ipAQdbfdGRsdmqkMxL
eDTbvQGs3eybnVYB34Qo+tKMyDx8HMjoKLNtWRG3oA0Kr58kdyl5f+Y0sIzi+Le5
7OB2bUPoOCgvYTROT3Q+Cqrx42hwaQ3Mhtd5S2Wq8UZQIpaCOQPM98k+TSQSazMP
5h62W9/0u5LGzOSHRryW65Zfj1d67hBOtiflHVnSVQAMaWk4xPwrv5U/lBJpopaF
ea9wjiNqEBfos9XAopgCwLvF+8VkfkeV0GBOe2IzPaFhLvkfay8qM6zm6ipL9237
pWu2CdPUaNoRvheyVSRL7cxmujO/pNZ4FFYDTlflHjWDYCLsVF7sqxXY5OWCEgAS
hae165QH1wkLWoJ1bau9ez7b1OJ7DtjQAV51Pf597gJtQ41gEFOPuPesNvJBysva
mtK4qwsd5Uob1P76kbNWwSJ6vFfQX/HUA0TL+8UcQ5XPEteFPBMmkhzie3eZ7C+R
C4/NnFLlToNy3zMhTX+IxuYLxgOVGwDbIRw/z0bzzB+dKvg3lVrpMx2yTywEuVK2
XD7ZOBXc/9wJsGRwGFvk25B4IjPgHHh/HAaHVVD6KRSXXR3eqBYa66W94mDbCOhw
vgI1Jy9eimKxxJ8EIc0wDaCuDflcP9YrOgjGG8wdfdQyXMInSI/ndMb+WgTSAXri
iqhwsB3LErw97laDcaMSjTKj1GZ7SWUlO87jKL+vGrC1ufLniw9roBVzTzWnZl7K
Fpn3xpWnWXrFBjT2FgJvOiDrO7PijnSUOwahhyAhSmZp0U1s38yiDLcbnR7ohkHe
jGBUboliyvOJy6PsK/CBIdswWwDI64I+WSoXSjculyRNjJDqoXoUBoX/PwYTzKKm
u4rJKQ5OW9TOkPlz4cnd+vEtnfHPyDUVRK/vM3Hrbqy0sT5zqzlv75UIAIp7T8t7
FuSUr4wZJdQjDI5jLsQIXZGqWn5bI3ItocSexej6cJZ7RY8CVfWoEKWe31dMamhu
3wwA4RX94FaYpbVt0F2+dQIiix+HiOBjZdpy/laRqLsvtfYpVbHi7tk42wA2xAPs
WYLN/mhMjwiniM8ZorZ+9icNVvswbbz3RFC8wJpHt8oUUR76H4uVm65P//EC+bLu
mlkFqj4exaGjqDzrhcmUqsexYvSoRFsTvNGVBhVymBtSEWiP0UTI26wHL6wQ9uV2
Ky2fA/ryBHbGA0XBB5tuemS+gOect+/DDLciNZV/VhY78AI73A77hG/lVuLEpu4G
UbJcabfUzZ6nDA8XTmAH+UScZwRlBJv/m7Ng4F/ApUJhUEV3h6gBHFIbsMyy7i4a
WY+1LF3mlIwxg7pk66RJTqEQ0ojlfenVgOKF5Hs7I4FcQmvFpDWA0TdlDkwH+Hfb
L603uUBB7bbyLD5eB7+7Kw1eFYJp23Pf/LDrxLxZ7fRuig3M6OFCuc6lNbcbgizf
VeSnOTIODyAt6abphNpIn0Sqs8Y0qG2VHKtbNswC/5DrFW7PoFsrWtWwbpiuaibX
50qleB8Dn19TEotolNHa6Tcd7PAnVuzobs2LyMJRiUkkmQIpdqtLg6ctGcrYn5t8
wgvkqjxSsGl2pcmmu+A2aeHYs6li9cigJo7ENXyt5KA4u1/uhVAX/YjMSSs/HPA4
qRuaSq5tfAJm1kQJkPVqXnCUQCKKUkFEWML81mUPIG2xVgi1CdY7/EFZBiN0SMTh
ZoqH8HPzcBhSn/nouP0/jekFxVYcD4FUkK5L190eSEz80koA6g4eHFWV+R6V8ant
uvLT2wMw3kq8kFDdkpB1FMv7OzAIN0GKLYwEuRTAcEe3/mXPQPZCHj+2WHTi8e1+
KQVKfHTQ5uzyoZXwb1aBNytBtH6Dp3lKKpCg2HJa94Espa4HzFAd9qjPWnGH+Q1y
uNIDKjd6lVEAHkXVQKJqWIxgX/hkESMh1hi1BLThRqfMM8qRhS7iiqec9ucxw+7O
tpRrySOOBWtQkZ34efp+UaufLOMhykA4Mmp26mDWnpgBusFUu/Xa3fzTnHxGACA5
N81gpl8+1z+h4+USCi/NJREr1N3kkmjKZZNOTvT5J+1F9tpI5Zmv12AriRWupRnf
loQ7dGSLn8xxAWefdxg4Q9hXVQ0bybldLCNit964HHgd7RaBSSGInTuKXWhYw5C+
l+4O3e3DHWHcIoBIFqAWBGsvL2JRPCGQHJD9rNQhFLPmIUqXAAfCzVjWfHa4+lw1
B1We+C5dHtdwpyBN8VeTKH6rCY0WuftlbDx8iLTze4ty34kdVPWKR3CreErx2Gk7
SPJy7KWIp6ilrJth95mhuzHcs5ezbiyD9BNc0yn2R9nlzltuWFwvYXY4pIGQPsad
yPh3smXrNThnxE7leVig9U16OI72t/ErnfvR0xQxwKvhXHB2w2821N/6E/Gi7aSX
oO1bEOnxlRaGBRgbG0jEekJemDrJ2YkgBWxZBMDQiI4l3gOqoBXCCJZ+xAMGqY47
hBx2gTshsJrqQQqMALxjWrcrVROrm/RQsJoLbt4gLMvmu/uMtDBfaYYTyJ2d5o5w
6GxhbwYPUKK8dXB2FJAg6f+360mhSFcPoPZ2kEwTcle8UF5+RXdfzl3vyzq/XeJh
7cykFeJnZ8WWxtzJfOU8PJx+RFo152hswOWeDlsOkC9tEWJ097+TbcCqz/oPsyDe
6qQ3j6lalHdg3STmxXtk9KElFQCelrY1P5FYFv/L9d7zpYVJk+A+9Rc4fn427Gbn
+QcEytI+FqkN18EcD89SjlcbDv89cSF/IRrWJ4Y2MDdANkdwRKMJZw1YbjFb+Yem
dID6AMjfHRO3PGl6yhYmzsKE7o6rgxLUholQBQmqafJpSMg9cwNf2YRmwGBXVVL+
g3+ZjyeO9Fq+yD8969l08xoosp6rScN0NwQmoVXM8LqDW7Gmcwn40iHBhrsRHOhA
mrifxrnFSWFLZlfcfQGEm+N37ZUgH7LnQmasLrcZy2uNnWAt5wI/7+8Czq9Qj2/B
Xlf988xngjpuZB5MAUmNoofWJHODdv+cvZ/nXN0W4ndRNJ68ykjQcYpYHalxmgAs
+O5geZbXb17K9Y80jbfX2kjxfxJ8QSJLuBHxPQdicbjvLRFdknWPFRm/ZGeWMvzr
escuZmNHSTyV2Hmui6b41gKOxzl+0TF1ipjNXGE0LEh4yfuIqkUrPgQUief2sNtO
1tD/88MLYPLjWq9F+FzumRr/MbPu54Up07tSYBXAT3kfFiVWSv65I8wGx60bSSQc
tBSIOo0e55p5NLUB3jCdJTfqYtNZ6IhJcinFmdazmmp/jabA7GOfZpAwSmPIbeUI
Tm6x7JxzJARJhWZE1sE/30JxMPtHuGOwO+B0gatSQExP7ivqQq5RU9E9m+NNMyeG
kgTFsC6zaNPvxc08PSdLGqY7teThQQHcoB7j2WdNfBbvPuF46JINbTDHssQoIO2G
DR3f6WubEu/lSdY+oPdJAnWG6uiCziGPG12jBylJslK0BXFssDFKIEMwed8Xhvq2
f9Mv8jPTg+jy4Ig4Q1WUitvikV15tOUtquGabBs1CRnglZbvVOYaJXVIWIQnFPFB
/egT/Nq2hvE9y1zskWVzfmp2USTRYnfLIUrIyJGfGtMRUAotuWpv+AQJl2oMEBtr
6PcM4idgCu7+IQnRCXRQAxA17Ec1gk40qhlLsLFYwsPi9Rv04VHAFjYWTDkyL8jb
NtnksszkWnzVtKT7O/2C7Yn1xxDvfVJjA8VnQfglbZprl9E50p5r9lbpPgCw1mkt
MqTPPqVTMAu5ZY6mVsdjIy4EO4G0r8/cr2ynjy/bJjJo9E8Bytvv81i3WESXih9w
gjfllXP28V7rfZBUDPz7XSC5/Yd9lRLAb/G0UUtwkodQIOGnMuYuIxYKxzjP8Axg
W2HkDsSQUCc/Abp8vbT/E/sKDVxyNWHVKusQHqKJo+rimM38aQEfQTIVIBLbgVmv
IvPEMZz/ZVsQWe9I2XV3363zS3mD1tgY/Lcckbx57dBukDpwCF1urtcL0Q77at7c
ZJVOIFOxMbFfLbuDJlasVffR7bSUJsWxvQbasP3ph3ow9ycbzo/HCZs7Rqj/c8OC
qqfONvRzXeO0xj7+6gP3YlnXs/7c7Mo3em8cGwzY3Rl/Es92KIIyeEwHyHGDcjVh
mPd7KxUM2LVFvQRYSjWUZ9Lf755MxlQLj4ZW9LqciFBtkONv5S9kukCfVPSawGzp
YysNT33t3IMD9WC3ScKRdqo2sAzAnXuAviubA8J0hD24rbOMDdlDsZDff95jmQgc
+m6ATrQ4o/SI8aBfVAU3FBvSL337QYoPXF9A/gbTIYA2H6jzKcUaRCOiHEj/ic53
+I0VNO1SPrsZg7IfzVe8UyHlgwUf7T+ZnaOzSp7LxmhVMBnLzKBYqVmP9D/dRS2S
8zaqh3CL00oKVy/VC5QY3uiHtbeWU5Ls0uQK9uqdTxGhUr5BC7Hqzh0C9w/CjYnN
WZmB2i+4lq4Yvr4aZLMz1KPkPSiVQtRMbcuFbB4+GV3B8K6RAh5/OcsYGLd3sNUc
2ofNtq8/F8UkPf2MjlQAXb0b1bPcL9Y3Ev/dWEmQ1/XKp5wx99kmed+QXCovKInn
tLFnKh78tcD51gmIX/0xj7ds7YwMfYVwJBiGZ6vHVO3VAsmV7jbJZ2ikmHyesY7o
TTJ3WO3lyztnOoSr7hQNHj0E/hqe6uS9/HiXO5EyPzrah00rVs9blUIxKy2T9Elh
xWpdcczH7k8WvPCMbrUcsFNLaJWCouUYIoiq3OA1r5c/cKy/8qHSOk1121mrrANL
04NYfmJQYm17J0VPbfij8JJnn/KqqkcKQ7w6xNMGA9vcxyOmCvJJGznAQo8Eicvn
iNClbpRQmWy/77UEQclxO7V5KldlCJif2CDv5/eKevaiJPuE1UP8XCTYEdlQ7/Q9
UPf7EChFe2LBKZEhiueJLOWfpAhl1AWeb6kQNyVZrVDLEJhFWNfi9UYf+sfwUbtf
Bje9AwL+HyXZN6c/1yiElON7CYvYDDExB+gByliYu9qiJR3vmEwlpAyD/xdtdYYc
3opqkY8cN+MAvFqFao4gTEbsbzbOvYqyw1e0MSuwE3/t/8XrFULifzZcTnfoV5n0
gcCxWYpdZUdJF5HpmlkT/NYpz0XUK5KfPWyTG3HaY7mxMs4Pc+rPONNeC8DXEwVF
aD8lX5cNCQFcLfbUY/Jm53e5iwh/0S1Rj2no8j9wQPuslHVMepnss/8bvwli9Ohi
pk/GdMaXWX9YkLGKnogDcZg9GmSUnmIIt8nU0CrynbBn/v/Zh9DQ1r9nqw7uatA7
Vx0DJp/80s1nIOl/BJ9HrHngLNnti/lZAJsIuPGXLF+eQMxRzLqw6nhhdxeLivNc
igYREh8vMJl96LNFZftJLDwSZBwH7E1eqx3SVxzo0s46/aecPPIy+JnjoCLqkrYq
tfx2xlg0jv5tmnh9PGXj3BYVwaKGFshBxJpPGqOk3zugaq+d1oUnUwSfCM6fCDYe
bzIcVUmyZX0mwt/K+hzjWoFcKQg2OKRKCcin2ZqOnLMrxrL4M9TFNmRMuzmVpd9m
o2Ib7gJeZN/cuH0jzY1kOSfJgBv64Dbu9P9czY/OFaiXNFh6YeTUyMXItITipapF
XqyBzfCrvgi4r5yey0+QFg47Gr0oM44vtCQy8iqjnMRSr7TiJdj2nYeV1mh06EA7
7cGbduCpiPmeiD11HBCxP3gAe1LmmLoijf0RHt1XKjRfJpVJWvF78UMvVn8V5S6Y
ipq/pP0mX/KJdOgkn2KNaQiSCQf+pbH3EtF2vg7XoQz7QnS93xHTbVQH2jomAmJ/
Ay09JqiZZ/kkcUp2dDoGOeuUqiz1HklX/1XRYeIJVNwxo5Tn0LDQxZOgeLT02THG
tQCCDT9wtDIygsrIeofC6zcjD1YpvT15D1rHmNYSBbJ0JGncJe8xVovbM60BonM+
/5HNxkh5jaIW5LwkzCwWP3oorbrezDsJGpnVmTPAeSdBFE7OF3aukr0kaPp48DYq
I0dKJWK2s2WsqmCLsqDotBoEZziIoMD3h6813rZwzag0KrqklnIgEvHrYSFkx7Ql
mepXA7qK6E8Z1OrkjwwSTtr5Tm2b45wn6NJgjp8ftrJi+e0vaYLBxpx9F4HoybF3
qhwgc51fyTxSGeLMjE3o+ZTaFQbMZtuRm4mlkyRPXHDpGUS/YhnJV/oU/nsyvX2J
77x9567cXti01r2lzoR2zHlW0N/hWJeqswrhEfxlKYagxbqBiIBYSkudnO+1ikPm
6ZP0zEn4ieJe4YXpLGg4q+4tZqmlORzHJPcMMmSB+B+x1Dj8G+mvGsvtxWICHZXK
XYtwcD3k4WebbYxTCIPpALR1B1+RJl418VqmJm4zCkzyPusSc8gtUnNy9/5D8UDB
/0MKrN4af9cSR/XnRY8UgzLswMww90hiZimwmsWPUi3aH8bSH4pC2He1hN/H+ue3
j19xLCV2dlWetalPa49FWoFvplQHf+81DLuQEL+3ABvDE66lWBB9ipqTOZ1tPmNv
PaKEZu+xyD3KC+Yy6QuaJn6mSuCaQqLsPBMfdKvP9FreA3a+/WExBJRujXvhcFFT
YXw6u8JQ4EHelyK2USAibojB+tUvlMtKnfP44H2i4fyC9hyBaBGUgx06wypQWhq8
aM+Pcxjt/eE/fLXXzjCenR7jOp9nTUIZtLx2WzGqKu4WPKxNOPCAzR79Q1STshDt
onxQVOaVa3Bemve7MoestyIMGuHXNo11+xcAzLgEX/pgriC0mXo/8n79EHDXjGSd
OMfo4KqTRKejXeTTZthtn+SS246UOcAk6VO7BIhMXP/hP+ooRFS6aSHGUEttqK/B
2nm7aF7m8pjtZ4DBOPqpcrBVa7LYbBL1sevKeRQmGqEzX+35BgUlQ+8b6fHqXoPB
BbVqwW7bmw13DwlEiaq0OBA2tUl8GsdwqzBVLRWtxy2Kccrh/f+GuIpluJT+PUw4
T5/POUnEBTY9bM7C7FTV+A9Vos+TYna4B9CVdA0jy4xA+mKJNBvS2uQZ9s8bsv6S
soQlBoIeNZ2d7dBqJ9lcG0qv5CX51y6C2Ukzk8exYZBDMQ1XnV5w2v/yiFDa2zM4
g9FMMqupdSmlY7VBzpeu5Ir+EVTxnHehU9lBreNl2v2ERuBg0j5sUF78aKHIYf/A
sFJCrdgPdfH/FWu5G6qSEcMjHcidbA1e/Sg//CjB+c97iSCXks6EvrMTWZf/N4Db
8IJakzauA9SQtAdXY7TNx8ShF52bbtHaMMGc9TvYQly2h86UFrozbPMX38OlfaVH
+Z+VvHaOQ1wSqirMby67jTFKUMhLbgM48Iwb47G81Ef2pek2pFHSZhuF+9syEF+/
38UwdSuDsUgCrB1vqqsxbhWQ4oUXLmzNtwTZPAqDdDH/XcsJI6R5oNaFUqBdXMMc
hlKunzQ01iBX05f1bVbXBZLIrqkZ8uuZa13iMyVCsYUNCqViqF487l7r8BAJbO0Y
dxqpO2UsX4U/Ft2GWmN+At7t1fXO2+iPm+CnSCJzgqz3iOam08BfDu7UhOy6H284
dBfT4xLiOGWqDjrZXiye/ovxd8QEBl8K04gEQW+M3crng3N/1XmXzz5GVGG4xdaO
vpLkyV/iitRVv2vNnL6n5y0K1DUKKHHUiTKYiSMmgW1/S/hKnJCdOTBvRRL42YX3
XW9wWtKPDQJyzX40CAaBpb8exYIetcZjNUVpMYvxh1SrFDP6Bm6b+g6ShxBvq0oy
rFnpGzje9mCY9msbgI/NGj2clxVF5+QTP1Mkl6rGgttJBxiF5QHZ0djp7WtWtq5M
8BQP0Lwk8L7U5M+vXcIYzTJNJa7SHrRjuTyFIFo4TS41cExv0c+CQpRkSHBTqsR6
YZSgC/nPXZKo/6fCPFWGR0a8sjKTVBZf/lZR86I+Se9rcfXBJJ4pG4ffIqEHJsH6
7EV/SRKd5UPp/131runhkYKjTx9jKj9b2IhJXzkz/a5TZ0zr9RnMEGHVEWDLVjo8
SGYIptAOw14E4dvMNUXKFEGnb3TwOBoI2xRTBTEGFkfkgNaVrs5jii8A0C03QqtT
6nEmdY4CpRNKlVma4BDO1Jsw6PcZLELj4hj6wQpvHdharcq5dAogRg+8Xcbt+QyJ
EZ2JNTLEc0Or+AmUWgjNKCZHLQkWA8wOpG+SNQouliL1RSLH6yY4QvUdFfZt1Rzl
Z52qE3QxDoK8MHjqMu2sCitZvS9fwcMxzfRANCuJo38pZLo5KvOZco1/a7NYyERJ
ivOqNruRWGrWuRABjr7OiP9YOoq7p3Xeg3FCWe6CMGepDDpZLsKrze0dzc+oowiV
k/l/PO0KgdaxlnKZnJ7jy203xIzj+kJB2ZdAlPm6SMQRXw2bjRMWyaTsMTnD6KLg
XL4t7KFREGBUxv9WY0JQNL/h35tSYPfKr1E9X5K2MbsBi3Ox8bBH+QGl8Gwn97mA
ovxIkiNFceF9TxPi0n3ddPh76BNlwWiZAXTJeXwMehUXXC7zG6O0kQb0tAaLt8i9
daKa6K+zfMYiFhnLna71B2vw8MLHc8il9zKvhRmmjTqp/11ST3MyjFgxMhcN0wIm
VRQjorlSEsYVoLsGrxRjcYONu+rvxVHmliNbP1OUOVeebpiBjAfabvh06IIAmLZ4
VOME2Ev87cjxTgDyikFitT6KGikeRf2599fskVj9v4CxuRWX0SWRbMhJ66yirUhJ
s09DJ3cCqIQCNiZHaLsLwRMm8j+qsbcF7fq/bMqoBlV8y0dOPvTwr3T7AwifZjaZ
Kb02k8d/N5ux0ZCuImdAeMMOkAZJM2qjrsqfqkx2yq+0VgGiDdAQrNvsjL4MCMqm
XNpIEyBmw0lfDbiBDEW7sHaxh2BXpQL2MdnqhWHfm/XzDZGkpOwylEty+Bj1E9VD
nwLP4qBOCRHVF32yDv5T/m19odLQ7+GAMgWFSPyv6Vq7i23+e+Q4DmzCbzBS8gZ2
IsAKhilGw8rVhRsobduR9RpB/ydHIQnY1QFsdQANX4ghVFJMTlaBh/ZybXinmez6
7sHYYjRjiMTtlk0T9YeL2wrcR6CwF9ifI+Q8aaZxRzTHHkuwVeG/6NHVusqqTg1y
UoqXUgPYxAscnzbS3mA1cLCPiXxWI2v3ImQT+OMt8E3/pGb/l4Xv5Rj9HnWmwzCg
0zCQTatwiDroIJZeYYSORsyvpwwkEG9pVSx+GBbdE0fGv8R3eJRG9JPYK9ADXn+o
2EqeeIoen4dlGcLDhsEAdyUQ54/uh71ynxu/PQTrEr3BybzPSgucef6/DgFQt2Rw
SnjM8xA5K3XOVl0LTW8jXWg2GQkVjvDyt1EKKrX7u9sJtgF+t2Uiv6FDJ5V8KWhe
y14u5ikVOjfbqDTF5vF8Wqxre5kjJiahiQywzKjHzaS/YOka62Kk/rs1MUTj7LfT
VvikOK3NuJgVxhnRjRS1fbLZx/A5odmWDQ6nqIoJFvvhACPGfWF5i93TXnHTPMs+
c9bblKHurKGlCROalUKEAc3Qx7l61AOc7xihoskS8OqFKT5Lw/+PnKLbFZhRUaKT
+q3C/H2zi20sOGz7rvnQRjDsz2bmja+66YDptBspM4ubv3aEK4pmW3cS1Cv80Lb3
Dhqx/Vudln/zXdWjKoDgkn1Njoe37KEFx9tke67/6je49ZCkLBHAHP2ac/L5N8lL
impEWoZHNiHfmR5UITpM1nYnEg0aWeZUd1rI5smHswVzoePU8hod5eHeUPz169mM
dTVVNr5mfWiQyp3iJAlk+X9YnnsE1a/3DAA1tG5ui0+foVCedPG3lfU5aMY6Sfm+
JjhnedULzFmPoMkPECpqIbSX64c9PuO4CGiyZR0hWhVMEZMD+/CdfUulmBP+g1jk
JjUoBgXSrSg4agTgRQcY0XPhn8Tg9jLLOn8AUOzZf7OyJ4zgMcoPmT8FjZJcpfYt
dAVEPZk6rcOl6MzAnsYeRDBFqj0qB5AdZTZAYM09Nu2nv97adEb5WvzYyMtWqzTb
HGcoYq5vzaZTZO1PpUUk57G5Ae5RXBdVLhveW0nANfIWTP3zmd5wl/6Gll8f1zUJ
/+7UIUviuBebmixtqEfm2KYCaJis6S2mzWVC218Tt0cQrb85lBvrmFCAFxQqPbBB
SwBONSQvIuVG5nn3ln/xZCM6fs+7EVU2AYKMCdTdWsP5wNeXR+O9QlMNni+Y7np0
/oWLm7nedEGn89DXrNxnD3H0jZIPrhtA6rQw2x5Jwh7WXSA3N9o2thZGm7TOH+Xk
aB9zE+BeuYAkh5PgqigKsj4vQUFIWNjOoAyzKJUBgrdvj/xTZW5SQ/GBtNTtTgGS
z0S92KnjVcEymjDW+iH9eABwxwR66+qA9krCpDNzi5/YoX7ttQbkdK+ID2OHUP6B
M2jiRWTm2mVVjTJ5b8c/jqAA4A1RqFR6OvZI+0zysqB66z+xB4irGLSuBWFuPpaK
SoPp3ssamxpEAohvwd4G9vEUQeUff02X354td/b+7GkDGbs0ZOQipyy2mg6gO9ZW
Jk8WMsCNZwZiRno7rm7qEsmwJ+uPdeEAU4m+ohIwKpzgrlHhWGowg0BCVaemtv7E
s7nbTunq957AATzQkDKNIIfyrulDxW1+/8sKDsGfCpl0xW1+j+5kPPE6O/jRbNBo
wf2eDs+NCP9rIQkvHoTmLjS4eMU0Nde+v5IJOohcruqmUdkjEYjrqm8i8rN1b2su
UPm3at8bwO9mC41c9JKCNB4EeShvk9TwHxTwlVqpfb5IyM/SvOd7qC5dt7veiJ2j
BVktahP7mRqPzqFw/bEFUxDZiSaynRg1xw8ZLBVNXRuP8X/0jJueSqYutLLh1o93
Ss+9SoZKmA6Oy4e+z3T1UnvsqE6mcXvBwrv6IiiprdiHeQ9rm9ay/p5yWofUDhSu
lAcIy6n3/mk3QHYDhJ9cEeVwjH5EZqbXPvA6tAuSbyABhjjufiRHhMFtoYaAUo+z
DqKzWnluJAYRwUTZz8uZboSEwzC8o8uva6nTaZS2XTnVaGgwDdQ3lfgubnKfbt3E
uDdGs46wXQmo9LGYDrDOEKeXpPqvcFhAYSkhumAOIY6kV4jdSrERKt+Uj8Za28y9
cq18gc98ZCn3rrFg8AuyTByR+X5qaxNlZ5hUAzr/LX/4OFTVUc+OrIvHDyjANUCn
7PZOpY4G2pJoCfJ/0kxERFwOGB/Tz+lneQTmSCcZA3c2Ee9ECfURWRa58nTdEaQ6
me00vUP5yFWzlJ7yDCuy6iJRqdjCo4gI36GYNg2PeFJvUEdarwJU/7MWYqEHGuSz
XSdi4d//UKGTQfhZyHM0eF4U9quQhO0gfm/WjStBMCkFqdJ0XTu82VzP2LCMRkUr
bE26ntiR1qMrHkw6BH2LUArNmp1GKxRyyCqAwizRNwg6r5U2tuqlEUiqT2L534u0
5XUX+seQjcXUo3gTHgRtzLtTSnnNjHmyu18UTNlewrLYBaSkfUvMeQx5qk145gNB
Lt/xpL16m0JHsTBm31sx6OYPhYWJec4OpLhfpJzOqWfV/9fEPvxauXaKgE2pWxS/
0DZP8AYYcztmKmbT/jyYJW6jGwZCo8kwyT2G4tnhwnGovvy0wekz1LZ6AqWDWCn6
Ua3dePnysd+ALrL5komDO08+VEwI5aLUzUDf+tQkbiTmZY/D7KozCU9rgSqUiK3u
ZMgbuBSJmUqVczNG7qCJNcW3ez+h3Gewz/LPzEmCh6TFig6C8ZQrccS/Njuoe8Le
C3ohRn2urBJaeNP9SYivgXPBNR7UArXU/bovX1viibDikg9Pw/V1/ypTRW6GO2Wu
Qi9vlKijNCDBEUSB4rPdqwjh6Bz8V7lc3+7KJkfN9pmKLl0kMCiS0v8JhJFc0+/4
8fDrsQsiWqGufngKzLNpNaKdSK2zKlX2gbANO5Bvj+n9OdfBYde+OXg8Ym0OuYHU
azwQS9rujphxPp9cJAOWlsWnGUxhCUZ4XQ+x5tsahohsbCXePyjlONaUh0UFOPdj
5+2ZlhNYeLeVq0VQoyEvQfa+l7Tpou7SerGVyUPSidVu0/ASNIKzqBZ3dF7U5GBm
JNn1nWuA7AeMdyXQRhmBrsYNf3fEqPzFPxU14nyrL92rr0MS+qN05+eI1YP99YBY
7vCOuHEwyTWPCREFk+Lg9sWs7vDmoUNh9C1XZ9p3dnyJUx5Y0oqibQc4pOhJiN6F
hRYlxuXiq6/EUyPlIZKSwSX/8GWTjfg3TizF2nM2T07333OCTWRCLsWDhEdZa4+5
o3x4RcXQL5GFUH65imhEEVRc1PY7w4VZNsdJfYvVDmZLt/y8HcB7zttLtSONqB5Y
glaqmReKnco4GWUbffd6lCrdRf9sSuLncDj/qfJo2952DCdN31fNu24wKsG5sjrN
AXVaojF+KhLXF1Mwp8lyjq5vR9e1CirjF+10GKyDsDWm5MTkwb0zo7a2rO6ZxTKL
NIESB59BgPS0PeEftC/bw/obMbE0947qylqsz5QSlOjzbCM61N327U3pkOQLa2Di
cwcaoVJfIjkS4K7hIAMn6JlWZBRpNUSNFYzGExaKwEZd206ZXeV+8SkPyn+/9abl
Uw1ZYWvO8G1SeaMk7tszmOrGDr8T+IIEamI4TwDn57VsSV8HgqiV+03Kr2+Qz7tz
1DKr7y4gm/DArVMVfZMN+V2hIkD85e9zZsXsxS2NOTxtL4028p0UFJwx42OK61Yl
cfGu/uJzQEMAzA11NbcX8fySvgvewca0o0G3WEptqc40lMvvEDXtq95DxMA/Ougi
j8+/POqcJO/GVCNp3cYkUjzRXIluDJCP3wige8wtj+w8IP1zITBWWGqopTemg9/o
HPrziX9GqAj95G6IGLS91n+KOK+Plo9NOJBZgNDcvIkeA2QRjELbKtUvxQ9h0l63
X8JrgcOE9hGmAF6hEdDkCVdEyu7i1xWg130vHp9DIY1Ed+KDFXSQ2gKS4FWHez8F
GQL1ULg+2qomqBSctUwlR5ExzW8RsI8IMVy7rwL2oI+TJnw/e58ur/p2/JPnhXoK
+uMGLOE/4OrpTgcGFUonpTQgu75a6SxBBOWZ9SFO9rmCgVQBXYmYcETiqqaOX715
J5wx9TTs8esv0TqKWPhFh52va8WflW9WfDnCMHnzJf58RE2c4wgruqxNX4cjSRQ+
b6n6uvDHeW6olY8mIxBwX8kZpgFR4oRzNJJLCeWnC2TFyxvR1D2HNcBfYTKMT5lK
oRHvJWOQNuqYcmWAM4GcwpQvnpFJt+za6grVqoTgxqzGb9+iHODHiMPVocoLcb2r
QJRpYbbFFa/UqYM4TdYijRSqapjwZJKw8nTfA1RkBjLyGN6c7Ulr6Gjcdcs8Lrpp
wF9Es5qJJDSyYjoXy4syjJbTrqmAv7cQE7zS3ehsB2DtRGYjZ4BQYguDJ6OlJVgv
QkSOjlj4mGb8qCh44MMkBve/2RFCfqSf20ucQysemD5+Ugm4UqNa0PreB7zH/LtC
zfu03psKpEX3wKTz5/uWuqc6nNqNTcctu0UCD/ybsY22ep2u2CJIAHTZgE1zEAVA
KXHwMegJenInLbUMQPFVQfj8jzhGHlA3QS3LzW86DfMdm43yC0SB4iZFlj5oflBP
`protect END_PROTECTED
