`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KIiLogTK91auS0saxRjygkExFyFK1y/cF5DbmsGyvTwbR4UHb+Y8xTzAFeG+ITn/
1sJF4eCpbY+mT0XTaCK3y0uRjShIF5gB0M0Q0XVJzPwMsQ1PCMt7GahRK9IhcPRv
MxfBFzDYIfHdOoL3H9sCTZBpn6pITViBRB0i6exRPIrFFr7V42lxSpKkbeZEvgea
P0Cyk9LKucYzJPCOOIWN3nxpp9tXChFDWGt97XocvHrdEd7o9mkM4WdWfEWhIoqH
d/wXBUklm1ejvyLmBis4GJKQEIjcIjW/E+gmzh63vVeGOtFLkt0UT3yBbUpu291V
59/75RJPnjRnm9H1x9axqk8JmVBSRN/R2gpNfd8KdhfguUvLOmJAS9epHcIWPR6i
qsq62h5E7LZ7hDK0AmIQZLDCapHhTehEDkd/wIYinTakFV6rlDXt1GhR8UpOXjJB
c+E1ycC3HN5KCrEWg/A22H4lsvJi11bmVkR0qQJAOI7pv8wtDtnGzanqDeGpboNh
1WxsuuQyTB6iReywcOWvZJBqzySj3eSqQKNiCp/Kv/atqy/NfHkPzYkUZNgUvKE4
MJ9P6aGihugYxY3kSevLt4A3AkubdhJVPOCdjIKJAJCWXh7o/uxyvsNratNiWLY/
l0oxkbxjB9tmnQJQq5G6kqTuVe3LLTK0p31A5hmgaD3p/g1U/sWnC4odLWUIL4Kb
ZHZKPbjVi8wyer0Tmn8JTITLZsesd0Quk4rEKdoMk1rHUUzdllVmImuKf/r2eAUg
1ly8GzscqZG8Xb5d3VOQxsQwjS5Gm3I+3E8xlKZyFPs+mC3+ssh9qQ3PqJMn+m1z
UULqW5305PIvf/Gp7Dt1PBT/hi2A+Ilug+bpui2YMkOTCr9+ZFCyyZJYtxM4bS/j
YrYnF8eV0r7gobMYe893pJQJuiny1AQjcaiQNoj9RW5pl5ia4LVF+LJ/HBparQ2b
p8Q78caKhtnxoE0rReHwDGhaRhn1Sm0E/HSoqPZHoAIbYmRDG8UUZocIuglTSfea
0kHjepy90N2V1O+jUs1n2lsZFB3zK2bGF0y+1qtWVpHhPVU36FG9AP5jTkO2nYaD
nYtTgq7OA+WxbmbwmovQzJothbOPsf64nAYI3UEsbdZy7HFf4jnd4vtrIDhjRVzb
ukXkLKCfblmuBdwpRCkOnlnNNuhMPYBHZdgeBUhTo2vuHXlzFNBU/bCM8ebCyWpc
9dnyy1+2uTVW9KraPCNod6oPo5UuNmpdLYoNnqO1EGepLSe/Ly2r2C1UGqrN7wrT
5ybdJ9C3wBCGJUoiAVkbG1zs7K1VvF/+ZL4XiMT/DlUMrjK8RN3BrJ5ukAoF23pO
ffdz0dbHi4lwiMVP0yILmJgIb8Y6FNckEH4yJ695UF+P2C1YfrKBBDJUNnNwpGVq
jAV6cgu7w7nEkDNmB6j7fKqbINQrQS5zesZMfegqmjB9JK9e/0SnGyyLq3UmCzEb
wVUcu8tLqkYhF+RP3SbCEb3Emy/PCKYPWEJiA940G9YjyWtC7RxDM2b7BQEBeh5b
VkI68IuTYV8DAfEuDLeZUNl3HA+6HQm2IhwTMc62wK9euDZb3cDs2+oc7It0gC3/
zMhKHfHH+c2+4z54UuJASfkwWji4c85qmT8oV90CLBX8fZa3tlpgJ+n8kzJLTeR4
mbxQMAAA/n7GGAhiEpXGYyf4OyzfQUWQpYzWx4+Kn9z8zF6s7a5iyUwnxbde1PJp
IMkEFN/IqPc/nzWdhyLBvSbn6nYsN62oHeyax7eKdZ/JmBEQ26HM7DFTsnDIqaqc
X4doQIQfQsccycIfgF46YcDz2ZDnq98t5vUADKiDxR0BoGywcGx1e9L9wY3zT1JO
aIlWnY7z6WabyEJ6gsF5pBSldCQ+a6wRxlBPOD5Oi9GHgpPhswy41DiIb+57yW0c
0pLKE1y/MFaRWKSNo4ziBnBgvyFLCOYhO+qqnJYzJofOZ2po3WYEF+P92E4qZeFO
vsZ7dYOOjd4ebUaFBgdrebMvJcAGpgkpSyB9af1KP/H448+U5dBQSYatGUAKfTZ/
iGywjQW/OeKjDo1TmXp17G+uagSj9irIpX0pdSsDAuuCFNc4CCd4Kfwu9BlRzVGV
kiiGKflhPMfcr0GCYCg+H8SJ8cyXjsfS38SOXjlkKgax+6o1y328fQZN1m9MMWW8
KtIHOp9SPpudkdg9uZoQRp49PxPDyt0Kpt5/TX8wg88+TFnf/Vc//vWnTDqni7x7
1jWNw+LIGfWYpx9ZYCt4kw==
`protect END_PROTECTED
