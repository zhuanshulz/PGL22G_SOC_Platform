`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yU2FRkE+NR0YhJBEwmcbgaNFIin2YNjic87++GlZOg0kzXslJ3vM4MVS+/Dpwp4c
AdiMM6tvfN2cN7uhEDyb8d4bd8IWUZCAR+2oSHtA1I4rIO5Mhy/1e9BUba2GXHbJ
qYoiXJS1n//jrdCYtSGmp4eeGvgQS70p7oxzGu2OXXkLNXpnzrqBhB5XkVbvMODn
wQatZ/h22zqT/bDG5jL3F1LS+sZBWynbLK+A5twT4h5fEHTPGGiZHGUOVj1NkTxD
7YM48jwEp0LviN2HVyuhEHTgGX0z0N5ts9Zg1SC+SARJW8KDMOG69z0u7cp1iGDK
LxXZzKTcRd+f3yRSrL4Icm/HC4JXGP2DSj3dP88gjjecuRxqwb9LcdsZYovJymH5
wr4kDfe4QuZwU+ELWEtr86eBCksaE4aapg9/2zV4mxeeTlQB04mQE37qVCtH3sU8
1aHA/+jWyIWTmDwgbMWfCdI/tiFh5izGYggkFut2bbSJYJo2Y632iAopahf9J/r8
ODB0L8GfR1XP4GMmKoPg4xeOuuvfXANVhmnNm6QHVyd7zsps4Vdu0ahP3mY+irnE
UuOk5qs9twkp4oi0JRSDlJde5IBK47ZRSZ5CtoVgJXm3gED49Ou2UoNq1Briiyzp
Zd3vtnCKyJ1m0YgFMS3U67K4iGBhfXtyP982KyBBWfsGIkhvJwsPQ2VHUEVHZfnu
j7RXwVgAUaL1m0Yy/MGzPJ0CrLwSHWrw3dUE5tQtfYH6yIMH+XgOqAz/P24+YYQm
uFWI0/e6/P8vY17fpMi5p8vR9c24E6DJ1k3/KI9VXzQFpGMpkDhxQtUdMfuUr4Y4
uJPO4XANZI/rwcCQ1sZz+50u+nS0s2NEWU3dLKnMYa9NtuyWxfMrWBpRJH2p02nT
kNpUqIL2CmpdyvzPfhfSX8K2h5aJYfZbsPh6vH4KQ0czpVULwROCeGI0uaHCV14/
luLOcySrQsni3/bDM836a+hWQx/qUTQ0UnGcfA6AbwOvEa6BpBS/zDRxOIICUAsV
0WXLL5b3V/VqvRvg3o48j98At0DIdRbbp2UnWzoIGHOGznjXzrVf0U7Dv20TjlnK
sx5EpxSuwe2lbnJs3JekOIO7W/NavQc9+BGzgtG1IvPDWD4Klm47GoLxAz3xe62f
Wv321aIfXgIyW980gKY7A2EncsS+2NNNhSnWKT39SzgNpcNmmTa2+SuALeF4moIH
qEHT9ZmTr5r6v8eqjSGw7xt6XdubwdFunMfqOXwPfHtVhOLKaUOmV4HfjP2esICp
mG3YEyJt/B7OtEQrjWC0m8N7Bj1GBkER5534WbsqRJLkkEQeeoIoFJicXwEvpXZZ
2fKZ2PBxsgn4DJwMTmOg5Lx+PvDawzPVibdJoxZGYcFvRXP2AfWGhtFrvq3j40NS
pya0qStUgHmVQLuVHjWH9ODL6a4tlQn8IyslVn+YW5DPMtTdRyPZ6nlY3aK0+kme
IW7jaJr5dxKAXaUx5BWP3+RUSTF9fxYbnjncBbuspcRSPB44Ky8Lx/A8lqc07+Hr
IzpqHOMPrwYdWgFk6nI43kl85WQ1Fy6/FVA6cQKdqpaNDO3MZhTYfrFqEw4ycSsK
rTTBmJZ5GrOWo35WLM4uRT1zO70QgO/PSEmviWuwiEEDTtKd7Qsi1X8dlv5jfkoN
gUE42SSJmbk1YsSMYgmX+H+Zjt+5ESb04VxWa3kmhVoTyf3y5cJA0e76qz7h9fvP
w3ORTtc75TVXWR8B54Pu7gFtoTNdoKE9XES7USWcTfS4DA6bFYFgUprmlFuaJxIX
6BdupGwGTpPxXEGPS+cX7O/Fd8EtJ0yPbteUO7y4yWr10iupL4XgktCpZA9Sp+tx
wZN07vOLaSFt2tP9MbJIRWuY0PmYDWOMvIK99p2jP/+V7C9Ou40LS9W5Y5a/TpdB
j6Ho8pMINdGWqY18cyR5FHnaYv6LKO6uLZw4P+WsD9cqSEypZ7NQpYN8Xvtrd6zP
ZfZmFaoiMAsL5F4jTefK2VaFKzVDOovZwdLtW0bYYgjZiuw0rbeyyiQGHv+nMIzD
SVGGfG3sIMqr0KpYe4zOynSxX241Wh2Xh2qvwT/CoVPjYtoJjLoceClQHvmZNtva
r4CqdFdic9G8whJBugABceU7+cyt/rb4/R0XWDYQ0wD6Yd8p+mphMpva2NnVs3vb
8qfDvrcn1K+/IhciPZqdKDSdcYG+kChhofu8KW74GZnbzhGm4Xwy51V4ZMvfYw4j
6AoMqbNIfkbjHwOI5jG1OGVoKk6k+xoeQRLzxGKaRjT1TQk6iTyflLyinDtUaoMQ
NAI8SzrRpiynJTyrFpcIKTNW6BT3yCI5CcoYCX8drxN4Wj5CE0PtkJXmhVyw5SQx
c3OFFFk14bXCYTmXtH1Qg/PQdkYRWmS28DUy9Oxk2sqvY0cZ/O++9oF3ERR7hGw8
V6dly/cevxZvd1EADSyIfxGPC9Vj6iJvHgzcI4Jn/U0txi1JjSmThOQJqiYV8FTO
iRx0G7KYssmDSOA+b/AXsuGQNlUPmk6eDV7yjIxpeByIKg2Ky908mBM1v2+UHCCs
H/aff5LcDJONK6zLdW6jSNeJI5hGwuI7gaInFO050Ql43XaxhKUKX/m3ra8H3+yQ
/BREwMCG6NkEeK9voTgQQFm8/dAdKJDZt4Ptqrn34bvI6h6m6qwErGIellbmlxI+
ebQ/y33l5x49nJHde0PdemJGpGgFpPilqKaC8E/GBU1Wu7YpESW94Df81UgJDqem
sRuhvhw71Kak2bTLeqvDRBg0zqyPtDZl1/z0uRbu/cYBcWa4Zp2ftQ83vM4mM+e1
yjSb6Wb+cWen9Fgd3ysTm+erlY5CirgLqbFCfRgoVvOPFXwpTCGjKR78UDQAktRS
XlxJikLXdt/fAxgOetc1qUkrnGgq6NxxdrKCQxWhJKdQMm9S4Uuzve4QJwl0q278
z8fRK1f5ZAfAyuiJkUn7pNFGiCtXDGYKq/2q/ZnnjmvkD3LmKJYUBhrZLZwDp9dW
ymMruagR0nv1t453TCyxTKdsSt8M4HDszpt59hj3jRoUUmp+HEjhEXGfyzCNbg5G
ndbEM20wSCzEgO1XCMAjW5edEcFDmitkbe0CzBGbjDDqDE6+/Mipx91NjtubzAFC
e7sK+JSxuy1ydBXBzbZO9qLapJ/L6t9z5/BuKCD2f7+HQ+mMvScrY+qZWle+Ehpw
Zx4l7fqEqm07P4fQnEioogO+bl7Cn7rDMLryWU5RlfssRpmhwlbOGJ3E239XuxLq
s9OF7CfXpv3couHa1Lf6VxJFiVx8MgmY1ywMXh0iOvvyHe8BYK7teD17rzvjr2wv
SPqFadQ3Wz4UyKBVs86+4bB4sIOeLpZlAcDGMLPDK6agdJ0Zy3ESKozud2RcJE9K
p+s12urCTuJet2kqQ/vn3pwQVyeounp6lZoQ5Y4adaS+palQ+wC8GFTP+gHwoXoz
N8LZtE8Vrx9AQI9aMqdCR+amHPz4KGw2AhnZwnmjICXwzrTbEN+5XhHMQFAOAbt7
44o63KMEqCZ1fQPbDNm8e2ul01nZUn2sAXf0qETroLAfsiPpFnB8i1VuQwnly4vw
CJ+tBnPEFJH8E0uaklsrEqRrfb81itIx4Q87ljmgvBoXU4qpE+33F/jPyzsoL/1Z
+QT3F0infPvvIxNneaQZ0bQAAk9p8E5DL0TE3Av/JZTRG0xpo19z3s/5rUM9dpnf
azpCtklnQtY1fAeAxYRigDovFQk/IhP7vIGylDlsS1B8+qn5vdZXkxA8RKY0FeZV
lV7o1UYX/iZoomkAUU3CqsOwr/GqWEv2ZLDiVQ09Ba7PsBeB/r1jaKDxbef67DGA
4gNhy9yq6ayogk1GFnYmyni6iHpYVAX12+0O1ZIfUsnP0tWxsZrl54rnYRflfmsD
XklimHkRZWKZlNfpTivsyDdfFzsFXdbjCp+Of+QteS1uRxX9XpuvURMlTmvmm5vZ
t4CgamhBo6MGe7kBB4XTrQhuj+CjZn1kME3fdBYczX04ap9utStQaRa8n/SAfcVL
ZPvoNEhX8we+23jghl5XJUKjUoQDRvVPZIcgCyI8ap6pIBn+Jp2wwOGgTFYCQa9/
0X9rPxRS8t6ReFhOC3Z2Vl71JpWV4qCDAocIdzekYmPCmMsEZ41u9+Y0mQQSkCv/
38YXuGN3boWfsXYI10jSFBvD6HDS/NW6v67LZZ/cRmd5HzjRJUbQNCTPwhqJaiUT
URo189dmCJnukSqmRbdN49jIAoLGZ+14uek2zWaGyPirclWE5Pkv6+uyM9y/eOMj
If+QYgpfIdEKSQWl53/Azb3d2JYzA0pflQpvnuVJLlrsSGDnVNKfsJOdNSOUMQ8p
mVby8wSyP78LTLCtNN1Bz7l9aRdP5sYqU67VpmgCoG5e3x1aoIVqgawPeyLH9w58
oN6YJIsBODrecvZYQM3A5o3gsKwH27QvaO78FZuwWCNAyqt13fkpJ2rbX8ZetbwP
JIxu7ATKsygrmhtzcXm295EnCBZLi/tK3jEZt/h5BxUP+hr7Az42f+lk7tp9eZR8
xdgDXGU4K5e5jk1OT5JVmqZp+m/CQcM5olyRVyfajArX7QDYSQbP9VgMnjLyQouq
u4ghyV0vgGC0TQCmtRb1eq4Xnk7P7hQaFTAoq92ci/8mykapPm97zgRiXhi9kTka
Ubp8SlxEYfcq6xF9MaZ23hzbJeusAAd9jiRESmywG8e3yPUaVBoOwMDWtHnHjSiL
OvNRNxE77dWWbv8DL8XgQPqYqBlb6eQ/ExSS/l2aadSGkvlTAhu+61fjq3lwnYAU
iv+jnmc4CMXafM5oI6Tpfn5cK60LHifuhWjfNmyTzFTggTEju1XHwPpAh28hzDPM
Xasy4dgjoksyhPAQC4XHTffjRnkDoan6TszIFIm9grjEGcpU3AnN8lP7nVYZVeYa
1YwyfsADdr+X5Uf25PW7o7wFHIZe6wK96IJnPHMhfE7L1RMmpMkUcVHA7xkBOqrn
sC2vGnr6Abu/LBP73al9Nhckrg1Yt2VzaapjW7DofS3HTnRVwGqCb0fXQ0ladWs6
4jPZevyqN8ViAK1TyCPCQNftGLgdVre7Xj0jmk+7dOkvUl93xMsE0xTrLri2FVBx
I8iXwmRluiJV/axMgW1sq4CgUNonoMz+FvmnwrNVCvDwatPM5kTFLwrI9fe8ad8Y
G/uM88+tUS44tjtbJTY+ksp6B4DZs7hIFOyrFwVMaRnVv6Tgiwom9/eK0Nfo1LHn
aWy1Q8Dlp/t7uPp4IfLEx73e+tCECYoB+aN75nT/lNwrxhGn8aeZiWGIuraf5ai6
/jjBVzNdwOaGxtf3OhAOPxMgb7D+poY23eGtZ1bEsnxGAI4sjDC6PvUtuCsC+ubA
77rGyb4rOr/aRUS3BgwgXD6SUrzT3OtlVALf3Ezzj2d1bM/nHKhxGIYw3HaACcDT
sTSxOLmAegWqPZEzCFuxRGObZDIWMhFz/OPxbgyuWXSyTA+wtzL51uYOiI+cMp2z
8jhHfrQ5OFx4Nj188KvCy8VAwg0wUhxosbA70+eUydE7OAEIQAve14L5GTM/r4oD
WZPzxyMLftyC2ag+vRqxo1y4AXH7EA9zc5r9ye5wgrOll5pUVhz2aa3Fet1dDJ5r
7e7HDWRpUuM0RbA3X303xbgDswqGTvGAlLeu+mhckmuKXG9YO8MJO5uDNigtFZSb
Q3VrKF84j3YQbn+g5DDnGNDeeTqEGChxwGRkWdntzBFyXNp0YNs3BfEAbcgECPm5
nkQc22yAtbqtKa4VUuOh6P9sfP0U1jCA+7Ev77t0EuKWermEJd2DTZ8kWQSU3ITz
0NoWQNkrJG8ErgEmA+EEvW1uDBfx1oLyHWqjFQt6Rjs3Oo7xA0cer3zFXaalRfDa
5p3Sy2+XRd044XxpKuWnL1c7VYBwscW5LaoQXkN5r6BSEpLBAsDPwiXoVSMSWUNR
7oPU2bzJ0L0l/0PNDUB38b5NpPAmGuIIfOA/6UGqwKd34gmoclpUhh6MgVVqLuhr
eCeBNrUZEwXEdIouUQbpQuTUg758+D+yAGt//w6vzkbIhV9/+xO6TqcKiB3EGOrK
FZdYMVefltaNOpDo0hvQwPsMJouXIcuMou88HOX+vjOFQkVqA/twQNihWtPAMOvP
t5NiW07jeLqMHW/PAYucvQRHK7pZL/UkmNQ9KhZJLgBBPA1kmDhljQhX7pkE8L+v
NMsmCEEdQwUNQsSA9vHiEKLEgn624m6kpeTWXEPTejB38gjhznb1sDQJcNl8m+oE
CVaylFZE/aepM9zM/3MqmkYoet18M0UjoCaerWUcSmCGQD7AkWWOhB2jFssByjpl
1a7zH3KckC4quOc+RHdM3YmuFabcp7Iz7cjF0cPyi39Q6X6CAwK20k+6BQfO5jBa
nwc+nIFOxq/YHmY6SP/3eI/Fa2yhwluHBZ5VjSNzkF9HFl7t10twcUWzjfIZwEeS
++PLRlPZYs6+amRC2a4E4WHy2nr3faQdApictBODWGQwphXW7ke0q/bu6EYxGqYw
QBrdNJA3hNOlQGlezQa22lVnyKLdgLNNpgtMePq5UxWc6OEJa/8YUfQ3afZj3qv3
20du0wRIGWp6mUPH87XUCGkLkT8KbWGdQWgdBWAxbkuAsyY4J+imIv6EJPVodiRN
6JVKWWmW7cPQqa4ziAd1GlMWumyTdqA4iMaBmCFxGn1yofGw0JeKv+h2bWA33Mj1
WTjKc0E7xTOWvPR4ZwQZVw==
`protect END_PROTECTED
