`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Y1rHAQrVRjATekpXYjDNo3PLX/GQeyaUCqjd4vPBo3xAOC4wpxSKQMBDOUmgNL/
EI18Tl5ahA8pRQk5FjmMua58THO0vLtABj6+GK8dtRxGvEp4zDvbjWf+ZmFnUijG
nhfNDPHenN1nJr15BHjdzPfuh238iXvk9rYubUTIkvQWC3IrFlX45i/ZXGAmmKO6
J/uXUFM3HirrEGkj42PeUSPrPCK31TTDuiAFS8F27+3/peJd+8jOI6/+zvH8FDP0
JIixw0kRBTr8UWB4AMNIzslYtpIQjTSOJE+B67snb7yzO16/gmTC4olOj7zrP86B
kQjpmHdIqwTjgsPUlxZTH597viwgmA+zq55+irbADXYs706nAPy4F0JBauGp1cUK
AeTDvx+/RDK5DCI0Sg8+CAMBn22LrezGEYTBmruCMfriTO2o+sONTZp37XQ2IZj6
PIKmk4j0Ec2T+1wKna/V5kT9CIxULBjgZw+9CEKpODpjfNKUKqz6ABRf+8eRXGOe
/gPMyxJaCu8wH6ZvcOaX/EP9+N1InbdKLFUBkug6rlSOYv1Vyynpayx5Rj/Zr24O
sxn1lXIX7IfPNNatCFEBWFIk2NrgDFE5vqUBBZpS4N8YetlAo9Ntxb7wH9qeYyr8
/Nz1EdC246zNJqIGu5c5wZi7vpsbFXkrsjFe/ymIl9jbxLHCY5rXHMl6cJJRwyLk
0eFcUJkKhpVCxy7YjTPS0NTnXnePmnjXXXmFmCJcGWzRNYblIVLv65ZPVqqDNVBw
FdFHLfKGaoAfjRS4T1rs8SfPGnKionKIKw+Wawx1opyNc8wRAuYu95iDFiv+1VPs
3TAHQCAjtJYtgKWNH/YTQEYSqgDfFXxqx8mrwquORWoR6q/fRHqzi3mWTYyFxcV3
EjkHxdBdA/spWgk87dDL1pYxo/QKjbS6xm/f/j/hjD22ZJyEH2ZVvF0rK8bJUys4
BquOxIpW5V5MftN/LHt0wjRXFUgZe5uwDydrReE2GtDpEVYO9VfXSfHqFvxG4jpH
oSpA4pjP9Ah6sQH/zaxxNryJUhINVH6lMiCilaZa6bFyYf0MDHSOrXrunY9uEc9l
vdSQz9kn60n+mKCgYu2pFkuuf5h7FwoSVYghrJdHFj5qidanHC0AKKFWf3BUzWEG
0gr3D7QLWD1qkaQ4y8TmKwDkVsuCzxN25PQUWT08bVKIypcavIdFZlgDSW1jG437
T2b4RfwGnYUtsdaGJvofBPsbovgWV3xAhZeX/QJ24hGy4zXXwe+B6rjzPHPYJuR6
QLTly4owP7cA/hthIFf6pWGyViVagwqlSm0HiKel06THY0voRztBpR4uRYcgZUkG
/mplu7GoovszSTYg6fvOcXthYiaW3vC20ZJtPyWxcuaGwfw/WvsLlKGmCwtBTSLf
Kfdg5C91xGj0cnpCNYntMIA6aX3ElYzLyZcgceBBbBqUjGdEfSGREj1ZT8OKY9WF
KWInp+lykpx0XNJTVGz6b3TjZJvaCT8ijQ+6yx0MeJcqWSeL4ffJ3AOX4MwtGvH9
u+w0blv7uvw6rkeNFRtl9kdXH9P9nZhBwOk8xVequAzIZmkzoq9IRdcwxqzpdYz5
EMnDxojMLEqIXT2bOEc/OBwsxROcKCwB1E3jQXUO/LNhdPdvuuNaq8cAXqGPojvH
VdpSXb7bJ8o/N5DQKaPHx31ewtLM0iu+f8SuskiCV+1AhLYQtyQi05ss8hIwhcr+
7hRbFuWIH4LCp+ccYAYgok69lL02X9/51lpIV82m6gPVget2Ua5AvBeVngGvFZwQ
hwwnyGHgl37F/u52OoSHbsDAWEtiIumgYlT8kqS69gxmcyHsDpraBEEx6qLoidwN
ctTkL1bKIsYWKszwMDWQcTJoCy6l1CP1W1SyZvLR13Lb7nyX7+WPCFrIKUyKiEQe
n3FDA5dbhc6JaT1anR7dfACQIXgnIo+IFjs2WrArIxm5T5cswwGzI6KZtJ3ciEDK
VwtTbBaQTsOH+ixTLV3N0Q+M5f7bRce2o3mLYQkeE5h0M0xbsGst70yGah5Q8mn6
9mG9zXhr0eS91WEkpYmBgEPhvguiDW9At6sPoVAZXYOGErkIdyJFTONdnMzrG0pB
vhNjVytIl/Vxu/cMqtziLwuU1YvUnzMwaq05uZSzOuh27CwXOzB+NdvVSl1YrKZk
SQR8sNbsacBuO4D4W5xOSTYRDasVRj/PazV0ibeYa/kBQzcxta7ZvT3UFZh2+TwD
tWQMPYmn8/GjfcLcqXVmLHpi5pZDZ4//npWcRS0t1FqEm09xKJiFvXcb/X0s2mgK
c6KjE39tuIsNdJh0Mh7vtn6tErsmuNqCNoIr/sh56z0B1tbT15bcwVcznspSyMpr
SJLR2bvh0Bu9GwupCwW+ULoOJUtVeNf2UJFd7l1LgL83Z/CetOLb0cTt6czRFxcD
HTutIL6GiRdr/wh1J5vFmulf6rpFooI+n6LIyFXci/nfbpT8eG7OHYc4i/xujiHU
hFNgPbJMdNPBU9kFYj0n1p3wOovULhO27TSnguUDrgWMZLeLoR6HREcCNfGxyJap
2I9OAt1Vvf2qghTW3s8IGLMP8v5Vr1/8T9oWgVT4/u3cBg8W+dk00T9F9XRvuSzV
6LDGoOVsy4UvFag4FuJdWm11pJPeUuURQqTar+4xbq2vK6HYPn2fwNWblJ44L8mL
9BMbAyCzzD+C0g7H4dxR1wcdOgTKtdcTICZZnyxrk35C1bFHqANTM7VDnuAjMZNo
b60ypid2UiRAWCd8e+btaD386u0OVq39gBtB0c6+2H6wQGZE/omap+ltBXohE1cw
Bh+mjwA2gzEy+2v8a8LrnRTniy9HR5uYCa6BivOdwxug3DP9rA0l4PJ38FKbnViK
WXO1v+o8/QQEkpcJbK9EZafINy+lE814d4XJQLQyUODpxw73mIOBf6Jzj8uPXqZf
OWr0xApmFud90NBth5pbFHw1IjT8U3SzwVncnFQsEoC9TDdO22inYPFOKA0C/E8Z
mUMwRdUAEuoDZa0piibbOAHIxDAvKV6BTZj+QwhrGZuJovl0UkXrZRdC2QllmjjV
xEmOVkZwovcXScPLYq+OMhEGdm9VR338dSITghmTjvnkR94/feq/X241KuCXTJFc
DELMJQgZcLrTyfeNA5ohBwMTknPt4GOxeN+HAUhNO5tosKNCR6jzhXm8nTOzzfkr
b2NILQK1bu+jN0WnL0+F+V9JCWP33mfwH+e2HGQHcu21qgQVTFr4aCKWNM+sDORd
NiNbeOVVRyoWGmYh+HYQucAT79Wf7KhxEgd/NQ48eYRSwFz0hVyWrXmrODjwSjhC
L0O0opMJNn72GLWbKqHpP528C4OWwLVf9CnRbh8+jn6F7zG/j/R65dmpP0gvbLaq
I8DLCHukdgxGEw5mtaRnCLk4Ur/m3rlA+fPAqazkTiavKCDAhSLk11BFt334KXuB
bNMWubjg9+WUvZ9+1jjX1Y74yErwCUdAqsCQoFUrvwP3rbbRKqWv8LQ8CKMhVfr2
bAARkzS2c4uGUZHOV04wNtfRGtaWgOyYFxMs3u0zIkGxmKsCeLfr6aLkLIAm7Byb
`protect END_PROTECTED
