`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LzqqpFOFt9l7aAynIEEzWsJYZJd11pTSrV4iMWHhwMoeur5GCjOj2afw0yWSUwTX
mmD4wlwz3seXeobaGNi4eEhKgRZdC0FbYI0Gy113OJcGlVzczpxUnZKHEx+hWLEh
b/+0x5jMnkFuPAV1Vlfdc7UTqYrdKUIJK1bg1tlrLOPJVfuRbtbV1TfRy6z1UTiA
rZvvr93FX3TkS/Mv6Fe+kT1k7S4LPzm2jBpHJgBnIPnXfvWPkeyPlrVZaEgUiaOd
1ANxK9slFvwTnGle9pKTENDL8JZSQLmO1CPxCVZ3NqROA+2WMO5V6PLczRrw4rQC
WPq85x9S1/nViWFkn3RnUS7qewpDYSAobwd7EqH+0eoboDFD6t7nSPmqzrTWGaBU
dhU35CW4RKSEyUZ7fM/rCQuZjPvwQi9myh9ZOS4AMwE=
`protect END_PROTECTED
