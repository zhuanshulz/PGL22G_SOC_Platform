`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0axBtr7wPoMOE4XJ7rUSErYidUEwxRDfEm7CIp9+Cso+oRCv7KxHkI2XYTf21y3y
9BONpc7g8gBMhoHDt0HX9rBg0xWsdSWfIuBZfTdtx4CsITgPPGhaK+b6c7ADT8yF
jQLFvbHP808pUtnxk8lnP95E+w2LsSSaQJJf0B9JoZT5Ld9dy57vvSfUs3M6JXTl
xTA3FiH8WDylSQW9wlrYvZ+fmMoQQtE2buBCCs1vb7MbWeaDkI8rDVkwo/DvmTN4
9QkQhOu+KeYQr8Ot5W8qwnT4Yn/UFGLpt9wJ5ZY/ZAZfawcpA+oarZbZQ8YXq1v+
DzIoY4u91aMhmqeSu3b3UJSkYlLMdZy+xxs9RzLIWnhDHbwZ8QcboLxyDdoQRanr
TBfixvZsqMdwA/NhiGAnDCLMmnLcLoiexpAANNSsKtXCrk1xckBKH8Bh25VdCVUc
5a/Ur32DelCoF/U2iieG5MLQY3dJ+yHvldCXrab2HXE0TX7IKGmmppL/OiMsaDTr
d3Uuvz1rDHZaxpNA4puvDHkidU1OC4LYHch8bAFTAZCab7oVhNlv+KxVz8QQmW5C
1p7/XPL+/McNkIgRymrIbSFetYFefwQRqAHEYjS+ysb76JWxFT9gPwJOtRM3zs/Y
hCzW2l49jS9UodaSzTW3caFgRHYy5T0mSXAyR9OmXrH+8pHVJ+MHp8m+9WPFSZlf
dJawO+c2sZmQsAKK+Cw5F7yddTL4eEcFQcQNMgE3ukxtRI45bumXv5qTCxBea6xO
pHhZK15leMHFpXm6DVvVIgQseoya6RUV6ORPSwj2eOSu4WDEHXgogD3Gr52uZY/l
GNxNZnUEjn1HRgx2uN+oTdqpuGOerahtsssOtvbyH4z8BmL5QZf2FEThB5wYEnr0
vb13lAMNdLiWGb1OKcwUnMT26Id6AUHNU7EUId4l84tptYvZdCccCvpIKb0Sp8Ou
WwB6FoFdlv2damy129T2iWjQZ1Zmxo0CiuYfNYAbCUsVk2+qzHG8UDFxBbr23+qT
Q0NdKtfzf0/dMLNqr2XjQeUeWrlzr1t90l1gXbVybgQmpqKkfDn10bfoBOdyOha0
rcgUluJ4rKt/aeB1riG7aJsJ4246cAsxpYqtBVIPvOkMCE71V42AvI2k6upxOuvy
h4ktr5LKZjdOE/Mrq1NDsVly836uBxzB4Urn0iBlVaBg53X2aVjk9EHHWwaDLqy3
9wYV2maAaZ8xcTAI+FWZMgidlw85DIbp6RbRjjeGvbX+aIArQ5MZAwT0zgrg8gjv
3k8p/QaugA7S9wLkz0cH6GvsrbXiiCpKGnegTPGGN229NPtBCN4QctUn6fQS6lPe
//CmGvLp4rjbismmBIpTgK/markWCfQQ95Jkmf14O9m3wMUu24fTbe624XFCavjT
4m1UQrct05Mtx8V6yQWiEbRf2YhbCKJutPqviKk7guKc0b7Llhb9kJiZtaDO/zJl
wlNV/XQZVou6KE3RqIwwKDO6qZR0HoirOZS0HZ4Rv1ywsW+fRkZUH3u5XCvM1Ph2
fKInccCE+C4mmRqeSKK24WsLIkcDqzHiCom5ewiolC1c/6+LwgGsJSdQcV8dpZO/
DA6XoCIRvHdjGSzDxGPzUPC5JnuhM8nbvZoFfbO+ROb7WjVaH3V8BV2Vfo5LGYrS
twChl6U+VJbhknf+Q/cYniEFNn4F9xNC0m2r9cUYFkJdZUHgHOr/azUuTJD8G+b3
Dvlffgdv8tBdiiKoQl0gJ+nkTqchCI9vL18bm8pDfhgq9+ev2Qs9ye2B25lkouKI
5Vt4Ni26ja89pigKIJSqyZH5iKxhSfDDzCXlC3S0z2zri/9vb7P70GVAWg7AUxkq
7MF0XPrMqLPjSkEGplpyzHszLToka5DoZt+H7LtlO0heXpZBVpPb9VmxEyNil7QZ
XDyP8wZdiWoww9lJ/s7U1wCptU3WocxxmtKBDLnQvgi5IfZ9QvdSp1XMcGbMOF2J
JhJju1RlLy31geSWI9z/w0V/qaOVHdAYB0qp2HupCCHOOEyaZQFNuwPxDnDuSBWR
xuBejGsu8hcQAdm3nP40nISRjEGJBOaPg/iBIw11VkscxHbVx0tvRTMLaNXA6QJt
+ugOvNN2KmvS6NvbLE+xIgcr2dB94k2CmTYruUI11Iu+cqMKzBzgiShKbNzb1U5U
xZpaRD67Zb3hPgONOhqnylV182IVsaAUw+d+eLC87RQJXLYbFqP0yiAC7KdkYr2x
PznlQnTIOOwpNIGyY42xZei4aPXhu6lj+MRTPaubZQWRPA77FuG6wKyWSYnkdv7c
7A9Dp2zJypEJVkahKcEx/t8zMSxnrBfyV6I3Rl3i1RgBKRxEv5ByN/1yO/GlqQn/
9XXq3PalMYF+UuyDnOsiNwQ97abITs3NXrShr3a4LzW/zr/kFBGbS1wW3/uVUar2
9S3Ni9gYA+vyHZd1YKF0j7OZn3qVUOtTs0bslIwO51IVwQnunn2fXWc652tOJ2aM
lepuVIl0XWekcFnQIdvOfwekqAygGi4Zjl0ooYNfsUSgDISOzNW/UVMpPiWcMwta
ToNLzgt0F3jcIJHcSECka3PH6R8P72NTQRX1F/WsDQNt01ecOwMlhD/XHaEApWQI
SBSClbcH4P3rYX0SGr/0q8IcBJF+2ZNCdoQYCozd+McPKZ61dFHSuW7v+DnfgYwb
K2Vjtqd9N2V488LbiJsXeac7Ekh7REyLM4SIGvPxvVV9SEOB8KPCEqbR8qBXAVsE
dRyOCNEBLuKo16AvuEbrBBMpY/A2jlHiY8wBXq5GH5MKVxE16bi7P+ZZIJhGo+fS
GpGDwSMr35wuBbjR0GqHB44lXUpgwPn1m8TYfNfo5I7jZAwKmE6FeSbSRzmiiBES
3FbKCel1hFJs9OzcDdU9rbH70aAWqyASydW1xudj9bXGBv82cfxCRhUo6/W4eK0i
NQ9WoC6bUD7Lo/3OvbEo4ePv6KAsyu+oH07GJdZdnodB6d6M2n9hyZttSkhULrT3
0cee9Pdq99KyeUZl0WBKlzoVJRS32OjHyNkQ9ix6nEiqpCqTuh/lXUwRZOMSnqcw
cQRabpIpn5s92bYOrcneBth7rb2OkAEoXUfBTDjzrIEjgk4w+oeewVylGbb7P4gS
O94TwETfPaTf0PL8vWD8XcfjrIeAaZDpCZwSFoEcAIkWxVl+IEEBN/QGSJvZymuh
WXCtkoaL1E4yC3x2uGDR9w4I+HVLZEDP830+KHphdltWhXsbFijX+fcU2eTK7G99
+pk2Nv9L4iEfZtyPE0PLZRYzV/xxzWM7QGwMVOYUaPfPqNv0OOGtSvPOlFQ0Gxjt
nfC3Rcbt1TmWMrE1oOCUOrEwmr7hjp3IVoMEqaHcL/YmaOz0BU3DJJOFBys5Mud1
ywSmbLRuw25nmRnfw65xlQF/DbugyGUxfx0Svhs4ENjRT0ol0hrhcrBpe1Itvicg
5ULDM5Lsi78LyPVYaEa358SmB/pKuaW9iKYiw9J0B5GOvDQRkuxfOmLTbm+WN0v1
qZirkT/zVnmRxBDQv1Xbsnz52hjYhKsETGKoOFV7iVjh+Pf/aMfzmwMx7CZCA2dS
YIOOOyAzqBd0Y5COg3k6ZU1lj6SHmxgPZNXuj1LEgvb2/jPla4tNmr1TLfWHc65D
8Gm1RTR9RF5G3DdQEgTM+Az9Ynvw/LmDRXh9VQEss9qMVAjGOl7b98F3/2ZS3iof
RSlkWzbflXWwpl2CjEUDyuS1Spt9lX3gD3INlZUbOtWda+dXmbaLI+UtNUAdnFLT
5b/WZb3fwgdvtbEk6PfAoitWxSTnZ7zVcwzS9wqLdxNXoHayRY/23yCp74vJwm3o
vc6LOZUdGLiBgNvavXhrM9pKjDfWXJqiaRL23AxJglSv6TcNHaQqIGT13oEZJl5a
R5XFJpJMITkEiT5lfTnQGp2NJjUQnhuXPhCjSrEEYxAjl35PEOvBd3doWgAlyhOk
x3NKGI4UCwTkYmYuvG5BOt+j1TVe9EOGQ6w7jEBMco6dHOUoFMkBen2fayG52WhQ
jsGN1WHX7mokOzJvDmjcfH6Vatch73nl+0foogF6YkFMwjM8AfOZ5SQNuOSjpw8O
tDFGoSs0gM5ZDzUQVf7SAqEfRICpXSoDMfwKDpLdWrhnGWTRyRr1+6O3zAfchpcz
gbDurC9JLLTs8q4LDY5P++OUilKjg0az3oNxWy61TEtyz1/0Td/gssHPrdoWJuEc
s0Iwct8m2IDh7DPYY5RL4vg0Waop1H6+DsksSvcFuXjYcISzw4ubkahNHb0yUqA8
hQO0qYKPZV7Jk8BLZ0j+Fri0i73zrWxcD5k5RGDsmeiwgyUdamis86DQflbijiw6
2WM2ER5GWW9vN6HNwKjH5YVwVX22kAPRjFfK8Mr62zJG6ywtQ7q5juUPDSbEUxwu
vO6Z+oyOhV/o4ThCLd86Z1zld+YeVPvFJWCE0bglnjLWKsD6rOXZ63TI/2qb7gcI
ZBiTO5c/nTNX4xr3X/D9VJN2kspLC7QcxlQOMtYlgG6oQrPloQppG1uj2oj9SDig
DGdorOMyWf+n1WdRisz4gubx7R77rx4kOOnCgQ1X5Zwtq6U5TLCKTRnsAVE6bF4J
FV00mg+ikzHwt8KPmnvIUUSSYTVFKhmBM7nivvkLv2QgzIugRn+gLlhdMEcol4v7
3VJ3G/Yi5NOwzadU+j59JLpK9KakM+qOJdgTN9yzvNhXo6OC/m2uSLzpiXeIv83C
T6m0ZP9fqvoBAaRPFYVYbOMAjhHH2VEGsRunz8ZuPDMUihJPWs47Xv4CyL2so1IR
QIwmSdk2kFdVi89PQP+yaRAGjCTVMdyFhwbYcx1tHoPZSJGUME9feNG561ayPO5X
j0dPmMo0DwVB2Fjo0avYwwpO5/TsBdlccyYoUkcqfMwE9eSi5su3BE1pGuIlBTcA
B5Yi9kUSRZ8Ri5qTT0ZjV0i2Ga/DFzTkw+j4eMnRDRrPDaghzW8NjoNxKFCoK10h
B7yMTzP71zjs77Pmu0xYSGbuajja3ipFc3OY8wHRzZC5qT5amNWUkHOO5T0scB2c
w8qghCCfLcCOnrJNBrWqDBsIZXI4KIvGmG4s6Cwk3kHw5qZ8bwXogmsMKDEu5Iuf
VhteZPwqyuWholO/M/e8jz+tqhtDV+N1y5a3bmMaH6iruMRVAHIIS/KWIEtp+H/r
+MDJJb1sD9t7j0DmivTXI90DeZMF0sEEDsSY6tilemPU+nzrZPtB/WbKFg5kwG0l
J5R8onU3yzZb48LyHGdt83NtgA224zydfpUgsVfybGoVOoUFnau4pzLNd7T5fIzh
XNu2QJK8VBSveEYP29HAgteR1aWNryznPLX7kTczbOwY7ZA4L99HWZXMq41DcFWp
0dJONiBxiwmDdt0mUsOfsf30QgtbWG1JJYwtDAZKPSLCPQD2CzzzZX1YxjE6m+PB
0DleNKkGfhAiMpesGd5YNGyljd9fFZPDN3glh/Uppn7/g/ZwHNdaAsVcAo/Zzdb0
U/5ZvgrrXqh+A4vB5t+FSUC6mRtsUAF7PcbCGzyNS8zj876kzLU75I4Ga0raZCec
T39/no8RfBzIQYqKxecIxwpY20Su+tgTY5jkx9t9P522xvf/G0tzbAtJ+hbGzzyS
BQrVLMIWwBPd3J8oyuJVRRcX/m1Xw0Bu8vmk0cwEbiu/2JA9kVIv4UfkDTzj2blr
AulMKBz4+gmU2emyGLcV/0fXoDSmmS+DOVS1Wo4eVNCjphkhzoQfOnOdxxF6gOoE
rByVGs7ZnzOHW3Hr4jt3HRKZXl/R2B8hpDBIzsV6YkkJURi91baX4fXbz5jOkQTw
tIHYgp/e7638SoxhuAdVN4ZJXJ6ziqkQk2lcZ9M3rjDMIG1biMW7udx3nwNGS83S
XNbB0qZKHXjz3FxUauqt+ml9Up01esaBK+0QNeVByCaDLYWQ2nj/YPq86hU5el0E
Jh2qetFqaLoEm2QWfAEPuY4erIyRg0I1bXr8iBnQ7QaYIh8DYsXW/IKelPBeV5UM
FQnO93EOIeQJfdt8mZX+UNrmCIVDG6WZBJGBQIq9O6V8RPewKw8eW3L2KCZ5OKxM
m88VKXTTSROzbyJwgxkP3uAGdlo47fItAjb7s9EbgAE95UXo3/2w4fzmO6qPKukP
56XK+XcYa+PwR4SBvUIh2q7/aXNtbTAzbHQL6ibHCsl5LzEua7QAOwVV268IGLr7
+gPMd5oJKV4OK9K0QuTsVARsRa3p54JFY1HecbAYMIiUqHtJiCje/4XeXgo1e6FI
Toie5TC0xNmh8ZdfnVO2oigHyq8C2iGhE82QEPhMigpQQNyDAz84lJFXTJpyBscP
iK1NhE3W37aGcFxqXqKBtIDjGjEdL1YmRrG2PdZmC02ECHTtsunU0BGifacEGPCF
Q5yj+9MIJbnIJrQ9bSbJrKzz76wx8AIjlLtu4CSlbdc8twV2q4RBEH8Q+R39Zbb7
kmruXEBSiXKyHN7v3Oox/9oojLlGDR7nnxJAMoWb4CKEMAL4H5cbSkTcP0YyHU8D
jgerlxFSOF8TqApWoCZhbc7qHjLSYh3mxe05ocDZnX4cj45/wqazPFLZoVXoQI/M
ph3/cK96KsZgdeSsfOT8qOYxr1DB6G/TFWtdprovZzom6h/EFB9phfd2Y2L2sKpY
SAQCsFpQKmPBsYhLnq2XIa/uytA2yoRQbxs1uBqandQ1qDjpOv9t6L3KAA+uf3fx
v5uJad1H/n1S59QDcF9s0jf+eW3OejokGxB8e+qQlExCq9bnSd3CDbh/CaDW/T1R
88epluq1lRCrNYSDG+d/lv1mGHSUA708g3YAvj9BT8iKyS5Mh+3X2OksAlHlB0WV
eVhJ8ThTfHW/t1ip1niYCEMNfGFlTylEQTU6hCZcjo0AN9MIG3VyYZ8cDJXp2YCU
L4F1dU8HvIunp0XHOzUWPgf3eh0iUQ1CamGpiHkQpQ7MOS849ugIf3Jwp7Ru5R+U
TRymeupFQhhRKjOCqeRmOyKVDbPTgQwymVS6BcWHaUXIj6UIW3jvtySqLXYMD8hV
H8biSF8s1gXBDYJlqrluGmbBwyIYKspBnMmoUP07/5ctk8rHm306tpwfMv2J85Ct
iDl9Wg1HlN004/Rg71hB68MQIRuaEtwqCVwBIJxrGkIaKYWYrULeUL65kLIgdlxK
r189KI+qLaUKmqGvif4I7HoSrd6K3bf5JrbnTdUggYGx36lhsODNTX13Bf7HPJlt
N+2ke8D8WL3hOCHNVc+Z418ygkJhV0qvxeSql3uVJ6E0A/f3rnuJBSziwe0QjEGk
NWis8NfYCyJ4h2EFaZT+MqUlrejcWRPcLmoApOyJPAt5OpdYUtnVgM3JZ9wNRAUx
a9caU7O/vKG6gpgRx0JnU7wrQkS8lS3n/kbeTDLF2wP+JnMcw/6C+6GIdu7hH2Qq
D817+urn59lRDMAM5u0ZhrXpWuHUj/Bs5d8pUYC58G5QMpilzl4IR4KiNKQCFPt6
f2l5B35Q1dCzCXTSJtGZDogG+rXyGQbGPynPucOCuYXkZ1z61Q/mjahmdJyV36WH
WyKJdAwIaIAm3eO8iuWM5A==
`protect END_PROTECTED
