`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ezadzYDflBcwISh/FwX9kTD4w8EBKkkDutt8t1S/d05kPoLuO7Qg2N/4bT2n8Lot
oIHkYWK8VjRJDCNONg96rEnTe1DAbV8zTlB5X3sOINjA0aIn3/X6Mqo+XxLFGISL
GnTmTt1hvz8khzsLsh0pCbCII9+zZsm+rcaUHG3d9Z0AZAqht3TH+nebr6eL4jbr
dxSKEKhh4vjkspKAHeT579DOpr8bjGL+faBotQ/0wMybyRoTkI66QNBriSsQwPWe
hPOwKFMAXdpb0L9ts+sEbpQkKoh+lzxqDrZ7q+FVYDqG/RT68EiTlJspR90rG7YE
JaHOiTihVJt1IfLBpP0BD1imgFPvVweWc2TAyiu0DqHoZeuIPCHBZq/EoCKg8+Ek
q7Pf3kNYqT62LhYm+w3sp/UyMmJxBTX9LejMkm+l8rJeBIzGGQidQHhv+CGInzci
wWL47k+j7BVQOXPNeP87vDZewBlALpmUmLwayFsKSSFB0Lm0VM3qhKlqQd4PASBr
xQ6AHQDUT48WbFWFiuT/yVX/2ELm5/8w3VCFxAZMOuqsaH+lAwpY0DAwqRfL0DBh
a1r8X8fyGYDizuXniT7UD3Qn1nmjC9YhPCo/zEkkEZoyBeaEQ2gy1Liiq3ybo72Z
fc/TuQXOjauURMqXgssKlN2Q1liktMBFvPIuILwm4ryiNTcWlrxqMsNPdQ8WHweS
yqkKBO+obMdCCrRknP1hlMDAHgugzibmhho3GCL/Ez4VbohDeulOwswj8JyTvm9k
RTvt3+V9C57p+ZvvUhddpsHgTLONI+RPhkNLIlzFJkmaroYdkI6xo03bB+pOge0O
ffN8/mSHyLkP9z5qmHas2OzqpAjn4VRsPvpgDBxXoyFCk3eLorNKR85ao+JKkQpG
M7sU0INbMv7CfjNU4X4pWgMjDrJxjspsdK7dLzgHLjB/O7L6mbDugp3XpxSd+nhH
GspLVfSw2GmLZQKgEGBurgq0VSRTRt2xl3nQMO6JgD71sKnj4aLKeLTZPMnFoLoD
DJ0lOzww/Dk6fzXH2YZ6G9stAUqRKHDMaWA79eGCMzVj8N3qPk2KFAhF6uMjUuVd
eXgNT5Q6Iabc1cjLTLrkQF+Ka8hJE/29jZ3fVeuiGzmCjIBjL7oqJfThnipjdUTB
l8ifblfOAWGuDfVFpVCcYt4VUzUGrurPQd4ys29RHSs/9qd4uopPEeIv+5EozTbV
BFUCHftuQLZoblMU0WJfGpgkKBJITMekIbjuJS/DYZaNfzbPTQ1bCKZbgm9gYKLp
sE8WvjA/vhF79ZrQt+RoscpMPwt/rzdgSwjVhqTaO0re4K6YYcs/6SZKe9SCZG+X
1MF1h6E8F9g6VgWRxPGmh8JSK69Nuk3LmvN3tnArJB9QAmBJYSwfY7bQbHJLzqzE
iG3LHsXMwJmF/+/8wmvA04WclPc18it8jlmxUjvhr9CuLKkxcQc1m7U8gKlViQFU
WkE2StXKQ4iqVGqsr+EpwfUwStJkHsqyIOT1g8/YLG5ig3TppdQzKcdrfsSgAprd
FpvYEs7vBPyLoF+L6eYOOkklwZHBdTi+j0pUxO9IlMv1wIH6csbZYQuoOd6oqTOs
RnSm8XnlB1NNQtjXidHKddwNwZU3Pqw6E5w98VlSf0/p8k4U1O7hoURhJTxWwi2m
yo7Iv4g1libx4Z5hwevblEMr9Zh9QR5I4wgbFIhS2wv16cFltJ7xqwp7hqk61HUa
e3i5zUNAwPEOJdJynNd3lvUGQgewlQ/LA54wLAnP5FAORX0FJfXmWqyJgS16Mm7h
8DyPwma87Urtpi10iq9wehURF1OEAl8vrycmvEWLw3kciWo7xAopwkAiYzNPd0uA
7kY8e+6EuYgZAixgXjRxknF7cUEnUUvLTR5Tm2nGnDHEVCAaQXMAuiB9BQezMonO
eyqK+lG/jkOhdrWyoLrA4wbE9cyVt7XZqcQGhZiTBJGINQRrZtrV5AXfNwoQ+Znj
Dman6ZmLJTZfxh9DdfDXTUZuNVt7zeD1kYl6DuWzqO4rEx5h9TClQItqXImXyPCv
0qFgt/g07JG2kfSMKJagjq+1TnR6Pw3gm+ovrRYg2gAWZVoC4E97Wtdyl19DC2Yc
PDpjsOLqXpsZhBjSSJZ4Rgc+B+qzu89nqRD6Dbev7w+HcbMYxaqwItKQKgBOtZf/
13s0BuUSM+iYgyyxf5tTjglcxw+i5oWPck/1hWMhBopT4aTmYSa5B5/uWfF2gAkq
EPahpN+u1E18Nf3yKFjxZcNc9iBLtTT2ZO/VvEF2Ua41fcmghSm/sDnoenzbau3U
En7wIcIy56yAhtom+/ZIUC85A/wjRJ7ShIIdrNOWin4PNvYG7280CxV2CZ2VBcRB
1zC8Bfo3UZVvFFGxmUMBHTq2ljFOFJ6JTcUofwUeMLcIincjjqZwEFCKNtjIHeTT
rZaxOTl7c5vMYoZJZNPbWoXUVlf/MmkDoe4EawLkCkfYUJke2szenU34VmMEq0E7
SFK+nOXrz1KyS7ggex4Uq2A/x5onkHvSQUmCPh2v5xlYU2740uLDA0D6wZ68XTD+
nUJSRdlF76KgRZvX73ORVphoyhIX8pCVSOXUGdHe4cdZCMgSqhdZAIVarq/K8kFt
ZB0aefLH0QrgSNHbazyJAKmLdQJ5Jsg/BiED89kDrMPq9XFECizrKyB+bOJQhfEy
eeuK3djE2THjWKOgPoXUR9bNaUoNY1nzNVZ5t1cMXsuHMlRkvbuHtKOKCGyYtkNr
eqvyTFOFT3qu9NQJ5RfMuZTseR+G8QhWXnvkgsZCXtsvYQuMgnQdObQkpB0QRBn1
1YJAyF2PC0lWafpK8KxQ35y8lQlXaUZLr7FQP86d3Q1JAbuo2G1E4G8/CskDhR9C
ZOx3TaAuVkvAxKaxRaFtGriuCW5uDq5UJY/W7Dyua2RFUm8CU3C28nyP4cs7lzQM
Ry4/A7CHTK+ejy09SLwhWpOEgfWTzzot/TyCs87rsuRwIHr+FpmWKvVCiYtLwUtl
gOcWnlMUmZz3kUXZuO0tLHb+TPNHpGwlrWysvNS4PCeitreyTtq+mpYfkzkhSMox
s4DuJi+2ILB1zZBl/0ZM7YC0502TvOpF65BMb2eTZinq/Pu9NPxWEWcirVkKgMcV
CfUgN46bUvyAoxP1hJHKV2CKUIkBBCCJoukoj/3MMmJMtZjL6uhkbsSN/tRpioh8
Ugc1rDk8tY7FFb/qumPQZY/8aIEDy9r0PpHfF7gUfTYkG/BXQk/MLXePByzcxgeb
+nfAe+Y/6RBou7bNuMrWkZ2eUE3reRKY+09j9Cf60d9h4eBr3FterM8d5ehhclk0
thGWm+rPiBytQC075ceXRJaG89Tac8bgA+9ifke9/qP+fdRhru2AkCTLguugagS4
nlaLkHLTsr865+rH47LSzOpGfHhUh/7wBEbvF1t0eOEEo/IeOTCRhnEDV7wqhg48
zz/UH6iz+tj6CLcAZXwX5VLl1A3bDOgWFRaM+/0mM4+CTrF6WARlYT2c90TUieXx
5auR9wnk6T0IylTZD97YtwktpgopF4xs8gFbf6igGofkQHJW+ASG4zu6R83+lHbD
Z4QqxFP9hJwtGoTYwRR/TYrKdEpFd1DNmZctc+5U6qEovAN9bK5ZbFUBiXknHwrH
0esnPAbYBbIv3k15nKRt2AAChcLhXTIxqmZyGVHD6sS5sil8lIBc1jcfIlgKw4lL
MGviLzSZMivaFKenqtrmYSkGEFRN/CKV/ohPoyxdFiwooRY+JejXBaCUJvCHaa7l
0NtCvDON0RRFmIpdHCkXazR9Pf+bGqQVOJ/J0XnV8Dz0RprB5t7LAs/dfSqlj1Qm
vp3bUJPc56zEj0iNe491suiQEzx0b7ReU1PkzKMqKqFxA3xLyXDW3T3gdrDqJRKm
Uw5e1lcZdlgEKfhYZlJ1QJvMle3IOF5yYiNvW4E87a+L54nA6qElFqPN50JmoW0Z
kdMA4BkA/5J4ESh1SSGlZszPT4raP+s8gYme+XTmjk//yM/FQcBkPn/Eh/pcoJ3C
OoC2KIOZLSqaPWlhnMthYuubmreP2krD/JorTLqg6U/Cd9z2N+joXw8rdv/BV9s4
F2dkb7sgFwAMNgqeprUdgQk93KtUYWr/xj31ucHFKEYwIl679J+yGJLsPze6VWE7
6F6Stjj2NiyoczL/10uRsxUohKuHJqoiZDBYNeV5jRJOtA1aOeMmeYSBCRzfHPq+
MkQfuMlQGjMg4Ek9iRZffqkOfFnpof6leF/piEPChI++Ht4zOxDy1LlNsjzkuYNF
lBwugOaeCv5OCn4NSjezCAKeGagFecl2KDIXrTBsjSM=
`protect END_PROTECTED
