`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j5mprW8hZ6yD9eHjYRailkKiwEhqHdr6pe8z5cC3N05TruCH54klr/sWX+pbATky
mFDFe8+YoG6hjbtbcvwqmepgGbQr+y4SCHgMxO25C7lrnzAkYRZZEhVpAj94wrVV
aaFlR3AeJKaRtc30x41RVjifyxinwWxfOUxA7CD/9fVO6MxxxkkGq98LR482Zj9O
cvCQV8rILfIF9FDsUqyv0YswITR3Wu4QXMiSu+Q2ne2HHqHrtpqo0vGS5QeYaZJO
jGdYogjB2XxBPBMeo7w8Hw4bEPRbTmX1ev6IOwNJKKumNxtFI7KYpqIvWzttJTdE
Q4vYGhgntLYJ4BwSKtuHx+Gc9rhgTYNbmOALJK0Pn59CJrzuhnOFbMCD035KcCAf
z6MIC+bCz5/lg8/DozWhQzAXQ/29zT4m+i8QUj4rtOZMBqCokWP1eXQAk39cu/pz
qdkki8TM0hyPsTytyRyBOLjfGuKfVGbaA19S89MeDt2ziKvvCQXctfHk7ZjLCVrC
teyvrPMHEtE23Y4rP7ViU5VB0pPSqIg8dkJIaYkE46RAtyZyhVgsRGX29AisNoFI
p7CgdMiTbaNn8zroAe4hEU3wu0MUuP2HhZXNXbkQWO0hLoros/IlCb9fhRnOY/2U
lLNIKt6OwKtBMskRuDgQkQaeOaJGwV0bzzzdaS2h5YsgLDUToLvfQwgL9b6+i2v2
545iZ72ffWvawqVd3ndk5jAeUv26WSrY4aG2uS1aks3aAjUITy62L4CjErYpbQ3i
RmumruCwWrUrQaAFZplEOT94/fBILtqIQn8v4V71bLxaYs7TY7fab/leCqP0HJT4
O/BoBcIkvMO4Sppnp64/OctRfP7EQLjYCLSEQ+0gLHxuXf1Tk1Kyef/jbWo3kHk+
93wOga7tyEeiRX+I4x+65fEo1DJdGYN64NzafXmCTk0oevzym+mnWb/Cw+79VAdX
q5S7qRvW7D0Nql+ZgoTGUqmjYfC8eDIv7h/59ebJzPgAeyk5DOxyKkTS5b5JFIV2
bMnqDYrmWxxN/NvHkcxSFX/CfdXwqo2ga6LOiVv7GV5H+1AvtZwRuiUcptgw1IZ/
f9b3pq/5TTbUj5sjyseTliIUEyoui30qji3WcXTtk51xpBjKbjIuygRnV2hNya4F
60enowFb/s9O8HWFr/dMC3HqsFgY7x8lUFcE5BxIeanW27mkjJ3nmSu5dNM4MBtC
sm2k00M0o2oMQBu4onCmISwF3CtG7mifRQBxqiWrlmaZJ9ZPUpQH8GiK7y80UKQ8
LNoUm0qNhA34xHqAjoswRIgOKHH0XG2tgEL2obPFjk5bTG/Ef+g1DgHXrJAQ7/BG
t39NJzv2VMCUID2RXlhHyeXBi+/HXZE8mNVEEjNFi+BuV28U7iTl0YuC0PqD+SAk
zE0jYJt/AJNFXlcFWYkqyol/1lgbz5BbK7YTefL5fsyNkVjo6NwbcWZ464gn0zzc
5U6SOp9vJMc/XrFIUEUJ0qEn6TkgKU2W7BoS3nmUM5htXgg+TSKPfeLsNRazTjgG
c9xxi1XbWTiVbRpSypRwRCk33G5czIF4PVxkEJEgNBrkRN0XaLK6QALhHpjyej8r
EeiimZncCTbBvwJ1WzI0n5rTkoUy0eUshu6RkswH2WS2le/fs9Cx9aqJyrYBfaOn
x9AeoyqecuJrvJ73CtKY0kPiFaBxBR6zK3bbwvS8RSnRRM2n74kstx715HTq5+3c
pGB16MGQgp/CXqufeObzaasMabb7RXeOFrck/GjVsM6ZogMrOSgpDikZ12wJcoUw
UQoy5rC6WieNQDfsDuOqUTF7le8vhBOA9fBrZnnNVHfe1tbNCWV7kThiilp4tmgy
xp1JdvAXaZ/4MXGwW8P0Q6ArY6sQkkBNHp/9JJ2+vyBUjjyEqewWKtYuRGZs5Cth
ED41CdhXzmgtUh8vW3DvPrMvJQo36lH7Zzy7Law2WSbXatTL94SJdweX7MzavaDt
MuMUgER6KoKin4FSRGfUvvNT3JGg49jMD5MTSohmyX6PRUkH4bDGPHxjT/AABs/t
ddrW65jQq1ZFH4SU+ZtF2LQVEXe51zLHGN+CUeqYA94gaKjvMuYVd+c9E97VhAUH
wAZi7v/l6l4Sa6K42/xh7E1crQ9LK65+nu50cmUtJHh9i/Pd6jwW7EIHLsSogYOV
MlYgRW/JriLJ9EfIZyf3V7ggvGPyOfjE1x/xQXMPkPrWL/3MMm6G57rYzcGZ7CJ/
6zafBLlzT3vJVjQbrDINA+9/OmTfkdw7dv/bhAQp4rN05KIpReymNz4D4pfbSs6/
lGBRuyeGQfrBN8CrIY12jpZByeYDCdUv2nWBCHg+InkXsoIfwHG4gJGsYZ81tSMO
3w1cS3vo84EeyD5aV4DKMYRat7JPXtznJRiRYf1cvZmw3ues5A6mnaCIUzPaa48Y
+N4eaXjG07DsjqYAcFDAQBWiHASyqEsPwuvw9xO2QAQIe/SQA4Ca3kCtlWy5PChi
Zw2/FvIUvpX7RYKrmFxWrVP5LkJcyItZHWu/YMjxLntUghjHBiwzcX9D/iI0K5Sc
uEpbVJKqAPgKtyrPppLGSL+Crj/Ek66s3P4DrkSjJ029kEt6MY2jNbMFnQyxHbU6
BigCuSXt0UNeZDNCbJfyKyNNZmuwpJRgMYLf1uchxaLO9a9vXufulxj7EhMJEdbv
4CbyJRjju5O1etXKHMnufbScsnq+vOUmZe3OC+KRr5a7WLUOtvkZMQbsxGNgojgH
Oxf5avhmY2H8MqH0dkN4GWcD26wW8+DOvR3R+fWO9UCeAQAnh6p5z+7yxE+NBLsK
jKL6hWXcadisNDWUb2+k6LVkqGROfD7D+O+U4qNHQwl8peZsLffcOlY/4ZG5GG1u
oMUF/W/cFRItVUjCa95lwsrIth+KBsQRqzQ+5I/QNR6bGSiWRd3vF8xhPEu8AGic
zUzVRyHvcIkA8qviY54+tQFetegMwwOqPdZQOytFg9GtsF1NuKmqQ849HEJ6dmuY
EYMbvTM6G4o3zb2jV4Mg28fmxEHFn2OYJaGljBt5T3nFfFf2Z+zCLS3l38gAuRut
ofZlGu2l3EPEqIPx1Knro5n4UfkdNEbbYu3oHQwTU423HcokSdTQsr1QJTujq6Eu
OTWUnNH+PzABSZWpoBb4gfp6CEvaAuSnQ/DIYO4HKJGSkJttWl061PV3c7n96PRI
WuSAuOLiSua5rvLdt74eKu647B1PIfWt1kn52RyWYhgTpshuplKGSIgycT1evzEX
rUu1XBS1qZayds6Kh05S/1tLSJWUkRYyD6RKzFOpXkVuTR/EvSCc4x+/I9rkRKV2
tEt5G/5DK4vd6wfTSC5OatIDhB2+NEU8e/Dfhkjcr0tLL9uSKOzmjAm0K8y4uoJK
XmKpQ4j9fzlOI3j/D2gEeSaXfTmEW5RZjR2URNu6YzshTgoipYsbfEiAeX8X+qP/
nB6bsritF48ilLdvmcw8KQnRTAhpAA31GX2JZ84FUxHKhTnjFxmS7GeNv8vyMhCu
y4VZ63WqFifKj8tHVNNkr2y6TWxgdwQLtoYSUvd4Ot5Dzf24yqROGr8MPVJok9Ox
+5upXHwKnDRCmYD3Mxm1KlCXysfSRoSxFssC37JnksFojMpqaF9qOKMBBElfpeLE
M5lz0ARWklZo5YmqNlkyfYil1KN0vHafNiNcFysKd6iUNaJ+fiv2bPqr4KvDj1/k
8BjQddnPYweuv3ZK7t5SeJmOkmruXscrMg3xOGa2/D7/ubeHQ++9pkHpoCPtOutY
UcBjFdwZ/JTH2rlgP1yCwSORAetytGXs3qw7zXxn6SDkH7g1zt4mVUR4l3Js7BWY
ETyVY1l7Ad1iw9RTfuuQeQlFWltQPyJG9YY7cF1LhypMUjquL0EMUn04jmtnQ3KC
ox84CtUEVHlRpiT7VBmGP4mtXO0O+rqhHEUr8mnyW1RxjySNioBNCqDn1MGzhee6
2y/kbY/ccxh9jsEswpFrz8b2FhMqDmHl+eUTrv9ZlLIPHiXuws32cLUfB64jOsUK
vUH5/66/XOAZFa6z9lN2cfV1avxssd2w/YX/aDV5ghDWcOkB5sXJ2GbykVJHaQBB
zMbah3YV/AtfJCi+SaoHVObKIz3nJ39BfCy/sTNpntHw160buHpiT3nxfZ+IOnyZ
/i8bqrnMZJqIhIQQCYIXNLNMdMS/bQRh0XhOLZTN7uJPv6rTfBwNu3tsqEeKIKJM
DCN+q8bsfB1AfQnFu9GrfhXkVnjCUDGIHJ/5D+zJNRGHD2w/IdtR0gZMI8bj4g5d
SiyTxysDvMtQoxH8xJ23Gw2fs3F5kaQQEhdspLbGWcwR0SWqM4DcydZW8r1qKu4c
Y5cx5jttuAhE435er47pptZnaGsq3NN8MUqCjD3JeQ4jDC8mqVApIDeio9WvqHb4
opiZEVcctgW4pWezoTcZ1chHH3kTmBzw9GTAsWLK2G3yC6mAbJYDknEqi8SUi0Bd
G2NSLnkdgC6rMT7f2awDXuuNC2AlWPMyKkFbUdzPEPBJN/D2Fg2y3GU7sT5LwgGf
dA61E1djU0QdbHLDlOX1Q6zZtUmV8Q0SUiJj95VRyt2a2NntOSfoGrjj/pwZGOZX
2TaIA0bYKk+ohJ9yc2eLRTDN1cEO3HzPk3QGghzPNbZm7u2BZYwZZ+EgN8tqKYOf
EpTrQW+8rW6jMggZC1r+QmedHEqV7S617b45JJpFnuGpgZbYsOp0Xgffnn/8uYS8
joORGO5dFAkOeAoI6kJ+c9cWabK4/V1hNyOKbVxh+J/B6HYUvSAal6Smz3ISAWPf
mk60Rtpxs2Lybax3FhUDq0Rw0/7f8DcuFw5ES5INY9oGMxmJWC9M0N5K4IhLmrQq
VhijvdlWssyPPNs8gbNsGPkpdrMoVHZ6SkZTx/5zWUvodBHXjerXwcoOlu9kzEuM
3GqT0XCQi5ejGPLycuvZLUiVqWrsVl5WOa2FTUjQ8w1LKsPweU70P3+WiZ8R5Zgn
HqfGkoid+IZpG0sev2aFiHsfgye1Hs68/oF+BYFDFkm7YHe4lQz8olk53DK3t/AP
E60VmEXm75v/vhJ2iiKnyJBf4rZxnwKhzZL3/SB3U7+tA5voqgktSqwzgfxXtbbS
rATW+NpJnm9GRifdQllE2HmhC5ESpSORVjAuCkMf4/RHGH93DcPaRPwlu95C1OP6
YxYNcH4Fp9BlYzHIXsgzA+vppwm8caQNEeMJN+eFLayhS00W46t0LLbyJJNN0sl0
ijmDihOzPymwzIKS3Cy/XPFJ0KDXa0lqsdNSPYLi++9HVziTcee7jrrTsYRZPMZD
l2ZHI8x2S9/tytAOXwE2oDsVsW7HGldqdMXDQH1P6Qfg+kr1dBXI0Z3e07FzWOm/
ULotSHzAclY0W/YNIy/ly2wlSBi+jbdqY8E4QdZCPpzmHlA9iViCOSw+wS0fQ4VL
zb1owgFD1/dOU30+rAjH7EM6I+Zp806BBUQ+rIbePtJdXk/UGaitXpXi+0XcLBDs
ZTwHOjj/hZniFKY3BcLdjYhnDu4osN2Mrd42GsLVB9YOkw59QC4L/SE/ULdwnBxl
FFDmakXjXwSF0ASrC7rbgRW7g/drWb56d/GBFhrWYvO6WyaEAzoTp2QhrnY0jG42
eLmsJKAGIpcpz6m0SOxTPBpGy+mzoWJ0ARcJMEc2ok9KfADcf4zTR1B95cyZS1Q8
v3lap0CSEVKpA1l+FZEc3VxpPqbpOJuUZ9IYrYuqdXN6yY6iVu1fkIM2VjSG5KVh
c42cho6cL9YAUYQI+DXyEkXujW6fA2wQvz+lfRTNxMIeUVxu0PjEcu6+HWJ4M9EF
FDKWmVBQw7aRgQhiU114RL8C5X0uhfUePszifYT2ARZUjt6Hxo9b4E/5bP+8dh1+
qvtqOLSjb2OkP/JHblXkrwrxcPBFAvmNxJMqhi8y7sEiOK9y0wwggNYvJpFfLiPS
pggYWvoGKP9ycxr6TlCZjqh650dgTSmt8cFx/cQzXI1nB0qa4+Y3G+MNk3acA4U1
Bnh8MxQ3cM5SGIMhvchlSHIoZHsqNSY0mCtTFq6L4Kmu8oO6Iv4oVyvcDttEDUmL
XLaV5d86MUxWnnacnTDAGsYF73yhp8LIcOX+AE/obiVUGchG7IH1aoPxyiA39t7A
WAKqKzG1zqQGTONnnz2Nw/A2sP79oWaoG6lQtx0irv5RqMdSJLnW5LBR/pP5Hmvi
MEEoWW5rWIRvlwWOhkCL0rnEmZ76B+GzECvMjqL+dzpmSKyHWDTT46OMHgoar4w5
BRWd+O6yWmRNaWRxlsJmHdYhezSwxIGsPW0XsVsmipBciM8xLQ7RiYPVlre4iJnH
pqB5gvKV9CpfBr144jUTD+7cJshIfMLMwQyzMWfzB3YW0+uIHCRLE7yBhTDdk0X/
FdGh6Y+RJEbPXLekZhXseZEv6wdmSMMZGSHgu/NTyJkzkthNrlKDTor0JZUs1aQY
BPgr7YycF/x+yj34f3FpFWdM6SHd37BepjiBxTbGXpTqBAP6Ka8EJ95RtEYduvwf
EdEeD6vCxFF0wD5YGVbCrLRrC3mJCESTso0yckCFJiA+5DVTME3voORc6UICy1e+
dgOQ1Ssjl252F9fEHgHvEEnwBFnTxRwuRny+7TwRZ+R8DpZJGiVWS7wwWLYTlpbD
xBKxtOQE3EWlmCobpkbZlcgbMhfkUVP4JUoWC+XnsDnnsLaTuoL+TYxcoB95rIAY
1sLV4tI6gy4hY7CUb1TxcxNMDQYzAq3uiJnUFUW9f7ls2yJP/VdZhgoFUQGH/Z0U
Ls6um4SjqGjbvfVg04s1nsbjQqye4gZ+1nuvH9NAC/JylSiyHn/7Qvy9GOar8G7v
h/evj/AFK1NofFZNKjBrLL8n2OBxxTF0ApTy6A8x/4yXg7w6JVx6KkS9i8jTw3nb
N4KE/P1ClbQiTLp7a2LSF4FMiWj9lJunnY/9Eo3+oDBtofHvVJxZCfWFREgbQX6p
lQ7UO4ezIXhLMBeQSqhqhXo0bVV1jGk3vKPnTAjJlonf7ocB6HnCdkPioOU9WWqg
Tcramt+t0wvp2bC2ZKRpe+hfEI/pJ7BPvTzzmctdXYmsXgk3RMzO93N1Dxc7LQzn
MbH5mQPYQmJkb2uRI/9uiuGgZxe1S19VwOwCbX+FGTm17lVuRl4G1qYs1ikMFx7r
NL2BUCT2Px4cGcCf6WjCanxwSrvvueXH9mqzKinIVu7hAb+KGpXiJjeHogLQZtvr
/v/T27VJQSxrBFj8L5lYsiJPCCHMy066tHkHWNbda5bRIaXI03BDlfLCc39n0jia
NmZDkwqDjL4ozoasjt/zv9zDncYqeaA5AYgxQk8SG/H/ulUiVU1akB+AA5MHDOac
IkNcPREdIzktfqJ/k0Kn0nQMIUL7euGfOWKBM+UJ2lxmqFaNyOLRwY5YPflb5WWj
1lY6b1cI8uwyk4Ex3pNCthixojfZZrLhTlhRZSB5JdWP2evDKhmP5D9qFLNlTM/e
97tVTG0Wdlyl0OwqjcyuTDkqUdERTdbFZlTa+5OtQalKXCYZFWwdC7Ep3ZAq1S04
6whKHixsef307D/gdaoVMa7lqPuq7sCVo2rwAlghcC/es8f3rCT9eSeB9tAX+vyt
BJunl4lIC5A5xsCEYgxwjZS/7T2DgY19+mfU8EN2MX5u4l8pWjbDoHlWkLmhZHDc
TxAuQEEzW+g+ScCfCl1oKjV9D73Z0b90W+tUKHHRfaiz60jxRwlNGc7mQHvcDh1G
E7pnRNNDR+/dVFpIS3wjrFqWeSaO2ozGy/Kfwh6kQIPBhKamCZMLbNDD5L0haTNC
2D8kFLDrsRRxDXmLViEUbSBM4wQwp8EOCepCrK+ozUtiNrJycMS1M76uHJgfXLtr
rTXJnq+rK2nSifKGmhIZljd85BAfsA6LolVk4+7UTuqJjD6wLlj5zLZ96vL6iRPK
HcAW7t1WIy+21F8RMtk/bT7iAL5nP+UoL9PnF704CvljaOluLiMJOIvVKwYVmXwo
bdH4m6Y1kj5XVOZXTp30uCDD0633D/pEa/SEjVNaTwa5N3RPKJZyR/UMqRUE2P+a
W4SdFVLbyCRpQmn4FrSiv0d4PC3NjukJneaP3xFseSlO8SruY8LG9sB+KQR2tPJQ
56c5FQ9np0Sb5rhGB5Gts+mlYV+Xr7QFg61zkAb50JzeJX/kCI5NPR4XsyOHta/k
ncxlDHjyuoXsVUCblOVRZKIkKnRzLS32ld9IaeHfBfEn/mIgUJPJEiZM0wGt9iV4
luVyaK4Ey0Xvwf5TcrecDMSxF/QyuAKt43IUvobNRckD8IzbRdSp8kIWtOj1fP0B
MKvVCcVRzfZWK2hrVUVOdN4icw7idHkcuYLc+3QFc/c2tsWgAA079sLMxE5kU5Um
25eLY7FO/gcRzAbmQ8nkN6paBnaLbiwJFVm78LDZOzG3/Py6sdNehoGHQ95CnbPV
RJIST1QuQY6OH0Q0rFwqrcRIfTVmOv5mIiz6iq4Mpnj4/BIXkwk6e6Rh/ZxfeKWw
+IMqHEgAY1NRFF6A7tQfnuA1qWzYdNBoABZEkQC8x2ANFciNmDH5rzHUlZ1roLuZ
bRX+eX+LKUCEeiqUGrtM1gc84Q7fVnF5it49NSJq+4tOFM/SSx2/L3MGl9e1mbJq
FMQYwZfT7cUIeZ85KY5IdTuMSiTyW8VIK7eR2JsAnG4/TWhNglOVC+nWYuL4y+Oi
JyNtJLbqWuxcl3fN2OTkUN+t7yW1DAcOjwLtCImF7hUWZcuQhmz2rlGmD8A0aG87
St4X7Iw9YfTq2dOKoVthiX+Ln23HeLHgPDvD98eaXvH+QNWaX2eMn7oSbuFJ+ydO
N4fcSHMfScECgOI7B21+p0HYa81vKKCGHD0cRnAQ+brvCtkVvadVHfHNqvBOVSWY
ZbwsOr1w+HUzdettVlRtqwi72fShLhAONHUXanIIxFyuY0TmzxnmR/8IT+WyktaY
qvp492DMp8P+GeUgh8g2YUWlasuIcspGKODTZcVbMAk0YKKOu1HXt7JPl8b80Plf
SqPRkZWAfbDWOgBb+CEixUoDwHXjSs0ijz01BoeqWAeoyO9PJ+YlGyzkMNFjnhxD
YLhrU9aKmbKtOE5/itxJJ9eUurUSw3hZzZ69Yd5CGqAMR/2JTidBRwIpCAhj48o2
Hj1etzOVEKfN50PbRJXckT6IDCNeZ9hqsYuINaGfW/Qwrd4h/Hi/IXGSK8rVpBFE
Ayx6CNMXbM8okZvsy+SKoXbK67veFnvYb8vI8JBAzf8Zy8R0v7bidzyf0MilAX5O
d/h6jCTFtDInsCtfbXSXeADPoqe1lCPlJnBuW9INloKG2sXgLhnM1h/RoPRxr8EG
NBpU6Ah0/eR85De75Qk1ESz5B8gLQUavcZYRh1oyDLsGN0VgjuzH+gmVAK/YVKUi
hzUUUSXBFtG4eBx0gLh12m52BNFNSVtiudHYosKjkU7K/4vq2K6uK0tjgcaDIczm
i+eZfSqY5lcIaYHtzNt2lrc8QbBh64kpk+9VcwyXK6dYDMlu/GlkGkwSaaW7/GiS
F639fLxk4qsfuEYpET1N+esqosZ23ejanG5NnOW2XfUYlpQ2TM/aKPgPnOpywD5l
NSdzFUldmFMfbibMSGrVQ7d7pKbJ/hZkn4KZIAXM30t5lrEAKK3ZILkimAkBpBV/
Yr7z6cDzyh0j6UdNbmQ3kHyXmLG2J+/IwCrnCK50gzLAizVWM9X4fQNtiLNs2+m4
PdULn9lCTEkM4Kbm257ih/zDwkWHvB6agNAminTQG8R9dQsaxuFY6CugSeVtoSsv
tPl/VOwY76CHdTOFvCkzlUVywL1evzj0k0QRjfOLgoqyCGcM52BbZ14nsi6ZRG8m
RWuqOZev3JxEe1UIcHUTUOrBHTlTpqoxlNM24qZ6dsxg5HHOKjwz7bSd1gsRYz6c
M/aQgtadF9kw0yWwy0nKmrfXZ+9vqjBygRfsBX4ijbL6tlgUkaHC+796siVFGAnJ
cmilglDEpaRzluU2HNkZvItFZC16FLRje3OFzZQanUE=
`protect END_PROTECTED
