`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zmWPyAjmw3nQPFGDqnw+BxX/XLt3HGdo5rWBYD2L87pOYAo2G4VxhSIqyWt6YOEN
ohGO0pHRFMRnz/UaUEryrpixkHFtSm71leLsnc5V7PquM/UsmpZ507nKJXZnkfpx
uZnSxp824U3JFMybG0n7ck2bRP6ZR8a7jIGt7Wbo4tlG/bnPAIKNAmV7NhAJneK5
ESZSicDdNi1ed736qXS0TVTrVY7EDGpF4uNhRqPAhwY9luqxMovheTPJfDglnUhW
lhL0V/Dx3ga3uKgjSw8dnTNhS743kJCAGV9nVNBAH/cW/+DeVeMl+3pwRP10CC5y
QLCgRlZbUi0H1bZ3Nxau6nwpr4GGrZa28RintzUdUFzukI/gyLlgSM3PU2nPMWjY
WxCAQtGdIye1F/Qy+18MnXHcdX2G5Cw2fyP6C1RyeKRYGcbTVB8EdMkS4x8ZvnNQ
fWJ5HEa6LYj1OQcoPKBLCBbJaKJPFSCxU8BTwDeSDHn5mUjyY9LEcW6ZW+kOEIyG
Htrxa0TTQ8DBMBZWsrLEvdloPEXfVbIkKzA4OlLEi2KqW8unNlrBy1IckH1zUp+0
nwu1fhUKhik8k8o6HeVolOsqIu/I1TQsySUJ04n5Y87U/TM5S23yJZJDsmqMeJ5x
f7gBsyc/s+bDFN+xRAJwXLF+IK59QdAP17MfZ+Rs1OnUJIcb9j6ynk5HSUsCQiXM
B9dAWdpiPwoKYIYLs8yRgiaP8OTMU1nP7Ef0rD6GL0OsFZ99Kd5jAg5Bsk5BVk5o
yUOKURDIQNLxuH81UUu95U3PzyUHA2xJ4TOzLGlL9sfKhjqNS74PMYhiUz6Wsyq9
lQ8qHMVflPOymKUGc03U8PbqliL/V0f4v40LMeZi53UGDXMzDZ6gxd2ajHqjN9xw
mlqNh9x0qiDasi2BhjfUOpU7kCpI3rZm2zc6GoS3PdgyRJvcYs9Sqmw4d0zZNDr6
ouAQE8LJPPWHN7DObFtallhwi5gexlcMksXCEHm5oK4DxRYikebtsQo3XgtQutCr
+uE2PhKlo68297kAszpLDWoCe8BG8JuAntv95uHjx9jkoT6YGxE9jWtBnm4WiVq/
BKO68ZPeGzHPvK3rM5u+SlvsIN0ZeYXwduLHbjDpkE5/cXVic8YkNccNBf218f7X
6TQDuIOExTYPiGN/BgGqjcpRgc81VZ89GOCbyuxJ8gT72B0o/ZpZH8bAEe0ez8Z7
jl3jIHI079Zm/12q/iW+qOFb6xrlkHR7IgQL9RATf7dW5RRfQ66rHEd/Sjdaoua6
IEr7rM+xRc/SvxNWFoNGtdMvrDX82ZEGKJLY1fW5hMi3UrkSXu3DxkDDrUnSzlMl
Ft182OR9aWyEsyOjjbik5EX55FZ3RL8zAejoxDe5eOlZNW7LT5fnmPVT0MJ50E8R
dUhcUFJztc/kvzNVfOc8qixZ0F8LTUsnY+xAZWfJpX7Jz3mfEelGIzBERqRt6TuQ
H8YA/0zhdVOkq9mPRQ3/REylRsT80IPYiv/bx9Pi8jx5V4Zx5z6HTM0+/paF+Gke
KaYJZVjv22QgQJGmw18yAmFR+A+1Bzz/otoPlpczO4T+vbUh1YI04K3HPK5sP8Cx
NJazwHb5Vk/hYWAfgM/bmxdIiZfXErVCzHGvLUEWv/BiNfSQ93g5HMvsKlN+qRzu
ptlzq0E2SkQhp9/rClJCpM8NOfDqtAUKuV3DUJDvPT5UM1GGN5n2nC3yEcRmxteZ
kiaAeifVLkk3KAD/r0R0z82W4XrsOwIeXI7D1v2b7BXgpTnQnH2MmMTjFqUSumuM
raaLKHYRnhFz0J3HdKcMNWk0MlMxd25gozF52zvPSTqDBqxSwOQGDAMm1TDkmo0P
nA8QfYwu10jkN/qpouN060SvgtMVzS3o98eDt5DWNwMzjyBI/1ul9M5GcBS57j1J
zDglzmHNxC5UB8g3VkR/wLm/vNtbO+TcyQ7E7K/u08BAVGKUgbZmhkATgjvQCly0
rLuZAwEOd4I2SpDDmTV5cSwbjdw8aFnGaGT4tt2XeVqIf44Ok3WrD55Kvt729YdT
LdsVTJGR2b8Tx+UdcI2Y9UvzhHHkWc6vTD8haTGaSwTiKp5mDseOvm1mX1vibLUz
AwPKfnEv2+L74qZ0Dh0eI4dyRgbkdQ888CBZ02mgqca3UKb1g6FPJXHm5OQ/pQSB
DrI4fU1A0IzRbKYWdC5xT7t4pcdu9u5qPwDBMxYCleXoFfbWlvsbAJHEzr2g1f6E
SX7lDJayeLl29AoivVmnlQhYIZh+rUMD4jYT9Ci/OAjXKCgwZYeF0JnutC2jLLi3
GoDZcHm3ZS1hVsOMyrQYgYtRHv95mgY+yZEacDk3+voE18/eB38p3N64KoeD6Ekt
hU2yplqFN/AJB6GNdxQQYoAxXdilwmioKT//CqcI2l5BVmz2JK6LogZW1+9LteQV
PX9xnTgraTVvNogPylXXwvOPzGF2KaRXKO/QZrT/GwmmcI3BB+DAL5j31z3EUbE5
ysgaN1uatjgSFZAUN2Klfnm8C3Pr+le2sus0SXVr/ymBEWgByqMRd4resPrN8ctG
KnrJOLL6eAAve6vKYEmvrKopIHmQbOHQ4yvUb/K+XGI+yZ6p4Qy0lP8T/AjIKz/d
6Zhsf98PeUq0yCG6EUDH2QiCNvjUhRrdliXCnD3sjTjPOoCOKjPKfUGw/WXkMipI
Z9C2ZsyT+aDdisc8n8TSTo2ICpoGP04acXXg3Zl17foUmpk3ukXihN4tiEUb8JA5
jz6OFtqTrfQ8ohdlQ/wnSgPywD7XH8DhldCUVURH6h4PlwPYW5OUhfY8hmS7sgn9
971jObekY6OyEDrzoabDyQswK7ca95K8NW/+k/u1xAE4ooDSzZqm7ItPGhKjiBbw
0AGSfFPf2/4Nk/2BxPA0qxh3u0RXStSgwP3O8/oS2K50A7uXYh2m9Z1pdsjk9PIr
NHmh74R9mbkZzQfI1kaJWBSP643daoV6N70DbefyU/IeVGSB0bLZI75RbzsFLfPe
gpevcBgg1zqhh5bMLYDKORBbFzcPPhUMP5Q48puZhgKinb3xzDr/pMK9jN2B0+EU
9V4CtaeruQXQ0XCVnU81qBDMT6C2FKaUFM47cVuFxSyzx2rLj5C8pV4L29pa07u0
YQCQ7h9Xc23pF+xcB4Q/MA4iq7R56LEFc6QWbzODaYlZnLE8pK5kVRRdl5TSLroI
nvMymWSBHdKGk9HhU7zCeGyVJe92ncU1V+bK/hIVVlI09w4Tiv7F6WZptOzPz2s3
QVsTp+I5LQ0Y8Xf6iKnwjlzBAC2tXgnZMNaml56GmOCUxjAj7/w4l7BFdaSESfyp
nRPt0yVxtsWoEh9xPX51Tpajc4WNFhv8GwO1+IRP9FuAcR70S5WiL2iDUvcC9jkt
l0WGo1HNIn64F4BkMeGRNgnzK8z93hRK25yxxkvpQhfk1PgvmDifZ5psbos29MB7
HjonYcgYucdobcgYPCYNZLaZzcZEjaKa/vBpoGCQbhlvHSgxbdR37usG4cfsOfnc
t5ekCpZRGKMYQ9Zg5SUsW8M0GL1VUgmuljqHeb1k/nWMzU/VMqcEwWUlq6kj3YEo
kafnjo/tBp7TtGAm7BMRHbVQeJX7ztboYAVb1AL08TqbjOZGp7NpUFqxp0/np4Hq
vRRpHare4PYhLEmAaNkwfn6Ar3jUCpm2lDDAjS3QeX/HLX0wMyQj3pSFqFSkrbpW
3z1wNFmcmvzWb79G+ksXLq/VnvuoCPXE6u3Thu2Rw3DLUr+YopuXrc/3axrMPxYS
BbdY/51tkKVdKpt4Wjhlv1/IbeeA74+Ow3FCmqIMmO0=
`protect END_PROTECTED
