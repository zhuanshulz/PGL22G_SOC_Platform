`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/b4Ans61dyQxoebP3SAx023BuHPRjZhsDDzXKno9oxjQtWHFdnOfok3WlhSwp9RE
AjcCARRs5QzsKThrc3O7LnN5COy52kQee912kz6qpHZb6LI1B7xRXcaq4v+y8Gu/
pjP321MNctVaY1eSVQIQq2aLud1iACr7da/Btxz7dsSPaliL1PcWdoWwkQ/ZE9st
mx3J2epO4F85HyNtRptL9DyqYcecvXkqjipC80zJzFK2//J+fyWfi7WExWXz2PPK
xaJmSRjevN1zG6sB86emEHy6sGZbwykUE9IJ7UZpb21GUuJIJSSrjF1bjgsOzvDN
J+RwX1hgUYj7WiTKBhCtoQmBKDCwxJz1bZ3F8oQC9e81JSOK349VBagI2NEicBYl
S1T6t9Yri7GP73yHhsOzW0D6f9bvY2js26iwL7VnbCrhZCyX4BwNnR2drtSEPOFZ
u3pAQGqzt02ii6GnlGkbERiW5PMw50wJ/yHEoyBiqNs0hBxgY3P6ZsG3SkjZVws9
5553t9t6S8dgyXJBB5JBGby8Se5fCY+XpV6ohVXq/bOqlsl2T/l1xmY/m/5Kc/dA
7+JaFC3BEVUrFylVoM8zctZaM6ukVO0kZJTY6M5HrTkGP5QUvfEwS+J6VwLfh2fA
Mah1P7aPdw3hYavTCt9RKZod+MolgxcbKlT/crEmIIk5xDD5Lpx1SnmGWrxzHAza
eDkC74VEb2Nk+Aaz/UUAP+pbaS+/nlFqlEYOR3s+sS7H6hz1DLor+JvPYDJdDBaB
/+QDlFdWEo1x1vkGxY0CEDcr4owlEkFNHko9Hsbb8nZSer0CsJB6GDlNBzW2NOn2
uKlsyywzYK69O8+qy6FB4NCJjS7LWeAXlrYqpNJhK4OJSzIc/cBzr0BlENOtQMlZ
82bbBS3XvcCgSU0UQxQJfFvssnEtDLPP4pu4X2BuvC/sXXUkW8OUHmlNygcJE90N
yHZ1SsicLoCMjz3ODccPOwfXxj5L7ECUh0Cs/yLtVhqKPkR7DGnZ0gsElahjjBt3
/FmVRZoCZimskEPAKogcrIJhPCPtby07SkkRZp1W2L+NQYv/JIRksmg5kwGgANHY
HIDdr3oWzJpsm1zFQWP1VbBgvVkaIKQES0rE7s9ucjVLOP3lomV8/+GubMvokXfo
U+lol7Q2JT1UOcKrdz7ezlY/cg15K1dCrc2yXBYpZh1N3e+cMHXmWFgtO2ZuIrlS
c84JFXgvTvxmT08lZAwIMXhNdwS3nx/Z3zTzfxOWMI0Ia9i98y8cChwjCSPnex4j
1KiYH+D28RTnMBVVWkWsmuKIo8sqGop05dxZycwsYwYJCxQm59paOXQCl0lWYowy
anlwHxEQ0UAvAhIYPyFBA+n0374+wlygLjQ21vjb+K9JqvZYZtFoVnSa7pdFYXcE
TlwjrYJiHNaW3nYPDx78Ou2QlUT+/mb2BA2Bqly1dVcYV1uJMow/L/Pfxqi+7b3L
hkDJS1rgtel6Dy3JgN3z9HT+TXN1DIXqceUxVahLzdEKW3uFRg1OsQhNy4i9mJPo
YfGnjgj/W9btDfc6y2Ee69DO5diUmsWDiejnV4xvy7hvz3awwPYsznTQrpjwKczs
Go179pdtmnltnlAvLCQVIT9LlYN8dI3LMJC13t/pK3lWCoC04PALVbFYiudntGY6
f+nNKNjDbVGwc8tv/j5D2+lDhnJKnPSRiWAVnmJi0Lwy6yqSW0pM6LfB9Nmw2pGc
HYfNstlvmHKClHWryTIO4pMefS/EdmdraCwVqqv9/nHw7oBvtTjq4/f8BVdODVlJ
KjCClHWdRNNE1NHYozKrE/1kU4CoeXzurlBk/vGnJbUEnm0C5Z/plZPZNlD3Fhf6
`protect END_PROTECTED
