`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ojbwaK6xOjVqjS1I86CCr8T6UHU65brB9RumhyihFdOxDMBLCAQHC99+N17zMaH
kmybJ6G6m50DkoiK02ftf8H7HVHSo9X5mYpyX3Wz4vwlK/o/Dz8RvtyNgsF/4aZf
z+kD8lxUT3ZUKWEzvYQ0xtIGVtL9jh17PMsjSvopjucIAG2iQJY+xEh9XeB7bWtR
1O/e8VCsL8gSbZYWO92XOTTzB5zFEewd2VZ60ruTI8Rx4Hyu68u5Gf78MRVFCt0e
ttHW/TTZvFCx9Rkfy5EMka3ZnCLAadPHTtDOz5pdMS+YSt8TpC9bt9Us7B/snUu7
tJzjCHQHGsflK2HWQp/eZfgwjkaI9F/hYPRciLmA2+hSFQqs4gcOBAgfzshCUQJK
J026hmKE1j4GsIOO4tBVkpyzGjot3eIOk4Wgenhj5bsL3KwNSGhD517t3lQd3Gzw
z4Ydf4BbP/yu5IcSnCA+iq2GPlmycG3fKp8m7r96IFDCVsa4ZWk+HRvCuVmkVLTk
R2tNON5ZaZtXNcEPA1GLizcZn7+vqc8vsr2Il3wK12UUyn4ov18btawi1v3fBKW5
jOE/EU002JebCUYt7JFvPqD6JsI0JQkcMAglQ3UFfoC5f+AMO7rzR7P7qdiBt2Fc
/MdkRYOOgZC6cXOFKgjGby+jM9HuHLSlFixb3pUDiyeX+tz4FQANWQ+RECzBp7Zb
iur6y9xbdempeotZyctaodPiOMhnWgZJi+M4SBzQ9I40szfF+0cMmN3hLwufbWSr
blCws2G4wGUR0VwcyYu6tL8Bw2TtBR+sQBD6mj3QkvBzjoP1QmXTKVHDbTHdTJBf
uIcbZmEdayeJUH+TKRyW8eeCU9sH43tPnCJnyJqMfYDJ/auhZw5bUH/Y/i+FD7Tb
CjIAnQ3nlh/OM7z4DCXPiACnYe8f2knk1XD8AW/TQtDKQ4d9wejBiczyfVjeGjfb
jP6YIX0fl/bDSDTxjBa+VUehg3qM7vKyMHFLIDfQpteDchKJc/4w5uuXvCypZIZs
MMWW40LZRElKCWZS1aY/xg==
`protect END_PROTECTED
