`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBbJDjafh7FkHINI3M5TOKmRkCnlCyysAaQFqlWv8dI4izdY3NHZrL6KBxmJSUP3
PQ1LH+zsqR3xoNhR7i9gNe8osvVZ4kZ07ZHrRywSHuMHKqprMrVzOGIXQxXF/i23
mU6sP3kgdHTzzrXKeajXUmsFmF2KJDBm6wzAXDZO9WRCoFXWaPxWQIce+5BpF0tQ
fP6+K6HlnHz9OvR7X61U+/5ut+nADsOWKKYc8V8OSht7aNTqr9LaWmIDrrBC4/Ux
siEWX+UveE5ru08iHDF3kw==
`protect END_PROTECTED
