`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uBGkc9oXCDrdQ+R7quD+t73GBzcqq8DB6xwVsEwIsM/dnfSOBzcGWCvIkVv0spzj
p0N4py2LH8VTvm4JENwFxfEgEFYRhUUmGWgcb+HbTPKKCY+O5z3SgHfSuTcX0dbP
ABSbzd54gEvOqdbE3R6Q+WsEcdVgkJ4wU8565Sbw1BmP9xN0xXPTdvntGG1WoFJv
kGBVa+HK2YAZ5N8pz+UjRq34aIX4lQja9ZBi4iUuHZziC7e0LlWARiG3rP6/MFNw
3d9inAIuU+GqQFzOagELTUYlSA+N+62LVP5QlZdX3KYKa1LqgfMjSIEtYde+49me
G9DgSFh9cHSBxq9rWLw8XmlpE4qtRHl2f3/FkDQibbEf6q4H1R8Ogipn4BMZABdy
5tjE5Hw7VgVdXPYVXUlo1/LlRsm7oenNBJA7DI6p5LdT5purpwbQ3khpBS33iD7o
g8W84Xyr96RvEO2w0RZQ0b2BqFsjJ2EUNfGOnryfZTzY2ay/bJXw4bASB8+4ZVgQ
5NscUzkHa6ZNcuz7Ryw8OS++eT3jMrJZAcmUz6hL42lucmAQNNSHGSVbyGk88RtW
5QiUWPIEkfkPzuJ4qdS7Ca5rsnUyfqkD0q/daLQfDTHvfXSyZ/s4Ho2pACa0wol5
mg15GxxtKFNU7/18DckSJwtFVW4GrofXkhoSrky/vBW8msGgWuMT9RmMfKLgotzf
e4vlfacduBjQaWUcEsmbIx5ngy3l+a498cF6TRKGOsVohW1URmgUVEq+spaR5G6j
LjSslGSpypK4TiYd1atie8uLIPB9fabYrsbhvsSylq6sMWrsD0QIMTmMx6BaBGWD
S3vVIJ6tHjhVCJBUtwC7uouS77pnj41Uawng9wQEkW9gXnF56EzqLe9ox84fTZar
16SL2iElCgsV2LZUjisk5T+7giyBB9j3c09lK9XHqsdnwMCEqV2Zo6DbmoF2AOie
lB1tt2hl3IAALcs1vTvHD9kBjZEbtr5l3qc34zScxaGB7LDTR+FHLAJWOWTDOP+6
eCXO9kzM8MkAGwA0NGXArd+V7NvMyCBbxz2xQxHsHHSgsuW1gR1/d3zbWMnd76i+
rHpkJl2haB655UvN9A2udQjLst8lzzfkqXpsLip9N2II9cTEDI4JaDWOpDZux8Aw
zFhGS+o1wiOzFOs1K6+/vM3iWvyP2gALHu2UwOkIhKeFRJD44hvpnLAzRFU6LfOI
nNJJBODSiW7sR//E04JRjyA7EetPH6cjWF2Bc6NnCIoOGOEM980aKnCdGmSq/J1V
g9DF6xp9lBSOPcGFG2IJqVVxOjHtRP+PReMYog47jyvdEy6I/Ydk7oZ2U88Ofgic
Io5F9X5V1/jR9oHZanmvx9r5yJPMCnj66IeMuRdvCkTrQKYSTtqfO4BLK+6+Tl2y
kKH87tVyC3C4+sLeVPoYF/8L4jVYPTeo+SnmbqB6leU3Ci15C0tcWhEeniQNWbCI
Mno+NBMzCgRVvmz8l1TgAxXNoCjO5D/IGRnWuRbqJMz9ka7N08oraZWj5xamsi0n
XaBTvFW4/f1TRwTGCmndFRc1jlVOzILV9Tfac8C56tfRWDtEsT1NlJMzDwcPNQ++
RigPFlSRDyX+EuCyjpFKGgCEiDQQNDds2MxBnK5XOT4HXaBIhu1zi/NcFDGPh94r
auujPqD6zCm79B8HQYOGQCUGdZ497FVP80Jrupbzv0dwRQO41Rl5RyODDXle/wTi
Pj0+FdmAx8nQCuEte0AcdoWeJHHlJsoveaLHOPusjpKNn9DfnUooGxU3sm38+fLu
ejc/I++nXwfJHXXEfroxRQ0WMII9VJL9Qc/ZxZPsn+JRenUa3d/u/Qd3nBokMBga
uledA2+U3TIZG6FbllCjlrwyo63ogKGOdM7KYRjMxeK3VYQW+pKZLIvReMkb+RNg
/x0hcp/aRIRV0q1pqNq3vv2sMKO+HBq4p1ZtimbQsXrUDWp1R/WTYAllhQ0S5wBN
yOeaAZgGjqwN6bvJqNjyLlZnbUm+UqhoMcM5CPAg3w3GsdH6HfyHNFUQAj136lMh
Be+cmeVNRRfl6F3CVL4AeR8ZvgwHRFsuQJznWM/QfEMhn7mSJMDkGUMcMgTQmL14
z/tTXOF0JEIHbQ4X4eCm9C53V+PyybqUrFBYw9tm2XOZ6Ra3nwYKh/xwwtLX/kDc
KDR5PjOKHZTeTQvwnLWnnarBzJKZBKFSrdtAV3dYYJOHa8kIQZ/Zu506el6PHcmE
6UYEaM6h6sBf6cwTsheec0KsFrn78VOD5WEG3ZCfzH/L8NrvrwJ18uckLEVuFLZO
AJS0qhPl8vjxm9ssrtCcRaBeLMPdL1PdPAbjl2hpi0qkZYZNAuYSNF/0wo/ijsLJ
1+DOsSwy6L4vFR+joqt0uoVBN3qHQJlZSEfkVn5fUlYlDQAYqieR4KTGV96Qxd/B
mRi8A021MvaPdIVSwkYfDE6V9BbP38J5qy6b1Ft0dmAAYSUY4GleitlT6MYNVtsH
XlSJ5/NXvAv9BUvQJddd7YoiZYX066Go5GNLA18zdx4fD40n61Zu4HwrGWV41lmf
9nau6ThfHvtcCIlVsozdqCTvfasu1Vgu7RjNUm6BFK/QT1NUZKHGZwn+1ojIxEZK
+7CRyyjc4tQux7g3nx3bJocuoHpWHWkkF+87m6JUzwjIGMhsNkGTNbeWE71jPTgb
OJ0aLfT4rpRUwzMygDHWLAxg3bXqx+bv1eM1+ZN7SqrhyegVw61RJ7lhG6lsk1kp
Gx1PRipoBRDNFNq356z3+BsZRBv9qfhdYd7Q64nt7gYsjiX/51SGLISLP1q4EDIC
lRLvZ5gejY48rVNsmKsM1Lc+Ch0V7yCufgD5bgfgyc2oY4r+WRqUZaApBR/8ln7L
gzRDV9WgjhtXjVEHITVn6GXWQhC/g+GhIy15+1A6WYb5MfhvKmWV46erp+qbG2cG
rYv3B9crN7xHHMX+wh59JzK0jA3Xr1EhRI2X0MyvWKiB2VRCNIr5E+/qgH1PWMH1
MLWXOIstbykF8oKY+Y7CrabXr0um5u/zRlD2gur2e0JLzrjZDaiGQF5aLruonUOJ
xEfcvvLDib71u+FDZ9ePElsPfXll9ho5t1BINy2Nx5BtlyEFkt2qJbf5W3ujk0qb
ybxDTlZREsmv7RB0K9toKEfdW309tswdLKfSot108+MhRlGOuj3r6vvTu+GJTeZw
WFkGjYNyo153Wz7hrBe1J6wbWccHLgScHvlXloKjjJPNz6LE3igbVMWBHqTfqa6V
tzX/ygvqoxLucuXOypsmC77Ra1i5iylEzGcI4Z3+HGTwkbzpOj/cOJOaAbaBHySc
lcaCgB5mXbXzcObDNVXy5IFv0lRSah1aIDlhL07z0O62qBrdolKhfmhhJPvlz9rk
o2Ag+2WuLcL1IBQA677PLb/eA8hsPZU6XzvsulVDXBmn5p8a70N7TJQ7TJ87qgHa
vC3brOTxlGWkaOTiuQaqSIHatmBkJUJpks6l1lVjY+DQpDiblFaCLmW/F3xvc5gb
nWDZIMZalbD+k7q/9757gEivacQqdx8lw2IOsHS9i/z28nb6cLu28RHkpOGp4jWD
m+btyNhwy6WCCxrPx/v07wtjXS5ULXzxnHiTWn2+2edYvYRO9z4V6X83igYQg5Jh
aUyeAnZC0yWhA2A9DWdGb0r5q9G0kAPwUM1gGaZDEM38Rl7GXlEPXZ0Fzx8OdXpr
DMKpfCpGQBPY0SatIuZushJ27lfRKAWeuPYeAPiK+0gFS8i0xlIVTw2Jv3OcFHPW
qPaYUb2vQrolg9lD1CrGseFMUun9o235XJN0LCTETI8LJKXqSwQ5RMA6ZT+Hy7V/
n9QFZjg5zhqidUFBASroXC2fl+der0RyOChFUE5vNo0Z7jYduLJvQlqdTepag6Mb
eUo2zVhoXXe0dc+0FFiPKoX+4gpaLGraAVHC6yKnFTv0cfNkKg95n1stP98BiP2U
2k4+RgzRmbqjDUgPS9hKrCQcdMbRvWCcH5c4y2hhfor4DB9eInblVQBNzCmt9LzK
Yx/e7H/lBNpiJE0nRYiSJg0is2s1CiZUZqlsNCm9Ld4+5dF4F3HKMcY2UEI/wA/T
hkmVtfSWh7+3TWBEWM09kVas+Ws7FG+QGehX1GWjVEBoUemo/jbg003YDg6W+cqa
FijsRXh3/uJ5cJXW7D+A8ZqTvnSJQ3fq7Jx/QVqk9i+h2LmSmdpnkJIm5gUiiAro
2+2uWyHzaOz6GHwSK9R42GyLzkaH5MGE5z15DQ0SeizXefhenm5GhYNH0XuQxKCs
zT60aH/Uf3tDrtEC6hFSMrqKnmVDSRhG6EgjVgDWBV8DDx+SrMBusKcYktaIZs9d
7hGadZJr5yzROX1B+X2mnkrRxjH7n9D3qYBTBwb/ktoFR6VXl5v6wWNjqMKIy9N+
K5ZiLzNxw/sKqkYc8wZqViI93uNuijNRCk2LostoUukOgEuIv0Q+/KCpFAYjIayt
SV0OLBmEigrBt4c66OqX7wzJxCM2DlJNBKZvpaTLr0pT2XfBLoE2adiamnIXtbgn
EAnStZSIF6VSUy1z31UrYxgYHQilNkvJSRd9wMwbgO9SR5HewZRQjYJgVZDHdE9x
u2ZA/l7C5llZ9x7Ro88oIN7x2uxU11g16zN9k6EBsXM2mn+mzp+Pwa9OxONLoq0l
GZ6gVqu7+T/Z9KRNkEHfVvmy394880WJQTluog+MF5L/bhvmkHquV2V47Bq/iNWm
FMdASYBK3xHn/LpDoDdwM5435vYSpxqGfryfJTSR15MJPr7MDLwBfKPtJhGbtxte
tLvmo2GzK2HsmHe/iGMZMRxYtxcmobxzlogzRuBuoAjrT2RP0v1ys1OSWZKIkThf
PPp00cDK2wxpCPCA389Z8FNYCGSgxzFvtN019nQxE9PfKEXAQV58lVa5bkdfpo79
GX4UiKxXfFeXr5eyJJ7hoAJJST626yZoTkLuHEnnjfqt0lEeGYFZC/3cIHy4I4fp
`protect END_PROTECTED
