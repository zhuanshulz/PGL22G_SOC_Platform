`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vd2dVIuOoJ3U9HtqMV1OxZ1hiOBOEbCc4XSSKguWCa3qkBLDWI7i+Vi+bkFBF+J4
qU0Y/TQyNFaEaIYpZt9UYcAGEjRJe78Iv2yZMsxvytHo5pWkuE9NmDvaCBzm7jPk
ig6QQGrYWGlTfawjZyDghVSP9CQ0BwtJGygebxvo689PdMTABOY1GKJATZTxkGDl
gA2VE6YVG2NdQkL/lsXRGa1mHGcMZyHU+Fm9fbi+u1JFPnHNTOxh1f7tF6VhGR0j
UHdMFFxFOyYXeZYuwfVhDB/zW6sHQXQYR7K5wsGfW1+yPxo4GJRK0qVDHq3H/7T1
DhVcsKSZefDrXKyPnzfVs1LdhAojrIRDkDjDFD314qWYaOAMilrM+XdAEzj8RPY3
6Bk/c0e5rG3MFoDEuvOMFtiNB0nHdsqzMzEVloMXL4NvNOHWokA0KQXLqellOfSP
OsadZkfwKyNCTKnsXrr/VOtjUUs5hmYVQzyb0A8lF6tPKxY2FerWD8GZxnEzSuKi
7t0iIYPP8S9a8a4g98mJk2qxkVL6ie5JcltpGhgnGRvySouSxBIKpH3Yo8BFFzsy
BM+fShKqAOp/7PcQ2L/IaPPqdaHp/G+JLwfwM7jQLoEMWCnLnm7Y+wkLlHWyF5Qy
+N4Ki+3JxphlT+LAc2woE6ILHTYsHxUfZI2/ATp/Oc/dfH9bawDirrCkb2sjShl7
H7tabw9yJH8Mb3B6zisVSkkZaQkWhT07H6RV5I04whmv+aB05mrKZqQqD6IKlv6p
vDS3CjqBx2yuAc8/2okAJJzdCOdU++ID7UQ+k20vpcNswl0n1XiUPfe91RQ3wdYw
H/gt/944eqHfOnXavcsAegf9d/oLx/Ar3g6wCkSms32QhhBgu/+8g2IkWaxHUYZU
mkMPV29M277e4PugiMD8G/t7mK7TkUkYw6EejUJtwRvfzmPWzwQmg1+nROjqBibW
dziEUdn6Uq/I+qgA0PFbJZWuQEBvGE9d1BobAbk9VYoTjq6bFoZKCl+dlyh2XpiH
qJu493ClvawRaOKKyMnu2h7T0zzQPNdTdwB9SDc+u7ryABCdpNzEJAYUV0bqXOzJ
hwDvca1PuN/etsYY1t9EkxVlwHry1Meb/FXUEZC21jtzlX+NRI6pEA1kSzESbSbW
0VSXCMmuJ8YiVgkyIlwDnii2SuURxFeYZen0GhreFsysvFUgKiy6sCJzlT/x4wSc
99QajN9eLGNXRzCvBohejrf82Otd4821yU9r9QHIuETECE+6WZfDgV3CS6cPIF4b
+5ITVNrJUA+cW+OD1nsg3/SN/tWLQqDbSkgOcWQnxNIfeH/5P3/IkdAnmNnXZZLz
HKbUC8oJ8hZRPCZUtiMSQw==
`protect END_PROTECTED
