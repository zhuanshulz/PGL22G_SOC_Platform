`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WajzYungcMQuvBGfxoY2JbZl4kT4c9tKdJxxdOKiBQuvB0QMjqe+L8piCwWC3s8r
MBGfsX9dCzyBUpIC2tNEM28gS/A5QAYmNoBbmy6QOYlZhFsOczW4m3jdfBWfec5Y
foAATtqq4hCn5jyD7WT3IXItjIDy7v1etPBAfnJFg+kB9J+MKGmBMFv9ovpZs6j/
RWW1uXYHAPyqq9dne1B5EgFTkupPMPsz3xzxqd24mae+A0IguAoC9Q3QK+B4dtRm
H6c6mIZnbXshIlMvdzwFZCaPL1JT5me2WvrmvEEOjHED0C3zcABLttJwHVZrpHsA
/+3OHfpd2QpIYkI6yN4P+9ixGXB0DFZvYm//kON1cGlDFzJ3aGsF0XCip6hiqIJu
JFK4qcczWDQ850MJHClm7Vw2Eg3ZTiPGrPu2uFVt8Hdgw8RsTBBzap6dVGwkGqmZ
XgOsBscKV6IaUnpgq0UEHJ4ucAvyIkUhGYODE5Bp/Ld2DTzplKO2Du87/jzlrRUN
l7qXLtlq+78smMkSv6W0WiOJlQKkpMZRmhI3HK8o3zQeszBv7wqUtzs7+yX7WJYx
W9p0HlijNTqchnobQPxtIlUWBTm5pqyCP6eAQJJQ2czC1E2LrXckRhNWwK+ukHFI
Z5HfzWRVgPkY6OzZEd31NyfxSV+8IxJlkGlZqODp867EtsPNR+yfP2MzRHa/rnEl
MhxcVhHHLDN3UbnOcgGxnYJIW6tMmzkRUD4Q54mooGKtf1ESZ62uwa/JMWIeRXKs
7eeqPsJ5YW3iPIhIgWMS+tm7DlZfMJFgWV3rnigzJxhu/1q1OWC5LqiKBUvIxw21
xSj7fVYfktQygu1CkmlhNS3CI3fRtouz4K/1xpi9GdykWm+p6cJmGazyuaOUTpaB
V87W+aEzI8hE/CgAcdo5DoWmwCt97fvVHvI5MrUu4I4I5ewBmx7a42M1pkbZa8K7
BdZRUTemFsvRIsE89RYSIElWU2afaJlyayKxkXU4S5lgC/nMY+8HK9CwD1GZv3c9
baa9Tqz4TJUfUn9aznXPfKE6cUNa+qh4nX0t3Y9IK3SsMQBNc7zt66noBR9ZVf1A
H/rTdr0V+ap7nrVxwz7UhT2zpkm86xs2/87AwXH3A97226jduBpv82OFw+uowTFj
aibsvrvFzgdDzGAbUSGw50076wEEu/HgGoi06dmTtiZugua7HiCuHyWyzpJHz1rD
bMleuPxHojNhoS3wLHWUcr20ifCD6skVQsxBUn4AZPOvURQUxGeOGZWLUeSj2q59
43/smRpPxBzYDt718wKzCURrbLcGnfo/1PWJFrdeHkR0iAMlnCXcdz6OeiUpyeL0
uaD7D50abwxRoadkxmqU3fsGz+67ZFoH+8Hc8cbHCgN7mm/lBTH+WZ+RmiN2vh+Q
KFfpYmRpye8v0p3WLCoNuk4ElAfNOc1FMgtF9TblmlZyWFjjKQzCcokUftUY/CiS
Tb4pd3CTeQFmmJ/egObm5OecVSa3v/IeZPUA3Df0voVViLt/YNeREUKx3dhioU3z
xlqEwiN50H4gylAa8/GhogaWLKLvt8EfcugJ2pSO2dwnzyvk09il730UGU1410Ux
N9WMEbAimXrG1/OriJyw0tjk6qiKzd8kpK0vsLpBfpqYY/DLfMZx315ijXe9y+vj
Sk8Uc0jV58yb/nOffPN7p58LNDr/SrkvbNz96zZSPiHcUvre3FVedAR4HNIOCrJa
XsVglamTSwWmj/DuA1N+dgIRgBrpn0DNey8bVDnE3++gYi5E75I2QujyiKseLfCt
BWjye/dK8Eyzs2i/X3sCPHI/+7wRceHroXEoyGqK16urpZMDbIWQlN1955pLoaSK
lvBqyurrjlFX5XB2ssipRDjt7Gw3eqfb3fS1TvKqdwAZ+u8tLItkB4+C4H4k7AQ6
FHbtCyCvPMzpCECmlM45+8AJ/kEjV1fZyvK+Ic6wdqgVRJ5/s1WVXgDqQNYJdDGL
tFVtQyjiPT0m6r84g2UpsqIkptmLIKoe+asXV0D3K6d/eauu4dUbmO9NnBpAuYOI
uZ1pOySfn9OCBu8pB0F3us+egK2h31qQs/wHSMzzuBKvKHjcmP/SBVvxoKDtAk5W
YZUZwc99bkI9jlf74dZVUcyhkH79sgveOiFWuQ1cgUGPrlDSSP42vTSePYJqY9kj
dlfNKH0DmlJFbYXfsfGkVrwq2H17kwZrrF/YpHyaj1ylwusOBxjpyhI58S86ggv+
GHWGF1k6ycIBj4X8S6V6EbIkJjp6jNE4XqlFxCrBK+RJOkzr/r1XS+jxYcNwqWig
e+6dYez9R4fD2JEfVmp02RFtsT9o2qNuTLCEUkx66OpsLKRexyaJutvR9l/GmHju
kiH4MgE7qIWIa5zFY6E4W0q7CWzX6rM7bWKcmMeSDOpr8Y4T7O3EysRGfZIImyCv
F8HCSpV3bT9R5reyPAgo2y2F2l8i7wl0ay1RzTQtjnxLUwW1fAElG7yeA6Z9YoKN
lCcvRwNLvEFNPWps5Z2AHodKNVRFr4tUq95e/FrXRAU+hFXi7AKAqL1yBHkO4HTa
7tgFME4n5IqxZEE7JqD8EPt2Yl3T1LCNHxxZ1XAqv6DTWBpdXe+2hFgW2l3p2kRm
iDxnpBxdWdhfHNRjixWYUMvr7i5RqJ6oJcKlAlSCBCtTP/BKVFnIj0Q1bxVIJDcX
jZKBkAjWJguDwPs4KzNufNXgvNhSZ10k82nzt0vlPT3KFvoy4No2+zKzh+uNMIeT
a/UcXNih4RyKJ1PEDf5E3ehUweXaKjvr5PNj734YFIfmfyuVCnP0bLG6h2ujgPAY
QVvreX7t0I/aKYBAAYtZUdetDxWP/974ANcBytnBRLrDr2x8bLz3T7mBCSXAAhQw
h6FvrfzzfjcEKMiiQNvrLAwNgn63yQJ4EL1WVjpLV+cIyMXHn90TCax4JK2FEgMW
6i+dwpkGH3fhqZYbATrdan1yh3EZ5ulPy5N21P7Hx+IIT2MW+LQeI58sC4bMq9Rv
2yS8QNAB+GHWypofZo7hDTtYxnUMAL02JIoY1eTpTPN45ykTwEi9bC6GyjEHzf1K
RaeBqA6pAAO8/WbEhdDsJMZ9RAYqikIt0GMA0yQIUQ0nlhK7XuhZ+s6BZfGkH+Aj
lguFXEdyw1aJLznCL3xyqg2ZPMYsEWnxb/ORsOjNZB58Q3yqHg9oG+gBRfmeoXIp
gNYYLUmSGPmK6rki5/xk8P7lbbFQkfI2MKoSxZdnOOSTpvRp+ChvhRNj9h/pQ9Sl
PxFmVmDpQVXMNi43YEQenyvd/hIP215TUfLh8eTC7AfYo/UvPs3e4xC6nih2di1n
kNnQZgiI/csCApKT0iZBfwH2pXTWVgyYNnI867VMpoiopUgHFS/W0q8oEqePQB2i
qRjnEJ9F+x3GGjqXrBaAVhUFfUxfm2dAcOE/Hgh/oAajtfIoFc6W1RraODIsFg+N
tH0HsvYTmq5hxqWJMaveTFuPqsWewiP5C1tfwsorrqAN5opZEsd31IwG94Nmw1q+
ncVL1cTNHWv+eGl94I9HWBBIR7H9g3VzHwQq97YfNhKHGj/UieiRKKoX0W4nb+zP
OhjF7een/6SjwcnVorcM/5azd+qjhdR+l0aPh4dsag0oU9YCeMm45zQPTxUaQP9g
9tLA6IxUL5LB86jdgz6tFl/hfjnLXX+7b8QwONBO1Gy+wIC/DJC1lFpz4CHHVVRG
dufpUbFFqooL+2tOOM16f81mLQkR7FItKkVggwkBCj6RuLqiU6+SYGbKEvY9AG+z
z8EdV5bXb43Cgr/LJgHBE8fGMi/XoNRKNqTnxVRhO/LvTdRM6HwQ3SLTBe9vuDyP
PGlgEqhru8d3t66qmdE3K3SFPJRs51noObTICddCmaCOR+DD28NdjofbIHCYyJmS
zgvmafhf6G4cnmKZ0V19lrl1O9I4VIXle+ZhFpUiqoPujuUKrnexODMv8D8ZoxU1
KfFgY5eBUlvk61ZdQfIl+5gjdWTrw6kFaIfEHhD0GWy5BQs81Wa68c+XZB/58jAD
AkbDdSI0jINZ/bZY++7B2hIYlE3zYLFrxTunOlhnpX27mFySYpKGoeaiubBFzHSB
9z6pI5mW+drqHkA8Nti6fZqHOfhxwBGaBtTTGluly/irqyJ7w8rHi93We1qSFlFo
Y9aRnvqmJr3VOkI6NHGM4cnjKIS+TjCixrcaVDpmpialTUumRsrhNU/UahwnPPyo
CeMjE8Q5zolCUOJNKCr/iQqrOz72bZ2VAl/yHk6Mj067tsKetfE8Ivk+0ZNPOJ73
ThldecUpK0USxip/bOaurTf73Hx9LKMFQvrrAlbTHEBHwxPW+nNc88CZQPx4C9TD
t9QRYrqeNbXApqoqE598+4KuSzmQ0YI1J5CtUvI9b8UqqoYhya+LDi4qMiXc7GHf
6pC23AeXaN70UoXlxSQX4E4x+7wHn8CxULlD/fCydMKnys1nbHtS6wtTbXzQJiLB
Mncw5kL8kh+Kc2K8TISmAuUGS6zpxvq35UT0Ae/cC3+eWWpPX85lkAEh7FgCHiJO
`protect END_PROTECTED
