`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EkETG5Lthcni8QojyvJ+VabnGD6CoIPO10UbHoZDNiFPaZjhW/xVTm/Xz+UW+kSc
vFF60Wb7rkivCgix6fYPjoXEOeWh71J9TOGvWrgcxl5pcItW3t978NMYCGp+dJVj
dx7/alv67XEvZC5FshiOe2lpVkuKbpD9I/AtTZYoyQz5ucrf0cWUkyB3fYL6hGaP
Hgd6E8BNrwTvJHXpmLNtWw1I8/hFHtWUm39sUrIa/nycn6YdyOJBi3hHeCD/MhiX
U4nL1wnhWM6L5oG6PAsuPSEPgmO2NxqBv8UaJ2KBslU=
`protect END_PROTECTED
