`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BS6tUAy5l3Ioai1eS74wNw6+B4ifltL4RnbVpSBQcTHyepDLA2uLDvelwrMYZNgZ
ewgBRY6u3dXtShapwAj/+tozgtXRF+e8VOokBkiEqMOZjq3mibZ/JKFeQ0t8aq0O
3mxr8ipVxrN6PbRWtWquMf8rS4iGh0ahyFM6ZDZ9STZjKNj5iFSGtmwPcjF6ll3G
MpEUA2/a8m40LPr4kkQy+L69Pyc4kKS0mWv+NdzvpfVOcWEEn2Yu+u21E/S0R3rg
V+GmPBltpKGNM6RfP1g6b6q4WmzN7tlFesNICPHkZXkTWWqLPtvN09Sg4a2ZefQ7
7/tTQPLowFR2ejXwBER6rTgXgZz4cttfVfB3chMjfjE8SiAHZN7H7OFF39lql2K2
DQ0y+xfQ71fmyztzwszRkYXjG20fkszEIF5RoHXG/QyIaNEeOgrV/WECye8v09wB
ZZpEAfa0Tein19qFuf2Ynd9sINPfxFMfNytw0jrdFlilv+exzS4pgVE65D3QhZX2
9o9E29GwvDdH5ipBKkUTUJiMGKIUUzANaGd7sMNWVJhZ0wiv65kS7Or0e0KS/Fsg
gkHD1YVFpWLDFt3qBhL8vS1RJwEGpqvnoxUCyQXhABkkYSJa6Z8iVjJU0jvXZhFz
hN2p2YCSMP21+3ge31V8RelyiAOa4nd6QBahB+HTzujdlS22gVuA0LfzrGaiRflg
5B6KSNZG0SzwUGQ9RguBYc8XwKZ4ISS31B0J38uIU42Af6uU5plSMJyNaVypcg9e
4d4fAYty3AwbgDlFpX56I7++Y6yT1rGJUXGzWQOR67Mu716UEoY7ddY+TmUaT4K5
CrEP8RHdMA2t9K0ae5UuDyHkRQ/hyTONLxDImHyvpnIxeb/IiPB0NLJ8/1YXehYN
lZtjF0U/hs7CRywIvrqO03kTeGKRtVHNa9B1JmIqJRBqinXhrXmLrqZQvkeDPUZw
Dh8LVO0WGXLu+7/DV/vQ5w==
`protect END_PROTECTED
