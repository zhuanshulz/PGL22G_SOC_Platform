`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SET/OqfypcaqwDq53dZ/Ti8J8p4mufjTcoGcoB2U22chEyipk616s+6UoWU2/RuT
4R6gK7CWuLiapj4YJvFypBGgFqLF2MeMGSlOnoY4g/cd1VfDPEft4bPmWtSp2v7s
WyuN13mtZDbabhD3PfynrCZYcxylwgh3uq0T7TvF72zW7OSexDhmAUZXzDtZ2Zfp
wko/DV/91cDOo0csCysf54PGEt4t6itfpJEmmcXDEsb2fJn0iX9N0BiCAW+7gs7m
EjbAAqsbaVa74bArjPMZmEJsPvuDlTewEZtuavnhMSH2+Pyd5KTdREtdyefPhRDZ
ta0D6vugDTTpS9g/vhWGaUWtoeLaWKRxRhzArvBFRcgZHuPRvmvXoye6pRaqSA/J
b6xaDvYCKPioV7iOmoGyACu7MtE1NzugyisqR0V+rqrtZyxHml1g0dcL1cf8oRHl
qqIux4OUzpspBxMBnGj27CdDP1mLARsDZZE6VOWUKjp5/2pPU330jZrDUKc9OCBY
TXgGutbgrGpBW02q2XrndtBhmfRQ8TgDJAVu9VAMD8zd4Dcly0QfiBlsK3pqcIhB
0Cj281moN8tggERR6q5t8mFbyDKPIL4U68E0jd0Len6xqhKD5VQKOaa9jzShsUTP
PGPbAPrhsBuxyCr36LB43Q9by4GIBFgmagcIAghNnSNsZDSWoL8j9zw152coJ6k3
V1DZ1R3lZMccEXgtHH/Y2uQmImRB5Pt5Cv/KMw8FxGVnEaWK5Xp9qDLYICZe7SDK
RyeRvp6JqvBR3gsGMA0K7475XN8K3di8EZiHlGKbpu+Ff4l34B5+XWGq59kLTIKy
dq7Im8gT7uL97WsY2Fh5GAlaVooHsvM5UHxqm1gR44i1RdgSa2Vw6cWDsVBezoUy
XCpmD/5OTuRza2mtKiVeMzqw9U0M65zKYBC8lXliL1U6hEZ5krL8eI6DI4ZDsg6O
E4kIj9EoaAgiEPAFDlmxtdv4WW1CFRvFbk4RBOifnns0OON92d7hspkK/Y1ipcsG
9ONN6B3ePArHeB56NCt9Is8Ns1FmSLHXbOt6/5VMIaBdluJ7F4P0mlANIhYUzXJd
hrwtMWeBAl/ca2Pe2UA6Y6r52PGOzxCO6ePzSLOr57PMZnDpu5QydOnF5+gMARl1
wI+MRXDeQbqYLDk6w2NBc4SlYCt+7BaUumAZGCE/Kl96VjM3UjHJ70sJE68rLG60
4PkT1EQHo34l2YJ2aCLjz4849lfPkxg61nFE2L6Mg/HD3zxA+roWgtcYg5W3NCPz
F7ea8Jkj77Ac8KA6l+LK3N3CJ3esc89Xzb31GdCTb7Y6OiRv8vmgchbFTOiiSgyG
UqALe0fht2p7ZvLyEW+312QVc5oqGcgedsBa4jTGqlTDV1AeRmhZnv2Ro07pVu2O
q7F+EI4GwXcUzDWCIfpmsgNW5MA6mWwYikM02kmpjpgsWICEPIoE0qqLX7DU2rJr
WAZQOLGO7dQ45BqKDXz8Ztd7W/QOEG0Q4gj3eUA8yLWWINJObIyj89yKHhFKc7Dp
/j7U4wN7XhaVP6WKaR0xhxXDcWuVlL6q8o3sKETMThmW6VB6yvzvSYk1DTHZdJuW
yAoU6tM/3beiPNg4z9fp3JiBb1pmWvpHFoxB3es8j0Gcr0lywEaxSrsliw1X2QEV
UmHgGuSunBuI6KbuJ4HsH/sUlNpuHVmYmrWi0tgqxSJg2cBgBGm6JJNlVKARQwmV
ceEE9HX7Wvdrg4PR5NVhBlqnLcTiBvHJdfFf5AN0oGylkdD3zJnyxlKZX6bC2PJ4
pR4DJLA0EWiWh2aeYF1lGWUergDugBgja7Uxo9RYfV5dO3EACbERynXzVglOnA3Y
3cIUQWpyBW8sqdFH+jdOh2VJwcDsi9qHrlgMsifWhRAvapZ59As9j+boBJwjL+GB
IK3jeqeKVg8/g+QLm3ilJ/BGZFQoABxeK9OGLIKJf+vzspchY67jfupy0KRReWuc
bx9EsYc5iZ/O38BCY1LD/T68lSoBOYo/DaP073XeDayaBhRfv7lW+qs5N2wBo0E5
L4wTy4He6YvW1bLNBIkiisYKdHwC87VK8vNf3i8CBW1rDAmU2cF/qJpOl7Yb/ABZ
JYnw+evVKcDBs9VKGjxkgLFY0LldvZXXbtY3Ow9YYze7j6k6sdfi+Au3kcnuoSMU
fQCMdo5xaYU1oQQy6jrW5hiDYzN4yLSdRMt+aeOvsE5vqzqr+AIvSUpr1nPSKhwx
t7D6Be7+n8xx+QOF1stewEM5Os0k9ZAWdVwrOrO6aC6rNzLsNYzkQVShMeEekk8A
gqYpBTkeTMc9gn5jAb/mCZW0aoHKaNpcDW9+7LmL+0WAZBVLECXrRkHKtN97Mijw
8Ja9L/2DK/lBhp464nwPNqTnMuiXmVCrB/Bc9q3p8uTDGBkTFM+IR47XI23LxB49
Rc3PjtF5z/YSNYqyrWF2qQQ6ghgVi6NVqoLnR2nf2kobjMYsOdFLVqBhVUJOpXWY
orjLoVQYbDnoISjOzQ4SxqFyBuwQ+ZRU6Gc7DwHrmJk/D4uSC3w2sncGUWBMJBZD
JLm/ftzoTqN5woqe7JleS4WWlEOA+vfDE7O2Geh2QgH1XtbnsXWg9VNsz2WcdnNh
c0m20CiDKsxBu48GfPfpWqBTLxQjl39o/5FaPO5YIHLpTABI9RXwU3tBR2fTQIsd
JPYNNRhZvtEA5oU9y4Q9oJPC8KJCsrklh0VZh3qPeG6Mx1MhWTUCYQ+4IT8zL1SO
bG+pHecFDk4r5jcFLunjkoJ2kIAsB6+YsD5pbFfMVTKWH/sgloR9V4E2TWXAhJt1
rdzMmoNcsQuPF/MMmkr2d5hTJuZDKOBhOgDLGOqBRka+YceifB2CT5jjwJO1PYqC
iMQvh70UYCDbcRc/TWDv3lnLdjMwOlSV0Wwd3AT/qZE0dQz6v1Zshw1pAJcaw0fa
m17DSGkbmrafQs9xyXw7xbKzZA4EjLNXQEPJTF8I/LIL+cXmgctDaVRmPIGbPYiX
a6DFY+uX72FRq00KzYgwUUQD/eVOpNwxDBzUIpMbAl9u11tiNRXaJ+m0CMtfw5xz
/48yeId6XOU7DhLxMYfT6+j5Up/E+elvwrJ2AOsmrAhQTu9jqLurzbVZNtVBVDP2
Z6X9hgCIZkHwGx/gxqQoSCdQVuc0Rh6TS4HSMiREC5RpqJBwWKCs9fJyMr4dkFVp
PSeXrmuWYk+DKPlVGrYP2gn4BDXn8/c6AMuKZsOsfu3EFvbNZctFN3Og/kX5SNK+
hqNNMkD/AVy6I/bwDzXiNNtCSMQwAnrAConwdv+uCVfdbOhES5fxhGIoodjzBqLG
OGf6sPi6dJubRH6QdE9q14mqC2xTlczn3CuZaV2vTtw2yuzX1aJ/XImRTvX/iMAm
tyXB5HiIxC59ospe7puhSIMorZb0cKPT0QTD/bKXc4P532YzQFSfa6I9bnuWhNjp
N1Llg/ppiK+d8vDwy7kfUd0uqF8i6aJee1sJS+chfb9Yp3DWiJj+j20omYNfE12V
izieEOuDEYrSiQVIhudmY/s2qlZg2X6LPH9Z8qxACRSb5QVd8OphFfb3Dx5zEqXw
xe0TIrQ4Kfd8A5/Yp1WrkiLXScQJjSccOodjoqC5U8Ep7IOl2hDJJUHOSm9702xg
efPE1iOH6dPigIutWl6uwyusJtWhLYz21dk6lXDEsmKe51Fz4RiC7fSuHi93hLlu
C2BY7THUCla4eDGVoHjpI2XOwPWxas/s8U8TLZxQG90AhRznVJe3hevonqHFlD+E
BW6hgBF8kzfDq+ErhPFRcw==
`protect END_PROTECTED
