`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
80S4aefddE6nLh2+jdWl4JoB2I7Ksyze3U4cZ+zGiilm+XmOeZHbbRWZ/cyQ49Vx
ffBz4u8Ni6BNmUOFrR6KbouguXSbOf97Hq87MqTtdWprdQF+OJ5zEafkAJcBn3sU
E3RHgD+AOiLlWr5wzAyc9E/NlaJYG/kehZViY6XYpoep2xXiy1O3shBw7FLFuEyd
vqVUdDGfpHHdJz44EWLOLD1bHbhR2S6NcjzC6BCwpdxJVozdAqV4VNGDItaCuDd3
yKmx9c7UucUg8BmFf3y8aA==
`protect END_PROTECTED
