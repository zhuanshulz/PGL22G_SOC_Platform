`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9iu1A+TTbwb8MgMEQGYsKjlX3Jc8htOZaf+vjmzJM5CEzbKdp2zGAFotFfWOwxg
LSYTWiVxnW+3PaRkZOI2dfax3/t+eSnCf0aET5RsAuWidwPTAy7f3yb57f8TzxkN
QejP2vuyO/UidFdGOuYySbpQutVTB5wqhrKkhIZDvkGuxMGuPHuGO0xp5pHdGZn+
5+UZ6M3NQVV9WESVG7+GJSkeMvZDcdUWuOtqq0I3vhxaY6pY4lvpIqjvUTFvclHg
J53nk0JygPifa8JH159bF6BeK6Zc84B8VEVE1a7JfWCodftn9z7GV6yMYjr6tE3B
D55Z/s47olqcbMSgtrJyPLRcwy+V0fYopDLGHPSZZUeQ+vYY+wmxCvI9BbnzoFDe
1xJJcsV2HiQIv6c5MJbjn9+nMwxnKpeHRYvkE6C+yeu2e6abcKo9ebWjsJ583yEM
zIN3ftH4oMRYxm+LO1GEq6om4PJTwgCx8XfS19zmVEUj2fgqizwFqbkhimghOcTj
MxBMFAVdoAic7FhoSpkx7++EGOkv1TDRiLNiqvxLVCM8GCOEsQ434stxp3zaUZSU
ej+zYDNU8wRFWr+GFTNy40YrORakyx4H5LI5ZHtAAmmjBB3l6GGJRLtm+gxifZW7
ZDGmvPfGjhsRRQOHL6r05nFJFDQ9oif7QamVCX27bH8jmSBnVsnk+nctV/pMXb74
guDEJprVirClZM8ZW5J5xh2iMUZRakUZ/GRia2OzdHEhX1P0zWRKETXdOP9j6wSu
+B6kSckvRvCkfq6ESkOJZzxW4JrlanN+lb6T8Q/1UmU=
`protect END_PROTECTED
