`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kyXHxAsLu2uej5JrHczD1DPNWzag/xDofxYWF7IQXjSMFsXK6u7gyqjnEU51eRQo
ronFegoBalo4tWYHRyaFafBmgAd1Ffwh3Obbf7qNbyFxrX7awaQdCkprwpfpHslD
xgV4WH+DJELPIsT5h5IQE/Y86SFDPBccs0iD5mneRmYoVk8NBeFnGh3B5PxJyc1X
E6AYLmB+7DbMrh6LbldM0JFE4+vMYGfzQ7fBcFjSZTz2yf8OkyYB7MZ9ZekBIuyJ
/9I825GYK4yKv76uAhmLJk73bbHZUFHunX/rKElFjDbrpp8dhMi8VxjD8kBvoR5f
iA2BnZJ5tkrZ04ePFxqmDt1ZW907kDn7ge73VOR2Hz2NeNqTOnaF7YtGZ5VE6NRZ
oFjO2ed24yXbLiF/slr4Jxml+jqrPAkzh8R019ymikC7KyAc2AbJJW+dD6SR9rFq
Ohq7r07vF513bfL5WrpzfKaYsj7+iNQqituQ5qi7ZSPUlNVFrOI47WgXXzTavYJ+
R/ta7ZdVg6EsUcp71gvPow==
`protect END_PROTECTED
