`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zkXwKt2t4zjR52blVzLN2rV275Lh8CmoKqqee1dSEhD2brIgDk/1MJH5WxVCIHc4
2XVLd8oTVULkGQ+GOTSc8SI9Pcl7jO+8KXwkLarBNMTkcCNaOnXY/hPBYFyptxeH
ZcBXGrwnYaeEEr28xEmtZawhPLgDv89QZYvN7pJmeJqxlmEMPffZMU6V0XWErzVA
VpWd1L2Hlmsif/7q+INM6QphZ/LliG05RKszAJGi5V/C4K5qm+NOWt9TIMzX6mkC
cW13ZMQ6HYXWRhjgR4E5JaFMx6n+UEB9qdYRFtIu8htu5kFd9lNJsujby57Si6N3
UNaXHfv+Y0UTXkREOK4HM8C1IWAwBSZjgOwxxusk4++Bnptmz1RC8BBxydTF+Ygm
PHZsL9J3+wgRDHApXW5vszOGsV2wtyiDWwll1SXQIn46mfCerbbzWXfxCLMG6kuD
jMVc7NeC4QGRYu0FqmpZa+k5MJ3JKuQSZXKXyfzY//Df+RsJxGHU2e7rTehB0FiD
Xo5DIWYF1mvMEjnb9kGSmq6NrRdhBg8LpANBiwKdi8AnU+HjtzdzW+6jH4MI/dsz
rgDZJ+MKT4LY9bOfaPvwJ5EjStO7u90ijZB4AcVdOO9LyzHSIZY2EByTEmqCqUu+
kNGgOiMHHnr3B/UUa1MOAjrLNR1ZglVFMgEzzNLOB6mqAkXXpKgtaCe3ynivrCn4
x+Qj0RYAsEH7ZYMwYb9TdTZPqlan5UvA9Jc2NgWjXVv7v04lo5BNM+4NgD7kjzUm
X2tZWcFdv7+vWKa/EpPTrLq1IkFsSYM8PBR99dE+WzPgkKrP+O+YY0m/n7DLE7im
17nFiZm6cc7X7h0A6CzW+VPJl8rVqN2w7U1DYHluGA6FE2Kw+34f7111hx8OGEnn
h/j8tlydTCSNGOfdmkSx1UjLrvow514lCxqTQFNEwyMBOZaEFNkvnImeCFg1DpUG
qpdpUkOqDCBanulGbGU/iJ8uB+Lg4YsEftJb8RVIgOPIOpS25h6Y1ncwIn7pHnjj
HT/sKN8dF2zJ/sCc4h2paL4StZUZtWyDhtgebJhpeWpwHzBFMNDyTxcLQjUWc/MC
dcvL1lzWxEn+NBEzZi2bsbG9hETNMThzRYczhDC1A8r51X7vFnLkRk0GMlLEBjZU
FBW2ElpxiZ4EHYAUAhjZj5m+rFLp07gnMW7KqT8z5p/P9FTKSFiDIMk2o0fJ8Rup
jlR8Pni2ukSn5C5XVj7Hxg==
`protect END_PROTECTED
