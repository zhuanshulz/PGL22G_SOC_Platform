`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/oZ3imMdD2qoAbZRBrAk8ei+dj2tkYc7JBBj7A8Jz582vBwl0A8uJA0KYn3G3r1Y
iMX0SUvvoS0Ut8Bz1VfhKtJN1mmChobe9bf5fPG/PkkfSqNZKLCLFIa/EeK1KT/l
8gaqfYLfDZ6yDB0Ghrem1omkDdPsc0mYbc8FC/riFq5hy1pRIErvrpWg8VHyNwmq
L5Qt1PKPvPNYcigSQ+OBngB/uzopImOhubfmBErANiq7sPif/8sqfrzutWeFEcyX
r+tRd1ORWQM+8UhhLk4poxf7clgIehPTF1Xqb0z/skZ6g+ha8YXBb9My/corlA2v
oJqxJrCXbnqGC4FTQUQQSWk6FE+244wB2P5PWusBZGwTEopPIoSURwpsu8K+1FYE
Pd32vvRn1R5YrWeK40/98hk94EO8LU7dAnLXuTh4sE43kwDXSa9L2ozoglmo1mHT
m+/dJobCbJWpRIWVlycaIaJLU63gXsX5VHVtOn30GHDuqpVwg8Fc4zeEPPlrBvrt
tLUJmuC1C4hj1LTmP4A6nBD5X1xgX4DIlhTUPsFj5q/QcGXLtaSK9Y78b8Iqrsrb
VHmM3frFtd2c7hFCjYh0XHgPF0WzjM4WTwr1eSRdFxIkeLoyI2yPpzUhCiN0W+V2
RWcpLoIekI3mtMyZ2SShW7AvkTVu6SFkn2rgg6ndsQahX9O0ngsROv/quInrwUAP
LPfNofiStnDG7Cx+xFOvlcGjR1GD6i1meOod1NUUWSQObHjkdi/ltAycbam7AWB5
OC7F+cuW/90J4ynSrQiZLy0VK7ZnRrUJu6GT8ljuMN5cuMLiO40dZr6efNHVgK2Z
b/yGotlj9QcDz8LK2FoQ7d6z0xIGmPKCAProVCs2b4xUSEWtpSSfokuTUVfV2J4Q
UPCtmUZQRM98+qx3rIGajinn9zWbMn3UDvsMtD26Zf9Frnr7toWmuT4hPA3l2Rzj
8nttLTbrIgKKvJqXk7fSWw==
`protect END_PROTECTED
