`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rAr29eRtqS/mw69ddPwWe8hXBqaQYsq60DKzdb1UBwtq0COrzkikCpKz3XvjyWY
6c06xufVLSJ3gQClNA6zKihDoWwBS+p/ExPWMt72zJ84QHblkO/Yj/8R+LoCmy4d
UK/OpbswIyrusOSsWX2h4ggQIQmO7ufnNOMH8ukf9oYmNh3XeFD6Jtl/NNXe/lIU
uSXO1cj0GxnV4QcT6b5oNnKaTcpRsPtsSTEekfu8cG9NojSoSLmVlWgtPv1uC0mv
tJC8XHHg+b0NyZ3M7sA/DEVI52FW1H48RPw+OIQU05LyXlsMMoAAfBaFlyvsQtpX
xiVnPCh4KUJ7akuJBQ8WsWNShQCRvlbtCoihIn1lNRm/zCT0jVjMsW4J2M7Ggixv
V21qJlU9h8sCwXrhxyFVa0z0Dw+9Jc0aXWBWXaMQeaEkB5Ouf2WP6R/dvupj4PPj
UiA/iaX+8VNqotwsCe4YhGD7Eeaj0zGkkwuoBnlm3fyQXNTMh1R8CnlLO1p7Ciya
rTsF59TvDDITFg+GhIfJLQgNIrJFNmwENLSVHbbJkry2HvsAi9aOFV4bqQUqeOzF
Sih79n2iEnyatIyIXUXpkv0GqVDPt1Ft9D/lgn0dpCQrMKJ/EFhJmSGBOoMks2VA
nAboh9qyAvfhGQOX2hP5jVDPjRV/lHSigB2ru8+2h5FbWzgPlpGzm8b24NC7LmJJ
gCSWTvobfUUmUiRi+fBGOKqS/2qBw8/3WtqSdQIiwDl+aac1zFG8o8kr+frc9G96
Et1fk1cglsr274fyofkJaYXa6Ol1kRH6q09McRwPgj52s4onekus41WvazAW4dg7
Vch8I3xMbhwh3M5Ke7v6yC+fkT3ekO6PV/SEYOM7NpVaXj0JzH0c0eMEqWDO3Hn2
Oz6xEB0D8FD58t3RaA3UcQ==
`protect END_PROTECTED
