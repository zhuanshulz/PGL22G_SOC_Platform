`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2YVLKHkS1AhN6alItzMdAGKEx7szhNCpz5xJkwtMkUwCbu33R62h8qBHyinOXqP4
c3MwRlvItWopEJ14X1R7OtkZ0tjgTQiyej7fDo2fceiGzPbqejD41BF37c2dGML4
wDs0Qg9UGMi5cAWaT3fCVEaDtyKLKBgkIKlEOmUj+Sj8he5FdzaYi8OQRDaJ/tZ7
n5GbfohUs68jI81sfRK5kV8Y5tYkEqHdfSlxiPMfGm4LoerOcrr2XXT0deBKle8t
W3u9yvOP+05f+Vg9hu6NFLPONcvd4tl3dkUqQlAOQUmefBlnpKN879GFOp52FM5Q
WWtSOob/rUJNQ4vVrw6zEf8auCmE/b+5nOjmdITKHAhd2qHM9d7ylNBwE84g/+Gh
OEW6bK6Ow+gIGs+hrhAbuFlrXPQh+RbjNlXJhYancD97NbcH1a6nGg9T5qy5hSSX
hySDV/k5Zf3NstgZsktS2DNDIrUqrL/JLOcjDlCUtN+GGGuBLdRCtCFPQu5WIr7B
VxsvRUlqcoepdWk5fIL84nrf8VpvDEF9OqW/Xiu3nXUj0GlP+gN6KtyRPbMU4/NV
QL3Df0ZZ56eYkYdmcUG0caFaLJ9SEO3l+H9gfZcOOZFTaYk5PRhhoOyWvc7rcFGO
F5GSxDQpaI+KBYJlQZdy6atUE3aerswo5h3aG3jXjng/v508Tqsg6UWCdhj5CanN
1a3DqjskyI/kRIoXMamyl8md6JJL0LT+el3tYZFXxbOUxzTsXPR5o2XPo0zLMmvF
cfmeOLq1iEyWqCS8HFPWqj0pTeG6gX++fBDLuKV/dy6sffcxgknVQa/0KxGUvLGX
GtWikH5SS3FCWcIkysP52+Wqs/8qu60FBr4UWwmeM8cIBfdknOmjlV4+h6PaaEH7
ohyauMVtdg4A4ZKkk7jiRcqaU466rbFkd0c4V0a360H/gU7VXnhnP1rKmY/Ynsu1
F2HjI7F4XxyovSXGxfDV4CL0BQWJuokosQ/Wt8gW64zUpIQIBoNB+YJjzULvQfr0
ZK1J+5dJWOFjqpcrJSdXsewA+b35bz+m7WBhKzNC0vS2I3BdILqc6UQj/66ZBdP8
sU1Gq4SVbWtyj07q+zwUzrWsddW9bdMstI4YzPJnGpiCK3UuePAiVt366yWTDtcu
W9D/8AAP7ktB++q3lBxB65CYGMTDGfJ9q0sN5LKWlPJmozEOYmQiCQ/jIynYhwy+
6cEM83UDMAzpixlzZAcR0YWcs5BPruQsFRtIL4YpRVeE6DfAdCQhxh9sQR5IaZvU
RlgbEJM6d6Fr7+Ma+hRhEGkcpyar5P7tmYiLkaP1NX2ecaKa44+TNjThr3nG/L8+
Q94kFuWwQCUaaLj7D/opcHLnGEvcCRVK8TxT1FuaSFvOEsWAd/uYDEn1cy42/4f5
uwLb82Tx9yKcqF5VtCKW7xNqCIaKZHZl1rxe43xL0YUO+n9REn7MAv8/Qb09j3Rh
PsTuUGhZLJh+dBIhxBRcbYiBXIo2T1bNPMuWaXJGLHJGg0S87c5nb6NlvRXvN5R1
DcWGa6CUZKUXMiHqvC0BdDMjx/GWS74NbLYDfHjydPjM332xiPAYKHmkyIaQNNFO
95YpLeh5VtvUJHfXU7a2V2+Cs3LTwPzQczcFuKLU5OUlwDuCMPb9v226oNM5Nleu
GQqSJmLWBiIn1GHWaIglp02XSoQriO4oTvD9FhEdy1tZOTkhzwxLJCfyQ423QPqN
5O1QXBSu3+9epg8KvgIIj3MTViP9pXOxw2RdHyyli40u5QutnwsWsWPlsFwr7DLq
fwMh1gbVoKAv5l2H09xc5BSdeMzV3yGvzyrWyQFTbzyYm+lyr1zrsnofg7eHGn/c
5VsEE14QFNFfp7dFIJ3TYiq0mnErz5QpRVUGrQOH60bZryW8orkHbY3ALAmhZbuQ
DbfiKwm9faYIvdZ5skHAPKKDz+xXUsH00BIMTCNTPHN7qHVzIRRJNuDYrk/5Bb6Q
9tzxMZ43ZNQgUddi9TvkatZGLjS3uUbStiuCF6giqSW0pp9N/zusq7ySPEjL+kNg
yP7EX2knR7xtaFOKTZco0smgwWsr1J/+sL+VghAGBDNKyIH0Ps65XCCV5arSLXKn
x+9CQo4//FNAdUw+GMFQ2KUW1TOavmz8mKF31galPhzAd9eqn54NgqiUiMdtElEA
LnpxwRe7Od4Hx06G+8Zjog==
`protect END_PROTECTED
