`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K++POLLfdfchDEQXSufVsTHbuvyaXbZaJuErvRrsnOPaD4RHtOGQjbxssDuInlfv
A+NbKENaBeM5FQ2AUq6EYnG1toHLo5Zo6kBhsYayPrZP7ueG6K+SE4wiXNY6aqfh
6NUgraS4sUpoRuBrjOoXhMiCcDy3HhxaodbzMIs6c2XEOHAGI4TE/gEGqX+Hx48q
6jUTdMCU47Jpc/uXZDqxDShIkmdFCp8uz82n/ZQVvy1397OeQaxGG/az41gRmcg5
o35/Y9+mnlzT7qDovMz23HUdOLEVRy4/gGIbqf6GCmOAqV5kxFKS2cW8GSOrlBe4
1DqbR5dXcW9ZK+DURfdsR0c29svcXBsdnST+WdjTg3tpbIsWSLYwbZca9asjmoXu
b6mKZ30UOsEERZFJsuoLn6mao5wy0OQj4iKE18fvBJc9EsJMSOWMzvDAGb9VWk/Y
pGcZ2NLGyidcbzbrDpFRMJCEUDvUR4uloqe+MFSOoJqIVcSorK6fW6hsFjFBmwha
uZt/cemeYoQxKDOxtStXnlBpgoFyiC7vcDcx3t9GSDuJ7Prkze5jKWJrmRGo5eSq
wZxyc9p7zVdWIYhZ8GMt4RRc8V6ogVcH5BDDfeSBQYT8Ccm31Ov3Ow8CYqg3/VaH
RA6xtqqNVBO3AO/ae9AOBMrv/PuKRd3KxaxbNXWDEY2H8HPX8vopJwYLT6l/9YjY
bi+7GAfH1frti8H+2Ea3oxqo2EkN6GmJyAH52i+YLgWt7nNhL6ZvpMdb5+775Yhr
eW8x0LtaTxf7UvAke1I9FSZ8bW2QTHjyaXzzRm+7dj3da1QczBbZPMYvKAJrwFOD
zWMH1y7dOS32TaNKMTlAYr6z2PZ1fw0G8/inI540zu/7EGbzU2vgvjYhE33BSZBZ
gid7kZag11gr5TEeYrAihAYa2wU3OovspUc5tpBVZnAh5yUrNfmDStlBlHxhpbPS
ZVka1a2p1mWvL4fhwUjF6k3uul5VyMcw4+ulfntnCyDT8pLxrfpp9TAG0qfQM0qh
sYlQLvwBM1x3ZRmPdC3KXnbS5gKMPt0Ncr6Qxyws8bhw78hg3aM/lOk3oLGi4CPp
gKUFEFHJYOykfYW4qt3ns8iRzuuEvszFu37mZwo1lGcmwAOLJs+XI15PCtQ5VXB1
Z1DOCyV5/pZGChvrVx/GOOYH6Xq9+yctbud0/CX5SFBQmZBo3G9LTQjzhCKHOvN/
/w9wFBN835LMv1UaI/DsYLbopyvgPCyHWFplHrLegEcoJCOPAagmU1eYk2FqrEPR
e6RzrZ8kdC9mEkjjOuFAiXMmKWxjOO5zNoteqJEOL+0=
`protect END_PROTECTED
