`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0DfuUGwX2rZM7S9mdgPeSXTk7/0BN86BU5MHInK1f4Ui1Ewch68nF6oECiJKXRCs
GdBT6XiJ8abB9+A1z0yM+F7FEqyZG9+zYPRDE+rAZD2P4qbPkFhaJ0W0eK6emzUJ
3/DDYIC+zXj6ineYk69tiR6M1UqqsDjo9eVwWQPB05Zls3SQ5+xXJl7NL+rv1qjB
PSQ4N8iZTxhmWLffn+fNjzf+bD5ygddnH4cySlCJTfK2aYUjRXV7lBwc7t3JcjkE
FnO9O8C+1LwettPy3jIjr2RD0SHxXquNl981cDtzSa0tOtACzJ85AgNwbnbqkgv4
oRMoZsnq/vyPrVrz1j2ORMO5NLR+hExZfQza2lEAw5lpVUs4XIZTmw6/SsPxYD5C
KG1RNVWSO+g3/REr8VHMUf9TN5D8UwbdKa0oEWKovVKQfSA2ECj0tnehNScSwfdX
FYHT/v3ehy3VniSR3KBz0jyi+sca/RYPgQVcfU2eTwKvT6bo5agJPS0SBcDKgzSP
Gked6+JqIZc4NiElt0xobqFxpjTvENrBvNPiYdXJNh/qM40ABnP1av8bzBnmpZ8i
THilpms72cUpktCvWTRqvedQ3IpIFwwInXUvA9MtzmgMxMrnkbr0vYUGeYoKSQN1
2icLg0G0ffd5gtyc6EL/+EshKAkwXtH4DsqIUWptqnVaOuldBTymNcGFPMzazvJc
MWlTozlZBZFXzXx0bYEjsDqWcUpqK4OUVrbAVdZSRF1eJfT6T1iEpPzOBsUHhoH+
jo4SLlaMmS/AbRzR+2sMP5/9878B9Vq5s0HUcpg3URX0Smxqqt8G0I3LKG2MAWA0
btjwDc21R1QX/8xz/2BYvOnYqYXvJ76LCzDsK7AcDn5u55STCspJWQw9bUOe67Mh
H7P2MRqw1aIh3NqetrUcx9pkLBcgel3Ef5vUpg3hxPQ1oxmiktPUFsBJzCXKVQKV
IXdXIfOYO+l6agAoNsuvCNNOk99T7O6t+VG3Ih57pGNWw/ZbG0CVZF4UGmzr5ZEW
QMBpa9uNBIA/8yKUOimT8cHOJDDeNc6h0+QuqHyRPylChiASzJhQVBGftcnLv6gD
x9tCW9wBhXKlPg4GpHLjFMaaC5j5iX9t0ImqQnqRlgf6us8bSj51aHWwS7aLimMs
d39rDY0uVEJLJ7lsTJMJkBuIedmAjnBWVb8OAVTg+KQXXNdjYR8Wn7m2nfwEdVOl
ly/3yq7zcPSylJ63fvvkI7Z2HN8q6qalIGnYYdEHWpALMgEJSgAD2f3NsUAug3I+
GQxMg9CHtOQ+GYJYxDbusHiWHCHfyoqPxsgMxixWn0uaTLfP715KA5Ac5BYTH2Or
eF4S3VdjxLpLaQdZ2oWrwXIkXcDLIORgH3qEs+u4Mkd0UhFXs8f/KhzZHE5nM3vd
xwnP8GzTiZJbc4HomfHu47bmHoETZ4hc6jGONYOYFnlF2Yem+qdkkUZlFVyBZ29C
OZ3e5F54xyEQ/5I72KV4GG3XGtTug7MgRv+a3tf/EuFb6pxOyZDYOB1m/hy5KkXm
hek+6eMtjRd82kxaQlifVOp5z/vrGxkuPJxogx1xo7PFxzwOB3yRSS1BKRF5dRuQ
41TVasdlYKiqzYV8rmuYDF97Vt3QL0Nd8mVarDMEH19t7CGXttAKydcJnP0Cepmo
x16fxntqcehqPesMvvOCwH1qnwwyAkN9+cFmwJodgPTDJY1XieKpr0VVL0ZsaKxb
r1D9VDjbnpukhcCUZuMZlRbeGDpTBe6Dbj/RZc8NS4Xj9AC3/ARzZuEAUyCemBEa
lqWwHDpqG7xqSLwqo6Cr0TQS0abxeoFZ/ax4TnonhnC7hDZBRCkTNDEOAY/lOEqA
DoWg6oVv66dPExa/AmXSWrz72WaE9Y9jSMnPHe0NcwryNpeB5Iya1fFLQzwMkNE5
m73clrT8jdb7krtNIlPjEWRHPnF3d8dUwV8SuljZ70s/DVUZb8QMouGS/hZskpHr
QLYyqTTpOW6500saaYtUrLlU4SvfSdSZIEQcsbNy4leilABPQAuDvRBlHJAtbd9Z
W2cHLmO81NSN4hxXz3Msk18BsTPkmb2g9PnA5I0a++ic18P2l0F8TdjXW3R9z8x9
cks5G7AA1FSG/crqDiT67yEcai1jgPoc90fNNwcQCcfofQq7bRRkteio4UtxZjk9
qXhUbEgP+Npzyga/K6K9icPnqBB2TOrmvHIw/v3ymiMRKVhgg7kzsEdUf+ogIl0e
m7W5F96xf64GN3JU1Q5ipyhwQ+4A68A3+EjiaaWI6e1CFoF2Z81z6ErJe0yoLC/h
JQaziaDbNT6Po6dLqc156+hc1KeHfIHMRXA2Xwf7iY5bcybYB7tISMIEkb/xko4p
Jr2uyCSMsOiwvNMA84sp77UbVs+gYo4Co8I/Ls1sp3vryVgDal1GlVNKnOrtQFok
kiwOz36GZnMLpo5rrJToiFIyuCBpvcxYUlhOlPzjCHnE5mbEmtmQFvd4hrv6qOTz
f84Acdxm8dTVVwcFzCGisCvTNdr54j+3vbnPyRV6PXZ60nJZfDaUqmTYOunfcap9
d0noYZBZrit9yIYygyDNkXb9+3mQgNR/LGIzeLhJdpgINvVddc9jpTnwxC5DngRD
ePMlDXyMzEHdNeiS4fQGYirgYwU6blyMyeB9YkmireK5qGkj/T/rNfLYnhV3c0ud
q+54z2vNvD565MZqz3+F2RNVfs9Jx8hGkF63ZpXf5ZL9JUOKIJkziRqgMK62VX5K
DZlvrO6gVNXL3JpvtK3IlUskwJdprNDwv3Hb3EfQiXX2HPiGzkUMPwPbIBovXXB0
gq23ZMx+HJ8h30rKadQa6rxI7ozEYDqoCItjwlFUHIyBckPoP8lRx0ANjtp1CmCA
WFzF51JBOCRkullY+x8SldcrbbYG1e/guozWUbb6WW2oWJbFN/wO1o/nEQyG8nZ9
Orzq/yKl+HdpTfT9QZaI1fg/w2OybDsnCW7hJMHO3yUhtk+HgwagcOKHfKc35KTD
LCUWXQ0QJzaa66sJwwLWY/i/OyA11+S2lXCWRklxwWEtx27ITtw4j1cCEqGZ9yA0
Fhz3pdI9nvxME0H8vhCP0uEr9QgaUa8Xx2XFMz5/DPKd+ILbP9L2uwVGLn0d2HeE
nIaP9jRWh/Wb3rcymd35eY0ZLem36ptx2AlG+RUm1ZMlJDMYrqe32fLtG/tU15Xe
O6dSI+FJlji9CDtOO4N8MgBG0lSqFnibkVmcgTDFSgI2kCn1tM7iAiWy9gikqghm
cOIW+owsrMDiFdd8id8q7tl11hK1uuxl9LqVkzHU537aL27c7Gwx0HBHPJ+r9o7v
v1CuMLZFHlztQWnR0etc5/9J4zLtL1gO7SFBa4AwVGpzw/yhDIf1y2fKf2mHlC0h
9YQAm9EutFNzdd3qzIGGdsPi1HJulkADMQzhGTbD7leWRHoWQAxpxvbUDVeVHxSg
mEcIlxazjprih4qDQGDXLZCo1XRJwrQ2SOWlk/iFaK0QqK8Bfjfpn1B7WLvNnWww
dUKiBx8WUtFomxU7t7UmRVHLUoTGhweGAxqpo23fkzFWY6OiXgsUyl/prmiKFRHm
eMGidOKJMuGjmdq2GljXeH6ePZMYleCbxVqxQH7fQ94ppSYPzry4W5MYT8IkaGGf
dexKU3KVKmxvmP78Cygwk0iX861VJVeaq+nUZ2JQir6bAQ5zeIrQouJxTKYMnZ4z
lFdKAUE+3NrXTYFrSlc6iggFREG1BlCYC3RsdrNj5rFQo5/p7ntzxP4x5oMLnoD9
L8dB0NU7Chd60S8p3d/VCzpxlCwKr9IjWRWt6Plgc9VM0I2dUczcTgJaEo3iYw5D
QUyUX42PUPdS7YwfZOlNgM96NSj+CUzcgjuxgPYL/R5F/AeW5b+ByG/nck5m4Bss
XyTFd8r/5urzuJw8I/cKpd6qEx6k3saEEG4EeiELijLvNI/A6g8qqhSdgGc7DhUX
pisRxl/YyOKUjMdNYGSB+ojUKeiK5BA4rMfXZlZukjDoEXgYSvOlUqaIKGsDi5ju
ss7c/d9m/u7+FRkmhGn4gWudmsvmp3B3Uq5JuTFNwdPcsQdfUbQCfcsepkEmjpMO
MIG8i6bHvMyfFK+8Nau9+y+3ILUCjQ21n5eGx78Wi8BrsLJ+e15L6Zhrfk55lZPf
OYQcokA0FN2oxKxgKhmDPujATo4gIJei931OViv4E6c2cd9jbLKjClkBZEafLqil
GM1+1fEW6xMFyxp5qQEPPVDs5AqRYJr3GbAlEA0v9qH45YxnbTFIG334ZmmNA28p
XgnW0S1xZGm3Xl3G1kq1K4mal4zBrH6Gi9foo9JJJO3pC4CXUIB/lvQ3e/wLlZNB
/SvVVdMxQmG0/c4frsfBBUtWPohOJejYeK3WXrkZyA2yxxlMjNn9Or20ivc32Xlf
4XGPhqPmgdx0JclbT3fbA/LogGwYXmRdRPneQK+PdaTZD/h4RK8bPJ6fNpMHtajp
Cq6MeyjUaDSJeFJvFyGtIbhIGhnPkbG6v6dWnKEzIArSrweZ1Z8wppDH47/JlAL0
RXq7cuRm7jrk2j785xU1l7Ux8oam8jNnFg/71Jv5c3jb0eykNJRErrn5GkAEu9az
DeDhw2d38k/fCt1xfahuPOKH6NFP58fL5MDN/Hi8+4AJJ61pRbvVaY/4S61EqeWP
ID4MCZh/SBOe0zqU0t0ARLltCdH4255SnypFFRAicH58qlqgJfqxmJsXDHHx9ZEE
SZEi+qLObNvOabCA2ixbNEReF0SWqyj/GkgC8PWl4Te9pMyk9WM5X7Ka8oYQO8b0
FtK9Sy7lwy0VA0gQxF8j6sO1RbfdMo818S/Tai4M5yFNRNJvGsJspZbDeNSp9tXF
gsAufMI2F7z9URKLG8FXCgo7M+PDSwIw/NI6hY3X3gzcsmjO/GD90dEGnXwPSYuN
WIMVm8+CLCvpFx+t4rfEVzmiu9FK6H0Rz+jzL88/kRx+P5/hRKAy57df+dgHE7O6
kbLzGCq22kGlpMUG4WV91awmzJeSNgX0Osy0tJsAbR+SbiyKtJx8WllQrOMZxpVZ
Hl8p4WqucdGfMRL0xBNQcx4/de4AAXtEx61BKqyU0Uc+d7AwIlLhuxMMdQ7b00GO
bbPb15ltFV1i90lDFSzylCplcpq54wrfgedTcJflPSdLoDi3TZYLjnUpw2gottfC
0/KB0aXseAnRGLwR+dlaUNu4EtrjjQ1L3ytb4TH7CXn+7ExPXHtIr6sL6XNAxDx7
Xo0lHRxLHsuxs0roCkTmXYmXoTaZBGEaJwah1f/Mr30Gj9cIaRKHiOyTQSc8snqv
wtIZRoD6iLq56v99LXC2vlk4r2xsIEu6jSC3pd0/RgkE+QyGrumHvo9ywEwaA6To
vll5KyGguWe0svVlDoVYRsFYBEJZzFdV3iOCrTm9yunyEkRGbSZhDMGZihjZmxzW
vPTULMqKOnXyhe68H7hyMsYCj9tAs1zL9Su3KGpPEnNygO18w4eGFtRynM/a8tDl
TNXlFAVwbQ7xK8OpfJko3uix+1EMiwVupEEAM/swMsz5WLOtaL/YEPis0ZBXhx+9
FLAUDuI3Os5lsqi6RYnrrsniALaowTEg7zyr/tv0Mk2vkTQaY2UbswmnvmqfMXSg
lzvdzl18K2aq3pYZrL8eFxr2TgV8swea9JzVZyAEmrL1uXSYwh1Jw4W4hbyMwRf9
FIn87imVbwgUR4ThREO4qj+tp9+hPW7cEazE0AwXCzBclw4NPeTdvrK5fmKuMEe+
AeBxTyKvH0Kzr3+qDsN0lR9z1EEmZegSCddysf00fh/hobGRV+Mhv/3MELciuM86
GS0rCS8KZF4KhtSRkNmIuHKCNBzKHZaD9OLW0ZVspE0E3N/MRzKgDwmUg/vJshZB
lUZEG0uYZeKZPJRQWbk/yC/F75UFu+iBba1x9u5qaiSwJ1mhKPIw7h0vW3YotHQK
zhTlCsyu6oHkTLYiwEU/jCwjljFKe53risUo1WmiKmK55aF10pjJKePFDfSQwPUw
bZj+0wRg8wQKNyGtR7jwdMIty4d+XJWODfkMu78wYLJsfpTeyD7cZ8dFTixjvMpT
A0EoB/iGCOOR8csw+loMAjq6qC9DZO8BBRY5LdR10yLjDRDYLCVE23BxkYgM+1hM
qSuhhnzrXnSgxmDavTgXyHGTKhjsQihRY9xIjAlpKIcFFHAvVi6ToEOsRL+iEMYV
cX9KEidIhd7Jntg+D/1rumJCeO/P6kcEb7lqqQUIrIKcfe1s1+CyiSeozMiyH6Mv
+piCsn8KsaHM1ncvXnnbgDXiQ9O83JE3N7M9p5JBt9wp3fZEDBKKBvi/3a/oRpbs
y9o/Hj37MoYLRm2PXKE1BZwtxaGMzXLYtRIEJDNc2Mqqba/H6kZ58e4LSmOGJe5L
ZLHuX2JICFi3Q6jdQw8EW3zkZeNWeNeR/kNHCcbkw3+VEPHw8qAwk4aOX4WEoTRa
WxdqRb0VIHATTkO7jHIDoT0+wBiLiK6d7sMgEpr+B9iYUj2SGaurDnkL7vrsKiNQ
2CssqvK6gTtUfQo5iRGD/CSP0kIoEazpztbyEi7p/YS5UdXnM297ERlv3+MYZ7kX
YzVKA9s8EbiHN3quu/avl+zR3LpnT2J4OqB5ji68hsmNSwQoSjVHX91LdmsT9aAz
McSSix8Nt022KX6CqzX3U/+GT65kpAP7UzKAftcZnWVRx48mSSjEtrDD66IZTAyW
sExUbIfTtrZLc5q0qX6fWBwiDmYpIrgl7zpPLP+3cJBdxLiRf3T9qak2EteUi03X
JFWpJy/0Y2fTRMUUZgo+aUeaojcewEWDEEtauO0FaSJ/eAn8Bob5oxfP0A82OZCL
3SyjPNxdKRvB+EnI4Ns+a1neUZKe5a/7Am8vsCYZNHCdEnXv1NokvL/M+YINwaHQ
6ffjSquw1+DeObWPg0pGKnX85RkFjdEu/Ksr2Fk/XyHO8dH9TnPJiQk5bl8cc8Fs
bID1hny8Cbp1WlB5rcKQ4+AFgpAuKeFeCb7GTtOkqsStJ+QiemcLH6dJRllwl4WG
ipR2aZX54Jc4ffM5e65VFP7lAPjsJIpbn5UAuVgtWkB3fUPh1OoATOhoR3bDvEmf
AuAtRZ0E5O5xXXjl+BphZpCcV4OcM9CbFvTvaqVLckcQgwNt3SHDDEio1IoFPP6j
YnQsYUb5vOrnqDI5mza6YENgXD0ytLIYPXcj6nsdIQnTkDvYQST/L27WAvrcRbnS
O9/Q2NF39MXkGXG7NA9ne0wYkKVErGW0SWyw6UZBOxJOsrxnc39AAoZR4+7QYHXG
eXpi186gTFkiXjSLT1vlA0EHxyf9xJYiY/GfNw+j6t5o2g61iyTfdH/IyQQhUzWv
`protect END_PROTECTED
