`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+O1hN6B0/kjNGWdqNun+JIImtndWTaO3s5lyJhf6Clp2482zyXmwKNy+xKDyGtl
XvJLEOIyAiJuXuqXbirlJteQv7kNt/YFeu3cVxpXAENZucJrkDRo0+k2h4nPmuEX
5LG7ncPXl614aZKmmBJKGH2hfmWDvkQScZWs9cDB1LQk4AQYAmnA1MQuBqa2rgeg
bMffCT0x8VJmmEByTdS1sAHl9riWwDKOiKs0TxzH3pKZPBg9f8BWr97LT44wRzpa
zPWcqFzVTJ2qiSVNdCcuB3p1MPdLkdpMN0E21JalNpEPAhgLuSLLVbCNQRsUzxlX
b0CE+esDDkHmUUNFUX90Pk+J6WKM0V3BZBFC8bbzCaN4lnuIUxiixtodrgvmqWmQ
QkgCHOhcd/NB+E2TUg4ureWgs0wW8hYysgAg0oPiZkcNdR3NYbSiUMtcvx6x+uHG
0p12Bykq9eQ6ClvuZz+2/2R2e2XnHax+BC3CtUVpOyWKIPRRlGul32Zf2JFzXeq2
v+Un1VY1AZWXZQgEWmohqRVJ9owuCGd2t/aJqz7MMOCi+HyeZfznOc0oLZQJ6xt0
16HTqJGx87uD6LZbHTJeLmMcyIBfuZFaCrEUo/TaCV2z1kDtbgIFfxMBXxl+/xyA
ioHw7QGTTcINL4xsYrSNbn4ssuPDtTiRi+Ng6yNBB22fPYVlcgyJUivsURLv7GXM
atexuDu8p6q/HuqJJhBNcRhs+T/CTXp7T6L4c0tUwmYwqWLJRj8SDyfXzGD7RG0U
FSDsMm+SRLw7UwwrPAvu2Zt9rpvSKKVk/YiG+/ojDkO9O+RBXIYeT4PytTfZL21x
GLJrSMjYOQWFKq8TyGq6P05tQq3oumQFXEbhwhNqdbvsN8nVi1/pgOkiNlVkYoaH
iRyAMGg7bOSy4URLktG07X8jqqhuwLXpwwfMqgTVyOQ2EdqcJfRGExQ/hZP1QYTG
McdkHFDMp8dMedWNQVgmMqyXdxDP0/QMYQyXwtsjJ2n89VyMHV+GnlwPZwHtMoup
LERoQ/63FCrDT18dZw3oyj9imPn52VrzW2lRjh809sGqbnw9QTaIev0h8vELC8rE
kU2oGphRysGPlY3WZ0FqGoJBSxdE203uhf6yjB7Hn3h53UNQ8Syxyg/zLODED2Kw
n+jYgVNPueAb8lJwwZ0UW42LHBc3b8/zgLU0LaNnQbYeCEYHJ4QOtKA2jN+ULs3r
W+7MPdDqD9F+TkkTgt+K2LZfnk2VZWbQQLPuYFqL+TpcLyzLxd2fp8LG80hE2CLK
jvfG9uPckn62hVIl3lDu9IG9osf8DCPm0i6T57s5IoOErVbqQPoKaRp5qQeLJjJL
gbhn4zMJhbpWU36wXxp17AStS/CQ2K6MHP1iMHc+hztMxxPFPBLQFy27iVJgBF8j
Fln7C9RycI1Yjg8L7XzPVKesqDHvl/LK4arile/R8fYm6U6uqY/KJRZ0xvfYa+YD
RF8UipdPHonG8kO1tHnu5MIKGSctnG7wBmADv55Gzokx01+jsM5DZ8mTl6ZJsz1Y
o37cPRc79lInXgvutxexJdDpD3Y5B2i9m348DwEG6DjraQ5JKVkNgCcNiABVulP6
D8nkEfQDUem7RL2CHT3PdFuXDI9Mno6UwtUboA8lKNsCBWOYoKcELLqtDZ4ji+X5
OLuDybXOpOFnma0pHzpgghmdrhEjL85LJdAfIqiH39nlsSjDAmEo3HDY7BkQbuGs
82HhJ8Remn5ZFUGeuG1ulxskCRaJWzYMRkb1MygmbSgSS1UGMknbjyeVnpcpExkn
0ucr7DTo5SF2nyCaArpVihU66enltUVGFWZ0aygjIZhZQXm3mtwss1hMWApX9wUH
X/9hW4RtiatT0TxnQka8rIlSAy0ebXVihquVH4VPbOOlGso3ufi49CSOwe+URBJU
DogzjaYICNU46+vrLW9GPTTMpeN0qh78vrRO9Yuk6BuqtwuhhHye2L7ei+/ZUmM6
UJ57zW0SJBr8zm0o/96Fet2Eljh/0wuYMOGcop3J0jr2kJnNePTJnCIZzf3bA8WR
L6yARL5eIyHFXw+PSK99sVLZgfxyae60EellsMm+Z/TXJ/w/5+i74aHA8mWl1g94
LiAKPyPSsk2Uxcg8wzSjZwDN0yViNl1F2O2mrOaq0QKVvBb7xUh4oIRzCZQqc1mU
XVG+wHwy5waeS6b8hZHIqeSqS3LcygOrolbuad50LK9ZE+Pevmf1UQ5moNpaIRN0
jd2u5DKOsKTkJpVpReJ/brqMFbzM7yuw0v7W2NyO/Do3JDpodTt/551A8ZcyJZPZ
vuMMifLEk12eW8y15S4n+sWipfOtRy2ebq9SS+VEw+k7kTOOUVYonhnOv6SJBmnx
RZGLaXZj2RW7hNGNLP5192SCdjYb/IRqkyuKcaxBav2DLS7bDkgdACrOufGO0q+G
yy7g/EtOM+edzANmxlmX/pbb/1s2lTUEBZ7Big1qSULoZNdM8b2+UMMvjdvf1eqi
Crlwu7ND7ovV9Om0EwxPbjZYIdclxuvEa65FYgnQGp7PohVAzPAQz5fphWYNbI1f
Nni/dL+poFX481vMt3bFoSaQgWubF+cId6IeeHdMSLofNEtlKnvajwS48S2woAT+
cmymDwJBlLediBI4uEfdphVpoTIAu0R0pXQ+jLmlNSJpdy5wFkke+Vfbt+PxGB9z
uY9+PlgDQRlqSrZkw7JoaWcQH3kjuwNwsB/bQE/z6rb8mbb5+Uf7EAoIvMHuPCV+
QofIKKRFYGARWya3+wHjs23wZKDjQd6obr5sOHrl3HMKXlK/s0BghJ0ELF5x9D3y
qMzXycI72bFU9hlB3knFYZGwE3LROVcKpEkbZyv0G5noy0ZxEm+KEHyw+sPIRbOK
yoPNeNMbAjSvZT7ampBMCg2uYnEPpmnZcartr0UEWljRHRgGhs+a8b02eWng1sLl
/Ol91VsFTOdPEEJouyNZdLGLRov90FG6BJX6BVZwKc9eWw6WqP4RCGX10Kx3RasZ
MwPxhRB+Azy4Gk65dxU/oQhqdVCqnaVSlYMUM0dZkonSotqL4EBBT2j5oO09vP8r
k1d6GU6B7np7UCoAQG3PZAO1lnqZpv8lB+epRXJ4kyO/mkfiHMEweEj4V7OBDvV2
PX13pAAVDUwx0lJcla9JVcE6nBpMCGPXO2+ODm5yUfrf1/SUKoC10DMh+hAbx+47
Ao6FQEZw8XcFcLC8wNwm+Bv3RrLDhfI9G5/iWcV9mB+Ro1Tz1LvbkfiwJ/JIIm+3
YMAd/WAmsxF+xy+n32YAHiREpHEBW1+05w7lB+NLP8G+0qt5zuw50re1ELADVeg2
DuZHfFCTDUGBZvvU3XZ9goahtUdm/OL7Qvp2lw2NjkksEocqJN441d4BPE4IL73e
4bgT+GkCQ5U+AfCC+TVbhhp1LnKMV+VWrUktsUdU3tE=
`protect END_PROTECTED
