`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FnQ/m6Z5gpZfRL9Rys/moOw5EoeWLcc+js2Hs0tWCNxzmQLPWvRExJz2Jden2x7O
9+4zx3rpPvX7OIB2O8q5Zv9BBOGvI8IDF6ldPg32CPSPDrr4lhrjxVuYWgGYlSVZ
6fGkniOyG8FBnWEu6ZxJkr40Y84TBF0rWQz7FAWiPAfDaOm2DNqG0M5DfYsO2ZkL
jyEP+W2hmZfTm7qLVurpTnfZ14RB7H5dukOqWYXW4O4XcJS3ZmajD0g9ufda8Ptn
l6za/NMeHNE1kLctVCwLC0SJlitXuQmgtOCH3gG4wrZBLHsVN+SOMP8hZQ+rgQUs
d1ZDwYzznwAbjxFm5jUPUuRg7W/wj48Gtb1o7gwUD4QQwyZQ4GqoqU1a2iyoelOs
zFfy7XEuZ8vAgsnrjOXJKD06VgRMHI8ffXMyUq/htrUEAWvQBPG3MALwr6XYB9/T
Xyot24pK6+Dwv+R3NZ3ieoYfZJcSkduuI5dF+6iAc+u7R5+8M2mSvw1I5X0n3FUs
/UC1d9KQ2zavq9Q7HGOP9g==
`protect END_PROTECTED
