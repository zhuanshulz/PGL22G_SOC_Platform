`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jX4fAnkNKUU1U1RH6fpmKv1Ux06ZY/GPG7iKEWSbxICrE1ErlIHv8dX3Jx3y9aVZ
hKo/YqZGKGV44kxGqejPWPa19753WwUlSv3+X5vt8RbpH2nvfSYEQEvV9cSn72ia
wYsVWKHXONm0k8ocVXIn48OKANODh0YJNyiexkwdwLlDMAhJar1ojZ3JJPXzkgVj
H2P5G24CnXQhZ/z/YAhNWe015wk4qoB4sW4slBnDW+zQs8M417HR4/6G6qaDesYF
8nEi1Ap31NGv6cGZHuBJDcD+UXy5N24z2V8quROOVBOBlxCE+q4ugDjvOjJrIiJs
VthRRdYhfEUa51U0MeUGAbYReUZNrUdRvM2YXUSm8mgvSMGjN2581MMQEk5hlUrz
Csx3yvYqhow37u5rI6qWCewHUFvTmVextb6u3xtSXOc0ljNIvZmfwDoP4W42xiRN
pX/GJJdOo9gztSpsbMJZr1lhTvgLuM95Mg8cDsjLb5pyLsnQqc4LhDCoOR1H6SSe
bCUBReRyA9JV1SY4p60n9xrT/NiSuJAkup1CViwgnZNUtqcQIagSPK59Ujl5fk0f
l+i2LIkHHFln8D9x78enwtsxyO1Gpvv6p/s4NKOB5Ta/CgwK76thMXl3YwaFYyzr
PI8YeKFiFsQ6liJUl4tWYbeRKqsItG6iQjE56aC89yd/teOP5iAhnOXQ21das3Qd
oDN8Nq2lZS2qI1up9K4WJt8+PvvvUoL2LzTdx2oziumV7d3WCn3060etgs+KSDVy
IRib1Hg8HOv0HzJnjftsBMz7so71+aB0Cf3O8cBsYiNfOpR/8b1igx+u0Fh9MXwO
`protect END_PROTECTED
