`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6XOkvOPYBEfZAe20N9ssw/D6CrxE9MPfqxMrvfE4jhoZ3LkZLObvY2YR2My9P30v
802B2W0a43bysRwgAJAkXqoLk6RjSV7/00rGE8m9ITcvJkSVw23sAJCa7vu0uC0V
SyUhJgwBsacSnThcq0m88w37ZlgZbr56Go//jky1TJIArm25OCeXVfn/9rOhI6Og
WfdEJ/+rse8YTsOwDMRbb87gnMsPxDB3LzgENY2ILvCGzfGida70V6H3EW4n8zuW
eg1hNQoq9P7AzwYXpDzqW7w6SWnBxAPa1bLpFV1knCLzb3bXM1351bRTt208Duae
sFMkwT+PAtprxGSUQQJMEmScnDkP0tsLyvqOG3sgM/QYFR8nvVytM/NdnGW5i6Kh
DsRdN46l7z3fL0YFi8NSap2QcRC8uSIq3ibwezKKRsM+p6IUJwGuWTyQLyWABBNw
jt/HZSz47RIjQNSSLMEBZ6CJ5LPJ8/0VZWOmLRYo6BrN/v/OGSHeGiCALZ2/S07r
aT2xyAm8CrD8wETU7kcwzCl+6svL8oafbT6bxVQg5drsc/ssWSYFQljRRbKjr0Z5
jSBfsV7Gq6ru5RndGTkja2P+Wgzv8hq46ls96zD8hEz8Zzz0J8ww++pb+umQ2M+f
6SOWO6iCg/1QV3hc2O0NDeFfbsvHilcc5SFDEOEclwlT+ITAUMeDN1bapbCAdRAo
qqrvZCygRysu+ghK8uNzOjincyW5Q91im58RlUgURxazlsN8HEQtDFD0sr6NxA8K
6PciMdk0CnU98+kuhDH0DkXm4Ypa5TvTcXW/1a2lEVM6jlZgAExdRWUI99GmC+kR
`protect END_PROTECTED
