`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7HrpM4qUkx/wSbU/gmKJSCDlxsZT7P6xiiQoowyNA46uWO+ZM/WUotXzbxmkG3H
BfdLaUHhJcyCMAKmKNq6I8ZGoKBMKF28VtspZ0pnASYui2M1U2TWPHvX1mQjZx4F
EVlNPelLGdTTqS2Va/VTGEVWJv4zFsFmZEycNxGUZW/mPqxPPjWkwHJrbewHXRTm
oLfDgbbfiF9vpTd3/30agX4/BK3dgZiE5cD/i2WQikzOLsYXG0t2Uxd+N0/UwwoR
wHqz8nwATRalulI5sTQu4mYim6WSED1//YpzTAJ52JyR+TNYCBmreBJUxjHUxSY8
7ApcklJf34wGgpxyJkrzD2+dzm/sPJfXZ6klkvkw+uwEeRrqDdvxkiwuImz/MJyR
nvUhdvrBDf3GYys2LLFRNaWzWkKvx16OdMm3lJrW075Z5EBev0cgY2+6AUQJM/V1
iYYjmLtt/CrM7rpjttDjbYow5UcCNCid59ZNEoxm54szAoei8B/XXwG1MDsP0vUl
jZS8hNm1E6QYl0j7t17G0CMRrNpnMH9+dk2Ihgc1XJxLcJv+LhzWb4SwGf89Ly8y
0fBnQFHWdO9BEV5fJ2dmbfAXZQK8LBoVpkqieQ4xKR8yBvsXNxKxboFZqiwZTfSb
YuFLq4ppR4inIduI0TLAHJm/f3g+9ZQAnWH6w/5/5bfGOg2QChYr0WnZRDmr7Y73
mKjKt4AGQNRSqHIRGuhpelTJGV3v993GjbDW1TMONSBpee3ZGU9Ux5+n/9MMBLGX
85q0irbTWYX4J2nPauDlvA+HmuCmm1lN0RRAs+n+IrGRB7IuC1bQRpin0SJJ3Sil
OyA5oYefRAIYpNhmmYhX3mMrDwgJ0pUTDTCDiPaulXkWSr8/mxJbecytI6/TXhSi
nMsfz6gLRQwq1buP3kkCifML45+5S8UcAxPiDFrboceBHopFY3GmUOr4h9bge46y
H1ReAklPRwSCtK5S6fLkQH5XPwcIauJrLHus4+4w+jwpf2frIpdSdQaGRTkAdhJq
bmi/7yRY5pzQGw+UJ5C50rE+wgfSc0ZtD5dcgVPEyUwnzd8H0WpTFNyFX92UbHDg
J2+kSFDYTup8xGqBr7tfoU9fZfvGU603ytYCNZ61io/4qeKPA+Izes7RxpifEWjN
UrX4iEWxGdh+vxiERP1HpxMKs5LdEiPz+Jr3BY+qP6tT6JrtbHo9Krjevm+eNzWb
U7xXKzqgJE43ws1PFPLp4hs+FQU6NMGiaUMLOddnaokXSwcW/ZcLOANUMgxCT1Qq
mnyPVjdUlTLt1msRXmXjVoYOY6ng+XPv3sGM49Sj7S9IR+WEL5kR7YF8XnQwoAbO
w1iS5f7ECCtPfp1LU2RE4nxfiO30l6Yo/+iVXAMnP10C2QUFP8QOP2NJQH+zDTBb
e5HyO1QHeBv1IkvmKdcUDgtIFkaPFY2xR+h4W+O+W0tRpcR1dZSpUdk2F0kAGe8X
gvpls4XXnsDXXarMserua3ZkvGjotT5P+TWN9q0eP6wSpqk9GvFUXkyFJWnN6nFj
gFbiGWbPPajjOVpNda2vxQn6/rn5+Hnw9Bx8nN88ZW5Jcph/IVuFEpb3kBooGDeN
EonoHXVxIdgLDPYh44JEK7wvGJs5z3h0fwkam20HIwRdl/as6hBLJLUxAOajKCvq
gfXmNNfe2Ek2IJ+WS/Ig1OukqJeCnCPrsodxiGh2I49+rzRcQ251j0A/tS1qVIIJ
lcGCPIhTBV2AjtB3w55Mf8wEzAw+WY+ETL3vZSwSHDvDrnn9nAH5MXm1BUiGF8ce
+aKXrichVdPK7eSrKaoEo4ymGYrcHf6S+MCE9ryUxVrzStBrYK8Dad+PUXqSADnJ
g9gSIKpbXyLJDfUktKdIOlELL18X9yEi/nFGNuzQ3OqJSoGrB9Ug2E9Rukcipf6u
ElUYtBRnc2H9HyUZutM2+/NFT7NdCWpLXi4pry5XmqqInfjRZCgUDp7kD43JLtuM
oNPf9PUzvxVej28CvP2ZiVPr69EK/OixjC2HwaG3RSGFtAdmBNVw8g3E2/O1AB8C
IXktlXFXJdbvABJEB9blpu3GYA3yGWThYK9g24m3EWBJ6a0IUsBtqKTnv/HHI08Q
HH9tlu4cWtm/zcp2EzbwnQ==
`protect END_PROTECTED
