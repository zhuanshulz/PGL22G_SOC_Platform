`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pEPbdiUlLvYrfRnEEUTKpRMVv2Ai0VwquztRKxTUn79ccjnIrT527dki0QQyIqoj
ngqYiUvGmvliO1PN3crtQ3YLJbMlDi052dDNbDX1pemgwNA5BXc1EW2zxq51hrfx
k1+j5JuNj4A+ERjKqbtNmQCbTxL6YrO8JPn0jOP8mVUsUGa5ZOP76ExFlziumnN1
DpKAzX1vHEUcyytyujNafDXTOnsgg1g6dX+SUkdBMSDaTN+5IAMoh5449KGJ3KzV
dIYQCeD71Mdcqz19TEPu5wlFXN1jfAqU+as96q5wg6IZvC2qzvkQgeuu0KkVGzrH
YGysAOP8/Ngh101qahbfqcpJuO8AHKIQ1D/H7S4jAVvexDxToo35x6j17beUgx+4
HZWbOI4OoYYzcdgJdb0C9WLv2XrNqQSgOegkhXXGjV0a+HhRSbDf6Z9d5dQv7IhJ
zN8GgaG67iu2tKCqsouhZk1Pau0ovYl/Pl28CD8C5ZFmp+HJvovNFpUfB8Winpuh
WWwe5xzEmZXov0IcQz8PUyAeRUfMAx3UzJBU/Az8f8tVsPqZlxGskBTIZyoh8I6x
D2oeuom1C6sdQ7y8Dzh23UTCUmZrOe0yGjFptghJ7R7nh2RIIPIx5aCoA80FjWlI
THFBMUMUqD5mZ0cPNh01eRhNkw6QuaxUatmv/mFSXUIBQ8sa753TKSdXK7oJlDbY
9i5uFB1F1X0c7QHXXWJ4rr4bD+1nnd1y1FGdyWNGq47sG1G4+j3TgWMP1pf3VJEM
TFEV+XsPp7WHfsyYS1wqRFAOib4FvrUJ2OAh1+Hzo1ZW71LbKGmYVjzvoNd0QvSk
Ltsu6gQYId2dYZw2s8Ah8+VlGQ6yQgYZG1UWLyK5KqI7fTW1rGqrKWo2vnH26bbD
ypyR43u06b0XyOFQfbB7Jw==
`protect END_PROTECTED
