`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pguDhj3mI1gZ/R1grlw4JxsN8tnoFZ+HmpqZYcu5v31k/Q4bJWUD2tvKtKmB8nzo
b4eIV56CWwI7fyNqbP1Xf0xpYkdEe15yMcTwxU6oXOJ9xKoEEF6M5qCSO9X0tajQ
VrV+RoGg3jvKtxfBGxhIwtt88RCmmgra9E8IlvevV4WtAklgPOm4qG8222aJfQtB
f6XhiHVATBQTRtLGlxd9Revutz71TZiTVhv2W/tLwhJslvgQMYz6cBOgmVc+2xy7
gES7lDUkB3gWsVTqyXTa4+kMyxDq6OQM5zu2/J5mOTe3nWJQ8SHnmLhyceFi1lEI
77Tv10jqFd89+eeAoex3MYsgAI27bQhp2Sk7D4SKqvJh9mr7EBI4+0BZ+6VXrRqB
dVC9qGY4JUku2ZJ8SHSIwlILZaGJKjEpotjaIZp4o7wnQTIQQWRE1b30bIP/QbUW
dgUYnsGl56CJ2SkEqK9A8jSuCNQkT2V0BFUkDjsOTlJMUdKh4Hh6hH3MwaEOyM5m
nkMUGbBMXckSgeyLae3qHE3KgSXsK9qQPABgn8F3SmJGfC1srvXHIHDyTA0ytar5
DjyxYGcb5KhB/2+TQjxpF/1E0A7MQIIfrdz1wa5exiH2wkWqb0u+k9EXPW7WoAe9
Ye9lNb6DGmCbiquxyYfjKWpp5SKGwlguifyUqW0+PB8zHvDLaOHG4xCg84GmnxWe
y8raiCq3FwFgDb+y37+HHqikBuQPW8VKlC3uuQC3rwqT8gKOnEKzcJZiQkrQHt4E
WdInlhuQk4FBcq51DAcdED87L7zh02c/dun5d33j2jtS7EyWjj5fSULYHkTvitzK
`protect END_PROTECTED
