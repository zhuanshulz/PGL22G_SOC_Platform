`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hg9aZltdKlpELGYEDQDTB5geU/NvqI905BIvdaHc7EgQ27p97Zq4mj4N5yjh6MES
rHApZsJcDAmTWevsWwNs3AwqAojwEuRJKpwQnGJZE7Jmn997wJKbA+w/mYPoGlnI
omYM2kz8UTwPTgskIL04hI6Xk2ptWUuk0TRB8cPnfwVWcBoU3PO00vTUWCQUIYji
sN+A7uMKJ6y9sFRUhGPYT1KxynQQfSYLf+eBsYvxquvqlS+43CPuMwdltnX55EzS
c8i+CLKtU12IYfjTOcgVLAjHhl92QuwIHo8Cju0qAqfjgyFT3dCZIvMUeYhgGDAJ
reBKfpNzLdGkvNqSPZkUQPypzxBHHbH2Mit6WJNf2JhZjXwMCP2rwk6apPNfiNqm
bCwPkOLetQdG2RG7ntQKhjNYvzTJ/LlaAvE0uCOdECoZnO0aHJSMCSfwt57e+fCf
5jE8fJye/NsET9xM1xtVSrJu4ln4OyBcaCg6UgnaV7/XmzlkONK+K9FspmNTLotT
yXSztU/PQXwJtOVUqQuSjNLuQj7lfs4b6bOGfgqTg9p8LQk44IKTzeErDv3ZrAAj
FaTLKuPxCnleIo2u6ycehuc5sMdE1i8j3LgUT76LDQUCGiPtVLmiGMlgkHXXfe/X
BVlBm+t2KcfSy0BODpcloA==
`protect END_PROTECTED
