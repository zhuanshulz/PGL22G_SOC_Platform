`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5KR3V9pJ/REN09BKCeWcWKEfM/9ugtIja+vZ+95dxzI93c0ksFhxOSg5447sarrx
zqN8a1koowYHWHQUINwuaiqL9Ww96fZUhxJcOB92cdLTFCn81oqLN68FBHy/RRAN
8WyQprqH96Z7RxkQb0ASB1u0Nyde9gQo9m9P1+ld/TAlmcRy5MqzMKXq/03FUgh1
ND/0e2msyFEiredANhP0velZbliOrT17sm9B/IlFpOYjL3kpbSkQOwz0iesLtduT
qUUO5/JYPwB4Y4wn/9/83AtQgyLCS/QdCOqSqqHW7Nneilhyyck+aEvVgz1qzvHW
/MESEXL+r3LL1HRKcfBDdK+dIVnUSaRKkxV9byAta16QQy/qeuDS87hlUbwNzhdN
Kpr72znrqLEOSp0hnK1tvfetnr19KA9auGsLKL21TWcAqaoXu5KmsfubRPcbMj4T
EmQskARnjp8WlQ4uA8UoQFekTRpYGb5rCmFkSakpHIqrZrId8+3y9i7LiuQTCYuj
5seU6CdVl/m/P/n2clW5vRCklrK4vTqBF0Ee3MwRJIIaOQLdfUOKNKDVVAQfPCH+
l3gAiQmiZ66sA7vAmJucZt40ozERZ/BcrClJZXNtIoVpoJQza9wEWX0YDjGNmnqU
TfN5SOVXeV6tgVldtPC+4ktI5ZTCpFmMoxnR5HPOtlmmbfz4m+yeTsBXYlpM335K
Hqh6/+0RhLTyenwQyNi/2ra+7d//kmv/LFxalMh+JluicswbowP2Oz5R2E2nFkuB
1TxxkD6Xe1FZohtshzDqVuBcq2U/fnCECinoCkGssNT2NlH+M7Mh/Mc0pmoaYnAX
SFSDGeZA70mtr/6ADddzi37VvmCRsT1HnQk2wKLvOPrOsMDFRnqxyzitd/qMyfwM
6FbFuGMcxb7+uP1sWmjXD6idSluBt9VL5JOafgZX/5w5j88DLyBzXVx2qf6Kk8m2
WFbKHg0G2rzuX/igseWbfoL49Bat044BKKdzq9FCcMXQFIjLm5F0lcrjPYdRBpKA
YkKPHR29Y8ITAwiSTA8LFRtf6Neh9VXfsKA9yruq19o=
`protect END_PROTECTED
