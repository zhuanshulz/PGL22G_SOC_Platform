`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WLDgJkfff7V1+PI47F8Du+Ov+J9uaGdICoMN/LJIJHFliCQeVBPJqFUPYvpP/rQ
WdxqH07lFiWMtXohbXieXHkEowJ1j+NCx2uDuOE+a/CN4dWVqVrhsRmJNH1mW6GW
QfUWbupvB8plQq9Cl+F0zhKbLI32CK+b8r9f3ks3DbF6ZXjjUVA5GsLC/hhSkDAP
x3VvaE6BAvnQh0WJVAvCpO5hSrzy88BkqzdFHm+/IKy4Es4e14pJedxrXcDvT2RR
x48hN5tkWnKIEm23tk0dExJNyG62k7Vw1Ptp710IYm425ajvfIOg6Z04diMvzTQB
IlOJuahIRoyfk8l78f5auKYBocbXVp08cASI73TZJWvwiHHga0V3UjOlVB98W0Yb
+b7IXlvh3C3is8PfR/iNu9ppE2/yIsVHh73xTmb9qotEmwn0/2K2TuN04TeO8jyr
UtUAx7+K7yimi8QNfslJYt45Ht2IzjickLOqCVvw/EgEFztpkZEWxRtvfNQ7gTrl
++BEbtiY8WivdHy5CKcm9g==
`protect END_PROTECTED
