`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/PfSSTcEv87SCaLrhttwCza/ozTggz7fYy7veuIR1qQpOdGfzZ5655SE3eBH+z4Z
EU08DfObX0YS8mph7rBgCLhGX3rYg1xKE4FYJY48uEKMYDjvFdzU298N/+3yr5NY
PUuZOSZxfX1J38jBQrcO3F7q7j0ho2CAQeSep7JRib5ss0CNFWMMB6HoSPt6YQCm
qEw6tcykSHvApDJ0LS/4OdhlCJTAK6mt18tFRhFp8z+0F6cOP/tYUHVpgCpkotX9
8FI2Pkiicy++qBXGI9WUD3+/QfeIis5Ik5by30aO90dzaHpT7kNc3oSGR4nA8agP
iSbZ3mY0ufP0+Y7ZTJaPTLCnYGrFjPwUfyofOk6h5ozOHVrV6Ybpakk1/ya3qMW8
HT1ymX9qyvljc9NmFagfaMhywG8KzeoOJx5ogSQwgV+ALDUAPfhcrXAANzLcCLDT
fZ8l4QiQWvqOJtMV8N8z49nZURL23ojQMRILtHa5dUv3PbqbV2aCIbk8IfRhbBJ4
gfVfK23exlPe6o0/+42Na9bpNgIJX/HtkDP4j0efbziJWzD20q+CLgtl5DtFBK/w
IiwU9HjcEXJhT/HLLVDz1phKXb3YMLhsqfLspd/T+0gaJfFDhRsdXgepAaXIN4zC
7Xt29DTREBhnFaI2ifWFN4WTdkJxoJD6TSKmqNqY8Uc/22eHp6hGxDkt5GjB8j6U
XIb232QtY8wjoqtm1FqWkc1m12NcxaSMBdNKPrxuoNO8JSkJ1y0FLO73f9iTDihw
rC8Y+cqOq+s7zF7Dr1OIfDnBTLGBzPihMzlWHJfrLrYTMipKZ66elPGHn0fET/gf
McQ9rcEgv14NS3kxRvXaYNYikdk4oJr+Ebn/siI9ZXxbzNWwdnqxR2tJz6PoFidv
5OUcoNBINW4/ltzMFPQSJJaoHbOrQ1pzFB3P3F51nrSEiM9GcJvHEKmomcBjop9V
1bqi6j+tr491gR6YIXYWsBGVnuMoiquBL/5/7XoQFS+vGNQcUcCZqtr+GpT6BKJC
51nPHx4rA61Wu2l5gH0mOYjsQ4/Yj3uCYuZTlt03lctH2t5K8HizKYKV3CRGs24W
F0f7PDIPPY2g+vK9PbS8zqMsXdCBxjaTVf10xyRI9tVnawRsATZJUdOddyV8hH6G
sVuDEuVDVGuu3ReDzwIWgjqZXkOwXtKjiOS3vEATm8NZjfHSUXJyX5/lXZ2AEJZS
ny6sZqKbBQ4480/gbcYCtl6FY9U4329tSqDUzBUhwo5TG/Y7+bnwVpvc/ghnrjCr
X9E3eG0VO/9Ae9xWS7s+glhcZ6yxJS2cwxHlheKJrXI3k2fJBpAT5wl3Z/5iR4t/
NRuMAxqm/Aspz1WmQYnSGGZXhEFnYBX38UShW56RrqG5T+fdt+dOAJh5tK6jYPhQ
7vXRtZH/+6AdmslCnB/1VbW/oE+lc/sJWryS/xZeZa4HmUQTJz9XtRlaRynQ4xhL
KDVlywFFMHLhXLOYqoNMJ+9liDxDwDy2E5s4g+Orctfvo5cx+axqCgIhOx7aNaMf
JQVBxuiC+FBJuYiJxFRodW+wvR3/jokdmT7KwVEWTwsQyF3gUqMDcAhNl6v1XxY0
gFCg51LN37eT8pSmyVdD/DiTn4sBCGscHDDjdTogUd8zM9RjbxdZ2XPyHVlE/EJ8
TNE8b5RbQiBuV3CXleA2s5ZudyKCmLOnM/VFs4ZaKA4qcc/MDd3GnKd0LoIzTpdN
dR3O8ftFZ9VgXUmF2rwbzekcSfNlg7edm419I6lgP9eNtXdYVv5imrpKGCl85TD7
8yOf84wbUnZDZ0p8bDHufYZysl5ojoY3ZdOmeFMgxChf2U6hcwYQOTJKBB0bCTaF
SX8VmDdWzbyZSh0v65Ud5k9g14njehT2VihwXi/63nUWMCRkic6f1NUWjva37m2t
Zg30JUWYpnCsE+rfxCDZxj+8F2M5dlspSGLsQ0eF8jPns2+RIiOarmiTz6n6lDqn
ubMPHH/VueV1Jwcv3H7NvXQP/DK1dmK1FFC9bgnX80JgVCQ/17qCyvlB+SqCIb/Q
m1UAqUZJObeomRIepoWaBsOCeetGyzVATFQveveLboY=
`protect END_PROTECTED
