`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5do0alWNlJg46G/9lX0xMzQ3vB7QXM4MVmzcmNJY4RfLes01JIGF3Ze0nlFkE3M
zAKVLvSQ2WLmEXmtF+XxWbqfW1vU4S807kIObmfK+XTanErJHdDTNiTLEPSD5Wyb
n5ShyJuq6YKsyPBk5wHdjOBgLd2gkL0Phz8CqlcvU+bb+ELvzieuVQ/exWKHqjUR
LsYOQA2Jqov9ESQM288rs2krnR5PQYoCghz8YseK2AclJpX7QUrWYdqp3gr4VKJK
iQDoInoKzABWhiW+bU8iiP8wXGENm1gDkzC2+AHY2iRZ3cmdUyIVeeJozzxpa2uM
0qBlj2aHKtMNtBrtLmsb7yI0Soij0uHDQAjPsWwgRgkWtavgugdruwZ7Qdg1LKwZ
KPuacccvpRx9IwWAnpiU0C3m3miydCPL7/2yXA9Ridyfg3Goqaw3T4OV+3e6TDyd
SlhkNniXT/AuIC43VdGjN+8yhpjcokbl4dJpQ4EOAh5g8xT+rJp9SyDjg/mCKr/Z
xaOeZte5kXZvgSHZriT58lOuRFQON2whQo85zkf7818=
`protect END_PROTECTED
