`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QjrF4EfxvueNr+Qnx6de0fgFFE5FRzPDK2KePRQ/IjUVJR2Kq350BdN7wRV6ue+j
EOzJ7b2JxhUBwVczHHb4FMJqHwhzlPlNJELjxKdOYUcK0q9HzEdQHEKnY+8RMOBu
x96ECiMRCTMowKzyy5Ffgq8kdBQhgo4ZqB1v4QJBcyUKDJYA7rJzh5+5lnZGd9Z3
32oQ2hgkj6lwgjrOClS9oWwQ26zpzVl48+j7XBMaVS65PBStCoIELjNqj2kQhTXT
te3uHGZCpiMYUsucKP88lQ==
`protect END_PROTECTED
