`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MhRU7QypcYDq9P15SwxJlMoey6vVotCNI189A4eYmAkTGcgFTpIy2rMs8JxBm3Ws
XqpLHAusEcGvPahu/hxu7D+XFww1wrdG0rclyfXajb+XIyQs0Y/Sb7aCo2lMB+u5
jCrNHrEpDidGijfrfMmOS9e+DUq7rAqsb9IrK9tHoKiNbvnav5nGE2mB2sihqR7h
Pw2ZPBS0mvqRLPyeViPG1t8LtcLvf20bnbE8rogy4FGRQx3H2xrVzM0cpqNLClu+
o/+PG3QIKlX+2C73ZKGHxvQ5fS/TTSp+ef1YoYjZ6ZCPPCIAEl8qUqlVoTYCOrFm
9sb4ctalmLaly4NjlBWB8fICryhil+VA/PPMnnzTJHw24XbKgF5ZbPqTsVvrkikr
5ZYu8aULxU/0A/cBfOIJrMMO3qi4QDvrq9jIyGOxKga0i0BMni1it+TW5IipLtuG
0sjD9rs9U/oPlJsDim1eCr5afIx6dFqUJbxqCPtuRSmwZwz7FZWUX13YvtoA0e68
T+MiXxLOD3vI8FtZ3usHHb6OIKZZQUXwyTR8SAd7Zv8NhvVaNU54vab5pYyHZgJD
HINaPPgPwG6WspzoxFHLMhdySB0O3r7Dk7RkX1tEvBLyB6RO9w0I0VvbaqdZrDPN
KS58s/gwqoiGWxuDSA50wCNgtOnEATcWJjtHI7MHZ987t/tC//pgpdQLYOaSIKsj
biquABafZAFqiHxUyo1X9Yvsusoh5AnP7lWTSH+bGRmdl/Nq15WI4dPX2QfpM3Xi
NHBWqRWUxDFKZuGczhQSioet1IYuSLfST4NRoqN5Ef6MVrYjJ3vQhN9DETpEZzzR
m44R0r70NtaXe6/sEqlkW+wLH+wwVfBTvhSca5Yq0sBPdwhQd/+Xdis+MRjeIE5j
`protect END_PROTECTED
