`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkugilcyCh7vZV6y6zGTAZo88PmXFBvexlUOjS1I8pKLoEJsNY0XBr9i0Gj7+iEe
QJ4oEXfycwnsrqLqF8U3wqz+Ib7yzBXuJe0LdinchDBKv6m8RAksUWqpDsha5bgU
NcsJVOlvcEkJSy5I4P4kRne9tNniUWpRiiGQehPZiMSSGJ/fwiQ0MqyY93VKMTkk
sLw/04DSG3BC1P/Yxn6uGNXfia3UNRlXfNZ131KGQ3KuCNtSMUrnZSrbwnVlRbEm
mywB6u6KOcB/58k2Csy2wX5b6GnEQku7KOxXuBFFSMnCjrjt+MKP7UgUnIzbrePf
Mcq+z5FcvqHL+d88ln0Jz1EI+Z9LcFNiXIVX+HDvAZUISkuKmjOSgX0KRagvFiqO
A0QxUDvA13OTmMyTnP3iQyG7b5NamrNJX6wt1PUqLPnV95NyyO1ltz/rUvuNq9iw
yXXU/xf4flB9fYVSqx3ZKflJv8D2CSYe63Kxim+KRH9TQdNViqnlALaDzsgloy7c
yI2pSEW4jJQukNTtgVXMG4QTtaFgzWlExo5sq3rOBpB9n+j3cU7B9asXdsgzACcU
5DwLj6py6LWGoNqpNZNviN3prI23HkvOWXwNmwBHhT6CkN0sgEB1RIxT9oisA3CH
/OQDZcR3048I293b8d0KNRlpbgpG/f2P9LdSbCyOUCfZoifhSH/w6Ub1r7jJf1iW
gy9LCJrvzREL/d5V7f0ZPw44MrG1iuDFK+wQY0UbeeAwQLfS3h+qnEkzhcM6xOt+
vh7yBy2c+PMIiN2CErEWNVfE2gmCDb2UB7QrCuXVP1zygFE1ee/Q8FvoNJamIuR5
KMSGkODBSzBaGo4dTf5VWECjdjWmD7yja2VshAqieGmiNWmC7ApUthh1nfex29Qs
blRXGENhULQarSiOGZM4nAjnPcHxgMJ/rzR6D7lj0E5nPe7DSanb0rDyn90oCYyj
1hvZG6vJbTgbhh8W4ujJp/6arsU7EJbJ0B3DiUdteTxwuFwfVeQKiccEYXjw3wIt
AMB8kmi2gNGFGo30EXDnjcXDAGCfeOEUbse0HdOnkZl03gi1TsGZ4xdLMseI0Amj
+co/IvVFtFVJS/Vfb5ISB634TT6ApCgw06gc4hA8Xio0xi6+5BT2o1bIDdOOqqMC
azvEreiFdj4JZOaAlYglpxZysD1SXGEXRpIwib5FN+NTseI11e7IhD72BsHdpA9A
PJHV82NCwzyllWIKwitkJqUCKODoc4CTZv2LQeI7iSdVvKu5rgOpRxMAF+o9YjlM
7Uk91VXcngX/7ZA3+vSzV+wl2p+KLijqc9c45HOTjdAcIV3epoAF+n4RIEwQXHbC
plAmtp58R7uPuQrgSGnfYPHGcJK1iOfnsRQaHvw7XcuFFTzCXulIPPjm3HZJI55n
HT1F9AD9eNUdXEWeRNuwGEvbgUk1WolJzQTCyz9sBOJVJVMaJJ3RfGkCDj4SNH3s
MT5xzr8Lv+tT06GKpoYTFM24zrGVO+p6p67p+1ayc6TCizJgLzLcCV459MDSADZE
`protect END_PROTECTED
