`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TuI5jvF/d7Du/jkjtHCeLU4+Lloc0SXa4Do5wpnS1VD1oGBT55zseeB+gp1mBZJo
jyon/Jjps9x8vR4nDye2zUdRcL5YpYhYl1HdGv/tYIoRPyLpbQfVUc9BIdy6yuMi
mS4wgvGt8pEPYBMzI6AAanlG+9HlyhHTBx6A+DnFxHtUsiuvTB3CDJjvWHzKgbWD
0qKHC2DBZ60F5eOd4p+uPCJwY6xITGd90uGNXgNZwV59lpXCU2Dj5KZRto3P7QIy
3OLXqCjDO9nPi6ELFOx0FHm/ekIbVlmCCcHyuW6pIjCBfksvw8PB1YzVQdu1nvQD
XbzsofJUt+dmue9k0muvTCzQ9zmR51zVgQrXXHkrjRheSzTxcfqZv2LmvQu0gq8c
UdGh1+t0ow9SUZDD2v7605WZSTOc8Dyd3ZzAEg8jaRAdBBlq2wqTNFI10d1hhopL
Q9OsfDzZ0z5m07pLlynXV7J4lSE1cVwxfYbPlDaeqFZzf9zruPhAQ1Q37YMTVNJq
DhnzDxh40IT1o8wHNn8TUoOtiDTy1/nczZAbPhrkRAJovobaSZQo5OqNTcmBGpg6
mmaahh8IwDR9qldedGzh1NKoDnM5p2bhf59OkrgG0JGgaBVO5gq5vn7/3+OTIpWp
wetEcLbwNLSETEbkIXrHN9kdRcfKqyFbA/1ltZzrVXeRj+/aMReNAyKsQIGCNrBc
ojd8x17cp6XUen18RAk4ERTjV5ljISSSTbG/cSkvurtRyLx7KZ+zwgcvqTBTypms
j4bzMmXumrJk4jp8siuLnlGgB7DIXxmXRGENFySvpWvVpdtix3YaJU9IHEZaaOOH
IZ1RG2G6gbCowB5wty/cvA==
`protect END_PROTECTED
