`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OrUZivz9uDJ+p17O5DQ3+pSrZPgizQtJ6Omt2eisnSBdrDRcRnsU6UReIS2iKxR
IxsXZh0YIEPn+8HySvE7gprBjRiWX6JxUY+sUwhI1bsgJFkL+RgFBeJedRTDmI0l
bEE3eW3v5V6qhPUWJVucsL/VCDJP7I4dYVgra2A6o4MDk9Jkt1TMgBWEzW19n/KC
SQhGlANQKIsNWrdJFoyjWxIzkmf9a3fzhwYvDc9xXy2ilPiwALM/74xdvKUSBQDL
Tis6Twf1DQCRfSyaRPY525Hv2B/wfq7edWCajBr3dKlZfGGYrcMpq8HMYVvTtXQj
USBAXlgZl78pZPb6IoGk72TkAQVMOIkJBnSRt8gWi3pmL4qu2u0DWhEqXCjaosAi
av06e34QdTXNV1U6ApfKcJ/QMUPsBMgwKum5PH0DDM/9VmVapqDELsc+n+GRHtZL
wbDncDLq/3YBOlgUx3Bq/myKRweT7ZPQf0GqI7S9CdERl64q5D3RnNdzmgd82vco
Efl+SkjVfktRrWgIPnK+u7g+htrJ+hsq431QDpPClbm3xMqftTCBkZeCc/W7W18T
WXpMeGugv0kmHyR6jrdN0kYxmGgquOawPGjeFNh94iS60F0Jbtlk1u9VhJ55xpEh
T86R3YvhhPtR3d+/YqcpfmsiXUpQ9Nn9N4ekdOZ07iOfZX2Je7TfRJ6PRH3Ucjb+
EfWSZ+GgVXJfjVLJOFbttlC4esyyYOtXfHNdStvIaXazJhH61I7OiVG6ughsu3Lb
U6LQKl2mmN5DdCqTv6TA1yF8YNJfbb1U6GdbjzL7TPT+NNUa+vVqGLp+Gg7XS6L1
C6rkZ4mYbs8N9Tf64/zxnR9qr2GW4PT3EyNSX4mf2nJS9wUlFS+hFriFPcE+FBRe
GhXqjfaNNoB2bPiROerfxi91u7ckY5xzdq30Rc7ZxrwADazjA2pG0MlnI2Yuxmyf
pwngFzJiw+R3kwDU3y9A1Q==
`protect END_PROTECTED
