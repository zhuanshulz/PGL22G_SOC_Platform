`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GHmnzLL1tPtNKqLz1vxOeh6UmxRaziM6AdpDD3b2jSAojr4gfHz4ksJtR5F+9Sl
6I8YiQjALConGO7jHaBD+zUOC2GTt4xmmf5AXWSHZv0yRIZTWA+jCn8RGNMR6Lkg
TH08QFyrNcnYGD9ruI8+W4K7DIX4THUr1+d+MTpJX/rFSDZo/Kay9Awt/9OOXjal
Zlo8yjE1gG7OvCLxDVEDzvLZM6BBUcunlCrGT/gOjnf29tJjUO/Tf5+eHwlS5IT3
o5QbmPz5C/o/l50ezO4I43pZDPNMLRTPtsNZPzi+WPrGN3cYaoQOP7zy8UrkYzrj
tp7qIf/K4Gw72gBN9OB4tQQWTYuaAChqR18Ht2kGguRhrJIJNlX1XJ108UeZIdqo
zeQ3RghIAitbtdv4d7f1IeG7wYsubCjjep1RzeJobwhqX69IomvIgr4xkYUzjdiY
UCCayLr/RNlEZOZwQgsCt0NCpaYLPOcz7hyb0mfCbvI2XLljNH64o3Cj2mBYRV6x
11/RNdM+fedMg8y0iG2qBfNDB7Ir3deusyFheB3mCzENCAypQm8tGyayw1aFUsEt
5JnAvZ2Y3EsOjK2pglve8GHb9h/b3oeyNq0EeDRaABZk0Y60X3inFvqG36nk6fxq
X05qMoIEbH4jrEEZ74vvvs+xPWDCZ0FEBJY/bSestvAWHEc4+1MfI5wnb4Cq6X0j
Zzuq6STdpZpKGdZGE5VGjre1PKfuaRuhcsgB3CyiFRi8GFFGoHLej3v8+3SEwJXe
MxLC/D2Ckp2jynQ7KciDpMMIldb3Go7p1N/HrhXdJK2RUawGZTkg09zqsDpUrJTZ
xsBGVVTLT9vrb1KAP6k0+ynd6WreUPI8PWsPBqZ+qnXppIXcRCzth9VZzVyEdYK4
qbd6Qg5JmWiZ4Bzw4Q0WAQ==
`protect END_PROTECTED
