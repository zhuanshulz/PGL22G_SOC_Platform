`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrWLcDO1oiWQTtelj2qVkc3y3V/tFYRoCZy1g61YFdmUg5TIodXcWYgFR1t9TVvk
UvvHP+rgMGkDGbjcFFt9K9fmxeSC2otFz+3G1D5L5LnwwtwQK4MK2JoBVMVTeg4H
t1JJRrnANWkBoCsjYlGQzi1EZeiVLo/DYqmhiOllrYrrEiSLHNTaK8ZBCs8q74fs
41HBCvESibdZ66H+ab1FLWY48wOR8sYBHpyfY5WS2fPLr51PsS7/EjIQIERoGJdC
63CxBx5X/9z8Atzv3Z71zYqw+9P1PyUfWHGMCEiNE+Mvd6/Hg1fRB7+uvxAJe2B6
XGaNxEuWXsMq+V0i5C7SpJq8lmIuRHk2jeaTo/oo+gmZGRaXsEKkIryB7x8JM7r7
2KhTGnvvhDUVEkL8VErIW4VpaA4FhSMXbkrX2t7me83bwOceQy4rgJP5QdB/jYL2
5z7jVMViMQt1Pvn8TAbmE/Gl/zlHmenG52AcwcBdJV86rppkT6HOpZZ8UscpR6f6
8m8a6ji+JDa/MjwStSJzLNqyUqDOJC8mwYObs68TUxwJSc8Rs8bjZ0J/4HJ+9YVN
Af6Ebcy740tZqzdb+Su8utVHdgjZhqvpMJt1bayHI5zwaSwXr0UgSuWuYasmVW8N
0tLs3gz0VvAqohOCFtf1k1k9AW0UkTQvAR2GUrWEmZ4jJBZiWGOudX4TdeHXaRLm
YTjbdzqV7uFyTtXHT17gwa/fvUzKBDmVjWr8kRSDalMe5L9J9B3Jar9fmQDZsvOr
yalXjylFJX/i8xi4qFQKU7BuIHX/5sNPkU1H3lgOQv+Hj7hDtWAo2gY6KqmPQqHj
9gP1G/T+gOdaDX+G9Eq4YR1cDm62mQ+bdWqYMLzQeB4RLfiC7CJ9q2QkyfhrOxgY
9xzMAea/a81hdi/BmljOTxOVBeo3U43DhkZfvWnmbmJ+kVBOCp7BEKv1IRJk0rfO
0gBVpylNq5liNUM+3MPtXTV6I+r95wm6FnCq+xsaizcRUTbD04M19lbPQNj1DBSb
f5NWrborkrxgmtQPAThtJXkHURmIrXCa4Fj8zhzLEJe6DVjpVSFR+zEl72pOdusK
tNg+BVuCCGHjmplwbWDEYa1NAbxTQSe6OHU7dkFNofiHaCHpEfb1ySVX4ta7s5VI
qv35wX3onOj0TCIz2TEDlcIjpnTKTEM0b23WWC2tuaw=
`protect END_PROTECTED
