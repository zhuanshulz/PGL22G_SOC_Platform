`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5RE7bpyjdVu3VC/VLK4AFBJOJt1uQ312evhFw8A9mlihdjI9WLwJW9+f69hCbODk
CJ+lk6zKLyPr+0i3UfCPqDkjFdY3cBNlypdPW4fkrlcTHG/FpmxFF9Y0E3AnNZbA
7EuBHYR33XRpKVCij03l9IKa3MGV9vyLlQ38pTpKPs7iXN9+r5mKuvfbEgCLR8/z
bmewxMXHl0URSW21kcv8oQdf3H0hbW+w1eh5zCiNKNA3BbWPR/XA68N0twVsaVl1
y8dDCUKgT5sLUMceACsNPh+MZD2QQCjP/m6e50HomPQmy/9+qtqmliPNxxcAXluB
X7HP/I/NW3XaPa9eCZ4an4Zz1RD4nTQGA0SI3ukN6oaElmL3wTpuTi/OXgZkTy7C
9hY3jTqcHssVnMrJeX57gKVc25d1ueVcZXmbOwgP8Q6KRNn0+UDrPpl4by3YG6E/
wXNbSW0e8ixvynJeDjh+jRn9HYnaLCkbuBmAbf/+h4FuFa1G/gtKjGGzQM/1ssZ+
iyVuWv4DZy/ksVPMQupxBXYsKlzJu9hhxlvwFkqb70v8zke6QGyeNU/ksUB/TEb9
Y7oiihHLNNmtUBOMwUZxkecImQdgKcwb4fI/R4Y/VhDzMbTBvHRIKUrLaL0AeRcw
njZvBUQQ3gTR9Q3aE3W1IN9w7vmi0ep5c73C7hfmCl7C+5GWbifAaoJTloA8Gzzq
nexurILQQ2VLLnxL6RJHrkvksHODgS+wocXHbLgE5I94QHV9oXjJBAgDpbuD1z9r
YGZMhbOZMI5mM2BDtmdp+U2+B/GO2+KBqabk648IBqIyM++8SiRmgySoReuzWzeJ
Qq+rTspmUzB697xf4LrVR7nYXqSBKVIlkoQWjt4TI6km5xbruPCa4xUogK8L1221
vl4hcY12Q5TfxwbKJ7bqNNNq8ecPFUrSUurO6lxWLPMpuCIRMtSJyB+WreyzNRkJ
kirJY/GU8Yy9q2Fczj1SHBP12IRPfaCvwOmKsJY60hsOurosSwYhR5MyOmdRDLCr
Ya4CKs91yBGDWqfVWaX0Zn1KYrKKFL8EsSD8cQNRSAys673nnDZE8GrhcViaQF97
miRf+WtVNhxOGGiiM/wTNhkGT6NmAnxmhvpLqOAjR7C7xWkUDlhP8CeVAQeW2Ubo
A7IckWwOGtg4p58j86UFap3rYfTx8Xml4OZ1aABdEhj7Skj8EMzo9OYieYnIAEX9
lnUkFS+V5jpfK/dNmoZvn6QS6werJO2CrDF8wr1rS5nhtBR5P2PdoZNIQ5Snl2oy
/xZ7xwlfPu0O5CtGzqDknf7QaBpbOyZShB670j1kO7KO3a/HlXI4bHfDXXo4P1Q+
PLBfo1MYTc7dgTlOCJLtsDits+PNq+uPih7kaQyVCNVvfgZpuHlsRocoNnX7t2je
uMZxitVVCWfrSnnOqnv3Sv5QIZ1UDVOhDooHhjarVpKIz/qbD/XhGOOciYTqPK4b
ZpjohZ5KGRAZZ6I3KqRF9lyHcnBtLL93aeohe5eMMMWEfHr3CuP82nS2sFXYkri8
cg/W6NWEedY0gxTOdTzBbJjcGkw9gfZqrEXvDsCIYh/weharihsgXLkmmzeqC2wi
Sw1vtnp7j5HJVCbvGj4RpcGPVtwpKNDIVxmsgXP+v7l9B2xJ61+svez+q2mvAQjb
SHaZOewmrvKCNkq29q1eWVpxWHt4ys4LWQffb/zY1y/6T6VxM8GTOFtQnKcKHbIW
nzo/3BZEcKfMidYqLwCXgbhPTN26X+OWvTusC462rN+ekkdS7PTE694mjboR2i8B
jlju5J983QOTHswB/UbxlMiEjVbHdQiTaLw1Lp/poLrNNLErHp6tKnjDT2zcj/SZ
Tpn3TQG5nyLOef7NHrYXsJ8fd+WuaSkUf5CdqUtxprQrtrVCQkBEg61IN9oK24/D
yyO0N46CbfsYfK/DTTv/9pg1/DeMZoeZw/GOEajzK7lqdOkwKh5I9dlg3YIJf5P9
iB4YinZ9C+hAeLeZbVQklQw4Vq3auU9TpdXE6JIUuo6Lfgjkp7Jdpkf4luWyy9LW
56t1WSbrDHIgG7fYgtimfvgINweNHgSfmn6TsL3Ig2EnQq1AABAqSvlzIeHwRgF1
IKd+DAM3d5QEBUIoKyagDNe1pv0yzViTgT2ZWNS6riN7BXyjbkmvgmv8nGxQdWRx
1tGo3ai1TtG3IEVPmqK43TiGO+U+fXtNsBU9b4F5Y2YjoEGa9w6dkmhZFMqu/TgW
h6GrUAYeVUQdGaj6gSHkImFgfhZhEWNbvtZgcZk87ZSpZtn5DMap1/PYG+G0aimo
7ADyTs752y2kduu7Q3TLBBwQkdbUKMCPrMiLiWfwPX2JldgDfj/sOF/hMWeTMAEA
AeA2mbKQUJDh31KP7kvaxcxzmRM5YYc1+bAUGbpV+DAVl2s1BMggzdcuTPeseaQ+
+XC9FBS+oMvOuaNvipZA4iSm/qPONwapc2PcGglu5DFV551zBHIkh2O/W3SLDwZ7
EIA8YWnDgvCcC1HuO77b4w3zkzTtUTkry9DX6JVZLvWOcOsXvDONHkYjCrOCVhd9
wbo8NibaQJ8djT/Ke/x9Fx0uhgjBGv+liS9Eu51H+73S6lYj9jN+q6QxcIhudfdx
nBzeHa+iYMOueA+ZWHCfTqZbBu+vtsDsPpF/8rF1j61mVk5jbnD06OOG9C8KO3SI
TP1fIK8S9hg9Ime3iuIZBP4kXr7vFaYO+OVW6p04///nDEpVa+LZJRk3Vd3EPyoE
XbfO06zOFZGL78RiXbqKI88XOCpwuvsgZQPuXG7VcJ50xosO2TxewL4cHvs7WPyp
v/WX0xdMqzVQhk0+v7n8XUoyXWbjS8aXRNt/8V2/YaXgGKTWUkeLbZ5pNjl5rizO
+WoEvDXwvkmGF36HcPFRMxKmFCuAQKFVxk0UqnQw+Ii60XTJagC5XHTU4lEYPRDW
7C05qkjLVMbyovUCvIbI8J71VSmxCN+I/j7r706VSNGHiYjJLhChaWpaf8xO0l+X
Qif6CfplOjLxAiZ5iumSgHhLYKWtyKZq23XCNxvQOFgFOb2MzUtN0FNCrMTx2ceY
JmPFhabJEGOeVABaCRYOB38l04icW4TsVln5syDdhk0g/t3RpSdXlSfxsiIcLSmc
iWOIygRgpbsUML7FAkoktOBSVXmBtniNTsiiFR2UhBp9qAKMatplwVllitqG9fXf
+L6+dAVaTzqQqcBUN3Mti69ZRhYb0itZ4+EoDHuUAUCRPscecgJ/4N+jXQZPz6jV
yBj3yy/91eDi26NoS7YX41iCrid1z8x+Ec1HBsV3mA859jQ1Lqh/pLRIrWfVO3oF
eDQ4yBMs7Mwy7W3I/B26ax7Eau9LO5h6xZZbX1PAb5xvg4E7PWVZILPcCddznucR
A/Z3Q2LFH5u03LrsvFEUgKZVOo7H934ioJMON/u4PbnajS+s58j7jF1T6wh2STW8
UmSC/jVe8Tufv2aFL57tPdNkFDQnC4RtOY3U98jrfiP53PmdQs6KktTNgfMOgApQ
CYrpifly207lJob/gj6vDIks2h2igUakuZI/NKSodMMrHTEW2iybmsBzNqiySJ98
HvgKzzkNgxCTXWVagon5YYIb0KZ6N8Jjeq/6pD3hSxZh3HAKKNv2DCLMfdB7VuVi
tFN0nOwHwX6IUGT3HmU0vt0rM4Bi0Zv2UfjSm6wCMbttSZpHSA/ehWkzGHWS20OP
zuUuCoAZlizstYsJSzuDDeXfb9d/Wl7ic76pg28HYRXwl3o7Dxd3jX/bLchK+hHD
FkSVC7nhxdda9ZczEIl0PtYMOmnF9XbhwO2b4JD4CnyGi6YeGAU+B52YJBRL1P0X
fV2dUmZDdJ5Oq9TakgbwB31Z4rZsSzG6NKjlTZE3t8Tlt6RNVEtIATBDB2ZeNsnR
sLGJx+RTfMQrt6xXoytbVTVzpQqzV4nF/m5qcteQgRUuayympz84+s3VDoJ+isLe
YG+i/4U1/IpwUugl+PoPF+/kJQrbTzfPOKILvllbf7Q5RdnuB15S0UFcJviJPXLb
1UUtw1Ggp8p94YtcGE4ftAtWqYW9lJ+c0FGlF6c4iZ3cYRdOrTcAFhjg3vl3chwV
FXE3TRM21c+bzGS1drsifLle5Inz7zA49Fu5PuodXrb+e53T1u9SSdaOCYVReDNl
WUWPbxckWLJIblQouHKOKtlQWDPeEr/aTlOt0TEa37Tysu3MdCRL1SRyBEuC0azq
ye7LvVnkKbRkg6irWTIjpuTRNBb1mxEyVHTqYOgXlWUlxx9ZdP6ay/CeA4F+K9Cc
EwN5CHYDxvJOh2qoLIdpoLC3STMHqGDitd8DYB9ZGqbNh+LQkzFydzrEF1DIbd2e
9KlnUmmsn/+KcafQNnIxleDRLJzK5Nu5PuDavQGlD8w2gFDx0/FwAZfv4FlhU/Pz
8nSzvLOUn7ylQ9BNjXHLzIOUyp5pM36WhOGHYee85EN9pv+yA+sY5ffZU6P6Xc6d
nIPQXLws79h15K3c3rud6mJ/tBUyCxwBXJHOwP0iUM3vjqWjBWaskmbx27FcraPW
lJWl0MVIq/8fW6KO4PA+0ue8i/KmjH4y1cogjarJSlJXDIzwQ0lVRsZQapM65ruK
iftie7ubpNcoqlZPoWJrxQsKp/Q+5bdHlR/FIf5MY8wjn/NItWRjOudCLcNqIZ6C
vrwzztwsgPtNkBQKj19VaubhF5kfd50cGT7SUJeiBBIAOaoE7LmTKoDjHFuj8+rN
TOSOH8KlLaR6DNxv94BWe0Wtw3/muLonV0UCKIpu+KdEywhcnriQF8zS0gv7EZEP
yvzTsCMT22h57xtqRjII+uQxYBEXqeB6X20KCF0l4iOTEAtG8BoOB+fKjtidZWaU
TlvZm1TsPLnEh1HFfbgx2gjdzJRBJJPD5gZiCqWFTZlhGRoMP037aUrIt5Y2L/Ot
1aMo8DAlkGuSssi+FEpSUHdxzXYPyzCeUSHldoaX/k29dfz5BoMlYVBBouBzCJuq
bi+983a1q0r8L0E9Sk0SCumbuwVNewUNYnp1rlky4CLHx2qXt52cDmsm6oG9qFOq
L5zkWY46+5ndDYaTGOrV/Oigc/cQNTggWOUIu3tfHG5Z0eDvnitzDvQUhtXnyf7y
K8RWak7w+gAi2H+MO3dkNu+/p/7Y7st7LBj6KXxwZ0KltZQxtz/61rmLYiite4kV
sxyPySMVldvyS9V4ZbGvNKzkFWiQzD6E92K0qJZs8zR4uDM8ZlRr3dyDgbWAxJJc
hSAuKz4XVfsRrjQLSEAECjrSJzafsmUHfv09JTwKJXj3xbC2nw+7tDXxXiFwRA1y
Wne/33t3HJuBfkkubjcIvURdlawOjTj4ThOuWF4uUPfKLCPAEWE/0K2QHZN9h1D5
Izwp6kT9EmEuI1sXzouD3mr5Pis5I/VLuY7UpVf7VBdgz7PJT+q+C7Yy0r30yuaF
oY/+6o2z+/Vxpac8j7C4tOplxhF2CJqYOy3b0Snvo7s3V3uzokUiTvjCN5ohbA7K
VYfLZQ/lX5H7POyPbTJL8Q/HEa06rjaXBYOnH66egMWU1L5iNK7YSZtq9b7PXOHr
X2yOHgJ4FKhZ/rM753NlLVN55PhoP4sWVk6bRfY2TNIEhtiE2EagByS0Ai4scQ8+
frd7bhvmtx9W4AKepCUbTVnnBLQvdrO+9c0anerOLS7z9q0vwjQUOstTWVGvkn1P
32DBRwJzptVDeKEywU/Bn3Hi5rEf+5w4keTUs7Wm7IA24/sRTpEPbrM3mNxyEBse
A04zNDJ0tsJFCrLE1SHyU9Yig2MAEN00d0z+suDqeSoF8wGoGZ6bhWF3CeDVJCop
4afY4mndv2I2kbkJeZndZ6wjGcy463+WA0xiLfYe2hKIPJBSBYAKsCRYnLL4he6w
E3lzzRer2bhAwQ37L7HiN9UYe+a4jJd2G9BE6Y0sNrIf9y17ircJxqiUPoM1HjRJ
0XtGALs4Y5ysZE/c6GRkxSTLBnpwbj220nuobyN9O4FdeqHsoeAQzn9Vb2eTPczp
j4DPuOeehkyXFB7XtUKXZ3H+cECRIlb+2hGXG9Dv1czV4vQbyGgfAUmObe/QWs2O
uBRNk0oTDIBRDMCYL0/cC68Grj/u6e2Pa7JxMlvORNuiOG8r0JSckYF/pa7mubQX
z7gQTZ0/TpZ2OWAXOktd6S+rioU2Auz4+KLiZjJHEFOCYlH9kRNqE9C7GErFBLkL
5i5b1k/8FnBMs+WeAFK6geZ8jUDFs11F+016WWZ3V6IzMMBDt8ImNIURgWQ7wYBZ
4xypVqEOoOjkP354+g2Vq323qQuiIDrIA3ZVfbiMOb6CaxDuQfzMbU457GUUecuL
`protect END_PROTECTED
