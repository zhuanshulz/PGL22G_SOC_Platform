`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+Lpqcavtw7n3Og40sRAOGJohCEVLlx6QZfursxjulXELnF6K5iyVmJJOVCwgADu
g9tOcDJiLKvQEhMKA6n+HSi53I2gBq7fHV0J0XA2NTHrRFKRc2BwgQHW9NmXeDiX
tYGMz6SjalgJ5xDPVb4HpyZQZGBE6N3KVSiFhXW2Tw87ivE60BSYnX86Xq1WjKZq
+76B+kczU5BFPIym9YNmviWDuejLZo5pTPAM7CkO5t3lHw47QBpg9jT299WRKxE3
QNslxcFzkE5rBH4xEk14/n8JguVrzB7u17KWdf9f0+VUGOdMj4JAUCTCgrivITgd
bnzLmLC+57NhuIkVtPaBFN8dKfrCABi4juQ16+qesMV9QE/4JxW8mxnAq7+7QmLN
upbaE6U4sVBkrnbDAa6ajqTrxMr5OKCHSFbKGYuyQcuXRC6TX6slchCGCCQvahN3
Rp8Z3KxDblte+a39koe++F1wAfixsbe5A4trFt8gqiHFajAu8brpEQhLb8ZmhKzx
RTQVaM607P/UufcuCTJp0Sm7a03PnE5ZUMeDxUhVRwdQdu0XYbxQUy2LyE8e33WL
`protect END_PROTECTED
