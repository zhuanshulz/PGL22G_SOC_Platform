`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uO4TlkWsbxkcLBr+gIvk7gWp+QkF3g289sI4EGvoe5OvAFxDb/hbfaf5qgBv7rSg
+LL43AGIMolLyqLs48HGEtaMlOnEjbc7PIksZ/y0bokv6r5NoQwYecSFyx0OGgGm
Iz+FyyoTFw4myP2dWAsgMFpse1u5GqYYjtBSA2Q1BXZNJO5le5UvXX/LjVh8QDqs
OL18RBBGhX4OidvGWPDIa6rzckRnGrXXbNdyWs1odIq4Xf8GQk4OLE7QigUB9Dru
rSvMMzBD5wf9OWHPViZCycuMtFNVHRlEmoYu6hNiHxgkVP/XVGCPtFHRgUbAOeSW
FeYvHlHzDulmqGFwlThP91KdcbU6Pr28SwAQoIcSxOWZua8vDqEIm50ko1oFjIjn
SZO+HCfHZ+fvexXl+KhaiB1b0Y+s0d15hDkmgIjDh5OCo47iSiFU4fw4F1XQutp1
o5JXqXatIK8UKfqttpbT6ojPEhE5vgXL1iIkF3YEO2gn3tfrpVknbsaqb1kPSxPy
lb9lqhUU7SzmvL3bkqnufLtOuYrDWacX+H32rpDpSRzGmnMB432QRr1w3jeIoIva
zeo55VCZ2H7yIHEBusaYFsmCkGTmq9/sJ0DgAz7Z3AsKJWuW3XXowiOW5O6aZYGb
`protect END_PROTECTED
