`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrUsUDEMSN4NZVXZnrNSxftiPUZsZWnJsHSpQajPKxvS9ECkAHwU4x3/Y2LXg/qA
FvR0ZkalzpSeShy5KUB5FW2JS1H4n1mOG/+hk8+Josih4PihJqShlUxCzShkY/6a
HEDC+iF912vhdBoGMFmsr9pLN4U2qxyvAZtGQELZfG7x2zDD0LILrM+4Frf/RqBG
PKU02sDoip2iWrfzTflef58aqCZ/T1CGMg+l6HysB41oShuamktI45RzgqVKdyJM
ylZhG7AG6KhyB4KV4XmlIzcCq+NFjMTr81Z0stF5fuutzzfPUMEkGJ7awFEawlJ9
8QeMXWE6CU/MtKuyEfj7tONPHxitdtCVjLsQPvWMX8Tiyo5J1yDlupriQemMXPd+
Euua48retqmfyt90jCSS6X8MK4tYBIafuCCqBD1HHhZBPFRSBwSGhfSEoalTnDXO
FAgUN0v3UUxL1IPawECBSoycCbZJE9mOt9sUOAPWskPbH3T3D+TxqgsYGI3akJaj
m/nDBNq1Y8f61Cf+HnZMh8ljgadc+SUcfggwcbgGzOrgZFlUGDQMkX36MHqkq0Tx
zaLTENXrIGwoQeSdMlmYwtWjSbq8N3LdgBD4s4yiioo6PvevmJsjCohFCVpUq2zM
at1ZG9SQ3239VKk1iSVOjqQSLub9wt/DoBcCfd4PZdljEwjCJcTX8soiLIuRf1jx
HBsV0QDRPhv6+Hv23cGUh5KodM+DF5o2khXAVisvft7sJ4QQt4HddOxY3GXfT0dk
Gza9POggSfSZTpu1YQYAf0GDd/zpwTLOue+8j1qAGOZLIC98UekWaxo+BBH81s7+
CnrF/s0JeDw8gz8F3Sul59qv5awGkLzxzggo84+gEB5XPPHyiOIj6cgcYXGAB59y
RVhWj45z+DsOoXBBghLFaPOIGt2VjZwnYaFBzJ3afTwUceinh04qCv+9lHjEJ8eF
8aYrak6FDPzlPPoTN1REKzsgKjA5mWJdGBLa8RhSzhTcXjGa652ufIh1hGI5w1i3
G8dC7wd4ogycqcBO0cu1r6Xrh1WIKrrFsKY1ER6D0xbxi4SCCODHbEF4i41flcdk
K1zaSQ2FsQ7SW0vQdfQEvnfbR2DqQN3OygG2NwUKQxNPFisx7Wy7lGZMsf2QaYOy
Rw9xlpxodIITy9tLfE35i/2yreBfc1XPp2nZUw8Rc/DWzfGX6UT4/tyiw2fk8cTl
MpiKq27MObqvwEwKsC13MMbERUgPSTeskiNl0M4qGtiF44fnT3/HkMsJbrkEMy5g
4eVcRQtyRs1PxCLCrJrLReCcAaRYMa8hsxwb+vJzBuEJZZVKsXL6EPNZrfAjehcv
qlu4xw3cAxLWhjF2p9SkMsGq3ZhV3xyIPgQ97OfqjPMI2KMWACU7m5lHLoLbVigm
Yi3EFcJ7EJGLokjRGfQZDzZt1CBaQvALd+rU9SvvWMbu1Mwa+tqtTBo9jE5zUmdQ
21tkQ75StuMjn8PFGjZldq5WKjO2aU+Wvr13PkfT1qWRcun2iEXjw1qot+Ky8s1K
DuMyvytAwi/dJr+2TVgYrzo5ip/9MY8cI5LNWVuCHypukp7t+/XLqOUCFtUIpTpn
x/zZQKl+7K8an1t5CaPUdVHGrE/0bXVt6zsVc74nMfN0bLoi/8gMlSyjmBhV1Hv/
lYBN63JTsl/ImSyz1mFJbmBcqpSIzAz7iKWnuoGmPcJr7ydutXvDkAsDagA5Cd8G
L0+DIfvkj+PO/QZvS/AdaBsR39fidibtgsDk4xw3ps1OcStnXJ24qQofDaSeEkCp
ekG2NcKSJDoE3PgA/yewA4SrefNgMoPhHPoohLM22ncRNGYqymUOicnhvj4XGoPK
I+FrIZ4/yM77gocxXVqVghVMVZmjCmUQTJG7Gl6nCHwUgXFRpDiC6kB9Y0dQ2E75
/hLrKucCydR2rWaU/N2bCnzzSCC1kNmzzOTTtgBStxAPiNhy12vH6/mDtft6jOXN
I2pHrUX4Lxn9drW742FqJf+kfV8XjPratNmAiiKa8NBt64Scu2iYcJMxh/rtApF/
+OHz4j7zen41NjNEiGx/q+M+XyxCIXKo1qe5yMzk8cwUBOsmOY36oysFxmNn3ZhO
xopNMV8hOMzo6FfAaxLDeQABleFAzatM0oSqWoI8m5kavB2AN/rxCIg0pmNNqoq6
ks3xGTGFK7A5gSpvb77d0eg/i6f2mmt8BpJLN2Fpa+6fQ+QbctGdo4JatMiz6l+I
IVAQOPcH3a1o+kraVtiaSrgpMzmtR/MGR3lFEWmKkBIPNr/atP5uGEi1lNVeadLn
qQb44AS0cZpENuPBzZvq2HqqSe6Exud/Nx8CmKlHqeRiIbvTYsgfHa5vxvNKrZm6
21d9T7eesgOwO0Ub0gj6iFuYIW1Z79tc1S6BiSs1s+qJE+3HRPKuyGp0QtC6vJ8o
1kxozESBGqI8XZlQU3PbxaiOdK2udXtW9uJMQ0Fb4N+NwH4NLwiv5Oael6N9vp2K
rpJHMWf6M361D/F3wfDqvk3oNSbqQXK0IJ9t97Pe3+SBy4estUmWz8N6L1p4EN7C
tftCIqmhYuyb33od9hZ6+gn2SrfOBvb1XPSa69c5+aDtg2FQQ73GFeRfe5HaYsvo
ORhi4FXHCJYidciwfhB8D7g5FX1bxQiEXkk7aYk0IZMXiyxWAZGBJReW9eWtdANQ
aAzgWBd01nMLjtHqxseQMiCHGZ70Z7/30cn2hJrbrimajDyBR99KKkjGhWoSyVA0
ffEhnKZn990EyfDfRERKTAatFz1nNnCYti57UaEaIaxH16aTSMQG3R7rVetbV2UQ
GY8z7arhfyflc1jMR5j4fbb/Ipzyr5crwbY3VNd2jBMro0qKEen02cCx3avoOtvY
KUF1X4mB9o029sf+RBV2uLT/dn2q09DWFm75Javfwnb3kPIYIqtlJRIHJS91MDMz
JRiFEA5CY9e4zQXIRT3k6zd6ph5U0aSNHCAP/+ESQRlAwSv8pZAziekJL2WjwGco
Tcxs1JJf4hmKf0Mbihnj7bjRWTFq0dC79yXi569WUY4dc0wDAgPqDJ0ESQ2sQYBm
GmG4jEr4vZRcZ/VN/n+Sd6DHP2NqvJstV+CGsVliwE6MvBYgGyLj7brEKJOfg6hQ
ok7cc/VDKvNymxmNrfxn3MlKScG5TNwzjltXQXnwS+dLx/EEXz4NvFCCRHaBjaXL
zEk8TuNNDVWQ4qFL0yDm2Cxle5vzd5IqrVaQTKYffNLYGwCHdCbhkSmyghcQXjvj
fH0w7mVM+mBUcY55INFxsDo2hdfU4Kf46+UZBrZpkQ4zVPUGp40D3VGJyVEwkqZJ
yOA+sMTRz67HjZmae8mjpTof6cx0SbZNVjhzzWopkDhJ71B0Aylm2kWW99hnMovW
iyjp4DKDYZNzz1zz+7FyznY82v2l+KQrV2/UnliX+LYN7squr11YPwcrov2oaJMi
x/6JVSXluhPjQqJBhNT4YVEVEs0hmQ9iabL5fRvqT/bJl+Gjz8HsXo1f8M6/hAIt
4eEwiE00W0y3PulrnUdDxL669cyoUToP58nx6zNgTCt5rLWRBRxK6GvmyPw8xzJV
tME38LbAM6St8H834bOO8bYsLczNGEZf6PLJ3qBauyqBprNTTz/qFcZPBv/N/mDj
q96Njso+qSSIR6K12ml1pJK5vMSntiS+5wy3YVmharv9npKUcKp9xSOzT0Cn2RN/
N6hFl9jBE4GHtg6/L5/SWETS2jLAnlm4NxVnJvAhDK1FSYxaBJ5/236gkciybmSl
WlN1fMgq+AbCqwAQbfXtPEJey5GTNIHlKjaJQoAq4dkMeH+5TgPPnUkVDuazbB7F
eXqM+tu5OBzRTM4ZJNPuiGpEqXzMLPNoKP5B5RgOCHoLB8mIF3OB+wnKhBtQvsLK
0l59J142U1PEoCwtqfupJ8Zu/laz8lWMl4gW9NNwR7wu16zs/1j6AqmcWhKxKi9Q
qrTX9RK4xIsiQbvSIl88UzAPkWmLe+28cqkaETabv2YVsAf/pniTOCQLSSw0qPcy
CwFJdw/OR0ZDstNt1PTMhh12Gx2beSwVyc6dMsoPiMfmzJ9h9LT+uR/s8kB6GuKm
LMDLt+iKb9Izq96L32Y2PgQxreUvzaUoEvJLBHVviFVG8Gs4MwtsEx27d2SR/P1M
VOnv5cCyiQXmT43dfOLxwWBf7asQmm3Dda96OPTTasNi4Lyn4xPqvY7T6+P8oqaw
GhV/wT5qKPrCFniw+NhWlVTNdS1ayZXPkSKYaPJuw/yb+wnQpTy0QkJ7UZaomzQm
bGfgUzXFtvpsV2XTVsRa2IxUM9ZKMCpiDCpcfnyqZsX3e7iRf+b7y02bwPZvJCKX
VA6XyQVxvGIkD6KdjkYjECqdD0QthRcdan40ysLGEXCjCTGAy4OU1ox5FDAt4z55
1WSVwik8KW362iTZMA+XAgwI0KNbANFe+BbvWa6chw5aTaQ/mLVTry2P3bQIkvLs
DhANXDMM6A2MboVtP/M9B8skqVMWekWpMuqCbKSl0Jye1WSbfwB+aQZCSkSb/sLD
kH9I2FHxlSjcmQv8LCoB9T/nXAr9gQcreRFLpGKnWi/Izv4SSWkU+nwmjMiawDKK
ujUH12jOOprDmSIjUlrtg0YMLBYkUTrktlyAcSHXM+QX3FnaHI/Xa05GNJGxhu73
peT9+w7+RYcvhfrS60NhnuGlZegBg1QdZSZPYMGnzDblk1eQu0HcChACKm1yCN+q
VdhE1fFGDLED1vgIS1vKENtYDq3mDKoXuahihI5TpLHfgw/hORKk2B7Yhr8K2u4S
+hon474Fbi2YUe6Adu4hNi4gWRALqMem6CxoNO5EpGgHxU/XuW+X37OoRA1zJnJH
cC0XauzdrjnSvNLOppvxozbWl8kPSWPrHhLGsd42KIejvcaCukXwX1ODifPcsxzv
7raPGlvy2/aSxvotPQexA8GMwFOulHgaMIhcoXRrnXDUNomvVjdmWS+FyzhJb+wn
HDpfyazgYKipS4f9BYvEX/lV4lF5rYTvi+O7hnpOkPrP2eSu31QztXEAjkt1nuIg
p8hJABp4HcZVo7G9D2W+CvxQoHtuNBjgR7FUMhWVGjcVK81gShEWK+c1KeyaXguX
u50u7cTNhp4dsWzW2LQDB+Tvp6AMWYyC8siR9/2e5UDDPy61zIE9N0eAROzFbjTF
l10CbJZvUEzxI25G3n9FRUnQhKO0M/N7m7Fo4gfsNQpTf+zKPVt/QDoqcujja+eC
lTfWSQCQjmUi4pjU/0NtbjPtqdEmuysy7jxlUblO/jcMoYvqTgZJTf5pJjieeN3M
1Pq0obdgBJnUS9mD8Qamg8ET6kic9AbAaAgezWl9zZ3I6Jv5/mJncOj7JeL6LUR0
rcgVyzvTrMbu8spdSy6v+PVCoSrT8RX14QlDsO/YUDBVChSOQ6G6KuSIHloTmQke
LzkdE3rDJ3v90hQMY+HaNf6AxQ8XY5bIgn2tKgw/z4jsUtr9gAkaDhG/v/ZAFqbU
70k2ZOGUAYNvSGi1eQ5fmKERxUqWCCu+iCucMUhGx7ztVj7XnDtUZQ/gwIPVKERs
mQA4VnRBKh5wrmE/wy9kLnkl3uCbrTM6FNs1lfuaCGNY5fHNFJR1D0/yhfqxuqIl
4r7g3gyuP9d9fIvoACUw6jP/fhnwkl4exaD6P1I7gL2XhmSoDw6ih1QK+5WrFQqx
dbRdo/4/vu2Wl9FZkzYkvo1UcOshNRYHb2hqSAik+s/xC59q+lbiDZNd1A0/oT4I
aVzdH8//t7WhnhTmuve60kSinh9pH25vo6/yWpbXDJFAWxSHd3ftyj9GKmQUrwfu
O/3kTxygp0xV7CMdIQbPJlNgYMXgZlPd2Ervgwy56W7eQOgGx03jJ1BqXbx6q1je
T/qFGS3BAJwTdRooPI9LgspXHYpZ1w5VwCdvvIPq2GasVm8GeRVMFDJD72anKYmW
QOjDhHldpWm6xFRpsWt5KUYbklLoLv5LfApmXlslbgAoD6FTaefdUHyGFaiCjUJj
TjI6dT+TbvOrkkPNjg37OEYZZeXAo4cVI3RF2jSVIWxiuBQYEsVylx4JzR8Cl/Wn
Rd/6t4pxDipy6wvEwyuJZRQ8R3NplGbmIPxL6nuqaeWoee4PseZyJOaLE9CMa/Zn
XLZ2inxLbPwDPAx8qY07kVPLxuG7dNp4q74fkbYHyUz/sEGPyZ3JUvovOIb8vt+W
wPhXEFNJ/22LdC4PCj2tgV+B6BrxilybBMugIIxiWDKDp1mH7pWhW0zuSdXcKuAg
s3Csd6cDalaAeN0kWnHOhLaqrLux9o80B7SregCaSLcShzDTIb216LN7vQRXqwUh
uUIGCq6XQkS2MQd9ny64foHXftVIVColEfo7hDn0gMDxQ+Pm6KQs+yfA24MtOO7T
iYf56OPCdx2Z1MuQ3E6srg795vo3L2d1RIN3F1W7n18Jttzp/TH8bRTM2FJ3vuPK
ynoZ21XBWj19QPaSdcmDsdt6RSGp9+BmqFcYfHTy3a7xN/xvet1P7t2KH8UEopfy
+RMfcpH3h9bYWDRQtgjzjKi7Jn/CdqMeLqiEZ6PR8zQ5UlhpTfTgl86l3uIddd4C
SHsss+8SIhFYjCxNVRJu1e7b553mk1Oo/MY1W7ubhR2V4aSXqzlooenvhIafiF0C
LYswGY4xse0Lru7S4KDgp31W7s1pLwZNxmujHipZEbTJFESiBJhtFQU0jooQtz5Z
1y2u4TSe4YrfOxbEv8UlQ5eTg0Xf2vyOx9cAi2/G2OTFY0BM+bTFrHBI/+6go1UB
zxpByfzIS40NknvhYiSUFHMjAZGlLEAFfVspKCoxJ0IUF4gz+enwKfrfA4aO4W/g
mHOzVlz5PIam+LqJDfHxbR8cZJFki0lWr8KU56yj5XxsDrZjagk3p8pR4TB6FXPY
/KOfuU6e9U46VN2q7IsjU6sGvCtRUoXH5ziPAXbsJw7QAjM3QZnqqFAGbFF4Bdcp
aEsnge7U7Mb5HrexjUHMJT+JykzNqmdTvqfQrhW9cVFRWfFju0If0CWf57ewE4dK
rtmJViC99f76K4QbR4Ffkttri3Y+LBYh3wiqC30B7eXHbZ0KnVMjJjoRexWxEDgs
Ku4MzVR8RCIb8kPvgfk1Q9HVcKTCDyvu58QlctFsalL3Fsgz6LkTLIkPIWG2XJWO
+7X3M0kRAtVzAQB+SWU1AHg5yChi7MuV33JxyXJjSei3W2gXuBzyPjbVaX8r34U2
ZE99seZoAXm/+IU6vXoOGhlgav4N8XTOQ+hYtUEH8ExGvDugMWrWI+/wptdSWTaU
ckdVUxKoskkenDY813ygFctLSMRb7qR5/57jIadf+oydOqUcKh84AmIU1s0ShAma
8k0QN36psN7zr+483MJ7i0XLkPCGW4jnpaWjld3Yj1X5aCg88iBnVqrzlbYjw4KQ
qp6+Shd7SOqNMjNyV/wZNgCrPk5W2E20B2dejSiVl6+qB+oo0Ew/z9JFsISNGDR1
x+emM5Prl8iUWIfHtX6dyCngX6dXPrBePnIttlwKRRKo4FpeVkk78sHCdAtB0IbZ
ajOvzlKgG+dxZ10TBfsK5x2XCSnDi+0cZwCQTyKoYS5yxiDTDOAWWyZGNQhAiA96
y0GyHF0boEmXFf1F+W5KEIy9Cvv+RzcWHBhC/BzNVFfYWYuB2UIZ82ivZlUz4wYu
l9yjsg3YkRUCqvrZME9f9cQOZ1PMe2HcLFEB2rsekODvH9mWkMIDc/SfDnxsR5CW
I4HpBxI3gUEQd1MS0WqGYD/rnI0yoIbJlWv+kfDIUbZv6jy/sSpV0SfkdzCKx3xw
wCB91dDDV6M/VqSf/iTIdr8ioUOSrj/90Pmdoh7XSzH0IY2n7eGUk186fMNDFtX7
uhQBkY/7jEiI5xQO5StGI2vwdooxzHc4F5XF8Gd/RMSlegwgD1iJMrqJcn2QOGNz
FBi3H4sCy64ILV6vOmmI7RrAMrXWVcTdTFWEphBsD/VDUpVxb5EU/+pTbnVcOmbM
0uvLCvHwwDzOflLE4iTSqTcBkokaEgEqd1LvAMWzmjVdGhgunrq06chNsqza5FpG
vjhqObK1A5UkkXgFsXGgfX6kNmLOjtsA23sD/THOCxMdf2TU/P64M2huwraVGBCl
/4+eP0G+wWm6CnsInBMZxeQXY3Hx+HzS2K0SQV1JNoZj7xuldKnaiyq18pziHX3A
G4sRVXif16lSef1IxiIerVRMTX9kJEKT53JrH6lxMFmfCxYpReVPnsg5tzLWt2Qb
ENb9CTUv9Chb7gHc/PxMOXVggD3wb45M6ecvt9CVXuuqorgxfzuCWtbf4C6KWe9w
Pte+vnbfzFWggGlsVP5L/c6sB/bjfT26lcyPw0/MZLq37dBCm+qcUjaUa+pBQ9MD
zl0gloqjBj+miuglsH9U+dgvD38vqEEv+NVsnoMK8p9yOEu2HAEyBaQlxKxA+oCa
80Mt10ouPUUEmcfxKDZ2q5ztsB++/al3UH3tmoBClRacVzi9wHq+KLwg3QNgXgR9
pAErvkCz7PrvOFG7W70H5yLXH0BmOTGaO0rEnVmpNysq9CVYxB4NVMNSE+AWnrKi
oaebrzBq5fFt2fcNDpZkj9rU+QbtJCZ3KSM0uZDXC/dhGBrRzpm8GdDFahVnmjNU
c6Bo+gN5LNuA9gYwoNPB++ALCqW4EkZdDsUkWShKtHyhtUOlqjzJ+2aG8JbCjNrU
bY6tXd1Pg65yVIUIHp9yBGQeyjhsUZ8CEdvWLrLoiZqwYNQD+q/3PjZeY0XH9dku
r1jEx5ZNhd1zKWMNhdMZ/mkHIxSbXK6ZLxmc3ECqtQ/HyqAXTVH1Je0Rw04RpGre
yVCtlcmf4CNRiDYfnv8LfuNyaHFOAZyu4T3MVwLBPvt3XafN6H7yf7bR5mPXpN1B
363HSFLF1/KIlWzQ4/ioZzcuLqW5ewhvOI6bbE2qFYCHfaFasYIwZPciP2Ea/ho1
wLYzyOviYIePtEUnHhTZiwRRWS0VP1IOenbpkL4yHOk1zFW88BMSNKnEBWJsHP01
2hNuKRi5Dtmm4M8GCsDzZDkOr6BXab37YOBY7LnuewBUZcgzdp6NFtkcauxNnrRL
Qhlr1WAY4K+ilMylkAIyX+k3h8PP2uxkYcQir028w1hzysWETKmpy+oS5YXMP9TU
CZVs0ncxqHI+laJx8q7WlicJyt6Yfrh8+0p2S4ZSGkX2+JBPmCUa15XqAwa3Vh01
6u80cKQq917THXWjIEOeuZxqZkGM922z3XwoXJPUFiph1EwRZpKz5hchyr6Y2z6O
jaTEjd5FYSN2p0zwFjYilxCzpgGGCVJwV93h94RMtRnZ69k1DZ8v8s/MRAsmisRx
/aihKqPU4nbIbtR+bpTEEiaLTjAyzpYA3bFVN4+H4S3BCT0LRO5xnWsCHY2d7476
YVW5IbEjVNDopvAqTA9roSvTuzMQ1weU85dZZFm6joBYGT5SflODYGqHL/CDbYV9
JqS6CAbDnfxwLZ0dgn4k3ETruMZZrMDVySxfk54EuW0+9oKIMZF2rZ24OGUry0y9
LMSmdIX8plIhzJjzuu4BxvO+xyGIw+P/A4jFgwhIMFFMdhosQMHiCqLb0r1Ll8+3
HnFTtpnPE77D1WiApIyn+ysrF/ZFfC91VB6cRJ5naOa4fuw0Gpo/TAZc2QUww+hZ
liFwU/GZAZE+o6dH93SBazI+ov0/B+dwj02aeHVSiRQkL8P54+2x1cy9P/Qi6TVS
2UYkuK/vq3u8vY5wnfIhxpr0iB9DNfx9QgRD8n3xJtHpR9MqMbO1kytpPJF8hkeB
Ox5mAXSR/3RaRHfdCrFh7NSSkZImCOTldkHcL3SxgI2L6hjMlCJgIXSZQpMzrJoh
LJYhvQp1jTz/W6uLMklI0DhhPViC5SOmbwiTlT5QGOafiHJsJSaEwWi0ucQgEhpY
n0EM+KZlNEWMBBrfDCNTzAkiLhbtvOvXcGVR7ixqNzh3UKr8TgRuocbaf4eR9aY4
uishFLDhwn9VBZl4/ZXKxRunPjL+5vXjZNU8bM2Vv8eGwSgp2LaTW1KXyqUChYCT
v9ELqdcmDQ6QOzpiJk6ga2Uah478e2yvYD0vBvaiNQN3DtFrEGj7WawFYkFhaSJ9
B2LUl/wOhVhDJYYfAmp4kfv5D9UnylNQmaR8ckJJLNSsQX+BDl+2RUzM3EU39fbS
rEB1+19AWQfZDjzkoNwc63/JUG2W+mS0UOUwEMSpLPdB5yyguw4REE961QghQaF3
CStG9cOVRl+HiGIpEwLhxrQu8O7NJvDcVRPK/lPgS7AA0JhsZsQ9ySiuDYayJSZt
7xoN5DLGWXQRgRdDQ+hC1gBkqZn2Ii4sE7uaRcmLUFdQhxRpCwpK9U+AT77IaWXp
tXxPpUwaQ/pRB6OJ2NjzgA==
`protect END_PROTECTED
