`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zm291Ue5GxAgdiWEq4g96nx4I6bzb+dMoBwmG776aiSkD16y/2/a8e42nkoPJOs/
UvUE3kJK1SOzOrT7RfYrb4N+AsPMXGGDbLNQbp3knSv3hgn4Il2DLkvI7ct2jSAq
WvjMaYd4tOB0K3GWEdUEHq048pLUPbySFDZQy9GPoEDd+1QGOsWHKnYnjeRY3qQ8
J8ZpMHSXsirMTT+4ldzP40oHlPfX8Sz+/Hq841NL93DPnMQKjjV7mXt+0norABvl
sUT1KwzmianhFAWjyqYZ7rDk9P+AFuDvjpFE+d9BDQTIKPno83SQiEqcpNHOMLdp
m/TK53e9VwHl+/DCojT8/EP4NVOnWZ8RknGInAI3cZFmZxCBE/zOZC2IoAdXRP+F
LLzSr75qnCPVQ3W4jN5yYIqPRVGke8xBWNFv7aF+CIPCjQgAgu2715PNCOmERqdM
Ypk0/RKuiDG1r206/OX3k6u2aajpJnWU09/NDPo71eTkJM2p3Gkx07PJzmhnt80Y
lfQ5IHVKQfHmTSKHS22KhHGgv/UjC289mOzZP/k0PELlwf5iR5X6L57jEmeFm7KC
WHK5gnTfEhOLo22XD7jresChQ4cOUDjli7UP+BUMKdbItNwxj3qTC4Zn6a5aEIz0
A04xsSu9bzIr35k9j6jfwLSeCZuV5b6yu2vipae4n5YWQanXq1anY3jp5lVQGphg
1M6ILmVW4NQld0aL3yMPqjUVpwMQd0dcViadz3gxcZx5gnn02kZ+wNjVg8aHlb1s
cJ2wYlHZrVw6ZtjzmnoEcqPX6IbnacvRGOG6KlhOUxzJV6ZVZjfgHqWgSNSgUfPe
BOktNdtXiwwntJO4FGZYlb0xTMmXX+dFR02gHCzC/BhwCXYgAeJwYKeNlQEZuYmN
QfZmnFe+uOuM1HBIPIw8q1fNwFcH+2IMQ132pLmBbZESBwzMGXXHmVMvV7fYhnRR
V6nHjtfnKC1+XsJXqiRq/fOEx99Wl9pPeXsWG05i6G9hrFdllYo5X2+Nxwdp0Jy5
SiAewnlwE5na6QQLRYIscslHIVZwVJRuN8g95kXV2z6U55ZItzDcGkUax4+yW0EV
sNgJkmH1nQ8ndcj25kVaNaYZFiK8HCn8zYZLhgjHakI+oL9zJuUz7KzbipIK6BiL
xQG5vBKfJpV2pwp2LarpedoF32hQxIbwj9wR+LMkRlkp6yweTE3/athTCOhDBqV2
bgXdChx/bvCxJ+47nzyOcxQus+5bA6NY00AXUjePYHdWTX2dItRY5dkPyryEO9fM
`protect END_PROTECTED
