`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61sZBuNDUoNytCS02NgL7/mcz2j6chvTx5dTTcuyMSBc/67LH8MQFrZwXXptY/kn
b5sdi6USKCcZo3OynlXcsDzh/Jhza4g1Apqm8XtbXFV8T8IIggG48D4OMXDhT9Sl
FRBgjLZ2qQ4FvhrAjmj0Tnn2hGBuKe430dXk+63siax943ZpRpoaUM8dThNcT/IW
DFJijn100WGJJQDZ8ciR1gTyxXs62WeuUELzyaO4lVlR/t4w9A88DrW32VaeC2lN
/u06vIiA7uPSTP8M/vRcF2C/Re0TxD7EuprSTt4EJ1v0trAuLZHN2GZ/HjAhah8y
zHc9r1TZmoNjr0E0wkxW7Wv3qyFW/rWevKzdBWynPojQmx0UQfy8RlX67Ycw0kSq
s5IsKE3CLD+l7TULabVdF8Pf2MrFOeouKqcxGIc6tcXCb/8dGk56H9XAl6+ca6Qu
3xr66hUOMYUg7d6Z1p/qLd7ZHn7+0kfsgXTPZHLzeoMvYSwGzPVHgN5h71rE+QhJ
QZ6MAFv9jsNkFrL3xJyWlokPy4nlZp7D0E+WQhMDcCKpx7pvRJxzZUDNF+WLB12u
VjOF67YPr2S0Js/Vs0ZqKoN9ZMXheg/XPCIlyiL6HMeE5bgzr3qAcCMl4arop0TW
kme7z3m/um9o9HQxl9xRAyI+Of2zSCKAQkeVvCziJn99rGNIIiuhbIaxmqve9Q4X
m1JyrVg67vAmdMNuE3Q8f4rikFGQW0mLyVReq7EUhGkQHJA9p/KnhA8865MDltA0
DZTdd1tOoKrj2dFZh+MHHBW0n9MhwDse6s5jXjJqR0UwBl2l9Fd94mQEGZlDYU+N
39aSV070TuJi+nraz39qcdYiTO+bsDZfm071QW6IaGW6p0e79XZ5SZwSHrhTuQI6
aoNBc6g4aKa9OTyRzf0Z+ScE2EOgxIO4zQvSL31y12b9EidCUeK8bUz7o0Xg3qGC
3Vbavd8nUCQbMAUZHhBn0U8olAMlfawpmAIoBbTi1VvK/HYHAa5DbhAWmHdcDMTE
oPX5YfIoSHa8NHTmExF6ekj2ax1LcCLAfbYvuUGiRwi63lyqjF4cdCpyeEWx71CR
zNRC6hNZHOQ3nnOr2RIW+P6mhxfKZmuLTDvvTjM+v1AHSUmKnkeH/FOBhZFk/mHy
4kM8DTKhSuCpVlcELLaI0KPpeRQOvyidRQbpCadkQuuMNNLRU97hWUuXMF0zs/0K
1tjPzDMmC2k4rDpyWrH2uF/n2D4uOrmjhRv92yPULMG2iHP/cHWsemtCs0Bcm8tU
W+bIPuIv9ldpcvefklB1vdSG86xpBKgOruKAT03CzsFMuHZIvDjqtOFffK16HOLX
FopxIiYHH2Q0q4j323xndcZKod7j14IVnoUaf4duFFBV2/5FaSLBeFUCMYCICuNg
J6VenZM0RKOvc1qd94qHXZer+yyBnthNcAaSiTL5ACV8An+DKIAQs1uhHT1z29yM
aK6U3oaYI+CTso3BaATeNhSP3H4zJgDyWbqsYEgAFFwNbxCE67mEn1YFp9tgAeHx
qisIBPjfoF9H6KHFTgPBpjdnv4XDJMzhcRzzzZPOvQiFS8U21A+xXXvds4yP2DgH
oELjiUH6z0DJsCEgnum1qWB/OYQs6w5xvVxSU6faMpccdVBrK3YsxZJRlLpcmCHK
axeXhG2mzWGkcbApEyBrT4qTbxJ0Yi/s4PsGcYGhrWz1NayA/hR6Rvt8oXQBb2R7
0ebwi/hh/2fpK5bPgu0o5ucHhnOT6rVaTd3y49gA2VeDfo+39fdzD9AGMcmbXL5o
wN7G1aT89DYKu1M46Xx69zSSF/M5Bl370ZqoUWKRrfQk2GWEpmAYg8qrKQQMzVYU
of2Ho6PZaykWUsbuvXVUGE/BVhlnHWvlj+/MdBqtPZdgOpx3NHXbhLB90fZbKpDo
uIP2du2tCQ16E35/dBS14fL4V6qxyi+txrlf2771RTzJf17ocfA+8yyUotvVoIVL
/9Xvh9jW7GpU6Z7kVHUUnLcIrp+WW1WglxwavvY890GLnETUtgNhYdGbgyTz8xpt
AI3Qx8O3WafTv5uI/g8TttpENX0D5ASjB4Ahd1gcXq/7kPTB5pOZhdzCNStHGuP2
msH0wsTPhZl86x/bt5UE9hzRjYHKsGhXffwf0z+vMb+n8R62GYnzZ1EbudTgarWn
Wv82fUxSvwF7uGfjRbVus+n2KeyXImZmrj/fqcXuM7X5Vhmk1L4HwunL8tmD0hZY
T9yiDHs3VNIWdzU4PtSQq9/r1D2KJVMPCIUlLj6ylbZYtCIPumO0S8rK1sWL40Rq
rT/7OG1QbekS4zqWHtYY8v+I48liQTULqtohyjmk7KLc0pTJlYt3U2P92lNt69eh
3YNWWqiKr7k/GbkHsf1cOV/AKCkwTuc81kmy8Ae/9rJ0YfcbxtEy6lw6DDWf8Om+
U3Nqk2GFKnv5pn3A2hMBxZyhrjj4tL3nYArPjHYnoPM=
`protect END_PROTECTED
