`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zaI6V5MGiUU0+ybM2UxhE8Ltt3Q+FIgYdVW45ScVrrR13eIzrZeyiOX1O0I0QPnW
R3/1V0V7gRKi4TI5nfvDLPVa7Wc0c3ozVbiz4CjMTPMB4dnpRiB64UiBtR9MUhtw
EIf4dFSDi7egsiAfUZJaVFSHfeHHgxH3CzP8vv4suX3llElKOMipI/PGPvuKWaAX
5VUttN6bkx/vdXmnAdsAkr9ONZIgc8hjTmFERbyvt0aL146qZciPLkHiYxBnwAde
UtthGapxn/4zBIVPDB1FkTFWbjthg3EGd3iJNefkVIzdBsiP1XotCR0RdSn8ggYS
naBGrL1i99JTe//DYZy4txWdUcEfLdnoi/BL9Ddv2vcdx5gu9zw5HvLgDpjKHhid
VVEw4hR/S3o/BidFpMmxExKHVlWAHEo7OjR0QKtywQSs8xDTTGCqb7j9jRr/Ds+H
pnItQIgTDI5ltvDw/AAEALntneTsPXm26h7m9nTYTyf0GRe6f9UVynQBG2eUB9VX
f9wKRQ3N16fVqJP4hq7mhTjulcoWInIX/woZ/aFljoJEWZQk4BuL77Bu2JJQHt4z
G7iS32MCrjQdx2aAiQJGiaL09PDW76Z9bC9ecFxUX9MG1aAhuJIzpUs9pJDsDTri
H1KlFXiGlkIMCavPibn2tsOiXxGcHokInL+IPOvwhB3+fRUPpbAkZJd+KXX0jGlB
VRMyk/fKWGL4KzykLpHMQgFI8QoSR1GDRihSIB66qPLF0ofR9knHKh7s5+GBMfm4
L3EETsHtElaL6orQh641Py+IZGvlI3cYDoYpNdvh4XgHX8dRMMa9+iXh0YgSCuv0
uhdrPiYTZs4llttqRzp0B6AzGK3SHBoQncnrKyxnr3nY2F1oxA3lcp2p6kJ5nS+Q
/KKy8lbWpnsbq9WNYbIK9w==
`protect END_PROTECTED
