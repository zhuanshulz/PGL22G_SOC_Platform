`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYQ0xcHtqNVnLsgAEdy4yDpPtfMxEsmGEpg1DTbiPwlYEcuf1SY/wL6ULEnHex1m
jEiRGAyMRwW5HGXTtSeAf1a7MCLiiaq9MBlcWX8lDEfKrcpNU+kYrYi+0rZmEKgP
cb3o1+344s8s0h0M6JYYNsYfAEf6X3CqLdBRZ56cfnBooCUaIILpDiPS3E4Sf5jd
fdeXk210avq7FoLt+4BjZBN0A6BpoOY1Pw/+W0nKHC2foumc0wOiFmws+F1S63cW
8qrmqesuLUdGia4N9Auwz5GDSnHLgeYWegiv6YtuoPKY1X/8Tw9OzPZSOyYLTZO5
Xrc8Q/3kPkJvpL+FqhRhf+8gehiRU0Pqs663UJTmdY5ZYvh8p5ZGEtt6x/+d/n7X
gHP2fa3cI4NRmP0FQkFCKSTkAcdKbdxp4DrdT2ksBCn3fCs/wc/4E6ZU+tnBPka2
3I7ccDSDnT68LHkvAoVRlv0mg09pj2l4yoJYzdaOZfmManrLlsV28qoDXvSs/224
xe5xX8CYr8HQwMTcdSGEFsNMDWWv6JNcXD9H7sanmIxO0oHC2SI/Ztri6sg+3vP+
yw2FlvoARMAzmhP08kiCskcgRZacOurDJYdpPRkO73+41vVhns1HJdm0uj3ZnUb3
7WFKJmP8SZi0mV8jQzgWYROZs5udQd1H5meudd/gXDQ7asPmwEszu8zxy+RWAMz5
6FIeUmTOIpR4Y/lALsMhFciVvCLm2MnjcOsV5jvAyHw7rfFJ+aWvc/7oDTUjH2oX
Qvjye19kdqlSZQyU31B9+TbjGyZtEUH4wT/1l/A/hTUyu5IrDN1dqujSTMHtiyKy
Rj0WJooJK48N/1DZm7ka7pvA/0GaTNz4+O9I/3n13LnXRyglxNb+ZXktUZTNgd8X
x9wLlAFlZGczgWLMnZOT2Kb9wxeiMRfIxGsgDh87HWsBJBNDLkA2Q4Cvm0dATfM9
4pxJHDOvr2rCeL9xbizR9ZFVpG03jntgTYHfJTQp6MZc8QakGKsiTAR+LgveLMIE
bOB7T/VTiSUqwwMB1asuwmckyNWu9fidEUiMkhyd8Os=
`protect END_PROTECTED
