`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeKXi0T2AFcp9YIguUY78Fn3SNwcw+BZccxx9cXAIwAS/FM8/yNa/h5x0TpsP8mJ
x0ZGfGZh6wmwv37EqCPDRWvRJgLNcsdyPAXn8tIs2WDNdgQZC7B5ENO++0qp+cjb
jBH2yCeUVN0kRElyAMrobfz8zS1aKNa/fA2gw0Mj4zk+FbmxlUIi9AqFrH2dEKJa
cpFLDU4Je4jHoD/6NkKsxWF0q+QIOliJKW+njrZfJB4NXDrJOHAjFvrbSDnMjtGz
2/13hWug+i5kFsaV6hV2fmGoTADYSbxwJB+LKKL6JpEbJe6Hn7nIvmfzQgPFngvc
a0LCGissegxNesgZeZXP5x7RlVCM+ozHsjkiyEEy7TPajiQYhHdX3Zh/uSPZAXjO
SzNuEgeER+2s3TZWiVheKfE9kQMl+pMYKKDMzrDcKxlHfTqniulYXGa3o0IKt8cU
cBRiDFOuzsOt6zV1QbKjKsUhT+cesL8C1+vqqwIKuh1PiqAmXfPPk/L1s7DSEqYf
XgA5Vg8NxP4lCFRNkiKyz+qCBcteUjc4O04vLKc3s2dFrzE4ZFM7mJB7q/CCR5E0
ojwo6O1M88EjWSpiTT19gT54jO8GGtMl1E6yDsGcnzgXaBM3wY2AuHyyuG53wRAV
Wr7zLX9jvlQtvUqGWUHLp17XlrjDaCznVkcFNfiO1yrHYVhc5KfiywXMewQtT0Xz
Wa3zOa65XK40T+lAF4PNBA9hlXW789A9g9svpuFLNA727nnOZhKhDrGkkIvj5Ozo
CqgeLOWFHYOAxjZmc1/l9tJsurSVmi1vQow58htmQ8+zJ59ZNp7xd2NhPAG3bgrZ
+n77QJhjaV2Inhq9kvlddDkloPFnT6y3NHF7YCKDMVldoW1K6Yb7A91mR9M6z4wx
4ZwdMPdsnKCwv0KbnrvPgZyW50pL+9FsAlqCpBvRHxxgO32PDkQt3eZqWjKkoGfx
jDsIJcviRbKJF+5PrQV4+sQjurEuOXEJ0Vmv3XT2zjK3YOULZ7Z8RaJjMCew/Zwm
EVKBVV4ytwF5leXw1PpUiCUzY2ioClUI/Wu9Lk+dTRQcGMuwfZshIDb2i9M6lsUx
2pS/IswRqaNUQUMFS3eKR2YNv8FJ2FDAeCbBUIT0dw4cXczXqjcQV/6cz3sIK02j
t+rXg8IAU74rJMNMbmFRiB6TLLsuvJjmcN4YEZxp0E2gw+FqgL/9FRyR1ufkzOrC
MnIvANZPoGr05JQI/06IVE9VDd88NB8v3gV73beMWMfmXPZJQ8PZ2YAxDWL73yPg
s9no8i1YTBEoEFVuLiQjebrZCmE8CZxSzO105wrdvi+lHWdHweKpbbbGIySTSt1V
fGQFpSbVT+k08Lbc54ZPh/GLN+rz3Ez4Y7ZSjmBLZLRDbHGbJ4oLNn95DsbiGYq+
Q6KSJBSRHvBfmfIsu0r8Xq0chGB3rpdsK/zVUb2CGUjA1ZQQklohbt+f2zT75r3N
FJgaTgBmVRulYHJmArmqdvRq3RXZDI48PcNpKe2EWvjuvSe28+3V5FtuhKoMsDoM
MO/cZhhY8+XRxfmnR9/Tkp3BOp2L5o5KpQ2D2qKgnxnfVOxmlm8/QSfdQg5JbYod
akemoU0yhDC9e9Ae45JrzRMonKSZnQolVx2miqwBbu9L5T7f323SeqlgG7rwqeyd
6fFMWVTqS0b6eSzmVRFKyuFOh/bZW7zNnGQO0gb3ZQL3dsSLbJoH1bjIEnlYyyIP
x3aD/MMo0O9IvU693rfaAmcA39HkJeBj1sQfG0TVSGeKHqFdngJ3t3nv3G/OU0ju
bg7YLol2xALawWhtPrZ6YRrUa68ZHnWCYW2CBb8JTk8VC+790DPSxPOAXOVTMDBy
Wx56vJwKvBgxSosHfoH1KMSQLp2MJ333iyZuGJQLKlgsjtZo8Cq8pOQgZgSeFV8E
DI4TsK52s6ZUSZ9Aovu1Z1vKuVXnyRIXweQY2z8ZO6pe+LUftjViTGOYDq5ibcUW
3iOHS12FhZMf9WTgCztsRPkuXe7A1RSXyHaaDkuO01hdnBNyLpwA8GfnHaBfWymS
5NGd5lrw+6UqVya9MwCuCNUJJx0eD7DgJR2BIYcKizyrfy7isjgsxjp/f3r26aoB
YyUwwvCjOdB43UzQ+ilbF8PewzdEcR2L9ex9s+Bb0kOt1Yf4sGP0J0ugTHrgzBEE
eUJH7OpUEW1AgxEWwZYnMr0XX2jZwxoRwvNWHom/fiDPI+6vOEPhnv15jyLmcH2J
p6jfJ67ezXEAO8A+DfGjj0AJQFCCLAOyx9JzCpZx7X5laEnlyy1aH52VHBwyB4xv
IXGQPLKxHumZz8yJit9BT2SQZIKlP10xLpkOgZnEtolRAVTXHl3mwlmtXyBVE82A
PrVHZu/I3eaPWGLbvxtUMJcAD+lGwYYlWUw0NalSG2bZ8FBXvnogEpYRy9taxiOB
0hc1AJHIpRfJ55ZMbz51uK178oYelvv3sZfVPUzhUVpGH/vCEGUdWZauNduBpnO2
LY0Ei+dVy8rfOU7IMDaAMWwKBLbImCBzwXuMoQ1/QUbpXUC3LEaOvJuNOoLoTsV8
HeDzGOq81KoERD0sJqRrqqRJQixYJ+LCwNuTMPZ6hwZLIneydZ7I+2LqI/nJ86Ef
mWybHcHduEuZnsuP0bW8yls01WfwUO/sp39cxHNE7antITZqw+VRzzEEbtO/zUy9
d3XEvf9B8SN84zlbpCKhF40YrieMXQmgOFGgFL+BABbcFPIQXaMtOBsXVKW8NB8k
Ur7WjleXtWk6ACqxETPtGcN+N3aRKJ/ehP2l12LjWtOcz2be0eQPmRT8aa7/1Nxv
JC02qMaWZ/smB4mV8dnNXtQqOQkHU56Re1EK/8RN/ostjU4LavuNL1kSRT1Hm2pC
PV/FsjGfw5zK/O6Yax3k8ODzMuaDZCEjWa84utZYpCY9TLJdY/7d9dhQsAFVmrzC
9Gi3lBRY7RZfEGxDg0O9Vy1yjPi7MiqRVCWQKw3ReyNkWQXgks/R3s9aY9ohQJJV
VOAuW5yMiAUbDUa1x/kEJYJ1SuhzSJAZCH+GeqiuDDIFRlr7oz+amn8mByJuVrGz
utMa64ovS0auqNp8r22zTLIrGOfilKF9zDwSQdJIv8jx9G7/1GSGEdjNiOFVM2zm
F3mfEeq+/JUlVc7Y2JkacYzmgGGfBIbEAgHBEMTeL3KG+ycQp3PhVMj84K5f/+Zd
wLQkslN43tiE5YcooCFIyf9aaGTEUmdlbvtTu0QakYM=
`protect END_PROTECTED
