`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdYiG3gE0xPNJQ6MVg2591uRW66z8qa1wTgv/J9lytr1T7Pmbd5OkFzW9waqGl/z
3+jX1zQCMwoeZHf/SjsENt8plVKoNI+l0fDY6FmK2pTCWfPX+pMgr3uvLvQlRdaf
NBN95EPx7gQTMvapyQEl6PqFLhymrWjpqWW2hLRfnkJ4sSCQNdp1C3dEfltS8z+3
4FW2uhHGvPOP3FMvVo1lmrFILTB4eMPqv5OBdpLw+enbDQEsBxIqoCe1P5kMBYoz
b53v4aa9s7XOXwRRp7b0W2KntYKh/S9DMPVIoWuRKl7DTfcGODFiBphFqhs22qyG
BdkVvaOGdl+VwAVCkkJhbTZaQ4HouKHS9j7RGsYA/CBOTVX/iBtXZ6mCcrLOgOOC
uJI6egZn7EyTEjtSMwBnQAfeDhhvTMl5TRsJyz9dZW42Y99aNaWUPwmBnMbW0Uum
zE6ieJ61H2IAaTTvNvLN1RtFj1puanAA/snUSWtHh4oMiLh3boxQFbtuWUgpd9jZ
aD0t+nsBEP08EcsrtNTC2L5YRrh2YRGkCglDxey7RD4K3xsWtmZ4kFnOZ1/6DL/4
YcWLdL3SWpJOAukUh78tuxiC8k2G+OEFYOoRz9brj3okYfFeHGgO/t9QOmiEurZM
9TISMX0M16kWhX/QFjQlCqpS84Y9en5WKxfbH096Tel+48sJIWxGlG0FkjvqZ2/K
pzQSwcDxS3qnxVafgw/zsL1ALJVZpRDMAv6QQ/lpOEXtRQMQd2wHfQjAZ/ndRqaT
cO2k2aa/P9qZqRSu+YxonkNwKLxql+Iw7RK23L51F7Pg5GPF6cL7aoaevFPDTMkl
S6gLmrCXVIS7sUiWDR+arNTBkByZ0MwPgnr7R2LANM8W0BkZ9YxuzOuKvSNAGeYy
1mYO7E+ksSekVTNKsxz+ZjdRcrdApMUIgw5wEzfaaMsjMNaC7aYmbI5XKE2HmJD3
N0hco7PCuQmHaU5QiypJuenU0V9d+x6muCNafp2hDeXlqpQvDqZX9bowYBk+S+eP
vZgGJcPOVz15b5UDNv4gzO/6eZhrB8qVcSQy/vN/5/kBKu2WEw/5W+2XqrSJ9lVk
nSQiNKTOM9bBNp38DmxoNIX8REMiDSLBOdKaE3GHCAWv+vl/50nJNMei6HFWcCon
0JomEkoa9eeIG/Gx/wfJLlmqGBkisXOM0DZNFxZsr8tCTMgzWENhwY3KtAbji3uv
EvDaWXMWazgNs5xtXhoNjyLTxyNLVZ6sSwRLVrkIMQ0bApXx/siK/65VuupEX1qe
MdEGK4dxC97krncTP+VaS8x1YJOXNacc3vYWQ8uNSIIagDV8M51YSDKlBE+Sg20N
rQgM15axmDuIvb/QOHeS109Vwaz4DrfCkKpKHGPRwSrV8JalPXmP/8nEW8IXABKQ
CKDAJBI8j603wC97Ln/dxrso9CxCYag32W7K3aygtvwka+LKeSCAulNIBpQuSnC9
ag8TF9Cfei+qmCkzlYi8QeNp9U2EoN2wV8aYCeLHiX951QJEXsaBDc8dQCP+84S2
O2LQNs2c53aTpQVP0HNC+OakX2+4SJx7ZgA1QWkadCD1NyR1gVh4aZNGahtq4dw9
wTSlxLkA8hdzEYT6GF6V2g==
`protect END_PROTECTED
