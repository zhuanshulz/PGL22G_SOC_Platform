`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MWp6lbWfoM0knxc4xpxpbsor7FCn5g04HhniQYpe8LWd+5XV9mDu9/qEN2vNR5gM
sGtwTAhC9cDyLy4ftNt1+/vltaFJ7Eoyu2f2IMRtuBFLTcobBgibke3sE87d9iup
+yVynjXi+5J0V59Mj+GYijP0irrHn2nTt1UUhvJvnYMrFVUOVaOF2Wwk2lPlHJnc
cINdahU5v02SI97qfs1PnOf0wzlukFiQ8vz5TZgF38iayGZdccKaZxvKVRDV1kP/
7ea/EC3MfZQoSdbF6wH2fuWwdcYmqRu1+rZpBg3ByraYe3Le3xmtrJwWtvEeiRGR
svixO4CWEw4F+38Q8sEDnGTnir+aykG7MYPh9HvBvdmXNOFteB1w+7ujXejTB3qP
Wi3lAxCojfBH/10V4YsnhxsoPYaP7yG8uRvD+sGZMFPpm803/914cSi9sqDIe7We
cSjBeh0lB9cZGGsPw5PXxGKJJYMysCC0OFN8/gimPcvCEMIpLLnJ2G5HnmOQmOII
rJLSjWOmO9J/y7MOJhF/IXT77ow6rqtwV2FfV256pXXkkZVL33CRKB44AL0Yo7Rr
zhw/C3NBEjlvlXO6KYxmLpbK7JXnlqj+UbEw2u9scoPK5qizpgp5HQ+KdGtgemsG
r4Dbtv1UjYAnWnGRUSjmouOGAa4RIX5SfBajs21c8tOlzaqyJ7k2zml1lUDlRroL
Bt+yGQC5AToBJ2hyvPdNSjPPOj/kyFMGrdVmwO8n7dc=
`protect END_PROTECTED
