`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sW6v4+78WJbikXB7Orw+/XZLMQrjJDglcz3Yh5cVcfhxM441KwXQ+Dx4YC03Y36v
QjA78G19VYUd2IDUAJq/BR31VpeNnaMGe5WteH0wYOLyxTevPHjT8osz+T1TRk1M
wfjvLl11xw3E91TsYmPKWX6eggC922fOZx3aRnhH1g/73znCxr1+ZxxUfhEOwhKH
mpam/2+AzlyDgyFi/fU5xQyUBcxVTvKIOdsnMJdPUo/NjibebtqeBJJYVn54+d9w
M9RpdkT+pvZIrrpFLotnnPdLdYAiiankJR2h4EoajVBErt/7mvu/o4AbRbofjSo8
DeM3snjHyqfxw1V7azOcBQSWzsxes352eWsak0VwCiyAUhy5ECy6+sznRNGiDcoP
XkX6N754gb41ADjOJHfcruMC2o6KvLZW516WasobXYnHCOGBdkUD0eJHQBHKo1pW
YiemJQ2xTh0og3rziJMXWJQuWTOtLrabGmjx6zjSzTIn2PANC9ZV56JNsfc4p11O
o61hncDaaTCvOq1dqp6HuYMU+THB7CTr4wG1M4F5r12bGq6WT7c7ma82Ko00n8eq
G5YLLvl6kOqoTtjCYLoqersr6Z/8N5eMjae5EFhWNEiRarLass9pip+chYJRl4pV
sZIyZMr5ugpm/wXkLicQzxI2bJL1C58a0BgZsNLjfSX5YxtTUJQYym1rzazo8LNr
CGu60yTgIDnmVzjuYz6ZsbZ6uBUIW+27SvS81PgRb8rimPNr0Tq5GbRGlviUxMy2
a9oyreburiznYGO+co/kDJbgrUiLQqYbZDd/rgoQLZutwqcomScsR06ZnpxkqoXK
bfiP4QLaKU5ar/cpZtSJjkhiCGqhWgDJRvX7ETlVfJFMl3Iu0+K5EnMTZcyD+uTN
Rpl+W95SWSp1PcjPqXqN3Tac+wKTNDKKJudX7Y5HNkQBgCFxCiS4oH0NesGf5S7n
+hAgMQT2vBlWYfxoO5faQQSbvvZqfmb/joxp4thv9SEARyj6kPqOGMCA/Ua6wy2p
BSP+SPmfFAd6lHECz5G05wmnHitR0kxBT5s6zatTL99eLFl3BsenexetB586Y5OY
GVoR4ZE+YpwoIKVklhl9IWMgUqFytwT5b6jwLanPFB3oktov5uOmeZA2ZE1AlAIx
H1Sl6k7efX4IDSu+Osiw6aB9e/KqH7VJ4m0uTG6hN4zG6Z69jnejH92SNNP0Lkhg
NW8jT1ZE4kgZUr/Dm0uMA40dZz0c5689T8WMN3Nn52ihxtqZW0Dfaxcq9RlL+tcL
UOBU47UxGRn5TAiNUSV6omT3Otj17KktAlD2I0P8SQuD85EHcLmqZ6Wj+NTC2mq4
XWs1TUAhK6t98cNXvDrkpMdzT6uqYOz3SwuHrcy86KoW1AqF/18FrVa5PYJazrv2
juYtbMP/NulbWFVqMjj0SKukEWlAdGtg6aYSka3DipvrotzPcLWpp+LwrlO50Qy5
odiUf3QdtYOybNg3slCZaeP92fC7+GDJFdzKc8qj7hrHkAflEnOPBay3/x7QtwYV
Pc/vI28DbFTxbBoIckUsfKHGxRyz5X+FdRAdXMO023bvAtX4R0OYZ0kv3I6QVJlF
8MGM8/BnUrdXJomTs+UQ+tX5Fs6GbPUlPhTfQHp5Dv1nTBdG6/DX4SMKPMNrA/gk
h8eecLCN7O6QuIrt9cw9T572/QVf5cPZv4EdhCypXHj6IOEZtm0t8j/2yXfgD/ht
T+pAqOhLV73BsLp8Q+CXEPvS/XuZqOSMMtlqm043bqmQ5PdrBk/fsPTdu94KIO1O
qadCDxwMEs0qgkb6fT4aKWUEHQ3KCkePUf8/W3InqRvTxGF/H/5QCTtQfmtXgJgi
nOFTAFLDjAiqGvYT6oW5yH/FjzxxXS8sNRU3kQoxQAD9jJpEsjUhMAan3LX3hzNm
r5Y6f85bXfNydXuuDUGeObCTHd7v5lzNmh9OWvEygq7QHdNFCXlA6UCz4PF3HaW7
TKS1L/Dzf0DhjRxO2Q5HlaiIF619Bx2kboTQV9T+nsQJpJvlV8iykxfh7FLR3qhi
l0RqaHf1h7q3hePeEpL/Wzn3sJ1okb8VIsH0QsCEjvKpDR9rdgIA4P0qoCK0ogX4
HF7HLEodEfdAacUHkIO6T8jZwzOhhFxTWz4WRIbMeYKNTX3isLJrBp2qOxELHTNP
X/VipZQNsrQv+vDxdtdMzg2sc33ZFvDJpMVpll76SuY+f5WMpK5TBBUriVy5wmN8
ubE/scBqB+/U6gUzxYwiVtgb9syKTPtVjbRkblG2hpBFXd2+50sPfmWfEl9xpOXD
UKYnqa38U1u7+ZpcDNWmqWqPzMLT/jW8Y1a6UJ8kE0lYyAda8Mn+JGq5RQzS4VHZ
YQ9wYBi2jexhfa7iqViiIO8CbOft//Rt8HJ/MzFSHc+nAMp8q53n+8mua6ObA5wj
uL1lUnVBo/TCYDYqJNe7sHcerrAdVePi516E97aHHSmG6T9DSKefZ5X8kHND1Di5
+v4Jwp7q/zYv9iwYEgdl9Dju8NdAuGKVwqKM5c+epPG5dkyiEu0WHshWWZEWzl4q
f/IXPKroyN3LEVpE+UN2Cq2BDLpYo0uiHeGzxFlpVCN+xrGtDmKJc7Acni7mU/GG
0BZNWE+ouJ4b13AamLlJSrKyRSeYUqgLJsqawy//EU2MiIVXohxSogKxj2JhWXhu
c9CFGq+0UNEdEBWRjpsi+OlQ1Pma+U17yyATLz/WkEhR9sbGX7Mld/Hy90MW9O+Y
DW15U4rBSxnYVKtt3Clsi0HBQAxezQe/QlUQ4GBLhFCudihfNtvw980Y/qquj/iu
JXKoPND30bIQ9oiLSw5eXqcqi/LKA5ONG8ruljUORolxJ/Y520kosveyoFNGiI2/
sSf/BgsfJhQGU8ndmWfJNp0miAlhvrjcV/wxUYRL8d78FhMi493PTFIIXzkpsLaE
RQ8FEImqmoArsZdAyI4hzgDyrrBrO5ypwOkkGEJBjKU9Ad9MGWDj+1DlIApSx9CR
xvCDuBGr1BfnljTuljQIBY5tJoJpfD2D58B+J6b92rv2mUxw+TNVjnaGVBVG2o6R
bl6+bd4wqPKdsIDUX43uVqFz116s21TBei/uB3vGH5s61Z9JkP5xp9GCvKiuOy5n
9tB7u5nHBUs4sabUYs7lFBgLo1hjXtdyG0uGwAhQ7601z/YS2WxkPCyqW5DTCEs+
qC+UIzFa6Ne5o1ZIINy9hLkyMYvt6SP5fRQrOqVfVO6C1dLE8uLZEWjGxFwrJoiv
Rq+i1zgfbuXSTPgGZnlromtLC+R3DEObSLV7EoJu9YANl69V5j73GyWCLYUXThE7
FU0ZPuTQnM2aE9mmQUdpEpvR7Ywca6iWNon9A0upIwUJgTGTjL53Zup5q/w+qaQr
rYS5EugBKrncEdIem6rSTddGMbhRcS0O0piGhmVHA9TgzAkg2njJ6ZXjFvjTtPOD
9P0mbDBrHbvHlEjYwLRXJSBoHrejqUtaMREefpciRKaIAx3toJhu8klcQL8NdwNI
QWUfBzC+QoKgM6EPmW3iuNCNknvd+X2gwWn7AhSMi5SBPLunUnlCfg6DjYF7ADM8
bjHh1KaSlOdTqUO0+2j+mzFSj5A+86RVT/6iEbTS2V6e/FwjaaMgIwufWzkbQL4Q
zIetUOGwcSGPlvZh/M0QwhJUXHk/ZDWs3g/2YALELDaZC3wY7fMSu8AoNNsMxISU
gTsNMOroGJhrSkzStl514XKD3IgYL/EU9KLSWSsnlWjyBehHN0vSTDf+rXFDbo2c
yxvo6CoqkQIvflo98P41NpmkXXywaP1BgQ32XAhCE61nSvW6CeTprbIPuiYlHJCH
rO1ur1YTOZZU9Qox4p3Z00C+dSgC3zmrWKjFvxuU4c6BsgtpPVbd9+yLzP3p+gKx
gKJTJJG+2Pihwk/m5tdzG4HqXfZz5oyYUgbFMhX9AcwsWh+uZhZSGDmPb7fCDT3N
g+bD1iefzOeRWYME8XFqA+tQDR7c88ezJDXlIOGEmecNrw7rlffbKV7mBViTojZ3
HkPIYZI5z9qrhcTPs3fUrhCHanmmOFcSk6DyKeg5TBI4btwUWl1GE9GeOYF0KIbp
EsgHtcErX5bS55rr88Yl90NGkO1HKmDpNdxhrVoRf81BxrmU48aeNgR5nfogULQ3
ODnmrTm1wpZJa2IqHOfiWtGY1B2awLTrNDhNZcWSvwRz4U8uofMAsaiubwgaxrzx
9t5TNdPgUUgXFzsprTzWISEtTC1v49zAJZkvw0XU6f8Vh5InulbIbDSFtZDeiwGq
jNcYkxJyeS3B45zsXH0vURDXwsvB3EO1SeK40uAt3hlsp14GhnkkswoB4922Dt46
9jZSGGZuaN1eLkcNhaaWYiildcytFRl96I4hov3UKNrc7wNTNBbFVgd2qrEW3rUn
kFFzX85GpTcw7/g65FvpFtWASb6gROq7k+cLDoD26qVnQb8fTGqCiK5v4e9AZyGQ
cq+cr70x6WPfMZPFuH/JJEe9OE3qDAje6sDxH3UhM7HIIWIi50C3ES8m+nOp6eBv
7JCTxtSQbWDd+3nX6DTQEdig685cjsA5hcAfXTQ1qRpOlb+uEmZIL9emR7XKXNM3
PcYtTNTosbrJYq3Sd0Cvhxj+lHckk26I1hMA1KW/Wu7QQmg6i20Pj/oXvtjS4LJw
vORDZknGNBiAfmLEV3x3WNawH9TFNDekllVgbn+jjjxD7yfk81VpWNWb9YE8j+VA
KLoHflgJOzse1VGBJutFOW8cahqK7c9/ympOXw74Xv2zknw9gsIu8Zpsk/QQ4K8y
HSkvlVpd1SYCMYwsyE9t3sOJjxCWos4K/9GTEFvhu/4ABPzdYdlnEXBoI9TYV4Ue
ZBhxL1QDGAcBiOrFzs1QbrW9zxfZRX/ZYWgNVfM5RDY=
`protect END_PROTECTED
