`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kdrPJzgabr/1mt7yQuZSD59+GhiYJbBg8wxInVZjo/Ot3pL2kPK3F6m5MSchuqAQ
P6T6bNfSkfcBC3pak1idO33dSe3YW7VpiQoPQYTV0Pmgov8h2sv1EiMca6nfDIEa
D3AB94DSzXKonDMkX19ZO1ib5FuGRAqwwn3CLH3q33wIh1sTk0bpN8mWtXu6s2Eh
USedrx4LCF02oa4ihgOud7m6NRUCv8BfnBX26uBCxUFfkNLJ4o8fNhlAeEPjETLi
wD3UIUHfKEM9lSPr6HH9L5B+loRwUa9itCi6SahkS6PekR1u9SldMQZgTFD5SRir
y3zo0Qxpc1o1JMp7Bk6Bd6Pw5PkJV7vj7nrRF/5AtCZFSg21wYek83mEVFFYh+2o
f0LWXYRyI22mCtHy3mpVxLcGnkvN8lcptCy8ysEPE9qcHlTZiGpjOoJlNTpP+giE
Cfb8L7UEHevLnS7M0p2rDh3Q8SN34lEQQnfcXIH5OO7Ukkq6J7W2H5xbRksnF6S1
LFybBCNsLxUB9VmOinegMcY73JoRY2jjDWBAIl3przYA9B9oTLK8zD3RevQ9NTVF
p2qPMYyYbcQUzYH7JQrYqysU+aoqCch4yA3Gn/rnpbUhWoCh+oCK+GUXWhCd/Dr8
laKqwA1wZnmknkpYBKbMvaJmOysMQ4NBp0U0GQlm3NtFMzAhuG9BdaZsjnAisQzp
TDkAon2WtJbBeqaFMFeMw3P5qGMmveJ8PFz8GOHWfdU43yEtllIre6gA8ySE068P
Bv8AzfCIGjifRR3SupBS1XUM7v+fLxqMjxDl+SEWbBhrQg1lRrx/+6aanWfPjTuV
QchnjR1INn5yXZhgk5KbU4wf51jdRe48gbmZudvYBoKI785dZydeqntzXgjaN88y
ZKKK+FaA4dlAmHncmx/47iOXmT0bzRJIcXXJTvG3u9tFL+s11sdkHjnwKv7vZt80
Tn/EB9TxZSF8snAUW7FM95iRoiCN1++CK2bqHdHnKyATGhZXOW+PJmHpAdCEApt3
fpD90td02LTQQ8a0HoyqyGmH3CRYBMy5ROUx20gHPsV1mvcG2z7Mr2zMxz1Zojhm
9btSR4I3t/pi0l+eE+26byI9yfC3DeHSPk+FBKI55osbjtwSD7FvTVPD6cJUtlp3
/qn8zeUxR5Aepo6MHo2iYx7RdXYc/qqPBRraa71C8B96qNOfH94sxRU7i8d920qp
oZMEk7maZeyIk6Jis9G1i8/PBwVH0N6E8iu44uCXBYYTWhKEf5ThwkfzDhW+nXRs
/aVq79gz8rQ2Wt5J9QZJ8fhB+QftFQOCPtO6hvLBw167kDlKANw5lINuva0XT4tQ
qrOTB6cK9UkzAkpNQyo7bP2VJX7t6BnlduMYBeHwQRpOoinhR6i2rQt24QRL+nQq
aFW31HQlfgMBNZUQg5I4NzCDKnxZztH1I/j0xpxJajF7wb9+1MGMoVOZOd1I1QeS
JdmVUZ+JLKwbwym9sdfr4NUudAEmWfVAVZvVUgnEKVPpnMTwokGMSPMDvzAKZD3F
B+n4cEEtFccYmxMGJNod4OUPDnLO4YtsrAbackUZxrD87Tu7lIPT2MSoXgp9Muas
U+QnvLc+jhrBMTN97AuL+Hn/2bIz/XTv5wKtdLGALArT55ELqbyJTkkJsJl4ll7a
3Yce9QdTK95DKJ6l6pYGWiqFz9aUtLUjLW5d6A+Ekbmq4NSs1qsOZkHMz5CK7XSU
b3+2bQiTXcp5BpX3XBPYGr83pWKTj1DpQ7b7bjf5BbyVWyHJE0oS/4NdSx3VZ14U
QqQ5UTJh+nXLZoiCdBpVXRK37v4tR8VFmSxuIuU0wfyI3I1DmEzy0SfuGAtlZsKR
GvcwxIZ4Rh/HOA2X+DFVNhy1NSa6UZO41CvTdm6mf2OwIoHKRCX2noeMzwt7N+OJ
HXT7exoAJtFkDgDly5LOlmuHDrUmV1hmEDLYO7W+Jl4jqgVT0TdY7RICNjFCPXmy
WcoP0+95Il6r0rI9P4CN6B3QuQnRPWRp0OXyg00sWtAiqgp3m0hPzOEWJpT8a1ll
tlk9e1DIJ4okjJWHDf5jVXSeFuKCH2fS2TonmcrmSVP8OvBBXK8Sj5reC7BfjYub
n515ZAnFV2z1kBmi4+U6PpJ/W/WO0ffbK+EdT7JIXJwNtf7U+cJhlPX9gtcBamwI
L+dduNVHyuqL02fCkPC6goKmOxFJyUA20RM/4mYKdprSj4joaCxlhHFmp+k6fY8+
NWinMZ/VFvT8KWq3/gMU1hsX38+PBYbT2Eh6DvfsyY8UBZruHp52JyI7cGsHbAqd
XI2hNR8Ea4XEx+jFZx4PwsjBIiSNxn3Ua4lvqEuom6TF7W0hB5/2p7tqwh1iCNYh
o/2w4O5ZCZomOHQ+HQVscyybMC2Z1zOtQupX193HsgA+Ylr2phQa5KpRY5coZvzx
ugpugnNWZ0gJU/Px/TijZej6KcCgBBqrDREnsDciE+1V9yKVbdjXBwVJm9OjSQ3n
6un+IacNuK//LwBhH62Wn0HBDhrb370ustlPmjpckqbyBU2Pu8xHjnKrPk8NNwfX
1efYW7mOuL9KEKpXC+syeI+wUAWvoNkmvMePsIntX7/EncsWhc5PxpZZ+M8eGLSj
WUrdreLzxMei3+sED+/pi7KlfLMU45usslj6jx/p9f8E66v87uYDVP3lRcXKD7dU
SUD/8g7FxHW+zVOIxoVytt1HDYPUaEONFcTHWDchBS4DXoaovNuRnHI6mmK294HH
Uw9M6Z8h7ud4LMi1KEJdGXkSz+BQZkHdzDpDMhxEq65e1uVBG9JOYi5vBlSz5JaN
4InHgv4xFnqqQHcFVzcv6sryqU8VTD2NDJuc7+TjoP0Y/4UXPQon3RFMd3sUh0a5
JzJ8B9qfpvzt2JYI+kvaF6pQZ+Xc+rlfkpkVVJ6gsFDWYB1ayqBYJglmRvysBOUd
Y5xG1EDmcmBnNbE1f3oGYNfoVntIPBdEfNZ3OWUR7DZUwDu3pLAqA59Cgx0ui/2O
HUci8C84QY3FE3zSY7rFJCOmgf1ZU/Dx11MnJIk+krOfBsIlKTWLxA9XFG6V/Aq2
84OgtvxpLYDqyW+yJajNrsYlFeoc7joyp/p9A4MrmMyTkrA/w8/I9eJeNe/zq4cT
UbplNn3t5HHDHEU0FEzEYULXjibZXh1+/6iXYxffoj8ejJO+6/E0kMi3Zb6Ble8X
5jRNThNJkbmAkWbvJlIGkV1YJMWR11/3k+JgPofSie/Ooed3C1VOt0wPGCOrjhq6
tmh9EPurGykKVFjb9q+L85ofLQ9nsvRLgCHkvAy6FGB5NKD/XpPZ5zQYMYjAVTP6
RwiGgenJp1B3LP2DuLQgnfS3FGjTPlMi0XqH1bT+4aqxttvsbJYWoldgpSvYUSuh
2bLCrtRoGWUcZNeeFW8aPSY4OGmS7GcR7ZYEToxNMl+VzG62YxO/DfSDSaJxJmv9
p+2w6DReEcNbIewFsxNyd/9CcVyozawf9CL2dWEbYaM5ATLNnlKvNdyWCyOqZ9U6
Oo+uiqj5s/abl2LTvf6mC0Owl7hSnkcNIrgcN5thtT7FbPsAkapblAzjGe6Wy0Qg
oLZKD04ZGIxkgsQZGfuZrJltw44e+KXX2FxGueNO7LKRfmBLbdP9vjaP1gT9IJGP
ntW43TJLEeFGd2TgOQLsaUOzfCZ6D9TBBmEjNmTU1+7RSd8EOCdEg1Y4Uqy3c8PH
AfU0iI4hmv1LEEGpJdBW3GykN29CAo0qcQ5/uBGcSHyLRsWuoCT+2QoZpsNUFxTb
APxrCSzu3zCvI3dsLH4L6ss/9h02eemAJ6tKeb1bxuoY4zz1puNGgR1+QUq2Siaw
5vkY00s7TuemPPODDizkmf+Q1PzxnaXFSt1U29AkxDPZe0pPNkEwo3HgBiuBIvan
X39jfz7tj87VhvKg/oGmbWZXun60ZzTuWr3sZr1SyT3+P5Ol60t1glU60vo62Byo
ICvHZ3LSyolIzCWxybt2faMvyQqWR+ivpSwxkJBWM8fdV4S3Du7ao5R/OPGtZe1h
PGSHsM87kAli0dK7GM6q2zc6Krc3Mnd1vfs8YbS0eyu9aPspJhGpE+oCQsrY4hcq
QwLe8tmP8x+uQfcTYvgNMN3zOlglMWrldn9Dxfs61CXcV3Foun0xaToQiCiRfTv/
/WJFQ9ydT9b2+gbQCNqlLTlMlgXKcP07PzcU0jVEoI2SDQgla26cFJIUm/8r4pMT
joPgJBbAWe5klyeh0eSaFeiz2XePz9RW5/Ju396Vti7cnHDvT+uVnKceAJ38ExTI
KYD9c3lF/+ees7hkKgQoATK5Q/B72qI+7tre3rVyMj9xF3t7kTHZwnHWVfYiXCAF
JqvYu0JPUndiLAqj0gIAIskrBMkszz/ta0hJy6wIC/iKT9ziQszwEF2Ew4Ci9kUc
gktBJwd5gTadYrikf3/CvOpi3V9XCNTDBx8909b7Fiuz+qZQs34WWiuVJxYdAba1
WabxrKLB/eXPsFYYqmlZ9ljG3h1zKaQYR9p3hBMe32JGEHhat06caqOfokU+TohF
bfXJfVWVASeUl7R7HllRDaMreZ53NibZkO0zWt4/8j3fwe4suN9kR3UxPWDdu/HR
bBRHux44aRGzrHTWVF8Sktt78vwUEv+a0dxNaVWg3bQav8ZVSMC8bl6rTuR9xiVX
Cmgz2mYquP4tTNLuFwwLB/3drPeRZrMPXp66CkmgF5Z8SAChq2pPtaqBS6yOZr/w
OROVoQjJBFxUS7StnwTw7ABSywmxJuYkangJ40wgv3saoVZOHGkO/DEDTkNH8Nfg
KqQaqY/PPPFggSHX8YgpY7NEOwVIXZ+Tdt+36orVBImRfU38S2ZCkxH3c4qHfG5a
ddgW0JO1CivmsvQ5/GIT0WhE480bfbgpzWFwxBX5dLql/J3EoW4qYVUv51VwhJhC
zPYxgwnbg/mwkbIud1wqewdX1v+3Ka79G63VwCeit+ABljt8aa2WjifI74nd4+LO
xCcKFsKl6ug0rUi+iDdoTm6asWFJmt9SNrn66VIuv7HwpOPdW6s8HV32N9ssvJFP
35C6xjmTqNrjKsuph7KUtt06FCsPSjWnB5kkoWJ21/BQKVUNhkXDfiK7vuP+bk0t
DWdkzS2J6y+zUCqo8/ZobmvZdg262JAk9ve3PCNoONod7+gBJDX1e9pho8Tn94aI
AUgn4inu+FUEXHe/HsSSDLCmqmUpNShleIbPt0QrRQDgmycy6RTzJ6brGqftGcAP
sYGuFBvy/uxGJ3EG1jRe7VbqaNFPN7Eim/91zBKfv17AUD4Pa3/gDaUBh0KXV0xy
hI74jcKfOBm8+CAsNQCpVNzHo6GeKfsngVVGWox1Lad44LCE/4/AxkbzNC9u1tmb
zBh/TP7KV73fsubcbdpl/ysR79E+3K7LI8AR9md0ehX+7PICwR6NTrorSwxXk4KB
df/SrWIKP1MhW+mj6bj8y7j2tzQoQ/MQKYciLHm3fKjREXTpOgTOcYgLCdE4iote
RRigl/QNBMByJ4A1TuTPqogZJkDnxY31ieNcB4h+tbVAehv5Y9ao/VgIZSWDYCGQ
p5hHqUrfueQxh0ch4TbVh8/TjaOOrg8jYOn4v7vJmQ7w/V35hh4fN7FprXEOifYF
VQkp/1IwzQBwnBgbWTqSv0ZfrrfJdE36D5gxHxsP1fK5zUflwvuHvo2AuuRgiwbJ
kgqnrGuuaUkbxOkCsG6ayxVjiYZqU7/a+kH1PH6hgDhuy/yLbohgi8YyW8mi8rAX
96dbZS7Dj3GuN161gqjoHLjJT2r+mzCTYvXQ84twpqWXykDLrshE6ABgLNByV1nr
Ty9HPd5BNIiqTtW0SyO/yN97deXVkuW/6CzQGQdDbTiRpDjK91F2jI5jzcSHo5pm
R3ytwFsJj+AgN9egTWnL3+DXQzWSpgLHXI/sc3QaJNs5+Ah0YfUUREOcugf3ILTP
EvnpZcZ1bt87mtcLb3/quWrIWC8NggSgyzA+TySpwCkoJIB/ljW/Wm8Fj8nGKkNr
fkYw6j3wLtG0FVpToHwA5VBQ6/Le3WVxN+5w0vaWSGFw5+fbFBLW8qtky00MtRaa
yzhtFsy16Pyaajt/G7vYyKCiQ0DVNKAkquUVqCAe0DScyoqDWTLA1QYbxHr8NEeF
QUAKLw9yG7dowQKS7BzoY2anXAC7YFFLwEAgMRKWq6qW53oNmotuyvEm+5GOq+kZ
AJ67CjYr3mpnW+M0+W84CDfpJSTuITFcI5EDiuq55fXPzvQhXzHPRNoF16oOicz9
+5hRXHCIsWRIVPSjGFlV87Y8eDIXJaFnZLnXcaxklJoePZ8WSwxMdtkYkl1TihTa
09yK9lBFhNkEJPZiseVtbhwkdhbYbTgOS9CU+9yUZCoI85JZPPfIXfGmvTjk/lVd
m7s76r6gZTzGOelNTWBMCvykUGkvsbEe7853BHpJOV7ncDN6fGU+BuJTGEEzKlOo
ZRyVRdKvYKX2FhbRLjU+NGwySnf2xLHP9wlkcYBtxeJvzjZ1EBMXroSDJoRotjzG
FputooJanbozVKxJaKyHnkBfX0O/QfjeGraD2fauOgGRou0IJHX4Lx5D9yBGfmfd
NhgAV55DpYTI7JhbhFe1SfYeXiZtqI6iomw7eVe3yosCXXVnnuCVJH9LhChIjshJ
yoICMdGdzEhGW29UuPKUTnj+lkmffe2KtadFMxCVAhFyO2zupvAjXpjtFY8UDy1g
NUQn2Gk0AM8D0qB7Akn9Vey9PQRIf8+uGyn7Aw0PaU4RaBUGpyrAqsbWlyhxrBUh
5Ou4Tv9MhgrNchkPMf2KYvxI5CuEaw2CIgxWfCXL3Iv8wZnBN4WJYJ1KUeLkHiuG
dFPuLD9W+jmh70A7HTlitauoOaSzapbPJdoPPRFj7XPPJv6wHa15ihc4lmBmXwlJ
T+ZpTNWG/4EqiT8wjOV/RCxFnH/cPahHXlCz1Tn1tL0o2YNrYtWJtQNBOvIi/x/z
pbcNxczpfxaofOWTdlCsYbR4gtvkbtyFZPwnpVmV9fQ3rvAvf6E7Q7MMK/YUzRFx
ph5VCK1ZelIecQjgaterKl9B/S6Av5wI2f0//VEevw4wWqKFK69y3lIYDGc/9Va8
oVLChibh2AZ0dFknkjNxukrAPj1lfNrayoBSorzRWAnJxeJ7w3Z1cSE2Ra3l42uZ
JC010Rbq76FX3gA+JzGA+SM3PMwzLXsmysTPddOcFoqImNE2uJVuO/l64mimQ8+j
J89DE1CL9/X8uDITdFEwYujUjHlvAZ35pLzoTtgQAKwLSy4m24KENFcbQ9yNQwfR
GyPkNevhsRfqeGE7c1aNEhuXTf0XZ3EBO4hWEujPjLTSb2GpykX2OLdCN0fJ0Lcs
SyiNnlR+XH9LcxVp1jYzI9TtHxDQ5BhRpBHMA+uaFLFFK8OhU6cWkooso6Lz29QC
EiFDX+UT7WM0/iR5TQu0BOeg0giu3L1QqjLEsBoH02h6Zi7d85UMa9LjCPuoEvmi
2di9csorQXiw3BFcGLSWNJBfjT1zhQ4nXCC069uAlg6wxto+aZkwNcriL1DPByGC
KX1DOc/JGiXPifSkEVmDY7QENprOHSm0C0vAyXZVFPKCiNZh9UcQxor2eF6ybIYV
pi22cC2OfEvlD3JzIfaCAvthsT8RSTbLoKgWt2aNHrE30MUTEISQRcP1opGBXR2K
mt7JmAugyALfWgye8msgsbAKTgfr2A3jq6lo75F5vGLJArXO29lWsEvGr8B4u2z8
gzHOuqYyIz283QMUJIpPEVd3Q1Wm490arBYqPO1HRZiXQnaGcBpck8wd3rkjskEw
mhetDIrQMPkIdk/zMsDVEoNLcYFTDnmUMZd8MxDhyPt2Wx1VQSJbQ9I72dHZzRqz
5pLvFxwyOfgH0fjlaqo6yjKqtgwh7Yz+rMnrWfPqr1TXMag4kCh2BqN+OGzQb11j
PbEtUkYrg59mUDvAeU70wDl4SNUOPdbobw83g1/T1cI0Q9MtFL40sytN2Cr42wZL
HlJfumTc8sAlnq64GbmRBdsEku4XT6lqkvumCBRuGu+DjA1juxUBgaiJnj2IuTNt
`protect END_PROTECTED
