`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a61I6clM2tAw8KubCXx+nINm+UEUfAd53SKyDkD7bk2Vc91rmDxkukCyNZESLngO
Tn0B/KXIj9t8q83c2AlFUkijDa9K9fH3TqFa0NJ8msCTvyexygIhltEIsaYY75ju
4cV02ad5mXaiZMZ2cvpYmu+aa7T/bYACgVIFfyJBYZfp8BeKa9Ou1g60z2tEG0Jt
FvR9wuQw55SIru0AwLMBWaF2Zwb7cTf2XDGADd+cbHvqDbRWQeANjMoCEQ0htfBs
Tc6HnAUemxoK9+DVBdumO5hMU7bH6MdoqmZuk2OEl4nhPg3XXNlGD+IRngD18eT+
a/VyAANshR0yXdRaPRvfHNUFHoQSbqqVYxaG37KkiPE/a27/W4fM78rfy36ZKIZr
vLnwZTiMAOLFFqWHGbcGpUIifcs+Yt9KNNMKTPLo3GkxJelMEV2hqWrTEieLtoba
LmoYJeL4OyAImj3VGawooRim1VX1aGX56CJyJd0RwcvIWp7sRunqBGdNbwN94z6a
N7ywmdOdcDcjkzpz28WIOuJHI4usqUhqjZGL//pokodvv4idHVduzsJRQH5PLZF6
fulGccaYb8QynCAd/iK3U5SCnHxG2O6lJrOxg0Wk0YpT7sd8ekuiL+nggngYegH8
F8D0jgh+wGCEewduQFUWJgcHZcf6WxLzwVlf7G2c0cjPJ2wE8u9j2rgZo1d8YZet
yWXOitfLNZwVPrZV1b/eSsJo2mN8PiAgUfoyitReddyNFOHf2G7spVx3YEo5/AKg
BjMrlvCptt+HRNYI0HOwz0BC2+sE3VDrbnZdrjDSIbov1F+eO2kQCaPbzbJHzOu1
VB0e7nvPqxCSQDmw3tgjJqOe5YKbVT/CGa/apMrrb8JptA8XvrbpY9jAzhhhQydR
nLvSMMcfiWTDRoufCVSuUUJWU4IZIeAsifCGEx7yGvunQ/GGs+saFCQd3KYRTLIc
lb5VulsIGDQLFZszPunDzgLW/vtKz2pjQToHVx6qHQwzzB2KcSO3+9JWmBLZX3R1
ctm8biscz5LWOoNQ0/Y+lICmmITOtmxY4whNE3QI5JrdnYZJdkEzmNU3Y2YHQkD3
SOocvJ2ETw2YqkykT9KsVeC59AD03eqqsbEwG49qKVTBpdTbuj5i0XrGUua3LL74
qSp6Q6BzjPRMpdt9l/jYzpQ0L/PxARKJxnjGDyYpK2lHWGh6gBzChBFpd5EMQ7Zv
W116fl7afcGvgsYn/ON4izoNIZeVmpIciOMc4GS4l/vimsy+NWOGJpYAjVTBj5Hb
nX4nbvXpeiQU0n8rRDwl/BFCc9VTQ6jTcHfQVQiGRKmp220uLusUti8DMNd4Vpa5
KkH66qsbD2niscj8zmvCCTAQ5TssLe2ruzT4jghMGjtCAMu2ee1gsgywnCyfuDTy
QECVbttsTsjwUbsYIV4hH5GwXyBjDg/5pywU0U0oiHVOwzfOTC4UAbu6SqpREgYH
q5IWrJy+ouen1sGNd7XgOQ5Jc2/oXpj4CKkQRMMy0wRbPISar3NFvnRxZCaf3I1n
EJXLgJ1o7+/7ELTjzYOthUphePIE3uGFH3dkRJyaWDsHOb88e7S45Orm97y2XJMy
1LI8ajgwEyonpGNfTqd3wYSRxk5iY2IB/YYyM0aOpUtfF7E64k1rzAb/uw5RsNnC
3zG4tODuEuTCJWJ8b3SeQ43h9i8dA2AZcXSzWSgpSOy9YDnpsTGeGl3UAtLs/UeQ
4164BYxvO6HwYffMRhpc+bbWIKEhiRYpH2M10Hcza7qSOhnXXDX0jmz+nGX8WmJ8
44D+bq6baLsBiD49Xp97BZvTUHuGbBAYednR1N2XjxMq5yztzK49slQq4lOGDtec
ypFUkah/dHQP3vlmwmfDSVOnrtC2PwF/Ms5Cl+GQdMAm0IYH5FKa3GsufInNeMEh
LZ859J18yXSsDlXzNeZ6DyaLwtEfz19uR6Jp/MeQgM+E3+6aOu4Ck9kC5q82jHck
X6Fv8KVouPbG7o3gHIcklYfQYUbLqsgGQRw0TFrTu2CnCAlI8ltYDcJoYE71Txe7
Q9S9c9GizYR/mseeOWdtCWNPecY2y3lwi6uyY9Uq8BJOdqw5k++vYoHANekSSLbg
ngnO8CHnxfxWVb+oBMoeazKDeAfdclTbaAlYY0EroFsdzHnS7ezTirreblOZVLX8
WJL1YG0YZ4uwv1s0ST2AeUSrT5FZla0H3UH7eZEElFULSkTcBxyAmrR4+CF3ANFS
9Zrv8YFwD9cLt3P2gYvBY/FCkhfU4JpntrKvWMmQUKzLVskuE/1hvRFgZQJSeUU9
Pi/4PmKFxM3jcpDevbHeV3jXoBZ39VidRpDyPMPyMQM32a96mLHc5zGq26zlvRic
E2CqZUgKebwPq29KOC22aO+4Q9bXnlIFUjdyVWXKNhA31yqSqWU70fz3lVJN+GXl
uuVhat4Y14Oi3gCx/Gu4BkQn6wiRvmUioOQY876P1cgTfDP+C2SiZI5PjT/08lRW
Yzg/b+ADwOULAElQH1lENbBf2i/cPP5tCJowdfWcrJ86RQsyMptL+6ErnYCx41AX
I0FoJ6tkCPOP9WahE2XauDd2zF7nDS0Jw7Rzz6VUwymDGI7jDyvk7Cy+lSH2/XUR
hq3v+lZq3FSdQr/KxTawKvOpDqb2BOTVNIzqzJSBjVg+FmAfQcXAvzq7wRusufdp
ip655ZW5/hokO4HPDSpZXACQhWuUWJhacAnrDbHj0AuT22hiOY7m/mD3NGaYtI1L
V5+X2/2+yf4Q3i4jBOEF4NI/mx6GfxfHmmVb16NjEV2+NH0rNJ3oABPGTItJPmpG
`protect END_PROTECTED
