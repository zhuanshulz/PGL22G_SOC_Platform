`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CAzi63Bnzv3McQhiISvyqYbPSKYDliPQP+foM7HBZNwjY4bTZXygDZPddKO3XSsL
UxTAcXuxTpXeEwaLBemBxC8WwyShXyHC910zmnSiawmwL4UDR3Y/eBHLg2IbIlkD
QH+3BGl7LG8mygfJ7/tDkZRikzpgrb84zmjjD/kJjoAB8QAY/ANvERmSMPpTuM4R
n7PUDBKy9fzneNSj33XJ1NDDLRObbV4FYtm4psSA6G3XOZBOtvxHwOeP0PYsgs8n
0AZM/+FmjPIjeJqqtgrSS1EckrJvQqo2NK/5Rb4faaPRLXo/LrDNZIIVmh7Fd6Rp
J4PBDCprfWMbvK+ySEPU1fMUxXYu9FdYfLNi89L9kcdWQg0K2e2ExwAeYvV9KnZ9
NEshEt6JYqnOp9xMHAMHCWyJAJ4IX2VVjQHGIZP9IFhtU0CbZ/+2wRxRvZfUjr3+
1iu40N2ZfatBpnWaIiPSjoxmTmU8jWpClO/5VUzIiPousWLG/KWtvFkdZd66yqv6
vDdEvaqj7kRoUMhnXzzVH6stMNBgvAt9FGF+mmzxImW7BPT5xEuBAUJKTyUszvNU
6XwV8lo6MUWZtwyRXz4NU3XbB1L+1jk3cluV4VEqSBXVEJ0uMM1ufVm2sVLtKUrY
pTYTq8wrkVtuC7WDPiRrd0oziHYhuAo0ZQN+SFvJwEnsrdzHCphSJgIA+wFCbDJV
8UwiX3IZ/tlIQbQA/pdEBlNflsEUbRJFk5rthPW0RhA6CmO9WPbDOLjJhLY/v48C
29dz4t/ptVDImI+5++Owe/hI7thJ5Ck8ks6+GOcbZW0=
`protect END_PROTECTED
