`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ESYaD8MP8ZvcV9MP7tS3n3Lf789DCv0EPLJsODE0/hjf45PoW1PU1wKuXV1Gaq0L
sBFeu6QWszRHF9QgyQ2bP3vvEjPvzP2tkH6kYNAhbXV1+NPtS8qfIT7ZyXSDu5N8
eHWVVW86XawtlOi+WnkJAvrj8p/C0sj6GraA6Crg6DdM9eakfZnarXbPibyO7yV8
c+KHyyYoxVhOc4G1HXgNBm8jvT6qz1EcPsR05waV18mApVOXG2m6VwBMMjbjmlW2
cMNfcZUqaUy80NI0sZeo5nU458S33V20hBoVsDVD1kpuBNp/4lBfFtTa/ixuHTP0
+EB3PUxwGziOzkYBzQjXBoNvQ+YvOlk8qS4W8aJVohFr9GgCQ7rOumtWDGm1NbVm
s7jPQFmjgx3P8giH/Mtu3f3noJtVOPmOfpY+eSpkDHSts9XnbC7RnogcwpR7xHQ9
OBniZjCcGS9smoUPjAiCqWCd+FwnZtVTuq3Ycthm3bjx5wK8FntF/xuqZVIH709q
eGGARZUZrIKQfRLkLa5MZQ==
`protect END_PROTECTED
