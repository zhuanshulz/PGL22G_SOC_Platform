`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocVIIygO6tY7r/tKlcBniwdfraeHo6dO/1d+WSYtI01nsBwcMZoDUzobriSfAEKv
vVWF9snCSsR1t+p7l/sFCJXx6FtnQ8UY7IJWkNiSKD9QkwQDMslfqEqTKZP+LQRT
wr8UwJ73FxlwmtRbt1/DRhL076ZmDjXqh34gwf4HsYPX5kQ7UXg3/wbMjhbEKl1i
EOGrmawxjOmPqQecXeNI0dSD5EeqIdIHafViwXKcFooEnvKoyeXTrg/w+d8ZaDOk
8gnj1KjMik41uGdQFXmlXzmPO/h3c8EPdeRyVfjJoGLUxp8g24JXzv70Lq2QmlBp
YzFC0qsoFL80PFJ1FZ7lUpIoWYGh75mbIt0qe+WvTabP4drx0G7GZbc4dGb6OH7T
C3i7COobV3jT772gPBoqXLoRLr2JmrfWamKG1gRczl4vCLm4F5tjxgwgN2z4ZF7Q
ZoKP83RI5UcUuQUm4nwAwGL9XZA4/dYT4oWyPomSDtfJK2lA+BGXoOIHgTva3ICU
awTOWnrngE0MF5FcyHS6uJ0jq2ZKhSVHzWm+Euc4ZwpCj/fV9cPDakfS+NVx9mAb
HEQPvdeMtfThez5HbRQc8+kJ7ojFUX5MP9oE/OI4BGvqOjTiFHhL3GEkU04vQek8
sR8TXTE4MhSMCZtPFGIRFd7NY6ule5FC4aTGyg6mTgUNF12Nv3+mp0XyzIM7cWJR
NaQZtHFFiHR1DDc9/n/B29hOL0fIEQiK7vS4mOQSP6vnBM7+6JLP7niyzyaIcrn9
q/VdVnlmvzcn0MQIrwc7uStIdp9WPTW8LhWsTkuUKStMtAGebKRm9581U0XOZnss
g2EFeJKAG10IaIm2PMJpZo/H0b6Y37l2t+UX7KR5VvFahMHMTlU4vhKw5IX+A39S
QBuQT+a87RinSIGxnu190Imw3TWC5ywnn7QwXMgexaHyxcYfVx94cCvzMqJ/uA9c
2v7EZE+CdFOlsfCgexh97ikhISpiO468B0bkUNsarg35Ge2lxkhb6Qrg6BGelIWF
TLIvsBD+OUDw3lWVGReUIvgOaDwZ4U6Rcm0lzV36TjUc3XFtIjW0UfX0ONEd7qIM
vllWAc09kXJiRuguaxqFGr1o3ewNlYHY7rjeSfMfYIlsHBgZDMGw7Nu79rUKJY5X
9Z51GqvDqAonns5skAt9WB7EGgmaYY4JhjDVfCdq3futesRCb1z0/2bRlFyJfEm8
GSlBGtQfF7lWPEEGPzvoEiYIO0E1Pz+kbDDB3KG6PUrAlkWA1ZVTiboqATA6910Q
my3DczCrTdgphib0oVdgIsvnX6pSIVH2HoWrFLxNw1rIVhvdhv3PCS50QYA9tdGH
wmhVo5v0YZN+p3S3Ak+iWt75emGwcAgsKGFUeh2j12Ch3U4g5u+5JIfjoyW6CBKs
T70dywnxo5j1EuFWpQofnacspaNHqfmDTQC/seuQ4uXe562IKU1DpxAE+vIw72oT
G8Llnk/5eIvVG8sbU2EfdL0FZdrhEBC0VAqLXInmPbvCTzcVpQwS24wKwkSAFQ/6
25J/RYg1AnJ0L/AYczNjg/9yybB5pTdSdu53sO8NqEHEtWlPCVcwuHgdgf5Tigvd
z6JPS9OiMROjGlX/Ha45Nyffc7iMHwvyjb48vVhAqh3w/bedK9L65TlFDhKUicod
x7q2t5FquljgPsw9ppJx5iGhr0MM0oOgixiOcWYjYxC0lQCp43QySylvjzMpH+v/
1XkhMs7lAFDwZ/kz46/lkd8ZN/atGhF1gX8P6QorVzapak/EgSGzlSkLZzGp92pI
xslXYn6nUvL+CUEVX5yk995G6EwFcUVZy8dxnERNsL/wirYyfHNdzI0V80wkG5eS
mW2MZ/zluP0S6DYDx8XUz9GrwDFCVmDB+nVApPhnoHOzDQRUoldc6TkCu/twuMjF
INmqFBoDlc1rB4pSKymYbRgm9yq7NrBSZhM0LAMy+sbubwrgmUGTzVOgoetdebnD
iY01VEbh43rkIO60lkX99g0NUm2CBsgLu+rR/3ZqDzY2g85khh0MHXXvjQeDojxy
mG6oZ4JrgJgh0U2Eo4qGFHmGw32bV/pq3NJnQL1d4VIfm7vMwEhXzN8D9W2swkBw
MbxO6fqj1HO0JB85gXfiRSkXNaMwSiE4NbuVK1hgro4NGz3YwCjUckjsd9HZf3Br
B9IlFdgYJpcx2XY5t35nkVNQsrXFXyw1e47u4Pozae1k/NVojpd6lQXQD+hnzsqY
uB1kqJQJCvmBYfNIxEiIFtdnSixRq/sMDbDmcl5k9XtVAQmgMCxAD07pulMjuJv+
dKPAca9jVIKAkCrk2dE80RAx4RtwSG5Gppb0hsBcUinpBgdYGPIlLyIkWufD+D9u
yjAdXKtRPTeaFIHjUKflMOCEdSiizEE9BS4sNbrsw/CEbzNq5inW3pUr5C4dqG2I
FLInHru5amJxSEZoLGXeXBNucF+T8sPFllp8TMzkxmOwOhWwOAULPpUDDfTrPxLl
XU/iGYWbPqmefnvSPXFD1y7yonRGyVwgPUz3yZ+fh1damlZVO+Mv37Gb276efZfU
nmZTuVm/3ZIVZIXC/M3FGurIrVyiCx9SHQ1xFH3IJnFGjy4DyrE/bd1fXzh/Y3/Q
okHZCLLKg61IJoixys3HLV5MYxmiqI1c1ZOxPgez1SEkdEeVa7Q1j4wmPK0d2rFN
3XZ0h+IFwtQi7XnYuQ2/rxBzPcdo3uW3ip1/QDLDlrbdTMgTepsv4aWHs0143D1Y
nmmM4lAnkT52I9zCxPKLns507Zv/0fkk+qQnuBzn/1AKRJJeXJDD1zygBeG/Crs1
DoNuIKZ1kX8JUGyn9rWUdlcwLBrEzk7tNzQ9MAa2pu9HhL3+YA+oRCsuEv8iSxKH
S70UUJPqyqFf0XKBjsLoDazlJWW87GSjDuJjm7zRZxKYPyJrveL3Rng9jWYwJOpX
nHua3CuQrsy8O5GGNdLaCHSTnHB92QifHECJExdaI0H8WFI3SKtrb1WsHOVhT1T7
9Ksux7EhhJUUQfbF9Fb51T723vL2UHH+5iXJE5m/q06+Js240m0zZqrcZY0mHCDX
/4FkFjOt4qI9T/DMuOGcsa3zKbTsKI2fN+v+6smByXoYLIJRZgb0eFpN33ldj/jF
pBPkM199bysAHMmbrzYDmwJCLVIC01qfdTDvKXmP0mdUHRmsi/IPDfDJpKwGOPQb
DWbdj02/fyPxOSG8/2OWTur9VwVMCRqjKsGxesSeWwf0BD4gk8O5yr7LStg8BDyx
eQvfaIAWc42mzHuqoKR9JHovq6L4ZS6KcG9BbmZjnOfX7R9h05ryBWuk8n/1kmHN
xRuu3Q1cKmsyPSu0e+vWNvLDtLJLl9+mJkWFzXmlLVrgR932a0IAMXqLbU9hIHs2
89XVVPl9tE2k9MCY3qvjkq08IBI+SturQKf3IpN3Hlo9chStTDOELjAL4QIjtdNy
fAYIDMYlMcNMw3is/tAPEOGsq7y8omAslCZbECUV0786yTfyp7ZnHLfmkFME7myf
JWkPcce4DlMeYOnVhwfgRt68SsJlYbATesyTogx4zbxNyfHjS4yCQG07M7h+KArM
+LAlnzDQa1iwr0o2tN5rnv4O4XZN7OHt5s29UFoH1Q6CH2zgeYXCvdaQrLrTz1mn
/O/buV35B1ukMD+Q1ml9dG/5C00PshSO70HyMq/eYYobxpqJ7ds5Gc1QOzRDkoXD
P0fSt37i49r5Sxa4/9E8XgRqvMM/L7khxUcrONwYt6lpAciTtnj/An1QFaEiehzS
cBY3ZCsXxzNSH+fWwXi8xIgKQz4X7FN1vjm6bwttfuSUJOfOQ8kpBAZyn1DSvaPM
h7+vUfrZWvcg1pJKAz2eSrEynyKc2WstDdzW6DoOxkhwlMvyvVzLtYxKCyWosyBg
6hqhYpWIzRn406qHVVeuR8PFsB4ald2Fmoe4o4gyFMQrwaZiU8wg349J5NHSVj3f
SYDLktSFsa1LCP4Srh8WW9dK5ZNoq9h8vOpV99lqxzZ2scONRja8kjJzlnWFVpoG
N8WdmhFc0PLo3NhsiPbIFtGTQbcdHhI68nHhKhATpXyRplGwyZOvbkchEARgja1A
97vprIn7JZeOJ8Jfa5vNXuzBvHYSBNGLYsq2wYmmR9FiyNaEFIamQVdPEhkc0sbD
bY4fBQQhu98ogULnMNBjzHRxrrG5Rg1YdZ6HjnRpS+XaOCHbsWu7WgVnf8LSEbnL
h9DWufjy06JfCCQUisQlwZlIaqEoPKOCci9WpRCZk0ykp2pufQoG89rExlarKMBG
UXUOJ/S/Rc1zYntnjQfKv94bK3Pd0yJ1+rx8hWcLHTLKgoWm+p/ZB5gNG8Hwxacl
zYg6HyA8C7wbN1oZWfwYPya70O8+4W4rP6bcJBsY2uifT5ZaQbbWk38RsSAJILFe
dbeagu0G2FGdwKXcoNeRQl1r9t84/x2xvWsUv+NgHj9QqzabmB8/1wzmWPFSnA9I
JRyrKJkLeTTiWv9RE7owNl/GldPuQ2c9MqXpShhlINfErMCp1ptuA/0jg99YMYgF
1tduwns4g3UY5s+6+U0v9hK3Mc/LcMU+DexhVMrmkIujo3H1jjLCqq82WurfbZwu
H3QZGxWz8xjqVU4ZZi/XoNYqRTiUw5qFXjSAcqd4zpp7ld+yaL3SHJNca/vc8Scv
AxDkOvnC7kE93WTpdbf/S9dDzpHyXr+CxVTd503OFbNScS3QUJOs5NEa8s65S9ce
mRn5Ymc9tF7KYcGXUE2S9dZZbwgCdtyerwIPiZFnwCIRw33ndje9qk/5VAj//kBc
Q4qBI+ADTXhW3djsf5OXudL6KPKmP25NkBZY6e6XONkhg6l35xocmfOBEnWSti0R
1xZJ2WMGBWU8E6XCDr3itIYcBFOc6Kn7L4GHhzyiBNsurP8VNY6ZZ7qn2Agp1nmG
AsLc9CX4ILSbIPTbC/YDXE9MiOXinyMNiQ4S0/GrZXQkdtpx5bCo6UyW0NqKr7zD
Gs2TEswoSV1GwHl3cxqk7kAg5P9XytScmzP3qZI2jxvbEbjAqVush+jhmrVatlcG
KDxNElWrAGDfpGrpREPy15EUCRhBoe9y/kf1RVp8agu1DkddEvETGKuLNqZ6Y7Nh
HZjWK6jXSWrvQJbVfBoXB368mD63ptvPqjJ1zhtL5G/yssDcXRr2IrxwSyupL3od
hS6pUrm2S0h192b96wQ9qd42/YaHfN0HHtAICEllvXKUdSwqFJKSm/DHvATwoRiV
VYl4qdTaSn1S2UcsaVEwVq7QMq0Eo9W70GiJjOLrBB8b742+0U2pZ5AIaglkl7Vb
hXtuWvDID1myfO1NyJ/3LAsWXRGFskz700aw49ghpVkdJ/wCzc0qdlAJotQhpP1T
Ufk/0srpHpwujTOJIo1+niQjbhk7bI5LUDcGuhLG0fhpKHAb/qLxmSf126VyQQLh
NJUcLSzxe8GeDpNs3EMvmbMyftNl1NNzWSDN22/ENgKjDYiKFcPqtq72taNK6C0B
TCUm/cog6KEKwUMJ9o+pohL6Whic2EaF71SdtxzzIwllfKJDlDeWDAUbyEjrYi28
zb7Oq1+BaxwOUpGNrWk1POaULzxKsX9IYTY0oQMN2yPXU5Mk4HaVwBpMDxmN5GLt
FoRUduXX3XSLtB3yyAEfz9XVmf7YFnFYoRWVe/nHBbDlFse1QdawAQGN+CU09/na
hc/lkdSeGkl0hEtSkbo8yK6Dq9ldDoLQhVW+l130rb4nx5uyEjCD9wLlen+6QpBL
3f+QZxMgFAcIZGdYMhbzyHDjnjix7syIgk+4mgqKILyq4wCgI8A8DEw2t4WzsnJP
lz5CZaCwpCLdBuVhJ2xgNENIuH0w9BJvpntrqOvnev367ZDeOB5EFvclhD0QslnZ
3E9P8pPQXr/W5LS6HSobVtdy1rqY5n1qmgmHf7GTxQcr9VTLhQGIkpItA3poCAiB
dImx2cLxgHBbL78eFBcn/9dXcXvpLFq3DFKN+PVl1c8v2cUsBOEknApEfj/lJEjy
+NFxQOECyyuXiaRbj676N+Gtj0B5ki1b3Ok1KnPfk3r+ubQtACvD61234VX9Nv4O
ktQc+o3xdSz664U3e1gajCTE82HlIhn0MKEvB/qDiSi2GK0VQP/L3Pvx/Z7lXcEl
T6m7GghKi41Myv8mCEwBF4BJs1AMxF2gKg7B11pYgZC6XwhobuW3wIAB2laehxCd
Xsd8vGRYyWJMJmsKV4p4FlWk+15B6R9sP5rH1xjhXx1vL4A6XDAv8O6vnYdlfPNs
I8u0rYEY4qNIeca5fmSs1M12R/g0Nj/xxPNSrTKZ+113YIt874uNRGqVlwfiEnD4
gONU0AEaZo9KKFSVu0XKmlsUteeHwhkhpxdT+0Zdhc0vqDJ71rVz5FZw41ShCQ2F
`protect END_PROTECTED
