`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bj+NplTevt1WX9i8xUKTGcZK7cPoL9RwmabZ/O3h4+SVKygGBA9RBGeeXksDn9Vs
9kfg8bi+tZLFZ4o3na9UjnEsBA7ux/huSLTgY7SgNowgeU00KnBJlo3A+8bhaGRu
TM8BMi5VqCIIGfKN8KSUK+tm+2mXw0foh1mCAsSBAWU4FfVyynXSUOB/JWZxMH5F
CIAwhzR9l/AoraBY2SpAN/SObcK6gRaKxnu7ah6BVreAkzFUaV50LCuCnWw5Dk+x
PGNBlJDNgOvXWK4FLLteXE9Cxv/W4r7VNpJv+f98Ko2nkBupYnvyq+kukvWd0GKu
U9xXFDGk7q1RUQ2wOeegJH9/z5Tv5XdYp3yEwX/hhBf5Q5TFe5TPCsTRnF9cmxfI
abbmBrbDB9rkmz0F/DbL9LCQJzFNfDllsHP6o6YditGioZ4rGWqCjckWWlwOmJi7
k7LsQ9kUyuEcWqREq8L5Nm1Ym0bQhvFOUrMgqxW4u41WwGoW/cctA9Tq3tRhXI7P
KX/KTaW5t5rYLkvzLJ1IS+kNUb9+71M1gVk20iZI2Ty0mmOhuzNK2mQ+gPdnWiyz
arKBNgNfegvcs1bzEQAPiYkmk7VqaT0RNxtm4Fax7d1zunO/XPEduQA1FQERMRvo
YZXA/bouRKz9RRh9rlg+e1Tnyz4/zGqAPAy2dHdlTaSae5wlfwuVdym3oqlfXqNJ
WwkzK4bWpWTfArpr4H8SN9NUo0VITHXlwDvlP1v5gkos5WKi4+vZRYivkbV2YW7l
TDnA8uRe7V6gupmiCZ9Ddy8i4GPvF1KvcflAm+yNJyfUkUaUIFMnj9v84EsOixid
QlgjwaYrFw1Me70mNpwl51EHtzGvD//7dlwDyCKQ4Uy8IaIHD4307oSSUWMbL0a9
JSdcKVFFU4iyIvidT+brOx3UTT5zMM78Ob49WSz+qLOCnceFP3g6ZJOb8gDiTafL
1riMNll89hTZWz8eznk5JV688CRHfiG0+l3MN0l8Q6+HBjghS/TTAnLwqkZ2e1an
w2P6Ug8mA1tr4TK3Fj9zMmzqUIozNZHIxsl/WvsuChEmAwd+fHgfAqnINw52R6l+
nqdMBZUd4zrAH+W+v7NGIY5hCkcdQlEDhG1dkwtMb1glgRs53wi07oaF3G7T3z7w
3y8pfqXu9bJAjUGHQz1dw2PjnpzIIfZfTOYsT3ccVzXyETKv2S1vCOQCsN02ieDU
6iGPpVlGRKvJsEs9c6II5g4blqx3JdoQOzm/VL4aZR3PQTp1bQyEJN0H5vn7FZPh
gIY07PDnQGU04xUcyePkdFuqtEIGvyk+hc58MbZBJeE60PKzwiY4pkelfJ3/sNCw
pylYMsk8TTDNLHjDSHorlsDcUP3RFPA/OMVUl78bI5LSeaZB0LyjMihg9g9evd98
MnNRBU5+6P0Z9C2dblUBoIkwDsqQWC4c589rzwXk7pncyyWqgbrextAeDZPH7r2r
HowX4RHDLstgBusMCr+kmnhhwQ+S2COcFR+ebWvAqvl6a5W0NTkmuQC8b/agwMj6
VPNFrxNH/M/lQ+ZxX8IdTO650vJa+G+0PStOPyfTwnVAuqRJi0Iq9J2b9/yPr12I
6fPn9MIhE1t2lBTbEqsIV0qVIFaA5eZHXTRHy4cmgwxsqAHDw2NefY3RT80Phlg+
SKw7A35ac3hsUuy5q0/aN/naoF3y8uCUAvGI8buQADpKd849T4I9j3a6Y0eLVGkQ
myLIyFAnRHRFE90fyfsriRLwKVY2jniw1WUrly+WGj9pQUKCORtcW3GiDGuEtm8C
jQM0FrPI+PHJs51WXX5YpiSxmNxmZ9UCA7DJOnX6WG4cksQAXIFdsuF4OD2luFPP
TMcD0FRa7nleIxD0bQpDnkW3I6/7I/Gp0MvsG1fXsA8zp3Hybn9VPYj+PcX7oP0+
Vx37UJiKuZ0CrmbODus92oJ65JecdtdyNKzhrrOmwowYUASKiM0dR6ZBcbHU2RTu
kLL1M1MQtE9P2jDInrYAUUTE+z56zyOHgDSTZm1d9h09P1cjRlCDc2euICShyU6K
dksiUn5cOEKcmOefob0zkh8vo+v7Sx2g0C70qKqHZMmHVHkIr5wkT8TlfWXKAdis
vGWdwQ/iPrHtqEjSRKf7duZ+lhkgStCPPCXN0jBNuTRU9mxCvDGvYirO+LkFuxOa
9jdH3bHcAb4i/A3MIqMrnv/JkHYZYGgMvM1tWkqands4FaGBUbccWYGW4lRHvNOm
5PMiTYyb+ht7sopovGRWtOUrBWzVS8fi2d5i4W+kfwazCPBqwzCFyxaDdB2Tk8KG
yHBNuOK64DvXZ7SIR874cgqOlwLi6XGI2g6iLnrBa8LFyyKofT73Klhq0SYtlui/
8EQKETsED5u9A9FdmTLu1nKNzkA8fjAzHgWx7tnoHgvLssX0GlhpRGEc9LnzHGK9
Q483R7zLITD8guABXLiJHLkhsbK7F1pMOn+AJ7STXnnFSyCw5lS9iuesE039x8IW
grMzyokNmUDG1Hj6GIFwpx7gW9HsJfdAFCWLR2WLQ7UN78NVgXR0hP9UcFUJPLYr
3z2/HYZO2GyrhQF8NERH8ZqXGrNT25Ph1Gne9aX07JdBWRxsTPpwgTQwlMteOJgE
3c9Q8hUUEc/eJ2Y5OR1m1CPdJPTkgkPYq4gMGkpWexoN39aBLKGtF+P9ayV7p0v7
gIrU15E/08nE4ooO4n47Xo8ldc8CNtTN1/MsyeSybxI5ucyRtRWkj8SVWH4zuZbT
oa/peCaHrKtF/bLSbXppIj05qS0DeGm+Jk0YHrDftFTP33Euc6UQGgobw7/h9OOK
0SRViO+01Ffd0DkiQ9cDwtuYKaSNSHxaEvpffcW51pykaxUs+k7q6P2wYvdTLgdj
xIL6MvNw8ERpwlkOMGby9CX1viIPJ7QL0RRNIAN2HrunwkBz3jKisCk19RrHBWTc
4n78yho0hdm3ik9GqFOaTOml6NP1G9EasHejgI+FAjI=
`protect END_PROTECTED
