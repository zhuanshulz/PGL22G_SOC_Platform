`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YUvr99mfveJ0dNWiP0FTbISpA9/us3cWziIMSJ8WRjsrbV847Wm85f8EjBrVGMaS
kq8q6k5Wxu4eiyVTbVFK7E4ntQBYe48hI7tumZ5urcLV9saLXn4IGg48I7d+tpMr
kxwKkLsas1UnJDanuKj+BYWdumLEB40bsLcAXJ84EMeaUCg4LY9m/7SbvYsq08O+
ii9iNKMDwLVgEIiQPTkMfEeo+09Q3ikyiNC/ARM1jployv0MrkL/k1Cs5zHYDirF
xXo9+tM6PXiAw9DuTOraNwa+BLBeDIMWcpbRx0qFyJs7HlBnyiuk+K+6OR2ZoFPX
SZPnCLDRkOJZvhn0GPXXbShaIhIS2N4AVyjHBptZGaxDjNjN/bsPvoUjUC+mnRKk
Dujdf/5nca2fGYld6tziHvYrpLn60uTTokYHLoVB8k3iIjMtKHPIg9TWt9Gm9nIz
/IG9t4nuB81hxIFqiGN400wP8DO11CfrQTXTUw0QwH2CZTqvoolnFJawX8BUcUsG
7ukiVnRCXg9c8rVHEPVusZQ0eYfLEMDBXWilLG5O2wEIuc4cOoH3M2TT7eYWVxNS
BviVdOwvesgCsnFnU2M7new3fN3molSD9Py1rqVDAPA/NCPMgdwJRjvmb+W8zxWl
5MZVQE/OAuliJiO4igmibqZMOsOWQ5mH8oulHUSOAl7V8x/AHmSCLL7SmNeN1+Gq
LcikqFZR7+YWZPvwKCOEAAXq4CWwF4GqYwE5vOZ83Hbwe+A5V1e+UWPdaIBmRYPm
TdsSNarCifliVtxIY7Jll5xyrl1VLn3I/16u4XEF0QqT5WWbq35fP7LfqMSsm1n3
BUm+HfevSt3Kw50rSh9DoBSWy8kOFQsINzikJo5nY5uP9KEwPpISX6qeJr91IWdH
f6Eed4hUYCKi/DfYZQ5Z3gDM26SH2qzH2uXs4TvH86GLf3wqIHlOeXf8YIXh08YA
HhaUNsbqdO8+KQ+dXoAo+Vhr6TpVix0GbShFcDzspgJDlqveqIgfcJN1/0xzK3Sn
f4OYdK047lWMQr/tL2NRc54JSLW6OeP9DtidIawrhrIcHVoLHIFR4VzeVXZGHeBe
PdHu9LeghOGQbvq/aGJHIltq7/Cb67SPZwKiLGhs6MNTdIheUn8jYi4UFSy3xHGu
h8oOA5+is5s+3oY/BS/KkYazfrfiECGqEjRfQ2/K0Rejo1oie8rkyJ4FiWb4JQdw
SuWByB8qEOOZ1wCoqpGfw60pzCo8xU81nsLUEz1DBE0niQEkUuDlNkrtCxTTrT8K
i1Tt3y7EYJze5QgMMcWGNELfFbP6VJ5x5Von52zAck06ZOV2MATUM7NXqtQWmOn9
PkiraCVPxKkucl/cVnhVtSe7gSH9DO+JpI/jhMOBVFzW++2OSyDxbRI5aexiCxAc
WolL0q5gAZo+GMaYs8i4C1YwhoDuEP9AxqcTvkE4LwFM/F9quZYWAfUmr8ahCSKl
rTpD7JiVnIxXbZ5SAKymw33RJhlNvj4vFmk/KCxuzK51h3kAJUF5ruN42iZTlHQ0
GF52nGH4agP9rbB5dfR02gnoXcx8BAnWsMqwPDsktzSLdj2cxDYDaqfQbhfMvMjq
8kq6vVcOGf0DSPm1SSySGQG2kIgfzsAbZerlC2v/BtuFlXbaCXH1uYKjr1GvXMiu
GCknblT/Ro3rIBEmOj1MhVnV7aZ+hmebUNxxoDvgBAOWdAUw/3i49Bh+bBbH0znm
K0hLTMa+4Ffy1A9Qd9R+vv9ki5UlUZUxt9Ca0tNPBRH1sf6lMfu/6PK/e0u0FoZo
mlzS2VXrLFPBacY2o/oFeDbIq9ykZr9PCgV73UX2YxCwXyHDnM3tSfSsc7BNSmm1
tWoXuJ2lCdAB/eKs7aYSOBOI1dzYCla4T49FmuMhh0GXjZgx2v/BSH0YF+/Goi88
wfyr95/cUl9mA+dCUsGRTFHQGNgJlF4H7QY6FMKzMKBpe5bePs7awlsXB5ERx309
C7QvIKRNPu1ba4iD+QcoR8tjPlGeN9pVRI3ceXZhDgxsR4VM5yEz5v/BuNFiKMiI
8R1W5LvsyeEv8zInuni3EOsPBJkaPJpmLR28AEBgdMAY7o8t+SSlHV09UH4RpvrK
wLOZQV8RtbpFoxox6adQs0iFGLlOnhwBVR6FgiL3TOyuD8CLxL0Mc3V9rABGC5sz
F5/m7mSH++HxnOdrdcnPARBlH1tdJUuU1sLo2Yjyb4xgMB6kqyqHsuocJWtoZ98P
AyImUI9EoHcVoEOnOCoTn7YnCsILFjqIQbrlldyMaFNoNifCrTitERj/Iv1Wenw4
oo9bSbIPdPsa+JgSFqU9+lxprOGSuGpNCs7RUNg36ir/i4T3HvHE+NfTD9YCAFFf
HeX/iAHu3evj/PLjl9gzmkuJUlJ/wE8Vfpzy8PoQGXL6qC/0qPIGfE0Ro0M/ccKO
KTOvLhh0I2g6IUEfCTqDYbKTxz3XLRxTT6WzV3z/s6J0pXneijyJYYZk3iZ3e0Zl
DnPKoXu5fXaKjdCfkl9BURI5Sr44xsojWxcVUMvEyucSJddxMKdSkhn3SfQrVI+8
IK2MySSYJ3mhpLeSQdT12qAwhUPVLXUtzOlt8X2j/U38StX18R9Q41MG9FtmpxtP
mFsxrTIz2vKHxGjFgqnL7+W5xtvJSL/d0JoRxjeNNsrViWSGSSdlThbavViCbtM4
ptAhWIuga3nYeWcQtL/l1/vI3vblNDp2UqG9rzoHyN4w0yqprpdGcFIyJNmdjnDF
3UrysZijbOilYBURIVo993Znufn0Tdm1FzoUD/paU6NJ/XQesTf6iYvoQ9uWOc3U
zu1oIMRHX3c8/aopQrgNlKZzMtSXQzaFuNO5jX9F4NPYsRonaF7CYlrpp1GmgYpu
UOmI7JLMyQoO8WUrX6h1kG12VlZRM7vAEWPfz4oaz6aOlT8S1ZKM0zAnv6CHNUdQ
E9q528laBL1WA3/MkdE7B6F7SD+0uoh5NyrY3IyQDfcGsFFXvXclAVkF7AgOubCo
/RX/mo/YmkC9LI/wELuI8hxRANMamTffaoxExn4TOQP3iUz7FmylYo5VAKte0iqL
vgiMlxAz6jObMntUBR8+5tD6h/yMwhQhzHhfO6cTwbwMGm7V1GBJm61SAvIZRW2N
8BavbwHy+v8Yppo5axHpSknukv5oTeftFnJxPvSBA7L01+Wk4IBqMtb55Wp3Ru+4
ANFKVxewmC8sW3zf1uFXeNNC4diINAEZQPg7bZS+s0LQxnmlIBnkDpV8JaXa3elZ
DG78uLk3P+gradeXJ2g73KLzBl/ioKa7w9QzqLmSKovzrtp7n5cmEHq4Z63HlGcl
PPPLUKsIkx1GniMKE8388aBFoHz5icwe9OM/rTbhDeVTTKzeYdvvRixKEqA4f6YB
cqiohYrltSVWrzsU67IPaJY5FSXnqa1aTCujTzJxVdwxn0lvs1JxyFSmZELcIp6i
A3o1h8IhwdKBxsH5Qe2Qqw50qaE6kwsQZRry1+AzLxj+KEP6IeB5+fWKHIb6er0+
8MYSpJkpBRS+ApHeSJEak0lwJ6lpoEhUu1Mwg5QgBHOlf2LJh8W64viq0OWZb71s
fX2VW6tjYEhlYXPViYbq60qNl4ZLSFMopJHTnwAD06Xq1S9p2HqdCxt/84nNJJJo
uha0nERbmxQCeNw+DEHe3oY5EMoKoN7jWGNuqmgAy/KsWA/AxOuR+MaGpve8iwdt
3PECGvlF/Sve5Ds4P6JpF7PsAquxW28sx3+35GHDRD0EK/aHElNwavp2N+FNiN3y
8gYAW1jTOJUhKKFICA8BcSF7wOhDP+T63u0xS+u6uZdWs/IeLKaSUiR3Tuogrya5
O1TjJrk9AXHwl2LyFIeXwul53S/zpm9NAwvR3nURMp2YalQorEw10zeAroGouB55
FYxz0Bso4OdlVKvZqDjfdzS6RG6Ne+1zsiKwa0AKZcBP0fDSfFq2e/3hCzd1mh8s
VmOJZ7nQz/9+32iLoCKt9WR48VBglQgY0a/UQRG6JvnIpf020KSvusVoGHmwQv8M
q72L1CVjom6P/4RK+uecIX4nAtcofs4Gct/rsQLp1TAPtDyHl+zrNnVeTsldSDvc
Ouu8RsKbzBiZwi7ug8zlWxeVBbY388AS6bbRov0XtTK5pJjG7yxoi5ERG9nA2S6L
bLAEyIgvbL84ipIUGcbXzIHmfmMggn2FE7b9lo5KYSp716O4CMZO3H0MMnf1drGy
vzGi5j7riHullmADN8yX09cNKj9SL8FrCrZ6L4d/hiWz2GRAfXW2eBK5hKh4Bjai
O3KfHbHSkQn5qTYFoFaPo65bNOugIHwsZcpK4FTTBZXrVKwr5vmSnjmrx3N7sQDw
XKM6snU8PmKd3MHEi/TimuxODR/Y9UsjmIZN3pnvhUCKrlgE6n0C2Vtsj6FDd97c
`protect END_PROTECTED
