`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0WbEZmDvQc+TpUfMZvL111G/KlCO0QuqxwypKATHORQxq4PWY97sYb0rNVmipVU5
xdKb6mH6JjuQw6cSWERWWeC+Qlg32hJCd60UK7foGG+NiNSVle5/5oo2uZkyGr97
jFicPOnXrHD7FdDnRWSEzOw418wWuqUSr9yUaZr6CrpNHi/Tc7l+814xizUNRS1h
TxdWgBwLTDNvaVfGDMVMwLEXf4y5lCVAHBjktEx2Qal7OfBfxq3orj3b12IguwRT
avNzXym/ihzWcf1pP7Ju3BRZoHIV9n7UCnaGclRz6nwkDVgdGM6gdjyhp5wZK8ic
dugxgL7ZA9E2KFljL6mIosTCtXCsXr41h5+kMoK1wIZDOGzffIRjeQe/ESFoRqI9
I5SvktMyL3WYIgbHj1C1OoFFoSjBUrvODMFvJ/UO0RxSx67U9gjKa7oYJdmPQnyJ
Kpi+/AKddmT/HZFf2FuUjr/OKvD0DhAx9jqzY0svIFlagsHa8v98tU2X5qGpT+m+
Or9PKonckVIgSykrBpv2+GTVQvRa2ag2FLncJUE+JRvLcXfRQho82gl18Xm4Hwd0
O+OHEKRiZM1Wg5koACkwyPSTasZ1X35qL5H0f4ymHdNFtNME5OHutvVLebmJg2OA
N5wB/cg8D2gsbwmUJ8BptI6r/viCY4++SmBapgsSrVUyf+IoIh4Qkde+sXahu79Z
vmCSoEMHMLQ9sg65mmZ9AW2BK/WjdpYQyFJX0c+66aZva2bHcDn4z/PsskY6lGfe
/0ZfePlexoTSFVQgxhi8uhp5JnfeqxDqmhA8eHlMbDRGfv/FYLuihCnRyd0zkXKA
ZJc7mv+QNMxafP+rLXbwLW9oc4fbW2DFE973MOBzXmNnqNSIstCXoMHe1m1mrPBd
yXzIb+3OVICxZkBmJrmYgr9L+HjDKAyyHLbq0/fcdwofvJH1ZQkYyauHjFGLrZ2x
tgzlS/G4JhWqjLBT/TGHrQJVb9t5wEdc4qNFvPSrn8apag3dqoswDz1WEy9zBS1X
xwz1jjmN81T8H2tMllxwsOIzo/KRQKwjtlocVkaggGQVxB4+IMmXcO70GWgG1cvj
c705YGlgcsMwdTGNgEn2ItlYh9FIJ0FxgEWSea3v8kSySo+uzFeh68FJZPpTJ8MO
AaaXXBHe3ZlswWt6mpcIipE4KEeSqfLjakRklFUDYaJ4jjLSX4AbmSIbmCp5c/C7
rCgsmnbj0LWDTOU5jotpyd4PMFsVvnUXR79lb4vQoY4DXm5U/eDHhk05c8te3ZDA
bYndfZJkZLduQ7akE60l3VamehY8VLFctVe2E6PzADuuLDapjnM3HpAzuw/W/ZvO
7N04h+nK2u57Eb+zkBAH5oOPArsJICfQ5Y690p3YNvaD46tjxgsynkAHjIW90m6i
fH3poK76UQ0eiQ7XY1tkw4MY2De5S2tDoSKleRh3/cqFqTC9seMjngM00z9u/k+a
8kes9szdUyfwdJQLeHeyBkRjo57AwprHmegHdlq3l5ZZYb6+Cy5wOicGYXS2YytV
hW5J7XrkpxyWgOiEx/uNdQhjLFQyBhFVPJZeJsNQUTxjh5gDkke9bFZu5WeU0HSb
QkRg4r0Ov0y3tGb4kF93rzyfgRkTIiDeA1vwlI224gcsEg+dG85HLkIboBegxAL1
8p9s8f5saHFbE8RpnUO71nc1+l+GAbqivbNVid3mrBfjOaIv7rkzqllHIX/dMGYE
7A2vad9dsTqdfsfMSkVwa8MsXamRgRprWQskXci/Uv0jcK4A+NIl69tRVBKrcLE6
/pEZ+sBdw1bP2lys8mQefH+9n8s1JP4yiggR88JPrHltkQ4wCNu+ujeIkYln/W0E
lfGUaVV5f92yHNmUi6lGKQaIANAaHc8dznkq/W/2fmvMY6WNra/+wk8/QmvXDBPZ
kQQ/xfGlFjbhtchZgT3tUgCEctriVdpJZbAsP/WhTo4v/ZmSH7CXe/CiYRrHBu9c
Br7+73HHXfGJ6AyF+cWNOroytLnLbfY2OnB34dxc5uFzweipqnzA86kLcauHY1GQ
meBGTz5gmdKpBIP+SF4f3ebbC95ST+ocpSE3EEd7Arm+W8+u+G7fjPgeovpeVAZm
C/yYc/wQ9SLT47AumBdVfCXlHh4/aozvex5BGfR6eYXqoD7kJfsPUOXtpXUaw0Ph
V18bUo8N8HWsuETbVgtRFfAFdJrHL/0i8YMC9Doqil0QC5zYDN+rxIus1VSB2S+i
u60wJqAVW/fuSoKjHGxwwgwnKaWUvriHjGVy8G2kUxLqVt0sRFzkFCC4ACra0qTb
biT+SH2cKzvWNQNWzwi7hvtuS52nOFsaH2/fPv+iS/OVBPs0so/x+JrtG7YalR96
/o1kaeqxKkTi0ll4VoryHJWMe5GGV8YHDXg+ebNe3bxbqqpIgSt5xL15p1xlpj/V
l1IrWlxkgRJUzDWgYNRU3AF4ej8PBDfYB0QGByXvOwaJNtQ3NRGZz6z6d9HYzhC7
6UN7BaQPwCpQbQ2Jh+RsOr43TTqkt/Vb7QR6BnTaNml/dvkVEwP5En06o00u9ILk
vjf0zZwu8goCUigpm6Qd4GUHN1BEvNAAiKL8igNYlh3e0crrTY0WekL2orhXNQSC
EHvQkYU+Ls7zp1Xv7ZQcMLisuE9QSOaGs3XW8DMQD5aw5zrk4ccTM1/MEHUbjYPH
Y8SypSp2xfMkvHX73uyeXbRAGpzbiBaawSNU0GTEMcp+f6zSPb4vbeG3Y397bFKv
O4m1zQpcGZCw/6hDgryrqUVRnk7Gh59Po5WfLcLMDIx7Txw7rUc4Ou3VpZ/8ND0i
MWv4u4FpUrF20n6GOTPod4MNVNPLOqVAfV3Q3ynLMS/QJOxR6YwEeoPqah4XzApq
9aQzpNVVTzWuVu/Wj7IgmKs8JldWk2+pADZgRzLtp7XKLh2HssYAkf0zyQ6YjXPS
bPEO/f2N9KrAEmGhTGcJk5Fc2B5c3SeROqwIRrFJRop/5jzxe9Mq+RqLpmPsdzCU
h1wHCQ46DdsaFCpzdlIy8H9RUdua7XoONNmAdzp33igfxB2wvnI50RfPa9GV5Zl8
24fvaoq0cyouDfkbJXRGsQ==
`protect END_PROTECTED
