`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
crSM0BDu+rpgQCP2Y9aw40mzMsUrM6Q3HXOgruEN9/EaiFyx/RR+LK1AjdBrYdwJ
JCq2XdJxZxEariA4XFnsnx3NcXTk8LFoP3tT2EmrDYsFdkAlX/R38fvtnJAmWGfT
+Jrrtk63Zr8Bokt/G1+tZR0kZA9DzIu5FuuYegF93F26vhp4EyNC6tLy88t3O27H
BDIi0IIFlR5hcvEoDBFq0uYZftF0rJCQokGSsoP1AfDdKV/vmRwYAiBoDbxgJzyk
MbVB3N+/5mcVW4W8xi796VH7UwC+J8B8+qt0AT6+3Njuv78rWVBVNG2rnkcPePC9
cPczwlzSHAbWBAV1Mj3iRj3Woycv7ju+6/pVQMNCRoAXNETbgNBap4kRr8QWbSt6
yG75/bQkP9VdhrrZ9vmWTA/+hNIrlAa2N5wDMwy4WeSfo0Mb2PS4+VOOt/y0Q3BS
FEzqOpyiw1TjG1mUiXtmF5hdAmZ2RnWSwwGqAIQpVOhro9VP4bFHSSXHm3n1LbXu
U5iiUR+jgkZuVUJr8CVNlzrW2V3ZpFC/S0omltRAJRdsvjENucjejdbKXG2H9nDO
6Zr/uuGnDsJVD9M/AJ790vJ2UG/BMaNT24y9j3te/sTnQBWnL+7vgWxChZJl17vW
5ZomzL652tLxtG//loTj2/A6MhUI9aT/6CS/NSVlbmY=
`protect END_PROTECTED
