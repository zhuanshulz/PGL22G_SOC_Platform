`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ToFSQJcVKlMMzNA6VluDDKSgchV+nZTMZm2H/f8z68xQnty0ZykSIPi+lvlEEehO
ew5a37AkngfK3wcpxy+UzcdEqAwHS9Ah/oJpfhDtJo3KOpr5kL/qhRUaMlLSaO4e
/I6VVIs8o6K6Os+KPI8iCcDh0cNaL64Tba9F5rDKDVdkm8+Rkh9Y6ioHDIrwHO1M
sw0J6pO6NNiL8314ZBtUGI/QCK5datsW5pjYqabusMzs2Lcj7E7dBhSVHSD64fPN
KHmjP5sF2/EmhBqsm4XkruJ7fQ8CMduyuwGssZX/n9o7U0qDfmPFooZRczHI2Hxs
4077XK9VuHbYvEkWz+DpGU3K6ppJquEk4xKM3+/CveSdXBFBN+NlifUEzzxgUhvh
ds44WwxfZ2BNeuatHZ9mg740VpaKxg5a2OtpieguN+LpnCLNTU8zWLNl4bAmedfW
FeqlBThI4lhlH0Zh6wLWteLBU4ksPOMzZvp31G6l2jjWw5FrgfgDXw/WduHug+Ky
p6aJx+Im1utKETwUhFKepCDKtKV8dnxO51uE+mDlVWM=
`protect END_PROTECTED
