`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EmaPrpPo1HbKTdgkiyO+Kx6iMYtVAcoGAYyeOFdZ5kYWyw7psST/AIMN4Jr+vgiY
zwY0cyq4PFlwAYMLDmi/WuB9DxmAw/vR2uwPzfNCJlmNuHawf8cg6DdLX6VkBwEQ
uDtqz27xAwiozrD2uP1rSQx3G6Q+DPLGRjrvbFxmMtbQEy0LbyqFRJ8qOMhtNYGN
a0TbB3qUIOA4GztYV9oa+9nE06J2ubzsaAuGTn2ocshbnxz7xU1ToK8BMvPemEUp
MdAUsApiw7OTrFlGAvr/qWVAt9XOHF8tVZnYlC74u84n24yErjyKnuLUtEzd0rtw
8KeDl2zx6v2CWnEIvGiGmZSuCLYYi0tyxxkuu2q/RWEKfwYeYjq5lFVTiwFvkxxl
R9SDuNtATr0xfGENXc4p4deHt0dybmEFNIFcJRlZLIvaxPVec9WBW+xkgpXhUttM
SBZFhX7/O+EqpY1XvUNkinGgUQXjbUmc3YUMOMXwinAru0hGEe6kE6XYFpw60ME+
u4bey05bIVIAigspPOfs86QT2U0a1Ow+5iF4Vem0fjpui3ZBwDcSNZX6hGk+YVaF
5sUYtp4HJPmOjhb5fKwYuJCqIBOo4wnhvgrtYDb4kLWZLph9DY7XZi+R4nc1Ijos
jkmvUYloK22xZCD0ZSN1Bn0hYS6AypKw8D6pmx6C8WEofiasPTp/EnxGdfKnaXnr
eAz5WuzYp7dSxlSYTD2DlX5GXyDx6yrlrzulVjtiX5yrY1FV/+q9fCL2naVSwhB0
mf1UnldVUtJNipdhE7ydG9h2iy1uubcgDo0x3beWfau0U3PsZqdg4FLLdhZTyGEQ
CCd4l4KwpvhnX3KlN9zZF9uwzZ9NGtpzxQG9cJpEgUOQ6GY4h3l6KtJB/9i5XwhZ
e0E7DEbqKMI8CN0ffGfhT/nWyw1W97LZRQV0AMOHIKX42ZiOW6EOsM9RADfL+Gt6
p4R1+YGYWJY0uNtoUiz9hdPZ1jPE0z39a8dkwQt2f5HeLJUppokJpMuP5j4FWKvy
Jf7Dv5Wile4a7haovTjAkauy8WRF8kWXQtOvg8pecNjrT/liRWeGCF75kDcj4XfA
kDW5wqX3hPd6eppdeN3iyfwQaKt3L0PbIAD0e0Xfu8XffwzD9rdPZ71l28RMSLkX
QLpMnBqLUK2BOE/6f0jq6i8jH+wyjNw5uuQwuRkJATIk3PUHGS3AXEByZGjxKo7m
K0veRDNOWxH+dgsMuSzcZipu8lLxNDp1dy1Knh6vHalW3LFjDrLJt/r1B73MkQt6
KPTT3GMtJXDvON8+YBHtuaW1yPb7Yuk2iUXa8UQ3nHqREo2o+0AsghWMpk3G+OfV
J6misiFi3kzhA3alUGn2Yv/g7jralJaKemxM1Cn1QyUxFnNR0a6MbDvyxTVJeTmy
1QCoZsxbmuaQwP775krwgZ2WJe0LsjJmmctGll1Oe8BiOibxTNFb7iO28jfNXage
Ro1I6P6cRVcDPVDXTMebK5wEyDhHV+2sKm/LN8e6jl+5TezAZJHHtwGnjm6HGuHi
pixMyftLyW2xSjKifzXLp8bOTUeHEmXlQZJxM6DybofPRkgB32TSdOtwae0dZMiC
luo+aI5gXaN2fSzklJLmzwGatm3NIvyX/F1EXhUz9zRplNG2ECv8QdBv5cmKW04G
L2MF3FwuJdHFD4E3p67abTbgZVIrrU+nJtaOUrlTaXGtHtgSg3AOvb3bwywCDPSv
wQ7Guxl/YM+m57YxIVxkVpC1m4BPR24QOTbMmhg+a0tFBP6TTgIdp5s5HI35fhra
EoEVZob6I2cF5+9NIjg1wFxvNla2Xw2gCIZXcKF/p4xSQVCzEhupsjSGVm0y/DpV
r8sb8Amek8WiXO8Mi+HdQHGMp9cYQdjjKInVHcfMPCMA70OBtGttLy4eAtpdCPNh
0fy6XdLIf2CBPM5ZEgyvsbcP78CfBZN09KbuDdH+wV+drbuWswBaIDGKnPM9DhAE
tN1rpxSTsuO6ySOuWhz0j1Eg6Fs0niHl9FGQhJkpLTP8P5j1AxIvpLXz5SV6fSWR
`protect END_PROTECTED
