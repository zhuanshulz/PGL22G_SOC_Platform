`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVGb9YBzHZXBBTydNQeMhqrc9wT7A/QUyswCsVV/if/Tq73YsET416i0Wl5pktGW
syp10dnYXNCwZLrWJUgbpj5/DdbGWh3g3UJW3rtZsocwpudV2VY6GlgUaYWfMdNv
ecF74NR1mDt4vtWlZtL9EZV9XY0aWP7YgvxfTlYpbqslUELzJjflV22ngKD2lYiC
w5kEWNFIYeMksVYJCkzF6TOo8LrKs/HRCSvEyS+hsZvdjUg2/zudEx8omPE4NTeT
ESBMbZ+Z3m5wncz/29ZN+IaoIoTtPy+2y/ZcQpmoKTcny5bygGeqKlaFV+kBf8Vo
rO/4qEqIpk28eI5MFF+HQiYJ+0uK031xYItvSq5fnpcwbQ55WCVeVe0+ONA8inCH
bdWEwdeXxUcbgpSNFzGCdW3sG1nkV5hR56yprFxaj70ZJp+pucB3+Hiy3hJrFgJ9
cuj3RbtHWfu3d++mjUMBWf5sPCMzsW++wqjhVYXSM9naoi4Aur+vOYwfm52z+wv5
HwqniZXEui4wj64GbSdUrEYsKj21n39IhbrlRyaassK7pZVSMx/6tEAszNnW/oaF
J2YaJchWViKU728gsipuzujUuYKSTmEXR396zsdex2ydopPJ9TKlsvbTFujtdmbL
O+DtvhI27KeYk7igQYKFBUK6SL6UujwvFbvg1eCyqTOhadVclcAJdZddRgla82Zh
uYbt2zjA+3LGbE9wxbKRucRyPXEnSkyQdDqveUdhkskYix2+075OG5mp0/muMDe3
nJN4Ap/tGQmYEcRfCk94ujwsfBQWQAQ4t2Ps/HhAweCm3OLj/Kt3C4kXVKlELBy1
QvaNcVK/DplBQ47cbGgRkcMW5y8WZNznXUqUqxMj9XG//hIRu4e1XhiZWD6D+N3k
8w9fns0MgeT0Ow1DCCYHeO/uuUrgcs8Wrtsg7R/SgsaBVSuIm3n57MQW1NAFIhYz
RyRiLt/2/QhKajn2BbaeK6GWydT7nUWXgROFIy3YfgQcxsukPMBFKnsOijL3A34J
+nBoQ0kHX9q5MB7wEgu8vW/qsKUFEj3sIarLLwjaR4GOWPTJx91PyHjdFo7ZV4js
RPkGOtGwSB6h75ijIXhz2l1SbTJztnLyibTEUcv0VElLVpPVk0X6iZk2Pbo5qHr5
ZOfQjL/LyvAKLHHanMmSRB3lMHlO6dXLVEWt540KKUjsF3N1MhNDseMQgcowv0Sl
skICCUB4y3bn9KbT0bC/icp3DVEdgIN1b/sRZuYeIfNA9rUIDobDtQznCH65F7WB
FjE1EhXhbaZJK9rPia84RqTt/9B729PAczzJiKxpBu2KkYuvCs0aZbWJDmoETq0m
qIrnggn2KzT9rj0RZu/d4lnND8Ldo7AQ4j01TCtOODtc7S5XjqgKSL7dY1sCfnDg
gnd1hinOhKvdH01bbYwxNjHB7M2abgsgAfJvyi3gBevFf/M7NdY0/ORr50BIblsJ
oLURkyFzlc1t8Wf04Or5msu5q2t8GOBGwbTjgIZVZVCtOCaaz233kuLIc3NpHQdS
+5nAIVTmbJs/PuMItmEcVTeZRdFUm+BiD6Boc9M+sRu2OQ/DCX9Rz++cg9kHntoP
imBIkk0WA5qepJvfso6IrJrLWes9R0c3MCHyAw4a5PZqNJorb2ZDv3fA6F5tP91z
IcCigVGGgoyVRALuBcnQN7mu86GDpVH8IBRIo7UPLoOaF/4ncnarHa81xao8kRCT
xP6NOPbZLRwKc4/wJctbbc8WT28xM3qaQ74uBknaslteT/s/GT8xY9kqaucZYhCt
2Ne3J5xa6QGfUINS1wmO/dPqa79owpLGoM0NKb11TdRHY44R7ZV6wv9rt2A6kdHC
oxkW2XZOY5r1mjBZ/jxADBNrB6CyWM/KNS27oKGDWdQIibdUAD5r3Xt5ZV7zkJRe
daa9ugiS0hRpgwQTUtv25OMR32my7BBGSuY9AeektSVh9sgtbalH5fEVk60F5XBx
ASTQyWbbu/D38HqxYcYuPktLlLW9iznPZOKczjcWGy5OQurh5E+vvjqfSp07JxAO
vj6CKPGEZwN1CgBosBDwr/MgVeUNKIXDVNEvHIrq0Dhv2D2SbNaczI1bUdJir/WK
HAjqzq/gXdr9IyJcQ9lqdW6wLPOoYBK4bwbny4wtWV1V35nHuVsW4wxgOs/X8Mx7
8Q+9Q2mOmmOc3ZZSpVYw0siTpUB6wJrmuc+zDJjTxsevzG1jKCqnnVJbKEM3zfp4
Ju/dboJekkWmYD4YmcxQoHEiD0Te8SzdGnCp+lXxPe0Gb6BMn9lRAcTMGhK/ME26
uk878T/PUllBEGlg+qJed9BvvReMI7bzz4YS42VPwyXhEo/+uVvyV72YeLuNhXau
1SQN56gulleBY9SrSAObT7IUv3RjiogeyupujaCPv33NSFD+fIDSgo5GdG8iA1dJ
/DMr0qgoKEpwY2bbkGNy//+u+0w7gm5IlpnaVZ84eLSa284sdy9FNltKB9mf+BZg
4YR3Q/PY+HT+8Ec5dGK0ZDiq8GzoWeF7hi47JywkZ3nlfDbpNyym9ZSychqTByF8
77rZ69rhMGtHqgR+xMT2Y6doWUbUDcg5d1QQ0Prbc1082e1nL2mkQ6oubxXQK1PB
L+SyyZl5Msm5Evr/Z0X1FsQtxgx2ECiOWHcEKHiOZSG7auy7Sjn3rhvdQWvfVMiu
DMKsm9aRYzmF5wSrSvG8+ZNa434MoZofx0SmErGbrib+JpmNyG8jsSSWY9nnOj8a
F4tmWtIFPvp7p7xI/wlX7Xu7OfVXt5VQnUbzmGL/09sFpbA4RuB5K4MSnupNxfNy
FsGo9u7jjdiDf1gAN7BEFpqdUwwC47eftEOeTBrC6j+czMxi7VCn07PsqpmUGfpl
e1S+/jHx6KMxDdZ4KJeK1uIVAMITRr/4C0EyYYqamvjrrk2LWUqsL/Nk8CNNPmuU
XSxOSlVAxe53+OprKfBwfq1ti1epfJc40wcLGowF37bSEoApCvfVmcPQzP4NsKUN
jBqBfRf+TOMKEoObg+8AwfvGz/FO4novlOt0MFawyEUJLaf4P148DX3Ui+BV8sUp
J1Q48LCWXXmHRQRskcNzt7SALVEI748F7Jq8dawbr4RJpGTOn2h90CytnkjxmBN+
S83cKvl/aCcUyiVZvyaySxV6UlYtiVp8vI9frfVeXzIKn83cxwDe5aVFLlZaFkgI
DZ9cUO78Fh5vglqMKn6PiMotu+8ymG1WcSqn4Awb3EXl9Hys9ckoATLniHdnFQot
xk/thof3vswfBvK+thtw0TbCHoll51Pl2Bh5t7X2WJ7epJVfHZwFWHMuE28xQ2t7
znG3cnXvIXVYPbM1ez3YGTwW9SoX0RpkQNPdMlue2rH4DRUVuWcEBaeTWPkYXF2M
IGDKZwcT3djSYPspDU0tW8s5fx5z4Jf1aX6oWKxJub8QCXdvZdtH+c8876Kna2Ld
O6P8NeJ3Nvs4q2ityky4/UNMJgAYU1JOqdDKCJPv3MWOtHayWlm2qJR0AiHpB/Em
ElDrUMk9e48GHlOoN8zbf7hMDXPMeogwRmkYAaER0FPMlChWCdCBXSUMdj/JLXPX
X/f5I0gqQXdKowF+yM7wDcF3W2N20cW046oQIDympdAL/JfK7S6yu/xiWtw4VbUp
iR9cQ1EGVlqwFxPaGclv8UQVPhNiTwYXQdJ8me9ef7AxtXJAqs06BqtBb/flUZPx
3aw2CnUbCILcjLZpLEGdbHFVO9LkWC2sXP/dHYvwM8k8zlxrU7NHNJL7L54YXLXw
DsLgJhTcL+rmJNV2Ck6KAoI37EpM+t6Fw8z1EC+KZ4LyAKfHqB+M7WnCufz4QRfT
CRdtZKic2eV+oxYshKL7hWB3uOVNMjI+I/DppIQ5zA0G8a3qZYhzQb5E7zx5uXyp
eeWRmX7Di8MFCAuMofcsBSv/4pcfeFkkzM+8v+df0jpVW5ZASTNrDKak3oxZB2CW
6MT5cOVD70SXOP/c6tlV3fGnHXd5hxuFh3Voc1/2rhurTOumNkXGIhKmDOchQtL6
hUZBKyivocKqQst9A7h12pzx5V91oWDWnjB/XE3dc9smGExPVUFDm56LopV8hDcR
UrhhRutZvciUabmgCzBsUoRRciS2PfDh+G+g/nnBcIlaaWdSFLaLqJKBm0r8oblR
OguZ/Vlx1O64b1JjUTrDcsJTks7m/DXl6fuC6tWKiJCv/rn6SQkFc7al6lxABrJb
4eYLZLTIgWhaoVMXVFO/TKxU1UOx68sEuF4XwSkqZ5PiETx5Db10QrYYPF8Qvw4X
4KxG+DTf369hIGng235dXaguU+8zK0AAE+v5fpbwQOeIYqui7fAZVRky0UnW6nuE
V/3MqJ8PjbfiT4QFw6Yglw==
`protect END_PROTECTED
