`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9G02Gek0x3BB5kjocunoH0ObR2otv3hznQFqVJklTH1HDeIr16taGlMFjkf17lJ
gM/1mNwaMH2iPQrp3MiBAtyaQWazaaM5kbr/cpoNArMQNUEIWJc2WEtDzTcieKpQ
YRbmVE6ZfjlvZT2dHOb4fUsQb6GpkAGTQkqpqOgCvhd3r777Aw7jRmmBNoKOYXR8
KIYmofaIs2kC/iwBrXEkLFqVaLgzLdrKMfJ0Won5U40zEIPLALaNW128GVlDY8kk
dj3HMs7ThlEJvsObosrKg1MbWjmqw9laSr4rlczHKv9RFvfMUVJpMw4VyuNyFf+E
7DYOQjwu3vh70M4ngEmYasm+Z8e3U4RK8jo30AWaa12Z03Ib8Xe1GtxK2SjgQ60q
9orGAU2jtYVBhAbGDj3hudwZSEPar914+zmaDUDg7OqmZH/XLsLgS+N3a3v2YkBs
CCTYRWVWcjW7qOXd30oswcuekcczE42I6wnzeuW91IW8tYzlL+motH/A/A7RTA7a
`protect END_PROTECTED
