`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
00KNRu08Mrt5UrK1rf/umcHNKyydYKkQZ9OsPMyawt55dzEvRM6wn7l7Tb9IleIm
34Koby3SQSWMJOoMa542Lt70poUGWopE8b9toY6H4Cu+46qfsN/tZO0mrK/uhjY4
xmomeSpRZcp4ZhMB3EEWjLDU70CZb80MDiVYqrioVpoN0FRz+HzJTZGAYM6Qcik3
sr0iFvut7pj2WWW/njXKvvpYo5uL5fkYYyLmpcSyXYsFAzGehfIql0OXZFLppHU7
FKOTvKDCyc50nRxc5Woml1ZctYxoYsP9ydfGS1INUqLqpL256lDWwWk0aS79urqh
hD6h7nueTS9AiakAISW07llABWSPhpqqiIbjyRsxCXoKZ2CqajTjQdmDE5C5gy7Z
bnlPVQd2O/gos+DVQxWJ9cOw7MIppTF067yruSe9UyI8D0JSY8dacYJTdzXsqU6D
USk3Nf8RXgTkyUN88mo4HQGqATSHr1UbHnlOU1b4oU0ypekzsqTiOPFd6Q2QgzqA
d4H1HpLnvh1tZENm5uyfq2zvc3g5S53HRn3+Z7t0aMK+IVrGUnzTJaaU3ed4tgT4
dkHwhQZgRH7p4fNwmo0WVxABZN004Sz30oMRUzfFMs7fE7ecJwU9P4oHDiqrIZ3F
CqQV+MxrkSbsNXi0QdqHMmAvU4ZgMuQKnlxbZjzK4QwrJZnsKLIa4DZ4hQAps/YW
v7/DCN4M6sdVciU0VKfwXGr7QcfDipTvdMTdEERA1Qf1DxaN40BNNM4oeer5K80/
szyLOUkC3GRdVGYZQoBCi/5CxesQ5aSABh929uNZVtg7ODnTLrRZqLHRmipHJAST
6X43DEH3Clwr5KQi6Oh28h6Rpy0VqWfL0O1UFBXWWMx3I82c3yoPuvIl0oDhPGIv
guCSCGkg0HJeMSmuZ4U20FaWpssELfh8ncD/H8svRr8=
`protect END_PROTECTED
