`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXFA6ddIVi2ScfddXbuJUFcGAj6bksDWmb3t1U/GteKfZRJnAaZCQesA8tvrnx2n
93gTDGIR0G29GIrMRlEUDdXYS3N9G4+ZnXjiVQEYE2+qvt5FnjW5ODFLe3NLXLrk
aUnHleZyYESKwCVL8JScy+K/MvfwuF1zRGDkp+z8T1Z7tiLAhPlpwo6OpNDrChWy
WmY3Wqjej4mqM7dzeXLHV44sYr3SCOPSSEzo2kMc1Ko5zatL/Ifv9VYba111SMtM
71OMnRKhxfwt6Tmii9ixpykh7ecZOHERQk4mHBqJOxF5kHcnxp4ixx0lle9YGvwf
761W29eY/SFJ4N1iwY86Ypfv5xL2tRJxuNahtOU4NTARt0QfHmPSGS3jJz0MTA1p
ouw3QDZEEl1oZF6FyOpd1p9wXwKfHJ0gHkh7+y6C2gB1RtqdjdDv0LpXZ0+OI7DF
daehdIHgfPSR3g7UFl7UE3vncXwsiARr3F1qPJYITOsl0UklwWg4LUX0O+47V/QF
zcIIwOFcU8xUiWWrmupdNipxBOTwr/whlTyOPBw7c91vFJ+F8qP0jacov/5oenKm
v9201aZ43xYb56lzW2N2fMEXuHuCx9XDCHAlG3k8DvrPOz5bi0PXmUi1+/T6ajd9
b1OKSaT8UMcHWa/3ubyGvqwPtsEx35aj7muQX3JwN32zqP8pDnCqBQenGmUKI3jx
avR6QNcn6+fmVPS9otvBbUpNv7wov/mmnlBuxMFH6XjzWITrrab27j1YoEy2GYp5
sP0YTukDck6zgMxwTs2UOcnO6oZCUlHWBtzA/q0STkoTwf8Uea4KNBE2LThhbrh1
kJ96VbWM0PBBEZQTLDTGs0n7LYE0c+nJ8tUexc017JzZJWTBB+zNfDLpi5Fy1i6W
EKH8L080UGsWEDTKmGGD9RphVVOvtS1Nn+3hXktsSd4dV/Ejv3r8DgrfJbBgXx6A
HyA7fnn2BJt6w5ksQx8a2xADLvU1v3Un3sy6juBQIE+0Q6+B+tP5ga1ap1ZmFDFe
RsA6UuQ4fVKLnMpXH+i2O294Ly2HMVsteiUJ1UgN9HTLrH6OOaYvNHEBTngxnqqh
NcnLV3usli/JtZAULO0cvRaaK2OP5LIfyO+/RAAiuuwSzgDWuoZOt0vd2Va7aL6W
OsgDY4jzH2WqJ5X2r3nVMLRSDUzxrpPLptTlVtoOOqfeIP3Y06oIBAcCPgkSP+aH
QxR/0nm8CiwH3xczvYhiM2bDuVTvInPeanC6a5YRuqzUIFv5IHkINk8tgkXwDS7P
2zEP3kOEOWJQqnse9Mn7oJ+v2UAQ4/3MYd8hISMiFDpTGqLX+uc/7HZdSBr7lIOL
eAcQ8xT6NrrqeZDrAbmVucBQhNaOsyoH1CClrPqY5xpTkS92gWOQtlOq3FSokbYf
oysLFp0d8APaX260J/qxSLWuipAH8JhF02zXSXwpAO+bm0VjCI8twG9o7D1F9th2
EPJRtR53JVZtM8W2PydUXsxD/UwYfP5bMl+zZqESBO4yWfSoPQ0M5O4RYqgZGWui
ialXdH3XTExAi5rnFkxMLw1pOp6MRqGyFBvJ25uyuqamoF7hfXTr8oL7T4S9V9ZH
LPy03EyaM3vo+fmrhN3RzFsBEBSaMSgWWnExjrDPHRj7BKZrluEvEDUzflFRo++x
28KMMDT7mTrtBvmWC/BxH0oBFqUgRq+7DHER8y/MZgaejHDwIgYqehzcV0OWUU7M
RVSkwU/Ppxro+0zWyMiBZPbPW8MGE3NNo6mkMZZHR29BhX3gW0XbWUhl8kukHW7I
R4sSDXEyBPyC/4om11TbyTgDgIx91sPflrJXeZwnvYB+NoLvYbGUNE9ChLSDFCxt
4Ln7ZJctg+8rqVRX/eISWMINjFs4PWIh1pCaKV7uTMjqpEHcDUHFjdUwbGGBqWYs
JDeuVGTYGAAXxoLjkGhFksgQWfO9C83MYQ06BiFWbNhJFfzAXO+NMMKYC/HJY1YK
dKVOIXwvdakote4bJxuqsuo/xYO+zEl5a5TcCx/Gc9R4dViGryULvcTUgYTUSdrx
JuVsn79dpGDkZvjaPyGD4rJMxWmsANUemJPX1szUSz1oqVZUP1BligB415OHM+5p
KEKe0OUs9M+VqsYdcUpVWSe1ScUxVu+qkZnbnsru5UvBzxR2IcKfBmkvG9xf3QBu
6CQ7fOMxuvX1PWxakJMksQba4dXVqc0hfP9uHwxiXQSZcFTvxEYaTXlvblDLOlaO
A2U5x7Zgf30DOGs4frk5rug8E2P+d+4h697Y1x2VbrlbSDIpsLZzEDw7iuxdOrx2
JVFa3b2MK17/iMeZ+jTLxPK7oYha+B6VlA0oR7vxm/PRecOvq9KuaVnF5mS4NGrU
WrVF6IB2XiYroerAeKyxu97txm9rmSo4rqP+QwQEYAb7iHy2et5de2PD8hKFbca2
nLI2BNatknvoGxyFuHZOf3AdFdtXyxr8c++Nrm1aUu6+7hfYzg84NLkf5ShNnFFq
HCByIM2whpouH7hQU0v51Sf7gTwCEvhOzuorPIz+9nwDeGsVStS1lUEalLANjfCQ
lqz3rz7X140kGrMKyv5RP3gBPWn0PauDjaSW2rekfElyiAh0nWcNcbioflAPvuiJ
S+hxQYBw8P9J9rkVjrGOSOTBqJMlhD/vz0/iFMxhS09y7SMoUojS8RKCY9o0XMY3
vOiJxZIEiOLSkc/vWwolz6FbCxZi209Q4fCG2yX/gkT0Qw+lM1a572KfZx2VbHAY
VilSZUvgQT6ggHtFgR3BSHft2oKwYb1vBFPFP3bdJJuTtG0JzNyKeDo104QrS5+y
ce+X0bwM5pt0Zt3LC7aAH8IMHJoc3CRVDGgKZqZaFWvmG9TGjeF3xaLKhJwhCwko
vnKDYLa6Lx+uH24tF8miF4iExigMcRuczG6Em2AboUS8bLTOXoJYEVhNxNM0nL5I
y3nC8iulzqHNt99L5Hjnri00bCAs+cpHxbvYEFN+0SSPv5grl4SqDM8dJLNqxDco
+JJH58AKumYVV2kVoeWsrndopLc0AzJ8aieWvqOqzEWlPdQ+qWJcs+cJ9gUu1zNu
pdWfKmJIOtFQ8NOzq/ymcLhudD1eCTOgxz/483AkN08/dVrFeyZ6ALhInfIAkWZm
n9jF/E4kLpNFbSzr/s51wZnHdlq0F/RE3KE2a+R0ZvnrujarHi19u1fI/MO/5t13
T/PC6RytsLtMEIkHxwo2xY8uXNSdKucnmZO1R+XHnBkhlCMgQuWKwGnSMEE+UPi6
9k4UhYgyIddua1CwCJKuugNRvTjWH8/kNEZWZYnzuIk=
`protect END_PROTECTED
