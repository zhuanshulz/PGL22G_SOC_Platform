`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlQ4oq+71ERfi0CzH6TSrvC3t2Yr4gO5kN5GS9J5HUHNiGrxKw5T446c2QHYD4Yp
Kpb3MFFsYJgThafSYEe7z7JjzRjCSQpZM4Ew1kigh1fbANcJOnbk7oJkkArob8CQ
E1qWJyGdwrLKccYTobr50m2vwAKD7DVCzokMl6c6h1HF4O668U0lN7cAf7Ludke+
EfnOMSZqtRNFI96VbDXpV2jCwTyVx/nmMuO6qViJuUloqb84JlBcBHPiavU7HU2N
gz77o0vrILvN+TaqZhm4S0OZBSlwf5EZVoTnZeEZMBPTLIO7fPmqB951dU4ltjTE
xPTj8nwUH73Cg3ZotP57unUgROwIMW8K2AckUpVF++iVM1Kdx0yERCqBpPb+tqjJ
KQzLYsTkerQswQFs2dBNXLbgB/g1zNUsTucpyFOcQMtPUk12p6V7ELF9AspnwjME
JS11XTcM4p9ZLdw0hHStXXmsy/MH9TIVYaWbh9cNonLcdO/8P51T6IBj0SeTe5+x
OHN4U8GHIAEAQcwirKb5kxCIPh0yU04oUGt6OGE/i6UJz/JfiMQ2cdJcQPCOzLbZ
T7EVKmL28AJs4JG5l5FpcMSZse6rdJJ/OShg3EzCWCa/iScNYLpgBHDhPEAmtuHJ
K+KLIN3sXahaNGR1N+cwM4Xoq6kOekzDwWICPb7VssF/RNkxDF/8NziSITzUppLy
dUYAMshWNoUaTJGEESbVq0lLGpvW8XApOuFjspVPyE+890WRk+S847EYhLlaqprt
LO3eNX3JjOsm19DJrT8mzY19tAeq4/G3W8JNPCYo9a69WKl0ejTD9ZdZm1bfy8Kb
cjd2HfzcukrcIcCQ5Lst1LFl34Wi3Vj4FMbOmy9IDyS0R88xb2lbrYous9YMe3ll
E2unhJgj4999eJ1ObqvSRZjtaGuJMSJeIx8wN+xmCpF6D2AmNL2Tydd4lBi/P7H0
mz0mYA9bgfa7dFOy5QotTY8/PBrAWEBO3R4GkQY0bAW9Qn85FahE5ul+fp8aWlAW
deyIw82fD0w4SYFkYagehqqqSgJKPrOWNie4DoeRM2uBIjxOHqxEjrDKqKsCnTH+
L+9O9HXvMbhc1MvyOBCS7WzpUEmyBe76g+noDLrZSneD86G1btaY+p1d6kaMfSpm
p2cSscsEh8ZvsECIR0gzzKpeaI7y0FcO/v/yJmb/JP1vDANzLVjsIR1wKr9E7GKP
lwvDd573m8EzKCkDP/y0dN8rzjBynFftFaR051t4EU6y8jjyNi5hh/8alB/yUtYS
BIJjF6qdLdTmwf3FI2PLm3/NpPDdUytirQ92j49mLnQhEUvdaDqBKmgLzx1VqjMK
ZjPrLbApReHnpCewg9xqKX1j4r0hKJ02EtkSHgzmLmPErBHLVyzh74SEh2YMT0XP
h/Eg8OOrsthU9kDdJvaNmyzLCwfzZsTDEWzvcogMnW8olrrB4Y4E704ERVXrD2ys
F/Uw6Wwa2VFfeSvtYt5hRc1tgZt5IP93la1dMhdXJGYq1xbGZ02F+KRvSLNlkwFr
LoQXR/+y+QcjD7qHv/NJGeO12eiatI6mUNhvFLysAhikO+rSTSDUYRNJY7gZg1yf
DwWDQN2h5o9SbP2j6frI2e3Yrrxx13AJowHnNsO9gbky4TGc5mq2imEMRT/ZSHKW
AqPnMG4wqSw6AJ4rqRJp8XMtrdiYxIJQIRoDzhnr95g/4w82+uGskzu6TRdiqdB9
vnZFgFMn1gf/BWTvEbeT36Vt7a4tUebq6V4cAIsuCvrO1Z1xqkgIRe2OLV7/io/2
uYTpaptfYyT/LmoJdY6scvTa8c0zfPrPq1NQmBOe80tI1nTpICGe5W7l0TWNdGOt
C2EiwW+FCt/QzkXd70w5nJjyoo9VIE46swqCcffuGgDnd9QX52+9vdeJaGPBR7tU
zMNNE09ILDqyo3aH+1/08oxZc7hf5Soitk2A3OGl4rGPtZvEuffETB97E2C87kbA
Hw/HW1vxBBt2JEKPmDMbb0WFywkCC0iPDRBZ6lvhtSUOXp6LoY5a+J+m9PN52rgQ
DcTGeVTTtZvKOswp6En42fUJWy8r2gciHkie703o9JhSqzvdiKskDZmCu1cvhWDd
iH0BMNPwKZMzIaHrL5ICiVJ8Qr14akwPEMz5vrs2sqyH8+f/GnMkFoQpAmt/15Y6
wJPBV4GfDpOKkjsSZtsNNfG0aPYX2eLcROvfhXifvmfewq/5huDe+IeLDt9vwhIV
4EXd34oxix9Oq8XTUehmznzAlpMIIAijwreZBj2AdzdLjUjaA6oUYfim0UTbyPpY
T8ch2d2NNvxsS3JGguz8+DyTaMI0Wzeh61vQ3SSkTPoKfXnRebM2xrhKmhz5PG2B
ri5h5/hul5/WsJ5IKmtGGA==
`protect END_PROTECTED
