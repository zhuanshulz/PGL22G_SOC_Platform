`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HW/5NUusfE14ZhXqO9tSIM0Wwaju2FtXiknVG/q8VppWl7Zh5TBlrBKpZySN5tgn
zTMku/dMr/iBJ61Jd5TSFAABHcK5qVK6Iri1cG4Luz3gVt+KE0yE0rytUW+X5+U5
JsYf4lkOji71Ojh+w5TFq93Lm2l5SJ3UvuDp3xZVBWcJB4vzDP27PNr5kijYlsAa
IJY4TXlqWx5pSjsSu0FWunASxf2NmgpWN2mECQvH7s/LAsi9KaDAXWPfbgPMGN7p
Hr3xmgkbf63WaoSOW1f628naTpodnCABZZRYv1x0Uv/4iBmnZ1kCDZp02ZLLWj67
UJm+bzBSlop/OOapUn6LuTEYn6Pce5LrL1xQoghO2/5moLh/8HPVqXK93g0+izbx
Y40+Lr4Vlql2PJ5vmF1TT51i/1YDXMy94cz01qGLzZO9rUQMYd4EBnhgGnDfXTcZ
X1MFm2i/gY304blcp3d6Lw==
`protect END_PROTECTED
