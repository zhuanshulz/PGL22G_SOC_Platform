`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CksB9VZ6lOra43lQ0uveJOT8pUOjDatb5dZJxyXX3Ff9nZTRC2NJl3qivYqWLwGp
MavmH+6+Ojla8eYEN04w7WN3PtUr+UVvkjd87ps5X5K/FSrp0N9wT1emxrVksHkA
PvL6k1pC0/zTbUJ8Z4UK8wRmdeScOgZRsGuRNho6drx7WWmhJIzWkc4nuZh2Wr+I
F/KHTNxIFzsxlD5R2KIO2OpEMMmBVHPdJad0wuCgaFf0NiSa4SFxz4GiT3wlhdDf
o4dJLt9BBf3BKf/SifKxh4ycKmxxlbwF1vBpfgrSYEnBpt79CFeIStGJpipWbOMq
Tmp3I8yokqUUjDoc8GW6EvcW5i8YDHf198FiO183dtgzYzF6pt/M91F+BSHQVXea
0IgakVbRIWsFAS1nYdABFmhUGzp3idLFclvJdUy0mTDScxkvi7hvGj02ZyXiTAJ9
5kAtSZsd2IUzhzPnuU9OydFCKEvl7e65U44qQLyq+TvyIX04fhnzWLdypfCBCsev
J6K1b5Tz214s4O6/Mvl14eo92lh6RkImpJkjeFwdHboqKDJhyrIKL5lrG+zL+2pc
iUrfTjJxOXWQCOthbxnJl574DQQ6S34kRgEej/0xkWGapzpX1/GkvEX5ktJU3Itv
sxfkFCr/NFCrv7KAYIZtx6YJU1wuOhskldgmhhUemkHfTt/plnx/wBzBPIqA9Iwv
E28CWWD49NwljJx75iGi9cuxqQMc4jV1sMhvBfjcomxuNdZojsRoz9yn46Y0LBeF
K9rds3LrRW8Zx12lYW61BdmXhYay9FykN2FJpTAJmTPM0oYkUp793Dx86h2d8qTv
ECQgFud9nbJSj5Uf43yjbzy9JDkJGu5tiDvWzMfbbipyrDAi3usZIoCmzttKCu0W
yET7ZQljBrjUzLs9DdJ5nlWXzn/V8G8y0IMg8aFlF9R+Ktpy9Ga7zDrQiMIBVjyn
B+uIYmfY8fwNgJ4XIIKa3HTm4Wvj1F1DXtXA5GsGVB9Fu4xInAfPOf6IJ/AaJWv1
TjDsoHk8IlyRWIxj6W0VjsCx1FMfGsvm/MoXPOPL2af3gjaF6Z9RHcP9fg8EIYY4
pBQ1EomA5ThcLcQ1hD2OVUmOp0VoxgWdOEEeIGrON1RJL1lAQFURi62JYOsT6qxL
BQZtaJk7qD1p1veOHiHtvWZkSPUmauJNNFPG3+g/Lwv7NR4jReQjugibXeA2WIge
yjcJfUICfIctHCkJ9JZnaVHV1R0M909+7aiM/9ecGHtsUXlmvdajdpQZ6lPmOvHh
LZCevkzXyrNEVDaBkrM4PMQrKu0HSel7TdFvQ6ZHIJkk36y0ldXBmm0OOvMctdUv
quDjYqwnaWxV4utJrCA0LFP2wY17VnyWNfEG00WCSlclCQ0i4B0SYCT88Vl+lYA5
B3Jv8aB2YbnLtPQjlj5yylTgHttFyAttuWoPqSYSS+DKbd6SEjZ22lT81uHpkQDB
834Q7I05aeM9X1/gEZwpQADWeIOh9Ha3Z0jW5ox8e/s=
`protect END_PROTECTED
