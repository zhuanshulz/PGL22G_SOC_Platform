`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DyfF0duZaRfBxioSZ+oRehzTE+UGznKcDxxkaUeVUVlkodPAclXLz6ppuI3qf4wb
le825/N6Kk8JkfsDAgIXxq2P0mSR7OXNzkJqlOEE+v1mPjqgPerud6uoehwASD5c
J5uvU3ImSoKe24lsDe9Oc/vWPBBhXXaLct1R5DBw/Vv0tS8DzTAbCmkzq/Z5H6Ep
TgAUPKKk4Ad2iYmytZ3xs8A5PWIsfLlNR7xEmyZydHKlv02HZHUaS1Pk5KOJEVzF
fb/KS86EYqCB9KNuvxOypIkfaZZquItkMkqz/hnX/EIZBusAcKV1YnuaPXlQQGFu
vNr3IXtZrhqbaMpLtETuMR6J2q8KeSayeCqyalXQqrsSxFQkNZYkRr4+c5J4g5kB
Kv1g7BBKjYm7Pk7cLBL2XZxPqkNVITTHoBy6rQEYZFkfgN4htobFY+ToW/XfTkMA
0DOa3V5Vx/r5INq1p8pAeyKGV6ZcmJUiYWb8R/HKm02nWHVJbn9yQRuOIqxDQrht
IvUs7Z4dFI7m/BAyIrh4O36hcShxIFBplqQqUW7QQcRXEl5v9pgnCjP0ToXyBJeP
prW8lFt8miTzrhVLEmcW8hyJhnbjosfVHhWKYpnvc849EuLiyAi/vaGChgeE/xrT
nRz9WoUduZbjUufb+CtVsORxGBBifrX7FyKHqbBBKBZqKmdjgq2tdYeUlNxyOIMr
KuTHDIaRSKckd4N5RLdR3hlgomVGBO2U4FyalmuhX/FivlP0MUIQjLp+mD8VOZ8/
O6VywYXOjVmaOYTZWl63T2bO/oF2oM5qR07tbqWeVFGaAbq5q4VuYQyZK4pfaON8
vVFPPei83+1cPkEnljekZqWBmgURrFWfwHbQ42u23tbHdg4AXpWmCzxtcEtiHajU
b56c5vhmpvrXVOQbsACUgyYUkrfQrnicY2QsJzpHEmm6jMsqb8TX+pcQELwrVXVR
QZXSsITVAltPqCC8LeYgs7crx1hNkZuUaVmsNx66J/e5Gev4GCd6kdXnmOmJS0PS
cmONX6SPIhPCTB1jXoHSkaYla8SH0/Tv4CfoqBHyseY7x2psafEjQ1X2s7yIsRIJ
sqYp8p6iQl9SLZZ18L/zRH31y9iZHzkxQg6y0H9wpFKU+CqtT0OXVX9L9adWOAQw
6UmTOraJdMsG6sB+SMevIC2FCAWi3Z1leMf5fApmazQEk/fHFRvgqnbjYFuH8dpN
Zyca0IYOZzP8oXFqeU3e9vIUb+dB+LA7LJqcVAf4fP96yQSfSawLsNC2GPb4w6M/
oMEWvlgMxLk+SNIEIaVG7vTCjryyfBeayqWXZXbd8hbN/242qSM2DmpnoCXwfR6J
nt/LXEoWfFj7bSF+h/od4uoxW6/T7WvFp/P3VNWCPGjMnBqZFJ4pet5R1n28JstF
9NMpwSbAmQAWe0M/g4Qnvz6ggjE6EtCHzv238wwMV5AyZqYW2bxJe0DwvK/S7YMu
uj3DQqxYwwR2Y+f8Fs0IcVp2NYv1w5xrhguX/GhX2v4/7luP3KvTYQ8fG9HlB5Kf
s+P1kjxKpQmiht9AQJgI18pqwo3QkAzj/QweudgLCd/EMdD5cwIALsQmskB9RMby
0a01yU45XoZpjpY2UwXiyF3VoU0adKXmf/efcwesfl85PCo4dFSXUIx2AOyNBLcO
QuSx67fEWeddDgF0WVBJ2GAhX3aSAndYSrfuP1RIpU3fHWz8aWanVx4gEjqmHmOD
G8kqWE9eBub4EC1FalxB8GlLU0KdWKECm/JN7XYVw7OLcNeF3rR3iLTqWmlvACQ5
1JILyPsB8e9311ACWQpBq/80cSdauiNexpPy9cFVFUn2FdVZnN8J/F1rYjnE9afm
3vZsVIew70fLCx5Ht7/9VRMMtapu52vSBBE4ZVUP5Elrhgt8sovkM5QQePdg4sFu
F/eGTHBVLjRLO+AVf9E2KxFb/VroEgZsLsg8vGVlp1HHmiYaO3awsBSj0l7+SEl9
lUKj7SS2luyBCe1YPGeMHWLDrQSibZ/AYhs5hpLlbCBA/Mc+IV5oXqRqYtWCAEjv
AFi7RaRiBC4ZsNeGVxJjNcvmtOeh42VKMzY72/YRtf0evmxJ/QA6HyxuB0PPNys2
a5Qy/CIZ3N3xIQXya+ouU6+c4dfF7tekeAzwGKllhDSWMJV2neVgFTLTYSSJfRGn
drjqUhIMMW9NnbnDu+5EBJcjJ7iFfNSMTN+Q/2ovsMrNcnWWZXPEnGstsyyBxUfH
214fFvtd4Y5pL02II0bMvFH/p6z3xZofa5USwgWsZ4xCDRf43SpY+aYPWFMidSuP
EtNJZyByLjXcKHRpo9IFqwcLQsnBacJ9RfoVJBsCTOlzemsL1Ns6qf/AkhxLilS0
`protect END_PROTECTED
