`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mLo661LXv6+hTdYFurFqwmqb/iQZ27+/Fol4q48W7x9Rvm+rc22mhnL7jR1hy7ab
h1sLfyO/QGQUw/ujl8Xw5guGQLAXhpTnumqUmzfpm37A1BDI/UZtxO0rUOlEc5Oe
pVq+Ndkd4CRUbst4IcyOveEmKD5wdRDIHyswdAKM/fVvh7Pb0IGDKBshFgfyMuvy
Z4sRIq6F33sb9iYGmGlLPDb5Zx0F75TuLyNX3ymZZ3Ch2u73r/W4NmMtMNipC3ik
PhPjo1frMbwf1/ubLd5Z9jVxfj/9hlPT4vglxsAxyjKrf/mpGvoYFNDy9tUD1I06
lWlNqufNUTmpv29cOX7ZwJErK+/N3z9qjkkNtLwW11zPVTx7bjiLBnd//PplHtvv
RVLi+IOc8cYZP+s36DFf9NR0pNE3lmZg0VbNijmirSseqDEzhirXBR4zIGfEl/7b
K3Kp8o74IpVAVdWHVlhX3qdxyirqVGA3CnDBsSi/e6zbOj/ExF0fTacaquQxaPZ2
auTPSZRb41qCo6m4LakMK8+KIjLIXKIXnYFey0Dy4gzxVaWKHd59CTdriltef1Kt
YAMEAqbNNp/3UUlihFlpZSQHGo36zlVdgPSzXnpr2U+35ltW3GKFEYG8wXVQBkls
D59K64UAkZOZIxr6mWQZ0+bMYIKFMvGSNkwqd8UxmlnMmQJUyPKxd12ZayINNsho
bT2hfvPqOGnNnria6WreHu17xqQgw1jn+t0hWd4oOaW9wvTIHWKWhnX8UF53+vYl
eiogqHXimOn/Ru4qjLKOeg3J0qQI7ArelFaYov3J+pw4QFEq9zrYhjrYtcl96y+/
0MmBfKmoyMpud2elPX85QIhibtxr0aDvZKFu1WkfQ+WlsLRQo+zYGxY2bJLqepSP
TL5wBRgJhqIFAzXPBoOpNV1jHZMiSYb2IXwNTAT5uqqbJ0yvscBrkZ0xCNQtoxxm
r2fOn90oR88RlQps2mFLv59cklDjKaPYlPmwgAzJBXskjdH2SF9PdnDLPPReygVQ
GGRmu0omuiF3w092M6UlWtdiHaoQRC3W9k8TjPKPnXKTdj+tTF5corxheSfyZvqT
Reul3t0rhq9A7ZR3iukbULtM7Ki5s9Kudmv/yErqqIvGwEhMCFbdL290emVxQejI
gO/7cq6V4i5tfoYCw/NX2oCynXJE+2KzbrWRelai5KhK38d1Lp7V0sSA13uOqfKJ
xHbRO8eZx3AwOz3KkbuVCiFXpYnLip3JzEoDVNY+CfyV7vvKKQheh263ypJboGoW
Kt9HnL3DC38eVNufgO+xRkx/NlXycL5EAxo/sX2uKIQdQG1QoekfxpEuOQlpY90W
dOZN+A9G8V7xLI8VyOL8/7qVXKaTSfiX2DZF9INjGhA=
`protect END_PROTECTED
