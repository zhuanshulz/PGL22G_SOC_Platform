`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ooztaI1S7CsqlcLAJKVjXHUmfI3FrqR08plti26gcj9UW3CdMc9AMjFP+SLukyq8
3mLwz5QdOJGgJrTuombG5Mxy092Xe7hkyEyp6Kj9GWH5C79DIppblF2GiwndbRgH
ROQ/+zVQAtZXlxTmtOfRQmWKNCi3Vdby0gVn0o9btLJsKN8fZNrwX5VzczbNhI/m
JSGkoli7lPeinLlLogPNvhU8g/RIoYeymcyXuH/lF2f6LjwCQE3HwetoYUGK1emm
8Igo8z2JEPMAHJvpSCSPVsrBmjZLsvuw9rM/r2bLJ5KINiLh/JbGO2N9HSCVaIID
JyVFiDPEsDuoWbhUvdjIU9efvWWpJiNBOr6pKL3GXu1dvJSEm7StoXEmbuxuIcDW
TjiI0NtBw+1+PlIFQl/28fy89KZ63oi3rqKfAqQFNclAuoAF1xLpPsB912HRYXFC
k5UK4Z3aN0eLBs3HOcmjTP2pZVMUyeL2qKC2iO0PJ/kpmNKPvdRX73OqcBv/1sPs
B2kbIA+HLvVeqLmJJNgnhNxwkkc4rG5HeMr1qIl22jYzmyIg/65Y9Lc6i7Kv9f/R
Gnnlzx9+GIUCy4yHWXGHehoQO8UuxlyGqvUxyxag4lUbQIUmDbY7dQ+CTwde7YL0
FW+2Z+vPcwfBhSgGcwsnt0FEENAjQMWMZzuNopQYJArDIFnamWcrtmrI4JKYmmWk
37K6/6LPquiGULRLYSgvWES8eettwR0Q8XvOos2QFX8cgAWAo8xnkBpNXBywWOOs
acvuMae1hOmYaXDPjjeKVwoo0ezzx3FUKOsCu7hGgIQ5p1kqDoT/CFGuu2FXg/WL
MzfOyqljfsx2gahJ50igNeGCp7VLiQ/HVwHNXqmQDeA/395jKC7Biux+Cu2U/0Z+
I/Fz/DdqQjhl1jLmmYud3wvoOaoDcH61KHa0k65Pt9uYmUUBxmA35YKNj15fR+Es
o82xvC5+OU47YOI5CYRFbPIQhToKNthsEZnWPdQ575A5szZwzBRUK0BwgdoYIuaZ
39RkN/l8Sl/2Kip7y+Th3EsKRpV9T5CEqtnX/wGKjBiejYmGnr13xbGfEr8xCOSa
gD3CHpNZ1+9ba2Yw3AP9gOiem/m4uP6AFohYyf3akmcaZLNlSu371E0X2Az8k+F7
dGRwaRCSDWrpROsEn5GAjS+w9S0+B+8eI3WEmO+a/L+EbnBqDGsGA77VYj9DqWrC
2mh3DY4VhjbBDe5IwA8D/Xn5ZcBTMBjGWS84npkQ7mb2A3xkSXW12bf+GpgQYjWq
PYg0TqIs5rJpLxq5MJIQOkyzVeyNknzLTgEHJ6CcPptrug48IFyDJUuHDKfw33Cq
Gd8vrgsx2vbohC9T9ln4rQKtFTlmREQI9HZrJvz8BaEl0CToBV1JUOuar8PXdKx0
1XpTf+g0EoDjFgzOxd56aEP0t0ORxFR5UMB/PUzfx2Dmk/oCOzQfitlnAoMtUzuF
ap80eButJzI7XfUDgj0ZbN0LESZybnDE2zimQM/MbjzXAdU86lV0z85oJd8XqHHl
VEH+ERC8I1qzV8THz4Jua38WLiBDGIBDrwt9Q52Ps6kNH2xhPSzO8cQZdlkMu+IU
ysn5wFLnoN8+Kp5fKMDh6lLLs+QyntRrU0cD5XGSa1PdeUH6dym+0aU5cCw8Jx0a
0ms+C6JVWlWPxl8y4GhCu2vmbJjDJeiB3/YRt3Fv4yxu3s9/Eu7aOioaBQhf/dcZ
z5+n1i6b37UUDvTzgtTwk1/4ylhPaGY+Ss6gr/q34XVrDJIEVmyT6ypj8ngr5NIH
+wIKQ7QgJREvx1+WItrj0LZi8tnvrJ0r2s0FubipMmLcoskB1iDfwMo2c2fM29Lj
RCRxPO6Edk5ASolBXzACYnt2zHoLTs+25ApGkRRkwgNm5WZzrWqfCBf15ZsxFG51
xTNM3DAnNM99+swUTLIhLbuAWbB15b9quEHQZVoiQE/hfNj0Gc5o/xCqc3zpYwfv
DU/sUqVQoDraugYjbgxlk/uQSVKthB1mCt7SSIO4+ZcrZNtFCjbvjcUMPPmwydVD
DxagCp/D67iSjgD2o5lU2yZlOhMcmDAeWWxee7cRtrqhq/RPp4qiJDk86/DrNHPh
UIYe/VURhNz/+1P1HK5dXy+lBF/WZziMkaDQdhSuYsV6OxR1za4/fdP4tPPdx9Ir
//yTeJNJpsHaOpHEjJoWr6rF6uykEJuR4XNpbIUO0pppBduak0AU0zVBPQj+F3bQ
THwAjmDW0A9MGbh/v+8VaGcNOvoQce4WbEdBnGWWYVignAJdIjGf4vBnhtYRGFoD
zusmt8ooU6v6yCFfD+lcbqQdnSV/poURmMmyP9RpSyDw/AZ1uAe1IRKR7d2am9nY
vxR+JCLoL6LHhsi3GMkiw2HKvWSMsLLQcY8kGoBSrAT9vAFOLJ8e1NzLvOcaoJ83
2HYLFS1as02LJFePgozGdvRjXdoQJC++nzQARR09i6vt3RVsm1BlfexJrnuWyzcL
P3a9LeU0fGsAul+seN48Nc5i6O+zM/bbO0Z+yaPgySgUVxncFKn0/9ALyplgLlhQ
uMBwbs7N6etfyjsQtqh6IXYShAivdIsZJnCRNWyCXerFXXDZEwBVQnLeeKCvfO+d
u5HcxuVSkZJffQRK9M8Oy6WOGMhgEh8vvcC2GB7eFPoIx79kBNoEHEdIEgB0TXUZ
Mlryj4ngEeq+8n1wL5JycwtcWxbyI5G+L3nJGrBI6zomVmHPOuomtXOjknkD2mKT
S6ikxVLoIb9bmKpWDI8uWFCrlHn+sHmMU/q1odzhtfIEtMd8wb3Sh0xn2Mqxgwms
l4LB0062JTd62Z15Qf1twKYnHnRw5o6FC75k0nThMTGJwbtIW25wM6e/hB0cyj3B
PWU9a4CRdjmSpg/S5a6l2dyCW/9bZhFe5lUB8QCRDXHqNBm2I9MUktSqO8PXL8DX
1kN9QT0AwBrqhtAjJi/lK7pb1+k3PwaWuTeOXUp8nRSC4/JZaMSfWWbL5kGpf3RJ
5p7xjxIeSll1xHUsZ0Hr7Hu5VmzGnsxsAAv4K3FcZkkjD5kFWa/55Z3nq2LBrV7I
MOVuSs6qjP33nKmhdPCadhuq1nf4NVn0k8d8m29RzsqkYv4SJMyac0JasylRafNA
rBglQxnKsn0TGkTCQKt0DlPGymAkfu0Rc3iqnfj0ErC4/sSSfVKbKoFxfCHEGB5b
KVo7EEXiSnMGs7yZcQMWATj5K5dAAj/l4zExGxX3V5+ZMEmFz4KvG6txRxtjecNl
sLpDaCcOApVr9nCVaBuHHaWqLMPY8Jn428ucGmU8L3PY0OMukf1wfCNJ1UtQc7ch
/O1Vy8XELzwrLqW0eCIPjQ6BBYAx4s+PUZvMteBZ6aSLDL2pjYxnt3EfmQGm1i+b
HjmrRk8JA+gz2rbUvPd5ADVipP36UcPDsHmnXe0mTYIE0J9RkQfN9oaOr/UfFyI8
xTzZ4DFyCgV8EPeW+DTmoObfwleoO5yHv8hCJJjWdg80feb5KtQ5NKFjngwSXXe3
e2c6kxv2KCGn6kyDKZJreRr8IW9KB9hm/gWNhwveG2ngcsmp3xsEzhLQK2i4LLGj
vV/It25emipwREZ25MIbKd/y8VZUEbTBO9W9iDhlf/8+Sd+MfFEmbEaTpZRQ+vPp
/+AdSrLeXQ7mmZWz1ifAp6XARmIGA0FR/fwAiN2f7yQc7IaxyhMsxuFYA1LQjAk3
vfAYrMjvylSPgyr+0rfHbl+8TU561odpK6US9FOZPen9CfHG1QudjRRkcdl3X3hq
HMB4bEWARTIuulT4ta1+qvmUGsXEO1Z3PKPu/g74zmQQOntxHpOYMoeU+xvM0t0h
Tj32HDedpc5RoWkc/RN3/v7ORv0vO5UpGnHvEJP4xtWbjISqGXguhTVgkRhIfXER
cvngmlGyePV/m35aKQvwxYrfwWqnarAENI/VlVvcOlJ4XGUI91BEVfeO75pe6A8m
g8YUuWkr5oS94UlChS3C4mCZIbgOQi9hbN+ZkhGpw4fqLO6X7LpHW5zSod+wEezG
PF8g3C2MGbesvUxn7O6LScLCczq82yLWGdEdkq2uYE0Pmn0IMSF78GOp50meNkVK
iW7XYvSV9CgxJ2/7FarhPEt6MohsMf1ImGkXWfRFm7X2+rluobUV+aZHNx1zmzdi
oBQ2vmAdAU0YFWpFD8S0GhQxkwVYfG+SMcQ4D26Uaivi7LuMBYUHywS2gEijlDVQ
gwihz4jov6En4SjpS5qL5uv9CkM6a/teJlq2qkGvROlloqMUhRgVfOqKcWfK9spl
NrWU8GYUtO6auE4sXRHfqpec3m6q8tbos6T69u8Wta4fGT4KPk3qwkHN+O2tpywt
NfaKbkzJ2RF/w2zevS0w2IeLKNlzxwovk7igiGR7epqZz2F2bgxHYr0zrL67dQ+x
h4ANpIKBb7T1AwzR45Tq60wEsPxBpkjXMDOJXdRauz4njaqbirlm+jTIVGe0ZQ2T
ERZMTcw/DSB28REUx2k5TYV69TwbJUygEqHjSptSNXJLL4c619GDRLPn/bLYdW9t
TLmqKmVGQRsxPRQVqNfr2+dp8W9UZ4RUlz0dPzyGTW055hVexcxYo8WUq9SxKQwf
Fc15zp1T22mzsCqNrF3aimbvy4Lyq8NmqUnXuOzsYJhMFc5uxa7bgkAf59CgC7hE
ZKiS3kOH6D8IO3bLDjMdJ1HRrD4DZ6X+Ci8sgu8X3oZQ2IQFFQ3pJGBAPAneRwiQ
Ka0wF7Z801d40uEO32jxQc26RhAtayYkedzWIHR/E8GNX/FDtKOOMUFSd9kqiHRo
llmXLpoy0RyUsfRHcevzgI+7feFGY2UpNsKrH9pwWydNwerC8/YklW+L82lj2bFE
o8raeTBYXn9qKtEzqWDHw7mw0Jy86ImQICY04A32IvqmrOfQIXfsq61rWluFVv/T
RHJ1ara7dEfuPExN13X21RU3xFfBDgnzT9SDfBiwoBMpwaTNd4yF9MFHnXR+ALg+
1NUTXq5pivBU9i+76KMlwNXUfV31Ate9h7eNV6EqxqtHGufts8bfoYCESU6zE19h
udVoUvf7mwWeKzuZLJ8iM4x/rkF2w+S89inKxZRs7RHECYzMHvbfpKtKtDRae0D9
Js+xRgQCET51zgsvnvgTJQ3XMGl2feK3M+VG1JvNF4CXpAE1ExnGlz1YCoXQYOle
4C6mbMCIS+wx72aC7jvEjgPQS+NWbgxuQBzy9EYT5iPeCBI59u//On/t88f7mVx3
DmcPXG986t/z9/JYpuJ9xetPXe71fEZDRXzrj/qnz2idLoVqRurrx2cOPPtlBWki
rR9nkWWrdYMvPZJmjt4aTGFuzUtI2ORiZZKL9RmCXDxT0ac5VYwfSjo8tzqS5Fvj
twTKUpIo9JVG1T2Ga6bEMygckomd+i//Rsas5KJNX192ZBB6ixz8T34uRAazcajs
kyiqLOm3LlAkKFwsBsc3Eka3jlzaruSem+W0g/7JoZrVi9zadfvowXjE8c1jl3sb
LvEgdr3O7SxFabMUsp5bldh8n/Go5eBUxu72Wi8C4fFNCUSixK3imQ7RfybKVeK7
5H2vCDIPN3yhyj4hWp6WSi8gk7OHRlGm/QiFu8gTKAsgos4GIVMI+bSQa3xkSjYk
uDEZgez9fMBcp2YjHJgKg8tPTbyegtu3FLa/hIKG651Sa0PIP4K3U0Xan7q1OJaT
RWjPZ+sWzEc8ou8TxJR2XgVK+M45eGHY4CDrENwZk6RyrXlEviKzAaVugvxWwmP4
DZYJrrcGTc8UhDYQh/Y2KHnkNvPyoHhdzoNVfYs/Ay8WPtG69FAulTS43mPZQJZ2
dZSjHQnC3SmFFc242iQov4pu16NLWbrwrCx/s8hpGoL5DTBa33gu/SynuhTDlJkG
QITuQziyrXzXtoIvpn0BrJcDyeZIln1TXBktBP1VY5XaU+eABPbvOJaaTaYfOmJT
YZrSkZ9bini2rwDq7lHcR9ilTCMwXq3wWVJRnZ+19kgIOLMpo5g3CU1GSDmm0nJF
iQRQicKQcKMvIhdb+Mua2RIKGsAp+3jkn8UxXAUJJx1tVUR6U1IdEvL+NE7yFthg
iKkTkeJf8hKcb2TN7or616N3ysfHSCZr3w8IBPW7dOKbcXzttrs/LVePeEaG8V46
y/Rv9SP7WcEqDykGdFZEVRcN+MHK0R61MMa8MvoNPA3wCt+VueoDAXI9ZVhE2i6C
r03+K1lEFvBlvVktt/pR2F0D9KC1Rwe03l3ejWmjrlRTHNENpdY+e3Ild0LZSxCR
ZsRW9CYxiMMDYLfTeNx7wddx9QKkbxcTvjHCQGOMFw+//fbQiX/x3H8T6zmZww/T
fFSMNIWTkHeWxIFBuht3gy2iNHp0a1WCYaQf1kZff3I7kc5GXKMqphPgIRdyTvvA
n2WnlvZsV+L6snO5S7xNfj7t0mMAeXs2jJ3pVerb9TrUlu20wUsvzt5gaWfpW3ml
amdbTIrrvKEQg3kWZRzBjHYF89enMHMjut5iv0IT+zL3vaHG6ldx7p+yUNXbGg0/
dzbc4Rb9LSDTJ6EMZr+QMVMvNpJtwnSzWeUUvqtVhR9zUjgk+FJ1mqtSqDUOUa99
BlyiFf7GigvmaO32VBG8xVkIe1NfAvMsvzTQjc8x9lJWEZ9Amm8BwWltu1Lynfkn
bGmcZZU/hRGh1QH4DdTesfwNkBRtIKKuljVmmTMS/T8FvXnqiMqChv+53QkxkxaF
YxzbtY21sMhzogrsn8O/qbEA9+Um+QCrdpv2AzmT9Ok0wTqdf2vq7cZeg7ifD9Cc
cJyfxTIS0yVg/ailNEVhhU7bRWsEGITdodtRaNp2rs06pm4yj/A6zpwmF3DTlXWD
r7DawTog58QaZ5jSC+cqisrqY02161XNCxSROSOMnhvPBlxisLi83foD588Xg86I
CjcERQMXmbKWUnMSRSLzgWuEZEta2YlMR1cea3+JOheHJB7kz0t96gt0M19FScg2
aO5nLsgowKkqocZv8vJP6HybNwEWJ/MELtm5S2u3VfA=
`protect END_PROTECTED
