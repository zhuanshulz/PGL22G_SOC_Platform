`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2F+06YTg6CxyTRePtmIW9m2gbfMnf6XBePlEQzza7PIuY5ypVHfKBp4MZqHRuJ9
UX6oK0RP8tJKbReRFMe6FE507BfWvF0ZxkeY8kampkpFZDwDsYeSMTqmIdDYtfud
COhYP8hhH+GqQRb7OLeBYdZI2NpkEgqlBpl3PbY5IpFXwrbv/MvGpBHl2qzB7H7H
C5ZrBlYiU7dkSv8FI2oT0khqmTpjwY0jXTyjsN4Q1FN0798XwX+RsyRw5tY6hwoZ
MQyO4Fhe8H98E0Auu1xWC8Gig4U52fFtt1utkcZDHnACbP9B/q/4M2C+W7pLIXXt
N6Mc3yge7MuHbq/jBFkawpnclpdh+SHIFOO8ja7z+0fXKjbzOjqSt0icjvxQBEx3
SiIh+dvAJnEg8CrvbT/IAnRKXtu6yKgDo/ibKb+NT/wqX6jzDB9Wnc2TnFXP9IWJ
uwmEjLiXcznb9h16IF9eSSISPZSiuWQ1bSHUEtCQDAF5k1lQHwZ8b/Nm67CCU0iv
hbk/ivhKXervguisbaqyArKF8heiLCZ5kMTxG+Ryl5utKFg2gVfunHj4LToUshrl
gv5SLKlkDa0Ezcs40rm8TJvKhk8ydYwlywQm1OEIGRMI1Lp/vztNnqyLokPhr2Ej
obx46jfpGcMeD2mwn96/mGZdTpH8T0SF8Yh/5UFPLfnksx6WSBlDdkaaSKWivJUY
iIi+I2Fu3jfrhPGH9AGgG0EU5DAFM7hCWfTKWIRiF3c4zWriegw9pBL9tq5ubMYE
d/Yzlk+6w56rAaerHFsg0dX8KOAByGH+e7Y8zgPDPPB/2IUATtI9cAb7sRRAbU1t
m1C7bmUQeIcv01t3veOxs1hFHjbsrOZjikYKkENBYTEArx7PO9Z/MuHrnE0mvHHF
EsTCll9g6mOXHzm4VDk9SsWKf7LP242o/rdqqRmsRc4k8X2rC7YF+YyQCh278yT2
6HVFirv1WL9pIUeX3qvlO2iZ5DedbFvfVuy4bY+KNv/pMEi/CYOBRYyccEYMOdwD
vsO/kw13AFLMMC/xHGmMr1m7tq22tC5O1hzhhCHAcpc6fMkd37LmQwzDtBcmNqYm
sBpDnbJ6q85FnMGurWmMu9ZIY40EOBp37r19cjabmqGo6vwMbT9RRkPnVDNeb2t4
CcuFDaupDs2vOPjNpamDeDZ3EOlU6wE4R5PlK9cz3RAYmPijEBD2vMiObGx+4TPE
lycCMx4aRUDoPQP0Xvf67KIBIl+6zjgo46i/leXsgyOMeopxii8ZEmbAJElUSn/q
eV9/2KeVsd3LaaJHvMcvIZksDE0WXAcQJKRNX4S7Uzh5/Q08NeurRD9Y9vu98JeU
9VqQBS3yTtw3doIrYfCMqLCCrvRd5/TjqdXyc8yXpT0Xdc03ZX/wkDWsmeFgUzBd
XPDWw+9qQeX12uy//2TIXjXw1svig8i3Q1U4WNuHynAA+RDZYvquoWqcfQugiUTb
EPZQSqfhS52dLgp4aHu1Y9CwsbHW5sc8uIIhGfKDmdueeTeKunbO3JPHBNXNt62T
lnavAammfLH7b1cHc45AuAwsUTOvJmTMto2WKdEn0Z475ZQhiuFtYsyPJXuZpCGr
q5olJmEJmvKJx3qDgkKcJPSgd/KvmqYAlEdpp0Ron5SdRnRp2C9bqcTL7+vp2xfP
6OhV6YKYJ7b1ZOZwOC6noHHDX7uMSjJVtPM1AxTEULg=
`protect END_PROTECTED
