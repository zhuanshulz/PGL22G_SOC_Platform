`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfVC2g4g8k6kFM6Cn8LSUdaoCZGM8gOqSFENnzmf8n/7tHCTikCEGcR7+dc7eXsZ
3ZswrsYbhRJwpk7umjIiBP2wKEG19a085I/B4y16kkYMzkeGkEQUsvNObEkDV9ZZ
xLFs0Nitl9dK0H1D8KYKaSVkr5oGlVnpnpnux04H+iGfBOhmNsrBFyPewFpRVVRo
N5HGsH8DthpmFugTj4XlFuZaaefBCGIrAkXAFzPEPIMS8b8w63mjFcuZiFgaEDZT
/9LfJvsndHUO4Q3kFeHI5VxX5rdsF7HMBmO1Yugv5XTjZJJDqO54Ebw27qLo37JM
TjHmM/C8XWmIQx5IbZCRJSFh63bTvtw3nPb4g6aeL/vvCX9Tmp33spxYldTPHuoV
rVA6Mq/nhIeX7ElW2AzoTN2qTk1fGE2Eq9B9CLPJawV9ihj4iCEw37IvrMxeZpB4
xxxRzNFqIS5U/LQpEDz8laUTxNQxCp0erhyM0Kf3DGKLbY3RjO0UsrhEwQAy6hWj
hmjL9tlgR3D0UV01BQWIIlxWnQCqU7dKbul9/dM8nyUjc6ObcJ+1/e3DKu0nbqHG
5buIJwuovcW9jobQDEPSPA==
`protect END_PROTECTED
