`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wXMXFL/5kBmkolEyTcUPq6ATngrzkRDbrI4xq+gOH/tfJ6HJYEYBSS6BJG+LGKHy
o97HtySxPG8KuVxpseSnjp4QM+/dvtF6QB+8wk6ecaQ9RWXBrMrX8awaQ2nu+iqJ
0mKPEom37R+ErJrrfriSwdNxkkFy5LDGZ7TLYMH2/LNbhBJrmYel66jv9vk+CA5w
hJ/YVlO2tVUtOregrEgf266bD8UZp2siosalatMozCjaa9HzAf7F8xconnI3t3Zy
xhSEUSlSaMEb+GbIvvVuUsiVT8DW4qmoED8aQnXlVZZfGGKmc0HPBbLKhiDWyP1M
WBoqk8mu0kwW7OtzmP2AErMIoDri3LcXPHn0pDC4sOMvFZ21NXNfgLxqbrhE4yoa
jVXIE/ieqWD60TtuMBnauEhBnFrqkRAfBeJDJrD0r95ELlT7J+6yFS8U51vPPjME
7NHaQSVxYREgec/0fkIAbuSppBpnHUV7vERqg5V4j773URcXce9PrCHnsiJVxGUh
P7nFZSnV/ta78GWbvHLuzmaoBdZ2g5PUtCg2FX8Qvr05DpBFsEgMNXx4PHxunP2L
7hsXgyyXUQVcOLzqNNK01QV8H5CumnKX19mzcv0TqNnKjBHVwtlUZq4PymBOZvVY
sG3MIaTa5LtjlGRIotehAGto7BszW0+8IKF3L+z9VJCQ66I7go00HkYmpBzCNLA9
CBbqhTYqa3gZq3VbKo4Z3NnC3FsLPNmDxe99y42ogOAEEG6yDNcqOUg865Ub6/Aw
uAiSGULhvzVrnTaTEDbFbz+HT/yIJjdEoNjbIeU1SqpC3iZ0yQuJRB0EsC0s+Nm3
5pzYOEpWBXkCUlJuRrATUgql0oYB+6GNHj6shX0s+7vGCHf4bbxGxjiQqpmVYEWy
1gIsmZaiM+kowOeN2Ob1jvDl7XZO4YF+g1qGDS050gZ6Eg7wEBBdvuus3uLzHWJV
f6898L20e03idImezhNu2/zP6t0PzsrY+C499kHulxJFWEDsxvrcjGwpd6NPxyGg
SFtiHh7f5F6AUwsJF+9zlzX1LTLWEpGWo5UCGdZzviKoa0Q5cEaoPuqzkF+CaeEG
rRpo69z4v7stqRPrkorNinoQQd/ME2LK37Ahx0Z4DQBgICbIdk6XyHdRrKAT+bNt
26W8nDVOhJND7DQuLIlHQF8JCXSzk3Y+lYHdALW4DjquVC6x/rCQe2ibHSsZdPav
HNomnlHhZMvHPhtdXenETjgOLahT7QCEDMGxs5IIGw9AKCv0Lqh5g7pTw5X1zZXD
unrkIOGzFNAs+F14qwSPaQZHjWO6PP39v8fwXDyJGNfycWeZs7zC4dRMyxDznJUL
w5hUCLGDemBNpk1noayd2rlFn9sUsP9RpqRmjcY/JXXbNiDvzD/b2SG250i4bp7+
z9siRi9c72+fWMlc6JxlmOk5wiTsBL9A5EYSwH7fJhHUNi4IUhOVL1KVNMtaISSZ
0XYGuW3oA8XAwe+PlPI5GdU4L0gytWYEoz5u0Zjte6LAt41UpnYQTl4o54FJtR/s
jdznd0ZddCdkMVgOOr65ZMlNwqUMAEL0ogWh0MVpRw3BXFzWJgLFa5Vp8zVrSOUB
TIS5X/3ROkuXoQWbamm7dKChSCvsOZ6Nhu3xC+rLtQUVE2QjWWY2S8Id98EFs5ss
M5rTuF0erdGpEpx9t2FBE+pJCQRy/jiLKGmZuvUQxxbkez529UBD4qoJ7QWeE1RG
kjXF3oNS59n2PJuL/NUk815hSQWfha6EZQ9jThqGMR8uB/2hAfYq0OJUKCjZWb42
U9aK4gjGRz9czuD05y5hZ60WSXu+yBelCX0jWbf8cc9bf81HsDuvgcsHx8ejhIKP
yXsXxbYIcIGXIibljnim/33GyPJy91D216KYLDChJAuZ4Sz8/DWXlwIEYyR43XDE
rWyMdjbw3eERFQnC7qmW4z6LT6cVpzP7DI3jwCp1DE0pl2iTGzSiAKxA0Q5LLRsP
eKmCv6jzz3h0qw/OWtI8ZiVN6BMy3lxdbk2mG+CXzf0BoBkhzShETK3uPYP6K7Lw
0R34LEz/V7YUkuqG+K9ezGXHe27+HRa896x7xaY++z/XfsGftuT2jGZDZhJrok1w
bX7Yk4nsiwCDdzbbfZGB3hKbes6sdD/TLJo1/oraDuwq5HZGaon+1kzErjq3Km/L
JChNfzwErXBrSRskagRvFj0wJ6k8daMd9DsRW6haggG2ihLZmPk/2ChX7eM9bQz9
pVbQqRyf0pJdG0zO5k7+WS32Z7H3VD1UFXKj+KLOjZAVvZJuxbyngWoNMdd36F0S
Wxt9aJGf+kiGhPmNl302ILAonwI93p6zEB7MhF4e5vGZp3Dfl38fnlfs0KDu2jxk
YjaTH+aunYURKJntrpeRJIU+Ak4CHlWwIvM6h4MihDR5Iw+FenobviQ7UMNoHdc9
zZ3hO2ZxMXsyJY5pO1Zs9GDJXGX3ZX5pbve6FikeWNN+cHZh/KT4ga96kHwXCiQA
Q9c5MmClvc7Ggnsy1bxJLJVEIwstC36Z+3oJXyoLZptxwfTOaCuashj1ONh6FD5g
dSjvygnGncXmT/6nBStsxPduqrG/QduPxOS6MmoIDJwRbqBrKgcl+YB12ZBbZq5c
WooNsoK6CnnTfCmUIUCqPb0yF3ygFl3IBFOi6VdAyxZTqUxFeoSxCjFMxXp0gbnP
zAHO45buCVo4KhII3hxU+raeMCB0+yh/geW43jZaq7BXRKDfO4Ti5J5OYctk3N4B
rIOXqETmqjsFxwFpUnS82ULZIfia2ol8TYfhXkqDrl6hGkVgB++koEc02OnbSCeb
EgnKdqrWfpiSbF5tbD6Q5JVN2VS+O70PNowGPs8h/mM3Z3bu4pX68oCZ9W847MPM
MxqPuRxbystuZHgVSkL1UrLvW5HIvVH1eYzM9U1fMU0rQ9Y7bq7dp8ap8d5UR2dn
VMQqi9tSZEUAqbVShpNO4c6lKEuFkAuZfddptb7Jlo8XCvqfego+NdcczUNyR2Ta
1uQfhnjlPrVvDso5aUJY3XEFjnuoViVAwpsV9ibEAGIq0N3+Gshn0kNF4r2LH0i7
sidk2Q1jFfPn/9x/MlNZSa0EI//d+/Y5vOFjSVi+GOu/3sdeyphaNWZTP/069Z3/
sB0afC7LSw5JboTj7O/0YFkftIhJEZxMSQ2l28zKGzDgjVIsumK8PTczd8AlNd0p
Jldn6jy/WpxpdoBgTCgMp2xyHmlhrcDNH9a7myWf/tXZ+jfm66XCb5H2HDN3hcpV
bzutBO3hJHFWg3N7G/1P8ArrNARmqTbdl/a9ZxxpjSa7fKe3YjcJ3s2a00B3V7F8
smyZyAWdDhGXEzDIP+n0WcSBdZ2WJgBtFoKGm6H+TSZqa0GmEjpehMLtnhQdKRHr
xGb3L/IMJ5mEmIslkKYGxd3RXD41UIpUJMitbtN6UCikNoPcfTLA51/KFT/u5e5K
EClEN2TAl0iNf2fTz1MEK5VsaxdpsB+D8qjtBF0z9+cA+cKDX7F2Y12VCtEn2TjO
Y4nkf1nogTF2UvuyrFz+ozgoy/3aQJUzrMZoxVY0Ql8Cnn0DCRUeYLzzLjJNwOMC
ciJD46KCkNj7TCocrV4Yci1dZSeFiDgFNoFwWCZFFR6XJSmXJ5TiQnQenrIAFWXM
h9fOeN9qmzuiMQenO97hQQ==
`protect END_PROTECTED
