`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIt1r4f8qk93qrCmPojRGPGAz6TRq/qjJj71e9pRNJWZqRFsMEN2VIOMGyQXIZQG
17VpwHVgGY/u6Q6kjLlDRyOzTrCoLkaIYAuzR6iACYe5gWfeiUBdgmjNLiywXDK9
aYOhRTZAofiGughEghuHpo/OqD1h145dfxZ5g9oGFO7AHUbXSUNPTYtK96ZMEQxo
pYz3to7BH8xUL64qYpb5kjiF4CTA6BPZq6Qq2HDBSGZ31mblCQMvgSf6F6v4ycpC
GieqqbNqfNVRNmSdkfqldw==
`protect END_PROTECTED
