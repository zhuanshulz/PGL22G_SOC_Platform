`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwQig/JqVpawdtiUjyS+oPDNZFxY1kr1Jj6+8Z6EYSxHTuEaW4MSjLVmn041O7qi
iZiOQqFdTi+XSbCWtU9pNwsVGDKao+ehdtAzkOLwH/Ma05OwCxv/LAhiXIsU3z4v
Q+QhMfPIOHg+fGFkW7Tb7Z0p9JBg0t3muF5LTy97lB6D4lIsVGHf3OPlJr+PqJCo
pw8DQoV5MXqhMKcUiQ7BKiiqwqgD9pD7U32x4RQL3SIEo73OP4ZpN3vhNq2jtsSR
uJ4V8MUUxleld1zrK7l6bTv27XAa2i7ZdSPJbSDZ7ge1OELdeMH42B6qGs/c7PnG
OfmCL5la77g7XLb5CUVW+90TYvl96xa9yiWvpbJ0JDpm/8NQZz3JzLR6aO1tJByy
Hm/JBKcOXsBA5cNeZAB8bXeVjrt1ReNaIQYOy8Atwg7prBON8dw/LNwIxy2DPouY
`protect END_PROTECTED
