`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rs28n7RQYp7Ij1qsVMHJbFDzFtfKKFvAGOqQDGSIs6KNnUxHAXdL91vpkCvAN0v3
pi7xcGSfIP7FYK7Hm2J8h2HpCXYB56fGLtzE/Sk5TrH96+u5rNcv0z5+N3pCnDgO
zEjreB/4bwzrSK80KGAldzWrXMBV6wCwcBHPWhYolYT2SBIGamediGGrbPkrVU4O
7X8Pvlii/5Qcfe3Y9EUuVAXGbyU9a9du3KoTMCvakr/7afEpTKMnBynBJaenF5/q
y0eRXeEWEL/i2SpFO0/4FFuF6AEkQ+mAOsUfAPk+6zOSoBda/vOvcyEzCoUgnFGP
T6VwBaHirruVujAgQPI1LI+d+H08q5rhNvzdqsCdNA7UDzVSYzsXIvGzJZ+KVuUb
OydYjArHarZqnRVcwXTGYidY4o4r8mQbaN4w9la3TEyp2x/eEczGm/I7qC9VNUgb
X7YWh227M2VSskXQyQCHadRXqqjKvK50WmgcI4NVgvY+NR/N+WCE0TBTm804Wpox
sOCWiW4eL4e+qz1eib9EHQ==
`protect END_PROTECTED
