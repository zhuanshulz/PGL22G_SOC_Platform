`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xK3ju8Pw09OmQ5AorQwTKDknRJ7IwMP6vKG/E5iq5AWqx0ky6IhiGM3IBG9aATkO
dhv0aI7+oojmkSwCH0NNtEkQTvz0/msIF9WQmegOkrBWxvI4k8HdRETUGxKaJtsw
kOKiUzhyUl/WhxeGXPcLhpIZA9Lpm2oDnLLqpvMsUzvgFVyFrITs5FETHeUpCJNh
9kJhcO3y12OqcpR3At2Xfw1SakJ9LJF2gknOzggqxQcYAWHISn/592o7pxgDO9kd
sGV2nLdkQhI4d4BAJzfhvanrp/st5z+tubICWyYOK4U7byMKRN3+tSlIlG0pJ7GT
zZNK0Ugd7REx7mMP3QVflAbqTmu4svb2Qj9PeClAfoC+KuGBzTT9vy94xfPEh29e
wFYPonkXx9/CbJzgZuSmUhOYVo/+LxDPIxEUB6+D7yM=
`protect END_PROTECTED
