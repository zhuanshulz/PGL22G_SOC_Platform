`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
diEXQlQ0Rb1V4WpVVnV/D3R7iV5IMhiyWL6tBtlJnpBGAGHN3bdnIQAGMeyKYo8y
bwLVknTqOKqH3dmMeK07d1JZcu8aLJxrO2pUJwsDfcVohKOLUgQTb+6CbceDFmav
Bh4U0fcIEVOeb5yeecGTS8fb+/LfRCbqllGzc5CISAqTERxBfHFq0rtYcxEXv3cD
oldoSnlDQkjhljAzZ1RWt9sSA728UFngVeeuGOUflxNBcwYKvhwY3wgcgcq3ACD8
s4uhNQpnmYeubGPpEJiHG2Pm/XwfnxcU06uq3DB/hY/EPvbyCuKXVIhy+Lnvav1P
ZUsC4x0ZqXZQm9eNnfDJ3dweXkGRpPy59jqi9Z1fDT8Sbqmk1MzHqZvNr5i6pxQ+
XklgZp+nUyoh3Z5lft0V7D+t3BIpz4iwu8RK9fVa0ydzNKZvUmYfVW389tKU/nRT
m/PPcbKuoMImGLnrzHFGUyHjDAouDcvqH7D8TdB4AMc6uiAQyD9KeLRP+FHwlyPz
r9WM2qZ/AciKOS7NMTz5IeuTT6oZnSBG32T3ZJqI17undh5gcgV260Zygid9Q9/p
ucUFsxxezqgrchs3tghHtxP1pqq2Gc5cClFeq2T++GRmL0zJZDWCtbJLh2RoScmb
2KShYjl/QMzaFKWJ4tssIJ4EB/zAOKBoRfj/9a7sMqxckGc/xmRs7vIzjfMgrLgm
pZsT9gg71wMdku9vuvuLqP96UT1Exbc7zbRSZ4cUMwrwCTw4cfLEJzdqzhw/5LVo
TwLkcyHbzvfkp49nFVm5mwtPEsBzyvc1dDBKKUAT2jdZR/FwlVchgqyGUZwPMotc
fWrjtrzE+Ezvwcdf1U3cSJlZ2+RXRR+LHvQv1OYPifPYZRIKhgx2ezYpHAZW4V83
t6jnYRHUWwxaM+d3nhlIFAAUOIbOd64uyFNf7uGHQJ5IdUTu6Y1vibi7HPYex11q
iuLq4c0H95l72EbJKx2JV4BdU4Wb3jafOlgotk2igVkXZlSu6hI4ljFUTsADbPT5
PSn7Qk2OiorFPp0KPEZ75qHIcDGki1wDsIoZ/6Keim8Bh03dm3BanAfnKw0sdyCI
o0+/FXQXUZltO1D44Ht6YilcWPuG7TbiirljXAdEhY69M9g99Juc0lYHk+UrNEez
a4ESyQ/6Y0yFdVAB+nma0S4wiS9saSyoH+guik5geZ7SLeWpz9v2wDQbtaOvy2eT
QzBs3gqbIh76KYLHEkQ+SMnvBuPAOaMurvAGZHtU13Zt3sJMyZ9+iCZfehh2gDLQ
bbAzOZGuPMbGY3AiJTjnrMbq7HElqLB/vZsA6wXokoTc0zjs5Rkk+6n0xJVepAmr
+41nIKc/QnpdoGriz2cj4WoZoF55jREAcuw63EplmQ/qlNdvUHutfl6dBFwb46U5
8peGEQzuWslGYq+YV0EhaIexAUpM5rM/WR92vG1GujkmQboipAO/fU/HcnGGgtRL
CbS70A3ZmZTZ5CgCC1LxL24iMfzw5FAtehLWH7A4vgRDPKsLaTS8LAGl3YMsutcL
B5v77701or5ErUAQtcCwthjpvW69yAn+BPT1yDBPMJQfWc4UJGqrlHkoibxoc39h
lW4cXcGB4ZVl2g5/2s6Vu48uzFP/VG8VOOx2jJPubWTWlzIEQCWteEP10qUWWbG3
mkcIMCs/Hm0aMstAvhcUGFL3/5ur/vrXnEndkVTisPEB4ZRFOLwK9+D8EQe4wSfg
XROpytKvuvMj+40NGt3cXd0i5sU3A3+Cwxo5yXXm6IdE40pJ0SEeuTzGPr/MfIz9
/4bvuz5Im402sI+M2sZdTGHyHuGDHlf0rFoUlxkGCTuQJCEVAKiaXF7Z0cK6+337
QDfB2j5a/AFP2fd/1ue+zRoMZkNiJv3P/q9z8YV/umy5MrLypCDaZd+8LBxHo9z/
gJECJ5hZYirMv0qoO8eCv8ods7NVlOya3xgtNi5GiQiCbEuOnSR7WtEUkCXeBBoG
vPwPQHnKHhKljSYZKWzFwx1jX+qhcJVVGZJMxPXXmqTEBNqvv+FG4oPSdmpXJsr2
NOokB1U+zT8UTC0cGBqVDHSYjF+NPJiLE+qfNm1ZWA8Si6eid4FL+Rnl5SKHTi2o
auIOHA6EtSAa7bUCfVYFV5aM3Co/AjD96XeC1/K6ASrTUt3uVOFRHd+FcJf9IGOX
gNjZ0BLM/EGK7MEkk7tSw3ikB/6vSe6OwpyMESzmID1mkF3ATYm241dRFlfPutQG
nTfNbHWFpW4Z1DiPYE56hV4VYrr+gGoTPGM3pBUmzvMnbgPZK2e7yRxK482QUELa
DoOjBKT/dnEyMEOeK75xPNrQ7+vH/rkdyP/5pGoJ7abL2fi7R9ZQDHR64tNPhvLY
ydkhLVDCvx65ki8l3FqzwTkU5q3Vd79fQK344bPpRiXg0iGuhEa8VgckOPKykx8x
HMoIfoTWhk9viJ7FhRES6FAzMqr/uLllbBi0MVmJaOucH5QZLpPqkYmL9JXZCjOI
IeQ2ZaaJjy7whec0wpHC8Sq9628xAv/GRdXW+wWWzYdjOG2n/dybBsIdD5CSmTyg
k852FkmT3C3RhA97hUUCljJ0sMuRXHxTGEJJifuMCMKf1dRZ3ikLaV2A5/q4Pyo4
1W8STMP0yF0uEOoIWKKdZUPaIe+r0u3ZVd0/KIOKDYaJNWpYWxcIfIY1WdvvJ11S
rbLMWQMo0E50UMNDi8DRmu42Oy2cawWY/fco62RVm9pd3vLhXDaTYkBImrTqCV7P
1Fy1wti67IP9ldOYZ5xpmw2VEynkOVC1a/67kc/Df/XcMUsFGu1Z07CPFLybZYh3
zeIPFXWnW3sW2dpMoMrJ271aHdlWj9RST5Ppra/YkQmxnFLz+4UtfuG67TqKH22e
FhNe9DCMbkG4L53NEZgsd0llIPwB0rKdNLqHXf/lCNga24tQs3x5u3GLtybb1it+
bjg5l2BkjZ0nt0aQEjcdjn+wIqmsJACP4h7n+wMoCH8soUD0nsXlw1MBVvWB5/3a
Ld8BZqZoCSSJdtzS1ydLjXn8v9WNFAe68NMCknRmnUJrE3MMpHNHwbzHFyGKtRPn
lWf+vZubXuP8lUSR/bl2oSNVa0axtO/mdu/e4zaIR37JpKXK5qUl4Ks7XO0wPUGq
P1ej7Np6+NBElFmmtpbkDfvGRCUj7mxBaq8Db3T0LZcrZzYbwo/lDYvpznww8TMk
qn6B32qivpjixKcd5c9VdDJ4fSZwpzZxvvsNwP9cYZR9aKPnC+BPqjuNU76VKekf
VHj9F8ZpPdyQfy9+8yX6EdCVJseEhf2dQAnIJ5CpjCzRk11K4QPYiPCEv1rcsbIJ
PkgVWhwuTsR7HsBQMuUfs147fAkN92zRAqjJjIwRPcDP/2G7MO6EYz9QU03e64Nb
7V0qep4uBGGsPmPrUQwQDjXBEfv1sIQVUkVWywxeWdflaWBjpd6Ja2mn6AHrK6HX
aziOrujFgIiLCQDvrU8GyaoFRAuqn7LTZHKyGpUKAkkkaLnDJDwTMJFycbbvKB6S
MUySd8E6OdRnN0s6pwzsjgCkwc1FlQHD4d32iKdT37CyguPwJ2k1tSgsr6biEiRR
2vys5QksBfK05MmBIu/bXLIKCNll+3PMFRw8y7f9ldvMAFDxppkHOM2VF3wl9bNc
Js/+RXGs04TukQtWy1T6MykS78KXnbi5I2Z4+j7fGfJEdKMoK/Aol03LIodF/B87
M5M0KzmAOZc54jqlOawRbPtNiinJV1lp+3HAPVtae6/Rk1UdRsktDfUI2W5lNn9h
GxamJ09hYz1p3L7Uw+7a+892jaAOuH2C8M2n4ngQ6gGRRrQqiHjobGfRW/+m88BB
pMRjMAF7CoiXpoRZAoyy2FvA34lqoXgBk+XvN4/w3QQJoePdj8+C4p9f3L9vK2x0
HldrMG93wBs/4ACzUybimo6BeY32526+lSdZArR5EMUeVTR8C9acFplFavh5BGPu
zb61cjuHm7aqLv6CA3z+xnzn4SoXa2C3K8JaZF4i4ickd5FQByG5NHKzmzWt7GKx
6WikTWHMB7vjRshgM8k+HJOmJcTHeXfvu0eVkJqtByEB0tSEhG3eFLMImI/asZgP
D2zAd0nx2puifKe9nILPqI//BPne3dJ4GDpT4vv2+8fy8UugOhBouCs+dum3xwhA
QOJyTuzhjPK5Nk+1826G8CP0iIx5nln/S7sVbQ8CBgSDh1qkP5iSxFJ/vg5W7zuW
S6IqzmKitP9W1xiqTh+AuL6vn4S4o1e9XBbDkLgfDNEHKYMOJ+0RIdAmm7HROQAJ
n8D5Y+9OU6xz4f911qc8wI1uTi4yaPrARdkisR4Fq7diaI/xFWOPptM7X+z517ZO
7GzPpSeVgsdeQWaNZtVE0IatBaETU3NY0UfxI95RVsmtY1jzQGSLzHSIcDx1UVUB
ATYPQa4A2qBkuc9Gi5PAAMb7RQUSlSYBfURfG875+faEQW9de/9I2BPRJhTVO+8i
q2qe4YQUuuSLPkEfbfxsYSnkz9GneJ26SDeOUOYlS/xBQea4o992+haNXwkl9kz0
ltbr8UETZktQm9rsRLKDzM66nmjDLJ0e1ilSMBHM4CnVSE+n0W9+tXjCAf/wLZs+
QC6gQ+m5vz35F5Ndp7EFJo7B6LmMdM5YV0xRnCF+cJZo7RPUdxry8mIgo1EQ79Nd
bhFIHEwh+XYY+DpCWYobCdL4F5+mC4IjrVU0RUf/0Zxd+ApvUktShypj+/qUyF63
2PeY6cNS6t3pKSsIiovkiwlP0v3AtUXEm5mv3iqqka0=
`protect END_PROTECTED
