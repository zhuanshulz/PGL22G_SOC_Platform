`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lYBh9MaEVNmfJDG3SjJmnBrpt+PfCozT+rPwiofSR0mAL4n5Qen+MhkTvEFbRZch
PqFcrrQPe9q5h3GrmDPWH57KyiauUrp/YnMXIjP3xRNgWf2HpO3M8AKqSgayPoFL
xcnpoRsAuHpuqBwGKCiSxJ/qaT/xtrVcBt6f0/QSfbJ9T1WZhPJtDYWffLOLlJnK
vmSZSfpNrNV+SV86Kx57BIzuVKAj4C1AmWCymwCLF+Xo+6GA8RpYmRZ4eSpje8rf
9baBqVb5AN1Yv7TOkNhdDa4KoqshwP/NxhjUSfWYxaKW1+kB2G08jz1huJmJjmQr
sjyq6hN1UKqkAw6bL3yp+r03BWlk3tQq7Ov//yBMy2KBAIq0TkFl4K/oLLYPEthu
egdFDl7Az53He0IMHoFU9By0k0VcbcSy5sEoimnmZ42WN30IjqhOQgw+QIWS+Uf/
V49X30P3p0pr5d17NWCdZA==
`protect END_PROTECTED
