`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Vm/4DaZs3+HBwnI97SieWXE0f+hjwwSRry5k7Zr61wwYU3I6xZrpyoj6K72HEnT
KmEgKi6tsHBJNU6XXSTgaw56F859pUyAFpN42VO59vi5scrI0wGgoWToD+B89zbg
1ecm3lRmI5VfwnN0MexY65oc99Gmzh/JARSfN5Xe6vQL/XCAd9zqzfMa8BNWC4Tb
0bvAWEOFxF+NPosBpI0J8lY/wSt2Hs0jqsxOVD48NyUmI/thnjYAYYF4ohE6djFZ
aUDyeytFx3EB96qwuLs+Pgkq4HI+r6Cj4CIyGzoVjfVoyhGkrKNw6f9ShwO/PLzt
oss7RzxXbqX/hRSS6o5vsfHBkQR7YyKMXqonOlF3cOOZvnRzSmdJvhBRY1erOU/0
KkDJ/xNtmyUfvmzEjebkxZa1NBerNbjOkpZ+lreLvd9vI2BvOgL7y2e9N21VfjUl
/kfv6tvfVJ8god3/iiZELC3nCaC4PdMcN3ZhkQIbg11vWFsALQ1aeIXo6YxLInHC
rwGOjxnVU0p068Rr0iNAc9FzY/SjNXXHpcUH0JBf5YU=
`protect END_PROTECTED
