`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Xa9MkOzzMdnjMPwT9Guj85qaUwDNxy5iOOV0GgQH/pBJ4LiWxkvp7IVN8QT68Nt
+iCPL7vzKdWV1XEiaLet+Nn+EOuyWqKex5xLID6EvvFmfFyn2PcpGKGWDDjfHlhH
L/ndrM+Sb3wV5y4YHPklK072zRrOEUsD0QFIzsMbNFdToaU3IWKc628OrQz9030r
7CK3Wuja3XiMTbt4xO92rFNcPj3MehPRI4cyiTXmT5MjCL64gsyQB9A8uvrmPkIM
jBaKGamtHwGFTY4AlBo2zv/vCx4wDNXgyZzpZN3MLdbjVxte8EGNFpFf12/FHLqK
n1iKPUqTtlVgmT5nQHz/RDfLALWAS0eXrNKMD492a831h1Q1n0oij0Fg1iXtKu6p
ii6cgqcX3mnIRiqi65WmvClDAoNFD2WTamjtBwAujFFBbLlmlM8Csr9Y8wBcvpyP
3dY0bnaZ8AvLNFxgiSjUnmva5l0FHl2iNecb4pbMw8FP+P8g8IprHA9jmCnRKa8w
x/zBvBsiSXwBdn8MKaZJ3rtisUgzYH+BTDo3RNSHjwsiNcPevHKjhVHdD5DUpckU
wSxYiTDM3MgRxF3ltQnKpwxi4/vf5YLAduRfaxWFxul7SOhnWYov6vKWW9gGIUnK
zYTat4ziKjOrbWAwm+m1Jz7TisDoZPqP6OU6i2IJdLu97O5s9+DckrNcduTQ1Iy4
mAXZaFnZpWaGmlZEFN6aaZkQTyM0y/LeY1uHMxeGz1VwvlY/ZR6roWGROiPPrJs6
pI4AbKflN/K2gkcm1LIkilbNAT8jaIuH293lUx1iTrNupQP3WW8EZ808Xm0CjugH
dAQsCY4BmVxFvAz7TrlRmv5uDCK0kogy7lii7QVSsvRH3HAHlwoZo+J+wGgQs8q0
oqyO/QCttdeLNyyjbHSiWOqjQ8lbaHbzGHGTqxqWWQNtVADLFPfSmrR2I8OQXucL
U7BiGKoDXjJTpa15iLMgLCeoFsnOFmquf+LP2i3/UsJEgI4cxuWXZ+gznsik1OfY
wwCYbhOE6or9SILlDB3v+IYQZhCx98lHDNZzoeqX4IFOOBsEAzcFeSvoaxSFD92e
taZ6mhDtkFcSWoETL8sVf8Gq9cDKvlbCUlx1V9+KisLNc2h03zgQf/g+wu2vI8re
PuatcApIL81gdcxeEMyC6NJNRViBU/ot/5TaZM631JP8JC8rCh5eR4mLI4oonGCP
9js+BWc5Tcr7y37H8028vDkObiL3yVquUCGLJWWtYecdTP99v64yCLwgyCDp3TBL
MbVpCXeJYtQce8cCtWgYoIVnVMDOpsci50mLMgDnyeJ9C3X5VywgL02pZg7hLp6N
rd7inVMcWIfq4Aze8haTPn0FMfCqusI1S4As+3+xqEEgZotfQo48N2ZCTeas9Xqz
+CIBSEDLDiuGs/5DWbfu8E2GsPbqpZeNiH7unETTrN2wH16teieRf2bvNHam0BDf
9izITaoKP/ivEAC8/GyIHLI9Bx2M7KlFxT+dN2bYRPz5CMdzOBCMcQ8/yh/oLPCj
KizTKojjyBYccyqrtUjHlQiYkawkhOmGEwVHqJGFqCRk24xbzPj13R84htGs1RPB
S7ZQ/NKDyDu5UkOf0kiVkH5nWLTaU1T4FXG5jIzLf+HAi3wSVI0uqLgOX1aE9YJB
Q+p6gyBBmhvo/22ikGfMm8KDAVKckV4RJ1N/iu2GL91ofMnUTx+edlP1mq53nIhx
8dlZF5LupuLee9aaqMmv/wWJR7o+Vo2OGGnmcZLZukMvN4os9dUpZZdtvxh2ghOa
Y4dGpTBsZkcOs+BL9x8BcoG4EnzupcmeHGLGQUU7eXSQO8xL/0IqulphwWLA7uXk
inUYVHn8f3APn4L7/bhL1thCP8UAOZsljlSH7P2U539i/IwlKvMOvAjoo2dUWlfs
T4oQma3ZWQdV7gjVMhVXSNpT9zNDb6tc5543w1igSsDCzUn/VXTBCaSx0nFHU40S
Iu2mMgp5250zzkfjTWTzeC6jWHTD3O8k/OX+9NSjwCYA/ww1RFeeE7sMyWZ+zCdG
y33+02I6p/EsGWVGoJIOmKt/E7Kqkz61Wz2FxRZGDwJgKl2JirZRlRWgtf6OibVI
zI9FiIna8UgkMq1IM3DLOQ==
`protect END_PROTECTED
