`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cb4mIyBiTmTsD/TvJbUAqggYhMTk8kPJVk1nu6wIZ6RK5Kl90DKQx9DNzCXldvyz
8z1IqMy1qHR9RPwM5hl4H8S23o3iK15Cs3D5wCgd5t0xoiFeEml3h2tRlMC5zfTk
kcVvPZ6FX/JgUsxAWxGBSw5UqDs1+5fmLbNW2JanoSZXUkZ0pvzUowtOJ1jwMj2i
7N66lIB5JZ2jNTtj0MqsY3JwzwR7+RYFCIuORX3X/x54dRLvPz9nluS6uaKPQJPz
5vGKe/UrEUvFd/tuiZqB3fHBlJZQjmvi2h3BAZGVRXmyYbKyDLXGT+Yix42EzJ/S
Vr1Zb8CDxNpoEB1p3SS6sl3vkq/kF3ccsIlIzPoa4xdxcDmHQ8Vo9GDb/dpHOMoc
u65J6r24MWSUD6xGL5kXWB92REDBTSPRg1w39UyMdI8Fo38xGe1PJCeF7akxfZUW
74lU/ASDj9nKU3znpEH7b6LSpgL1s6qzK7OWFrUZ+tBS8U6umbAPwoUQuopOtEx1
dvkxy92/R8J6sbNGCd2dV20smvfWHQnF4UBI4QCV8Kk0hUw58/j5UvguM0B0bPXE
Cc4Qbp+7S1kVR3Zbafz8cHcIctQ77n1AwBgmdQv7bOi+uMmO8KzAqN1WXLbE7N6y
4uruGgfnSCA1mRQqiD9FP/zgkz5Dl9GjzH7WyWsLV7XAhp6dEn+a65Z/bO1p97Lh
8Wcm+6/yjIgXDHdj/4OZSTMpXayL565XQ46oWXRGTUbS+MtB8Z67IPSGOlGj9fk7
ORgljhWDg69O9yVPS/STco3DaXX+nbuS4sNgFuc0Mzvr/4r9y8XD2US6I9CJVmoP
wcVpdMT+ZVxoCRJaMB+LQAl4b1cxKGxI1VbmodUHdnhYlSXhXyANol1CnArnM+Hg
h+SDIDGXIetAkom5z/clMt71km9BlsNxfBOyrESS3YUr4FYeN7Xg2AowSyRXdznr
WKiF94u/AU6SWh+d7zrsciE3FO05cMpEG3LAe9X9qQR8qFkwzJ6Lc5nis9S1lvEK
TtTuL53brA5ag+4O9548jRYiFFm3LhNzwib+4P5hX1xtdROQq33lq+/VE4Io0Brb
6g7YRvVjiYPD6f6FDuyUIehsxyadAe8zTOiGtG6RXXAe9EnPys08opet8SFDLRqu
i8mtCotOhnLFzW6HddUFGw+wcnK+u0aeTB5/546+LGBlLyzGT+9f1QbhIp/YlZJD
KeZcC7CrSeA+sk78Lb7YTQ==
`protect END_PROTECTED
