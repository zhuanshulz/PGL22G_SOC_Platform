`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GfuLWe3MXsBSsa5B9FKvLyxxWRA72WaLAkWookfRLHMfxYx275AA75Rtnt9wD62T
1aKKCSoE3EUVJmjVQbQ+NI1R350D5dbXuF3vjViB3U++SaZllMEP6mvLp8wcz9kQ
mpCdZiWiMhOVOy56C9x+sFtgwuwf3WX95MZRAsbxX8QdXMp7fup1qurhozoya+94
4TAFJxZoRtpmRhtNpo64iqtBtlIERfpiCVOjc8zJx/JN6Oz6FCkk9bU3f84aASGA
WSahMmkFbt5ZIbjSviTq0deb5u6kemcAfWljeya/UTb6kwKkYhS01igcyap/WMMJ
QXXtT0j41jF6GODk4+Z7w0F+gnoZZRZnzqpVZyIa5hZUomjv9cYvPQPaMTKvuEKH
GaneCGn32+9vovbTWHrC8SxyCzPjlZM1y3l1GCdODbKJLhkcRo7ghbuu9jyJeJWN
z50MZquZWTq2mZNRoIimTGjrveO0bB1Dt/y4oSQtFRTnePBvjv3fDCBkg6K2mdQU
zeak7wOvFl6WIEwXfh6gpeZhExRLVKG6oH9e/72jc8kZ+ZhtvMOojc8umWn1eN1+
asUHbAFdBIHzPXgtM1qayw==
`protect END_PROTECTED
