`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHe+VbCnInuwOUhhm9FFmp99httvg2lOxP4v6ILS7aZGj9VHHHfiewQw6/jnHoVC
jF+GB3AjddTKkApdgcbInP1OKsqy7Lj2KZKnAfj9twVZHqFO6jB8tdCf+09SYaqP
YwDxOLS9Wj/lZPWSqFrCW3nnAy5jCppO9cehgtUbx4PE46sFGO6BD13h1GevIiIB
Ju1KkkD+QEE7uut7RuKR3oyZLonqvfdGy6MjkGptT6R+rTrgnm9ZTeZ9mk+fLxXw
IPrOcXUenkCPLH04kMyCCZt19jtCUsClkfMeJRHP/6jEHY9iKZ1I57qlrZK0Qn9L
fRXxO86jNksHv6P7MfW3ua76KseoAvAGfSxahCp+P9kNsdYdaD8pzyDNegUxa6gL
EYdOAFq1xZ5ggHJUYDyRRzshmoDjjqBFJ6AfKmqH5E64GqBVqnYCksf/C6FQTWmN
vJ7O5jXEHiJ2UXaGgNzc9OiHP3kpWqO8PmUeh6ndMGyz+ywNVVu/RKSncTDWIVAY
1NnPXHtE0nP18i534szjrs77+aaahUywVfzsvFAn93JpsM8KA56s7Ku0CFP/VgzF
8SO5Iy7SVHjbrejnYWkG4Dt3Vz2MsVcCatMp4d+Narp2HS3fkIO/8f6ztsAusWgD
OKZqYz1M/poNmLUZ/yPkKrfl/T1mIx38I8joS9hEcwje7w2OyZXzBC0ga/gDTmrC
+Z+kk8PKlRBdjl7BOSnMr0NKztqphgydj1jHrY7QLxcp8m5gWBu5TXeVMtoE+Gg2
mb7vmraqlgcSBFK8ncySoUAnWF75J4bIvATjJWJ7l1kL+iPIxoQCqAHqW5QlPS3/
bdqziSsDCurPCNY7MKnveKMv2kSNRs4k13Luyv0Kmq2VlTvB+hzJG8ARGcCve+qA
1rrxrZewl6sm/4boKC14fo2A7+4BuODkN8Ks2+qu1Aj5XsvLVBqTcWc09T0MX32I
`protect END_PROTECTED
