`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mxCurwJcbJOUseRgFZI1/z2wY78pG+HvOJCju58cxXIxQl7+C9oo2W1Ri8QmWH1
cuXJt4Y6zHHJ26VWpybV6qwJs/Vo97Mbmsfxlh8EVkigRiShjw4NUkacrDahXihS
mep445+Fyw7J+T8lH6tkV3ddnpumOSwWsP9PLm5a+fTkeO5epededvGuqlb6Vi5z
2yXsigruUR5/eoU9VADlpF++pdkGtTagNa4MgrBrHgfPNSlYPKrc3Hwltj88chET
bDZ4chYVhCvncAX+SEsnL6qFIdTU54XBF7KtL43M+2Bfk9G8cik4ncoNZlzBS1rW
MlYvtkv86C6ska4CnRzw0xfP1vP1WjTHY0OFo1t1WAkL1StRU5nX0DY4/E/qCa/n
`protect END_PROTECTED
