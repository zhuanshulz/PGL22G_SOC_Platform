`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rEhZlVoBbQxwcomcaYhHh/pfyvKBu7mH+//fDiUeMIJff1liE0mwZiEfFrsbP3wG
s/aWF9gHuas0ecEsqtT99fgK2c8p2I7LzOnqYcxKHA1p/Ib/QF1otGrKB3Ym43l0
b6prvIZAw8rI7QVb5FBoTSo2sKYtyKT6xQjpsbbob+FQMioYBu+Az5EjoHGb5cuN
Y9zDe70Tclbm0kfWZX7RGdO+zPlw53cwkdhOk15HC1bf1fQDHY+yJ/6gDrqTbSm6
96u/Qzxyp5dZHnLjqZ7cBY18d3mEGPwra2sjnwwuONRHO9betCSI9xnHPZRLye0p
iWel3MEmtbA+laYdEpD6Yc14dBCcoEEOKotNS4bMPX87rSchY1qSC6qJKwB6b7o5
F6DQq1r+fv4PdPLrUiuxK2Z6Kf+i5kbHUY1TpK4qkpcQ4KWiJeTi9WDZhkdEeIxT
6TwvqnuTX1vmMe1vzasnad6LVZw8SF8RKMkd259Qpob/F1EPYPxROkQWj+rpg6e9
W1jLTe6V3lmM3LiK36s95+pJyWvuF1v+s/edLzAH6V97+/wEgmQgvdY7LAK+tONY
7tW4BqXWKjYwqI5dcpXZpREKk8XGJLkJGvFRh80+omArqwsBX7EMqwgX2xSIGIqy
/g58WL/ceqO+hBlKrcRXNwbzPBLg3Ih4fUmi36oz4BBpB8yvvTu8GbAM7wV+5MJQ
R7Quo+wIeGqOIwGXrzcmz8kieBmsG/M7OmgnEyDUuyIP3xZoGdR11X2uZc61hDgn
nyRpvqeRpKmy8Rh5pvZNQBoZwpbuA5QZYGukelJjfcYupf3YJgjwnFeHK9hHvIqB
ehRjko5sQ1YznhfXeSArg4xFmYV4GL1L0T56aLOSZge4NHudkkKbwNH6HzBpferc
t0g6BuhbHicVC5/xMPOvlFEA5ckeJITCsBXGSw/7v6c1fdmCc8i3NV4UlRTDY5hT
J8ctkjYfRp2w236fJ6GmDIieXyFStp+tLpOBK/9C6HxaUBuWlKRB3sbLaGlDSoNr
O5LaGfwgVleR2DXTd6mrZICb2YG+pyrbC5F+vLcVsLSDI5GwktoGy7WyTnyI36H+
/c2trLbegFcZtz6WrWoVA6EKeBOxSo2iOKJb5c3wdkk1YqBevZeckQNS8pcoh34i
HCzp+ieFqhjkuBHsivJ/p16lwPdg8Kh8Hp5uTcN79KkfY/Qyq25bsAXxV4pRpA4u
3LwpRCmXyCwaiZGrYr9Mibr5HJvjGLyhSnVK11cIvfx34i7/Zpet21vCRJUSKnzc
tXCJnrs0a+ayTCEIVDD+NvKaIPSWsW+Ut7T/u9SdbAIaUBpOJ7/jwc7DIw5wduQv
0B1ktGNMfGOyOM1j9nhvA21d4/lEEMRC6XefbKCUtigG2+xIiVPtteCRBId9sUrU
TWXZBjfEsmAv/Kp8k2vJ0haHzHW8u6vao4A4ABAChqM4v2ogXRFburIXbZhFeNH9
Vt1fE/UupAEwXHfzuFN2peLv4fAudKH8vktJ4XNgSMzcVx5t6VIAL3KXYVmjNgVs
QxpN1XP3VaajGWJXFAihK2m8mK1oSR9LNP+My7FgSHH5lRwDUZ9N1HzX1rmHoXwk
5GWWULl9W5G792KwEu30rWzGQLOMWv5S52tqP9rzgkuu7XWK7ydP+nMIe675428V
ZaPiCBEB7BqacY606qH/v7HQj7Sv9bGoI5UdTBHCjBAlpIeyDnzj3oExr+/kA/Ib
DTvwmrqeNHQGDESJN3Nctvcvv1g+bWMiAJBwkHUlFI/0sqDMijsXC5eGfCDhJf4z
qkK+hKft6NSq+FnTTALCeUn8wGYGKGwloQ3pAsCrWH5AV2Tu5V7+6MIb3SghOxJQ
1BXoHJS5L7kS08u7iQcCBLTGCImMe56O792cfX38RQvS9O8cb1jWNS4nkO65u/P4
9G26iuOZCGQrmttVEcOWgyWJDz//PQly3tnx+djPku6Ov+JZfufxgRBmLFe2BVqn
QVZaMcZnTZOw7lnM7xr/pRzWM3fbzBw3LcySHuKq+QHglcBuERSXmJLKgxbK4jGv
uV6fjNW1N0kL19FXxP4I7n09lsOP99DlWgwlM0aa7LqXYC9EQaJsSUpR811JPDA0
1mbfyg+6j9dUKVt3znmUaCHbHuxZSp+oviDHAZI3tPtIQhw68ZkqSwVvuyY5FuBk
w3UcBBtXLQFGUWGieFT9TX37WL4yP0aGSirkIzR46M/nKV+CJWYYvLw32bG9lBc7
G+9TPnq4z7ZQbFmc76kDgcEIsffNzk1mvVFPLnrp6Uq1FGNiPI0TLJYRrQtu/iRz
ZMyHa6t/nfclF3dh+amITZEA9/7Wpekj7GMl3bhOx1TibOKG2RTe5gU198Ywv40c
SHTPlHZQiZky3G++1y05syAbnOIq4WbrWKjfeWPafJp7fpZHOXHkyM7yMyT2def0
ehZlhmkpz0oSNgUplwjdqNP+/vUDjIUuPInfB7/51plIWxem0KnutemYJfnhWUux
qvafuntWHwmrWJFaD45g77Cfo/YO4lHKdjcxV2Pk3xmli6PlA4ytcecoOwewXIdO
1Dh7vrcU33KaBI3qyt+dJ22A+HPBEPteZrLuWPzaXKDavWwua92l2LxjRp8p3qIt
FKVjgf81TFF1lRcZ8NB/2ZrKTlSJjOEWknkv627Adod7D3iNEZ6aDIByMHJpmexZ
m3ZMbSCUZ7/Jz1dmpRgO/WFuY6AzgyJlcBbaMnxlBtMVFGiF/H3W9jMdmj6irj6V
SrswWkyIYq/4pwyMhq4xuYiS62iFaLIDh2ir+LKdlqLciCUZhFQr4wIU953FRM3j
oK4gL6CJtJTjr6UF7/pU7JdmDRztcZeQiALJrHKtJzbQPnvufkkgJEGczeDsIyPv
oanIB+3OkIh/OZIezJ1BLZ+iEo+hg/BSOeL7zHnRK9O+JF7XLh/AWXUjvyJr6z5v
U+amL7JWQz8k6uSMnkVzcN9hFgwH1RJb6d7muDudlxyIom1Ta/LQKzuCVRxdM7ju
LqfMPr6o3msvnGdPNbgEruvept1McZilMlpTdatiC3n7G4v+xXRm00oYZC+KwCiq
UQCIqqBgqR4GAH20pFIF1+oOh4mO6JH7sUajLwTCzFRqVRr7LXLmy11zlHkPXRHN
s5Zw190i8wx4MdV47Xk5mGTGBL8eXqYpUb9kdN/9wqUL5gzG3/6nc+j845resTRr
ZXmxSEfUVcCNTZZHCI4rWh3KucQDMp3KZiMqQQ1BosBTO69HhGras4fSH/eWIIF1
KSsUOgHjjnwBTlOyyvx7ztQjRKRUG1HyiDU6lwxx/5yAHGu5K9lKGhfIwY/UMj05
ya2HYLvIE+BjL1vxWBkUJmt/bLHlef6AI4iBLoBxtQlvy1UZEsrLJqKhq36t5286
Epg2eaojpMTz/za4LEYWSvVRzUcHp9BBNTxFoJWLKhk8Ci+U6qsvHeN8r9aiCuIo
MyiFFc20vHdedzI+6IL2y5PvdUVonjSFFVOwDZ+Wy7P86OIQPjcdtoa9Q8R6wf3v
imXIVt94CxT0Hob/lJBDrTaM72qOTBjbcspiY3sOyaBtzuH/1YQPs3NWARRVlRBI
EuAuBJgqjCyvAXxbcYE0F3iXDLsKb4z4GPcmwjaQTF4IU4N4pTo+bSjzaJ/pD1V5
HSwGPj09GzHIphcNZL680W7WzlicU7PAH65uvvTn+CUKrLqg6LdkvLXJzzztTij1
TxqDbyTv+yoOhmRhLBJv+wn/fCbb99nLGjXpUc5Rb4d/r5N4b1LhwqR1SCam7r3b
810YFSM0rjkQxRquGTHE2q6bTKUpJLO7ACgjR5bG903bylRyS1ou6b8iwrRcfgoy
8/3nEYh5pfbC1DlBFRuesDAJ1BSSw/GG8Tz93B8XZhilieI1/xeY1i+B4/N9vX95
1lEO1m4IYNcveB5R0dFIK9ZyHItGyRilSrxtWrUeuw93AceQAwgR9ySVANdIVyn6
5Vm4jU4+J1Y5gMeG0BTH6Gdmb2ANCU1iI8+B468jRb6mc6DZnQtcqgNmbMC01gzx
zP7O2/i2+0VK+RfW9NvnJ++n6SLZV+y5t4t2J4FWMkmzE+ryRZopZ3+yjBPZVb/o
QvF0rQ9nsMlZbja7k70dFOL5hRge4KIdqovoy9yRXzpVLsGk2X6stzLnwwfxyi8R
eTjqrdqdk6oALmaP7wOCZuymHKTsm+6U9K1b5NPgkjRZmfCCotXwgrf/BOXKKBEb
dq30a9sl6nqQEW6N1oeYw+rRkiSyPRgiv5jQ6FmXpRxcU4j6kaWyIDwHRtYu0iWE
T4EDUwUBnz1IxJUjcLgNz8mczOTUjKpDnahB9rPeLgDQLF66n126o6Xa6ztDR395
lDY2EbyPeCQWBGM50AV3tQDRDMGb8V9lMBWz9IR63mlGBx1CgF1TQWxz6Kvbmg+s
2LrETGCdtE0vncbDu1JL4+I+VNbgJdaBa8aKpdX0fU94vjgChNWkaGEhAtHy4Nxy
aEIkdJoEoCh36Odyj19GUedR3nt5fA9CDH6SglIPOtCJB6fey1UbLzSJyzhCclrw
x8DcEfksb+1yP81kpeu+NlywZKknC1vR0wH6IVX5RhhM1otC6U4v/3CL/uDTjRMt
PSkxywuTdvtyDL9sBPTZDwtzwYU8jSJkJA/JZYonh9sK1V7rkWEygOytZlUi076G
sXAPManchfcvHjI0VhBLxeINLTkb1rBFa0Wr9iFd7VBOWgIW225KBwtjtrb2IeAw
0jDiE774hdyvqaUAgNPVznE9LPwnpq378SnEYfoaDTindwgyMn+K88GR3roxB+A7
R0QO+Wu3WkAzuwVZjsrS/7dn3mhb0bSozrITjrgx/M62mik+jAF5IUDzCDlKrfHF
YGuzBGMqYcv/gHj4QHT+p16Olt+exLiZ+43cOEUMyM6WOLkWQzarqD8jtkDUVEep
pUguSMulTYxT0J+kj2PxvLQKFBmBh3SvKtEe6O1eO9a3ZGiqBjBGGwB3P+EWk0jL
A3uKHiZWM2on8C99WjIQ8Y9E/R3Kb2VQkB7vUxq1U5ZPN7p7+K/TptdZqzm4Rdvw
NWTa/lJ03pFny9fB6fAwkw+8vFYrtdmP6Z6ssA8fBkAkwXiNA2MMLq5J1f/UN08n
r8wIOXMEeWO1cTan/03k0nzo9uBoUTpNzIDyzCq141ZhUT+OrVEG1SWt/s37XY3q
G/7yzf9njaKTwpDyJC3Qld+meIGlrVjbfsly5d4qz/XvNZrToaqQOBZ/NDeILW2a
40roScFwsVHI66pH0ZkW03t0c+r+phxlCL6npekbZyRyK0iInCgVxyj3hF2XpYcN
k1vpweZROdoz3dK9GmDKkipSjqgf3fTxQ/KbH812rrxqH8AkEnagFLRWt5eLPzo+
2csJZssKztLXyMqhUfrpulxmFvrr7hxL6bogj8AcQU+ZopUfRu1znQOCpQEAqiuU
HbFPwDsCKpB3JFaIjqMZPDUCgfwLiO7Yv7qClMEmbK3ZuaY3YSKBLRW+OPYVMmxC
o02NQjv7uUl/PxMgKEQyymZd9En2BGZdGGDjHF+PjAOB/AXJ4i/OZ5LghMPViQwF
xw7NqulBDRVAdLKPTjz0/fB9Y2u/7SMWei+Hgcs4tJyp9Ul0bttKiVLtjJ967wTT
Yznbfjz82bzPVTa1R5WXmCJwUEIPqNfyMlX+OHmKv0fMOLjkyNLU6X8lMeil6Kuj
+dRTrGrUKYu2qNOd4IK9YI70S61WZNmsMDS7P/0SAU98tMBpjtEgeeHad2UqY8jy
rtTSPcJ2q3QwBqpD85nTV7ahF1p8NYrHfOgxQ2v0D7iECkBxTBqauLvD2H3UtLcw
ZwxkEI4VCjcsYusbFcLmwiG2Bc5ECzf1zXUjTpWDONSiXIlB8INo2FEd66eoSc4C
0t1dNK3UHDs2smYF2cc0qAvH9eyU4reT3vmJ5VsvpNYu85n3vETGqKEkx3XO1aeo
UASQ3+7UifYFlHmfNmjeMyllyvk6s9Twc7kTcm1B7/Af33CsbNTagB1NLnW7jfTg
Vl+atnE0RgWlgLJRFkL+UEFTkq5u6eHC4HlMwe3ykyfiLqx6hJN/tqR4TiIVxFQr
2u3Qi8Ay3uulBEVYaDWRq2gtMFhsF22osJ3+pmzcF9Dt39bOY7bNK/z5eZaUDD4b
72pDsmEVzlxabENK7F1KSpUw/SWYcgMfyitS6DIK6AvU/gFcRi1aNXTWqjSdHbSS
sJSufSb3PjZPWbw95+CnRgvenshI97rUnAbVJE58t4dv+ofhJfhb4Zl4SdHQ/24/
olS7247SpCX97lccyij3gIIamkzw4yTDRvwQysZl3hyEeGh4wN30Rz586yeL1oxE
tTieZCcAaE/Ezo8+9Ni8/j28Q+rmtw7hTC5b/qz5aLtno3gC3dQYn2Q6+Qo1GadG
w82W7bXwGLM3yzfe3nYBgtOoChuwcfgzMKb8gYbfSbDuoH1hNbniOqiK+Q+HXtyb
+E6+4U1b/7+bX5SOjuQiG5xSt0L+ouck7Dw5+oSk8cDeapTPfpp8IemwfFiPNzo/
5pG6rl2RamJ5xurDxYbd1SzvNk4InqbnxqVFc3kiKFy/PBiesNRmoo82wRqm5GUM
AWX0xXdN89/z37Alb9l1dwYuLa5nFnA4FOXRjON3df/BQwVl2iprdokiNc/2Da+5
UKlEHcbyYN81yXxE/SsVAk1sfuq41P3/b5F8ggGLkatmxaPgYWkOkKw/mlu9kvEX
2Ac/QzAR3iA1Rf56Yhh9XpCNMbocJNcbB1U0aaoCMql+Y1sO9nBjHf94gKL0SdXA
aoyu6t5M4k1fd36QCkGfeAOp2d4pZ4zwfXiChZJkeD7RA4cDpod6d9Tz7hbFQ9eN
KMRz4SNW8vLtTJSQ48eAxDl96tYeNSsRccM/XRgKNDPCybvW80lMvccoIM5nwu28
M0xDHOxbl9iHLyc2zync1fNQkRdezVfadPAyKmqgvbXTvJjSQdaKPCI0LhEZvPdp
kIdKAyric1eduDnFZjzCxxkMjJ0zNgHs1zRw0O3BYFjXHJkQOko3ydXuiul7TE3z
j8sbpCoRCGJrLqMSGvGMZr3hN/3BcolrdPbaxziS9++6brAtBiCYUBzY/Xgp+oSi
3celMFr4Z9sHEfNDsvAfCc6m2WUGZBcG1Fi3ZKDnfNmEqMMicZHY9riCfeIzczaB
fKHKqRTouGbF96QD/x5RMsKI/Yen/BWOg+JA+USHGahQZR1M64PYDgv6BP3UGnpj
RnhuBZXH4b04bvo6J68vBlqnv0mVTmuc/wQbIB+FugBJBUgsuOXqixagVhXR3qtk
C21Oc3xqTMMvZAk4LYNVJGJtGUjB9JlOMQYhMryoydiJiT57aG8Pm7t5tpIKKL+T
RejJi0XgtkhngwqM0nTNDGe7v9WvhGbpLacxyYVxd00y3Qbdm/vbux3bPBQNZQ2y
BZ2D3QrSOPqcCD2JTGyZUst/3o2UkRsys1EHV5VlTiWpwSFd/uTCvEaVhj9GTLbt
DOs08O9EeRLOLj+vZFeXE1GAx4OOA93X614D3QLEoTm8emebqfjjTaHL34pFpUQ5
8LpU3AZL388sZrBITcY/tWhGBCQ3+a32HLGkKmt6NoqasqZ/2FG7g5jM/dl9aqLK
42h1PCLzFo01nN/A6Tebk/iGb4K+jIZLwLOUr5BClc5J+xUcUPeWJ+3dc62+uGys
68Cqp0yN4dKGtGObRjZwgChlOr5mEKNNWCO+XDYx8xXOQSuPya1AFZ0OJ3G+6KPR
NbGJJVs3JhJLvIF5kES3qYJf190hrngYel+roDDSSSYHVaP+zS3k18175TRUZ5WY
iVeGmJvcwDt46gJBcw24p4LbWofhuG2p0G4a0Nidu6V827LsGT+FQa9u3w1MvC1P
C8YOfYgsbmzW2Lt+E4H/qypfqWhFkUURyACJggg1cwA/KO+dODd0hDVczVCEXuUh
yW+YNkb4kwitVZWOjha7x+Q3VFeKLNiUx7HYv2oYJCJJfSdbJ34HAAqfUphLICl0
ei3sgTLClNoLjO8MEbEfsp2gfz5dC1Ancjo2jL+pwPYSiNd3iZUy9Jw7iISqdJfQ
E2++8jwEyKnnYqwdj7v1H7YAexA7I2MKPZGPufUs4Rw9nN0ntqt672fp+qPtgDcO
EGoEB18agLnPMtu1zOmkyd+5qeZpSsfwtQkkagGwuFvYusj2qH+DemSJFXydl2Hn
NhKgMKlV89aG9yVPSCnb4XDVI980/XerKRrhEtZqvRlnfeH7jnjA8/OgXDE2DAbd
KKz8lpkpJGuXUwtAUZgWewNg1EoZ/p4cGkhdxCYstX7abVFe2ugXXIBfYzDQFUZR
aki4ECNrEnW4OJr+JT42QedPcGU5YUxGImXqjEMwLInpEAffge81745zO6N851hV
TYfFXih1cUsYB2Hm3YrW35fEUqcbE2QQFgCFYzniBh3gteSfDyrLL4/dhNSrf1uW
5D7bI4zFxc6Z5Fx8Y9iqJ7OclnNHK26eL3rb3rpoTZx+5k8PDHzRdAFGK4B34EEU
qfa7vCQEC76M16EMa+rx108qbpYeXPjF1cV0R0avMlYH8/eiVAF1+fQtWB5MCOuL
NRAXXAEXg3Gkvghf6WMHm5N7QKM1r0kOja5yHz4xi28L272pLX1naRCzX9vmQq8P
mLal19kEFqf0YhIKXQTc+cVV+pHypT8SDbj8wP+Yy6NtuMG/rsMp37eaZZRfyR9I
BYnwMVoJrolQrQYUWRTrwFY11/XtxS2MEpv76vKZbbEQUywrr8jMu/OP9qcjVsib
97NZvYHJfjgHCid4aCu7SLe4Mwi6xQBB3mTffgZl4qmJmdypwFjopaU+Jw2GCCXA
Fbwj12i9hS64Vb0M5VNH13UWSRxDVNUr0uOqyx4FpgJckpY0emcm9NcncBzRd7Xj
WhRuEB/fI4bd/TcQCdGZPwwsY0vDAd3ivBQkTRGC0kGiR1dM6M6wKJp2miK+x5a5
PJE/uLiL8EKmQKDZ6XQ0zh/MKpZEWoaodUhQj/dH5BLSPLMpYRlJDtL4GjWiexRV
hIKvvLvMtXx/TKEYblWtNIlZ//dJodTBbtsPygmqPAdJ3LFJBIfCvg5Y3P/Wl1zj
KrBN93KPKur0DkHem3Ig9CxRfI6ae/8ycxiP3fay8n2InOl52XjcG7HQXyflXAD6
uXmK4aihSWWhC3iaxJfiQBDtsEsWP4S+r5Yo/LeHRASH+6Bk/MdsnOhte5WlmR2+
qF0FFA9WHgYycCqdKZ+iQ4ZoLSW0cm77SsG4a5YFX7WlT1fd9o7d2maiBhFC2iTF
SrB2S2ZreQmPlQcZegDD4+OVXRaLjfcsbUujA+HsT9iVjEz9g8t0nV2n4qy/afmK
OwaoRJw5LIDvV99RqYCSDiyMYXWCQHemuxfK3QcuSVcKgmpdetGzHgwos54fx7Zd
T/1xrF53eHx1GZo//M5xVFahB/xChnSqMgHT6E+W6fVpFUnDkzvli0vU/L949QTP
16FMExX/fP6wdS1N0FbHRwIqK7LFT4sz2KoUfhqmq/8/qyM5ZMFeJt6oxza8/fAy
Vl/ieS0zt8tQRj1F+rChIsh8CRQ0F3Y193cNLVdiLxjNWWxMRmXUJFexlo+a9Nsp
GN337hHCsSmg4Z2zloWiKP74hYTflo6tkJTxH/n/2y7M+x0WzxBfiRoidDwlFwk0
nAyAH0c3YNRH1p0OpZomvFEnYSPUU95mWT+qp+OTOjkKziLPS7gKpQx0BB22EcVc
XypUcKfclb11/PCDpXdx1owY7ejOpqQ4t6Dyba3ChVNA+ILqoKz7nmuGseqttmZX
ush7z/zGTa5g5XupLLuZXbnLQ2ZltdXSsedyJ839i5kfmP70eUko7/DcuyVClhY/
oitB0vVXfyYIYLsJbbbsWgtOb/3SjDSgBkHUGQL5Vh1025bkb6vL5PgOl9wbD5Kz
cN2QyLeAtMJhLaGYSdDYmu7zkfo/7vul9b+I1RmClDuwPTXpGSU2AfP9GDcNArDb
nULMPF7wy203VUFXgfjs0c/H8vBPY7iiw8l8vJ4pIMm/V1zhNBmmR8OKnPhLcN8X
dFGZdda2+PJ+yDhxD9UMjXcSl5Kd0thwKeVtm3XRm1lIqa7noeClXXjBVbARYkaC
20u97o+euK6YhjjuS+k5/zpbrefmdXCr8DNfmQItnp7+Q2UuhXzVttMAbp3kLsYV
vX1x02KszlbGMqKVc8WUr0G8V7LnOtX3X0hJDcYoDLhy7gedATdbngCxID6WnrH3
7HuRwKPO9JOitB800chKF2IcedY7rluYc9rllUPVRH/xyFzVs/c++gW0kYtaY4ER
o44jK31d+dq50UaoHV4J/BtaplgZh9KgogpUUAv1slPP6yPYI9OaIKvjxC8TuuE3
UcWH4sKqPsgHHt8j7t80P8qZxGqQpvd5ULvKcRwtRIa3QVVpXMRysyg9DfRbGXcA
squJtnPw5PYCaLVuxpN8I2piqAx2vnCqLBm3oEOWfS31Q8Z1ygTsodcYxW0uUaLJ
YaFVQDa1JCfkFSDgRHN2RnAJyJmqUWvjh3yMAIoCYL5cDJElvpvuje/bSZ9A1QvT
/N+rPof9OekTL2C4QzWsgvhfGMQwA9YEQZ4us9TxJX6TnT4p9apW2eHpTH1680hI
/vt89H3epzJh6JKpV5FsyQUuZagmSphdJFX3VzAlniY0sXylpHaj47aeyGjWo1js
4t1Iu8eYzQE+vNJp7nuSvK9/CoVb/Az3tfT73izqClpCpkRrtsHDFDJPCeOzwCiz
mDbaARMdgYK8A9tUxgp2oyrMrW6cJrN9JtH6J1DWcEP7JVtDNyA4b4rhf0HVoEdc
EuqkYKQHksNs5ir8p8zbC2YpZhLckGAQsnCtzOQXiTJBV5GHOh8LBB9Lftyu2FGt
0vlHG3xIl5tyvJb+GRi+Kj65HU7PDwthxbXmfcv40rirwxmV/prduhYfDThkuDdV
WL5aJJPJHx+CDJNfKCCu3GnJ3zhTTXkVlRGWtWBoPJCg1uDa5lSr/MumOxHnLPpp
7SIzTi0abpvKSMAw+shd4B39CGnh5/J3HdHldz7zYTIdKXKdsCdFNFpHXtGMDk1L
FNY0JcIcf0kiwZFbnBN2eAmVFwnw3gH6y1C+Pc71gU6b0mC0gyFsOQJ+nFsjUXto
2IotsQV+T7Hhmd8KpaJWQ/iT5sRWCuRwjzJIfg5lGX92vDIqmWHv1s1YOLVFTSPq
Z1JRj3WAhZHI7GaFvu8r++u3rcWm0IkrjwW5SZLTCcaKUM6ZZHbHHYXJ9DhsRvmU
d7ef/DaXoj67LE0tBbJ9oJsoXe5vAHEEMPkq6Qq70AP5xVLsLmeZGeHFvGkOOyL5
CNHSRJB7ekvptmI3TgpUXhfromLd1HlJcA6t2D23csTULd2rUZuc9pQS16AqZo9c
AwiqftHVT/aMFYEOpi8Pqc5/961Fsb8r9qOPJ4THF3DXGFRC7beTP1Sc+W/U4WfI
/CW9ImWE3vDEBCypjYs9Etx4Mucn3sfJdmna6A9itBNOfFymknTjbDx+Mzso3E5T
IEFxOiXRu8XQFtbnVqklQ/IKBSl7tRGTSwFtHT84iUcir9QkpIbLY0QcTdkmTLPo
ogSrIgeXu+dBUDpHaDIxnqY4VnTsbwPGwcm/lOcP+qzQs9/5tEEEw10OdZkaJrdq
BG1mmi9JKGumEmjpRAM4XkmqKb6x+2WSwWn1gN7okeAQgbmRVQpPiEdRijYpl+T6
XLENZytlaKAV4I7dA623hQpH2Kes1Ld+Em/Gl12xflRIqDIKCyHiTnfiu+ezbvdV
FNBiu0Ew9bTMAsy30Lolu/PCf4EQotnFdSfak6/GffSVLNsYxmR3biFK/kR2tWoN
C+29xw1Z1fhXejLBTGhKEr1WbTucPTWMBT3d9sa/G4JUmDgBbFwT/mO59yQSqqoG
d4e6/NM8E3uXzpkvsaCkfmD7CbkLjwmfGCOqJYC2svG25NPCcs5MECnIQmQKjypg
JF+C2ESlfv+3PAwYDdV2O2WSyTyLhB1l06/wNEiJESrd0ogqW8ugpNW6lywQzi3i
XN/e6UpOUZAYqWgyex2/5y0zbCxrDaBO6MQkdBU2syDKkwFUqbv7UHUXGOeZ6d0+
VneHc3peTrAZ5qtWHHo3Ehym3uDkMZ/LZw+mN1aJEZY3AXooNagaO2v34zxcHv1w
45IBPOmPSi/VkW2PqOB92YsppuzEOaPebKDp88Lmezl517F7i082jPZ74gtr70Mc
v7QJftC1mYjvguN95UQzEU+uh6s8svC3DiPjT5RKJgGvAlI7p3+jjTGSLC7HU4YE
GgyRVJ/jExXC5kROt/Pioe1smKQv3hGVDkRzqe8futNukeH6uRHZvVk42zuZ+RoS
5OEdgLkzyIKDJdmLfNElVeo4WJ320cQF+Zaulf6faG8UUTsBtw3fxkE084eehxby
z3JMIlly1H+HbJea2k/K78jBXTGuf1A96fBnZGB1t+pnVVVY2OjpIdNo98m1jpqU
O82sAeHF0UGbkZ+u2pxlWP2ft5jM9qOgS7MXYFFPP6GKyifbKhJGYnv60DtzUTvD
+PypcdivMzm7jGxtualpom6kWSC6Bxct/otVVIRVpDGlf+G0nOFPtF7PAXqzI9lJ
zOY19Zmi6q2GyjjvCjK0FoWNgCweoV4hhOTQWD5kylseVGvVAgomC05PgCpsGeaj
5PGAmcfJICN2fskBSAcMLLr2zH0GfhwoD/YuYwZ2tSvmTmz7fQrOyE5AL0PkYJV0
csuWmCtKLLQaHZhhCn0pDYNmcN7686pfuZmXIGOk6AzfYiGa2RtqE0qKz96I13QF
3Stvxmx9t9Jxco7tFoyxcEZncNzcWnAhjrFakSwonc2dAgAZU9YzVQFQJIqoVlem
8Al+CpAAqQQcKcp/QnipYPOj9jN/CQBav28t7wwTZT2BY7e2V/aNGcuGRdw3ufev
SHg6sy0ck0AROnsyiND7EVRaeCMjHGME8o3J1/6EuSHepSaGeyUcpkwF1cpXRs1F
PtkErqOEEOvE/DLkpTbPlqwPIdBC66KbmYB7GIYfLsGZnfZr8IP7QzGsuIG53sGQ
xzcHRTj01ftYNEAlIzUP+GbsGrw8vT3g1fvJuB+CpqHiTBMPCUIwnftMlmP3E/+H
7pe7xEnnezZqEor4C/Nr0pwF7NlYKPRSFoFcqepBOOUeQXVoJFiz/tZ9eNx8UWwX
zIf8cIyFZhSCTbE0z57X/g33/rEsAZl+JdBo3oRkZf55A9eC2X9ts9U59ofSiHhX
nlqJW5SXHpfFgzoq7F1tvVj1tujs+KI3XgdtsiNUvgV37a2gXNCbx3eEZx9dEcgb
eqVKY33qGstMg+pRtPPg6k2rmT5wzrbrB8M5CwWKPdGpv46io3EKLVslIQsYeynH
pMGdSw8vyLlLsVUSAYDzwQ+MCnal04RMxM0BgHGWJoVFYcCYuGBkBzfW6FZTNvj7
owXnEUHLftryuK3J7HUdXEZbIrDJyb9/rmgpuR2LzOt0GzDPrdi2XmNKJSahLX2c
ufzqXcnR3TrRvPquluSzIM3SFHLksoKSAwxONn0KPhYZ9F7K0H4QNXHGFhE+C3YH
UPrVD1+EgdZfw7/n6wIcErBeYlR0kQaHwVXGcVGnhYWmiFTfMavM22+kq8FBBtR0
cncYgSPaf9MEL7/x85kBY4+Q6oPK9vgapT6tvDZxGeZTjAXxqeHkk6Kj8vyvnvT6
m6XFax5TiVAotL0vgePsA9fio/19XpIM/UQ2oHncdaESpKO+pRlWcx1FuYehmuWD
U3Lady1EPXutEjjkuQUwbnSQDVSjqGhOROBpwdxdMBazaGMRuWXLkHY7MdSyFwea
WfUVTKeDEtyA8obSPhR47BmYSflhXrMbvmtYWs0KCtnXxQ1I+l9UXyO//Wdf7HlC
RB+3hnOw/VGd5dbY/duzjVWLqe8h06JIzp9AFNeO9YrGamXt5CVBuyDeuQBylw5O
Uwg8IC7nQ1zxYQwqAxGr4nMRMHg8ePf+Y6XL0Kidoq4S1g6F+dWhu6u5Wi57xmXM
xBnwgSzQIQ9mpdlAPWJR/k3hQsUu/pHHhMUnFria7D1aIJJcIRseDkvGytHR14QI
sVZf2txTyy7chEe/VJXGSH13lxpeoAPBRE+3jmKHtFbwHUFzWIrNieBDepa/lzH0
pQF+SDcS5au+Qv33VZM0Su2fw0kPO011g21jVRI0R4qMzQkNQ1pKWVRoBlixw3qK
aT0luejmd5p5j2ThLV0A8JVdGdhz9RzwI1955D3iYKXKGKssyG8MAlZ80D3uD8G8
kDXWpu6kSymF9yRMXO1S3QtiH/XF9QW9KgmmWx6K1xQex4Ugp/O1yI3Jcddok6nq
w8kOE67iqKjzN8HYTfh4y2aAXOJwoFVbrFfqiGw7IRKviHpBVcY54XOoOOluLMp7
7Sqp0nNJ4CdUj1fpNHI9A0undP/oJGpSd/y0Vow91tmF+ctshx9PiCZYGDAEy/4q
GMhiVHvK54ugUEX49o3z6ogtWx2OOhxttN8lfExrSMXJG+SXNkcIRRNFQSsmoaZM
7CK2Vmy/DKJqZ9w2SUzEfCLozfYk1RI3uGUx7lQTgGK9O/Sjl4zhxl+WJ2ClLYsw
7v2WZQoD2PW84XRpP+SAqzX6KEQFpeRZoESKNlaRLGYWxrprxsUTtcJz7ZA5+uI/
ytoh5EuRTLcTt5M3rGXlQvT9tVtPfnHBJ09JxFjKJOv32F/qLbnmsswQhuVvpORn
VnkwGU+07S4kEeCibR1DCRpEJP6qKiI5NRtIW2B1xBbBKLN9KBDiyTlPv1hJoCkZ
/OjlFkJSgLmKb75EgOXP/gOgdFjFwThG9lQztnkwruz1YyEGNG1uw9X12jElQrdK
1sDPULae0crEjAVZ3jX8sN6KgMiko8CppIJJsIupXSiluoWBB5QCzTzO9xxMX3gG
WiEdIS+QqeQuG6z1e+U49K7FKVnz5cvFDkJ+z9Q6NzMXpe7ss2D3d0zT4DNQrTSN
mwT3wA78ml5LbJKc1EyPvMp2MeTSlGKaNjim2ul5xo1xjG+Dju9M3ACxJmMsC/cP
m6lSAvb2EC0qDvoua8c3gH8dMwPrgrDO+5Np88rb4tYAf5F5eS396jpF1iQoYdkt
R5LJhZs6Y+lVA80L7R0wQRhCcnrm85qmi1L64jgEgF2YtfQmoMZ4uIOU+9mAOBbk
wKInlfx0m1dxtxsuMOq0+hArzbWxDFieW1cUBQ/aNliayPnrHQ0Ktdi6kutGUJVF
1dkXJd9epQASpfKwEGpix30Nc9FfuNDpXyi6JbMg7hBsVLLZZPYrxbKP9BcWP+9D
Gub4luc1miyfUZiDSjdHzMGzv0tPoabxVir8Vt2PsSHA/0KB7+WTQOsRdsictBiE
66RMWYvr5rAYCTNMy1x5XZoG1RpC2iN+VnyW8Ct2F60ZAGCY5Zv53ZTC+abX1o6j
hDqWD8AONue9Hx5DIVi5rTjPmR430bUn7glmlsJrpISeXk/WVURgDB3yi+wcN0wi
ZUuuOPZDf7QuE9yjF+GaQUoJnzkYcRKoUvEsalSm+YTckpfemykYJUfGROobLwV1
4frqbSdcpH8i7rhYITIGJnMGZP+tLi9wyS9wKmyxD/NdOdmMlx+kfvn/FMYvAVeh
L1LosStYNBqb5xK4sWj0nK12OoX7LcCJedC1nwBBDulw0lNCHwavaP36Ukitqtvs
7gUxlmnsH3ofHilDLQvlgY+RLP2K27LaEqPrQBzvAqzStbRt4qjK8o0MWcEXwmTh
X1sHV+siQAODAf4ccokGThiVgAl1DEHu5vAdhu6YviBrg9YGUFa6wzUXBhb6WMsc
olwJSBYod6Y07XAZAj6GX47T1xf78VvDM89Idl3CrBbu4BiBzJ84NCkPV0Jey5KD
xkTZs6R+lLCQO2lomFCqRxrBYKx9dCLC/Gs4hKf2fDpMrGtDLloryo9Wqu3a8+GT
sUFfqGgfBSYa9kXJ+aEB6/dhTL6I56OZLUVIrO8Kg0ZnmPvrReq+BRnVE/8f9nVj
Mu/ioDg23MNCinz6IiqJQEfXeCIBvRznwrLocEvCyu1dopQnHCOfopv/SIFjo2xT
MJ75cpZCF++4mdKfv8P1/jy4WkgxXXo+dUO7PL4+X8Jy8xWWjDQXl6MYZ1iiEUNX
9AdmNNL1UD/JC1MhQ24V8C5kmzgvKx/Zvyqu7ggcyBHYe6X8nobjg6sxDs1MsXdr
AIudimrh6GMQd7COB9SPajZM8pEUsHFlTD+PA1jSjbLyeUTheua/g3vpPqN+QWua
IHu0KOvS0/T9CTp7aRbBxihQIYRYokuGfDKoejAk1W/k2t2AD1txGYg7o72gH1zE
sZrQ7GVe/zNIpCcBB6/5ifs4m1jdrBlNPBQx+z19j0K2EptDAzTAnUiTyInVoT5o
Ch1oJ50Bach4dFpHMpAmKlkSnSavqBBXILMSnw1QqIf2FNswtS65xdfiXTYTeSGo
ieTWS56EcIWdETxCY4hIPxDDcHM1410ja5PQwoFrKxcQCqyu1yfTi6XmdDUa1N/u
bVnCGMhSqQG/7PAAffEvrv9UddkSCokVWoLnfpelh2xf1Qp15mxLpxR2ehpPAI2i
gBV5aTaPuOhCJ8EGKuQExPTXauZIwygUPhKwzY8hCKg6FEzXYk14/6h5ymbCB+uQ
Uae/eSm16kDj0BalGGuEyq17ptkLdt5mWj/+60RO4thawPdDn7z0K7rXojPCgJNy
/z9ZmGJl6A677p8P11nLsxWrxVRiNjHo0Lpom3YKg6pviUCGCMpgSEkP82kgcoYb
N36vIWj6oRzZHmVwA8RK5NKUngD4lK2Q1uYyOr8Rcu6roo/oHTAz88oABUr7SkBT
i1nuDr9+GZtmR+b1bBCJUcxVoFXJd4g97jOfsx9uOcsIlGUK360biBz5NvtjcPiM
/rWWseeQjb1RMiZXNyJmfG7ITlS00ia6giHGb/51llzlyHwEiYeIfzMChftP3l8E
/WkvTWwv1Sz491kVt9WKIOEYb3O91u3gabW4M/QmGDols9ElCLKRQ3gqcPksR5Uu
mfqWLkW8SvNUc/3Qrwh+24+xOqpUPqUG9kX+XxH2vIyiZj+j6DsOkFJWQLfC9LEt
yyXo0g9dXixZD9Tjlcto1voC9/1UbkA9nXxpOWfoGr1gs0nfzFneD5kICwUt2Scu
QrVY4g5ub/2dzEsz/fNaEum61E6wYtQzJT+FJOR1CHzfAgSnc2y0a5UU94nWRp5p
3jmmY0V0979PERpJ1ZDh85Z+Ib3jXRKeDr7sQcPdAfjQ/FNy0n1PvdmrV5yYQM0x
9HuaVfESkoIQqRcUX0gZiPKk1qGR3QPKE79vySmAwB91I06oxvQxHwwZYoV4ThAN
ysTzmAt+dP+rPgQAqfISBdt2YnsCXxaedL911TumM6rjYKQay9/L10iZNf2XbWHD
tEviXkANMNpiW1Tq7c5PEp1k7qcibEOqP8xzt16tGMOsih3m7vrR8h3TIC1TgEQR
rlKJlCf/P279vOE+DghfK4R7CfOBaMC82P8J53+TU5FVHcPbywiEDsFR2XWz9Ydy
l2BWht3PtkVbxftZLNuNhSXZeO8hMohgFqq86xpg7S6qr5Fc7iYXUWNDC1KrrR9O
4/lfgNJqH4CuMWYuzZSwm9IEMSiRP68AF/jj453K6A2c3nwXfA5XMuPFeKI2dUY0
AbSQqNA0R9X4p/GZqq3GyyyFpWdoxtn37c5VOMjUTznP59xkn9hr4NSLE/cHIujn
sEyYJFjBrl+/w1dRSmNL+Gw22rgVxgkVRR91L5FJZTftAxLvggBz6/PYUrY2hWb2
k1CqU9QAXl1vA7Z1QiLb2EBfnnfIYoNMboIAEVmOHwTa5uEMYViqfcaznbTI1S94
IhorJIgmXltcAjC6mhphdhi757a1XP/vMcuIS/UVCwlvGMb4zpTBXRRWVZEr/RKo
tXhRTZbqk30dBE1l+mbkZo9ezO3hBd6ImyAy1o8Vkm2iktVv4p7gjYkxsy5CdYQj
cWLPQWM7Msgyb0eeNyyzJgTafD1l9f9OewgcWARamI3rU947DGnxJWDKE2xQDM9J
4KyK6bGRpMm9SfggadAK4soRBl67U5Qdhf621VKyoSWEkzvaGMn8W3xTVVE0wYMy
8lkWAebAcgH9/8CIoXLRozJH2TcGe6JQ2i3Ehv4vmjiQrPTBqXDrBTMeli/bram6
JBqx2F2dY1t6nNp6yvUIiILt5cchUsmyM3819gqvOmIZESDQBnWWWnPJCrdUTNL1
RYliV10uga7B3jr8bnmn84YP5AVL8IW/gHxgayRCQdZrVa6kYkTfZ1YKxt/t0wDG
9OVmlYMwL6YK+RC72N/PQ12EROP7NskudUzJXmaoq/uNZeWcTFi8029Nor57Tza7
YnZq1H5ck3xXaZceDjlZHEuQVOCxz3Kw7B9M0NEx+XYAv2vsyW0QZaX3EryFfnin
zddHE+Xd8y+j4BOPrZCi/HxBDeZU8eB5+cWfAeI9AkxGWw+abLZdBS1XsHaBRp3A
EQB6w7TOy3RVygy2EJNsvf+Uc7FdhgW8bDVTbccZaMwS22xbenkMvUhbKvrw0N6k
oZlwtQ49jxtYHV/Xt2mLk+QwEIQAfPKVeXjuwJBjgKgR+mYEUhjfe+jiOygPgqcP
EhLnNCRVpUK2FCjuC+zC901oldU82AHyUb8siFym/oMgjDkXt/D/+zxiwgIBswaS
YmAYOcf3k2hPcxQy2PmO//WY72dW/4FVdG0HhwWSVfUr3CVMBHsRvuvyM+ncsIMa
wG2ZD1uFQLNlVXamFEGWlHV6MMxvFdeOmgpRuRDNJPGcTEw5FKcxfOnMpgFs5kPJ
AYATUszyYRJKFe4hLMuCNB7BsTPOKVXp1+8H+kgRQrZN3+kqWPV6HCgw0DZ6zAYg
gXZKpjnu3kDXoiPGOMtCDGQ8xQiaY4nAjqJdNcY+O6JeMiDsYDkN3kPHoK98D7ha
8tOCvVkS+iPxg6Bd0Ep2yYnT9D5nZmFxhjQYkcBYofslrsJ4i923qW7sIpXYgLi8
VfHCU9SH68rwbBnVduCFem9l7+tQYzT1vVo/cTVh/TJgGzaft2UblliSzFECd8oc
iqk7o4p/5gcW4v2Plvc0bga4JIrMT70GQj5yUHkHVHdxHb4zTyP6mh91wl0UZppE
ab7jlSWZ/yBnkYd3uOdsgE3Po+lwbZrv7sPXECZYIivJvEDnmht3jslxZnapQuAv
6H/Fbo8K0U+eueGKhGc+m2gJv0dBemFHh5LCU6+LwStwQN/Y3Mz9fU7gZZk0f6Hw
62Ux9USl1tNwZ7pCpKDGnKGWaxw3xtl4+/5RFmoZgOUqALTIAnWQKJyOm/stYXUP
TLxjgsuQAtD2GiJHaPkKYbu26wXs/1VzgB3OqpYgC1bLrsW0IxWiDK81KkOwVoF7
TG6WMwqHvtVMJ1O3JoB/NbTHfzhSdAFzEp7Kb89eS4EB1YYnn74t0kJHb2rfplbW
oGGE9LhEgrZyHiL84pfAwFgsUVbs6VDf8YTw1jeMapN0HmSOCNqRC2K/yT6ISaGy
/3wt/vo0IhFzfMc2G8s6UGVZ5Tjbbex31+3sHs9/ie8FD8mEQbgMW+LR9Isu2E3c
iNIkqSh7aAvH6JKojyaY4YVMf8CIMVEvagxbNsLmH4kQND2cemp9lod0QGl9MTni
R+QEjtfpUW68KzXKz7WoOhKRIc1dNY7R1UtKmVQ1Qr3TiMzycUkxc7UnhKqXNRQR
mJMUPTsJY152GGy7Xgcn4Ypcwz5G9NoB96o434O5HN66NAdPEilZ76WMCBoddzVJ
kNw5T2vimtnipa7M1+mpZDawermiNBXmyITLw5Fn8VsVYHWTscb2/xWSdod+tEsM
KC4tEDZJSPtwRaq9yU1rELFzr5TqLUyqmqOT6CmBqUO+QXs7Ojm9gEVI13q+rrbF
feV7GFXs3W5D6pzTs2w69w==
`protect END_PROTECTED
