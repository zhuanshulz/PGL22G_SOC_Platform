`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UMvTJSJu6u5628zfbLQ5qG1zHPDNYymeaeKz9tcmnAgJ75dHeusBhGL0z+Os2GD4
Fa3mXp4g2mz0FXep9Qc2jgoWLPT79YormMVw8Mls7Rs4HIlD8WrhXNjwN4dDqsRl
0yvKjXQnedevYUkkqMNcgZ3rTWycId98fhBcb3mJBHA+bn8zlnpjyzRAQ6YOGrmi
TPRC7OPla4nO6AOlVI2fFs7NS8AK1dLHZUikTsxo3IzIHzXWCmt2tof00qlrJk4a
wdczcEbVtlrr6yc9Ktvmh20Q5JW+XFPduIb000YTJBjcbrhKerGxjp8mjG6OP5jq
wiSuSBE9nzLnuHKmViSNMA==
`protect END_PROTECTED
