`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6FGvsZ17c8ZAx+cUr1CfrLFVu2AR1EaTjl6CBoLlCfHX/M5qQg3KcVmki1/c8BUm
KLChEzq2wqX9EtRAgUNX1CqY4ENZERGBZfrCuXuWkoxQnuuLsbBQSec0scBeA//7
3lc6TB59G5ntKaBORH65Y2JKS0xsaM01cAvIU3RY3o9jKwuUiT47g5unikWClQS5
ZTTOhw/mXWBAfkOHHXuOGymLEo1gJmWpyw5xhRvQsQi1PWUZ3x0Cs+CIr0Bec6MR
jYNooQYdB26uuhSZvPdjAYeUWI63Tpr5uW0l/AOqqg55EsivyMujbN0A/Crk/Ddp
J1/H/eA6r9KqO5iAcB1yAatNRVn2cQEUGHVwBvMv4Ifu99LOLnXpksIsqykSIklt
dDQKDVu7LRPQs1XasnpAe8vDOxCXanXl7107N7o7cz6sgZWVUIFXosgXCxJHfV4h
5kIXnAzXTDdKvfQrzuGzbFI5IYl/8rtvAisGlaJGB9WxLSB3VvMn/0mtM1sb+1Jo
R7JozgjhE6fbrd3DJMQa8FVQu59pecqb4tkH1eRuju0apOtlzFTXi7xkjPU17b7J
`protect END_PROTECTED
