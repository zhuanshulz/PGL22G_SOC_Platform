`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8aX5uITzQG2xZ12fKbwkMNKcr701YhX9wPm2UQGswzEzxtUoRhDO9EEEiu4JltX
I9yM1zIFLxLQVdPxk6TPUVhLz+gc7GrKT05ypdnydGVYO+XL/fQ9/ZiVwGiI2bck
LbHAhKclX0dtnCclBO7UrwqgnsL3jQkQMj/YgR8LdLHZvEbTLm3RPKGMAa6ypIqw
DgsjpFnx5cKYCOQca8CHVqU5rXfabh18wrU833tZUJzaSpNvLI99c5JuhDIvpDTi
gRGIL6HAxDZ6pjcVfaiankHyWX/ViM3Zqj+ESZ8LFUdewuldRLmpQohyySauJIAC
b8CBMrsYzXIR4tKM7UejjSOlIPkgOTiDzzMb8D0mRDKDgHn9n1szi5/PR6TWmAAh
Z/vbgVTm6yGEl6HH2z5U0q+vcGkfjCNZwxAEXeE9AhvRLdGVu5+wOCBVnHMd91pG
W0cxOrjsF3vxVpweoH8ODEfsOoEFx0PFdO0Su2W87KUXcl+lKP+waV64b9GKN9zs
RFngWvHB87n0jhLfC1CoFod06IiIDjI+LIiq6z+Itkikkvg5/2jFFbb72znNKJaL
kQ5F0A4gBVhnOHjA8GkFgRnKKwpLUsYAV7zbhZ52M8RcXndGSSRDCFpl6clwmzuB
6HNYHZjTPkzpwqhpeavH/XnyVZNzQ5abuWEWsaDRpyfHuNpaCZyX8fZKOETlsnzm
UJRTtzQlIpC9qH7qrTSVeQZw2HE2fI+SU3+VFEapMGe3RF+6KHaXTXOWqTq2Ava6
AMugp3VGZh+lOEyxhaSbp5Wyspq2bta3P1p0zxWroMs=
`protect END_PROTECTED
