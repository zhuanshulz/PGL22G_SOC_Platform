`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0tBVI/MBOV+g1GqZNmQ7KVYT9BaJ7saIOA4cLqjsZXI0QY07NCGVZ3IGnn8OPj5
Di7HOAFu1+3H42uc/gSMqkALgJ4tOAEk00ZtHPmKFhvipNQp9jAmS6VYLG/H/c+t
VTMIPhE775CEGfRM7oQHcXS+oyC9bkEcEKxPVM5YkJ8+J6R20YE17aN+nRoo/bJI
sIPXyWFoW7l8yO7VQTq5ZqSxEMgrRGuwx38v2opMBe5q6b/Tt7CUd6kJxSCutMgP
mAXuiO0Ny/VFy1bVYwg7Ca7x/3EBl9Qgi9ORxzqEVQ2HXkYXeZf+yttZVnUY3FLq
9yTpaRN2I/vSVGc8yIv/rKSXqSz+ENx+K2enyZBd/6V8oxV8UTCzT8hIiWiQfMPi
BF2+s6ZY4+glSmk1AvqWAx3rFnbh4laHkThcSQywVPmRQjEMjxlrV4ZN/1NiZOu/
14ZOnMpHc5zUHgEpVFtYQJDItuFuvYZrPHYWc9j1liGK66eUuKyQkhjxjY37bUA2
mln2iT29y/I5J9S3Ma1XcXkS5anzJFgkAGF1S/1bySTcgXY7wOGn2HkGqsQiyv8N
HH2cTYQTrE7wL1cwqrzYHvwgGLcTiaXdDnuaWeBBQyVAGYhzlWzHo6CTzAH/qu9c
9ahEWXxr/cj3HTmPDfy2yRuz7m1qzuvRbEBPu/8/YNEMoBKdNVuXKvwty2o6tCKT
pM+jHicTL2tow7kZTo+PeGolXLdHAO7GnvWzyjs3xT23rC33PNAiumqy+9/RJd0U
bCsFZjIbBx1YY9h4mwuLBVfZ/WVUS+MWFMnuSK2YtqkMhUpnkY6ywtn/ybPat1X9
inoieKGwq4o9B8ZQdQOYU/C2rFtViYEjfJkGqQ5nsznttNgf+bszq+nRLq3f9RAo
KSp+ZT5+nALEP08D7/mWNjM8VFxlj0wm5Z2uHuvIOYkn40KTz0JZi0lyapGDB79x
i0LIF1cdazGWfYfJl4Q6wx/8Kxmvp+kZ9lcDTVLdA6mrAm1ImE7E1HjsRy3nfaDi
XOy0qXWFvDQd6Tm8Lwej2/FX0qVqzA1wVHpJhCEOtKfeRvk0l9EYQtCvGzdg4wZE
fwVGczuah+Yt6Maw9Fm3vo98pxabSivunsBNDLxNF41d1w2JStVB+SOvFPf85jkc
0OA9jSmbf88JOMf4n8r1R0xuot99Zmr+SaQ33c/wn/F/N26cWvHWWoBuh5Io+2T6
BCliwRsQWc3JvHaAAq8D9/4pPOslmLV7xWBpOMMIWgzq2vfdqkul7lXDI/29YhMB
iXFw+Fnr3pGDnm9OEXGvrf8BgAmPg0F0ei82Sbt6pFG9bGnp+nNdfVFakUC2+t2j
G7CXUb741Wwn9YB93zEyJ1yjzcka0XMSY67a2M/rHMfx1LHP7ZAhgnYAPbKgCIP+
pa+0dQRy9VJu+9ktU4fo0BSIoqUtcJx6C5dShDDeBMgo5264+aDv4sP4I7seGBU6
cN/GH4kheLVtQ1Pbvmfmjq5TYA7/4ydiOoVJfmth0rGj9XRn1Jlg5CGIH+tyN/rw
0ebCed1p5rd1Y1rb2LEO7Dwcgyjelqd7zb4PQGm3s4c2sGWAk+5odjrNFkBk+Sal
EovSY+BGt4zrQb2iGlm4/eSK9ep21NR7iAP4Ki0a8dBWFF/eH9RayDQShuQtFHIH
ZHdqFpAyhpcmZDMJhrls7eKTaSrMfuVxzDWe0PAP6lZOUN45kAdwfEbZsSWxnCe2
/whQBIjSB8B8RpF8H0d0pJrUx7y8o2eCc8gt0CKDg0j6AR0+RVgP6hQ1nrURHOx5
C+d8wlepevuIAofmp/hlDHm+pWmeL94GQXjz35MgryDFmO+RDtt25dl0Kjp6JNq0
HbQaT6luk0atIqiueK+3F4r35l+YUJw4Vv9ynH/OnpMedT009MMZ8hMqa1xK4lss
ZrmYzJwAGwFndM2fMJDTz47ldbZkQZcqNsmnUolrnNaYlPG1reNAoHQKIDTVOvB1
l1C275VL0a0mJCSIBmE8GFoHC7EFASemIab4hHa5BUlGyOLjt6HxTK+5/8UQwHeP
Yw5/l9jWO6+tEjK1wcTnHKnBDo2v/YIyI+ByN7WTh79PK1+/DjPTYK2I9p9PSEAu
JwA37jfdkeBPogZA4xzwLgGdpDndXp3aIoVFzippvmsbcOAjzqZNkhRZ+tC1La7Q
otNUR4zNJiHk1E4aiBDCCMjXz3SVO9s/YY2FFeo/fqVPmnDeGsg+t2+ViR3Ud+MS
oW2xc0GC0BSkW8hARGqjIE/Wt3zTT7coGmBDytDHMx5LXBix5XUAGJNFm1qTzKpR
BDSZ+WopIDhk74T9JxxG98Y9jsR2NMCZZXWoEx0Qucs5uCxJb9zrfkkzIG//l05T
lyk/dUofn71wtHDBEXOGHWd+F+uiZvDlz6uWpbZm+OMa5nGrO0F1SnmzAs/eK/Lu
lYw/crtTAdE8vbHWHk+PZPJrMBS0I3amUkWmQRRLAgiS4XweMe9FW84YISIU5lAf
sX8l0HcrMGaEXUDMhTNHXf1SMba7kXx1EKO/gGvUkwxv58Qr2hVF+xVHofS3YMnR
E4nlAgk9K7LWbj435xXm4SpbGo8XfwaenbdXOoR3rpC/LviagBBXnb0dCDZpR/d1
A3Z+3R743qUBadem5Vq6yhimaRhMk528CnCq3tnPfKnaZyvc69JMA/tqOdCO1kBB
lZ1tnu2K56tnL0obk7EZ5RP+/D2CDVQ6aZ0jIJM7j+33AiAVPMsVAi1t2KuLrccM
3zq4vmnnVlTlAkZpNCu4cKGKXWicodrt07yXyjb+uPwReuUx5marA3QoYghOsrML
4RQ9pf0jFY8WvKlBfxB8Ii0VGns5gzW8MDO8fDnoWp8QyHS+6+wJS101Y7ctEIuY
7V/s7C7dHzIMGYqouFo7QPFo0w1urgOT3clVYYxc2omiqMZwJ3fN2xMNc72yQdwQ
fX6aS8GxYKxHB1JS3e1NezTrEP12ZECZSXxB6Jeh0pUa+IBA8lUpuuAxqMn77XZl
R3JfWCIuFeNeRo/ujywR2KtVEVwNV4sA4ULQTDJQg08gQ+aAR9dU2FbNWAmTEW58
DOKf/ljjPLT6pojzpbSOP0V5IsxRxo2giYZzlWYPQXsAjFwNNhdNQ5kIrAbJGiQx
nDcGIcTPmbtLZwBEPkQL+TBy/yX31R1f/bfj3nVAImV9GtRhHSY6qo0Iv49UEIKP
qBKuagzXQtb8eQGf+X7ZKGY7n16PNP/UI+g5v+tIWE3PD07REYwjIF5DIJwU+Ip0
TKO3eTSSolCyNw0bLxu/wURKyPDAe2eeBpRINv1TBeX9cFW30W7FCWPVXcHYoISV
f2s2BPnxio3Ir3/sSLu/Ec8IiH1MY4OtL2KiUmHUIcQezlnwmTz6+D/CJIJnqAbv
0XNiWqqmhrw/HX28X/2sYWbigwhGL0iTaD9epVgpJYYeOZRDbYKDnr4o6dp0XWdh
cSAuZMvZqKtVmyds0W3/PjNX63ojk0CKIFe9cZ7y0nBH/ikqEtppAVwbu/cfeBB3
Mzh269Y/oHHqH0utPCjLV6wViJh5O4/I+FlLsKaQqZmeyugT+Uj2HuP0PFh/Hpp9
M8IDcnlsS2MLSNrPXzNEeue0jOD7qX6w0DH6r/qeLvo9e3j8Kn1Fa8R+U3hEGTI8
WX7ZHREgdNafQpupVVrKcGXCBkcnf5YgHdKfbffBBu818bdMgQdCJbP94Zm2bC+u
kbtRYzEPeZDn7fcXm9irgaQ/MeYf2yfQMeuDsvNmbX1YOBCzvdszvlQYKSBb0v4/
ZKoPDSe/uWdkFYlkNRz5Og==
`protect END_PROTECTED
