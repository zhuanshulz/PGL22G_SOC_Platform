`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
haBjQxm3R0S9Ht1ZtHIzIXRWe29TBi7rE/u8FMJfpnyS/zLn/7naTgaQ5JrhzvMS
DlDGuH+10LwklBP4UrX9IA2nTI7dxNY2Fpb/vuH2VLqC63+3c9898m4eShDSIQWn
iqXqE8jdmw/Y/LOz00EsvWDTJgX2Dqc2OUDfmIZIoGnHqOQUhWg3sf+wim6sglcV
CnZUn6XQOXA05PTPoO1x6+FydFdf+5m2Dfdq+/E62YBxE/oskDbPzFCpY3A9ttIw
6DitvuIjAq8pGr/EpYQhtk6ZTYJofd+EVECGXaYIN8wRcsxiiJdU4jsLsseXydEF
OciMd0plvB0MQvmfkSGgCYYQoy7NwIWKBVcC/ObcFRTGwJE2jt3AJUN4fpowwm0r
nh6VCPLFTJ2Os++EY+llFgs7MZ2obese5KAnNNwWc/waZn8Sgr5PA2SBjHytCt/z
JiUrqUpzq1JxtOxKREPly83Edxe+m+IFu49zvK6eIjb23HQKez+G25PLKQaZW9WL
posTq5YoMaofi3GXMB3ZnpkQ9SLYy9H7qaVVvEuTzAbv3L/y34PUin86Duk/kAIj
ZjSuvH/IudY9A9lYSbYWWC5XQ+eezU0+VMmZg6o1CqBlv6nhMFuxUAxSUpAwINMI
skUAcTuzBMkURGP819+bGvuAm3LqNw0XSC3Xhz1OncBy7+vS3gxvgAvrRvQVKAi4
puaGkNqHCTJRn1nhjp1SbUvtnxm7EEvzTkWruQTp+0fF66SD4KkZjfyrhYHMB1dT
ZWnk0PuiGi3EasYaSyqmr3WzmD3iqObbEDR7+giKlvLop/JoAtt97BpbiOfi9VjE
EXZFKW1wIYlU1QCIE4d0haEOtd9YHHlUn65VQ0yPd+RSj0QIoobEbrAsb1KwAHc0
gRrW5ULrBbmHZ6CJm2ROLCfyL5RSPObzkQxDUvES4BnaUWCRIfrZ+calNZxhs05u
Hb/8nU+Hfl82vpRzB1eqTJwXlq2y+dX2g7QUyuonJD25ZY4C7hWxxbQZp5G610XU
h6butn9/f7S09AtbUTxjz+e5GUHGRHJrW5vLkxF0wDEp2V7kYKWJ6TJZMp4uctF9
0UYn/3GT4bZdtcXUz3Jn7SNfTp0O6m6HirNPmq1/UVwstaVaLltyloitJBRFVLzk
4SSLtT9eW6lX5eCFJ9tW3hzGFqvsHQw4AZKPJwsnxWE4peTSQDI2LTuOES2N7/dB
PxDKZDnUr+cX7rEYyfZ4jW0YVLoKUkqKi0O25xnFx30gwD5ygppAB3qGEucNee3S
B/PmzG4xDxYMO8f4K4DdhwuP5VZF5wjT1pOOFq2qiQVApSLk0AB2LK7IwcJOke6w
fw121PsobLRLGEydaOugN03PEjn99Lq/Bmhnle2MztJyxe6cTHKNlW6nYdxSdnt7
AetGbmpea7frdwtayqQCr8IvGJgt5sITeuKzAvf3HtWzpOmwXmTbyvLaQL22SxvL
II/8d4v3bI6kfGTMm6Qn2FflhZ/FcaCg530GmeYIO/4piiPM2vhUHs0hB6GfPCbK
jm26aBRWdtn5QFIqHWEQewbMKJQSJSxHm2aIgwl5YgFljqOwnx7fL+KpPQ9ceQXw
fF7hy3eZCzwRyGZA+zJPd9oAKRBqmDKpUalv1mA0FVQuwxk9WY9bvgPkmvuQlggI
hRvLrVwjaP6Qj7V50CHZal0888dRMVfDOUiv3G8Plc+MQshoiHL6jnJ14kQq2bzN
KsRGbVGgILTmiz7q5+el4jY5FSmLGGcdeF+eOekutYq6fVGYvlwh7Z7PgUBgAvey
4dkvnP6RA4a9XxVHRUrGoiCmb/e05juxERL+m2SufZOnOMxzR3MWVxoH6iZam6ac
1HaMnbanzFcEtjfd7yNzkgJqVf1RpWcOogZ9NKzUF8J1oY/idtobtipJ0kFhjhm6
VubFjo1O5hB8Z32QG2Z+DiCY5e6hgMqv69HZgwztyWqccigv+zZdH1FADWCRpqPs
a+tvpYp5LXf/+uZ4akm7lBVsS6vD1z/eUjSRo66hfljP6fFsrP74FCpj/Y4Oav2j
KP2HbqkUsVMjj1Za1K8FTxyoIp2KMAnma02CIABuNxui+iOx9vbhpAXSWKCGMi0e
3SrXjlFzHkS5MEKf8U1y0Sqk0zO98CQzFbc1iwVDW/luWcYN8RU1EqzVHYEK33gh
c1iylqq+7dQy0qB9TZzstIU/bIE8kWKUR6CavIWojipRx5K0TJ7BrULdRG5W8wwE
Pr4tymIV2R2oUmnPgINg4NKgrHW+tew/RPHFQuiRR7HTuRvKgAqod6Kz7qDwOSsc
XTrgh5pxfrSF3zCdF5Byk6y1YVXeuuJIZlOGDlTey48inHWVV/anE5H5zpeirQcD
uiPNrqoaiGM4pWMZB9DClmNIZwt8lBf+7dXIlBMDDiFWvzaKrJ15sWaH0qiIQdrb
uDXS/e1wki+Zw08/LbKB4Rab4BpvvDYgPdjN8ighi9SfgsGx79y8487zk3qMqPcr
fkJq0oqY5dAywUobCALn+wC5XsQCFN3NRvBRJam/DS3CZKpcfamYDGxhHPjMNWrx
nwogDy0sViGxjZpS7JN3X9Kq9boMyIfOosgg1gyMdjRFqw9bImwvInSc4LsfTsIS
eFjGmbwtFgKZhyRfZazcJoj3WHq8yS2/PbrjQbVVW3EtbuQvwezajlbkATb0MSxp
XgtZRzud5v6retMWnne65/1FPHC4viyxvUSDmDJfU9S9ufPyIQNn1epbkpBvhJL7
GnVs/azrVlaepsB1oLj6SNuRwLYvgSmzDnxH+KEh6GMS0b4hyvbGIglHQH2IN9+I
m5WcX0IwoJDJ2dIesNpb554g4jMm1H8GREjLLOalm1azHOQNGFA9Uq+gW5OZekro
XhOkJ1bbqloyRdW3LOGG6lmBUP6eQD57yQkLkjOtO3EQB1LUqHkZBcw/VyJQZrBM
p9QstWqi+HzoNzSiXA7KGTpMBjZK31Xz0yoWRZdSx0Ki1E4xMxEwOUXe9MymbZwL
ui9hCVjBD+8QTK5mloKQf9CpR4G0b/pjXkPQtobReDsYnaRbTnGrc+fgu1q+RRt0
zu3JlrNzsOoF5tx5YfcPFzgwu8pUyG1lqO6TKQPuBbmi4iO65y4jm6LqtWjnX13H
OzJzyY1nIChxSYElqTRPEYvNl7ZIa2tk1AEGQUzeSuKKXnqowpHZZbjEtShRRVv5
0JppJQsD35ybdf6FAv7hpIg9J+Oj2+WBk2l0gkl+muGbs3q7w83bT8ezruO4vz2N
IxfMsLQcd5p6cmqbIqnH10QpW8CtGucu78D+1bLsTlLzagOwA8DJf6i3EsBzvd9j
iGZGXIkQrYA+OSZoR2LNlmpueyvfkWobY+hBiC3xoH/WcZth8dCOn+O6OV8zLNef
sdR4dsaieUhC2cadoVXx0OzTNa9Br9GQHVJpIinll1ImDWpyLoYNajY5JxTtGGQM
ADImVtzgxIe9tX1931UoyJaCVE7oNcPOpxZgA4h9wCVTtMJadCsxAQMojL9peUTc
KdQOIPtIPU3PAn2nzz0eGvMPTp5lGjoJaUD3y8Isv5TgXG/FlvocI7ijzEsV6D0j
oOakuHHLPWehlJhs2vOrjPqVV8efSr8STa6CCTIRICxihGo/ruBRybLScf26g9xb
W6t3MefvuPVziTfiyRUuLVy3VpJK+tyZxaYUNfT0YPd7h9eHLvwcq0hk/X0fEnvj
X4b83jS2XsRZ6z9M2wYgVC1+RrvT+LADT6L2q1ppXM67a4QTd6mMrMad5oWFZD3U
MxPpASa00MqKfmiNCWQ9Bu0aLtwrYIbrRwDmlPKBVXhtCXj9QQQJVC8eYayB0f0r
H/qcNNGEb8fFoIOOTzQnVbBBDVt7Ah9GJ8+WFSKNCwlo8co6vFuNI9Nn0v3SeCua
aIZnDJ4/T/ly5wVMtth7pK/Hia+EJyneIgWfCGB8t0ewMvl9jIpYp77cQlMPd7nu
wG+E3spUFDo3lWq8gPo3TnUY/r8ScrtLNoHYcluPpKaDw6OkvtktKCohMbV3PIfP
0B7DKkwWTIAcXsTACDnt2rSCyNtHXn+irc1U/HO29CnDJkti076EXTmh4h0OCdIg
2DTNutehlFtU8tZAq1VnXtl9ir/psqKuel0ZMzSBo29xpWtcyy3RprCF4XGuFBdF
kCOUXLxM0pWL2bZzImTB1CNwA5Sc0plouFNZCN1VG4p3U6cJue8aGNfWpeF0eBRk
fE/7zPNtZdPVHfvHkgwFW2AV66GGTJFw9pOwqzft0Xp/lcMPko1FpmxH6HtlIpmX
LhL4OCdP+HDVUFM98Roeap7m7plDyEAeQr9QbapWN5KGZpvTdX98vUIBX32vyE+d
OPq7u2ebvpIqxGnUXy8JZER/pH/xbdxi9M3yA4Jf8xl5h5VTa4vBLKMB5la8s9ZV
vV7Y5286Gw7KPG3skT1AV4CiVN89txRVeD+U9d0UkZG+uNKgBLNOoVS3JjQRpktP
48Rd9giiir4kycZ0Nn4MOKce4bZ3n21a1tl8PuKDAXfP9RRsNWv7A6MyYkweVE7z
bEtT+jXs0tAa6AywVOpVS84nRcEGMqt3wbiKkkD4i5HT8ZNy1EJJ04iVtKqydM+P
aIKCZjxrk1fWDvthIYh8HCCWPxDLXrIY/KRDWdrIjGkAw1nwIrvA7xLfXnjFxRYa
WJXDRx2z5VVsBZ8ISKlyUtRKA/lvaFZhzSmgWeBf+NIkOjNi2Ay89ZeiNyc74fQg
387P9TH/PJW/fXwQH64/x7IDuMAgobnW46lMFDwReJIdgcJMFyKTy2MsSdA4W3P+
9/EnFoRHXFFQqGLj504JNjvmj5NjuNsxE4eY0Zd/r0wZJS5WrHfSgntN2kL3whc8
MJ4JAW+y/cNdw6yi9RGHfp++InW5WuTvBBGUDKPTieAh6Or4O741Mkhnb8kg86rP
hHQyD1HpzrUWl7x9J3f1UviH1iSx9iWpkH8/ZdWCdD7xSAr/fHDflI15DbKJhSMZ
Jl5wZxiLxP+KCGhzDZVTp71wh7fqOjI7YKbalYSwiGQXeQqHkGdhf1IPjeuq5KVF
m8+Kk1BY8nhG/CassC3uArSjpU7+fhU1ZKcBOA3mSUzKyYiswZ5fP6gCTaVr6ycT
tKo/05MB+0wzMlGtVELrSPWePOn3jupKVF/3bIjeU/gpQnosM9OZPqLilJOnJDyA
rxZA0RpERNi9zCqQ27/JPFBEoArRWsd+IfuAYgqIMnWmznnRoYK+LpYe78eKsr6+
/9XvjJ5gaGyqYw/bAO0GTleCprYCJgXpZpmOc9kf6wGzIUTzdjPBqm259IYQVcWB
7mEQbStVFcULBVbcR1GPsp13s0eMvpyEPcMjHgek3wuafz+YeIqp8i9cDTq19mYe
Fvdog+Y3qWwdx1dWuN7KBXeLo1UZLBhniJKU97I2VvcJXFuz00QuKuoBGxq30Fsh
GB+VrXgojgUpux56uDu0BgYYB+BEzARmHk0P4t7SrJP/LYWuWvGBwzKGRFAVihM/
T9SQuQnmiv5daa6fRfx6IrJb1m7pa8LTM0iGQcrk2sx9jMARXSEqJpoWghq5Gys8
u+dFnOwGUvI8jW86vWIQWhchpvblDX3gjOTr1OZRc9a0VMMRHeDvC3/M8zZPSMqc
2pllmb/4tVS6O347Jt2u/XzMadRVkd8TrxiwuG3qUA9q5dNyFnl6w6t4CrgS4q3R
bBcSH9eQstrk5mquOCtuHBxjMrxSKeShXAaaA8vBtZAww6F6M65kgbcewaOs0YQc
55HGmh4weWKlpyp5np6xu6Qx/0NR523lwv0c8DJ3e6twMPXTsZk0froVbwS6nNGn
EPubJyAwKQnzO8q6sqpzn/8/eLWyZ2WC8civiDuRRH51luzJHybwybLkp7VA59mB
xk0T9XrVvGxpEo+uTzxSiSTt57PIvloWxWWybUQLkZYGGyvsngsxDCahaKBo1s4B
5Dw5kkDHXpFgsmXP4QVB1OekXbahJ6rpLAWDIe/AeILuIfkSyaWihVnGXa4qIhZo
VPuR3T8BlA66VpDeAH41oc0lBjklRJhwG2KD7o9y4HD3dH9YL+v/evCUQrszErQj
CPol2RVdFu7FnWr/m7lcTQkEPGYSuTaO2k9LsKn3l3+QAqCxg6pbjdBnUOqDpeXS
SOaCvISLBD97ubXoTnJ24PhEi+9uU7GofrZRzDpOHcaAAjFzSANB4RB8Glc0J1O3
uOgQIddHo2RyqVuYwwtX7PHasokfjzU01QVjhVP9v6c6bCr2Mm5Lf2HVnbUul2Ok
hgPAodWGU0WCu/IB/4eWojtJRMp9931YC3CopicnCQs9VgubmFAiknny37J5XFl1
JNmsSMKZo2TZTuBoE95SIqjShvury/wGS7Wa6QPFbebppLULAxpEbKVwMqPT6qzI
+Q1voK5rgubNvHyknBZdczdQJyDVRW2PGJ1SDUyzlUMV+DsPBDU2rjpzdthO9bYU
hvhVtYk4ZYYHJdOGXknyte7oPWS5rMkdyDy7ykTI7lLYgluAFuIKtz9s9ovz+MEY
aTJZeB88OKaNKVcaY+lhK7b7qVDPVo1u6DLx36c7DPmrj3SOwOltCH5cPiM8Emmm
yhCTgRKFmcYbzp01uM6RdpNGZfdgCZ67D+Vnui/NwyHdwbuPwPa+JyEGZzmp8ohj
Wgk7QY2FpkYLICypaHdAI8nzljDx3pXwGboHlUmi/7aqVdUJdooXQgWv9bKMuuoA
jo3Eysr75hNLB9shfZhAaDx/vqwGzNsSEg+fz8ZzOs+xFc5TjTap/+dsHED2k8XK
fZ5aScZu+BFUn495OLLUzqli+GXQEA3qCbtg4CRnKLu/HAVGMcdyH6dmZ4+Nxy+k
w4tII6GLcThVK1zgFZbGRb9fD8P0hXiJ8zNTT4bbLVLCTvOjyE7nDLhMExTjM2ny
Qg8ztUCABwcfU44X0DseCZJqBWBtKG/m4Ph/4iquZAYLg8I3unUoJrRbJbIAgypV
sgc+SbBTXosCWAj7NxYorBZli+B8BqeBHkfr+hjSewMAbvECpQPinvvxEGGo4Thk
30X/GPDNlBdmGSPsPtN/QEr1N57sanAzgv5TP+VpKXF6xrwTQ/JR9kfTVPzd9ALK
HCrWWjERLIN/f0wslFilUVX4Gl9JOmMIfLue2A0erzfNm+gvVikFJ7yvuJcwNEzk
LllxW9/NFtMo5b+QqJA53g6faANyZx8NDGahJnrNDmoj8+6BHeoeKDh/wN2/0/y+
JgHXqQTEQUO5XIAIzWw7BtBv3PTxnqh/isufh4FuP3wdLlFZMTx9Zg1AIox0I6mQ
nJ9U52w3tvecEK9Mg+P60+IZuphvbM1zgyAQvEL3QKTFIuvo7QFYkuO3NJ8PpHK4
62zrgMqjpoCTiYQNcmjaBi0iyHWo+8BDqUIRUADSh0/U5GynwtuyuffUEs5tTe8b
dK094mU2YberE8ovOG6PWJqgHzX6kjGy0WTpelsSYUz2riU/DcB7BwCJqkOzSmLP
1wTGjF559oSVCbuZfk3Ihw+ubKozIy6DmoYNU/z2A4RnZ8rg1ccRqlzsbGZJIGCA
VA2QU5TXRgFfQhKyAkJKIgA0EOeqvhecBuFB/zjvEnK9puNUIDJijJR4nbHFjiEJ
PfSHlBLuiS5VXMw0mO9zq9zCJDPau7eda8r3HVShzP7XpUxQ8MRpLCxAoH2gE1iS
ksAbq6fITPvGa0Xj3Ge81Rd63uh8SlL898TDG43zsbf+IHgU965vrqQtn4Qjt44M
2Iz/b2D4i6PognbPCib/8hheQRIEiY0XU15LjPoy2MPZNe7f1wELEHiMUgabij7z
5oP7r4PJ7zmhxaoz04hPTCKkZBwyZtCC7qSMq7rCMXauAQkT7cM6bcaIaHszhbAH
CNGISXPoa/RWGSVXqJNTaI6I/MFdvf44aPB5CUCtv8sAhYZusMs7i+DwAk2ZJT18
MG+Hcvd9XDqoGOOnWhgRCtyj9oM+JvSsE4+mDtl9LQ79ZFVCtERhr3YJkys/448+
HA2S9/IsgVIwg+r0EifoiLij49NiU2nLXgTuaIO8k+RomtW7qsGBlruR57Vmo/H0
shXI34JK+lBUVva6StzqUoGb2tRCxocHWiG70dy/lmjrEl/l2M3WrO+FYN9r+ERw
TLSufSg42MmRvCPcU/o/M1CHAmJZ03+aeebfqz3evWc04yeR8TXATdrraBZw1yWR
sxBBeO9SZlKqiJbL3jHAJ/j7ifjq+5dL6Sc5DBbNbjQWQrDNXfvEVrW5BD0Xb7yI
svEwa61+xcgsheuVxVKaOERwTINZLRFgzH7WjuvQYnXvRlHo5ww2DRDRCuAbakcM
8ZjxYU5m7YXXeGpokExtCMrxMJHR3BLj7DtilId8VUfAM3SofHjgyeGcMCcW7tkd
70ZJ1WGXLd8sP/vSZcrJLk7HjjiYF+jRfpOC/EZDDsNSwKwdqHy2VsUe3GS++u7U
k0vjCdT27BV+wrdRKGUIcHFZ3ib+vYOsTPbv9ShDyjitbBVZlJydqAoX7/d9l6Xe
LQzlg/msaHiSLcmLc3SNcWN5/Uj6/hOAYWXr7Qd/dhJY41avA2zN5lTMSYzfrBa9
/+81wBUqUxQ6+QI3/F9q5SDETLqHD/mVjj/Jb5tgb+VZk1LnB0MnRPYHQg8XzGYZ
`protect END_PROTECTED
