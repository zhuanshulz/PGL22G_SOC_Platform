`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSJgtAt74QielbLUzBF8YJRe+C5gXMux7bBqqVyaXmPfTAgP+yaVFZamQMH+0E/1
+eYk1ouphfLH+9VP0wWiQaLK0uV2XluWuSVRunahDywLKls5Ki4qlXEuGhLFrLpH
NuVhFVu6H2qyg0PNDNLoUXEoQBi65hR/6bj7N2h3p4qegpX35W6k3AmcL5c4y6Qc
/5m10z4N1htq6ye3+2XoNZprecBTf4zlSIlA6XB97V+UywnkDZ3gajQ5C2t3ZCm0
JLFjSbVnPoWGTlcrKUWsMsdRz79royOCJAyGRYGUPZ8ZJEl34lCxoTxPYf4/xFNI
WUn8h5W6mOu+ws79QHaxrhSkSvH2cYcbOMINt+3uvT+Q6p8JK3Cwqd8Zq/mQuGRI
ddXQnYVbg8i2p8379RuWSGJjcOdpwegug/3xxUhNe8D/ekfZafdPqey2Ovl4zxF2
lC8SdU4100JX9zR1ULnbW7wdalZFbn6isXLSV8hyhYx+FJdk5uAkZK7OkcdWMHwW
85M4/kSdmCxAexXyWqGFxpVlA49wQIMpLQZvWIhu7uCmOUtxxlwhvmewqLLGMwol
XVC03DWfOS0RDgLOWKf1IuwDcraAZ6BZZFdBXG0UNeqQtcpXr73bihV2UkOJk85R
iqlceg4WwWRqp/CPFBUmeoLk2jDRAsrJzHwKW0dq5XulahFdMP4HngnPyCiDO0A8
xEdB41JHXJvud/AVFTTdrHU/qyfcpOZC37uXWXtRai2KydDNJr9ZpnERaOdcgbaE
JMvR4hafbGiFU3k0oZa8HV+C+aRTPC5XwlrqTuxRYGg7QU2rIKpsZKHpaahf9SS8
2givepTzdIBDiW3PoAlQ8QsMp8+ADimQYCnPzlNFAoG8xHx8vHJkNikteRq8kCAF
kZPY/Qk/laPZPaXABuU0z+aNhtbHyK0yt7OTaB2CtWsWutmcKduIk1abvJ0e6gOT
NuCSUmKwmEpwaDLHGt9u8x8SZCinI4oso9tooQXUp9WCtjXPzoM/loTkMpQt7+wD
Osh/y70dnXO/UZiew3N08wzVhS+QHFShpjnvhAqZRlRz/UIXkH7E8+FoOqS7/SCM
e2mKUyapnT1/to/qCtZyVeHdfB2+QN1T3HBreNzKpuYKfz07+qtmt9uEN2BRfwrV
Afsdm3XrEpcNcvwu4PSubt8fcavtwD4sFDK9ssfpA2nQ1SCy7yoFrjJp8WBFWuBq
EZHq6IQQAf0IlWYy0P3b3NUfGapl77eLLMc5yzeKaH8qZkG5yIsKn04bAhnZ53sd
PXZQh1tQGJvu7dqo8xwJUE5ug0s1t7Jn+h7FAu3YKAundOeOuLGAga4dNLHkG4I4
LP0rrjKP69VzTVzazyREE7SobEoOqGmDQDHg9pbXA6xu7daZ19qf0XRTXUcyQKUR
BLiXz/Veh58srJtnRQaDDcUTiPNtorRZNOvWIfZQ5n1xqAY4zzNkimkhxGY187gb
OQ6VD/rAiVAooVj20sM3jCePP9w3Vkfx0rgVZ0M9yNQ7eI8yBDRMcZXebxac/zCA
KdQY6rWnOx1fKS9aSOT4z25L0CAfEfAY4wSE6STzErmbQoNYrqOyelcBu8x5lfrB
cnoXQm8gi7dc7Y8NF8vfDYKLxjOtVQw+4Z4b575C+k9raFpAfXIMuU09/yZHTcn3
IwiAbDqlsvFq1PrRRtRibmrQVhEjqc+BClmd5Sadm2EPHuPI0+pWR949gZDuehll
epgG8aPC3uFyq//RHkQKfY6f4lBC2xG+ssb/JBvz7etw8rUi9/4X2yJ6skxW7JdS
CmZzLhxJzmOtUpZtZWCQQxp02xuu4LYeEaRDPnWXmvH1q0l5fqvahL7WYVUIHjr2
iaPVX1J5RL0+IjP9CHiF6GeIE9bkN9IFb4JcjiSkug+QWoZY9DtRrIEhfuIilzSE
gsokgs22tCLEONOv+TXBg5EG7OSF7GLnYFiyKLRR4+gx1xoRfQ82IL3i285H2Wpl
WDX8Fj5ZIoog2/Y7/h2Su7mCwxjk5oXUSgVre6AthQIPJBheZ/LOQKGoY0cMMpAO
Ezy0yxn4xJFf7t9ze7TdltxGnwiAf/SO04lEU1ia0VAV7oue6Qw4/ULjGHQkC4zS
zBAEfCc6TqJGYS2DNVVneSdOVWEu9124j0LF9DrAFBW1+CUdRYzkin/dkq9kM/OO
Sy6Dt0GeEJbArm7ya+YA6j0qkaJGpOvAN95lBRz0kawV7oWsILyGJ2VBtcW98gw3
aBcAYRKTo/cTa3+vrhQwMdZXtUgkEQ19qL2NdQhdzztIasW3x1zRO/1u2phTO5u+
CQEwfphtjVjNOT6kqazNMJVKTO4TKYwgTTAGxt86qmnJzZHHbLdNZU/XmG0Kp8uG
6wbmhJ/AhkBwV5sh9NKN3vjDjCgRjCq7tTQOI6KldMQZbalgrQBsABAMVqa4csr6
l3ajyz1U+xq5RzUMKLHn4vLAmODaxJTN3Zb1GlIi34EaMyuca+rS5eTdh5x9uVvP
jBIuj+xUEiV2ZOhi3kKlVauCoW5Pko7ngZ0c7dDInElnuxLokMFFyoXsBTM8VI01
+6PCkvNpZ2/l/n8pzH0UmV4lJfmtU/tt/4lrjHWVre04aBBjkOfXQ1CbDMVTslK0
yVuTQpEyNi0hm3BWLh/GbifAyPm4kGJuRTLz7cNH7CPiZ1xgbd1NIpV4yvkFRLWW
BOAf5+gf4DhnUrkXBFMJbhAUtp/ZFiv3vnRikx0rubmv1Yc8oBt14/xoT6lq7qi+
SS2zhlOvwPfVL9BwGeZnMJKDGmQjwZjepmzGMCSVY2tglXaNGfgkCQxfnTPCre/v
oR6AkY6i1+FYfleAmfWTxEzqBUKKAk+6mqMIiekj808Vt6gL3mim5aeLO0dvpcm5
saaaImrFisP3u27vug4/Avxw4Qf8gGhJd+MU1wWsuVoA2rMV+vSGmB2+Y9rajkIL
WP5j7ztvadpedQRHAZMNme9zdFEMCsAZwluTdxVYwicM3b3ewnLaJxVa+Kk05hVP
k8lXGwGi6ppKl00Nw+qghjTSiRpvXu8dPxLBjVqd2setpF0y/oDC3p7ABNmJH1Pn
+iXaqhOH0Woanj5WMkOiOalIWRI6Xib/768NDd3bM9KG6hs7FUOe+8DBGcda625V
nlmN0TTg5c4R82jru9FQ7IyKUmSyl1SA6vHsQ9hSy98lswy0uR2YnnHN+3v2SraZ
Xc5ThlNXJmRsMAuMxEwWrjMpsT4v38i48KFdsYss+Z8/fDry16ldPMjJYe4o1TZh
nkKW/RyaEKTEVHgMbQU/qlW7OP8uJrPuAyRz0UF4rkL9LwQQ1ISd72QV2fYXIlQF
QOJYpSO9z4Y8cELNfyINbIIhoDnH2uj79MRzBt7n1A5Jrv6B43a3LLe6kNsJ2TWp
zbLBHhj3toV4ot4K65DilZPW5i4Pos3qna2OCOz4m6icqJ80/z+UP/TzRVpLdwo1
IHixI58XJ6GiLIuAGJXhYYQpku4KplX21xpriQoHkeaGCP+z3TCqREDDHJ+4ucyQ
V838xALBByEr+T2Auy8rBtFNzZaX6bVfT0towtEyYdLHlABJBIozU16N651TogU0
GbIHCO5VUjxPd+JKndX12Mw/AquPZLoY96RTrE8bRaYHyU2zHI4fNM07OqTax5UG
FVK1gcpu3JRxvLEqOslet08BH3jq8IM/X9xwpoU/uWW6DzlODK9lKw77VqHh2SdU
NFNmpZmOvxxxNCG/bESSNLGeiPo0VzWwrMUOnRawow0O7aCtpHpLYh2TRybEKMuf
G0ToBeMi5LtKUwdwm9wRIFj5A/SusUFuRqDrAmSyR3dN0dnOcZ1Z6cF/oaVV5zmr
`protect END_PROTECTED
