`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ql5TjK2eoZf2/K7/nCofUBG3B0aj0qdrGl7YITqDcWTI0nY3a673efZOfl/KApMe
uvX4wE0OlyjhR+QJzbZfrHHRt1Fx+EJ9iatZ4mHPM+bJSpfia1xqMB/8mpQc+n/i
kdpCPqzSWLM9nTPU8TvaGZEl23YS6zOoCVRjva+fQsIY4+d4luvlEN66e6AFB3nR
5lrWIMAVb4jPDPVZEokiXUjZAOISndKDhAxGUfHI5OqbOQOpMDnt96v2gK9wJ9gS
QNfpTkNXiYXTc1ehVwXxNkdGQI9X+GCvjsZFH24QgoKKiYWkWzb3ade9iSGYVp6+
W3vckxeeynocyLM6hD4pZJaXrAcXewgzyxsONmkBOV4fbSzIoQ7Zyo6SlCsEuJq8
9OWEb/pbfyw20eL/DkSzICFYZW+nc/W5cV1DnUAcYvCF85vNU8iMK/jaVC22LgUj
hU1EGUq5p7FKAMaQwdfDevfHrxs4Aho5HgM3a2/InmyBuCSj6QS+26ClYtwhSMMi
0cmk5P4n5v0vQ+ccKtKjJm9vs064Nhu+O8G5gztSmYQPyV3rOMvnANYkit9//gym
QjDOR64LmdSPeIpq6bwbMFWpOxxC6duc+WGi3SJCYRaqbXHKamN2FXwbvToQvR8G
2Hk3GB0SgxNKqwFFLaKKn8ctLPwK5oKTkw8K1ItRnrs8E6STJq65+sZnGwHnuezG
`protect END_PROTECTED
