`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0QwGq20bZVlNta643M3Lq2eMh3/0q7msRJuscZLG+iHIhiK3uGJ0WiN1/Ejl+U2X
GKYUQjv63FJKfuHVckAVAymZxe7fb/QSM6nJtnx6vzU1/z8us1sqqQKxIeUYZ6K8
7RmRobQVkNn9rEgYhXRqm2/PLyST3EAkAFflrvLfWxLEaO5YdcvJ6RV+j+sGM92O
DeInW9QDcZEZmBUQAbkdUkg1cITlzzznrQdKSn9p9cKYUvp4R/ZTD9O9zPAnRbwi
ttkRLpsul6QZosLsBYkKINbJpJz8e2s9sCaSQCzgSRMO67Zjlfpy4mJR01EakwXR
jOLoULi73FDboEscukOhPz0PdMTnFHqK3Je867n9ThWyBEL+KpBW17dg32UfcEG6
pofNfftFlJRyxFu5Sfn9WG3EB8M408ut/BzQFxlYkSk2BA0J68AJ6axewTksmcWx
0SZXtxyildXn9XRMqyWWA7rCNAhb1XnL+pjB2eRnZOKA3Sh1RQBrLa3Ef4SgheCC
WsJHWdzl4gMeezmuTQLWowQS9MRtxf5UBcUVFcQC7gHgD4l4tfaIv9EAh0DfhLXl
IX+FPrEgjdD23HxiyPfNRx4Bt4u0o9MBVr0e9nzOq93Z8W+7xY90VN8E3sRbwDUC
lHfKPCubI6amD4Af1zlJk0bg6GgXP3GR1QNH0/ns/FVCx6hGCCvxbolzBBFiHX+k
pvligokviD42MQADI4E1Qhm0qqwhk2XZWxGa+6VpH1ueHobh0PNJZqC7x6oTjV9r
3aIbIJEL+ebwIb8dsM0p6dk2Qkgrk0fuhQJbWDquxL+Q/eXp0hkoNezM42dn8reE
tl6M8vDWc3nAIira2gYZQfHDxMLiYtKaM7X6TJSCJ06YtmL3Rwg5WoSbN/DKhxp/
jb1rGJVlsYqVRuKVE5uSrd6OsbdSIrlx5wioWKayPNLN76yzWm+gyMiEjEmfBAOS
oTE2WZ7KCD0kxa4/7cTVQGlFXyZxS40Hcp2buIfhN0hRycIJaNoDNiW5kRwJ7cft
QnYHV9FDOLjDX303PEcqBmFyD86OxTvpkYhyd3hg7g2UEe3Ms9U6WoWcHS70Kjj4
oxU6aKmEJ8I1XViVWFpus5k9IlZJ+F8Ap/qRw+Rg1jf0hQmrVO5Cmp5YaFPXuBy/
a21fV5uCiJk2KkCrkDgcmmDyjSDEF9mP76OOwMxz63mzXfhH8yhTLjwzuQ26Toh3
MQB7fl7acQlm7oD5yXvdnQiqdGHldutObrGtetR+jGs=
`protect END_PROTECTED
