`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYAWx6zIx4FdFhSHZY4HL34OF1XRnTI7m5pRdtMjevclAjJA3tmCbvfafRFt9sgQ
WxoComT/PHbfMHNsFPWo99unH2rcLZgmYC6tgtyZijJfYbAA+zIe6syOrCwdHIZN
ZBepC0cP2fi0kbDtVLDsuc1WfN7koQwqX3XxfmCjtTZbtui4vyNodQsyjQ5FVvOj
x0Fmzavw01QCdxw09vGt274LVAZkfS1xpdh3W/vgJ7K1HTbBPWIVnoUuc6VqXu8k
o/DaflFN7jJh411wHtrJsfkHAd1L6ikfNUS3wVLOtkYjAMLwaR0iu3wjOvmOk4VK
5Z4K8vCQWwJ12jgRVXFqKjZDep2gJhpQoZn6cyeqPim2hCHV1ztHEU7GiPov1m6V
XT20kX8PIZi1BP67kDF733Wz090WNGpv7l2cxANW3gGjnxynxh0nlTlU4W0g+PQ9
Ex3Nlq3VVoZdib1plzVHOxnn1h/f5yUSBaRUBiUAFrdk5hFoYCQUH3ODhereQwX3
mnOPXqFidwGRBhIGu0v7FcprjHBySo8aFDMFFKQF9QMVT8DezTB0a5cC4h53fWBu
MA7Mzc+JnhHaT/drJ0p7HaIIUvB54ancDz17RMMzyqh5VNcvHoG+r1zQ+y4USOdX
B8JI9+odJt+uilAiW1pGWDqEW+cuBM3fQ7gFf1FE9T1OYyM1wUIaFKMq6krzTvjL
l8qJjwxWgWLOo+XH69GRTe0hkpaNQvmuFwypX/SRfX0sMhwYuHuj3Pnpj4A3L/tO
jAy3WOMO6R1mfCEE8rCNkIjvuVgMUpqUKwewaxFdnaxR4MnbI+7tNb6rA7DoXLD1
gtJudCWvK3lirYoqsXIkbB9Qx4RRKteWew4YzL/lF9mDDU4sMd8izNYBcE3r8qUM
qx/T3r0P3iu2cPnueP980ni7SJScqNeEJI3QeDEKeoKVj53BIzNtt0zjRGak5iMb
eVKN3wUxFRVpge3c2e4n9LjgwxZPHr1zKFr4qTxuU+3wNJDDNn8riNqzRC1sc2aG
`protect END_PROTECTED
