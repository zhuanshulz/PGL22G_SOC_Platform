`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gfs2eD3gr/x+8yvQnA4KjsQ1PjCcn8fxKOPfFlGz+IOTBA6aHrqym4io91hjbTUf
KBB1TMXgADSnKiOxeB9D3YRowo49E2xAJk9Q8VxNVB4qCw+Suynds397T45x/P7O
Kh6cRlZJXsHEitz32B6ovY5SjMcumeJVOO2yguKA7TbfSRCM/SrKMLJSi0pqpUqV
u96V3zXlWpDLAHSZDu1/2f3EzPaDU8NfbXY41+xVoljihp+hIGCkdaazNGz5wMKx
If56ARx20YAU2rTLucHQ2/sW/bBdasu+K/s+v1boTjGn2+B9fU6nQ2FVF8pk8hhd
j7yvWFd8HUFTsRzQnZWB/A6UGJFc35AfOF9XL8dkfCMF+3CiVhgXKzByzAl4FNek
oNk1qO+RsieSf62xYE0q2GeaKHNstpiY0OjnZdN0zsQfCGq15Xq3yT32pmd7C/Da
hFzpoQVpjDdcLwFG2j8EQOT30KTSEk9SwDlh61YjmV41OrmkaVr7ZyPedrYxTFua
UjRjtGG4RroBjiuKrzpq7VQ8+0cnXHgDjM87qHUgYpM6Moc4Ccp6KiVdjDKipim4
XI4SHBxNh2EQCEN9dIp1paSgEdql8Eb4VSgPlMA1YYib/H5WuD2HWCJP6czxDPmV
krBBtWykPwDSahZnad+Zxbg9eQ9WsdgbAO+xEDeDQWFfXzVfMHYP78VLJwAXeKf6
DUlc7v6OI/02zbEtjXKbN4o6WwXQZhw5CfRoN2Ww/3AnHkoAVqG9BqlvU5W2fPla
ZfMfS3wciBh0KuMWZeHWvdKshhIS37nf1n2bmHSzCZg=
`protect END_PROTECTED
