`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/cIImSL5R4J9Mva7F4WfEyXnqiCV90zx5YKIGjuTHDLsOgARM0Kets7N1jMOixdp
aSuTY4vNhSFM/dkVT0lXPIrSyGEXx8f7nKTR+H5qWc1p/7Hs+/aYy+cQ64RzVA00
k3aiMzgniYkwHn0UM+KUXvBpIButLwlOuTK/MlnMX9LEKvUUtS/juot6HU0/tT+1
31bwskzSgS3WsAm6d61ZOpXVTWmy4YfTFxFxFEJmUAXSU9CpGZ/tKJSotFDmJ4ep
k/eKiwBwVekBO6pGaoAmdoO08fbl8VPkchPM8fDjVSEuN1P/ZM272XCdtosJmeWe
wg4cxolxoQfbj3glVP8yZx0RwtH2gpHC/Aa7ptcGFehFM44xSoZZnWxBztR34GjN
x70RoOBYA1SiSfxNxbMbR27GTVjj7j4QyU+J7WAdMpUEz+xDSHgf6ifrr6kEKV5k
C8sLyyLdSS/v9iT3fO04RgU6/IPqkDBWCqf/CRWrYSdebRXKMklVtr5I9t/xC9X4
U+6bmVVjjexO3v112CxAwuvj3AS2AItm4zIMAgsfrdmf0d1I/D32TO2znQNtMiUV
eO4yyGSD2O9DHi0GTLPJ+PM8+9NOQAFcg9OmgynbugFoXekF0ruZQfbhZ266uSmN
/jbv0JnzcjaYp2Id1SXKfbrI41nA9g5szDQhpRDSycmYYhryiiH3KICMkawbT9Rr
mAAaubeRnHH2YVk4xgd5gZ3d3gbYKlVJZm64JI/Uv0hiXq5nxvxnt26QmW8CeGPo
G1Vf1Frz5kKL7p+7i3oVISI4NtIVLocQQByX+2ePTMwadJQIaZmGSjwttJImWSmQ
6HSV1CK81OXanwKdgBV/v3o1WwWrC0Mpl7zc39XRMoRARIjThAz4Qkt75IgdvWAm
0JJVQVXuf3pbFfrmBO72eaoBaIXTaMTw0XWpLTSIkxkeM19KQS2P6bCwBgZU0fHU
c0Hh6E5rVbRL7Dx1gIKOWgss44zX4CSuYPvi19ztleqdpYRSnqhjtXzMTGnRsknA
b+qKe9FhOjwqOUZzngvqCJsxN1+8XNcBFVHehgwxgLqvifA0Qnld9IwG2EQ7hua4
cYHhBZcxu7ya2jzypGr2DzM1y0UPM/uFdTzL0qxkYo6C1ANe2tuVjmjNCMOBCkQY
rWhtsb+yzzUlqbN3SgNBdZeKlndYtV10u4sS1IwlYfXmTk6RHu8OOfSZg/KzkczV
9kxo0tsN6GWHVxDxn27za28DXnVzpllWAOxIuw5iRfSkN7HxDLsPDUkUB5vBjOV4
buNgZ601/4iN9TdthW/77GJJkAY1mpbLMR2bwvQ26MFSh6JaEhx9l6qT59TpgfZ3
sUG9SxFLeD88sngePVoOJoNZXkM9tFDCZz26J5w05BagzUdHZJcppI/adiZyLgSW
B2PLr1X6sUBBwfYJs9Y+NwVLgaXnZFKnTmn8AyqOstQl8bgLKjSnPuGh9vuSnD+5
wpaYuIg9C1a5XvD3WN3ldOi3/+PjYeHDuEm6xL/4IUHf/GC1s6SFFyQJ7GXyxETE
ymDNcIX4AfMxn+R7xz1+4qUX2iJoz4v//JaXrNqMgschBlJa5HmBk1ngXQTYHmrw
I5tpYjMkQaCloNTux+8saCOYlgq4srU27quhMJctmBsYnifC/KzsCFLkoNDMdPdd
CWoahBCOKt7LwKoSrBZavLNo1a05CDJQe14D6oHIqEMb+nFhbjrsZbV4gyvrz4E1
z9XWtXU72iRcPPiMd5tRHXMyXG5yjMksyidB/kR4Y2HtADSNv3nL5pencpM+5S55
MbCU7iV49NGv30T0Yt9hu5T0NdlshxYgh0vf8rOym/qjKLDysIFc0+40rh3LzuaD
mK/6DjnidrEA7BlD1ifYmBgAI+RWxq/zAfYeEHKbpE/R6j77wEwvJM25ubcAI2qs
gwFbw9k5Me4D2fjewmCSZLOp1IWSMoAB+l7aa1VPeFmOKotzG8oIML4rsJNCiCTF
0zeXh25dLgd2gCJLaB91PFYfTiZVya2l8eOAsjlXPrU16z/foldxIpEAqA/7t/xk
TVK2Hyv/I5tNHpMnungdcn1vWIwj6uT6IwBTUZ8Jk0ScuXQfHcZ/++ZR6A0+JZPd
uXJe+6PqozqZDkpfeNPAgriFs4IPdYUgYzbTx0EdJMqAmmgGTKUhshqPWMdc70HI
jAQYw5axoakPywhmK038VQ8Hvva0c2SuaTH2FXzIBdK4YQ4brgPGuPBh46XToVqh
Zl28VKqHCHCzb0E0++/+HrcqXb6Yd7B9jd9/J6sKjVg0YW7Oz8slyWd4V1Omr5Gb
NI1md3Jewfg3kLOhO3SYpY6k8VvR1mnfNHx9cws+Np62wUnkQglbW8z+uaC4hekw
2F+LbenV/JJC1eMimVmuSFK3ZCSDU9KXiSl8V2OvC5/pBAx5g+jIVsUPHW/9f6S1
OdkL/tHEUg9GpAFRcibjwAo0oXOJVWJ3noOJBnaCSBoa4J2phGc6K7n02OAztH49
1J4FBotCm77VxH3wHMNu6Kl8u/3cpzBpkckvRIq1Fx8W7URarnX2SH7UN7RyUOeA
5NA2oB1oU9eXB2FtbzccO1oKDQBUTbYs9yp/Ei66Ny3rYO/+nSvqzkJGiXnl8gDb
Bm32r5igINQXEC/ERI5WSI8QzuikCKb4rW5TmelKiP2OyBi99JDpCAVy2f9bfOsA
wODP2VcMNzYoxnrhGWN+Tm7xDB99NztGo+Xd5h3NGtx++1virIH3tjXHiKQGb3m7
d/TgVWnmzhbL+fv3ZwjIINRkI1xQYWgWc+Xqyx1k3nW17w+CBVbYeTrhbkFxdlX1
a12HPKlgi9AdJzXBQp8n8uU7q73SvED7BCX+OavKvhk9WnpX1sjYUwYbEaAp3Dpl
ZDqXu0Y6guqoiri9nz4J3f3jRKgYiz0dzBPLzH7sFaEm1nj6x/d1/XeNMySwC+sF
kUfgRDbbhfXNbTu3UIMAs3JCiz2eGk8z+sXaqeQOryCGfxf+h+3HA0+H0Wr2pAll
NI/Jpu6OAFNZWrhlJhNDRdP0z62kwFWetjmZnMCDvO97Lelj33MT7hlXiXz5kywN
dEb2fZle8BU8yNkVBk57gb/Xm2uz3SCFOG9l+7jFBdBl1N7PIosb/klrYZNndHMD
i920G2EJGCnL2qctfnIduK62Byyq0q2ZK/UVpBPEBSmWQpZtNkcebgqYrNfQC6fZ
sduIgBjZvZup0GbAiG/Fof74huGvRuhy8eAM+PgIIhhtMiFLhcV6hjKt0MRMZH+D
XIbFRdkbUG4fBgIYmOi6JYe+FsEkiEL7XFSbtMTxIvNPPR0NitsnvpPNaQaFyXH+
0xrTgWcZWMKdN3FkyKjEpcje/SU5IlQ5CUaNiA25zq0hbuEM5P8BpNjLd+y8fvQN
3tvnYO5CaSBuhi6CAlL+SZcr//jtX1GiGL6xY7Og13ZeFgj+kx3uZ7n859LXOlK4
zxJa5i0zOX+EzQICl95JN45Y4jgRkFLvO9pk53eHEbVhTU41hZkh1iz3c7DjdEWM
p0L/QP+nGujpFRTUYKOww8zj+Nx7ntY6qiOtw9OBlKNsak1NS5iNKcYSUPLNKvdU
7GCapm/OdDEMZMA8P6A9yr+K64Ygs93bgQaEgYkNCNq4/o4yKt0GosIX6mQ1HFDE
BP1YpB3sZsu8TqMhuCZ7HLSfPJ/8aM0qJfx0u0NWKArJFPbL51REfTBtwk29Cukb
d0s1DpsnW8+qQT2LFTnAFQZqaa+hCLCyfbxth07xtTzcnB8b59SVHcgQyQ8oya1Z
0uh61ATF+XHaBvl1s6as6SgVTFax2v37h/S1vcqTnvNLm2HDKlib7UPludyABzLh
3Ot22CKL+Y9e/BlF2NgT1P4A0v/l/rg6xgHhLM0IxJc3p4Mi47VxFG/70h9JS3WS
z3VA3REBnx1Vq1lEVTd+E41j3T4r+WT/6182kKEmWQqZ1Ze9fdJ7djoTdSG/iE/F
2CfPiUbSLpjee3ZnHWQq1u+7bjuRwFGoU8844Q87x3ZtXiyYqvbXf85rAOQqjCj/
4ffeKumwqKfOM6k65OsZyS/xfzt8vW3BnC/lNyhUuVilceJPIGVShsI5I2zdKeb5
vrszIvzR4kKRM7QKHmO8heCxLBgzBJhusdb9h03ApziqkkyQiJ4OZQSKTg0EI5iW
JRKDo4m9g7YZ6lex5iYgP1RO3chh2XRP8nvFgjesj1iv07v0sEtHeXz7Yn1gD0nx
/2hHaPpzwVL/Eat8g4iFyZpyaWkoLwRMytM2Zsa0qiKPvOtGzDUwxi2oyflaXgO7
pOJH4r7NU1ptLe4I/essibUsTbqrtJipv9rGY8FDXsRLFPXWLqMEdlz+pJ6UPKYt
DcJAGWOxleNkvwF44FdamoV9D9B5TVNM5giUb8Wu7kFeGa3i7GXxqYN7wprWh4SO
B9Pd6p+eQcw+sPWvBRFwjVAFWej7FmzFcaT6oi1hW0UYgVsyQ7VhD6JBQy5S3v5+
Bik2brBl8OvHGK0bnHn5d3y55gUd3NC5cYwOU+YBWVnZ/Q7YR/pOYOoVVPNU2upw
CzOMZh2ZgAwbLw8Y4fKC1gZDHwoFkP7gG93vPXEs3IB9frFGNVgnJQIuWCNa5Xah
YOWYW4j7uJ9BeFdHLYOAEkgyIUTsb6HoVmYZQtQvZeZ+BPXEcWAh7ksf++46GYGT
6DZYcXxvvwEXdPrHS+UGBnALgZMaZrunx80zzDHeJE8eIe66geBUWfOWTAMOST4l
l+IjNeM0+qt+66sngGjFWXgLasg6PsYAe294ZI09fIuflMkvrObQay74L3S+Yi7X
NhNq8d9Ofep+WW7XVgyGR2s4Y1H220Q7im+mg0RWctRCLrznPez4GYSn9tYANE1a
J46qj4VN9XHe+oQwi6M37smWO+MTxP3wUYFB4rbQh1pMNUlfz/bbXoYZtgr6oezt
5CtgxOKOPq88HQMzAio5gOhXFls0Acamgbb4RMXRZ1/gphtszNMKkZO0J2TAPogZ
1wXwVvD7SglbLf8fbsvt5YMnkKRyNzXeUkhBZsDGhiXmtzt8ScDQdM/8GnbXH63b
8J0alyBDNvrorMesihglh12ZOEf5y14QDyr0IkoqZkzUSTOYN+sxPZKKcmzMRTXe
kqWjS1JnQiCWW0dbs+zuGuTRPX86IUuv1dN1+GgjzNj/n+QOTyj70RZ+4atrGXUV
bqYChIRw1oNH2EctUsDtielEVAOdsDP6ujzsaddPbZtxgvWQKQMlJkWagswcqQet
KmJNYhSPMBm0QIQTwC45SK9HmAHCv61WfXP8rBIan0otWR99rhvewJ8QshWlYiUQ
FcBQmadDX+zjp7wvZrn1gAhM/pWD6WZl+FHjUuy09i6yOeQRfU2SVmrW3jkJDdhU
AtYczIN+cvCS4P7EUVrpSFvTI0DMydZuhh/9RXqm4BlaSjX33TRTc1SuzR+HJwbF
5b7hVDodGAC2YzOHlHLEjlLRnFPbwDL/8i/FihtRcT+RGHwyUwW3HB4Ii7VxTRxs
hBS21Z2YOASJaDVPQ0RVNeWfefatm09/7zNz6CMfMIR/hsQRLEMuzWtZ8HDu/iXq
TVwphVlA+LQ+aYXnnMgqlgrw9sQlkmxeG3cpL/0PXenoRftO83RD7GJO4d9hxUV2
/dPZs+e/pWq4eGmFRv0MPQRe73n1SjhiurE/mj3aL5eqhHFMr8So3sgmAZGLlv8U
f5jUyPfA3oMye72gM5eJInZGNhATI3leH+PFmB3bC9p53Cn9XtImuwvYQDxNRmpI
hbVaan0MY/Ko+53TIOQLzIFREXB2PN4G8C1mp64m1NvGlkkphxRK0cT5VXh/dWdW
V+OmcJpukWO1JNUaLCyR7VzkC1uoKF/KTD5NVUT2Vj1fkdJ2l+aFhBnJ2Fa0kYjz
WpP7u5EZ4kQKTiM8wkDSrKRd7Plmxd6NB8IRajLmjsmZna/ISatjQHOPADOV3g/W
bUuxxbK7Ry2mquFc9NJ+BJXyiSFE/MajwvIbIHRak/TfPFGXPbQsG9MSxuvLRAL1
KmWp7TiEK6/00qJ7EdposQ4VO4Lnm41EM9ddoGlgRTd8HsuLKpOzSqfL7phqmSl/
3eYf5oXGvFh2h0fylx5Q4zSf1uHOxj/BTZpYR0JFHOGkzheccll1J41h8hyvKU0x
B6s/9Zami8aQb5LCMyeGhx7kt6WDtGQCz2NUWQNq6Tc1K1n6/OJJUw+hQ+IJQwN8
HJjTGag/v9n6VXVfBPARQq8cVILSWfIt+B4Eu67tjB/dC5W2ZH6PJ0x+a0vGM9Ia
BQeM2CJZUI2j+FAwO57jE+GMs+HQykcDszs8SCBxk438PM3CJfOfpO1w6bld3LRA
a/KcuQmoNQUwW4sqeRI45VUca6N74Cjemmlx/VvyyvUuXerxpVQJJoLhcZus2Sqy
spy1XWHnXWkutIF0busmIXh7hoLWgftZMf5tn8W0IaTOB9OEiHc0YuBUdtb97pyC
4yBWz1abLLgqrpTUFjVow6RrH/CKhOH1kLj1UapXU2Ed2lJq4iJ5kj8rlSzGqO2P
fOlWn4bWQbThilLPreE8qzU7VJa2l9PvJQQUXQMcUQJdvmTpqpPl8btZ3A5JpqEC
3ngkCAJNCppefzzwErhPBHTHGuFsl7ThT8r4WuAX9FamgI5IV+H2txitKy2KZsUZ
6dYddx1j71Vgymsqgae+JwzL+9jYxnFuFrrd8KM3eh/3brz9yoc1zisH4FwmeHgo
6gtCD/YzScbK2WmxloNKA5lZeOH60Fm3I7qZ7sc7VR2L7CRIxR68diGyIB84m5wC
M5rGkY3IaRCGVl9UPaLHoy13Hn9+FYURRpaXC4pJqZJL7LCn5kfPwosOTP53Bgeb
sdG4yWK0TUkOFJ0NfbQUICVtB4f/7UfGquYWnbJiZqOSWX46PAGgmw06fhkW4ouy
T9oLwRfdaiiwWWxpTcipMtgxP64qho3kTlVOduIpkKhXb6eiejAbzVUys/11obOl
7o3AtX05H6pv/qT1fEh2S7zBXZVlvaFk+OJ10SFM4WdX+xvO9vUI2ujKLJslLM4w
vXlC5882U8vb82+bJm/ZoWZ8gLoKAbbaILCR9zpXgXTWI3xthWx5jGgl/AbycKJV
eXqSbZVDSa/t9/aEK0bjO+KKpr5C7q8FckIeeNdtH4i0eZhuhd+WDdFABTltjWUC
kDnIvwe4lF9YgEAU8unVxlX6P7NI+WfiQgQO980G4OMLPnp1hSROFe2C/5TRw+cX
9tpIMgWuuOSIBvieQ8i2tIywTygBsEH9+W4IYe04Fvj9KLXMp1+TQ+TLQa2wjW6u
Ig4XE2U7dyWM91JMqZdPSM75BHD9Wh7noFGBlWMzZcjD9zYh3sw/9F+1wpb4EVNm
C1LxiLLPH3/OKEHQtFcnTtIpgiNWxFdL7qF6dalfydlmy3qNggxbZitFchaMZds3
1k2f5F/nOARmrDHd0VVQMVEO/qXJMNWNGC0sQEI94XZxoAKhOMgP9A6F1O9qy6W6
H48cn3CDXGN2jMtq7iQGqopScx7qHuj1U5UfKJETxeQ8VdoAop6DKCOLfvZ/rLJc
ADK4onxkW5q6f6c13fTti2xzo0iG+UlKYujb4B8REvee+p6ol2y4MZejcgvVIF7+
`protect END_PROTECTED
