`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yX2c8r2uhQU+5vAPppkQVCEzt4oE9FqYcHjGbNaYOkXOfRxC81YoQvDuWwIjqTMZ
yBTWmWMMI/Bt4LNhwdi9iHJheAw7/OmIQeFdQ6PZngA3H+WOBs3lAmVs1YkGYhA3
dz07AePP32nzF7LzS9cIBPS/UfhfQ5+3vXfY0MaTEFP4ukg2LLckykWa/UjtcEN/
4rjoVAZZhR9dPpI3okO5vlXDNdQ53VaI6VKYNcbNISpLn+lggFoBwKj8JwBgXXRW
MbYi1F15djvmMnwXNr/72FD+byizXIW5jQhouHDZ2s8uBSSACgA0W19+SeshoQtq
rCLh4AtoA6xku5ikZWDN6HG7Qg6gWiyWvvcLvHScQkDl3R3xzVOxg98Z4ixCuYGP
DlIC2gnGDm8fArmSQcmCGukPamEJpd2OfyK3l3SJssO0HE2O+KNViH1a9DHhAr7W
`protect END_PROTECTED
