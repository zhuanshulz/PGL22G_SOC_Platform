`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zd10/0ZVFdtqLZsHYgI1h36Ckx8TWmM79yr7YtqlMrKzOkMgPWvgwQtcJ+fGwvw5
ORQUk4UagX9ovpsOJpdAkFAcjCUYjGwS51S1IEw3fcFlaF6LSe6Ku/cvI69vG8Pi
TMGuC7X743uB0ZrXk4PWhI+EDj5k0zfUXAJsCeezkAt4LP9C5j+BuLaAdDrqFW4m
nDLItFwV/W2LngsfGTR1XCQ2Ywi8ztOk/esidBeTb8dVedfjJtQ3cdAt+UeDRJ4f
aaembCD+/3Z68Q2oK6T+GFPmlZZwyOnt7SJeoOzJ8eiYhUat6tW7xW8k9+K1NQ8h
w574FYrbagVjdtwoaWp4MpVnaOP9APefTrR8Naph9JEcD270FBqM/NuyTANPhwTM
TqBAiWmR319FZAtCO2Nto/WMWflCnzhQJtbY6omQUUtUQALoXylFhst11A9aWs9l
sHpicryauomZjQZQCq3EgDPUQ3w9TsnQkSR/RrKBNhf2d9N0JC26OgYl/vnI7Xvb
dS2JzhbM1yUv1MmmDpXNJ18c/CdHDRzI+Wb3FZsHP19xFQYBEo/CpzxbXbr9N6nz
xB35MrSINAd+5ABLKibTyMxigt9QEFZJw+iGDzAn84uoAPqSH3ExYscii8lb6ohL
lzruWpkJZDEaSVuK/o05L24np8YepRioNThaN2LCpwUr9OjK4I2/ezt1w+rca0d8
A6mN7AhMyz9k/v7aizwEZqXgxH8Ak9rUfbaXQj0NiHlE/R8w575tkXZBwsnZ5lNR
wLN7pKnycwKaexNlv+GIFBIokO0Tb+CWJOfNbRJwmR1G599Mhknw/K7NHqDbXuw6
ObQSVglZxOqhHvIdNZnN8Ajp2pkSsM2GLm7PziTM1A+EthybseEeYTdUpeThkAfj
XviI9gL1D9bqxpSrE+2gFLcnC2D/StETQAaZ+AjrE8WoGsEIXT+NDEWMyeIddkCx
9IMjf3N+iJeo7EloU+L+Y06j6ABsviGrH5Dt+Mf059pcgaus9+ffndffDTvmhDlE
6POwtLUwqWNGr516thNhRmzngx0uNGcHq2NkQ2Wgig37AcTedSw4oRYGwq+esvjJ
0hMHWeNxXDIajUSvtU8QEC5po38RJgJQKi25luIMQjz1xozpYvajyJJvoVxWOTHH
v+eW3uGjOOMqWz+nNK76gPBOa1JMzQx09jNy2U2oKFYZlBnZthXGGyqNEDq15tTb
gbQozLuAd8kWVcIgPUGZW5bXvqNMcmOkzgd/G81gc/XSmtL5W/i1FDQhMjTg8tOR
r+fdC63JUhZBspRv7lJiOCcZkgpDXoeNCDrb/PkGySmvgyVaWrfe5AVZlmQK8+jd
nM18jhZccT02fH/IRPv9kcEHWG1z1IvGY7T27vPD8Oh7VNVUqbU2gNJRxPQX99bf
fwl5RTWTAzSE1eU+XXSH4iIVKJlrkEtUePXTCxBQxLdYQVkzFr3x0WXIuh9Aojcc
x50QvlGg4Sk55Gup2mVb0TsjXymI6Pmsmqq7/rhP3L34h4yU1D2brZIPAuIlAgBW
ExOZAbIbXY7BAdC3tPDfE3/1mSqwzsT0kdaWwbtEnF/pdKva/BX2uNUdKGOAu41t
PHQmIEweUxyxJ33Yf0NvzPfKFhMC1QAFGbRribkxZckDCjsfUfsnCS7/GBHotffP
9sRsESJSpiGapbfsTmTPIgUiFbY1jzPMm9AiOjJ90a0xMzRVeappP7RTR29JoPxs
grC9kq/G5YoUNK99Y0Cjh1++8/ZNVXlB/S0zjI0qMlhdgjc0hGVozWeBZRSt0XXv
M1Enu2HRbGAmNgy3SDqpNrDd1gj+dYlmCUSyS7T4sS30CiQX/gc/oVSKmNShHkyy
DvjofbQo5RLPNBIr3Hfqswkv9lT/vyv05QCQ5WUGTWPPRX3JOMUFo2PfsN61vJ8x
8GBZoTCgbQMyyW0LaqrkBUSzmNtQl4bt67FB37JoBRYzH1YUULP66mZKWXcsbbip
CdHO0Mfx7Vu1B7uyIpRAdnImWHJ8kH01IdQkXE4UVHdPVL0zpYgOAiPepGvqCyAn
3JBrn000PYyaa/R/gBwtni+2w80BbrY8TYu14Mdgd31d8IxSsl23382H3t4PBzi+
VJkJI41CNA1OfqpgLgMBrVmmlckgH8V6TdZC/84Ff647tRJivsY4LROiqNFUAxob
hg7C3YctwDCT9jgqKv7no75L5rHe42KgrlL5K+Q9JqmiTJUIncLuD5ptu3ddIbLz
Axy3ZgmpVKE+hSbVqJCVrxXYT2hTDX9KrYI6BE9WjimDri3mh48r/V+goDfYgutu
WqI5HAE95FF/nzuHZxCTNeFrKjSKbGlj9jdqBl+y8TwusBKENwZkXFWTBtNO+ADz
XNItW8Tuh3EdWkMjs4TVJYvhfmAMblGs77bnydwiA8aq4lVZJzcu8iHRs/XSTF5s
V4RNGJbjxKkp42JZCJ4+tlLV6LbEMubLl7tHaHU5GDXswJVl3uI14dJZECqXhJd6
f3Fu63zC2x5bJMSk3fRMPMHrNI8JRWU6wxzIiTbl95nIPWSpg039ulU6T4wee38n
JEUIBUKZ/W+4aZzJbxkpjVFsWOn77Jth2rbXPDaVIxwQj6zAXMcvfinz16RDQUQH
AziF92ZwRBZpGDeF/05byajDWheSF/c7vSoUmhOavjcJkzjDlGjTY7P0t749D6m7
N2GnVLwUVfNYXm+koi8ePXAKoq20gkI8V/j/6SSQYLuL0o343jFGHzZHmFPxatOX
e3SpM4qn6B3KC7CVLmTz8jpM58zZ5bk2Ot9gieSdxlL/RNvoFjddfyZtNqNZOiby
BQzGP1htOkHGHX75Ayf1SbSab9ny3rxuwvZfdEe3kwqa/3hbO7vifeOtD1Ck/Uhf
ZoabArKAbDdNg9xnhf0GY8GsiH5ATFsGxNbbkvWFVhhxa3Him6FLBJO8CxHroB9a
quHRvfRgE1Y7ekGyYBwI+Kq2vi4jP8YqsvzRfrbZpvoD7TGHGJMfnr0dMTDoez9d
NaVZGC2wQzQvLfvo092oOK/SIAZ+njmpznCpbOMxqbxPrss4zdLlHdmefY311WtM
QisxqMEdthyaayAirxQMO6vWgABX1ofGQ2K7MPAinPU/47xRI8vIIblT73ijbTlZ
+kiapH88wDgrq4GT7+lmkWwaHnLLUEora3XqVnqqV5uDtHFwDIr2BAd4FfmhRVSL
wf7ZiHv37U2V2HWxFEQ5IfVy8podP4beN95eSULYhKBVKzdAGA8Jj4iiEdtMTxy8
XaExf+rnHiI97o+jCM4Lt3rdXD1pGQ2KW8Ng9Dq/d5nqguYF1T4U1QyerWL2nkOM
IDyYl3mjL7vgJ7wzjA8ItLMoDQhWx2d+AhAyZKyLlfw71FcqHpiCkR+KM0WUR6G/
rAX1DeWcwLiLumkTPFcNDXGXEa1KaI1G2WFqxfJBGgRv+RZhZjt4U0k7t74iHmB6
hk26E+1/VtecwHK9HQ36qf1bXzjvH5UIvYIdVQ4GQO/dQJKIMYXseB03e2xIda3D
oHxJDapwyMBLVEatQa0yVr0IhPHp+yO9pOI1EAGOar+wz/TocVvp7iXCHHaJVeOR
g7n/k+DhilZyIO1B1qkDaxm1BCFVp/kcqS4lAosvmNYjTccnTRbQSkbHDhnEdyen
S4Ji02dCWXQCnw9Agk7Ud57r5t3U1ImYRyys9FIgl49D4o/Y47C9XlOWZphXloSr
b0Ozi6glYJy8OgyMx5wNfY0Tc0Zu8rSEIn0lC8jEu9inoiWnN4ISsCxMnDo6WHOT
HwHYfXhM2hg1UlhVvLnhonfdL2zoJSGg+mu65YZW4OHXnHXuhh/6yFf7Rt9w4thN
j1DsLb9uQgXh35BM31avWefHmnJwA3tGzi+WHDhnHKP0SXHwqeobHULScxNUhkZE
9R8lh1BrsVhqpNrhtBtmRRy1d+H6DEVndVo2QqcuRh3I8gwBvOVJQOG3mlCH2QcU
W7KpJF0E+WeBfHpmoPJFVD3KSH1TvoyWCh9MGjIyUiKZjGUUem9evdScQPuJKl9/
fo3sCVgAakOIrwUZqOclcauJWwTLk9pPfuslgu5a7jE=
`protect END_PROTECTED
