`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbqcHRkegFX8NQNpElOfMMv5RKMQmYyh4Pil6ZcHyd7EdTnkCwy0fDzTXonKSnnV
jBaC8CUvDC2BETnGy8PEDd+WP+aT86ZID9oxQXpvWNCNt6umucMfejeGnoTqLaU8
GTNqqgJave18XFtAbwobzZ+J4uLfI08Yk27yynN7pzZ+Z0CHoAW0tzowxeHgOIGo
eVu11qb7zUsC5IQdD5V41nzb16GT192UNGQ5HU8Naj+3cgNNhNR/3rZiHYDflAlp
cM0xnBMghEQ9dUAXQrq3kXk2bC7Z+XPGxc6N6Z3Nbf3AWzLXJQczfZ3y64Or6EXh
FHtV3RSUht214lOrBE/wpMmmJAJDKJNSc9cGu9mYa+TWA2qsd3/G89TQ6mMDlgjC
nHs/cZ3dw7tkdmJUP68A7m6uaF/XqRKeHojxW+EgYtCh3b4srBQMSL7mWAoHJtX2
/h3pLf5jKdvZnWPLJeG0Zvr978bBWGelFMKPM5C0A+z6UQoPnF9L5bH+gNxFhZn4
UcoiYFs3CsGPaFWqTkC8GRL8W+ZGHNCnU1gxyLzldI2Amo7IYvjiUFejFXsw/uym
IZnGe5/UFHQtpZOO0bnk5JoTXSwdDccFc24O/UGPfhlm3XAZRUmuOnMwOutdG856
wQ9hW0UyCsGiIMSwL9p+4Jxhux54lFHxZwL//T9KFoPaTAAEPpahKn/C/yZWhwWL
t4Mn3eW9Avjsx4aCYI8lAzrsWM6YyoI/BA/z5hbtdxM1WAPPf7niCX/+qES6JAZb
n1OujJkpMBN2vTGCkbk6y6zGOUG9L2wnqeQ3Ffj8y4I5zrcRYiM/Vd5JEmfvMbbP
cjDsHueDf3oEcfPcBSbzwf6aom+QraFmOB62Y33hfmgMyv2ZPOfMqxVtS0XE5AoN
AKiRmiuVHr9TfsWQgkNFbZfbQoIWC4HxjWV0oFyDjHIaOd0CQ2qyPDKRmbrn1G/G
tkI101YMtDc6UFvK3OWNOYn2Y4tP+3+ayg3tiutewhwW6xwMblq7rDzL9hS5+yY3
/TCUrWy+KBQwhO7BgjVBRlnfQJwcnWb8/Hed1RuoI2965lb0ybK+20dYFoA78pLl
a3strXjm/hh5l6BAVJCnH0pPyaeQj3Yx58aK6pqQvZot1dRclL8V8zVVZ+yzo5ve
6g1DuyKuO19yUcbB5TWqIhtzfE4fHVwMS2FoCuOcGIeQ35cmVYbg2UR89Cq18fw1
+bg8/cYykm1K+tqwVIDtvV0pfiuh2dxO7NSJEVrGgyRf8RWM/tbh+uX9MlBUROQb
BCUdcdnDa11TVcwMXCSgrnTNRTzheA4+Yz9oX1jOzUd78CMIOmBg2XMQ4My799Fg
9tzVUFofTtAyTMi3jmPw2aToCwUJzFTIEMG6+FRe4xjRZ9ma0IaVd8Kb9WzhfOPu
laDwgavFy/w7vLFolIlQiHyir/WsPtXBMgCxyg0DCCPsjWgMWp0HxXbzZ00Kmy3W
QN7J3CPlbqaJwVhgVKBnEka9Vw/C8+syOVdW/7dFgTqS0qeOBwYZL2uTGTUKrx7P
0N/mijSzSkN3gwYsPYfGBPJM3/jhJyVpXOqkgDpjGD0DX0tU6mRW8L3HRLd7phVP
Xkz5omCQWt9PObfrFI9BCQpxMbTo/quzWROp6B/EEUsakoZs7fMNMSNLVpFwNLDT
bYKcYb24ukNbXASZv6iuu7Frs8JuUpx+9ilFS/8+NL5lI1q4LHUVwDwYC5hLxoDU
r6aCfy/Ow0VtaHdMlk1j/Rv5bDiweOjPXEfYutcRPmzszkC180ILmytDyEOL3Yzq
DWmcqWFIapoTZZMHgYfom5YMul65YwM9wK9UCVNMothh0G/KgfgjXKb0/2uXU1GR
glLoBLxE5zFz6y5Zhtv+xTW2SpLj3+EBFsnPQDCqmlKjfIIY1E9XxGNF4n0T4+v8
tOF0l9zy1082zzRalAhIlW/nxgudWzQzW6kSoYAd+OXHS9ukxoCzx5YgAds0VWDK
LauIjBraSCXWb8nEAo17AyEuOkRGqvPqvrdqZcetyExxlTbadF4Q0qkpl0zicEd2
e4SF6hF0dyi2wZFTcfYPKO9NUSyjbu0PHzvt3h79RtFBZLowKACyLGBkbSQxsBcO
6RceF+h4u1nWf167bvjXNmTLou5Y9SZU6CO7SKSzGnmUqr8phGJFS2RiNN4bALXp
ZzYr8a1Nn9hk85Db+hx0mXAMPLjfD2s3ME+CF7ajsGwkCBsN3WX8tzeLTMVYh1vU
5wGmGM7smjQLiq9OusX3gRg2IhFpxNyYR7hEgKGuWeW3KV+zr5xkAOwCCaAJ4+OG
41WBJ7iTsbd9STtSMixRFVpyaqBRDdGumM+9zgj9KwZVtsQJxXprnTTob5VuPj4P
PXBMK0hOOYRDxXf1EHaD3DGe0hyRMuwf0J4Kg5J15rk87YzkHtsf7Q7y+5sXNh/R
27r8W/u00zzZii+rQS9RqDeeZTpBx2ZFkPtnRUHFOfZPkGYr/KOmma/qf4FcBjPb
prmK2h0nDbHbRdQZaJaqtv18FnwN1I+Bbm03DRrbjTFR0gsCmPsGW35HpoHqaib7
ivCgnEdslk9QO2tHRKsMcDZ1EHPn3FO/U4VSw+ypSoR0m9A2jYZpW3GTzFW3UH+z
P8jvE2YDhTP50OuDpeR5gVk9Q0Rr2G32upXNJHiSMEeh+QZ9+xqbVKD/XBYld71n
758o56a7YwyZTq+NLume+DfVi8ArjI0+mS1esRfLR/e/MGLP/C0xBmM32CToLFKd
DzTrw5iul/RjN8ig4Bp0+7EY3es7bzSCaRR9h/eNkwMJzD0my6qXvGJ2iFcpAt3Z
FJeMHgoCT0+bm7WHK2G0Gu/cgcw5SGdn7ueV5LQ2jkOrEjLIgLKbCp8wVkanVwW2
TxZKmJxAhXSUvjejlQvIw/AQcMCNrQFkwlsn5lezHJvHFmgkKyvvXZqVvMlHhbM4
cwfGcb8btzTAnD3M09UpdnVFZV9fBgVmP7bMZMpr1keLN/lZrYLkNc2SR8mbDp50
fbqDLWJ7o9R9HTy+1m1+B/o5AOUjt+XLHWuM8jo/vB7DlXXx6yOIyLL+4LbgBhpw
xt7moGAcZU1zHLytcQQrR4YQM89otIU0sx9oGJTff361z0OaLiW6Nf49O+9HUfVB
q/rhZf/SOynlrG/1VYOiBLcUzMN+3auwio3O0bd1A6juYNllL3Mjq54AwGfv9cHp
FHdm2OWNOjvT+1UYRxY5XcesZ+ZRoSr+oOlFV8muqxm+sW6qY7Fhg0dGEDBxoO/p
yELnUg4pEoQN/xO2U/fea6M47RAFzkbIErpSUT/jHRx+iT4BXYSeXCaZdjjMsFDi
TWg4OxoiqAkKvnroQXs8OnVTVIHDBX8RJtDOoqjItiMbm+w894QGxAB0PvumtzKc
RoOPI0mo19SUZDfusRjQqutt0f8skNVf0v2dtPxkR+i8JmgOyCvnSw1lh6AhpsED
QNCKCzuarfgBK+k8YANLG5zSr5Cb8xfE/gjNl6A0ZwA04AcihBa8WUm53RmVPVOd
s7b6DleGbIfMINoi+pvGCpWY8hii1P7Wjwdt27mRoL+TA4spDgN4lMapME3+CLQn
oU8pRcQbrq16oJ775bABmCzWbhZ8I41sk8idxZSKNUAnCAKT0Jx7JfGOoH0bb+4Z
k8M2gnq7IpM3lw2kM+ukcpn0nogf2skwHj/MEgGrx+x0BhraPJucs3gnchBBwOdc
V19vQlj0KAiaTS1NuWSey7I3Y3/f+w+bcxHMS0HVdBCOAJvd2zpFymFekXg10T2S
xkltWQ83GozLDKsVvCKJWELaBDVtFNL5N4gCIZP1yXQkAca8/s8ag83ILha4im/4
8/L1YQdqG1r7VLwaH2ylM76kS/aHiWboKMZ2QpQRJTkAoCtz0PZy1+kIhfhBhZ3T
3iBWOmEs3IyYHOGqQTD0GJWMa9OROpjhcd4lyWdyad7TZlWqIdWJwjHMALYBcL6k
Ppk10+lnt4yr4opTdJzXiDUD/SxRdd0Wj+GKgdNTFrMiCR3jXuHRxyGhjoo/XM0t
xrIsVZOmbyQxMS9yk+UBJgGWwhDM3Kim4X7Yj9jBR8I9KC7Gi4T+s4CIegZQUamb
RifRREQGq6GVlwxExv17h5CmbuyQQQrRRx3P7KzIAADOcv1qtyde16oEDQ/ieaJi
Wshxg06x8Y8cSNn0LQzGktwHzFopP++qkkiwhbbqF3NQXpwbKqfxb2a33Ov+OKbC
ulBaR6CGIChm55RtqxF+L0PCNi0IGjmYD4Xt1ONzrkNcg4TlEqJhB5fubkQRNXli
r/KWH8tiR4y+IeQf9TFP3pyCXCcMXMPX0K6gUhN9/wxPcxgprUYTeUjuw/jsPjN+
175vrEjajrfPI1gfO+xaeK3anzh8fpT5udEUB3iRabqeVtdRx6xpPYSuIUR5djV3
pAN62rBF3bj/Q+c+YXumiZuHYFXQJlcNlq8g3y3ZcJSmEszlPKNjl05rFfpVwJuy
GMe0gp9V3G+tV7c9Yg6/xX5AtdNCQ8z5jByHExwTTWd2GYNe7mFv9c90HZuSdzaX
huxb2+sfOjc6ybd9WSnWtDSqZEicn4k0rjuXtvbcEofGCZb/PFdCONpCKQvcQwii
8algHhDc/JlId0VqtDxmdJS5a7eJvay6xhQKLMmohLT7TSzVmEe0nxysi2Anidln
NbGA5gLJQ7/hWdZWN5STRR9p2I95bb2c6tRym1CWzJs4/ZrsgKU0sw0BXZ4VHyQi
vL/aGrC43Y4cvY3+7gSnyw==
`protect END_PROTECTED
