`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NPjNjzLJlRjijxwb6lZETj2IvoSEGuafoxgqdmL1xTCvXJKNH8aTQM4yAG8kHqZK
tIdV8SU5ZkPBkNAcjrsHlTcXnjY3kBnPqt6zUUuv8lbzIU5DRpW5UqGaoNITnKU6
2O/fjY90u4ixphaB40mRHhtNGcJu5g3Zi8lAAfS8NyUzjBQaqFtt2jUyMGGrrR2H
2PjJ2OwwgZ4tNeZfOfva+vbgXkSk6DBRJNv6HyjBOEF7Ma2EHgARaevJiF/tik/c
XMpeseMTBL748z+U/NDBchfP/pMHY03Fp6mDSzAiWZrYmP6szV7iK7NbZfOAO01G
PLpgAHuHeHfZ2W93Mxk7O2dVR8yw4fesGntG9/V39ahyOkwSyuc1Lr+Scfolls8A
p4rq/i0Ds+FtahKi3vkO1irlZfJMTs7DQ77Yu+12TY7jwnbiTsWvEWx+jW98TIjV
pd/3S31w1gGjOLBYJmfquhukOuKvHUp6vTaCG5lxmTPNuF3W5vNiNGLLBbWsz66v
s3X3SHKNO/G7TkdoluAydBcXlWYQy7raBC/35aDdK27GBJXz71vvZvjyDWHDJ9VN
vdwKkWwypPatymkOeF81JrrlkHmHSP/PxM3RDuj9l1A=
`protect END_PROTECTED
