`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUyeqoa6TV38kNraITmuiFMklvqMcr0PcNBX5u7OvdoIb+I+41FuRvsbC6QzVwBx
TX7kD/CQ+CFltqzj6tlgZQubhG/PbnjoobekvGKWbxV50gdUBK/93cDBPMpgTZ10
ZrWbYkIDHWn2sPyeelvo9dLO4Q2m024ADmeuKIpDL55cqQi/AVnfA0IbvE/lSU67
RV3eKjDw6ENNzmVYRgebm7F0PhclqtXqvUkapsILxm+/FALajl4J+YN8c/oIp+7a
HxlbMg3VJAkHmf1E4NAMLO56UQ3T/gmwMsTZRJyJnzYJQeCOLq28Qm9HEgIrKQdP
5itOJ1AMJ+P/jDORee9oyLBhp/R0fssOQbY8FchGuyQYg8tHqfG07oQj299kWCRE
Me1a02EUaPWphwIhDh+np3L8Ro4dUHfRx8Ydg75c/SbfX2rZV+fn0nkGp+NVk0Lo
2m3YlfNObGFdqovYnn2DwrcumgXBRfFHye3O3ftBwtZFwiYeTQ02/3XJtbLw4p4A
WYgj5fZzGC6I3XTiYUB0+jGlnclQgiFJuHXIIWRrcLhf6/LlMO7kg/VJ6KJ0hjmZ
Y7e/8kkP9YUz1xQWp+AEydv61hGwvdYYNixtMSzexglI7eTY8EBM1hBxZ6MSAs2/
6hlHWxBjiUq2TElKFeDzBRewDT4Vxv/iK+ikL21Dbhm8TkiBABiccqvwEEYePS9r
WwHKvFgaudqsuQiIDQaJbscolMaGDIIN2KxvuqbuD3MmVYs+mKpUWHizLHX1iX5y
prn/3wQ6MJW6x0nzUfgG7YUTUJ50Zf8ENfAyBKaAdG+2YR87C0rdUYSIVSXzxmnD
iJg18PrvnyoM4xGq7me8kJ2WL1GBV1UyGjb0w3EGiBqdbeEuAeplxN8UAPtuTsjF
X0pTbzxuxNm1Gi8gigwBGxRUrevIpgb8JymzGVaeulRcP5P5W9M1BCyx3mY1fR+F
g03pXAO11BeYQqOh+r08g5b+f14rizHxn0652GS5eF7Vto+OzaDyECjPFF1j7F9Q
ZoR2lGF9ruzCm5OUndHSNt6EvxW7I+zGuQAc3ywgBR6AWTybbL9Q1ywoKzku4Yhv
TQsYGKx39/I75Nwlkb+OjjjcUiSXKujJQ9OiCe5E9zN2K2jl26QUTuvpECUBKa1w
afp+FSvDX0Zx1BLq3pBuo7nxTrlOh3kMr6tkS1RVRrX/ElezICmF94+kCrCa80Ph
SOjo5lV5YnRZgCxeXS5vI5cABsml7XmsDKtkRdzddofIh6+fxhZr+wlmIa5dHZhy
IQ0rG9qDq1mPoulaqsodPUVb6A3FAIGl5OXuacMErM2Hmdh+FYAp/Xu1TlzI6TKC
EtGiIlBqiobYMSJ8xilLgnfPiNwddjzP4fn+m1CCp4mY1jeHgI1c42x5ranfTBom
NcYCzWerZbavKXZuszbbxkFT92Tb2HdGWSLbeAHohsg7tmLar6vcM/jZFSGHHnsy
T281JmuDIZFO5NQ6W7YAV1UGQJsL4oCFHYxRjw8pweKgmtT/lrRZXi+/jNMKrMl2
LfNkB6XopXhZcLy01UqSzeCvD4VKuaZeWOBeuN4zLSSXAGiCyqLlQETpUbj6Fsg2
d4pgBDSr4/rKkdwom5ozFKpuw0lYi0k0qX+FAwEqRtEmLxcMWR2xECfZBAK4gR2G
orFg7hYTUKPHTmLdhdNj6VV9YPqLDQJO4Bvq3+sLmmB/aebM30HQO6BRLgCp0Tn5
V5WWnjD2EvxMyPaIIz1PvhOM9gA6eFJX6SGZSwAvpVgxmmhoeAG/1HhcrDOJ0y9/
vdfZN9HIRZDthmVwDS2AEiFFohC1EmBwmS+3lWc4vzr2z740PCp9M9ifCVmMpVrE
l/tlyx8kIafiTnQHLv03pzT82noGp8G3fC/1U3nqmI/px4LqnR7V562158l/KMif
ACQmECZOYd12N8fQWMDl43ooX0mxUq7XtF6OzZUdtlsMMr/qWNEPmnDRiDfoCgqB
vXJ/X/8FaZFF/ZPIWmztQoiuiJ9icSg7wfG5KETq93HXOOZzNpZsKk22Fk6+Z4b9
MU56lUx26Ewuyc9gBQXberyB68e0RN5/pJb5sChVojqoPboiuSOjbs77oo6uFgIN
aqYbUUBcSM+E/d/kIBvjjspOhD8MYCpVTJKVpj3ElgZMlHUbA+5eNIqr7feaGewR
tdvhyx3kVaYYJdOEDpxuir7HUUMB/KOeCAILhQnEm3UUTdHjdN7kxTTkTlQcZjTu
qRsMDKVUwQv2e1jBcxjlyfvqxMIkCpOj/hFIqYWXtylc+kpxt6pIJy1qWjZ1zrss
diNDM4ukKKnD7HlUV0XjaBQxSVU5+honomUbCeCZaJMGp0ztCRz6TV6iNiduKhXg
qbxf0+JlV8lsv3RKqyrza6wYbJDgKPKRZGB1sXBjk6giUSJLv3z1nk04Rfs53llD
eCHeU9S1YtMPm5MgsRun7YP8Aq8ZubFkL+F2iIa5Hk9iJWVjhJmBFViJ5lx1scJC
VGGZEk6KruEPADSxnc0ctowN9QpDCXiWc+bgtLIpFu4BmCnURVF/mEBLRw0yJPFn
rSV/CH2IGs6/ZZy+MsluA5bowIu+xIo9joilSpugc4TXnX6SHjk/Bo+vYkA1sLoX
KPoRzsEGl0BCu98gxuQkG2P6yvuJ/seE2Gcw0JSWZDVZzsQMdnAHcC0Ju1VKYFxW
1kKoDLD+TTWveNzmMoo/29PzbPvda94qeRBgM8OdCKN3ThPlTAn9kf9EMQITpIs7
QerbaeXdyFGIMhVUcX9iey3eyBHwif41zbVPWrrOLHU/ReA+D+TokhrNruSdS056
4iGQb08vgf3NeYjUj1QGdZ5qbuhePMCSrXHTJGX5uAp/QznuQW7nklrQ9pX9vlZn
6oc+GXSO86PEnvqJfJvLZS3MsbdC/Isr2c3q3nWpuKmBzVrAbLiV0TZ0moP9fm/o
C3xvif0tRheE76T5y+CYQ/oBWe8clKZ+25F1wbZEwSiONKeeCr7UnvHuH3oR+GQv
FrSSuAOzFqVR53JNj6w4PTSdRjPiEgG4wi5aywG9HPlj1ymWIrvKuR9B0tmRHjXL
/QTTcmmFQ1NOJAT98mqZEbgWuoiA+91bgFv/nDU8UKI1pRNrhMpgcoyWlfSQ4zZQ
TguZOfaBAStlhdrX8W2DBfEE5aSJunpjV2bDnh8kHsQ3ln4W3ACkbw7KLpR/rdzx
ce/ofeqzkID+VEI++xjYRPDxedlYqtJlepoW/7K7qM7X9AkSFyOL1Icur0V0zgJ5
wHJ3js762SxA2IBwSUE08/mq3Sy4DhHCDBMuE1g1/ooAix825xuA9AYtxuOWJCnO
g+cgP+NGwVbdXpOmc15oPdfQ5PdvE4fp0jnpry3pVMufoS9MU/ITskA3kEzI7ksM
Nlwt0ErDtDaeEcdphspWr9+1FoyQcKnKs4aNqoHV1q2GyeJGRhb7ojN47g6E4TAE
q/Q9sURYsup5Ne3QVXW4yTnenVH3LKfwgmYrX8IdKmW4HekYaM9u+zl/Oo+XiyKj
RFltRAjDsri1gFmuQjT3ElXNkzZrzS7GN3xt73YL+aDx17l6trjBgK59hE1pRJG8
LL99dKoZewpiVtvYWvXUeIiEmYM5HTzaGMAnOf7JGpuRvZ8FCHsRXOFxJZgt1Q57
NaEvZihdCu+0Vr34ABptjsryxaQTeyWrxBwCXvYsI7PVSVJhKY+rEl38XjlD0jcA
tUb4iEstdJTT25dVUFtJBNCAJe3chb5mGvSL4bSPVIynAKf1lAjK4HkB1daspUjH
e3TN0k/pj0yle7nwPM4w/KkpyaKaq5nqRPIZ/2q8V3OX1JcqTaxbBp74qhRbd30W
wihvFVeUtKOUK9NZXFkpin/BwdLxwh4iq/xLAPHhMYdWIS1wCeUs7SlSPt7M5kR7
xVAtEwWx4o2wYqByjUIT8gTU40WWRljMvSoZazDcYrdYlxyrQeklvClTmTiHT2z6
o10OC0McC8C3SrIGE4BuP5XDOoo+sx9dyiHqiSHkSc/kvjUNQUD/OF5jQx0LhrYK
1i41i2JFJHUFL38L5qdnBr2Ew4RL4woFfjbIswucTsEPT70dk2xViaA8AG5OGtsS
B6YLheHsx+3iuNIcKIiPft+Dsg/2wL3ieN0y6zs4TmaPc7hrLhPabK29if6Fr6Rk
dTUvWvRsv9qY0VHHEFWWDTQRhHE/lAnwC42I3JOpYVv4Oyl/JOeFMkPr8HWxlAPF
oBqtg5DYSdn/nIlSCCayC2GTzbJJnhp9cs9j62y41Ip3w9Uy/FjHUqHcmflJP912
H9H9jh2D/QwflQYeYvmb3AJwoGKGzuwGT7/rBeY6VUqA5Ai4rn7/igBtRVeagN3X
oov7/6qGJxpzRFfOz5l5qOVkVUKcY7IdYaEGl7jWfNDDtxeSlzCwYaMCtJGrVeOp
G9dBVRSfQFNpuPLNJSAm29fKuTyXHUX2ZWW/M8L/r6dNBTjUjCuO8B+v7ZHH1q/z
M2pM4YXWMVsGFyHFv9ezEbTZFtVFNbugJMMkUgUj+M2kVmVAtgeT5pfL0JI0oIAZ
0601+1BZJSmIPyYDEbBtRqGAQYlRA/m51ZwLbBVsMwJP8cOOhhGf9sigUMXSFs1m
CB8p5hqEeeVL9ijHCrwTNdWA9LEdNvM5blFNm4wfRTZ1uHml+3BMDZ9u1ACRX9+Z
LNKB7LC58YHwR7gl5BNiYTv3KBUYO3FcOJM7PJkg915+j+0DSDrSREXu6pYs/fgA
gAnvDlQcTdUVm806raikELnjxSw3It4ThDErj7ml5aJXWWv24VPOaxarO6n2HZDy
+dOOr6JX6psnGUMTir/0NOH2ptrf4zgAKen1+FJXo2A7uNA2H5RisghgHBp1oXjq
unG5gYmhppPK8nLpfdmSZx1VoVB+bC51rKFeWC3B9EjVj2M/n3v06wnqeuEYnVMS
iLCPaaB95kBYxv7C2qknggyWjvhS9IkyR99FRU847ABzgGXaZOAR9azKT46Ai79G
MPVvj9ObFgxPS2Es60oXsEzv00iSmSR9GLuHxOHMETbqYUHuV4Vq0N61dWa8FOYv
x7emgk1o+4OGWUmtSKXgCaA2kQRhqw5Y6e9W2OJq5K2Y+3MARPUV/WTPFkEs1s2+
otQQGDZU/aQOrWe+2nshK6Vhwvex9vyumSwugMn4MvpZKkYUktazUxwpgCLbnluL
s+yHLgibSVx6nPaQgT1hyNTUCt7HeAPl5Ra3qt8rR+wf0DaS1i3In8XKhsS6kZer
pq64Wi6K2wr4mlSaMVUg/iv30t2+HJvYmwTQClJnGIjYW1sPDtnWv6aXPUzUFTKT
FX8hq8SYd+EvD7+By496ZVw0FskBiBqI8lilh2si9Ux0TAPqgfMVts6aUd+QonRR
mVRlIJryxHhUXqkM5il3WhDjpOXpWvjBUvD8//W5LrBEiZfOx0gzDZ8gdVVFYO72
U/Rp08nNh746GOINgE4XPQi59E4NPqW2cTSB2xf8DzrgIXRillw3UPPQh7Hhfua3
JUXt7a+ORcUFZeRjUbJWlekTv5wo2aK+nx38apjS5YHD94JOpOaJOdoMcChoY+3h
SSEN9rNelQvsl/8ykO0SBkcfTAxpXdDUqKPeiB5uHTgPiohzxDeDyiCu3FpPWjjA
L4zamNp5SBjvXTJdhRuinPN+YTvsWvh4N9pWBqe8XHFpRKvKxMMk5tw68c2FqUH3
DkF5Ygfn+UdteSeelLJrhtkuMwb6YZfIvGB+zSzmfgvjemliV/2cOQe16C4eLYWk
TZWVEa6eElo9/Ev2RlY744Y4JwVDsHt4pzQYERBgKCP+p7XHdU1+xH+9q9kMWhtJ
ud537FUcmLW1dqg1XXX2XoQMgc+Bsrz+j1EcoPeBRLDfOxZZk7ucXZPz04ksUen8
qzZm4kyWuIOcDbfvsldQzcnvyg3UPT8Wo7BH4InhVNuyhS9jswzwMts2QtpFOlTE
n6ECsPGmOSwqiu4RVR9luZRR2wz96U6iNk+PsCWVXVWG4BBKEs9/3nHiSSkXxpEW
9nTBZNqsAjaCc7XHXoDKUXEVASoESWEWiaXS7VX3WAtY8FO4kMUZqhEWwhCPgt7/
+aPVxksxty1DE9XBSp65m9rOx8udvDklzfFLmVWOz4uoRR9FLquzuFmg6GsvRNIl
lF0aKuNBoBHG3iUhO3zQG2tXE/bEhHlzhim/Y7gOTcfYCRgu6JFEILoqyLFnQ9J8
HH/z0mHr8MCuecLCS74a0hY1iT79HzUXAg1p6WYv5xs6lI6ygTrTK3arQ6Yy/SF4
JwJlYIC0bIkqoolmeW60QjFQk0rVx+GUAPoVUR4Py5XcvgOVUrZRTmT1gMAUUpmN
JG8CILtZVr0Upf92LIWFs2fCjFYCTjgwGkN2wTqWzDXBNvZhOog/dIC4OwsEpKVr
sj4OtLVCCpEhrvqx23FnTuCtMpp6w6mhiqeerTnFEUx+WFZxR5SKk6JNtinfAV3z
wX6oUYZ/Hhc+SXuPGiKNskt/FtvH02hqRbUHbADMJTWWiU2en0tPKGbJKa7dTui4
6OpNZT8LKXjYyiVeaJje6wnbbbK5HAO1m/pgOQ+a1n/IYqjU0oXdDJSs78XqT3Qp
SWWVvAU+3R1q9EFXnRhmwgPtqAnLaKR9qdmH3VYKN0dQ/VvFvfb4ME8CD+rQd7V/
ORAJ3UqqPtxPieWfLsTWoNwJe9S+9mN8Mich3VQe886We8UVOYGvUHQ045Rfv75d
hpk1CZ4NfQzo+P1Bw8NpaEhNHyPqDFtPqMJDb2qsBw5BlRqwPqKVP9jsuYQAmO9/
d19hPEiJ4XH79CX72nIFmFjo6d7U1M8BLvlPLDIcqK1tKnOEvHaqj4uNEBb+IUkj
g5r4SR3atrt4Lb3/y/nurFz5yQTAtidmQO9KZbf3f9MA1x6FGmo9rZ5ySDiQhdh7
DrdT3Hnc/ynQf7jyUtwhOdvWFTR9Pza+ei9QOg4XglM/s4lhHF+zUKrUbC5hkuI6
+hiXtWt//8ewgbIkxLvy8GuPYjJekJO6h/smoovTuySaFSluNtP3SD9mIZGmZsWh
FLo3op/HFU4kbKYo0RHhf0wOHAyxVIZVTRMcvPHmslTw/1vf1wMB/Qb+UJQHhgZR
z2u3RHs130/BurUeaPHSeXYS6hwT6tYH2A8eGgGZeSUfl5wOTJF0bOtOpGuqc213
hpI5cU4HQJiHYlR7PsZS0C6FhDm4TwX8oAd/IwKWrZ3iBS1DKoMybV7IbGBjG1mp
H1OENm5gg4q9v0zIb7XUYAq++OJJxZcGPZrhFS0QOcOP1KtAmcUMbj0C+36Cvuk6
2E7fT94jmGkijLj6L1LD3ARpNdAfz7VMB7ECVmG7xDpPlW7x17TfvpKK+DMja+CE
X0d3qaJOXtaJwUIhDK2hbZwiQ2dh3h6Rzx8p+YxTrH11E9Wuhuz09hbG3vpD50q8
YxqkUN2OSVUKl9VUdL8Xq4taymQJZYrOmqRYSdALgQhqdFu2KzmmwWcREV+UIZn7
gm4Hj05t+GZoqZJ0hIYu6SlO4Y+6DzH2QHJ43UP9BiUoHM7L5iPfPSjWeRJqxqp5
xh4H7PgRsQHQwPes1vH7Dynnexqmv6IUW//NgpR1pK09SVTmuBe/TlPGvc3n2WLw
trB5GfcO2H1mvJbYzkmSOWZB8aLFte+i0mJfJgd0g2PTiXIC9xWheDKX8TeXOc1c
klthZ6EuBJbmB5kjYdCdNLi8HgvqKdQVE3VX0wUVjZAfzmcTWtt8cxgqdZqt/M2j
waBO1hNidrIGzqOJjEqluUkb+m/pcgjOuo5eYFe5laSepvp59q5O3jfQdLlaIE/m
Js/KnROoxz5+SOjLbE1O7ilPeDIOR2sxQjQ3CJuKvRWaDQQj3T9Glxvr0wxnv3cK
YRmdtTlYf6kak8JG5PloAIZaTRLIbvdGdLU44hlORDNXeJFkDKQPVD09BLzr1i1b
CIBrdLftdCqCApK0/hjjJA35hNJg9VpRCf46FEPiVckxKrvBMAlFJAbAdUIzmfdn
fwNqUE7ZFjxH5tWftTRyV1bVI/Xp44wW34RchLy4sBPFZPqIGxQEBIvW+i03cmCs
i/mkr04u84qo3eQQ5CgKOSWucrUdocxYflOwtd7EnikuU4f4HvfRPnNOoKL09wi0
CbX+pZOyfuZye3trQlncwIMau0W2wcoDryF1QbOg9EGVYoVr5f3W1enUKkHv308L
C5gxEr5slDxCzfOqZlPFpO5y2mNoIeIigtmyRiuPxA6DBG6G7gFuC5oAKkOiYtvW
mWfdTq8kRy2bP7mPBllPSF5ASn5421pNg3ywTi0SdRzdQp46b4rphJGTuFdPx1VL
FDHdj3tDpdqPibCR/QMgT0NozkVJIHWe4d0duyuUlxihHYEysd2G+a6X4eMxUqM+
9/2ecZgs24pW/b+W3XiWxnp/qcEAg3gKBJGoyDCvReG0s5CTOz+J14hwgiArh0LJ
fTSpsd49GuxVedlacDJYOh+0Hj7UXX5d1jav8FQmFGbtS4CEjHBOeVkbaNUa/lsr
dUEQe6QJLcc2ueCEd0SJs9gNDF88hhLaQRpU7B72lEDXh4Nv2rynuLJ18GSIu5wD
JZxebdHazDGgtNz93rglBUZnb7EbdtyHUsPgQ0mBV1X01QNZf/vWTIplkyh55iZj
MUC4PjPSY1mpX6ydAguWMV+K23FXatiYYxYfJ4rxRN2v6wHvdLjXMTrHwUlQj3oe
rc7YtXfsqn8lfvErmHRfUiyNrR5d0fPz29gTADQGnBjdpzlzF2cSFnT6WJmv7wpn
c0ku/wooLzhYNZ6+mbU8YzlQ5fOYKgXLHi0KJ7v9jLIct6IdiPVX8fxqYdffLlmI
ycJNvgXZv1D5274K+ovwkR2DCOWpqug5L95KdGEdb+5CYtRqmFTPT43OPIOEVihI
KA0yRIeC4im9BgpjTTJlsJb6s1VVjCKXEtJwBTYhMR4zQI8N4RsLRy4nT7CiyAFn
Ek5J5HyPG1dlMvtkrauEFvBWSjRoIxJwPOGZil/ob+mNJ2+DOHQssSPDWnisEB4R
/s+xDNNpP+GSdzWUAiHCvRkTPKkMy+WUfZI7+uMrnQkg6oFNFd4tiq/MeRko8WgM
rhHyRpuPUQ0hk32bZg0tN/2aiN9YZR3DFG9SHrflroCQ/eB+J1OX6QhkPA079Pw8
rpjPXt54rd0bIOoEWRDkPmmOnFA86UC4f4i+Bq8q/6cS2w66vfa9O2fbh6YPWcEs
zV0DmckmRm/LHKo2Cdl+8SWxcw9xpPGaZHGLOJBzFy5zwUXaap+mQI8fWHYdkQNX
/bD7XybAnAiJ8bScvNC/CLCkMMADyYLvNcYyEsX15euWqG7TsmQy0wQoAB/jCrmv
ZaAzfS6STZD0ew783ipEvEMCu4BLFrdycu/EfVPzV0OiZv0LhKfATUSOdZHTzFhD
vI3tOMPzczKVT7Wc52CXkQ786Hiz9Ao+W9iDkw9Q8B4H9xW3mTNziMsb4XO0Wg0Z
A7sjnLMANwlSheMDPL6k2b1R4yUka+hNbrAytxnVf9yDS553p13m64fxvZYkd2RI
FPT7lw5Id6FY3IZcjU/Z77XUz/h91NMHQfPK6XKsij1ICqKnh0CjjzCSrMtxraqE
MeNEm0b5setewNkFtzEeKnM1mGg1X/mhROfphtmIwaVcp5qYH2sIA1BhcAFUKH2L
H5lC0YZkeVnZoi2VDnPXqQ5R18hW8oCEOKZhVctQ4ghGKtgBPNvpN3Fd9ymG/Y1Z
lbk3GhZUWOkOyMsBDXJ5waSWe3OQDG+JDzKWtc3HUzbQZpeUPsLct09OqD1rQtzS
4vbXahVVzmcAal3JNZqhE5R0JWR1c/qpbaPzPKPR4l/aO/TweEOKsrfvT540O69q
X6X8y9eo+dFx89Sszqmryzl7QeAZ1QjDRQ4le3bpTmUNaFDlOM3qtHsQF3NTQf6B
reN3PdmIScCF4c+PY6aYbW3uv1i0tOiJXlEiXRuBfu+jjgsJ5sFu3qPGBt5p1zNj
9+zdjqCI8H9OdyCBuSk+sHesodSpX/1gucWedPYwEK/nA0b2Al6gf9Sf+oepoU6w
aMUpI9AGhReNDfY9FcdacgWMhIHZwX3MSyE8AtGMuUTSdmb8YP72FsmJvmr/UqKR
iJ+PCyh+Uj99TWgOUbc3i5vbWk6kMJyZKg6Gs34l5Wqrq42pSPIrCF1hCwv3nHoE
VfdMNhplbHGJMmJSjcsnfKZ2LkvA0LSj1u+UTuWFS0INytY9TlS8r0PjPxYpnfcW
mIfvqhdPOlOE0AmI27QOWmpMlwuIcQOBGLwpvcw170uDcS3uAEtS180/ZxP3Lc5p
jq7TIVfYFSmXemghh+2h5Va8QYeFyGDzPiISJjrPUhlsuSzJoGNysxeXWuoblszg
ZVlDoJRCdK47c0RXddEQRLX1lJ7eKgFqZ152ls27lmVPIEbQ0QaKkiQPnNt82bc1
FXtWrdAycy/4yvJhA4ebIAiOkH57sCJnXau/Yq5D/Vpg3cfuCLwYF/mVAgmCvjd6
zqv+akgdRb+LMAm4Ef8EW9MG2kd0TjQtfp/D5LJe6wS7Pn90RrjU4rLa679s5LA/
L2EW1NuVjvpfZd0MKPceydZupfArpOARc9qrZSoh5jtUQJU6/uX7/tNvcQdoEV+f
VcIkiHhKW3X14GZUPTgMF4WN81yLztzBmpxes91mLBojavCx4jKbjVHBUKxSk+/2
oR7UNb95kxJb8HEN9mxWFjnGw7fVYaUiz5HZ+LwD2ZW9nH/6fnIfNvCjkmc2hcQZ
IStk2hGute5yqQTnIYSDaz+uC3HcUdMkWUQmscaqiZxl87ZCLRfhR0mfV3MagyPL
FclJg21b291cBYwpj6k8w9ff00LaVTtqdlE5oWXB3OIDIgz1Swon/Kp3nwiBDM5I
miztIWUAYO6oETWJ0NK7dA6oD8ARDzmrBi4ZQxew6iZkov3/t3HTy2CuE+QRcl6W
0381JgxQepEyNIxaqFfHSQmE0gj47PhvAGI2KcxPHrd64ew4GDWXWirPlNzeYDKy
yHDHTdjCs9ZVGqwq2Ep8bI58jufph9CkCQFQnZXM2tzOSdbhcniA/ip9vrXtGxex
fgn5LUZyQfALkbnVvdOmbwESGxDOJMR/4rcLpVQj7Wqrn+ERIL5audW3cuYZLEyb
Gi3CEIQMTSkCW4B4HvGizOH4fen61EXT2zW8M7KuV/WKGr6NoyNA29kutkSGVz9V
i2tnGoC/SeRX+4bx4ze8VQNGY4kiWhMBBS92sG0CWJgLrBuLlWK/smJFZSH6yoJ6
r2F39wVg6V0CKUe1p8VbbjYqT+eOh9VO2WDU7VwtMyzNUUZU68MBQYXre0Mmgoh3
MlfjXy+9QYPQbaZVqztZrW4HKjAqPrGbli5Y6fdL9gZFFPUwlOIibMCsOzI2R5Fl
8xvtz4GwxpJVThEMKT6RVG10cJ1XOeLLPONgssXV4eYVFX46OGyAT+QnawhP/idw
Khfh6bA5X/9nqKy22s3Foy4FyRjMEOKUwUezm52Fu7RJobRqkyT86nNRgehEwEpA
W21Of1UqzWYPgq0fHXabYZ3pg2M6bulbGsoQkaTSKmNJ1j1PpmJZ84sRGTWOJOtz
YElgzfUyVGWQZu1zpOgbrZERt5+6xQ4PkZr9bDeX2VOr+L2cl3A149fVrlIn1XUh
5EdOglIGgySQNGvTjMBSeEE6fgfpBRweUqWtJwk0DOmdUjctkPUDqnV5jgODOCWo
BMVqIgDgKjLvyCZNj96nnBtQOSKIp/IxDmeycA6+iAVEs6xsTURlzkqzE8f4Cosw
IocUYUADWJJmGoniE4GJ2wUxZxgPscXqY1IKu2fp1f3SA2ZwVqR5ZaPT1gPTM9c0
3CRIQOovDKLlFdfCCNc/+2jm4YClzWqH16E6FHoPBTtQ+bQIlZEDubif2+u9m/Z/
+jgKuaXUuRiJ88++q3x9+byyUoun4wTXlluwNtcMTkQtKlr4Ql1pCh3f8Vf8BepZ
Ja/f0wPnvlg63WE6cWEBBc1Cez8mPR7BuvAz4C6tPa+XFQfMLV323FeE+zz5llC9
j3lDCfDQntZAx119+I09qdUelGirGec8M4kH5XtrtvA2ZUGa7BEKwJV/LcbiT6I4
vFwCp4ZTVYMnU7Mf+xqsz1vcqMPkfN4iurg3Xp6CDIMo3jeDp5ZTp0uj+pg8LxQV
VUTrRHrW/Fyvu+D7O88Orv/E99kHNHasZ6gKAw8bcrm0Dtv7s9uTcazb4rgrEoTE
StL3UriYDZTiwixRqjd9JtxTMGur1LQaOwnrAMMS5coxlvqt+OJXjc8MEwyl+21B
C5OLtDvHTF4XV6Xp3iyLh4BQSk9y2cwRA6an5/k5HAgfRc1xJU3i3h3620fJZQRQ
gXe0/IiPV0AhY9qLb2xCI3PftnZ30e/UvlNNvPCSNRSDyW+qs0l6rdejo7ja/4NU
djM5gX3YjTJ6not2Q1U2keUGlv3eYvubOIl/U0Ht2fcldGGgZnI+g/IeZ2pjLwTG
d+d7kSlvOQBpnDrasjZQM/Ba7u2G9a7lufmpnA0LYZZfpi6KQ74l8V7EIfsgN/C9
flyuJmnjusowEiN7SHsEmCETGSNRnXT6DW9s9x9TbfIfQqt3KMbthE9rb9FuOVXy
Hp06YK+T20D+mB3I1Q7GFjmjIx9mbog+sbgfVlcwD0gGHx/axYj6cscYE/OIdvrm
tqC4GTCRKQ7JNE5yVvL/b5yCYcGzpMsvdKrsX1Kvrio9a+fJkzNlS27HhXQvFDMq
hWtYXqTL7hWzCcas/YBlARic7FiJwwjGwbZTG6OOUC2aEk4NBtM7JG1sN/Wd9L9b
ElctL0ms3itRgI5HrctZ+xyaOh5rTd/PExPb9rpHXBsCne1iiEnN7XJd0db5dIE/
rggc3MWKz84dJpp3F8d+Eurn1bLYYVfpRz/77C7dvBIOwTmbsZNerLCIPZSUX8tv
LhFFLbwrAv2bANs3bZawzOuUIEoXAL+496W+2AxDHufTLOEFO5hCt8NiIQRrvRIW
D072+fCpM1itf2+cjJNSHP+OIdQw4Of/GYkQnz6FiGFP3w9kCF5joc613vAYGwOk
DEghZpov2GZOvFlEA0voz/ORvvwHsMV9CkJsT3uRw0HECeE4tvW1zYXp6Kkahf4T
DJPCuYamm4DBg0F+91svUx8+YRwsbnwaEP0dOmqxBW0QNb1K3neXB5XvjcgmkP/o
KYFHvNZTNzUtz7nju6S9LSjipz0lvss4r4eaLEiz6rQ+v18jgVyAQVgNwZwvNE2J
AzepYhfgdTVuj9hTpwqSJdZ7RChnAYAg1SMFcKqB9CH2R5J+IrUZVisBm2R+i5MA
NhAZwl9Jm2xHQtukmhGR/13A1g3i51mZsAu/NB1d0gzYipuFDanjcq7fR93CIksF
nuO6GXl+oRukLmOaVoZUO25ndRReSyVqtn0ATdRm3wdpQ9HgNGU2jJzr0/zuRftR
5oDJty6pgFZ7J/QWqxRaN5OZ8ZkYAbJ09lqNlsMKILEqyu5SkJwnsPDlk0uHv7Xd
MUM4pE/wmRUSVvkZizXCazoMgIJza9nDxnSVen4d73x3PbJetpZnVIsuINE42jih
8/dO0ri6KzaAkMEDUJOPfVwvRmFVmBN3/AQMBTpx+8xHtgjlu6iwrQbqF2gt7LCl
AyamOCZQppwHGYER6qRVpLlyMXDe8rzSPpZQb7no5IhAHUknJSn1UP5BaYWF4YoH
soP0/L7tTH7jdvogzXHi/cAYWA1c/eiDu0puS8mBvljwoSRVBPh1kWEtCNQXpvVf
RWKTxzGQJY7TE6e5gc5KWSD7/BmCbTq187jzWmdzzkYpGTW24hoz654CjZ/Hgs2u
OmFVFzw0oFrn4lcDEE13JtCDd7q25f65BpkbUGgGhafXLz0JYRopn3y9+H4qa66x
jyzwIX+Ic3PMByyUNmR8c7kKYA/Fh5USuIn5p/qPKZQkFIm61IZI1YYKybttrCcU
OOuFPWmMZX43vc7K3FThjz54WWAJoUpIPD0JD7xo9aMNQuvQ5rlNtvsaWNt6gs9W
QkzLwUW9qerrItQEXnLMLLxgMnyQzi8tJObpIsHPzHXaETvY5/By92Rfsv6TytPc
WT88w2UdPKCIDgBr9FLWNEDsE5bhkS+NwtKivw4P/mf2R3HfYIPOTQKdVyedAj5p
E5mAXLkngSzT8LTxPC0y2IEZ5IhxzYMo3I2Zb2ZLhBX8+VoPOk3YBZvAZuqIutDJ
Z+tM5jqlFWCfCVVWNGl3xNOIz/WUjRHL37dSFZ68NgZgDNw+baEIgZTa9KFIqv/d
Z9JY/quAjEF3/4iUJN6ObPKsgRNKymDMT9admw5mremm7cCiQlgpZB5huaKWyyNb
frXTXo8LbWIMSfFOFKsgjRqWe3OXaOt8KXiIkS6QFUh5BAMxhNmx+jmSqNm182qE
NkEN9nu086tSqH/+RSbyelypaqYo1tyWJSL/zfXsgpTbDSWOdCkzvhyBUMnxCwyr
UXAqgVPk0VXsTh6k/n+Ne7pn3InqcvWiOGztajhOjxz55H8S9VToIAnUn5URRsHp
y5Vy87e3GKwuS6NpxZwUeIYKZ+x7FCa7n879GVPdBBcE9HG+GYei4PDxQJjRUIV5
3TV8R37clF+hQsJLCbqDJ1wRr7Sp+KOexnN0rmxcVmFFneU1ots2uH3UFjrTrL7L
TsGcWkECtUZqrzhJqLfg1BnZg+2RJcfA8hz64Mk6uxIr/W238oZUjLj7gw9HD0qf
ExqgcFA2DGj63PXig9JpQFb2SbIotCBuQ46Tl5LNDFzM4kO+wa7GAjtWvWp5ykxS
7qsL/TFNmoOPCGGIn9H+OAnfp2Zc+XQpJVDJNU1Uh02nLB30k+NyhRNC59anxHl5
ntPW9jRGiEXzo9jx9xjfcVtd3+TEE/bJIXyClxDOGwxwmyXGt/0JDMFs55f8R6qd
7op0T+aiiHCT8vOvxzPjC0mO4XFI/fRN1jWLbE+LDXy6nEFVtD4eJwvIw+0SfO0+
fWrrm1A5hp9TquSajOPGKRG1doVRBogsyZzBbpta1q+D4SR1Kb5fq+dsoANS4RGq
oHjoNhCU+ccYpHBNCJgJ4BYj+7A+OmAhF62hfalbwDXPcl7jRceb9vB5jY+OuTiW
rb535TdUuF6lppwYsf6hjsB7GC4ZA4DgEy3+hDai6WyUgpxKXWlyNWE3LdcWXIb+
+Bj40BX5e/bjLKLbkoXDiak72hUWul4HxBppw+4+3sKZkxMMUAQiIHZgknYAT4sc
pvQJBJrbv15q9a1EWRhPNXH3BZg3+lCDQhSUrA8u4txYtB803CzlF0FtmvwoV8qw
UW2SzjrjHt3/AiI+HkdmODLH7arFY6LqbPBAZT2hs83grd4DsxivLm3aWuz6YmM8
Rgps2dsGowGDmH+dMCvNhUgkhSfJakEqmVVfDhN7q/boZH/zoY/ZsPkvJ2GdaKEB
gs8nPRJUNcBsJcvjiqMD9CgHhg1GaRwfvjbMgJFwT8wrnz/r6KkaSsRbVFviARLz
wXohGibokQGONVshqjk+hc8l05IYHRGO0R0Vw90cdnAD//JYQh1nueJBesbgWpns
qwJ8NIG6w60Fh9xNvvk6JUMqPRwBHyUo3c4h93NPgTtIHjDpT/e8Lmy9X8u4Furu
aiELnIZd6lWa/8tsWYjW+TlGXEeBvQ/jK2X6M92w8Vl31Ds0TtLqNzE77JvuCvKp
8mQwVEGbesy/ayfM0RCGRRDTZDvP1D/tTP/kVspvNGB79eoKFbzUEHycgagjPQ3v
4dIsKCmpTCsa4kHTlQ1d9ktzthrlrnQhlS+HUclxTNlrxXrj7NBgwovM5kl8PJSv
44IJk8cBDH/CPiUH+rTzE/JNfE7dVClnawidF/MTI6suOa7xVfh6OtHCC818uy6P
orExoG9Y0rwQQGevEUvghsvBodKyg6ivDhFfxYIcr31mUHOo10XSCVx+XnQzBhLJ
FG9Lby3fonskeXUvIUohpaHEyE434g26YkuIO3JYEr1ByhsEmVPcvE3+RL5mpUop
XptN3l1IdovYPdORRTmx3PdmcLBaSSvnP32iOK8nlz7doweuPWXTEkeVRjWYDQk9
fwpenhqp6yrdWbignePfxdOWaulRoOY9dLRvaNqmZicIxZJEE11AxpdR4i1yuAVH
LJcx4BgIm4UOtT6n8kdwhpGN2z/vJAY9cNosaf75AagdKwJ+gaKYsZIppYfku2tF
uGT+P6CLGVlxCaSPytZxSZQPLyxJdKE3dciaZT52WofiQu2zDfj/vpLZX0biP3fC
hcbXClW7TSW8P3WMumE6S5aZpSrWlZQkoevUc0dcrgs5FMZM0a0l8ZlVRF3KOqCa
QzvFTqpnIVCK31ET3IYlWZGtEG3feDQv1WgIvF4N56AO32ApSZyH56sdfXxVUQDe
RxMOaP8/6SHuEBpn+7lSP63iLqyvr0cDtvbvkX+Yoy0aj6oUhbCgS0opQ5ouZih3
0062iCfflvPQKFHNGBMELgukEL14cDfAP2DnziMzohugNYpa9nTAAW3rgIxKRbtu
UKMk0ACiGmLCXV/3H3TC66xJ/pXRjJZHmM4mLJHMmuqe5sTExcIU8HVSgf2YvlY2
LcqC7FOG0+biJO099BvzymEMpGE7WATJRcucEsRdACNN7YT028MzGbgZ2+NWkosi
y74a6mqiWj2nBzSabxqmFALmG9StgoA6jo76jXgsXjri4OzmePZTc4ypAGiD8sfA
FBChkGc/629hI5LkMva8MPYXYpXxL0ukO5U7N2p511RP+0EOJ5ryP6u59c8jYnJX
oLvBpoYFW7DrWHWSmSkLKQza67mXQlTrVwBmrRAIo3lAYwzokgoh5fi17i4qcxii
5Bc0KV+ZTpVmB8FUERG10k7ootqeBOoygnd+x8X/CoEdunnoH1f7dqAdqyChkG2x
o4MnBj2UA5L8VYJOzIZ8D396eUShM/NDEPTkCOfJutBzhe/7dP/sVzXwVrq7UJVA
vgqp4BnJcb2CHj1TUcQ206KLuIT5b6GC9AVJyIW3u47/eEJT+sHqcteA0+Jnt8Fc
kWdJ5jwfmx0N/5WtQ4F/33vNdjY4YgE9Tbmi0TMAImZk2nimtSF3eWyLR7fr7DHj
vfZCm2K2iviIT0rSaoeQ4VSsfeSLoNc+uCubfAOfCWm/j0VRhpkZn0JbuZtHa0Mb
9OD2d5BR9rKf2UxDmEGd2cQr+oTREYK8ZTQgRJLf5FaDWGQ3uuQaExczxrLsXiiu
I/3JwiKzq713EzTCYXG5D+qslk63OD7VG2gg2gce/TBTTsEA4RQgxh5hFOXMTwI9
xVp/RJvJBlsLQstFmRAsymZwxURZwFdgH12Nq65gMZJZ5xDm/+gaWytAZuAfk4gI
6mt3a4KOHr5QCYQW+XozkCV0V6VpbSE4bxaMBkaz/CC5aXtCofh5xaxGb5MHEEdv
YfgSXe5q74lZitVEC3Nb3BOS0QLrWIjkab2Wg1+zd5AZdPsDTQwqW7I5TnVia2WB
5pez4q60sgeNNBqt4R9xpZEvAAcGJsNpk3X/+wWm90F1z7XwaMCd2weLgh99Db55
A9Y9IfQegqudbdRH400o0WgsQJIDKmN6U70ImEIurg181TzaL+Jt1Fj08HwepyoA
2Jk8DWsCv1VbhN+1Nh/iNV8odDrGf3TelAgSxHEPD5J/VOv+gbC/uY/Z5296Y9Mm
vftBo3hAD3zS2+rbFeFA0Aqg6rpDMoGFxqLOJDXQXds/tz/lDUGtxzTTnW4zUCZd
rTkRargyGgKs9Kfk7CD31f90CLp19cEraJ+GM4NlA1L7VBKbj+LoQGWuJNNBN83b
ApaBu5veo9gpqqcqRpeoKyT7tjzh+JlTpz3+t5N/V/R23Ar/j7sSNVBvWBSETyJy
zrENYXPirGkrukl3qF3FGDFePGOe00HZPCC7OJhGBP4qcuUOpdZHBt+HcmX2qS91
dVw5DxFJeFJFG+xzQKIRFrgmh24rCVnaCcUC4xLlJwBCsQZpANOex/vTBQB0dMoP
1ZsJ0L8OUSl+xBm9hA41fetiBXZ0uxNZaeaPio1UpYMjzKTexHgvczsuiwDE59+W
uXr/IAoTXvzC09e47hqdMDCu513QvWISgxOQkZIOLhEX1BLVhKJGRkdfh/TgyPmu
HEbwuzSEgzhefeiRN/cSGoUk/wDk1wBZZes4OMHEHUTPpZZY8olhpRM4QjKMpetJ
UzTo6t/wJRHFwptHaurAY4x6IPQH1H63tYtapLRblmf7jN1bQ+S7lg9YrC/vjd3/
ceq2n0wlnDR1JiWWcrUMcagutHeaO+a8zvfZVMKpk3efk15r6MnH+3OKEgzCEqhC
temaLtEBGuRMIR4wvJPWfEr6T4YQEBLiWCJ0VP06h2fzC5q61IXn4Jucyt+eiwK+
kkOFRnMO6sBSCphTuRY66DwMQxVk3TpkpWWOui/nihJeceYiKf6eYPzRU+beOKSS
pT7vs9AWTFJdMf5hvU7pGzHrsNrWG41vY/35Ws3NLs0jGG25Mp1t4FHQs1Gj5Q3t
DQvWBF2YvzilWxl6uDiQrh5EKuyLpXC6JhSUl9DrTuR9gkJ59VKh9PjpYuBNWgO2
blP8z428rWyuLMK3v8QkLWulSsROC62Qduorh9NAmRtYWbm1udHG0u+yJFrZwDv+
6lnoxsdMCyav3jERNWWSLiH4z57Ihz6KsgD/C2BMfEER5rBvXk11Xyw0LrcRn0We
EiJk1LyXt0cjABdvafhP2QjPTjqCLmob5t2d9nH85x917dv87/zB2kc0s5i/yK4a
zSncqvUIG0gyNpErStLcduS3kqDr+XfpuUva3mVmAbiyqINXPP3uIMiGHRsfT4nY
Hbpt+celHZDkACDI6NxV5f9s0xasNb+nsPpA7BHtKZuhzUlFFcv12ny1LFrSyuRE
FFYqdTkZXJHIryiaRdkp1PM74UJ1NRLwedXTTS0khLw1p1vAFDl/blc9BDhz8BQK
Gl2wbMpq97Ay640M/445FEDzQUycx1yeSQ0e4JIlUKt5A5gbrVwKCRUf6O3OBSk8
DE1QZM8X4b/0yJCqqGATsU1Etc0+2x+ACSFP1TDgcRyT0uAIDXDy0sxcfQeZhRIA
55thGOpnRqmvhYrubI+oQzGbZ57NpctfWLgJ8bIAFNQOR/+6jno/TzrBm7ZTFGSj
F0so6PuHLbFzGyBvBNJBzSqBfJnvApawdIcSUpgkyCN0zeYmEwLq2xcAVWFoKsTW
cdmWZg0+tqJ/PX8KC/PfHTSQc+cZ2kAU785q7jsIfPKM6UE663K5gDvX30pM+VWa
BOvI/dhex5iyBRW4Lt0I5VYQno0j6+2th3kfbaLRqjF+4uyWngjdIfJfbb1UWDMI
TGl0nmmIFvl0J9Iwy8fh4Dtu442WNQFUhWn6BJE/uOmF/MZsGH1YpOgtHZtnvNBG
8X//FqFi9frNuUy9K3x+tRUhSnnrQcYay7GDgs+n9qJHeEeDWZSuCsJpuCOmnFtd
CUwHMxxeMtyD3yPcDAzGlUCYutCsnvXOH/iiGFZSfjGWk68QVGSqTA6TUvAlXIXm
hVng+CipMEpx9brJ0TO5VpG5KI5YNzEX9dcTvLSOQtGQSofUKStGdT7xB4/voTZy
NhBKWHT4XdXF5pyD8RXDh/kAkNpbzOaTXGX45w+NGw4UV/AIdBw1mCP4fs2jIjeh
KPgJY6iOygtyhgpqGzGpdnNrD1vROp390wHQTcTEAhPGDUNPJYj9OXX9bSu6ShFL
u3wHO/Tar99MG2zCnq+mIBAz1rJt/UItJSs+tnpW3TEkn7Hrj4g9phLld8GhHC9t
HNs+TqUYEhMoGrEdydGWuK2/q3Uw/uPz9gw7p2d+OsG0+74ou+PlvHO2bgx7oUo5
/GolF88PdEh5LSQ0jnF7cOAYS0t0Ngx5+hOfsdHGHX6mQQxhj3zrmRDXNX/R0yKZ
7R+sFGdbsu6bM0NC9Uxrm8y5q0OBa9Ce6UGkpOT6dtCkQ8fL5wbKoZu5Nh6OkdGd
c4Z7pA+sZoVuq2K+vw2GjJe6ms0N7fGGHVLrwp9etQAYkoINqmDEVfklgvQnp0yl
p3R11lbdMQFNMXJDpB08DTtI9PGyMFFLqiqVL7Sq3pDjMovwUD0tds0ew69PhxMP
+v0AuAH53rmgLn07If5bN+KRfktakh/pju4dQzT/HDmP6CMjeChQAoRGxMyT8lLg
F2PQaCHQ2flAPOta67arUzQQTSOkErfJWfrQHuZ63aLCZPhLx5/GvpENtDuW3cm9
Mjp65NTciT/9DKNlVmxbDoraZZtzbPREoYkyFwCahrnU29f96YNv1H9QXMLCi8uz
SJNxphjGrq2e6L4yqvzSb3MuT3Nma4sH7leBOqNET7vJhKXz7WL4YdBwlugrp7jG
ZDB1c1npwM5DhwxgXveCz5X532YgvpfhYmlPpg6MC0lTiRZykKICA09A1S8U4dLM
nvpuaVdr5coGdDpFnQnITGZwPVic2hGFgK/7zoc5KQjBVTl83hg/LplE8iMdvrwD
gjAIu66lM+YJyn4m4LzteYYVsTDQc7mWbdrcruX+wfEINE+1KKDqebdz2LyY0VHM
nUP8r/ubzwOSfVv/il8mRAXVTdlbb40tlNPecQSXAjAp5GFuJKata7VcbqUxy5OK
Wzr/jic2sxgjBVjzCnYi42p0Gs9gxFPEdNVxeaX6yzhKLxhyqgzZelofP9QMcne5
xskQAJB+9iKRRxy1eIYsb5uRCyYjv22fRjhEMze+j6UtilOYzzPKIj3NwO16wJnO
+heOUaZXaVTj+0NC/3kcO7rXQQOllur+6StVGdgFkY8Ms4FHugkJ7KeV7NviwKoI
nSxQ6eoq/MT6WnLvRa+06muD3/9sI3/Iw2KiB+3RGHgreUpkPKkdE2doaH6j0J6T
xoXgtdwzFW1TQrqkW3aNQy/Tv9I/+iM7go0Uv2OdnQkafd2h0/Tl3OBrFiBGC4mb
u8M5bVM8c2zad5e3w9cwgLDuz6lbSTmd+WOQHa0K8ZVCKGErUnN+3IHWq6GKncMn
NzK9Fu/GIftsucdojEPaPRD7v6s70rO/p7Hlvrwfr715Ix1QzWk3T2uwEl6k1Uuh
ggkg/H7DPm6CEtuznIYL4Jq5Q7RQgnVZvtGGD1mB+9u5fNRhcIv64iu41DntkvjW
+41rCr4hw6P6igS2hKtZ42fCsnqJTeTLK/7tAiuACY8VcQwdWbvhaEIl8+amirMS
Mc3Q1cfBLomb3Cj+FjiwIIrKImrr8sUhMP/Hv6igyhexTFDJ7YpSLLtYdV0GG7T+
WmxiAIOTSLqxaDcXLAUcUX4pWTVK8Dr1pFqdP3ttFvIAwtSJLmGlaq7KyY1sEzU4
KWy+956BKJeNXmwdJMzzUA8VkGZ/6y0X16xTk59um3Uv17yfrk3y6f7cxYduNMWB
x2vrzt9U6DAghBQbIsLsY/ThMJAVZCuBxzcHTOR2EQ4aweeij6FraxM5pCSVyfZI
JYhqi9R3sjMHnKp0U9MWilI91tsRnQ77+e2J78Yd77C1COtZPornS793cikv8kwX
/mtUo1Vvk15iJKv33jQG9Iu3Y4GJa3iuY54VR6MoW7NOqy59RQjmnjlbtH862iz0
dNbsU0lUQIQEQEqGw/IPYEqwMBsKtOtHPysANmlvJxyUIWfz6833Zha65g1s4VWt
di02r1vKZWjPBrVdWMPEMzpHRNW9XFyU3q+lnPEBeSPJc+owz4meQXS9Z3De6xg8
VsEUf2PHYKK9e/ZzXtGxFRO4Aa/q47/BXyTitO9Jrem0gvLvy+4yoI98CrVh+kXQ
y6GKJcSaRuSIsGqNxPjMAZGGPjiGOe1VhLg2oQV9LGuvLesRWYrALoFAqgdve5+k
re5ldGe7v7tqQDxrC8p0inpZqf+FZEQEIWdFxh2XKlu6VXDR6Xp+yk2VvpkNkMHB
8kTOUh/oG1wy0VJiUkm4rl2eulYwSPnL1ICbVkqBPPa2W0rjjw+RcyxoD+r6zukP
Vbaaj0DiUsIVx+EXgGDNgJ+wSk6GzTne/Ek28zw28xx6gpUsCZPijU/8wt4SX7vr
1pmTuvWjrej5+Uql3kyvOZRZzxUl1uPnmxmSLXb5mmwppEeGN3aA0IIXafOE2Cb0
9QMAuRkW+g8jixr630IJciQQAG5qJqAl5vyfnjYDvYiAkDogRWxB/8ANfQOWEk4i
RXTndZiO3qj92Ik/uJqLmVVsfCOjAfYD4hhn/Bi+WADS0hBRQiDnPTQ3BDEcgIJF
Nu82IF1vfXK9sFuKyo/X+z1T4r1QE6LM+AY8hJcnwG3e6UpqS6A51m6ffi2E8I3Z
9jmiQCL2BL3uiG9RRFYbFSYVEEIlciDPhxYZ1OXVb7lXdqsX3iwjTI0k7XMuEzCC
86yKPUfQoN6b0FOxc+HqYHtbSiXTtZ/8EVm6JXTFSthah0zaHiZT4tDwxdMXq7a5
5YqvFfzhz2Vmt5EJii0RDsx1NXskjGhlB6nOOhZCvVuErC1YphtrHs1JLHw92P4o
AdakIlmofwKA1fNXVMyHZPO9OoLuR7XHYM5fYDAaLLZYTiO4G4qh7NbNDEi2nEZk
xjGY11fvbU5fw9cO/fan2o54eTPTw/UUvKm4J2gWg8Nw1EG6mo0u2t9uHqvSxeIc
z1HQeBp90Pt/4F5eI13WezH0PzzncnUyJSQg/PDuInJIVYbG4qvnQTb2Kaxid3a+
fPgy9BwSHlsQ9YU8NvuRJ2nF7XGkzvqG532j2E/uMz+egPqxtzkGsssSTRXuBg88
0jhdsJDHpkuOiW/IMxmcK+FDAjov7KfTNUxd85elwhJTkkGsl8U8XZXA31wsfWxx
Z5CJ5daK73fahe+nzxyklXcm+OEPNVnipeyvik+yfjq+0eGEcCHlt4seQZW+6Pyt
PmLAbqrWkT9H/D4WyIukFzPgTJSTCwI/x2LPtyVhUHZuwjQKkVErv2cpuNZWxDae
VQFKYx0vB6eCXKfQ2KNne/MCFTKyomcqHWqJBnjHJVaI9Y8kua/3Ya7Qu4zFBQek
i3RY+U4G1GVi62qipO5Hry2vENsdI5b9niKIU/FAEIcxCsrbWpUt8ldzTnxyAPXb
VL2SR5IHECvGAdhfinmr5zuBDkX+f3AIpu0hE/J3s+4VIIPdmrWHIkNG3ts5C/q7
rveyDSS3BWspYD5snQg30p2NC5y7wNbShPirwxvqYpLY2EkIuKuBjLXvy+yXj3G9
iIzatChlY/v3X+RCw1lzMgafq6ltKDIsx83CU0lrqmQx2uXbS8sgIRIZM5oVmhmT
j9h1AqJ8MvifHv3ZywvRHCXTE1fTPlUkPHtTjweoyxd6Pei6wYxRpqqnS4XLHPNq
se/6dS+Bk+0GZ4OqiPVlhTROJTEpFsHFxR9RDSe9c8lEuEdf55StWRDbGRNJfgTr
fYO/k8aPTjoTiirAOky3bU9Cj5cYHdu1eXlZBnNU/LmyrVtipGEgIjdJXsQLcQ28
ctFcjZKnDgykH3VFXjbVVybV8U6FBi+VDz/HUCuQ03KDmFXTUES9L4kyg7EG6ZXv
awPGur4nqjUF0yF7mPZxTi20fbymte3uGtkBfcSZyXY4F+2wH1AYLlgNflhMDhu5
53x4b1ocgdY6nPmlIDaB+dCuU55IRg+gjcWa6RiO6yRBKmEtGIHQfLgVJhR0ouPu
woomOmSixpYIDJH/h7INbqqrBAvVHPIwZfcmERU/27E5N3aIMsMYDiQURMZewHyB
ISgRVROq/e+PcoP/GzuIJsHUSUZboncFgNaqLcPJo90PDrVZmDi2MMJOXfvwJDwc
hyu5Rq1rWeXiLhFJKBKMlIJ5vUILmQlG4JjocSRK8glBN8BdwMfbT8jW0WHKXaI1
tie0VxXv/LxYpNrfVquR43WMHA/BlUuR1zLC0R+BS4khIcsP6yt6GwoMUPQnPGSY
fpF4bf5a07rz0nRHA4B0+tgvPnhNoSdpSPF30PNB2FhLISEbLUVl6aSOBqFvXXxJ
7xrJXVpsL8CLR/JGEbO/hU4TT3N0MzZM16P5RPWxAGdlTqembcxw1b9n2KfT2/rw
AH9N6aV+/5lTgUidW6/05kW2oyZwwvqWtwHl/AMFEsAe8p0GblIrrUgHUrDcj9c+
sGp7nEG6r0r3aUZkIAh0g/7cpsgyummcBcVfsggEHTHezmmyxQsT/Tlk+HYmMbkc
RotKlUErX9yDGLzS0ikuWgXpoDGtb102yEyZqXbaOOr/1jtz77stjGRqSyLNefVR
Kz/dkFZkcMkOsqT3GXe7LMq3Rjjdkku3lsSlnsWKVarx3a1j+1xfT9+bZJq8rG5H
pzZwcjQL/iiixNNnFfdFulGi4K0dy1aGrCBy5JS3StBtaL79o86ggkLAtUp513xZ
7aHx4cR3lMKoJsgMNAG7rWmPMspuYsREenRRahwuKGpnq2V2v8kVtc1MTymK47BD
iTQV98mmH+VjbGCMgN5xB3S3bMcM06hgQ7jN2FOviZULmrEn2glnWEQ+lhmVAnzB
086U0z687tAboBlrs0fsKcoGlRv/D5D0ZpoCJknLFbHlAOspP+0a+fvuUS0YNSEj
IfGnqOkxmZN82pc+ST+v7YSTniOilYa9vgwPLLGiYUFkDnpxfiXSOkmWGyh2d/1N
N6fh56KRiHCjnhwoBInBBeMVr29Bc49wUukfPitXHHzfZCeCd8GT6/DJrIQKPWkp
eKbJ5qy7WrzW46LsQexs5sd1U3WyKaqIYooJhMtsKjWFPLhCgbj6dS2THzjWC0bu
pBB++mT00dOnK3KFs7gz4VElr2TSxKZkzx1urNb/DEqhRliIYEaRl9W+ByCfBo/e
CpIMhUpdSpu5T6+PQ7Szf/Ed/SYOcR1x2K2MXQgCHBwt66+C1OKRkPQdKnVXNggL
kYNONJfD8dmYfB79lhUkj3W6qxFbipfKe5Lq4nf01ahcBjVwug6z4lNsCMWxcrJw
qmi3fowd8Ex+P51Ec5TF1dsz3wXS4ovhscFVZ8lrYTa5E0wkoQYCSBfz6RHt4/vz
fgByppQqJChgGxQEjrbJ1JpiHAI7NZvRHJYPCE9P94oFta4mjBX3cLeBcYP0ngBc
qYQoIYtoWYYkXa2TTDXHri7GrmIikbXjDCnnDGUypWmPQBzWLQlNdOb1zakZVDOi
gw0yw4h0N3X9/BHe694yzcHJzm+kb0HMgHQ8xvqO5GBgBskRxZkCx3O4yWdrdxEY
WDSoEl/zzzmmPVtXWNUumIj8LZg9iSOEOgnryVWNtr7MyltPiPnol/JDdSu8wVj/
6JFX6V1oMT5y3Ub6Cuv/zDQiF18HeQekPEeS3qMrIrbA81feflBD0Y1w4ZEUYxS1
8vNAoIu+zq3OEFPD56mfm3WMMqU8t8Pc9LrCv6B6z+teCS/UC1X96o1uuZQ1vJd4
ElBvlcLFcJpe90QQ+KoPwPhI/4KuWs+p5Dc6yusj1mk/PUTGI3k+46LCsVH4Ramw
AwVS2L4Eaqi5LWrQHFPAAghKwKIGyJdQM/gbCMZ9onyvpM6OrWB4JQlZBTKgu653
VmPXBFatOhO6O01wBZkaWuExDoyQWAdrL+Hx74NArQuBJEufdz1eejaAVh3q0PsJ
lO+wbfWcZ+/3DMsCwABdnY2ZnntWYhxT1KHrkKYDaHR6XUTfitdMYBxOvo6YRosN
N3H3P26d7TfBtBpiaYEki2YyL0gwXUdx8H3MGxYTSHtjnt6Nfgny7F7kqad72Y5X
zfh3PCuYIpjkld2HnpQad9ualFbdIS2xuvuf7CvSLkIAHUKxyp4IMKusvJ1RxWIM
Jb/28le6eBnqhAWapZwhcFBkqM+ZZM8b+/tVHmv2UPNEO3pPZqmswDVWmNP3sX+N
JK0rAMoBRqZUmNzp7L7m2/Cg6Vi2BRObjKx0um1jKXjr0GgSOiSX6fB3dsz+aBeF
en0IuUgyeLDa3JNi1iHCTKLn/+Xcy6oRMJXujgKDbXhmu5Lyxq/6p+sQan5l/RbO
CtWoT3uYdjFK4+trpEWsPdh6Nb2ptCvarp84CYBH3aTTOpZI091VvVKK66N7XoNr
pvs6fVvGLc+SWDkdwUyDLz/ooKtXlCpifoLSCJz5ww+U/MFAWlJ1cDf1DOCm8iQ2
94Fo1cigMy2bR6K2drWfDlJ5hn+6DLOD5zu93zd5LA/+oqcFX0NvIOax581nkkb3
GA8jOxnVzyvYLAptHYjUIW4XqAT9NTN1Rr2NVBx5VVAQA+geRUaKQ0pFjpdBUdYJ
E9SnV0HBFUGQmT+6goIRgsExFjqYX21b1z9uYeU/d9KACKRwB2Jjs0KHe2zz7lVT
AP64iBJ3M+Yaf7XTLum6LaI9FkVWegvePJgq1Nc4RlGM6pbIBxUc8puJq8WF7rLX
QScoTSgZN7lqwJ+AYi9vZ4yfQrjS2eq7rrC3/wvYuaRVtYr/uNmsFJ4v556TK39P
JcQDJx5qJXqsRC6yXl7twdMejVsYdUn/jG5TUwzzkIjGpy3TkqqPuVayUj7kh7HM
CNh9p1FgGbZXvvA3WmFQunHu32eIprDoocwl3k20kuC/VzMBFSGzmewzweR09Bbr
F9Hog/OgRGxzfsNCW/JN0idGjD9E+E72r4tOtT2A/TKEHlpr0/A3ax3JAzSDs4nC
LwRApieh1tXzYii+DktyQgWLdWiT1GC0h0iJNrGbJare82XqOvegKW2gBVNTggL9
pLI8m1FX+JhPhr8cOssEtcIDo1YFzinVHTPZXZrXl3Un4257VlN3D83JjJ6N8oy/
0JKRRpnP5yXCWJbsQeahTwTpwLesJ0hY4bAa8DmLpTtXXm4wJkWsdCXQ/rKhtEXU
asEuFhPUQR8HRQuoxMtfxwi9lUwXhddtp3LKmsFMEZSbcCYB2sGjnvF9OqsSsmNu
c1F2cV4vu923gU5m8iTkaaJ5dj+3OYaOGt8xrQ1wHvXUoCFivWZgHC+CB2ORp8Ln
+bk3DHiTUV099hHAplWNNqS+c2+eNVYEXTsEbevcfqVHu0857n11ArQLTRR4DODX
AfdEKbXauCENmCTCB7G+kddAV6WOOPD0UJZTYsaQhl7B0lrekrZZytYXhpLNeB8y
ZahRz5k28ujxHQOcQCwIh4qISbN6570WMUcsWhqSdhLFx6EHMi2kXrgkVrREIoDo
uS/MNT3HHFChHkA8kNM9QzEywLE2E+CV+0VqGihDrekGH55fOSe+cyPoUv1vidoe
G/s/BCYMSP3DdkJNpy/kJiE0ETBY53nx4e/qPRRbsPrq4pSV/SJ0+Tj9Qhvm8Zjx
Y162zV17o4ViYmE95xEG57F6rRozzbx6VjpmU0DYmWnldUPuEp0q9MiD+GVWaeoY
khE0567KeGtp6aqBErceEQSmq7ptZTEYb/cnIATCh4I0jRsEZS7KKBMEAm1OSkSY
DXHOgCe+yMiutVLHVXM9PjGKmXgnfLMLhHZ+SmBkNN+x1dO5zuluOXTes+axYrFR
HFeuFkdbjC6nV8Kpca/XxJ3jKzEOt+dhvZ9rMJ+TKRYW0rAMDmFlqYSWmO873lMG
pgurKnabxoF3+JApZz5UX8TVNAmwZd8Zv+sjQ9rW77qHc4dtPWTHhQ9uXl9MQtO6
qJhQyNruwyeuMGaxjDAwwSXWv4uQi8KjVvTlgqs/O0oGnClAvfwojU9VuJwD3WgG
RSXkkNSpJfuqgn96rPdNKKKs7MyIRbEhUGzsPBlaM9f6JJEcHrOggeVVIPev0nh3
RHQ+xXljkst/4PZAg89RLjiQjJWNqrrhHRrGbETlfn3ASA7vdyIk8q1BITkEhpbz
E53Ro/H0fhM6DXQssIbuRz3Gl51a1pB9byeukOY6S58r7XqgBSMITreavWLO7l1/
WV9K5ixsniQGEeuF1TxGAl4uqn+QOl5SoJFCMpBZI1kqR4QM7ELFznNnt/DkU7Qf
+Xu4+7vUXCqCVvdG8y18Oe8kxDP2ohDl8/fHX3us8X9C+sMCceL8Tzz+GeF8JIXA
MpdJE4WULyyykj2LUW1n68ZGQOGhrRbLGUXA6F52PjD7nNzGWhzHCQYJ1FRSmcuD
jpGHKzVEyewz+fX3tmZYKpAzNqmwWQCnyTrA5UdAX3bHyMpDRsC3VeyRW2sb5lP4
YsLO9+nS/NswG40aZkX0aRRPm4pBH7mFRCjhnCw880h7XGwNI/KYrPj6gL1cgxAN
5bjQJDHmGvuhDNdeD8VKCr5pGzQeB4PxCSLN5Wjmvc8HarqrgOaS6wVJE1+6WD25
mvpkzpsnRkYSIDdhDCwbjP4dPm8JAh3pwHTmNAIlBbk7nTcAIAgJR+A6LAXT0f1S
yEM4l+fWaIrChVm0vk+CAx5vqJhBl1pRcyZbCYLO+EAJ8FFP/2lobGLdRTrJSjvw
fw3CCy7Jvt1uX3zQI8aEAaoSJLi0VCll7TCm9gXdYHp4wBqaBHlOlNzSCbb1EZIJ
tKnc+W5SklxUF9ZeyP/m8Q0cPvoK4c1cWcVr7VIaEKIinau3nYJFupVFenj2fxx5
iuDL1EyzqnJFWP8p3LKl3iAWZel2himo9BBjGZqw3NUc/0IthyQYR27p2JUdPbbx
WQObiBNnjrN5Mx0d9XQfh8lcD3qjvYpUQ+4VwlzeOD4sj2wcjqCvWnxJK+BhtO+G
y6Ok03pHBFzhvMwbR45tXOK1CmpzcYidZCqBFxMmanGwori6mfDSHOUF+jIWml3g
A4QTBbOsRgVbr1OpqcF3JGyTjMp6M4Be1KwEh6aypRjavcQpkEzoO1UZ/oFDQsil
Tsm63aWkVx7xISubtFk7cYuWwMxPDd/MmkTK7mZ0d6rKkAaOdj9AXb4ew7ranAnc
LwHqLwkBrcNN5qY1oJAWOVzv2FERihm6uV8DlkR6BvrUxVfW6sua3G0qP26p4xGq
6ZtHsZFnk/Gpdf2/nx0vp1CH62hNVo5iR6utf8GfgivbDxZ0v61DlSG9l5YtLkQh
L8Mensh14NDPvj3uywDBdVrrOz6Zl2r9iNguulco+Ki82CF7THKpubBlsSII6QO9
3Wy1t2GtvnMxItkMJIGnfagbJyxAhmSBSgdZd3s9+i58e6cPHLD3unpWP54h2dj5
5wlHK+znr4140jUhA+A3DMSOn8s8LkcHtf1pcG+pYkItM/fl8itzyXJ7EpNPAdWt
1o/IjRwjXCCLErTwTlUbqSJPCqKcHeZSE0p1Ab57Th1q6BblYklEzBdBk2li7rAj
O6fnFS4wCF8W3KmB1GBpcwvkmm8/2UQCSzzRCfpzzok+3Gs4NbacpT7zgVmIrOTz
kmy1zdAT3T2/Hz+Q0I49ZS06uq6nVT6iiqiLy6+L1ILXGMUysL09fdt2ql6mPRmO
gCCJEA53pFefqa3RZiKaewtIkjNnOF/j1D15po0LdC9MxBsOkrrR87qz1ZJZn7bU
I3efEo3Yr3fs9c8hthEusVarvzU1DrsbGJgFFGDSZ9kbXr9O0Ywu2XEk9icwOar8
AAJnqvNQIUcZ6ZezbjcwVzVR5DufI3+9Nfy5vG1a0PDjWZqjSY+1PdMf7JP3zJYR
15AGSPx2ZjIxB0A3GZCRTnRNUb+rUtALe3dXeMscrWFq2wQgsQvT+WIBV52u+kcg
TZ1yUU21luwM6yT+YrhBL1EDh9kOosbzGsCiJ66azZdutCWDQ3+J/BaRQy+Bz4r2
k0wFG1rq0t1gddICUV6WKf9TKZGs4BB/64bb2jjieAEkXP/5B2cedievPOJtNinU
WjuEEjgQ5WBnQLxoFWRjtiQrVFFwRaGdKkFEvvpN1eQ5k4YYLSL/EKQ/ydAp4Bn6
+avkwXF+rax90NvjrrwlYLaD0wQbE3AVZF22zaAPE6xIvZvqleNYfb5OT8iOC/o6
oXqLS8VojElrSR2I3XYLkzCx+73wa165U5xyFoXzE5nrncp2qDpz9UsrcIah+GCn
u9sWM685mazPMQVyLsJgR7OTrHerRp8fCEva4Wg4AfDLI0792MRQCEcJP2+W0d28
AhdhFyojpw20WnOZ0aFuvGed43DkvrciSV/ZBz8v5JyOjdnn8/fDlujv0dOTYS2A
niRfZhYPj91RsFGyvSypYCF3V3gc2Nf9I60HFoC/UoyLlSDGaK2FpHAiOzSfY3iC
mxhCDsyJLxWNW6Y/NdNsgtl65FTh1g6u5qqeVtQtJD+nQLV/A++4yHEACFFkoLmm
JFHNa6Pdoiw/hOWiYMGyovnbOHWCz88BZKV3K64DmKYt5n//y1zIoxeMHwBDf5zH
D+ADeSPG+PLMYNjAgCZHGgpaoDwig6P0Dkr4bqakovBQD72ryjNjxzdS33vKSpsb
S8gmn0pyuDI3TdLGHe+gf0GA/zjFtvbl+P/muTL8ZAAxZLv7qvW+in70GebgFJZB
1qhytK7ps9QPIC3Gzv1vv5rTiWaNNYRmL5g2PxAp+tgOR3q8fji4/Qr8hy0VJbR1
sAals13NlJcePLdthGJM03h/6fSoIS9+Vj/s1/POwcx0QRw3EdGr0ha1HUBv+nnB
16gJFWddlvOdsht7uxrLPrsjnY2kQka/7fkzXCc62fRgnc90d4Jgv1ZmakIiXNT0
ll+Z13qtTxgz/8etjVnnItrmZDGWU9qQp/Z9T38dn8w/Qw80AN38Rrv3g7J1aC3y
iqnTbqb5BrHHt7ZVmwdXj9v9G7yYY7NXkU/tcTkIMDnuviS5Ou+/DxY2pUKBUA/7
1g8m840supfLe+iRC1NhIgwngTleRxp/y0Eduh/g+kQRubOpWO0k5i8C1+TPK8gZ
wrsW1vAg8oJSktMbuvkOCSFkfazRsOusMp+jg4ctN+uxFMqQE2ylbkGzoVPB3fjA
T5Z6afH9+xz6+8Y9Jt14Cm3Bp6jZ69WbxdmOQk/Pr0KQQLGfdKHiMUDyY9hOblHP
tjcszjFjtqBbvjrk8V1OIV6zazACSiA9DButb1R7HnBYEBu+PovrazScE4wtomds
WF6DI/U/ZWHkeIgGUtbTCTbsIcURhyYkpD7RzJTkvME5qgB5Y3yKr3zsE0MnAgDk
06rDnHFf8qcDOVVd37vhj7OyuX3nNLubkD9kCu+sbfxw8jmG/+0u54TcEu6q0La4
MIJv1sgA1VSJvSKEWEY1k81AFUEzYx/GiQKWN5JlsHY7wPMnFAjUN9V9nAH3bXgU
j/LbhSBMAiTuJ/lAxw2NpydkSTqsGvn7C4TmIEoD8dZzQnW3bqjZdFkkjr+kyODz
AD2e0YWJ0p52xWuzIT3GgVSaxaFal8T84wEkHbOMXVjusST6qljYDHzngy4v++fl
FVbrMVQj8bQnAM8jnT6IPfl62g5Sa8YuW408nfScaJz8P5gi9WpJZCYtg08HQpNS
ILb7/NeuW5H4r6ETtEAgXkY4d5eGI0dsVNPDB/qD2/hHlrHLznBr8BeY0szflW0M
FIe2x537/RjGNNgMoeXEgU0raEi96Ki4D2898+hJjmEOhg+yjC5fKfgL5/LFgv99
w4gBDAJHCp3meNlXMM5thKbWSoL1hSCbtddWnJVmMloOqJu/40L4vNin3/5sxGYt
URZjrYtImNMuEbagwEiFkcl7dY/bNU4KJ6MekkqlcPF3DUtll5z60WgdLd25UFuX
mpOab6gw/SCkVwdirkBxjh0wi7pAQq4gdXkKBldMiLIVCZZI6CennRRcRK6rWeTy
K6MVZIsbiSlacNyF+lY0PAhbkxY6Jt/Igar/Wef7K7L7FABp143poK5t+EmaNwfu
1mBGsIrSmtLsTjpAv844zjU2I6KKht8oN7jy4Uqr+LhYbjqaUxY7OPTJcH3pCwUv
G784mLnxikJuomgYMTjziZUXH9+HRXNUbw3Puo6QTKLbF3j0sQMVSXAhAwQVYuNh
48s5DAX/WCxBN5Q/o7s2k7yBSDJPo2G5upRx8B7/AgX3VTIgNQhgQh09J+vNNuiN
OLKgHgRZmZLPHhSyzpjYACn8dK4pPOWj/gZFq6huMYZnh7TZtLTjVxgf6qlrLwje
sr1tUAbobo7b2HgbRjuC2iVP1camrzkgep6sTA0zOXCe+NlH8WZ3D1tupuJFbW0b
xiYCMhzu5bGohB/tghJULY96253VDl162zuUh9L8cTFyjVItnhM+Cq2xb4qSDIIg
g1+ZOXgQTVjyxresA0uqqZNwvSjHu5ejOc6cQ70S2B7xisF0XWF2AMYLuNrvuC0T
z+akzvOX7VXI4TQwibz7SXLPOIGFMRsZlyxE0L8iRY6hhn5GQ0TZ9Og9OmttDeY7
JkJb0BrfTrRvfW78LArB37IsO51PTW8T/940n/zzDar1uRuDNWBUOXQUANPUsYa/
i4pC7IiTDnP0cQFv9L9Yvt1t6tLVlWDQtubd6feGHrPU2mzSA13te7lQIqo0RjXG
deqxUjJN3KnzQywJdbPnGInqUou29AqoxsLKgF9cDR3aW88KNl2zsyludjqD2EV+
oUnRNX6E1cnlSlPECm3Dx4dxc32GVJY0gQ4+iFNI3p8EwOAmtJRRGaApZ1tr3V2k
i1nZPcKcW3uXXj5fVD+KK9bij0/22UeFmpVk3FVw9+UGqSx0lhpWKseFfOaI483V
6NJoHY9bnPawWrsOihaJo9KxUsddWNUF+1THqrlT/xN2O8iqz49OYvzvb9H/AqHb
UClTRXR+Xz/TXR/WSINJBpqb669NgpnXwdYZm1oo+GEkEa54uNO5e+sCnG6rkPCP
NSa3yWkjyjB9lr0trBJfsreC+4eysBTbOpY80mh/leFltIy4l4KFbHkvy0NN/sdn
mRrITGh7dTe48lgbhMtbo+e6Iy/vk/dAA93Jbp8cfeRbACdciuq+foovMCiy6KMt
8QAhoZ7/tsSq43drnwoBocrYpOp8IpEMI+y8VFoo4vKP94oii9fTcRVmoclse9N5
IGBjs5JWq6FjUC6nrYAuhZbvS+JCxeiO/5bSzvNSR8oMRteD4xFS6klce+OKhrgK
uQ5XKaF2rUuxCz49ZNY2eal/C93emiJ2/3dKWZut+NeXT5mzzsTUhDEWpXN/kbnF
HMU036JqOp/f4mqxcfWNPu6Tp5ea3pcvbxcIXliNiM1uO9q3dxF8x2mv3/m5xUAd
cTgNao/UGSw+S49GaJE5n1aXV8tDMPxuNcX7zvFMLd9CIWvLUxJpWfs65RhIP0yO
FWzaOkW/yvr86iGJW1KbPv927JgbuSK5917JGMPFmbLvdF8jypa+hMsd3IuKTKvt
Lu2cIO0WQNISO63KGi+NhtZrZ6Ea2PFsibMrLkMj/KuP6cBw6MilaSH8VGGDVPqc
vliYee+dgWpEvSoysbm/lJydCId4yfiDziBFNpcFu56jKroJD0FbUAzUilF8DWji
7pLoOzkn80awhYX5CARtURpsGR5MCKfAxjOpW+wSzXvrp724L/e/JU7sd2CJZnzC
ReUXE1MqgzDUHXNbnfmnkh6t6ifUWy2E6K/XfMraayfTgBya8quWDRG65srE06MD
MYb7YwjWdGazVcnrJa4Dmkxf4GgNY6p3CazSBMwc3nGSuSqneDYGcfrqozlYONk+
ZiWa+drTTplCqk4gWZop7ne+fP5yhOQm99K0X14/u+f8O02Oj5N4Yd0PgUEq/fGJ
dSGfMc41YissGocJKc5XLrdn/W6ZeVttqGMYBEmRWXCN/WZVK4ImKQnWYK09nLBC
t1cRg2I3vfHi1TozCSoHc0VLw2LdoPEtymZ1WJ1RMBfygwpLdZczLPkSclt4Q5PN
pb2krA9il6nhObcjMdL7iVHM2GjCn3aMw7sNnSWmdQ2XhM7TSKXA7hWBWigpIljd
DqR7JyPd5o0/H5d/nQLMFsMrQEbYQon4uCFHzddJNO9mJmj4fBLq/jMjuWULFJGS
oBKWJeS0hwmxLdnDAKB+Sz27O2WOe+NcHkBPgsU0VexzLe7guyofru9qxSiLtAfh
0Pk4tUrfep5L7ZFISSycyV7ctv7smIrLoPoZ8geAwTtV3MBFRWdt+KFuQD1Rw9Hg
vL42TkVVRrmhOGuZ9VBMwGr7Uwk4Bc2HAtP4m3srzorHgMU2+Ed+hTc1XOhWrGwx
4t1il31K4Gd/gjEljF1JYRA9qGhX7btDnxVKtoaly0Pr7lGK9j0LWkI31bNYg0nV
lIM0PeDy6IIdDOD0nYsy4QnxwZQcJgMxbAmn1GjwtkWh9uA2NRLa9Cz7OyGo2Zgb
slBV2KCBInOPo4cWuRiG4g8En6VHsOl8dPW0qpr808iPsyOvFC5cbj/Xbb9/AUwJ
unX1nfm74ABC18vsOUKGJNIT84RQJwXdXDhMxkJbnH760TNveFr35eDwvXtAMEBf
jiJLax07Agmpd+6DBwrOiT3RLZ1PDlJX+s2unpy20roh04tnxoPDb7eeHX8daXJj
jKkkFRz8fwCpOVtrcShnvq8NRq6suoGEjnWftgHc0JCAh0HuRUD1jg2m5n6e0I+d
PqQzvyZCDxyHMHhp5GJm23S39YVH9UcyCXMKJThq68D+xrAe/VdqqTXSDQuUAkAy
XH6yAKkgama/VUK9xm2GXSa4LcRNmHo16hTAUfJhGPjmiTB8maYUGodQnaJ9dFzT
wsiDEb/KUZ0a8IhpTPP6AdFpRpRe6NWCzVFR/veehASPgPO88PKKmxwXK1RHF0eG
uXEbzkwMiMsbrDPpOqijf8o9SWGov559/3aU10QE6/CmbHAZ9ZWKOOcwYE7s0yok
OkRbVsmxQrVE2NJu8OVFfxlJ9gWNPA2sG/DPvaY/qjCRrXXqMBkGIXZ4v0AxY2vZ
SIBo+0V9fKGGP5B8DX2LR2x10pDsJ1G2MWNgbpwY7TGwQQ8LTwgpuvgFTlp4b+fy
qES0DBebgfa3/zCu7jsPkL/w2Y1Ptv+N4wjrOB+tqcoDZcvyM9uvUm/mqxFyFuQP
2vsVQQV7p2r3UBFurClxSSxJyIkD+h/XUH6ViEFUEEgwiv6L+eiUuX/8zqu2iCpK
qvwiNEiyy2/PAzmKfJEPLijQ8pCQpvGfVKKGDf7lgzu9nxE1d2Gfh0S1BzOFaucc
PdhQEDPEg0gD17apkJBnPdcQvQphj2jTa2uDSfR2mZ+AeA0oPrNdYNTr1nCjlO8B
jN9F7OrcoxDCjZQ+4/MQhOM8fnmdxnvBjb27bbYAHyPISkJqiIVOAkIwRmIPmGsR
houvLCasGaA2oP3hv2PenMtXBP2YP7XMO/JphpfcCu32O6zQtJIwoVSYlRiuXw2e
PHU2Pk6UPszGY/ltPENzRUQskl8rs/Q09JjPbTAXL/n2OqJv5qU8xu/moVJcz8SR
vW6Z4tV1s1E+kdABG0Toa6gwZQm0JWE/r49uBfiERRgp4PZC6N28og3UF5iAHOs+
aAvofJ4MZh4ceF+Dc3CYbqII6dVlt6xgGTn0185jG2rAam3ZCJmIdq/zqblNb3NQ
XL57bIFvSlfYTYe4jVzE1JB4liAT2ylbRGy9/osotP2OgiAd6rKrDbf2esYquGQt
yMkpuYU13o1ejSilf7AwcXZpuu3b8wESmGVGswpBNP3PhNfuh6ULdjtF7AwBdcW/
b9skjJwtl/0syGWYI1975yMHD/bck4Qlv0UqAYJWurbrFC9yBxqjJIWCjdGFfowk
gpbGhGa2Z1YJi+5O5Jeto1Fu3z1wOapMKg6+ht5Lkv87XDqJdHlrRoE9AfEIqpKN
bp/69ugerTIj9ouAZn593QdZ3yUXaw15e2enFa18ALtbsTx6wfd8NfozJdtNcXGA
25hvPg0Vanb/Rl2cQFhs8XBHMewxQ7JtFuNjib1k7+5MSPXvFqINovWN8c02R8/o
RaX2fAMfYll9Sszu65gb8uAPRsFFSsZfSKRko0IiFVRxnSETOUreEedKWLOznKgz
CJvsywwnIWOYSgKHfZNMY5Om2MpVIk+3WAnxxu9NPrrl8Dr4GQCKJCKRLJVEvnPY
d8QeyN2mlpiVLaFJ2X1Axl0NREpF1PwRTpjwJGkJmyaAlr6TYwXklLSBeOMd6/iO
v7qE1BIHwuX/LkNhAPdVVJ/KA2FvLik/14I9md8BNtnMCm7sxirgGdVhlxoaeR4R
7eT2PPX3HBvZD0uIFzdIULH0Y2QwOicq1xId02iJDjazO0Hr/V/gOhnGWMAiNgns
QBjI6Y7RwUgtxJhWnjMXsnq1Cp/2Pj3zI61zZ/G2W4aXVdyFR3dPVh4tceNzazyU
q7Y3rFOMkZ7dXrzCwP/eK5ZdOQvrqtFcDHoUXb4g2roLTfhqR41/FZsX3As+sk98
qreLVn84NDCDXTlLg4OqNe3jh7mSXdmUKQB8TwNRKwaoN5iZQI6nsutJZKHrSSwE
KiZhO17tPJotnTFVNtDfmMiwxjHYY5ozWj2YKySchRiLqcMjemfpPtaM/QHvaiHp
L3AU6HP8SzhUeJJRlKnTYRFgh5eWHch30i5rQ8pP4D5XPS6GuSmvO1Pub6TIETph
WH+OsQtJY7+ue5ZfBm8fKxnYbtcNZPp1GCxJ+4kvXfE1CHAsFPNiKEffBOZAZlyt
ls514uCtJV6NlhTIzpl6ie+G47PYLdPzdX+U4M74BBlabofIPmmpIzvT7Yna9Zot
Z/tvJ7/SH9CYycMtDRMt+dHau/YtpRvJUkS2pkZAz/1P1UYOk+a4RbAkWhp0udyz
nmc/pCO1ylRpDHL4ka6CeGVvcMlaOTU4eePNB9yZxsnGOL2Zkfbdu8ppHCEt8HrP
Yne/4CzdBoEgdvTWwrFVUodrhnvAjVRz3UHZXZUbXu8qI2rOrAnNXfsTE07J/2mU
lMWMuaM3rXK070BM6XHiRuhYkr2VQtuE0zmob++Oqho9c3c8n7W+9a0oU6Y+Yq7V
gR/wMQi9GYbn5B+4wrLwwM5a8Ouh6291v9tPk6lYkPEQYlBYqbGTiVuj81hHljDY
fq/3JLHwX+RAxeAbITsMXKEV3vlqjMWPoyRNE26+xXmlt0QyTD918PfeSvjKE8F2
oHTct/AytY4A2OZrX0Nv8s/RoCixaLDPkMpOgmzqBsnJU+EQmcJzIU0XPGwTB+sf
VQhgG4aJqqxYqugjXcdI7FNYHKRI7tMifnuK+OuQP+a7hjIRi5jsNOX+Gpl0sUsp
a9i7IV/K8dXR6L2ej+YsBIvQWtxD92L8UHfiWsua9rU1dQO9Rrw27McFx7AT9Tct
z5PHGBe1PLUym4ShlYUhisewzAwlEDAutkQ1nLFlc6bVdvniSLWa0CjkdJ12AjmW
SO8SmkCfHQpvfbtwCq77py2meXt37mw2cgnQi/An5dFl3Evbd08Fcupl2tzX/pCX
nmHzKfZwoJbucxb8elu8JUiFir5bfcUJDMKsYYX0iIi59XrjTBUQf/9Cc7N7j2/u
bnBCtqEaLo7E3WqWoJU7IIFQ0X+UMfzl8Cy92ho6DZ4uACXh7HtuZFX/a4jZJTh2
UNjpXz6t1vwjVqI/Nm+jC1PpM8imviK/pBEVyTZpAfVt2oxloKE6BEdWqYNvg8e4
Tu8xw2QKDGu0Gk9oiHdTBfuuzzGy/m3q5KDCMRrQa+0Llx64grKumoPsTQToySSu
WGpFMEO6YC/NzIM1RzZGiUbbikByAr8aIjf4qXKDqDU8ig4KkKDd9Ax6p6OKlOAM
uqyXsFonCpOZA9hbD+d4Jw2o9TwjyUQLn7K9s4HblWWmMJvZfDTNlhBl5Aqq0fn4
dWJZWLSHEvtKPGbwqKJX0JwjPsLeIDY2IaFpfxESNTA35SpkhRnR3HZ8LgOL07/Q
3pIKGtmzOCzWFMWMtbB5XTKl5Vp4RSFR7vyZxTsOBgDjKhkJ+mS0JLvtNS0awwfd
pMumcTqTkgsB31Zp1kPqNMHVWOQDCXp5jpXN9i3Hy/u+kBO2zovOf9mIT/bT0K74
fYwQYPE2svZnbkey1+wNIVhMcg27bUtDNblnB+NmRL1xX3f+pDbHU7F7Cp3RSfBa
ZMEl7TX/drJ2HrnKdKmHfu034ZEQKq0nD6YGNJGZmmfMUCBMVkW2++Pzo7I5voeA
huLDWhX1NwaoP3ZWu5Wq50JHZuCCuNitHEDO340IwxksgjveJei3KsRK+48SwL/x
fGA8fqywNiv4TRD680VDM3c1/ITRv/9TBCpubIHLIwGZgSUblByFP5UvjH/7mUdj
xGbuCfRymiOr9hyRTsWLhR0r1R+oEdIQJ+vCVVlRN5YKvc9tKk7RLFWIZ58zO/oN
ULE7dzTDohIkFvht23+HaVUVtC33o7k6R4mxjP7SrNZAE0Q0+6U2ai31ZWS7fuoY
5huSdHwvgomxfd42fIn+CtebB8IhEdv9qd1a/qqTZyBODHj5nt9IBSaarpwbnutB
ajXbcILx0QofGCoxT7dP7t8WqdXaeze3xhI12HtzeZqdOXfzJnkJyNgA7v6NvBay
o7plVOwA2vgFo/bh1k6UXGbsyyBPn877Mmex631ZO7E4BU1ymXpIjx/KgjJM2ncK
cImxNArz/flsKItgSBqT1/3a560slvfkjW8EKJx+gf3QOtn8VA2vDkr8TN6T1aie
eMlbSDm69vfgYCBJ6aPYRckBL3ZA8zRyZLk4rVFfDb8yCoRFUh987sIQnOJwH71f
FDTfkJ5wVx7qzgjPRAkygl/M980v+gkBx7HB68r9wZuyv9Dst/Uy2QgBnwgFBJQW
gjkvDUh9xrIegbv8vbeGnReBkx93+TWAWEmK3tt4MBHad0q4aRzzMDjPYQW3cXfk
XLKru1KJq6/2biA/BL+3JTr5EYyh7MJVX/vw7jrvnfSi07qhXaNjLXOnAHKE8Lv0
b9l5G196stNXbPv68g7PGE9WU3ZMSIoN6Cxe4kguXZXaBcAY2L4tnW8lBCo1xK3c
GMsXlFPhxYmj1zgYh+xaHPNC+wyAsGL8f22iz1P9X2g5EIYAw6RIW0jeuFrxb6Kc
+nhZqgwb8d/0FX6Wx72lOdG95j16H6SrunrQteAldIQrNivicSFrpeL7hJTrXoeS
kUf+fDfBshtRJnejpMjex4/2tB/oqHMu4MIuGXIEtT+NTDSwmXHS7lznYMD/1Bae
Qlag4aPq/qdCRsgYZ7ofZVEJxBQH/W4cZTxHpR32w8EZF9a0vm0U0pdDxxlmJjfP
es5X6WdapB6Hda6gyqogzSSw9Ynv0qDO6gmFXvnyCNyuv1PTsuAdT3Ph3QE3WFyw
VjX5nkD41FdjCZGciDqUAvESVSxLWnuMvTp01qdtwA607TXej60Skxv0na+trC8J
AO97+RdIVC1eof1LNbER11pO3neld92Fop49+CmBrnRh4CxA1pwGsRWMCvKL0Bq5
BsXCZ57MZnZBuo7gZSqu7474LR1d2F90v84OElP6tbPP1BvBtca2KOShApYs1LpU
39sNfLSiOcway/vvE1Bb7SbtqDqsn574E1BteLX45LvGK3sqIIb1g9L7o4WcKLL/
x7nxhA7KzIHeCDkwGOovbPYteA86qhj57eexHC0ItdcqN4nTtFVxEjVqd9Ki5AWi
cE2k7VB1c/BocEcLkITQdkZE5BxcnqaPAsSRZTUiYb2SA0Wpj3LjU1HGEJAUyQ5R
dPS9LkSJas0Ua2Xd9LiDjD5icGb1oKBydW8XGUQqzGqEtKLdS9Gcr2nln7p8XYi7
m9nT9rQFbyGe9x556ldCtG1+YMduC2XmGZp4Yf36F/WUGLeHLjAaRjmkv3DNHCcC
4s8lAt68UxvnI6GKbL9xROSioMM81WxHI48kRAsTb9TW/fiV04CzqdCCSb8uwN3J
nHjyRnBAQCIv2lFH6krC+Cu7Z+x67/W6G6Wa4LXSR3FxDkRWBjN7gpoP0mIfeMMH
MBq3Gcfgn2O4Y57PJSd2SJKn0w/jqB8DYssBt0V0OrbVoEZ8AQ3cx4Qa5OkGttvv
g6qBIx9JyeeTgM3STk6EfcPVn8SPbZ9VCp2pZMw+ffIj4J36EXQDToYv+MYDrTTj
B4xDpp+KTQmTFG+j9OKPVRU2uqB7WchBqYjcgLjGQu/s4lBTGGUyOtNXUPP5/4VR
CC2JTfyOMBhFmHfNV9oc2+V1ozks8/JwylDyssTwc2LeNSa9Qtj4rrXHT9DjOHYX
SsyKDIZ0+jLHKoHFroRbsqpDdTI/OLfMfzVQmJm1T+KXbQ1CmoAzlUuwO7jz/nie
K2Kuv5eqNbiN6Bz4RS3+Sw6cUUMq5dOF2lPXZ7OZXh7kNbKnQd2GgsOBrabbfjsd
fgQppxiyAZnI3KyHh0pr0zjdCVtOO5EzR3AmEo27xnPZBeXaz4Pue0/qF++pIalF
VJHFI1Q+OqS3oRndOQMWVj2ePj6AWCAwPVNQU3UNvR9rvBSYYU4voVDnVULo6Nbf
mM7XeYxeJf/giGpAM9ufxDWoBQmEirQHRnN0jTraoih8kClyaqx0UodoUwMOgGOX
nmEOGMnRYRQl6stgCIisVSlzzPGHknB8DEPikpkzgWtYPeL8E4ZSqKrUwMOSl0qQ
VsDo2QdCdGwKv0HCVO2f/V0C1E+a/t+ZBh5jAuSw4ySXlyTqAzci7J0LtjOn9i7f
sW+fGUk1pH1B/QZlt9J0wd/BMjyGW1gbezyQIbmLRdS2YN0pFnUAkyKEzS2O6n7/
h/8ylThs88GKDen/kCbawMk8gZMtZyO0cFYIglWjEIW2yC3OzU6IyOd0g7DR3B4O
5bDOjpOrL5+z6CjO0dE1f4UTUNIegO60+HDSALl9vMlCItmap0ROn1/AO3jYMAYA
vSWOxmxc6XAA87daYSnfgl6uB4VCZMHA/dpC2kOeOQvbR6kTN8MWhcxX1jJUNgql
JfYoNQ2NER4pni2dSJirNpcrss9YthF3JIsY+Oxso3ERBChuQlTnhNgiqUcClVmG
K8kPew9tqMqEXKdlYvk2dXsNH8XsTJ4N+FxLF7jxZqBqoxNJMfhh6kblGo2bKwR9
BLxbElcJx90UxNS24A3xW1jtz+U3q7kcsgebft+eBF7qvgw/yIEvzkPADjCnmGwX
3/RGOTx5XEeKgLe8tZYHOxW3dT/5MrE3iUXL6Yfs1TpsJPZccrTtUcgCym5/U5AK
9eVqy0If+MSmm2aFotQY34L6Hspp8gEA27HsSKpqy6h55Xy0IyoE03CFfcmfHwmQ
qpoAQs0gCJZ/hK9EgiwwOLNL3nOT/vScXEWLjhpGzPMyY5t4pZv0ZfCj8qw7Fa5O
wtbmHUDm/ohTr0O0LvZxsqDogc3J16ApsJGPE6HPP6lOrGGpo8QVp3Qx04RmXFkf
imLLrPlUfUMa0/TiClMNowJsVPM2SUd76dkczf/iSeVal4J+P+vaO1Bn95/fSeOV
IQqWQ9CinrGW7z2UnStB+R/OnjX669vc5eipN3twduDC1YQOI2HkWNKDkdDjSxcH
prkODXA3zNzjN+zhAX4NiIpJICyQD6o5YoKI6Adxl+/DztoHfUKI19I7CeNkR3qa
zkNps4FTNF5CoZc5zuxAw1pe/PCFIWGezO/wLAn26+YkILT3anLecQvrzx2+y4DR
4I+ZlN0IHlmmROzmcxY0OAI2iezKJCHQ48DIX0yvplZ3Q8Gr/iLoKfH9qd1DJIpH
NXmY1QVQXqY1nXldUsKNs6MOO83sPRcGH4qmGuvWrf6vKFX2qFLBqmC+E+7TQe5+
vHDTU4jtrJ9NcBDbVps3HNoh1jdvZQWx2UsTbuDK9ePMJ5GRLzn3/Q8avg2l0xZa
oQ/iluY35lFWylmj1fnNV+77beeNi0Gb6r7LlAMwkn+l3pgaRAWruu8d6NXQXHF+
TuTBAIBK0cwYhp0O5q7auvAgEPhoQ43opehZr6tpwmdP6dHXJ31z2oYdqPla6JwJ
OK+f7y5txoXieTrssYrWlGwR0uBcwtW4G5vTmjycD25CQ5Ccrcl8W5QFz1+e6x8q
7H5xZB4HqFgYCs4HEVzz+dKmBHSKTF7i/bATQgXdJuNsx0eWVSP16l9mak2epXyN
G62vhN2+s65xGjBD3T7IBtXwVEpFWhH+mgV0vUG0CEariiQpM1MIFCNnALCnizmR
4yZqI8Xdxhs0qr/TTIdGEGhgHCYQjJs1hIKpVl1s9O6is6nPJJoAkQ3cYQh+9Tjq
6BIXzsnSJdyn19A1AUNR+kY7quz1jWJQ0In4ucKfqRJhpvsq79TnYrqMjMj6ZBML
aZ89jKPH1649BnLVOlB/KbrNSSrK4uPHtEz1FEbv3Qb2SMdE4ZGPQYRtXGYKpn7q
1ELSmTme9yBJy4zhc1P53VAYKPpAiyYbQMooOdaoGwPIAZpc5/c9TaxKE+Em2W6e
JzNtJQBIIFudpruOkDzek/6/kZlujQcW+FB9gMT46dm7BSZvUYppm3beWUh7bPQf
PWibzVS/7HheKVpJFilJQepF3AHgrLvDc0tRENIQyehZXq24ShJdLUw/6o3aZW7W
/okwH2hs1TwCbl18Kx0gW0HFpPopFps0fLHwKKh7QpErfF33NsVxoZIAo0ueIInV
Olj5ghevM1zizYXXK4oXxTqLjmX/iV36QkYEe+CqMQJAv8pmL7fn2PEu5BNCIk0M
TXn/a5PnJNh1nY0TndKOUZy/cGqQ1i+2tEYVO9YC8lKELRgTyqdjeVyVPeHKP0TR
6lMVrEXKhvH29rgmB9UZ6O/6a3iEGSXCyV0wO1OxwFGxAvbte33d/KFgjiVwO6yS
1UL18hw1H5vjne8MDkFfhm7Ypujo9nKZ2u5/4gy8pYCh4lHJO5cEpZq/r5PC58N0
9r389KwbBfj8sQFwhvDKiZ+E7f8Bq439BraktfpmbOvU6pj2FNP54BQiueByclCf
jOdrrEIL4ptuxwLJOSdR0kqYBseileLRcKN1gec6II5MVptFGbDro5Vnj3BIyYD8
Y7mX+jEkjpVHd0S6kbzqYRyukAW67sDE3/3WNbbYtmHZuUWmXA+4KSM6QeIRgC1y
3vsR0wRJ9MnncOFCYms5QqKR6TFdQPwh5Zyf7QPFD2gkpxkKfYIyfrkEDP0A3ADr
ZLHX65sOomBPZ1xpx9e+AQ+N2svkn4tdqSzh++NwcXLx+FFKHFwJd6//urO0uZmf
0TQKp/mV7AkG99m7Bwz1d26C+oroO89uOXEMiUWlqdpY1xDY4EZQGqo8cQmuMc4r
A3uY28D+Pv8naS3vYIXPsJbXCLrdjPGUop/s5xuDEBfawz30JT1PW7oFdgH/+ZPM
J0EL2SSsuWpi49JsjfB3u7qRJbkq7r/d0hpGfyEk6w7fJUxNILW4h37HQtzgfthu
MDh8Rje6rYzgQ048aW7UrmiLFgDNjKCDDeCRJDMKeDpVlQImYxcgK8vsUUnfT19L
a+EoPLPhK9Ou+NUxeDB5HqWiUsVT7ChZ0fAcSaeNFL+hLr8vFZiew24aV3plkvba
b7yUcsKS9Z5dn05zoN3McbqfEmoO/Ix2yzigupoqQt/IeECBjkE8NRFPzfoDPoW3
ryozcbv2+XWp1POTwvG73cjC1RkM4V/FzaJjdgZbNr9MjGT/VN7E97soZGXJ+DG4
8cPtM+AsXhYs9ccfQSb7EDV/gEitMdy+/Ff5De8IJoc7WFnWIvf0oOm9y9ACe9H1
9wbTjj+7IrXbbZxgIcQGFxmUG9MqMYxkHA4+qa2THLoOv0Z0gGbW2so4f5JU8ggH
1EqDq981/xThE5Sjfjkh/3cjk7sp8+ccnloX6lL/+HDHqG0C+yNzYjhIX7/lCcge
62mxWUrecO/a4GEH7/UaNhmVGAOoHKFB8yZrYxJ1Cxjq42On2elCz2YGKK8eende
XWDxzqGKIOhR6fBfHKpHuq/rSDgvv1pLK+4qNULh4bX0IYcFm86tNXL/gkfPdYkz
KzInAprOnkA1HWuonKQ+XHdNSfMmjVRT2HqgAi7Pbdb4HOWO/5qKJT6N/Q0kr+gT
HHLdMJ9Rv4H7x988DREM25/XxA9wZC73ZalJqQ5tmGregvdzaFGBoIHXp4lj+6EG
gizdkRTRYahoxYaaDgZT5RdSUwLqRi4poErrNyhUJJ2cCorDcPJL8Ugmabz1R92n
2+RYYWyERctpoSzsM711ZLY5cbhqQWx+z9Njux3k/xseFQUMbvFYlgTpEo0cMff8
aC4RaFqcTaStz1mIAcwp33/KkIQmP0rCXMGK1HfVTP3n1NleZcX8KXdJFa9SvluU
QAxuxHcK7g8srU76CQFPAL6GWKEtd5JiilM42SbRA5X3e0NFTXY9EUPj4GbXFJZI
091r2r0Hqa/oj3C32F6Hs8l9p65qapQlb3uihh4t2+PFIs1wKkThCARAzwBE73p0
+DdQ/qqOyG3oTMnhQxik6hqeOfDqN5bjhzfaeYV5nWhjP/XrFcW4Xc7QhmEb46x5
7/nNLx7O8K5ptnDOwLLFErMYKH/wx9PCQWRExHkRICPQEjoAfpKtWHIFpb8RoKk0
DgIH4a2ETew/LXAuP688sIdRMo7/7xbX9Iydk8v3IbYtmG+naUCQMci9wB89i48F
cT4d+MVXSz914FLFMeURPJCgWXIVFVBF0FACiw3NaFbgNdgaq9gg5qEuZeNIwNK0
m3KRVNXOpNO+QtSBskoHJjf1FJ0zwobD9MENcjcVBXH328Jo+CnmOPzvXDyow37M
M4cI1rRLbHXboNnLtxq9OR4oXK9ozHXkRVnMQYdyS8DNsTwHtEuJcolcqMk3xi72
/IcA7uyjz/lEt3U1mqtMkSra9E1FLlRyMnltLld199GTYmLI21bhPlU8jYIIHGy1
fw9P9gspwyBbghDrK3sP9XdTZEXOhv1aMa9072I9/pWnPpAFBaU1iL+pRUJPV1xg
eZ2NdPdTD2PH7CEcs4bJ/UH7ZipvCBmkyViT5SScSXNlhhJ0SzsknLdBwEEKdiZh
SZ9cfNvcFUWEjmWpbDeNsXMHZrcDR2PmnOtOuu9LQ24OL+Bh1acFd8P+mkHH67aP
kjPCdaw1J34mCQwWqCU4zUJBHJ/y27WJItx+VzeX3qQAOj2gCs+ZCLfprHHPRbTV
pb103Oe+QnK0JemT47rl+eoh3kE0N/fbRXV6YHTyNH8JXpoN14nGBQ9xjP2e1oDb
EokXJybiDKg9ga2lO48ZCXKjPjLjbudTbKcD9UfnZKW1ee5vZ2STvSDgp/SKGARO
CaPCQCRswDtCVtA3zGhkkiRbjPkyZIw7l2f0TQd+Z/qT0PuiJLCrtS9ID8BsyAv3
8HymFY/AaliZ/jLsWzgFf32QvmP59GyOlYtNvD2dSAAfQRqQaLGfMuWk+OS6Nss6
lzH0iB0HA9JKd+FTaTXPySI9SQhpHVizZdpS6S083MZuu9trY4DuztsLNKAImMAN
YnUUZugTIrVk8uUskiKrrHtlsa75zYOotDHq+Y0im4rPiGvCc6paOLk5xSkH8p7I
UpQT0IktYux/su2RAk5OCaGDggZTxV2q/jtqgqYEEo0sbdY6tNxXBGijKSbh+rCy
9fCV7pS3r0A89J12sJ4WVFEQ7qk3JhEKFEXOmJTX+eH+pl5vLUWxV9oXbs3yjHR5
06Oo2UhMfdMC+JuEPRlXrS97eu3XCe74N2fE8J7Jl2mf2rSmeYRQ/cWR05m9g7rU
9SrCAjBlsNvaeRLCKoZFD8DQgERQdsoaNqJ6hAOU71vLdb0ZBDGTZDg3ZVdeshEp
cNVQWQhsoix8CKTA2QdVCzrNrNdd966AeA3PnI9mnmz0OinFsRJ09QsssFerbXkb
xFWciATIS178VDPsKgaErUWfln9co3DPQaOcOGspvlsnDFFQ4zs4uWLK7920zhs+
OY5twdo/GQT+nvk40Dqf58VkKe5e52HJeo7dzO3D+K/jpFNEht/nz8itbaCfFQzc
dd0OrVvriWiFYUSmd6jAafmzVjKSvHc/FcmVy+54PFjyWW0U9CW8FrNd+9HquwMn
kn30oatjak5S3on1KJDdYMjPIu02i0zhVy7Yu6GARsyxORm+/Cwlkf8kgAumfmEn
O1xl5Njt0udz44f1gXe3oXwoKfeq8FYm5+DsQPXuXq0rpAnmq2hs+c2QuQ+VuEEQ
JdqDFd1Zj+M3bcEtM418JNHmF9fOXtbO192sEe9mHRvKPrHMu/HvNfJGa50garJK
UPrIF6bhSbKtabQAzus+U/K0WV+gvUp4BvlT/nfbIVMDTLzK3AmdDQM8ujFB3VZP
k0K+eVEMy8OU959AvCiS78bY4X4dS2Nw7SMtNHSYIAGkqTC5z2DPxaKI2fcQ+V+w
hBnCQkjJx6Mmc1OtgUnWqKjyPQUhfUfq3CBpYh0Lqi1QkhnnT7pDe3+u0TFhhACe
K8j8MWwFATPmoOh05cOqvJjRvHtq3jVhAMBMtwM13FqFwHGbnaaEWBm0cZWYKuNI
c9W+AFxagsWpjwYq8UyNpU8Ws3TQ3P5KehRONT51ZgsmwUJ/6B+lJ9R22usg0TMV
zleyszogxrJ2lYo9WU4tcHfntzbAasKWYEHoNTRITcyqfwyTNV8shjWPq7tHiO7t
hnKbdU8pWQyLeh1RDEAkWr8HqQHeZudVUVtzokcTcz/WlCyjIz5Pl1nguGUXMgU4
B9Lzm0rSu/zQUKujYvX0a6YKGEj/ya2kOTiehXlgvOfCozaVsYFWPLnUQGgh7/5J
Am6hFpAmd8p1bDCgKuTwXXpFb63SGmPb4TyaVI4coSiSkXMp8s4bhsoYEtyJSBlo
dU87Wb2034tmgH2Tgch7qhJGd4gFzkTaEmt1DrJtqEOrPLSXXVe32T7cIMcEwmtv
TAt74SkkuaO5d2a51Ad97yTof2sQsoQuQIbmICKzkq8IhbTEr4WhzISphJ/IhrMW
mjieozGsSZ4BXVFL9XqHcukhDqllDGlKpRFKcqPhza3ArPsZhYGQ3fYz62Nu3rqK
yZ8e6fD2usOYXxWZ+ApX7lQu51cW2d3CZ0ozutzHkj4McoP/Fjxr1rLSy/DjUzt0
ZkPQdAzEA6uR23fNydnmsUigCNJPMP9LNd9D/cK/spJbVo4Mj5Y/IdzLOIqhyIcH
43RLfAUKMVNtbDhtlSQzkCW2zptytxx4zrmA3BTiA/FkVUTyXzauBUyv2hBZ51H5
PjapFH/SuMYko1RnH6SCztf6HaoEYty6C0laNqs21G51HTX/Hm22HJFRDyTzyxmT
T4mIrFT/1bIXdQGL1PG5z+fwy2cjadhflht20miRypVcHdvkYPVBx/GBmLAlH87A
p0zCvXeaBPJPs0QLEXeg5UttxOH4zNGUNS6Orl+xWTqp/orGtgY/GhkmEdt4SaO6
GtnQBaFIuDlYOoGdITd4p47T3zzBAPGpWYHMxCVYWqk0MRitA9njzpdTuJh9/AXP
oATSEo7qD9KE3CzNI6+W6IQhi/svnSJDtlJTf/u5E7+fclfLVUd0Y1LX76XWWMa8
QMWzQXtsPJUu1SAcARvHI4K1q4zytIZXgMTU/tLEGG1kzDK9HabKUYaE4FAk3PVx
WOMkhZJDyrY8+WlP5d+HNg8iQZpts6a9sZYQUkyemMiloQDQAuImfc2KA4Ns3ibT
JOTcwoSPXLNS01Z+ebMG6zKyN+taJwPuKXgrvNpqGuATcQG5rrvF7gFKkcQdSEV9
Aom3+2Dzpza5558k7c4//ijjFcqhuSB+HNxTgdllizbIWmg4b7y+Lwydjt34pT9m
c7cUgZx3lqehSSQgA+9Y98c3MuQlNBeUQPWrD0EMS7v5JJYYiGC8vTwwUsA9lg6z
7RBozKY9OSWXGHUrTpU9vocqg7XVv+DHN3X+zF2wi5nWgOkTH7NRqFInXwTfSywp
VCGzdPiKNOoXG5kZ9QLuVBGcGwBpt4wmKz1HVfMDvoIAySPasXQAlLW+1rEWztzQ
9PKLJ3r/dX81QWgf5nytYpkelzPjBbigV760Yh1SkyiBcbjqJauQUrrwe0dsehAE
5OcesqW/UB+S+5VYnXopKzxU8SHM3iGiHmxqU0hBPmxDhFK6nTDvxDxrWKaAdgyT
ZhjHDcXYFfZm1ERxlaBVfMgwaTq1iftAyg9iYbHWmVIZXm/viIXopvdSZUwlNcn9
6yESPDBhHhvgBMaIkTwi70qQSXM5K5tNj6lTbc0v25ILYrJMYo4pQwVE/FKwJf8L
tjqrVTvwee9g2udLgmASbxMdDKKE2ZIQLtOHdUWv1UQ5TC0t2TNlHctLZyMdocvd
T8FfY3ay+UmVLRyxRtsDPoe9qEBrKU5fPlXgVWkSYkMZEx+qM5YwriRu0r+jB2+t
/dD/R3yFpptKsDvVcAX5wAYwN20d/ElXF8nMm3C2oiZfxDKKzc3JhUSwkrIUDZnm
V+KLP7NU2Jadil0MMDllLGvqflvX/VUiLibadcS4ECZVHUUAyjbL8hzuaJCfthoR
3pWdZmuK+IQY2jl7FGl7DwONtlkJ0ym16gBMq3KW5JF4PG8xp73j/TtmGYQ7XmZD
mRnYPrXmdUh2AIdZISe+AfGGtsa4u+YEnm/CEzjSNrU7rp1ag2TRYSBVyHXxVI1J
NC0bnbFeW84s20Vh5fL6vzDv12y/GeVGHvEv/+UQwdM/Sp/ejpMzQ1CRVkeH1MHR
QXeMuf4QdBABLmU5pEpqySSupRAjU1ACwB1wrhEY6xZMNxyeX8Z4eTQo0p05fAhQ
FEiXs66mwt1BSN48J43gBd4Cxz2ii1Ry2ekRdNmsyOmwxWOhTkOGsuo6DcSeV90b
rxLzb2FMuRGkY3PhiOKrazWcgJBgzlblC5kCr49iNp4Sn/SsqTnPAzlp9azldTA6
8b0l4rkM72fxv6HJkwXOnYzSA1yovmDgODGavXqcFr31gZEV5NL5lieDAV++VdaD
XIZouZ4RmParSrtJ6bMrwONjzHiOb8n6Bk1VVtc4Hi+qfoFN21mvWLdL2wLkan14
kQ7oqPandKz2gLGwC3D79l7d1R/UonmOVYBSjafeFy7l/IWyGAcCtWOV98xEV+zJ
Mhdp3adbuIfbmhHHepUPkDsGz90ovLAAs6BxZ9kZP+NxxNKfJ5z/u8bhWDweyuIS
oHsNoF2bH0KRhl1Ac0OJN0XuRl+qzbbLAz06OrpJv7rOmIY86KHzPy+1N61Lj882
tjMvf/FaJ82joS2lOuZrNkjaFKui3DR3pxmeUnvDAwG8iuzwcIEBrG3WNHKiu3re
TkvuXPKyMcCmAfMBmLP/vfOLjNUs2cVGVkV9tUc7cFifXbsqAvHP2NyI4UiHivyE
pobzxP8q/bSbTqBEw6P2FRHz41yr/yun4tILJtSSL9svHfZ0Rc/O0/CE3nhC9ENF
ZeqMNbf4gVm0PwofF4N4Dw9ng7t/KpP7bpQZzb8e7MiHOUZ2eaSzp7DGMrW/p+LT
4gYuBS55gTIYUAA4Pvx7Cml7hs+xloUQvtH+prQijvC1nfcihnXVewuObFClsPC/
o6YM+m4HtIu8qeDWw46JiovHQ5XAHn4swXWAFCGZsMCftmS38RcOs4nRkkumBVPo
Tfxa4dNAwDv9PyyAShyKtDbyKzRAj18SeAh1UoPmpFnHw+c+skgOk4HcZAcXjckW
djBvvG+pB7phzyMoBSvKuck3N3eKqur3Y1PL//rRB1UyqlCesRoIwOCVt6vDleEe
Hz+3DQhYlqmnsaxffOYxa68lWmfvb57pWVMkRr/hDSQ19kGgMV7EhKBugczWJYEW
LXYi8cA0JwR6Xk5sEbEhZ1GySyoDNvrMRJREbRWoJmjKBMGh9y7sciyRo37Gd1Wp
eYguYwiGFtWiHW/9xbBy19dA/eU+BapV2TAhHsrxEujz6AFDrTB3nCiVg2bR6b1p
59aFk7heRB8LnqRZm9HlcTVXS3cPVhCMF+rG0SNYbZiNrzxvO150gVWODhdKqSCJ
5ARwe5nWfp1CXz497dI2ShyIv3xVoPjVR6U0MuCKJVHYqihz8OMGDWCPnqqY/0VV
Yru8DReQF1RBzXhJ1elKFLlkg18Wib0NoaeTWbofuA4wiz6DYTjRHwwTmSRlVAzx
72Muedru47WGVDLA71gFK52SKtA4eTX2BInJEn95O8LjvZctZ65lNdsmYmp4kxJm
KlhxVjL6o3/ZeYgyGB3LjIy4Hbzi8mqEZelonzjEA+/4F4PdU5O41nJJGN5LaZjV
uA0XM1zoTuI50K6frnqXm7cBpqDd4NGYV3w++JRgpRSSyIJNWFryzhIrLKkpsSrS
jaEwjchSgEvjX51zs1hZLzNKaymhxs9r0kKIAsA+939NsncA4h1xAoo8XoLU2niM
xYnLhKE8iCbhe0s80OWwCq4rkvDhYQf9MheK2DpOxI2gkTCuZG66SNE37bZWotsS
zF9HQFe13XCGSWF3cdFmPhvglskO/X/xcZ6I+0rHSc0yw7xdi7KdhZJH9oSXRfXq
T401kNB2+Pqg54+3nuYkyhA0E8mHuvAyqE/deP6tuUPMVoXTjkdBz98oKe1aS+Kq
NrE1eGOF/+zpv10FnQ2yxjxHWC+On760/GAE677AolK7a6rGW4P4xJZg134mHrnz
xmibjVXWN/0pmStccFuuK4tbbZ4ca4lur80JBb6RjEdw0bLDi+WsMv/1IkPbcPpR
w2H76extBMmWhiEx/dBv2No4CB91GCsM4BFgoXELnlPu5oc0RMGmy6I/dpQMQagU
LdE+l/wjvsIvhM8rKMJubk5XI7urzQeaFpuwGRQnH5VHUrkFh10lLDA10yKGRl+s
O491UjuwLKMKzzXQf3uvwqiAcC+Ky5Lgp/hvx9iIW/j2GHigYLm1wS1Ns9CnVV/S
0a5HFUM8wTKMeWUCdw38199S7VYp6UjZ3kZG9PlX7vxLjyLTd5/8E45sGesuzZGu
v+2/bszRMopOgEYDQREIiYAG3kTb+z2HZUix6c0acrppByDNuaN3t1Ls5NPaHhXA
JSVzZ4Eq6Lh9Z+rt8jP1hiRBIzBX6edxD2RhVfFGStKwkJVHZviQUjVFzmJLQC+G
tWZJ/1MPUoJq1D3RzrisT1drvD4BoJ0jxi1IwdJo8WiUKCOyB+76Lm7t0pWHxrXP
pmbcc1B8EQ5yqtmePD5XyeYAPlhifrSEbBTxyfMhcheCWyQzFGMRjtlGexGHbWAh
LxvwTXALDxALIqLCxkPD2mInO9MvbPPAAop2Bl1npkycFhJrIRRQ1Q7HCDIQguA7
2JI3fz8ZQ/S9/msE2pN6A/p2iQ5aTjgBcyCbkNd2OGhc4OE2oiLtidT9BA0We9h8
xtbROJK8Fj1mB9ZVkUCOvkZr608Bg8Yh0Q1/z7qRJoZUdV02TCNuUhgBqEOVFoNC
+6g5CSzMkUyFr2VX4uJLCi/9yWE4rvaT1bDf6WVSbSXPBbqRM7yxT61bc3CLzv5u
bwcbT4/Z78oovZs0d7CGLitOXCr49vjsLsfulvrAgGLHWe5996oHSJgy84LgJjuk
VktFiceazWFxnkumuayQ/GB+pULVtt2sdylGkz5Z93w60K8DEuSbDyh6UIYOAO5j
dQAdTuvcc2kPkeHotf0+LiNQpKr5br0WwAkG61T2szi00NUwp3IZoq4rlXFE8Ue2
bkiRTgwsMBP6A9S/rtO5vH0CSEsyEtrAB4BPtZ5RCWslMkE9WgsvTb3vQPFHuWVe
MetRFdgtksoysejg9rAC6kwib/T3CL+1mzCyw16WDcPAQcWf1a6m+mZSjmStERfL
i2dVz/ll4fAnnQ757gQI5w0z9W9RMIxav01EdCaWr2JKHUAOj1iblF8Wzx9WfA0D
C8Vl59s0/JNFHSntvN0F+/nct+7R00mipU0JIOzhWXj50AG8WXzOC2hi6jnAnAcC
+OKnGDGBVPAzMS8T2PR67b9Gfk4BvDX23jTdGVD31bQh3ivxb0BXxEo6ibY+sAO5
T7nDcLFZR50cjUqfCbyV8iEg+N0umU5uPL8PrEitr3tS+6SzjVXu2shiB8X5SaLJ
QnbZvBfBeEvb7VmFr1LAbcr8tC2TORF+IhPFsLzlVWrbqtybB3ggWyVYSox3iEQV
q9LKi/V50qEAbbbtkv6hWxYDCEeM/lRfcfhjcf3/UcYrkbKDLX/+AzfWjQNbTu/e
RwLWRYsF8oQxSt3H1UPSxB7OH7ZTPD1IstRCof+YXxq0Tn8KpkjHNLJedhomZ1n+
3V3eYBh2xFlQrPjJ9L4Nrd+oSbvkUj9Z3jOhuvynf7F9u91j2lpjPIzKOXuVYT7W
2MgvAEKHIF94+dFdi8PU23kpDIo+ep4o0T7yBCPSfRrqXl4ffzi1ofDAXXRszD0b
HJLiHvzOrLcY+T/WHbwRhUVwDkTsIsJiHZas9Wk4fhFUTX4yCFwD03SNjwnFwP6r
OLbtvxUTvfysvennJfWzHDMirmh+TYyouWH65HYsBl/CmWJxZBR4jgBFOUCw9IPw
cc40CQ8nrLYT6niwsU9adlGL+b5+L8cJmuMgcmt32I0A2qgvNsEg+LWvhCSHTH/8
Y4HcJmskA5RRZqw2VI/rbfNOG0H90+f2VW5hyMKTd+fOPtDFl27xDv1C3ydA3FkI
nvd012dssYCVrRjb4Z9KerfShaxyVsU7v5KBVSZF5VZYM2AFxuHcyCPfE6oOKJGm
/wiRCeHxu249uTIOuGRfGPpKr5yVPNNxvtDsyqnn2jbQWAiFaLUERYcwl485sV/F
L2U7FhANDBLVlFQ15vkyaWKGN7KMryPDUKckiCRzrYC4WyY0F+3VuzhM7bgexoPH
ovT5z4mSDGsVi2B2ndcDrQ88DqhD+ckB/a1bPXVaRgg2T3RfbgsnKbvoQFNPpQwB
pZRYzHv7XIv3sqJBoMHvXyy22z5l56k5tSI56JfO1qpHJPJm6MzdhknaK2sPmXe+
FQ+a77KvInqrtZ21Vg5FzIIAj+WVe1zJPapLzdw8PLn16Kx1rzRtXo+JeBkp0D0r
NGVz0je71XvVatj+IaJWctSaqyyIN3BqkzL53Fk8t9v5DYfDii3M6mX331suchP6
PpTrhqMau3Cd+WILfEmG6HC909RYdkdRdRsPpWJR0KSAaldTTFOZbiZihcRVrroR
dSMyhW1oALpu3b2f6BjYTWgpDcGeVXI7JtGlHhXAUdBzTwow/GnTmtgn2EJc8fMy
ugIddZ/78t2Kfp7eedcgWs4iMOyDa33Y0TqLbx6v4pefJG6In1XJYaBsz89RY7zC
FOA9klOyjDJyf0fk+ofWYwLSfRVH0aw5nN442C9i9sCgc+XbhKtwc2nt1c2aH3ee
M55gbKA3tJO1dqwtAQ6rfpC+TZzbd55GqINQufrXG1GQUrHUhiXxmG0rO1pZMlck
RzDTYXiudvbnLmnFxyLxz4bU1HkDwGJf8cgvWKKzfJHrS22X+cQVzkR6sxLIhRHv
f3dAy2YxNwOy6UGl2uPdZbbW25pOwVEEw4kyMR4qDJcorY1Q4k11fMsjzTfMIUu6
sr07OsCfYPnsOI0qSEXoxcvVX0wINn9DfGfeG/jljkll/1V8a3ndQDTmTv2BiwBm
6ZsEBCv4HaJw7LfeZKo5NGhbLvNl75M7mOou7IWt9ebY1EXVGAJzTh93dA1bEmcy
QsVtqbPcvSSYTe9pSJ99CmnZv+V6gybMZfSBLQSgTED+zpkK3uPdVC/AwV0rkuZL
PhsxSEc2GuNSnOeYbyC2nUu0xAtF4jIDs+ZijyclHvHj2vsgJWTjoM3zG03p6Pd3
5kxT1evcrg3KMtx5IW1ume2/qNCxxGVdOuDL1t3xy/LiAu9iwdG9XAXbaz6gX0Ai
kHd1kDU4Cc50/9pKrnyntri1JZaWPd635fN+CpVEJ/04zGfPNgIS7A1G2z8qvTr/
YoVEDI+Lgsm4JmqM9Nw8wJEL1QD6u75BS0hDvqFOk0GXVRVskbJWD8M2bIw5C0qz
ek+DSj5qprW1lgW/AuB6SCGGiisgJsXfvZXNbvZpJ+sMXcOMdr0gydtUsy4beVlF
ayplAuduixxQL1rdWNzvJAhNn/uT/oyiddVS9V7A9JI9FGNGgqZ3iNvVKU/AKL0X
g0KTPw481R+J24KBf4b+d+X+3vn3Qz+SmAvWI8e82Is5JE/l9JH02Mz5ilw7RoNu
/GGRc/3pWDb51pcQz6ix4QC8wl3gx+3l6W0RZ1R8bbLxHjYWLuMPgM9PMmN1X247
HUrm5/ei346GYvFyq1ci1FzlzRFGg/TP9ncR8XGZJf/A5VtK9vAt6GSf21ZcThhQ
//c0FGhCnW63dTbzTZ8LQYOL7+i0YhDTyvLQaX3+IO6LH1Wgev1LZAcL2gGIr/jV
lDafDmyCSPye/nZNWfY1+1Lt3MPsbDTKuvpjcz3KCQU8ZyhKk2ZkpzpzFoPBFRfw
r+O4D8DUbsYbGHBRfW2zHb5mXdOZkYAMqPspod3Wcgw0gcRXSC8Az5rqzx0zPIYo
M/KwBypTE5OhvN7vbXUGas0lwaax5QRgEuENtHoVtBb+6qV/F/mS0Ow/7J3/xyrF
sBaen3pnJ4jr71eMnqmgUb0ddbzGfjnDdauggwjOY9iwI1fx5vCJsHQ0qdJQvSzt
/p791Vbvdo9h2ncFBVLvoG9IAB0u3WPd9w+t15cfSGB3xVslvdwml0NHUQ2k4p4Q
mApUGtR7e+uXNsddo407TD+RS1Q4RTXDaKS1tlNaoRLisIVl92ozGevhPmyMz7Hu
ilaRN/yCv6lcDH21yuVGNC8fkNsXMHdKZtVgRMv2/BFadHA9Bp7A59nATX4G6PY1
Vo8blJGZNaYIxmTut9u0B7GLI/HBT6hRO6scFZ/TTC80mBJwkDEfoPErRPtLV5TL
5UWE9xpYhdlWUxApp8YnOElASIF8WJspNFcjw75eZ0QISULdE4Eb436bKTK1Cdr7
RnstR07Q3nIW77vw7aXAlt2poVppd0pw6ks3Cn2K/mbV/e7uA4Ou158Fb8ZvD3oJ
1N94KZFmIxNaqwihOAPsjI/l8HHAloAHS+gqBLPfLbHmArlpL9tOYlCP/hqs3OFO
lU/YKW2Kca2ao5MD0P4FqfUQPBL1v/0/xe5hZRymmgVJBaILBjFCziNXIkR7ZScv
zL7qGgSFPq3egsTwChtNVnKEGmtUowbHdNkqrB29tm1s3pddP24uPOqaOqN/ZrEV
4iL+DOvxBW8s8Oa141NCCM0E8s8sS9rnUkgSNMqjq6f/IO15uaM8dDnjsYXQKeXG
REBY93Ot2B3XUWmwI2M+h+XJOLHPw85SKMzPqsBagMM/SvWCvhUaY8qFpHeJah8d
VoeMhqr8zUCqvFQKRVJLq3gCbG/ZEPMIBRF/b+0//+nKbHFTWKb9NuCgXGBSyKO+
c6OcJqgwnR8vAa+P+VxiEQ80TkWZTdU3Yb2HTeBij/89xCfgZPHmf5N+vGqIRWOG
Y4Odo4HcoLLdtC/PPtKXsoPmwRL2akBfOuztOUQq3F3MvXFeSI/0NxlzMsH5EcHX
9dAWfNHttbFQ2VChdc9LU3BrVxQA0KnFo8dsyvLtsp9DUyNp/FjqEtrCsZIpi4z+
VjJOUVVkN9PygJfbW69BKaxTpwHvkritBjK+WwyvYG36uNYjUMk3pPZiAwnzxDU3
zohjicH7ZQqFCFFdX/RvylRlCjnYYTGXg04+fb/rUREtXce5xwpv3yazOilVpyF2
ZRKfSTo3hJ4FbhmovmQRcI5LtQ1gMZUzao5WJV0uZ8QKeZgXHEmyo7/mQeZ9q0Tu
iRPRMeqaz656JcKRTXl5xM6hYL1vCHjeBNwxzeGglnlGwz75UTZamv0cA2d4ZjC7
jfWfKMUL2z0DhW+nu7l3ysungvGkQ1QzWFPedmjvTtZFdEdI9FZsCEDrqeTI822D
Hg4HZ5DMY811ZibsQxCJGF5DKR5/C09wviAY4K9iIuc91h+R5muXw1yBlCAdIPOZ
m/mnWapK1N7Rf2vFGQinTP2R05dAivu3yip77wfv75ADb+d+bUMs9IbzYl0Z60Mn
nW3fl1ud5A0+sHNfy1Cw9whlT1Tu4nclpds7FWTCxWcPF7EHZl7Ii+tD8u0xxzMa
7pT6xKfcerYuuznRmAmDS1a1vcSaBUAic8Vo9MjHLWMfXjreNZJlDqcJ7ERR0Y8i
rQpe8bcUJGrnec/6yi48Csstb2i7h//FwdWtFcnQ6slmd5/YTWJZvTNVWLjf8b8U
GG1GGpvtKOyJebWFa5/rNho5n3+PCa92fTf9qznbZR79vF3htpjcLSZyCQ72vgjk
w1UE4yP4DOVv14ES0HB8koXq7HagPtQl2bLdToxk/XByXz8Xt8jNpV5t0h7K+sMs
aMeyVroq5PA5rq0so/rMMu08oI1JRVYRYsriPx4+/egsqa6ggCI0kFlnHSH6ZdD+
m5534A5lGQcJsXy1kIhJQ2g9YmdWV4vTU+/ntXIq4dBxgaeMaOPlXC8Ql7/948Pb
7GMEiWRhtkFyK61GreBiVeRZ443f6s4H8uvoBS8CEar3A7Wc+5iH+7BIoN6H+QpI
tTJCbudeA+woU2R26X6FcwIWLnLObOscbbfbnxNA35ga7obDiT77Fa01LowVzM+N
4EX6Zgl9lW8USx04nvoPsGevtfEgf/7IKkvwVbdgd1Ca957B+HXo8hpt/BAsCM7a
w7ue6biR6efNup+xfktFotVbVNi4zMlIK3DxXKJP4g5S1CNqIH8msq3Cm4bvwkKM
giItsANhRV90ysKU1usBpATIpWsgXNbJA0A9jBE05pDxCsYCrVKKVwFEnE2Q7o8c
3gNto8KCgQRiT4Uoj/K1q8L32UFpJjcwsOzkkh3ep+yk4QQGLcU3qw7gpiFGBx9J
qmLmgwZ0e8SuJBqIGGpsiu8GZM7wIGf9jtIeEEXVg0Z7LY2JM9DI7HK4bQj9YUtQ
bhlhKePX7+8w3NgVGhoYaFuQri696o9UhzLNlNd/6ZhHsiUkh9vhZ6TzClHJmp1d
BSY/VWmT50Fmjz9FYrCEL1eLgw5S1LO7RupxbUoSPEc5DO9HV0GXA4LpA14zQktL
kPK7Utqd6/IDwnlDT+Mz0sLSbf8W1a2gpPRJKpOe6n5p/jFtPlWHd7f2KZrKQsPW
ZGr3tN8eEdE3ocXzMpyPkBPtgWzbMxXtKw+ga01O29e3nt7YdemiBKugo+9fVWYX
ptXgoA+PbgnCSG4IWmFL9msQmEgjx4uNZMWRJSbMWBDedwHGa1ti5sgq5A6il2VX
KE2k07Z1dyTgVTEIsDNtgDvvWwZS32JqROi8Bmr0YvHGoVApU6gGQDf+Qdg6Tifm
mWwVlhkWc3Jd0UFWwxMliktk6ajAf5qbJ6f8ntCGFlOdJaVuM1NlVwu+wmEqSkHG
aJKlU8yYykams1iuTwibKdmodFzHaFyc/AuNT4iIGBIM1+B+lkJzp0GmrCBsN8Oz
mO/mwJKfU0IvF+aWw/72aFzYq8uwrFc/hXJbVLfY49gI/y6zbbsAcPhdgu8isb/c
Fe0mOwJztqCqFjDqalY+CoclB2bGBCv8KsKInU/kUU1Sddkk/F7Mlbd9tz2lz9ve
frc7g2DCGhupDjpFxsH/yI4Y8D+n/kZ3wvpnAUcLkxGSkLILSTp/fH1bzNVAP+3Z
keYiOknlUMnFPdwoNJKQRUCvN5ndvTmyMI34NILhYl/TAj4vz4tLg2wBBd57NGD6
ur9mYkdwRRJEsaxegvE1ZRYg6oR8J9CEOAtuAc046aYUTiYlfPwT28RUzmVPdrzr
faAzM/VPlcDIECwCG0O3mruphaA5F/DEODJ9uTx02nG/oXaonAL4Vg37ElD6byrF
9bYj7kIHBO6794cn5KEwSIGHGhvoa4d+c4lVw3QH2j4IvHKfx7LnWTIL6yxxFHWs
DPEgtR50+O7RowukjlHgR9QI0LOpf0IjXfFVHyxiabY1oN5ff2IFGQMI0LXW+Rsg
V65kmb0WVnNsQoUe9GPEcxCo1id0I9k5XIP6xqxD3yx/SYJ4Fn9U12eS790PpxPn
dXSgOsdAHu/kgMR85MPTFuO8w/RqCLvKvsmwFoIsOh2sfPZDPM5MC10dNn8gTGEN
2f2XzXKv+vW4sVlz418CO7AzPAYjJIfkwkRR8EUlCHgL0jUWM9DW/4Lqm82JNoX1
vyYOg5egShALsfov5Eb1gbil5zAjJOM3xicIv7NN3wl9FG14H3BDr6+2/XChYw9o
V5WsMjk8DejoWhd4xc8MUninC6LsaSWvfMkoM9djK5umApIiPsqtxHIS3QTbUWa/
kmcAscpHcZo83ujy/VYm6med5NkYxc1FxQup8RxPt2Kl02tVvi1eMgUMj3CFi3de
yWiUgpi6slSyQuwn+wwcm8o5iwrcbZCQp+aIJJE9PXHeDhUbRG4zmQUxPlap7UhW
L4qoQIqzsE0jdLYtNKUKtKojpTlABQyUegLzs5pov/oZ/F2OrCN1KRYFzWw1MN69
d5vimSXDolWlnzjV0FXow47uZGypfxrpk3zZchimZ+fo/ZRvhOldnhOO2gr2hKv2
V4+pjlBUp6brgY/dh1jU6Ij3RKDkDZRy56pLP2T0KR0SqtV58VvWFLkU05jV8rvW
990aF9bPl4EscGNcY99nilsyJyk4zfNBITL8TxKgJ4PhuXoE4QuXI+znYUTYN5qP
A73HZoEZh6D1Yu4ibY7D16esDdJiJ/3awAqNeB2KIisFKux2jHXHJy/ku2qXisLy
u/CEn0tvqM42u510UuuypJJ9xLaVeRW5fQxqhhhvyvYuvPZLl0nyAyovCHZ4aWYs
va0ThXkNgE8uf2bmfsHvJJhBaL3wzwvVGhogl+e/xchkvm4PtfCPFE1o791mOv6i
/dDpwubqfZ4zzrslRs/Sy4OXD6MOV3PPcvwhu7lXQi/ou3hEJbNi55HX9Ac+ZyG4
8IOK4v4vLkkp5pYg0l6bRX5B6T3HmJmyd2qyvBPyUJl1/iQGQEpY+Iqqvhe+3UFW
q0JxfLBwsuS0tJKWmIDjkctdlvkRtlitbhsw57q0MZmUJ4iw1Cdg72Zy+R0W4rNA
BePQLqq0rpmTzb8xOv4GAeKAo7jVbbgNWgGo99amp32LW5IIBuoDOVqMsZdN21kF
yZCGjxzewN4veGWOp8bKZDkBbHOGrBEQP9DRbjMFKf5hNEYIybF7j+3sNl+otOOO
LmMGv7E7AiD7OWuXI7lJDPzJ142dWdaYYGMARNOa+PVjdZ0kwKPi98sGvEsppk9X
76T5YSnTEW24ndEJw5dY5vq0++N112++XMZtlJZGx/9W93s7fZWVNA9P6IpgBpod
uMzuRsW+/C5G/wVYKzbCDPMLojaXWvGiSh1qGBxbcsPZDLtOjkVGskB0Fxe5RNKG
/dWLRwWKCwipwXkmnjWrtpE4hBDejbEjRFf5M7VwXoMjfo2HK3DBcG0VQTaMQZmY
L3IqwH8I4jBdVNVXiqsrvnmCCAc3qb2bQlHhE8i5/a5R+DMmqGFOv4j7r8EL94z6
Relf2fjoJMFteHAiimomkI3FM5hyGvDPjHYld3wVivMImwYCZRVFXLLRQ5E6wtGQ
+v96Jl3GuJRGJoZyJohNJdocxw123A/LUQEBjeqvdMhPOn8SsriANWtl30gRTuhZ
BDPejialrXiWATX+yCNoRaGfh9yxneAqtaSopMNUoTgdMOBglt6P8NNoxPfUT/bO
YgFGBn0VYcgeGdsxy3BHZzwNfUkc6TIInIhwc3IrX0cYIG4V/nue+hhtaqQlH7t3
XUWBTI+DAIOfBaehqHtmOjAONs8btyOpDozoq7LhytZBheHuL9KQ37u/qkKRauN4
NBkAr5ACYbmTJJlRhCZ09JlDO9Wcaqpy9GWYIWKR/oJ68idN4Ua1P573qHgQiw+R
Ky08JllUNQjUCAPkweQboJiZP3TAHXyV7ez86IlwICECastysZckgj44I9qJuxw2
oNy0OZndCArNo1B6FjEJ8AIzcZFqSOjMH8KipxWgvwAD4c3aoIjZpSBDEYZoqJW0
QIBZ2ANmu55XCkO+GelbMLHiQBx17dpiZvFUIz+WKDSnoln57UUOlWHq5RxvGBWf
taje2vcitM1PWUFZ1bQlBQfr48Br8lX2im2BOsqFCuy/o6+bo0u/lxvwEpy+MEzY
IvfSKGy3SSiwfnWtO7S11j6Mjsdz6sKUipC5/pR20GVBVq0KM8SX83y1jiywAkfl
CuqV7cwbuygEU171wk6tooh43iZ4dEwW/4sQtLqobo6yD8JztHW0Vz8ND/03cQ6t
2foDzU7hND/ODamVJleNrQdfgdXuKuTHaXNOgNr/v0SgWCjfevSju6lwmNgtQk6j
5BJdbmS8kenS25VO6S5szkYW+qCVjPPUqeJb83tyNJXN8Lll1NnQvBflZU+MLsQP
ynFTPbdkHtl8BHQXrKeWkNfqt7DfH2ThREUkZHfYgKjaLq1Xr7OvE2DRS9ZfM5vY
7oSpzNzcjzfak+y0SAGsSGoX5lYAVDgHHq2ZcsGOUqxNrNVa9IVlRrQ2G8Y64af6
TwTNP5ac0dboug31oDH7tUdBkwQiKapVWiLnubCHJqTFeBEpx2jVm6l+MlkbIVKW
F5DLtrkQ5PIiVawoIZ6d9o8Afkb05+mT0EDBGiRP6eXPc7EsTcLdNDLNOE1zEWPN
WAKzOI3pCKiHO1VHU33+QOEEOvDJmogq9kw3pF+UCsLHnqcplsfZBMRvi/TcRK5q
kEGljZezxffx6HvqT/ohMleUH5/3b0qC4h2khOW4tHiv6SNJxnIcJ3WzSyI7YVJ1
O8KKfjzun60k4QPhESFXahmXaEj7Ds5uAAVGayGRHMbMdMZq2SAnOaoG6AJ36xLW
IlkMwNGWbRXdySUpMzH0O+/fWF/D3vemZY7Y3bY6ZO97wXAZwLLVVIJBdmVNtKFU
SjQyOCg6bw7+Zt0kljnFcrkCTkgTr84kUOrHHrdnTbn/EniHNjD9lIP5imMXxeHD
HoiqrSp3sWxbl6Sj2g4rbzMjR+6e2lyrubt3xXf81IXPK+nekqd8sNznNrExMTst
PXVD540ndHirTj6aJ0qKwyv12ablvQVIh388Jw8JSHFbAB/VTlO/JjiaB6Y4xQf0
e5ux3NZZ1MDOuJnKOfzwI9Yfd0k8AKUKp4ed55NXpMZzjtAWA8FB+CyLmgqDXJs7
d0g08Sft6vwD5LMrIYE5Kjk3CLMDxPZKSMerz5XjTEMDLPxmMUhm5L1s+uDwQLy5
9a3fIR0t1Lr5KYmu/9ZxQ5pPzstgRvm9BzOnEfKxBT4Bttqm52C0+TIJVvjGSmbk
+fX+xql+7p6+sKVt9IjEt3Dok/YaCLHLXHCjXDF3+s6CSrh+e1HPLuZVFHglLLvW
B+oB/86Mu7j5TgOJdpsYeInb768K3FwfZWKtHq5Tk50t355xXg/jxXx1fgRKXpIU
DM8UI9H5qP41CQxrgtiqjVeq+9qY8r1YNFmd1uRJPeuUmm/i0ZoRB191aL9PTmOt
OAXl0WI9ZLsgifgx7Ik5uTtg3YQqacUCvZX22Qx++gd1raFB0TJjpCd+/uC+i5KJ
nX9tu2jQT6w0zUg9ywole8BKhoLTmvNxTwl3Ckt7xCqBjxAZfGbh2jxMTZ65c2Eb
w6ieqktifgifCRcEbIhgHP4uX5kzDsER9XautaHIZiChgvZDHgcOnPYwcxgLCqPE
PCdFbicWvwJKdUkQxh56vdsIc+wPgfl3ABGErKDdmu63HgPNvb9l/ByfNZ6LEixa
D86qj0Uw/WCnY/xjji6k9hrXjsov0KunQYv/PxcbbWbYqyxUE9RTyllY/zNL1Epb
d2xKsObbfxJfN5h+JTqGcuBq1KtyaCSzJngloSuZ9L0/4xiHjPDj76kJQiuiFw3V
N4tYi2NNjz0uyjIKOaAo0+b6brky+WELtk4qpjGeL2h4PRv11BVXIZ7+85fILBeL
EMG1czYuDgDzq8DTFzN63rrBHWrRseJMvYt14xj7DtkHFGCwHBxsIE+g7wAOibzR
5fGUqQ4PvHI0xUSubitFZnEHUcW/zDD1k0mXPlS22rphgH2NkhiwTekQbkaK+vYw
WOp5knBR9d6lX0xoDr1E41dJ6hv7HPRIxr0x1bP1bO8o3ZpYmiplfXok/zmNttQt
ILZW/5w8Mwq5vf+7Ge7Xwqi/sRre+rsqdD+ghc80VwnygPxX9w4+Rq0+hsL6Xw3s
e1H8EpIMMss9+FG//dkbEn33ijK22e4oI8duRNu53xJV1MltIKqfN/v5L7+/Y54d
eOnqPSXKLyV1oUdx5DzWgsrTk7X5hQmJHjO5J17DkvID/X+tM/gKnx6LBAlb+N5I
4p2hz+LKnbBH0S/EG9V9WHqLHGS/vW4ytik81k7RXpeYxvc5K/ELAOoTqwjcYVc3
+JD5L/wNDtDGK92ECLncR8ERT7FxiHJHIggXvFM99KbEhbboXwaH6l192Z7dNi8O
gKp6COP4RpqxorWt3A/w9SN8/2ZUVzCEMDSUfzvQUm99YS4kfUQtUxrcRwKoi+sG
hain0wK7zyeo74X48mMKTmIjDYFuwhuIiPazMJtTpjMx7PrwTQBCrJDOnFhF9uAo
vPdFH7Xdza+8aHx3eENBfgXHHj2Rjhox2ZFZOZzf8xc//158yrf1ZJnVn1DgrNs9
x0lpzL6mK438+HyTfXMT05s7qaeUuLHhtJXPrjxT0ktId9RUgh/k4SF4Mk7L5NYA
Q67zn1S9sVIhxMC6psA1fU3baa6j7q9nbSngbJbmB74QvVTmlfsMokR+0a/5fLo6
4w45IGKErjeEAiURfzXKNJRmkhs0Ntqti0EoBkyrF1R0mip1KMjruHKT8SFof885
Udl5y/IBU3k3i7lKxdAqR2VmtfF/hWhXDNeMZXLVdIKFQB6zqk9DvfV+to7kp3/8
NMF5qq49LM06C1pdkqf7OtD7CuKKwGC8I/QzfrybyxyZeDtRheWwdiTD6iMzZM/C
9RVzliRnhJfAWnHYYn1wIlX4IXQ6zKi0UL+gdf2TlvGErVXWQCbiTVU1sHzbuj61
dQYtKJnIJFhRaOco5e2LNF3sCnJRcc/Gn2pGPg9O8Z9/32x8OYFaUqA7HRBYI1eI
RHnK9FIoBdqWD4W6KviBCfLPlbA2mXAwM6qZm/L6L+jiQedNwkB4s8b2/unsngQ9
dX56X3wnmk+Wjgw9uJjkM9gF8tpbs7J7FUnBpJQ+R3cJKuQJ/5b1dHdJeBhz1n7+
vexpMm7ytNkLjQGExgOtzoQR//HAqcSb5kXdrwXYm6d0lMpcEL4rsj5RfN8QZQ6E
ivaxMgn2vkahtFbsbTp+5bgeA3jcnOTyU/rAE+tnYHTvEA4xZ6+Z4I0XE/XyhhRn
mCSVCm+Vk+ooJOFrNeaEqBmIj8ZOpbU+9bjAjn5sOdz4o7hZ3iDFY+V9ZsmLAuCn
FZUG3KcTx4pVDAysM9jLZke6oF8RpoSdF0MmanTrZTSHg9ErJ5pm7GGffvPeaabW
8p+8L7WrgnA/7ry+ZBXj6R1mrI7ZJYRcACcXQEwMzDVLeAAkWkhjeXsGtw1cXjJ8
AcT7lPMk+1PImw5EPWMpt+vHbMoNNG0ZmF1H982GHc9IifCrOhpPF2v3yVJK723P
7zG/vsZHBCCPnpd9uxQabweGAsL74z6gPoZd0wjRKJ0EYGl+O9vluWGMtlcYyqT4
EEyyp+j8v/BuBMTOOCZEKz+ZYeEyQWbw2VDbRDneWDd7lrndB5t18ix5Uf7ntBkR
baNPZ2APghp4MMZrZaoGLDKn4xscl3oyo0FA6BI0NSKPPRgoFA+TQuCwNa9h769X
UdOTiS8aiTtWOKh9cf6dYeANhw9TfgKt8pe7wMOiSCT6XT1ndAzuYDHCULFPMFFJ
mwvZbY9VpJKibp0ThyD0fvtIFkuLVbWuf74aoGIX4COqmdPavdYNUHdzGw6bAa6J
qgZ+nbhwkedPI66hNxsErabYJGUbH6nsu1lCZH0Dz8HZ2oAJneeU80TV8nlaALHT
skfRdn2yH+AyGNhx9j1SwIiJCBNdvNKQnPQy+6I8DDldQ7GEmEIXhOzLWc5oj2co
lHvtO8eC72IAwmbdq1XGnv74cJeHpwnVuMZ2tEW5ttlRiPqDuUFOAkRbSO7WefLB
VBeUgwkQEdF3h1na5j88Fccvbh53874sgsl1ieiRYRG/RrA318IvsrhcyBxKaI+B
jLGws3rcL+mpGt5LZ6EuSPdLy6YIWBRVllYkJxH/6q9Lu0+ud2wi+8FzDbyW3E1q
Kb9ywUI14ClPo2GyZCCQjvRcjqPw3RsR3Io5TFxhOgIbWk0JD0D0TG44fiURr3vh
syPRikxohidn2cejs57MTURQaCOgRf0AqFtxnKURFKOG8cbq7WyQqWoVOr2HwLV3
j3tJqK7KGXLcM65NQhrtQp9DaM6MxrHUfN1ZXxRa8KV5415VCy4G6AuSdhcypVIl
3nNp4UGgOU5GKpM00m8SUVHgdv10SLBRGC/AH0iOFFCyPbbIUu/s3THSspf7BnRP
jRrr6DPkUA8rYBFcjQKai08N4bTBGyABtW+Iet/DtIdD8PHFAUfr6+sM2yrAA5Fh
0ibYxFpU+bsz7/7jJ8ZErlOV6Edld7aVN7wKuZnx/4++0hm61rT8uvhpe13cIg1U
voGfIxp6wTW3e5yPGMWZqDJGQ1O9KxFboz4Yp73MqLzbGVahuZY16lMHpCmj+xxg
eOjytx4Rf0uZQzJePjVYa2RDjtWbLsU35KNUhW6bYOmR4lSnb+C/tpwDjtq6QFYW
2DigtvseL9mn8g2d50Jfoyvh3hFfDZbjU/TE/55xLhKBG2o4fzxON98c63v/pWJk
cSrBxcmbjhQVyW3x2N3EGCBN+DmrJF+PSXYh0OVFfdbV5fGOy/a182AAHEMwfhw4
pH9bUDrSOr2p5CVjRRQKgc/uX7hXR8zRPQ/4mYjSgxnuwgzIqHmE3Xqybk97Xcau
0fKNjjqSZBrpyJ/emQJmqXRClg4tyr3dcCa1/c3rFewJ5oHNKGl3U7IjOSogO6OL
ULt7paCj/2siO3AXBeRbK9bpnSNhNJuOLmqrtwftQw0a7DxPYL2LzjXePbq8JrUL
it4jhuZO0EuXRSvwFB2u8RMnnIPB8+vms/70stxA8zUey9fswbfzzy4nk6cB5963
4pVdkJHviKZWQ3lkrDi/VX4zGeCeyEHuIFjci+OgHHiGeoBrJfG7D4V5kAh25brf
dHWzSPLsXuHQ8HvJyn3pzo2ervMf9Tyg9IYRU6RmHWETJ0Ug62qfT20AQ3wPzq/E
kKY2AL4j7yv/iirqBBQ6pfOSSJtlZnJroAFocnEsmmYJ+azh8NaCy8sn/H1jKdKp
r75BH1UaTS72PDCarNGLo60onFm6AfY/RUmNZDIU3+gXvNOB5gh40Ph8ZqjVGy0k
SZ+2n5ZyIQePK/L3Y0OHVQlQvnEUGSCdXJzg0gYXSEalRGU7CUgTlzT1+JaTw2uH
V9vTDroUu5rSWRIxT727JjfcM8Wzm2Yc5Ln4eCB/gu5J4ETh54D0tDV18B50u0aC
JozsC1alzVq+L9HaeRulQOvnA97pf/pF8oYXsI41HdU3BvLNBuPlh3t/w0FE9MP5
S/DWgwWXE//F+FhMtGQgN7hzCIs7VIhhfZeFfEf5BAijLMFXd8jGRos4wJGniU96
v/1EzM4JTI+eoW4SNdjdVF9q32AkV2vo6FPf0O1mz1x/Rk1+fzdx2d3NGls8N5/b
N9PZXWszqgV1caswqk6YRyqdN4Q30oZ9wBc3S6CjRmq+GSiAuQKuEWLG3eXFj6TZ
X8PUVhM8vEt0qR6k+sldeyTafWGS2Jbc83I3wMGMLz6y8Zy3kvDPV9uxjcjDKjiJ
DV13hLhi3ojXxW3TIDxide16PeJ1OGPGcwo9gyrZ1You5j2vN3eOHN8GNDOkLBob
PcVMSydVt4y5R5sdLKCUo3M+Wzc7kS++gOieRokgHIqoJKOkjvuZBiOWvtfChBXB
qturpphZn5usztqFIvsIs17wHezzivJf/dUwhRfsF+F5JoIYjSEu7Ma6LQfHMKUP
PS0RdF7AHlZZ+/I6KB1Nic6v/Z7iBl5JMECDFVN19s+7aHbN0Q6h3Q1YaCn8dPST
a6tVA3auvFXf6+kYktGN5slAqRBbSkxY0v/Cp5HcXA8UzRnVnOM75yMjkhPglfWo
SqIXEM1vVcR40+VJIJfQ2jbkC0PIKd3m5cBauK8/3leZZq8nPjUzTQ6cKzL5G5zn
6Xgpvxnd4iMd8XLgyUS6+3NzKCYdAH0USmv5PvknvxFym20r/p/+r2dxK3hD5j0S
FPWdAyFHdlxQExV7udD2TceIdb5Rqo6qVu9hv2Mz+I1tF3jFqD+LlfZcRLCo2Tp+
LwTuAgp9n/H7S6L/J5c3bNyfyhNzyfcB1KhkkRxshTJvH8oWDvDDZqw9QUuDpzYw
GJViHnDhZSIo8inZNY/WipbwB3VVDiNojzn0IbObSVIDR5QeH3OPnQrA7QBe/+yO
1l9bbbsn52in+0jNkyIsjlKNng7ZtU5HS6WYrYoRenMBkMTvnOdtZ/mK8CyCiAQo
oJT450I/7GyClEghmeMFq2xa7QWxqkaXMRdzqN5VaKC1SewUoWGM5IMJw6drwPid
0xotKH0KyZnzKxmUpxgQAZYpAkuCqkEUu1yV0lRLIOdwNvuWOcX9OoUL5ujle+be
Vd1Fh1dRUBHr6uBZYI9WKLrXf20LfQk0yq1tnpTepEOM3WCyeLsdE2fmVdA78i8b
Mi3Rk5QI23ZPCpEtql4yHiJX0rULZ2OaxVxemWTYTvDn1KEvMTe9LsB73Nvts7fj
kPOLm0DxlA4XhWE3JTa8Msopf7ztr7/375FJQbd1gIIrRwoT6dKeTFL1IX/HQf0j
a4BnKYBYLEcVCJyCdONLhpPLWuU7J9BLjAOWqCUXes7ldyMJIPtYwILH2k5r7HWa
ubxjfY+u2lI3AT0GB02Hch3wPhO4g9rDu5Wz8W80q1QuY31Wo34D7vD/pdPuYIzI
BckryvWBkQHCPxRoMi77cfDOxV8OaJULD1KJ0YL/uvkkRMOV4QY6sntvfz1jPCAD
eD4essUD365MH0SdDFwT6iScDqmfRW64vbsqdBZ4fCdyOxjHSQNoUkO2v78Daac2
/MQ9GtCNfYbM/ms0cD4eU9WcfqpGC6zSsDbAJYdmxQjh1sOnITI2l6qtsQlDaMEs
QtajHt5bh0p0vYzDsSfwIOM0OGGCqt14xsycfOJOk9T7FI23OE1VK/t1y1n57pZF
mr4aXjy2geY6n+JkZJVmS1zXjzqTsPeod36RV84AXZ+uRolNCR3W13ESI4ZCih+n
2l11O+TooLguxVFRYLKh0KBxDfb6q42n7+nx5O5HQ1rCYuE4VXmoSkAI8nb5kq7V
6y+xKmNVtZhrFiEvV7rxIhSq094oLaLsaBE+DHb1A6hZCTJpW4kkYexEX4GjRrmN
EVUWGkFeMnfkLYgF2iEkqH72TktEws9A49xwH5spxQkbavpImBiknmsqeZ7fKK7w
AxQQmt6SM5/iWISbbiliXlMU3seMOzxN9MKD71aUg7tqDEpR67yihD+iNyAoIeQn
nnIjlY8rDfLNgmTxlNm8iDfs0AEGpjr+PDbQsGPtGVujjrztCwZpNe0nf89T9/jg
4xfh5W6lTwWrvX6jXQgtT9yUQ61nBJ2WsVtm4e5rGYbN4vX+6bjBpUEnh4/E7Skp
udq3cT2gMCaBasao23HOHH+dV/efzVbgodUrNkiJJTbuNCwNrJ91LOY5FOALMn9u
QySTS93UeIa8i5vFxZQtj1QDglnrBGxG4MYF9oMMgZlRrsJlRRQKlrnr6TA6K1gH
LrqGhL5FjA70cIbqNoIWwwbjQz+q+tBklB5wUnhCxJyw1efz8Qx4EwVI5Juag/1Y
N5cbS7UwVQzX2OD66ZIICLmKgWeg/Pj75WdH9L4NyCAB5lKE1aYOQ9mUA3jELox9
2yalpSmtZ7u+l/V7GxbOrRHWDD2ukMD70xFJS4vYuI84649T0OJKsnrVUCWAxTS/
SyHbmTaTi3OrEzTOl6OYXIM4ftKIaRCX7eISdBiAJww1ZWWccqVtQq5tFSyvtRrq
64dDqxJrSd5evJkiVpe2LoboDJrW/d1LamghlnyQNZBkTzoEM/fdZwzy8VvcT4lL
7lMjnY/Q3pjzwLCmy+Hsfaj5neC7cTsdnWOzR+OuFtnBE/UdOWONqc2z5U0X6VBS
hDzvAtKZPHStODqfTKVWdorYlZoBQPE2RpRFuq0tGRvLc8WvDwAj72ETkes6uA2y
xrpLR+NckcSPszv0XDfQBCBE3rA1+uV9JGxLCEQNkUx5wGEwYfMTQbn1AnRjgbSg
2gAGyv7Iu0xR25i7wEK3SQWfK+hIF0gEeQpcwF2uNbDciofp0FfGNrb/aieV3ttH
RL0uXj1V9O9gKLKdGR6lzb39zrZFBXf4lp1d1e8gQlRGTJF9KZKfKHf2VV+QrpPP
7aPSQWCPaV+cAe2n+D+VXhPwIIgEJbVtnkeCZp+TCeuVlui7GsR0cJYg6mZ1mPzj
5TDsruSpHQe5gKUcneqIoq/9Os83DEiOhUTksL7WCCA+/UwZBK9yK9RVe0nDtRFK
7feuHL+s6k1fJ/EGN8OiAOBbBNKqK6xNL7AKuB5LWz+LEURGXc/SfqfzaggCiHw8
6pnjrsWJc1/9QyVh73iVqObb/JDtey/DRU7oOyx1Uxt+EBmTl+TchUXezdbXm32K
nkFxc3A9iVjDRCct+jj8A2jfXswaOCXXRubCwe1k8FlOUsmtwPj+TLp4tX0hXcjT
jGG0WaK0EEJO1HldAwYVQAUZtHFxsQXzsVasH+z7ZYbXSOk/MPCXZQVVFCql0dl+
mGkORCdCBnQhH03wmaUhUCNQK1T7P2MxPNT7C4o/1PsiXfXgn5+SUl3i9wAlWzNa
Ecr4c7pAClaRSO7YnklBmSnnJYHwaYJQSIQHkGIP3Zcdak5NWgCLqt7n59Gja8Hi
seRN8zZAc3lpBRuQIbNpY24soRE/IZ4mK1TOh9muBuYUw3BzxHvS/Cy8zry8Tmu4
CqWe++ekYRsmHeLwtYSIuVkwrqCDU28g6iOGdlfi20fwmcmRD8r4AKDKRieDYEzj
R1zzS0vyQIOnIN/o5tLn5E0oDH7QiyHa+sMm/rrGE5BhixnHWZ/auyrEIt7BSiXG
dzX5kMQ/cTJ3nNUuCXQy1U6P47D0OW5W+tuQQq8Fj96Bd8k3DhItKkUmizMqg7l3
9VlP/kBZ2njMR02Tjwp4sQeDuxO/5VeSLh1PLfxsF8xRK13E2DZs1EwhdK1jYFhV
yLxnPGyr3iKObFg6W/3RpMOCl9/GvRPbiuTlLvzHFjxShdLxcHcbOxdBVO1rXlDs
P89WxSC5c2XECCv+rhaNlxLWk+vDO0eNv6ohvn8IvlHODZiGODiWRtygnI3/A85p
Zo4PXWH8x9w6WUREM0B/d9K9SO7lwJ+nBT+8qRvvL6e/DqzZXJAyyf0QNyfimMWY
eSkh9jfYB5xd9pe0RixUDE8BHyJuqmpR1zAIVradRRI4fxdGQfN80iGFcnj9aIas
qjVNf8EwyPbkabey3njKqiwO4a3uB3VJhnfcIbZn2B50tMtaOyWq+LLUr89nnY3T
F0h1n6/LcHnRjx+o4LfD1oOkA02rOOBhcWmZc1KdiAsndkkG+5XWECmb01qVoOVz
6j+yCEPlG2UvyL50CfsJwh3SUK7Vds4h/8pI/5MgHWtuyCtqxwhogaO/TBpMDeSV
7FFscQximsWxjAFEF3wJ03SiqFAe/aBk+57YF7K3UXf0siUgmsF/j/SIJsFK4Dgb
Oh4/gO6Nt7srOT7e1W3XsRfPm9Z+BjX+rkJBPBkhKUM6K631JQvqSJyD53ZwMmfZ
gw5mk0tBYWycnIEVVsospIQrHjWCT4ck+xDnrt+2n3GMNhbG8Fi1WqFDeX9d3GFc
RaUeKuIJYmq/AYsEa80LlRhN/qy1Thok6nDs5EZ4hNzaEsOrq1lAziT5wIeh0WUR
gny+64MCMoFKYfUzPoB4BTv39pUMQui0S/PHqzApN5GYhV6kzrPVBnSYKHSBK38H
nGdCZA7+6fdbKjlar1DqLPI0zWOMhUx+D9Jr3a/z8X3yElWmY8+QzCFKSXLu0o5V
oU5z0AhLzhXQ+nJ0cFkVGMXwdq8yApHDtm1ztYS3HKS7HRaQNetBJtKUTQVhPCBN
xgtbz0xhsa6uHMPPy/sfc0sqI0SP5D3F5c6UKtomYRlhXbq3Wxdjvk64c2fBBJs1
hKJ77DHMGPVFMtH4rUQWuM3NHbmqXcih6c02mVEFiImgfgyKK3Frpy9LtHYWOnWi
D35ckRR8Hax104N59xrrKFbeXnuvyo30i3RY08Y53NHLXvWY8FCTcTav9yMxF85W
u09RZHkMQ9OoaxhQOYdiF3CRfcFKCDZClsLNnHlDn/7FMkrkIYjt38O+nrntR5aA
0mqGLTa5alUxCXnIWqUaf3FGWgK+C0Yb6CD6ffY9R2zDqIUaafo6i718Kjnxs2FC
w505TN6EZKNVgdd7IAq6fag0GmQ4MrREYOuJ/isrN31Lw+wCM1gxztIT/8ovvpbb
bsH/dYTVGByFdSxaj2bAjt2QumKY4etTKT/FNqTFjG7JYVbs+zYN5/d1FJ1TbWIh
lcUzHgoP3SNHgGHWFksL5XHeNVAAFW+SZvAXSd6x4gCJvgdeFIQPmMZqbVuK35+b
fqZvfVkZ91SskmsW1Ot+gfSek+ExctJSTQNPityDYQOkY7YztFSkobOiuDMbvydz
5ZeCVMSbQOSwSJBb7QK1MgASv2c9R6rXv7fD8WtRxhxKYSO9sf6XKD8P/1leDIJs
BHF8PMu6YdKME47SOOP4WXOTw8lGMP75qSyrPTLo3d5aXp8G5P28QSUao7ZdwBpp
acf4kEZ/llEeImC/NbkTxqxOmNVvz26sK4M8+mVnsrM+B5i3Zh0D7Dy1V2Pfkl4A
N/BcmrZE6uFFCe1Xn99TE2SBMqY/8tpWH75KRwAJw5mXcU2WDARn2S80nHiC+TIE
JE+XCfKGwpyRjdfFNlgh+XRJcPGnLyC7G8iAjhvx7KFi2xb79FQAjJq3U1z7tWZM
AaubFPfu/kqn9KpZOtCITTuaypfdKx+6hk4zZMHKsAfQIFhMfkBfF5VlG1MtjjAW
PVu5VW5q/rlYHRR6ZmPtjRRZOPg8OpSHdkltEfEmYuB4DZ9Lr8mpsOOzIznu3vSM
L21iUGbELRv0gJI893AFg3R0S6hX9sjLqQqrvv8K7DaUQeCgc1UcNLTy1EMtNnsK
z/QQaj+N8YwIcUzvOSHkreQVRR9aMB8Y3nf0utEycW4wOv2SgqJF2JZOVLwRyABw
14U1NZ1fZjphA4oKrc+xAdhYn0cltKpzmk1E9Lbr/m3Fv2cFZBmq+xBS0/PUbEn6
ZrjEZ4xufc9w0U3T196FnV/AeAAc3NKZpDSDILh0DdxS2gbXQ6z6xmDzGJ5ORaJq
Plcr9aLMHJBofD2zbyqFhyu8bZ/Tyo8dGkNMXpQrXdZ3LDTuPu7qKDEHzV1L+I9m
auby7zPRKRuaMALHlGKU7Tii26mrWCwo2S9ZA8M2pvz5eutjHN62XnopPuhelwQ4
OUavvIwZUPnlWZp9muWTEwHxsTXm3JjeTIk2lbMb0TRX8t7IIuoEFykn/7mnchnb
E8YvRQBv4oR/o/LSiupWfzBwgJWSUVmqw96ouqU4jLef59bUnFs4c6R/MmPhQjWK
o1PmRxX1w03XwTfRF0b8JTNkULOKGZ3woYAA73EX7vVAhoEsQXBniRm8FdTSIvrs
X5PuSOQhb4uOcBbTrU3hZFlCYnqRRtMmKp2EnVGA7WZ8mW4pHZhj3C8tiUhJ9A/+
6FTI6sZRYodeqjtuXDeQb4LH+JtNlUDiwVecuzsONY0+vrKEdK+IMF7CAV0CogFB
ivSIhhzYxlOLvSVXevYIG6db0Q4aACQH22LF+DyZn+TKK8dxXoJhASXpKBjWRNLR
qap+SXi+ck2jF7uRx21UdbSsu8VbvshIh5JMz5t6le7pAQc3MxBYGSVxh2eZLU4o
GgpLhEK0JBzuGggqjz2fbL+pGG0/h948CsCLr3JCZW6DcDwfmTOEVhzXjt5b0gBB
yMB1OKoplIKmsjQYT4qPYV8W+gWz1kEByTKwG1AckhtA7+KUE3dd04Tlx0qfU+GX
Xr9FxtBNaSA8d5t6llYryDoOmckSkBzSGplHjVQo8VTDHaI12atZQJqe2V9/jCi5
r/c07v0dcXFSY8NHUgjX1eYisML5AfAdo6IGS+dHYvqXZNNueyPJZ+WQ8+K8T7vH
6Cy05x68bSZ0SdSFhKWbF66d1XC+jtR7pFH5orBuL7tRNMJjcjXN2cGTX6iTxQNk
tfhzaNFr9liVCSNJ0nBjfemKj3iBlJerShmK0S/R8D3JQKLubsr+UXy8NnL6wWA2
o9G8mBan2uDDhTvDoVTDtYbXUFK5l0WlQ2/1pU1mMH7xCVeXWH9WcRxwKbWifkqE
Se4eC2OxycF02WmLgEpRClkdwskP0TaMq/CFANOyvLoVU9emk2dr86iSPp2FwDgM
UESSz3lsoa9cHFvzeij4nqbVCiiUn6c+C2vh/IH/tuQR5dHzn7XM+Lu0tDvc1Xv9
G3RcFZXjlcX+eeQHYBMDbB7Ei79ZbI071z9khZZRmRZNxDCjo85JPr2KJF5DTGCC
0oidnhVXXbS802UXakb0tUg2EQNssPCFw5Jg2mKswvWuv6CUj5NddIIsOr1kmhdb
5ajGk/laftpAM+71KaH9eYYkaA6dRRWjm/u5lExMx6rHTkt7+OhUvYjGSqdNCHAF
2iGnb8RRLwjQ/SaWl8+8rGjJ+iw/StHpl9F8TxUS0PNza4yg99wiEJVTiHL/bUBf
6764FD/LMCGnOiHyhzW78cx+Yf8ADFEXlaxA0DBWFc2lmn0HBaPSCPv5z+h7nMad
XfeXPXKvZamjO5gMlul2sihdngXjoYYLUwQNqgauaAtnMUk04WddNytwRHdjiVr0
TA6WaS61g644aL6Lg+nHWZoZzZ8DXxkiqdXoD31XkTgtJLPNw2/T3to90tiuq9PI
meJGW0Qt+1bk6MC1PwQ9XAzJ+lDNOr8bVub+xuw2mikkuWJPFV1QHnuv4caRyLfS
U0be/D7NVuDuImxuiZ2arWP9K0+jNyzfGe4rMTTQQsPDyHXfx23kAFRgr0Q/Aomw
GsjIWx1lHp4+1HWSfLiXWP3G46W7W7aBDw3HeKFdjXlbu9QbsObMGfJ2J0Lk+nHw
BPhgXNmRKa8Y6B403oO9Q8pKYvCOno7mCOHXIbvSj2i7sBTVki/wnCszRaN3xYhc
Z8b1uFEigpFKneiLHFpzzySsuRu7vdkrpKespssm2KIOyyvUY3oxW0p2djvAUoYm
DzQr1Wyel0pJNSGCY+STyaO7WWFYxsynwzt+Gct8Vnzsim/rDqpYAZQ0Bsi+X6tJ
5BQ+GaWnA0C85X0Ir/ExmLVk+SD/6dlDYSDXxoy8vOc+Nda6DHI7iokUMjkC9LEq
Od3M7risqI4yoJrSwes/1mG2oXi5ReWZDjpKalqZRawamHClJbEf6nlUOBI3IAgb
cjmyMTtO1/5XHTm/bQE6Ofd4V+vC+DYhYNLdyBOBHA/RAOzc7M32ZUFdczk6Umvk
n2rZZ1M1MSA+30Q/X7dMzQNYlUonckqN+C2rRcNPdJiU+8yKiaHJZqEE1p7poGS0
qk/8mdTuzNErqwodFnVgF/zYxa4v4bYj6uuWI/MGmX/RRwLUnQ8JFfuGJ0HPk+rC
acXc38543ZUz2r4upXSd0h02BBpzkbAqyunQJQtcg6EyjeevW5iyj1++6hIO8IKf
BuaQYmSCwR3aA4L7gS98Cr0KPpRirrQV+Ivh2tnMeaSD1ufgVJvP/oiunkWmxZ2O
AXQBn7C9HxxYnN4aIGhUtV/N59p6e/q6WY8iVQxT4J8kLn+3nzek3pH9hsVwUlJQ
PMexO0tZYmczE2psbSPOmpCTDrbQdNGxc/K5VMyOnzjGRvgYJ/YAGMywQpc2M5wJ
lF7sRSKILqi+H4KrWIXCPLAKZRfgfwApmDCE84mwSb0OYrUxnmDwRJfEjIuHpDrO
Qk25GdwCupJ15Nab5pZhU88EIRRuWNHLXkU5uM9mHO6+a4fdK/GnGI/ixcLQZKlU
MytJmukiqMnInN8JAYGYQHdDkYwzXuy4PvDec5yRfzvVP2z72GAs6N+C9CCzznxl
Mj6wcGgoYHVlrb/6Co5M8ho/NKJU6SBm4dz980zQxzyEHVKCcmFqMXdSVj7oftNI
doubmA7YD0w1g77145T2TzVAalo+eqcDEmo8IIfNBTunoNWqEoQJXw0WRRcVP3UJ
gh0EmZdm9tEP9nkFtuBCIgQlQBMoR9jQkBshdwgzVRyUJcn2IcJ/AkH06WabKfRP
VWg4uIPAT9HPZf0y15h3rfAlvFmJQcJ6s0U/DJCXp8tTsFTDsw59gtsaC3rCyYq9
R7TqJaqfH2OOe3QbJD3WRrZ99eoxbx8eaA7KubBdjL5ysBCtxF3Mgw3r1GHUoP0q
RaJzw+C/1HPyR37jef6/phXSOl97IsVn7p99lYoMMj93clPVeJE0H9gySXUTkobv
SC78HEEjpP17br5XWvnHnj4Tp9wLfOWnSsazpjyXWnvYpVtaoT2UGWrvufGF8vh1
jzxFrTDsAZIp+xODmKEiXUiqoWibZUgaI1hJA92r0UTI96YH8xCZvIK0xP7qcJKc
QS+QSnOIWt8cy9972u9gf4jtpX+IFjVlckjVdEg6xoczR3ROFisTvZn0uJ9LOsOR
bmyHrTRa/DStrpJO74DL+NMV+ImFOeXJLrPYGS8V/WOGTqpRXGppwOCnuBpiPM2A
2HayHByIvd6IXWR1wXRT+sl4csqosQEitqVEG4qpJ6dRRExRKG0UdKWn08k/Te3Z
Qr9lgeAsYKceKN/ARED/RWiqQmao5cswYRUx3Um7pExg1088S2OJSXUMIF+PDoRt
NPqxGxalr+QZM1pluMqG9GUzOYpM4rTOFpV3fSa1s23kKs2SHSzm1TldPuo1jZVQ
bipxn1SzFj+3ou6Wb2bTaIGyrWN1DfOUBrTN1+DOZY2rk2Ocnw2WeInafpIho30E
kz3Nsgzc9kfM6fO6tM+1ViATtaMel/QPythXdx1e5W4vhNmWsOzDpZVLWVdvmL1L
LufzVZPwtB+8o7UHYidg0BFW6HDhWmcl5+yEZkbwTSaGfvl/GZp+x5OgAlwNX9AB
Xz1oGWD9lLRrqPxeQcMFEkxR7GF4Fsc+zfyjA/TYrNMD6EzRfVxK8o/N9RIbf1Jq
+I087QbqN+UoZs8UJgM3JuCwI57KhxaexYWKZWCU4lQKD5Of7qpPr1CXf/NkhuFL
X6torZ30aqsO9oD0T1fnyiWlAF1vG6///z+CgKpX8dG6ZwmtACUX+B2wxyKh0UpO
JY0IgWsGfMrlUJr+sU861x4zo+sf/35obqeqr6i0S4NRQQFFt9xtHakEcAZjIdIS
eWG/BLT64vXI9rO1PYs5ZvnhjBs34asMk6oef5PlWT4qx4pGN11k2Itfrrsninle
ykvrtvF67TQl9JwVWfIZI3GbCXq+SvbX2igdsayzqjEqY2/+UqlJh3LBElEkoTNA
JBkYC/g4E+7pHm3walRJ/A0lzjrlMTDZsQuFHs2gH/Y5+Hqy1YymUwdg23h7hkSW
3d6wZP4HlEPTLRYMfebcNNmoI9STAq7X7nfsEBSluY/U9jy1m+Tj7b5fT0x9HDAy
myaX+48lhXW3SmEudR0FylTwMZ8jrtlhxo+ZiYrNV3kL/Hf6EQe72EGNCNcg8RKC
qDdPXwq3arqW0LiBhhz9awcmM/KuhsPd6wEJCWAssshN3Zr3OzPIdD6f2cHxc4i7
7yaBMCsqna6gy9UFB1T9x8PIkplkkKvNRWGTap0+sGdbM0qDM/6xaiv2awzOUbEd
wlG+p0d6H4wRviLXgzsjFm645tXrH7HVEXqHUGV6jCaaXeamXNzg4vRhHTooBRf5
jvjodhYJNcHx+CxNXi4rSFkKex8bY+lYE3IJTgjnPDDWihT+R345Cwd2+Iu3UZM7
XY8Qh+WlXPT4/70WnYm3x3Vzqd+oEcncJnAAS8JZ2Shvs5jo4KHW7c4scWTdVF5/
aPhU/dMHhWd/W43PYqLiOJUGemShNtZvF25M1H1xQ838VI6b4iIMsJHwUA5Y6s+U
4dFCDOhuMHk/nNw4OPTD50Ib0IfoPJoo9pYtgoKHPLF+6zlARnMeW7Dl8+27TLSN
O8lzF4cggn7h8qIrjNuzpfh6BznOZXbgYPhC9NoAFpj7VS/qFE3ChISILVqONWMe
z/0KqCYIAPNR10MKe3UpV+TOpGkjZRKY8iUpi7evEaiZmRIH/M/m911C9RigHImG
WJOHNf25Y2XgGr4U08jGALQpG1yA/wtJTNAaLfyPKiSM3hpbuIm8WeiWKZI9hgAj
41fu9rPBaedjv8xOIukiBjgzpvHlLL656Z6ekQ6zxUZlPl9YDErSQsp+XYWxL+7X
daQezCyWR4vXZZWIclNtEmqUGIiWNW2+Zf11otSsNj7xvbCNbVpoqUjpiepK2i2g
0Vt+YJbBYWJiGHfT4pLyUpvLq9IOL9vzeClDqd/5k68nO9CcFXWeuC1PCNzWRSMw
FKXwOJ0IzF5P0Z9kgZJjnu5paCEFrwTQCCtzQQg8vFZMTh5dZm8uws4WTN6w3mX9
Tc4TxcQRgBeavtnXm2f9y/3STIXGSkf38fUclzsOZOgv0CxKpgpQMl4h2BhPFAFS
I47s8MjT7zRmypm5W6Esw7XQu8eOcfWBrxZ+w+xqx4clUk62Vnp4VQbgTUAOTRE0
urF6bSXQ4SgzB+t30TvSvQtWvRvxHl2wY3OuPBgxyQxlzexGN7/t+PeQ+YEWN8+V
CgGS90fdInm30Z46D7s9PJrT28obWLG97nx3tU+tGCq2rJJULYFvHTUHXGLTKAjX
pY1Ai4ILg2GioHotDZ8NhMgVpfkcS61P+PHox6zQSzbzjPxvMk9Q/ORFeC8/2qnb
mH4tLQQY2w1jVyi/SKox0xooiAy/eHbOh/3ypki89ibPBLvSkoKYMTPiM8BHyOrX
SG1C/keqrDRKtAOYy2i7VE6hQrYJ7DJ/QK5oBQV9ccPQyebLJnz+8Du1Wjb9Mmot
xD1zyuBj2ZwNojF9rucKZ8JHv+9At4jPgamwx7b42hxXGGIPz9F3LyD0x8CO6iYO
SZqncXFAhG+rwqfhkfvcgKRSPLO/H1mTev2jDB0tBzeXUtK/0blZnbyetKB9daU6
lPJMr9jIkzRRbYiZbuk1xcfYWqo6baJOlw3xBp3NQe32ovqJ/QO4RadtHYBEBD8p
/9hqoA61dw6n2GjY8XYIsC5yBgeNOg+W4L8LTX8vLDMVXrQww112KVcBo0CutoxQ
UMZ/DnfCDc1lNlaNjFpweTkXtpigp3KaqkzfW470LqAW02jxcEwEQN9lbU6N2dir
OPm5t6SrX2M46pQZsYxvIrgZNYKI5WxBx0J2HYZBP4CKjsSh67yvCNnigicxpDUX
CshZUZ7ouIzcBCNPGTwwWtg24/s2rqU3MYApLViDzGC6DQEJ0LLSH7X9DAEA5dcP
ZBwbjjx1oFrlbTu7URCQ32j3W0nyqsJ8tP2hBNZMszEB6mF6nhlDrP6KeJOrD9Fv
Oid+kHvH+M7LylDntrREG9ZX9WgSKB2oXfH6eho3A3y9ImjZSijJh5Ukv+OzOdX8
a+y9LD0ZuP4E/T5QDJT6jGALkj6RaMgf4wRu6sScMddbLmcVztj7cdGIggOPOSYc
0aMpZyg9wutyANaBLUxqQ7vMgZdS0LU0GJ5p5RDJsCXbFwx0OKJl/7/yvFHvQERt
yp5ANq693GlIrMkTUhQjjxVuKuXCxgR0RMiVC83ryPS2zL+SR2M3wkbLDw8Sdc/b
UDMt5DqcpXgF/4lR9rhmX3cnfnv2tm+jY6tnsqDX7Hdp8j5O0ZIO4eKW09w+X0h7
McmdsZeA/iVltK5zch2iCK/aas/c/UhPdtL6ezreJdOR9N35abQurwqBpFsRQAcH
FWHN610I4tQbnm4uKbPfa7YVoUzbHDkIXZcvW33eHI0z+Hhb7RDuZYGyYufHUI6j
jJPt3gTW3R3odIZqQ4g7LbIBQjM5rIx1giPaiXBs7XbVX/xDeF1q8cDwv8MblDS8
+lR4xEHwrogtNvuu1mJerDq8Y+V4zXCNDK0EQj8w2oCgw2GyaFItqEbPoOwtccIm
CIjqGc1OA1IqcNFIhawtdrEPO+yH6PjAW5lqsvWz7pYo2IhiQJN4P06HXUE1TwxD
EVkVr0u0dVjm3zAu7z+qNYEqR2K8TPuviib47YLvXLDwFglYdI6BgmicHPjxgD7T
BDwgEAPJi5ClA+NBc4uF7TKeoj9FhgfIxLakMHX9Odp8LArqXdw3Kljr3mfSYYcA
4uMOEeGe7BRTSioVeqakeyo8OXO6BdNSLEJmMTEQlX66tRm0M/f2wmIAR0VA9woe
SnW79rULCC6MWOCMCEwsUwLJ4SaOfzMEN61ksPBpNG4XxwXCFN5FFvpqLYyrudy9
QyWckLdAP6QQ/ZaBh5JBDnObciQjAar57uUcinfqqni1OYhxMvSex824I+Aeg+KO
LtoSmJKPUTYQhS4aU3Ya4skr6oM/QDh2Wo1wX/hS0OSNj8pnjWUlSfzftZUE037b
6iw206uJrwWs7+W2u+BbZNPiSPqrnp+3YhIGb8IpfVWqxXwgJau7vh+9ucZwHKNx
QM/wrxVa1kkzWlZqn3koNUevft8CY3zCWAspBM+BKmhMCwFyGTyIofzcXGWoBxnB
3o8UTmF8DFQlQ7jsgSo8dWJStV3C1RH5ruIaaoJ7QAEb2d5jBEUCRoyX9nsA0Hop
aQNcZi/gph3oN6Rm4pNQCe/WiNABQEimAxwg/qLvBXTK+2gH0+LpOOH52gZIbdTe
Jbx0Hnl0qRSeTuBYPmlCxpVo3h+IKrjkq9XEs6XeMZmiHFLFDT3XTQC47Pjn5cbV
c6/dfVid38uEZYnSdVooLn7IsqwDh8ebP42z7uZWsUuJHZOPNjFFtTIVkwNxaqkb
0JHWve6mQRImWDt1j739yzLLMkaik8qhy1FMawRn+uSQVxQDUChYlNDkVkCTKaQz
S4r3kkHAVc+db/4ADWsKU0mQ13Ycufso+rfXRkwmbIrsWLfZZvBf5tP64FC6KxR7
Bp0V++QhQth3V/Nrw6NjRBvy7A6YSIM+o75qtkZ2NfNzQGqJ7g1/0pcOHsRdIzB3
65DQx9cgKteTlPouN+KpMXj++Apvzi3Se77foV7PCeuUa9G8kVb8MD57x5TW+YTu
3vo4IZmKTB3f+xwMrFOXW/z9f5K77EUwOmCBZeoyb2YbVi4eZQ84N9nBVQDaWOYa
TpuQF+F/fX+RaxHgjrZTs922gTUh1TZvo+Q5rwVZXC+G/ZSkAOY5Rm2+09Ckz8PB
UUq6/9EyKRKi5XYDQFiV1ow1y7EckVbwemVAXmD3VMsyLk82vtC/VFsAIIC6T9PM
PpYQUXWGiGGQdFcf0y+AQVhrBuXe8tTXZxzpwjWDFwgWCyQqMqT5BfMZIliQhPMv
4qAoAHaV9b9LmeYbqvHe5QHlYIgaQ3Q/59hkYSoY3gCy2Cb4nTZqRXBdY81A3cvt
UQQklSkXZRm19zji+XUUrxR40kkzVz6J+k4cgba+RCPPP8MklbvnLRzfhVaBU/qy
AnsKnXdAX7FKsN2H8EMn38zoCbI8M7A2sL1SPsEhPpTPFRAYckWQE9zPSuzon6S6
x2++OZU4hiW28ihGaR5Cv75RW6SXdfuHvkanvejtNouTVGQlUy5Un+Bpw+woWsir
W7hsIyGgfTbBX9Dqco7s6jbSUFcP0lvDa6JQGfGMR8hP8+agWo1+thAxFXV5E5vf
2V+fdyg5m55/bbVo9oos0+xoCLewW1Jye3ptfG592jPJKk1kzWw1vQ1hyuQ2Y9JC
7V9R5M0IW+W80PmTyljLH5DQaCdp21IHgmuc9Lp9y5iIfhTR/+Clb2CH0zWbHbc6
surYg4sB4qr7sdlz//yi4EH1ZKI+z2NWCr5S9YZlxEYno/5bQsx2lBOMgJ1vuzk+
CDgYhO1AiVRLKvDbreDQQ06egNuFHaKdEbWRX6JNyK8bsVDRqOyLzOpAVV/7C6sU
Yc2/Dl2hCxhcZzFr5JM4Bhja24BqL2bI1sSnStf8MshzQUc3qCHqoEy17KZnRVZM
w0Nj7OR/IT5WjEDIO/JT7XWRuJ0njTnkGvsyLZYzd6n7ZmwrrbCZ+u9fWpty8wXh
RgV0x3Txu33RnJRxdGnzcFUbvzMNkgAEvYI+Pr1R/srTZsULinicV+vuFZKdi7tg
xBODBIp1idwn8HsfpS5ykUc0O5vP7maQZKiHlc0tAOHdFea2LhY6bDvwSAKAR/sX
GT9y40vagT0VzsPkNfZ8H77L/XBxKPhKmR6PlmdbUwKo9PflsCkh7KWNkdPzLjFF
+fpfmemADNb1hSn625zWVtdLh/TE0m+6qqK/EGCo0dO/+X9lTvoRqt290XRSDnr5
mV3+/pgJbBTLB/2NaHIQsp2HNu6zsweqTNIDs28O4qWNnpfpfPwp+DONCa59KVj/
qZpuuXdRWlx18ps2bCEkJZ7q1oKaddXaWGpM4oe0Nh5h4eirDl1/N00OQwadtMZx
R4xs+oVMzqSg/S384wla1hrxD9uAeiuZe3xqNdE4yeJMnzU2NPvuN1YpubR4Enec
ADT/dVXttB7zwTnsgLNVP14beo9XV6ODbd4+6UkkWRwQVd3IJtpjZB51grqqLOdP
Bgm5mTWjWvi+UT8UoNGjUu4bwqxV/SfuiHz8epLL0vnRu7dok698AlCiJgLDVraX
uK9b9dA5FKOIyF5MDpE/+AXbuFdYLW4wbFit1v/f8yFgOMs0WxARjESJ7LojnfLg
LpuZUujT6V0Sk8pGVMA1P0vrd71jrmhmkx9tHIXv8YrA1wRSoJtaWoUpSh5K99BU
nfgElN6363dlksHyi7Lk7SYSo2WQz4MqpvAT+S/thlXti+beD+evgfmY2riB+tP5
hPgu4cvmhz07/6n8CXZhFLx597Vcd6DkqgPUsN32i8ETYkVYhYdimZAM9H4BUKo5
AjFy2feNRY5lePVk0EgMIZYT8lXk9o6RVq+UFOWa2t+IvdsGsdRdqtlogf71R4BU
qBHqkeoBPNZjmc0Qxp8S0iKu/Rn5cIDgJqFH9JboV2bEfwqca5P2QxB43zNrywiK
hKwTUAddjlS0QmCS0slw80928zQn7trojrluZgOCAPLd2Vdc38wAMaMv8FzS7Vqj
gZaVtmxjNPnAUn/mBcLdvDr6oympZ4hypXE8UDToCTfla8afV45eSvhpr2fsKVA2
82kFGGrNYR2vp23fWdpaLjFezAuQlliSI6+81ZhqWfDFuRcf1ZxjLPYRINkaxE7E
dVDQp/Au3avk+dpFscN4pkfWrhdW80yVsEb0BnbpooZX5rJ86ZI8bKDgKb6kQ45g
MJleQ6cV7c/BFiADZwPEn5VxcdY+kJFA2fSnRREZZ4FtQ+dfUXFjWqDUqoFOIxD7
QOZmifU1cNnrrZ2WYwOXKZgGP+NS12lrHMeSFKWeeDqaehcpehlC5oLd+owcDSq9
D4DrgtuJCRvUaoKJeA/ld1B8Z68uiDd/4mPTg0MYJFsnozA9F2yX/ydVZq1tYzaU
5vvNmgDzNnU3nupKZYKrlgsnUT79OUzgl6vbLxaXHXnRSP0qIG7O8o+QC4WkV0nE
PmPcaud8rWHTfUZKyEUbMB15a3a42IIXRsnrFMq48//waZs5sFbR9Ztl9d/qts4I
TLxrm7deS/dXOWG78HBuRRCB4gWkR46GBPHgKPKg0ZIKDl9esBiC3RL1nE9GN0RC
AvToMgZpGxQyv0ZWclK1M4zTVTc/zuLi5DGIQJVHGx3arsUki70KIgV6znUX3daW
5B31ifk9qgVgAaQAuiFWzo84j8bet11GbJS60pKzxNcU50c92A31J9vzwkxe8Xac
uS1w8bNjpMef3ZH7/KgHSYPrYXHuhA+xykzQW9XuLVgj4GMe3B3c+dtJ9TVUzGSg
cBdiN8lliJlncoshGB0o/tElT4jV0GM0IQ7Yrn2N+tWwrbEslcIBiTrzGkDYJtXK
vAAHwUUbzEpa7gS5wHfsZpGze7H4rbbfqClhECDDJV1MPYY91Kb5dxgGOZ+5eHbY
KPITY3UnHLkQOmzko25/LlUAa4ADwBkaDVVqV6Cw4hxDjH3SlnugShUYsOIKXsvh
68wPKqtrwmAzvJzQYaVW1QWchBnKbf6eHccLvdgkw2hgb6h0ZcPkXTnBAyDnBMcm
8nJ2N4OrvKAearJ3qZpkKT2Xtcbf+WqKCOybMn4vp0w3H65lMA/ePeXvYZac5ZW2
3lbY8VJwMV+ajr3298AxHKW8rthrxlPRAIuk7s1OusQmayFch0uN6SNKY/9lUD+X
7gcOe+eC07z2DRJnJkS9/y1MpbbGJvZVFnI5GB8fn3JieykWAWFZwS7W15Q2VCwo
2hI8RvQcVb3irxzD7qbjfG/vF+2li9a4C+1ZHAdA9QZXLzVDtgvF5nYbL7co8Y3Z
t9guys/SXR5S1z9sXaEWn+kJlmrvMHiq23WVL/4c07CYrXUZWBvXTd/kjNPK6LiD
tLI7KPgmpAqS5wvPbRWhafPdRO4aN5O5nSDBBdCtZBDADSmgU0t9wXPSiPkQlFPX
roJgS6VZvE+xv4n0+p5JErZiF5RxbtSEtf6E35p/NdK0ReO6WbJ6iI05mfobqJL0
7FXrypkUTBExno+48AVI+xKN+fl1BBj8Jk3UTlAC0xLjENsI8KEZFbKNOfcSP9wA
83C0MTSiAJ6crus23+M9VCfCqNRNkUfKoEN7F5LeSmsfmzchpguMou2nvYy66Bst
d1BcQ1+/vwiJQeLE6luibw5D1R0j4lyA6DK9DLhOrt3yHFKcTLWFmn+eBVoVLoPL
brj9pn6j1TWjdLzMQIRxtjHLnHpqw9Zd7C3N0m/mVLK28HhgX6KqxgqLyzoO1owg
Awuxk7U3yYOkAcJGFsSRV9YnkuWtJv54ytFRJz+orVE4Vis8nQnQqehpPgNiBM2/
uHIKN0082rYCDG5sOTc8qgjpQtal9Jq5oU9Q1Vvg/91061AJYS2PP2jB+wDpS5bK
eQ1lk3U7cT27Bp3CTi4AXe+NIqBmTM8lsaXMMkZBr5HmbGkR5qBd2ZcNmqkxUiMm
sG8P9iYVt44QRVOfLthWbC8HQfgDPof4JJ7rjD4L1IuyB9fLSNW6EsGe8a2YuCpj
cMbvEHvUWneY+WhfHVf5NVSa+hBFatPDPHa3wZypyipv8f5VFK3+vGcj+zVpDzg2
N5m+tb3QrBPPJ+J4+6iv7ifhzu3PGtJq+6NpYJ077I8gvmeG8RJ7frqa70PXhlA8
qR/iidQUo7dLibgCvRkD+M+F5e33+6XsXcikA9flEUwC5vokH9db2U5XtjAc+Qbv
YmJ5omdK/0sgOsyjgtprjg+RV+YbKi+Lbvo0w+M1HnvxY564DG9hwb5zgVq8BdA4
AZHrOtUWeGQCTqaEA5zT1dDtJxXeo5y9zFHaXu2Z6r4Zn5IU8Q+cn3Ue7n1IkikZ
DJQmLwmCZ6XXD3NwpEP1F+SC+dR5KObmNuKgfyvB29CY57JtMADIQEx4CTPLK4P9
XDe3tf3Gtapn4098JoF+sDfsDJ+ISdxvv8fwnF+BqjT+Vtk2TLjSeqSpISSeIvAe
BbjFtCnSmeR7KtfxvZ1xu3s0slUzeVvhg9evPOSFviZwaSz86OJ6vzbpTfKR+mjQ
g+tRi3aHhmij3P8uCBslCo64kT/X1rK5ALlE989cVtGev++b2avSLS//k9pw6gCE
EuMse6ssNVAux7SPlPb6Bs/zx2irv52Af9QiX7/7/THFCjW10WHMcGuSTp2eLNM2
BaChHWjRmCOvKk8PE+fiI+PC6wKhE/yjLwDGeRGxLHdCtTa6DH/p6irvu9MXxq3G
oHz0qtUsCobMGaHgk/Sk/bAfP9AHy99vJxRuxU4j2XVu/oYGl0jbVENVlS+11phF
jjwRItZ/QSkOQxW0FKvRoUvxxjR/zcwYP5q5ooqTu1zx1aHMiwzHoZJ9w7boGQ+z
2/SR5Dl3/7zaBJP6MeIoFKS4nEEYblibLGJ3CCJHNcWJkM+jTe+ldTxIeD+lOsXM
1EBbIpACDYn7pdjvGXrGZ/69p2A7HKdLPZq4AcY4vFGWp1YESFHmzwR0GW98fO6I
xJZml8kU++1B9P7oezSoYGtlVNkZ1BMyqId5cs82M8cY8GmWeV544/jiictJleUs
w1PP83FYmEndduM4Ra7lU9itUZSnDsMYAwOe5rS079qMcsnaAKNOeklp7w4q89Uj
TA7s34FOrUuiGOIPLvpPMXSoN28Of/mix4RnO48tJZQuq2tQbLzRuDDzmipb72aK
Qy7uJs1z3V9Y4xX2uuKSpsETlYix4CSWuSFujxfFLxmeK4JX7zzDbjy803BIY8Er
/2MNkayQl00Y4vOoIPx7wKN9z++SGEsFGfN7tmDBnsHRRHlg93EFxghmXl6oHCOo
YyG/jLtS+P1rPw5DAY+vV6rGZ8iNjh1gqdLMRijVfhl/ahnmF1Ek8gpdYyb6co4e
8YsAS2pHH2n9Rc9IIaCMl4TsxaKhGhDpoaae4wyYUExtOGYB/aWXD2svi4xr438N
lzZ3wHIKJ3/81EDclBdNbAiSqHRUmN16lXOQ4kD3oNRDRFJYqdTqKNtCd/ZEpChc
rbrsv/mYFlkMXk7LMTd/mqmZlX+36/x6gISmhM86gvg3rkm5KYRI89HLS3TXp/PO
crNPSu56dtbc38e6R4qvrjmrW819QynyGBbv+uyc+xaZcWuDtCtypOthjUl7O2D8
SeH8/WcKS0nQKRAVWnHgT/dZV92d5yf8V2V1VX5X7dYK2+n/LKrsNgFgswDjuQNX
EhlyEuiQ5onsCpprMZ8ytIuFi1x/5lUdO85lvOmZDnG0ogmWiurQ6+mZw8uljNrn
2XdE39/ipTqoXCqJXZpgt09+PG3sv0cOxyO0Yc2N8/7zGU2HQ5tRHZFSgW4KIrBQ
AmuuJ3Opnp7VwEfKaKVMPgkAT91oeI6tqbSsdoDE3JHDsVv9SRRSqS7wXn01L+c2
bJS8F8rbFLIM+lnivB5hLNdeUrETRC1dNIlPP6S9NgYASoOfzX4ZZa+rmOtQ+Qo4
F4MjdKhNSIFWZUkodQc9zRv+bjEUilZZQ/aTXN9NcizOyP7rVx0IoWfcHEvN2atU
cF5hjImNsKXOBAyd4XHprXGl7uKwrb2cofMs1Vgv0TODUrxMvMdAn8T/eE9+JPtq
Y2jmwueL13lIw1OI7xbkK7w1c9EQUEbtxLOphQfp0AN4LHY/aG5WQDdE0Hay3sQQ
+8rEuQ/BSwc+AGAgpzxk7CBGRhOoZytOsQHmBf7xYURb71lzUZ6jkDP7zVzZZhLa
G6gnkiJ8i5oKc6igzwLHL7gJF5TU4Gt9fxBf2FEZ2qN2RS6JKp1wdIOmUYcz4PWP
2yPxf90sbfRFAaLmSXGqu4/pNWfVtFtYCxYpTL0Pe+FswelidX6fL7f6wfELTPf/
XZi3eOJbRMV2FGXxkOgFCYqd3E0T4FVCN+N1FpkhYCYLitZ7XPfZ+/4H91n0gMkZ
PTMG6phqk/4ykQrNU8LE2zQUU4cdFO4k0yZsJRp4WGQ2sr4v9dXDRrLMGo8MWOme
zsBGD+/UR674ouXtWHnEILP5WpX9xyQRsGilXlL6ywHyYXIhb2Lnv/U3WqJGf4Oj
PrMUAIbN1uSutWPhkiYvXjoz1pAuZy/K05r93ZhNfXch6nepKJ+Q+Ci5CSCTtEXx
ZCo6rfCcjqAOGDmrmVvbrRIRKsVRJJTEEMugW33fI8nU4VOcvDe/zzyOwRZuz4jR
iUBgrFQCyJGFrPeAAAjS9UFBCBituQEVQJjgjECwDjU5y+BIFQBFuFZWTs+sKWTg
T8NFMPhFffCrbaaKR0vBWaySLE6A7OebRDZELlD8ATYUME2YvCaJRzrfCJ+081Eg
QvDiK7CWF41VaoQnrDCkciFgBZBQLtgJ5YScHhOdCWduUmOd8DUt3Q722LJyVYVp
35/T6RsRC2v5gCsBiL7W6PiTsYCvKCThNMbKqyTq1mc4NSANHTaOxoZyOsAy8IXI
7MIpIEfBnxSEIdzQt7xGXVlPOnKnETpIbINttqNrIR1ecfjyPv4AWAGzCbHN2xej
El4imGGOvPSATA/czxRgrc0tryQJvfgZSavuEJTvX8XYk3ogJR3UY9vf67hQhlWE
Sok4n0Q1n4MK6DfiTyGtbAIVpCXH5lr7mWqljBhbrpcUxoGsOh+1nLjno9zPCXDx
Q7V2S92DkOcATH7qJoP/yM4Y9miJGkMKGNDkqRzIfl1nJDrn3vWfgkKIE2iW7r/T
4SKO0q4PilT9/8P9Nkt3l1T8otbZFsBVTWCtCdT6GplwCmWub5yIYztybUtD0O2C
jcKt8DEpRv5QCPQkGSFSOIK6skN50JxFee1kaMUVP1t42zeDdOUVBMxeo9d7SIqd
DuPmFy5qiM6EKc2G2EMFJzbZCmwT4XZoZwHv0K+41YGF+VTliyj1jBK3/jjJY51i
1Zf+nBnkOlTbEuef8Je0VThB7G95jXPMMYoMkmlLFvSZtzD51TMj7SQlMaiUe3Bi
IaDpEQCyWi7ewJcoPaQgSnrEssaxW73OErZC7XjUiPzUuV6V5AukNdz3fPOmpvv3
FkxXZGoJMKOYDvHu6/fRqqz+o30fpjVn5RAPWwXwNukSAWR8a28jJuDKI6HvDjPQ
9kNu2pOyueoTDeC7BhiRC7mMfLHoeYr8GxsMxjFF1sRf6XGf9fMGCE/iKYc9/shG
U1xcPNlvb6cT5rBQ7iwRXlE/EHwIi7NutKJTFT2ce2rUp8drHXBRrV0kd0jgb+2O
m8eBH9cg3ISPC+mkj7JINZwH7SEhoPkZ4fKSQrY06KrTyN+X2TmSzBLmJPHvyk4V
D4tAXhUEdtR0sJf8lTHpNlWMdRCu+zXw7WwGCsEa5PKQN1E1DSJZNV4CTxGnc7Sp
DFT0f0sNUX3y2IH35hexYuqCDo4oOk8mw9IJTXcvtxISvEP/O6SiHq8lU8TV3Gp5
PIZ2ueFAHdX99G2zDWx57H9dpVQcyqEw8wHilHRNaV9bDnUQ89nta8Hy5pOqLyKU
vq42pTTyuSpM2L1IQU3Cwv9vK1OS0yTMnx9AyWsMB6LSkMjUpwjiB+KjZHiQwwS7
uYMgEKV0hVqxDtSh9GaGOZ7uPbTja2+ncj2y/YpySc/8Flq74h4pUD+HE5pN2qaN
n2YHVDf8khRSIC3e1JqJxsHhlkGx4oOno1atlx8Wf1isx/bez3Sb83rl4uEaEGMR
5Ts/9uASvTFtWR9/XGqKUEzvOhPaCaCa8aHD27erDsKE2p+H5Ba+MrD/OO23zstW
2wT7Tjk259aeCyijmGrDIFOOrg3gkFqw/6XB0OzbXTB7FZO+OkJ9Vozi5SKQf6fO
+vGAn0lGS9FwYhHDDVO/HT6RqMgD/XEjKN/P+ngogddm5JlMqQdauG8eJa/DLb7x
WXINDtQqbQ1+oV7ILUrrHRzLFgf7sTYoyuGjzr6A0DjsDvfj6H7NoJHRVMC6z4Gs
PTPKnHNFzz9JRdcx0Snd5Y5n4qnVjL8cdmS3Cu/rkjxGk5CzdE8U4H5lT/y7wsNJ
lFWONMj5cbnKWSVODWInj7KxcZqcu6UfOrQ3NY5yl8g/xitz7PlRbAZu3eLoXW0k
gJdT/332J1H4TDWdaXPNlPkSL1RKMwqww9ksfxmS+1/ycFoTWzD+14kueToQZ7eo
mLL9bNLP1b0eGngsrONOk7jkPPK7x8rKFHXaWwhhY2OgI/ZgYH6ln2Omi5dpbCg5
5oH1Ni7C8fsQ7C2FUuJLcFCnIfHycXdY1U4gaaApG4ZpoJ8UhdzLUdwWy3pCHoLu
whdk7IR1RmNS6G/Jr0tNRd8tHgqhOTgD2LhoXcOZeFXDPeRUhhrahHAAQPqKI6he
JBSw+oHUyq1AXftbDGXgWNc0c/PvlWxquAcJD09uoMmnTJb+RJUN6hc9qVK1zV9f
T8suGLKYtDFoio+6O1vWy0pZkQoV2d5k5v1zu0cg2MY8nCvSk/rDT/CwvMQWAmsw
h31X3gr4WqLp+iTkgFAwz3HUdYgNl7uadLc9CVbFflcRIa8PAabdZX6g56WSUAiC
gUyCyLF/yDM09C3ahM1vE4gzs38630uicJIppe51bPs3ZZ/DQzVKzSAg2HsQJgWV
14m/FkDhMNutdfemjjgtGrsnFn1MlOI70HMCyjNYLJVWuD4PKcdItUlxbUDPA/Cj
XrU0om9ngTwEfgm1Ec/q0MOoIPSDlu7JF8GvdRWBo/YmuLgkGmEZuGFazvOgkY2H
rmbWDAbEcPaQtgzFdhbf2jHtLQiROZiVkbXzqcd0CiiV4JgwRY/taxsbdbOmcjWv
oMlNKxh7GFDFCs6AaCRoNu7Y6mileRkYH5pJYkJdWLON0ya71EPZ/VS5MyuSpbWa
+VIJhyrIXJGRI85gJQvUzrZRln9r1/XRWE4sxalb8KdCl/2Mu/56LqMXpJRYX9XU
kdAL0LWhkj487LkrzbEJXkuRmQIzSM+mi11DyHUD9SRVERPvufo24weRQz4SlTIg
Fc7/Qfz3gWNqiiu/gTqdtFgtmwKyXKGDVtYi1Ju032ZvK2+8cl0Lzw+AsB/49bXb
tr0gB16/T8GkUef9uxzuvrvJMDNsYln1OxRon2GFlaS7Ig1qsxg3GRdoQCBNdmxp
IM6Cghs34KtNOR3zQwlBmiaPqigTSoopKeRBVYkj6A7BAubAxxAdqCr+wddzo3NY
jH88oZFa3Z+47gALWMv/+ZcOoZySOxw/xyXh+qzvpU/tUWOovowbKwBdAsgT7I4k
WH3//pk2kRq2cN0bTRwbiF3i06ujL3+y8AtKWDIBMm03adbHRonI1aqWMuVaHnve
yQEAhZPay1lgu3u3erhCpkWpisLkC9bhYok36JiBpE51IgCOOzJcr0eIcbJM1pfT
SVV/Oln25m1XphpxBO5nJsjbShhAZEdvTAsUqzzgUHVwiKoJQ0M67HrvlYASHNQn
vl20Ez0cxx+pyMEzWFPRIXbq3UrDLW2xz01fpd0xZqRuPVGEtJ+zQpYmayE08avB
OAPjwJXZO2qsnoytkCM7bjSrFj0i9pXdxC5SiTa0+DqMF/Adt8H8s6DgM55dcLg2
LIEiq/3fWuk6vKTIZZNNE/wCb9/hLoFK8t+lo3ySWLsc1+DryVU2FLu+uuYK9fCD
MRo2DnEsrveeBrDSF4/AootxsjH37dhVtGFAgnyw7vrT9i2VuFMP3vDtC+KheRSW
aN1NiMQLPl9gcFqrNx2R3C7Spq0drSKmIDY/xj4VprumQ4PkfNUPlvTqa4dX4qpn
HCty+wjvMjnywU5ZwONDjGC8bEdnPNNz7f19TvzpAu/JfDu6AgDYyY53wFgYvNM0
OYNv/tMkatCFI/TtEm6VTyavoYdyhauDRlrWEJkjMmznNT5jMZGxNlV2zSbMo17N
yjDR5pUhp6p2u7LEEp3v1dEpiY2Kcco5Gjmo/+HEl+tQ7VJy5MFtBdp7N8WUenb+
3WGmsGC8O7iwLpWtHOEIBb2z/GWBP0hvvOCcI0acDjoOEYm+Deb+kB2fqYXofnCT
JPnlxCtaBhmhUkEZa6ttoPZObQcT5AEptIBt4fRFabb/8WrSw0/kOQck4TSE1PIe
LNZE2NJ3kSHD7HWYdDqaS4HFHIOGBQSMXvsWrhanMZ4EtDLJEpIBjtalntdfzivB
dt04y3stvr/fnAJkA4XC1LFNrRr7ojFqEqK7GL2mfTdwJco6uISrar/0qMQEEd3S
Yzw+4nuTXYEjBsjabnKbNmMGF7U4YxIA6JonNLFmxnE8MHwea23ruSWWKLz0wI96
qhTcigpCkQYrnAJqucKOsZBO/uCY2h2ZeaI16HOfnOcvkRHb9mRF+5bHeipqgK3M
aoAlKbzgFBpYMdYu7ZT1yzNfbwXJjQG+u9Ui2PDJP9By1YG35SmVBQqq2TMTqxuB
UjO3XpshmP0ghk/IH21DuY6fYcLgHRZHP1+cpQy6TCJkTKMp//rgW3cpjTM44K01
rk/dR/fqNiTT4EB5c1ZxjtDH/csOQ/9zTOsA16kwak0pskEvNDDcDtugYFAygFcr
UcbtvE6f2oF6NCJMWyzZZBcR/VqtxNx84QQZAnEKN4fHLSGI5Yfo7ALlwjfLpwSx
KBdPFn77A56lR11d0hcdOO8AD59oOQ0oHnqRLYamisiccYe7VBa3+tPCrBP4pF+i
6T4PujylzL/1XU4vWBlBdqJEOQ4OO7FxeaXaQfv8NXIok64w9O+DjwjunWGELvRU
61/mo5OMdoWr586+XOJ9Dm9Pt5aFIevuz0OomMOd7vJ3U/Wyxea6avKc8KZnknBm
pMiFY/gy8tRf3NrK1JHmCnJdeL5yv3n/izyZbuTzLqT85oa8ljqnhF+WCvH0xLV7
FH5sNWSoH+c84UVpElWW2dQH8iTVQUwc37XIsnq0c7pRFPtjd0hFQoda2RB+z5hl
7oO8Zerwg23uuAtmwWHEINijEbk5DE5hhvj0JCLDqu6x1pjlIrlWaTYayE1OWqAb
P4CEkOSgma/pTeWyEGJXVD4Xp+GeCr6Yl1QCjchKY+ZyBBwDT6P5SM2/FtNAVeVc
DV7mlT5M6RUGB/fL+J8k8l9q0IZuy5j/GWq2yltojnsWv+iqAYcLfR7h0OX2O/dC
SNsh/Y8n54mQOOWVUCs1lubwKnEkF7SOedysfXKMYcEPrIoGEv/TJ5A9/09U0oAz
fTCNFzuFsOS/Pe8QBB3aHvs7e+9zBqvimy0zpzje9uR4IxuTWY5cPiEjNS700UtV
NxTPmTgNzcp1mLTWTIlStSzFLntxoxVFAOQjrjYA8TDRT0r9kfTwZdZ76QyZYCrv
cyAwCT90g1J9ORfLdyALIlmaMTYGyqfXmAx0qxfQmhG1HKfmVyOEUFgB/vZW1srl
2ZPONkEQviPahBVKDRTBjP4I/VmpLCoCbEbWrejVColGM0FlVZhxEdCqxys9LkN1
jRZMnm3km0FowrAg55ma3oztEBAWNWZL9CvVcp5wkocFDSNdZrgpUcM84EvpSNxx
R/doh6wRe9Newr05eqSLn6ufdSqXsxpCIDrYUzZTkxYMNRwkoTzKvqymWvpnqKUx
2lorIlMEFATYrko/UiReTMK4ljJ02etHfBh1rzANaI+8Jwamxyk3idTbj1ngzDSz
5BqUEZRigBxe0k7QHeq0rPIKtpSNeSjZAJ4c6oBasjsxZCajIJKv5QgI5ijjyRaq
lbEQHf07ttEJaRSNyCxiwzWRFRnLKe08aKvz6ZsL2uVlFOb+IQ5Sez/zMozMy+Gl
r9uVMCsDNtan1ySvS/nAddgC5GKb9B2kfA5RWCbipwRs2uxSHfUIGxVY/sVGIsQ1
rwu/v1dB9ycjKNRDLApcbW7sVD+eLolQ3bYoon5YPRPmbRP+XQFOB3b4Y3Tn7XZs
0ADDJgSO5g6S0KkbuLo0NCfyc9dyYpWi20xM7ei7U+//dqCsOo9lyi/pfQoDUnkm
wHOU2z/vrIZFnZxMxn95x8yS1qEdRDYqVbVAQPGQNwzhwbfswLMTP+wGD26D3jgH
LcRg2sgzAwy8Q9ENhfUhOJ/14O5TcXQhhtuMqC/L7QXRg90knNBbZdYyquSARZCZ
1jNsJXKRWU337KLlTOFgMtapVnWDF9WEYTyozyDoqVyv6tAdGV9f50jsPje03TGl
eoru4rEGqU2YmLLLBSE0oJ9PZ6WHLQH0J0pVEgtCFo6dtySBUXsRgJmkwItVN2/8
nBa2HtJ2wC/tjz61gClbiBPUm20MKvD+LLm8/087kSwSYLka/5svm/xqYL/yhzxC
ucH9pSUP21t7DnL4ySyy3mS8QPsAdZM/R+QwCSKshOLGy0CVXTlgPxbd6J52AcqZ
9dlXxoLNZxf9KYES5NDa1xhZB7SGnjPm3oMbmEDDW4ToVsMM3BIbCxllSQaWRB3V
xXGiBZQnjpHEShauXCb121eAQos7Die301oV4mPK24tmr7F2f2bajUWrfETOFSDA
H6xuAlzAicRnG8vrimgQk7+CFs4JL2R5CVy3BNlQR4sG7yzSgr7+wSySCnRmAWSZ
z0JA9PhHJ6c/y1/51SkzXCenEr9FuT9cJY/+V1m/XWiy0z4NOr5ljFq02Gic/3Wy
rcX+KyYUbBvkkf4OgV90cEtIC+RDR91aEX47jwT3NuSPNRAMeWyQEpuTPUy1MGXv
UqAlycp+UbqbIsAmUIC8kUA2mLSakFei277MnxJJD6t4KdGqTMATeHb6EQyatdnF
MGuLxVvh7IGexoc2RpT6LX2dhiA1SeU36vEcpRAWVOkO2SA7Ej15m1irJwjPzOQ4
0gMvo6Xzf+7F0T1ZeCoRwTMCU86qH2GY4zmNYJqfB7HBzzxHeV60MkOBQG3DtsqM
c2HLUAejZ/t/7yoNZ8JWfm3F5ghM+i0ThWmetgz66clHoD+Xf3Iqn2bPTrLX1J9f
IdeCyrWe8jAch0ilfD9XBEyeLHqwyuqvGTMqXqtDtX8z4UhL0qmiM6xNJa81ba/W
ImoBkIcsDt6ERjuUBG8MRYuJlfI59AYFjzivNeuz3EHFhWH/e9pOdDGqUFxmbg16
I8C+JsM3MVZkxBKAEvBV/SwGoYLkgoZfQwmcLallczL1BtGF/D1W5hqaRX/RAM4I
0WA04Ip0R38x4nzoG2RzQGvUlsQr+lfx0FDKysL3zO8aYs90qTOxwOp7HI076JRg
0iQcSgz0DIJ6Sb1Owv+cbg2GZd+HMugBwT4pdsmVwtrm9aWeFYK8DQ3y1zKY4lS+
HR4CJkjqkB3jN+MzoM0/1e8H2W3hMg3Y+suuTu2iucuV3d1EBjjV8B1r+/loj6vn
XujP8Wbc4HZUhDIYct1ri+PvrvCGdqGKFPUxsq+t5zKep8JQne/r9rT0YH/5jOaE
ngcOTex38d/KU59fuqBmOj5TcJjcEwQTDiUSwMI39Tkk301ET6RX8VWFoff9Alv2
YJ3BbeMDjes/XcpNeLfVvdHumB7Mju64LIHuXUqt5VhPu7+REeEWpYsl04KZDydw
kVaErJypqjnqxtB+a+f8idSs/lt0QbiSfSKUVU2Vv8NIzIhk7szkHcRIik6IEIMw
Mubw0qvVN5oMkwfuR3egj2pzQT1IiG11p/4iR+zYi5fXV00cM03nhe+UrdXZTbOp
joMOFqHA6tjwA8wy2g9maJwO/MAgMeDPopHcNJgZ6PrESu+K2QCZcF7Nu+x9UBIb
oVFD3MOIwAJaWUlFLJB83/gmAFSNGc0cg9EO9Zidb/chH8PrqRfGeK0yXHju4+kS
EyGa4IAGufJ8P4pMYmVsKLPSKenOnJ1gziV5f4ngwlqVS7AOlPyPIsuOTd5CoNtT
p/fXI6ZBJzARfw5snx8M+MdAWvNpi/E7S4Zm1hCWnjV5OW8Go7m05/yLVannnPB8
U6oI0IlB1DeXw6MPXw23A2CQbd/mJtF/Xmi3xlOAmrLkr3S8V0rkpxRnwhMI/eOf
RfN9mNFfir3h0g9fgUTRFBMNjpdR/HskHzhEAyiHXfivAdbm4NnIRFGJfxuJAWhw
IeBBF4Wk8aYPCdO0LjuJMmQENNE8A2myFcNDUZHBrTJPW93CAo0SqwRe3+NEs7bW
V3Klxt7uj+iaGTejicmCAv9ajFEKM+wazoMRYGw5BZ9va/ORQv/KE4Xj8soos86u
3hF7qwhw4aFb/cOcGdj8XPCLK8xw22aC0G7HKyoNGL+vZqQAw+pj9ieWbKw2YZn1
+Qb+QwOR+VWFLMe/DKn0xx8dG3AZ3V1yxcDFCrpCeTO44EtuxbixqyK+BwlRCaNY
M6cjEiVMvu5uAghXnMFzxcSy06ftOxyBlAFcvIX91q3+f03hCSfoSY2DHoAcEvg+
R142wXxS8Yki2Ln6ohuiUwCVJ2vJ+W66YgVxID21jsZO+azOA4wV3WboGJXBdmE9
NXpC65g+YZ3vCrsL4ifdL6gmsO1u25uwJCa2Mj9VdrInjHuby/WT+qSrHvDDOI4q
8IKExXSpCev4wiCNwsBdwuM4hQyAaH1NBnOcbnAuOcJkPkOF1Q+Cu6XmG5sqgKep
+6QM9DQBENhv+7TnEOguH2DwHNSrZ0KndeZY+ysmUR7hk2927+3tfONudyjNp6ce
04EplglchPyP+aD14VrXoQ4VyHJmsJMvRcNEC8Sf8HOAgyJ61teh7Xup9KyLdxDL
2Qz2T2CjLxPHgL/X9moF+oWxgb93lRxFif5XYcpPRaO/CQBQUtbm68+SWBXlNF2m
eix7eo4V5Uoeg4dvR5XZhOhGPeNv0VOf85wNAj++YthXEGMYRLgbkA61pdrkazvI
NL4L0T4cLsC1Xo30L5/yAgrSsj/C5O3HRt0pRrqHDvh7FHTNjv9/fmh1b5hNKYRb
`protect END_PROTECTED
