`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dcd5uMw64VdCsgjv7IS2gAe7+MySVrT0DqTFGr7N4smLBep0yUBtjEJaQBX4nWXw
H0R6BlnTQehbTKON0fw/NpSAAAVe2Z5BVkhhx4bxPzKqX3kCtDM2bPQu9KO+0Ys9
olEshReP7T3PJUiEw+N698QHDQaEca1IWr0jzUqDfTKBNr8W2fxEZtiQ1YPgcvBL
WJ5FBQucAjLL9K8JeKfvJPS65w5OhgXMpTjgqma0n9lmItMEu9Qn91//5Xe/WYH+
1yOjHxyDAE2f3BWbiBirpaTk+QTJ1gsmylZP4mefWHhSSgFGTbnWrloYD8ftJriu
DEUK6kPf5yd/IzhfosiR7n1Xl0HoNvqIkVCC0oV9bWtRfOuFeg4n17jqHuQxZWSz
1UhM2XSPLU9LNxgQHLTtu7wE42iDlBS81WQjOlUqY5D98DvOmVfdMw7jsK/0biPx
yjc0HbGbCiN4KWJPRHDC6INy8srHfS/AT7MXiFcNInMk5pdKXX3ka0gE9kq0Ls7B
JEPbqAKshPx6f0mxQbMMxrkiLKBkx2a6o3EW7lZ+20sURNcNT3VfUlVrq/GHyamJ
xkvIe928sEc9OU6OXlNrtOWO+samgpVs8vYsmNYpZBwVJrAMsdUJy2OTR1Qi+dqi
A3iZvXNFrPbsIz3Bi2U9NBPmApkQ05F3hHU6u90D3dBRAiX5W2FDudF9OuNpf9bH
SJlIu13QKB/DKIzh3lIZq2jXna5cgICqlWodw0xCy/DfA1Zus/pLgOwlaz8mCYjz
EHw2K18gcgsA6qfGCsZ9JNzbdIsYGXPTExloXI2TSAmwXwjx6CFotYtnydQtiC7k
jSwRj9npocdqfCruXRwGZe3SJBr8UvTWnr8N9IXO4ma0DPQV8zJOqJ2B/mxNW/Gt
B0ZKPhyW1CM8J9RlXg19u5dayEbBwb2aEpM558Q7eimKDCXDSo1WOjdKU0bEdWbO
iLGndhQT10tZuDwtkbTaqNjeykAn4apOGQT6CnHR7KSmSASrvu2XnTKQEhhILvj6
MEvwUsWdOnllgH5u1cO0swyKQGkV6cH+ymyQDERx/f1FMqMEPRN4YXMlnIzXdfsF
edzffMVyQ+eRxCMWCwvZM2hGBZ6gzfF9I0/fGW+ZrKEyFtMHX0JeXEutaaKiCfrB
gB4HA5OlUvRENeUFBSkTk3N7Pv3+Axux7PMSMft+G+rbhZ7aJ3ZxRvgDsZKQIZH7
ddQhe69tNB0IY7AdmMVymrWbOJJZxxwbLbc+OFIOYA+c/AHcMOUiMcW83/scy3vU
rvMJL2htvG2FiKpKOmZ4m2sy5CNQp95EUyTgyk0yoQY=
`protect END_PROTECTED
