`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O6cVKJNlwGS+REeTwi5MvoL2a0FjyQnTrZwXEI1PQjjOpHsnd0SaGXmmJPr/5EGB
WFgCO28o6S3i74p7kKElQ7EeQqy6Z1pop8Trkdu4kq+j6fch+S4IVcFH2tvGn8Xc
lUcnO1vR5xB4fJzOFAJRfCUu8zC3AiSKk9qNYa09xblK4WaNKzrksh5xPyEew6eY
2R3lJl9s0p0xpZD1td2c+CG8aN0mIk+YEJ7OFxNfw/LENDCho5hmvPaLOd1+AIPj
SLgXpf9VobDFtPTcRxx8c0JY3KBztZpFLu6ZW/8+4l62KdzKcHcavf0dII61bByE
OHjhXCYabI3pA7ODY2CnktQUO9VuODHco16BB2ArXGZ5H3cLgdWue44E3+OxB82b
ssfYa1dS7V6t/kHw1oxXppe8gU4zzVh4cZHuic1AD/2WJVGyeaZDeBof0Vtokzm7
jl5pCzSuwUS0QoNYxAJefovvFUaoDL+m2gkLQIyfmx9cK7mq77IIpGUQeoa/IPZ1
GGRKEm3yosxpAef1HKfH76pKwlf+4pmcSbHVt8RQyE5y38H+zXZX6sgGkicETNI7
yy+d7m36aY3rggOEYJrlZ4ODk3y0qamBdeu51xHg1F2hEmkYQ3t5JGlOghkOsYoL
hnQV+NjxDva1GipYquifTDuA3ZHrzVYEUPWxKPUKmgv2fq61/KNDUTOAY7acxmCt
Mo1HN3onLHOBlIoe8gSj9/50oK1c/cf0/D9oLLhck/VyerleGIawv2yIFdwCJz5a
Owwu7l6p3YS2+2MtgVRKkwkQrjd8je4AOldPML0UgsPWDmCXQOyydsSit0NcN09C
RfbxPKiMdd4Ja7aHnbZ+zi6HznyH4j4UhXMcD8HD5EVWiLpvXJ1Ae0IpJHlXRNnV
sYjOn169VrapozP7N+xbb8+3wKkZSfhP7jCSem2SrSwY9puLlGX1/smueLrfwXog
lRdDOtdvc528epJxpkSwPhMV1tSCy8io/yEPABAlivo4ACgXZrKHB9T1OUa6Cw9O
DzNJ2eDjaJWHzxnRLpVzsnyjUW5y4JP5K+a6fIikfl5bVGPJ1oiGrV6XL0i5BVs1
PwJtWTMj0zxoiRcFOBLryPdM1i/cH8Au3bXxRg/J84Ssp9/uzAATnVxGnB9JUSbS
rvUvqFASyP49fUP7tSP4WnGf8HsQ79YYdA9w8y3SDtoDPXcYTipwuWT2OwbPm3Ra
M11JhCfr8LTzk/eiTFGPXhtroWQ8RweJQKziE4mJFuXqAai9qBY6zFrCtlYpkKih
3/taG5da817JcS4aato5b5KPrdG4ny1VIP0y4tLU6ydgC1iuQq2u8KYyZ6aBhqbw
mZ1eP+jQAW74C+dDzQLca1UCwOqpztia1dWjvHFnkC6SNUOi23rSZFZVL+2Jua+f
zg/wUavtHKWEnDxHNa9+TIKDqLx1dPDwXGwR9Op0i3sN1gw4i1r5FRGFRhXmh1MD
G076uusq6rLuch+R9UBHaXbDeToWXFywRpjssPu1za0hkMSzmE8BWfdeDGDwAa4e
IMn/9g/Ag5zNfD9sxsS59tPgvsSleiB8nFlxFY5XqjCJYXL34xfOkGCom7EZF2ae
E/qwQWhOYRCYGrk5paIq1fE2ERL11kpUnhwbMMrCuBwEqNe4Iw8JlQn7WB1rRM1s
+A3rbHuw58S1DT+g/9RESE4+yNSSwweW5AUrpvPDHt0eD19ZJwusbwrlkvrGDAdp
apoRuH4rx6gsgmdQqz/wi1jKHzc3a9WC1+Ljkt6coGKIaIMY1am5Y9OwEevmyitx
o+7Erw7DXU+bsNVwHp7rEm5AqMIDMhg2V1Ys9UfkmSIe5FfvO65j/AjPAh81EuKH
xW7LmV+KrrCmu0L49SeUrtGWc4h1NiXPCgdAHqV88qfAXYI6QUCgOiFEQG1qiIZM
o8k/hBCQNmwNqC9+JUsWBb45CMzSHvejtgfNRkZVJAOJeGb0xuTPYFP5FuOz3S5G
ELS1QRufaRAlDorzAnaR5MgU2TG4+ekLKwLqTCmbBaEtoV/SfkTVxMOmo5Yi0HVH
WziLo2s3sUmXJalGBUQCgE71gVt2kgw2/eHP5sJHJXwH/XTUv494LBU8XOz1LrRG
HOhvvFKXv+ecsayei9GOCLU0FVlKbeX1ZJaaS4i1yljPlQXIVs3MckP+l+ELnvhV
WA5pK0Ml7M8OTdhqQ//+F3HBNUf8SXF6JEIfNpsEMkJa/O3w2WW6UMqTY4tLBBCa
FHaijngui0hfy6+vuunOZ3RKS7DGMIMBZmtaCbQZLpTIkqpVR07zuCDuPXM2IASN
bbMMDmz1ycMt0JmE1PUUY0hGQpyO6YSaxheUQ90vG+aAmsX7rQdUO9XjRINFY3h0
5/Aan4sMnTR2AryidVtQZ2vnVWzOgxb4/Ds1sR/un1pPaM7H8eojFtlkl/t+2oEA
unuOqZ4o6WKkeyWpdOtntIoryiI2fJbsK9l1smyYa8HwEFaxBmJRwOiuEqNAe9vE
vT6JV3qQF/3L1HfTgO3UkgsCReeNFVC6BKUPxftJeSz/pMTPESRDCmzQZB7vSJJC
AA6JoNfFklh9Oi4LlDRdLrRoemvty9xthqabfsOnwQvv79uABLCnMw7LAIFWdUWz
y8SUPX3bxjDDVZXDzrXYRnUpXcODvVTkfvcu8t7u7R7kC4svCR0Uc2f8ywLlJ7Eh
kjL7imNEdNaEKqELfgJor6EbjQu0vJjWixdM116bdoTPOUlH26b1JjPSblzlmm/M
bl/2IkL+eGn4s9y48/E3zop1RtCC0Z4E5flR/AiTBlUF6n4byVOY8aHPNwYkPGmO
x4CfT1fq2eEpWXNiEOdwvS8EZ2xTgJUS9ZrhJ0Qf/btkPhJV/+wVheK54FlGo+Dw
8stc4HL14nrZeb1j7QN9TFhc3DFvfX5gHrnIjUoIRoimeBfJKe0wWwOi063RMAQ3
iF1mWijgnUurWPvFlGBlQJzk0yKB8/hgeNVFDyuIM5vCRWVhz/FKgRIBZYYTjA4x
kPeEmTKZyGAI4GW7wBMvpWKVxH6GfP6Er2A5Fk5DqLb3SfhnReiIJznhPy14qhgD
NVHsRidNXnRu2lb7NiOVTdsoPb3uqbZgrGTe5lFFbiib1aIYaWhlRlGpqc600I3X
SXoPUS+KM9IzA6/hfLYDt9tBaenC/Q2qTt1oZLQ7rNLS97UKCLBpqTTXJuKRimC/
c63KgXGoO+xFel/0WXSrKVi30JEYvLqehDGkJlrQIpgqN1nFnwkMXSZM0UMZ7GI6
AVRjY8z8rSMypBaRN3InysKkFgUsl6T9qJUIYjnx6umPZaSAlnr+L8yMbCB4IfHu
hVbCunU29kZD2nTpIUSQIirrLbl+ktui1YaxzaB/4qGaCrBIzAvrWRsEN+Kd/db9
5xRNpzCHLssQdJhfihpRMWv0LRsq2Q/xLADCH6jKAtemseRRsmm97vhbdcYBFOJX
LR8xfcV487m1LEfWUncBcYfvNX1M0cx7oORpFA7BjquoOmCdyU3tr4CbE2erIRmV
kzq/QMVj6C7Gln1i9a50n/W4fW6UNmjd96kPzqxX/XbmVVSiSa+2yhog7P2ucr5F
UGLoLNNSKbi4K64k6pRxJ6cBaSId47ryU7bWr2+0UPEd3jAgzQMWkxhVXMitBhlt
ZnXHR2Fmckd5sj/mfp6UNx4ZYafrK7kOIaMF/HxJ59CEPS/C5XOayb3gjHJ9VHxI
w/4uGw3G3CUdds6rY+yyfHHQRMQ6OnMBnZanjkVuj0Lut8GFYVSJwmPFcUV3A/MO
YBJi1LDwQZTLobTxW2L+UmNcICUmEd8bigXIbN7UVwrk23pXj1xVZajgqJR2vIJp
nCLi3VCXnk2tJKDxz9qG+Q0HiY6MusOOXQWTXaUOauQfnCnCsKASH0P2m3tzJ3yB
J+wKv08mQGKYWi5fT/qsflaHGrKhgznx0D35JsLD5mJ9ABwH2drZwc9gjFSISMsV
sihd+iYHQ0tlk6vL+Lv1/PjNmdC+Z7OsbIId+q/1RrPFeTMuXcHAV/K4wnYtA1WU
pHvHumbdd+/34IeWmaLiC9vE3wPrDh4g1Up+QHXWVydAW1sUPTo8EIWQGWj3kgTp
UWk50UbP+T9QWqJ16gs83HmMGYRIGuBmV9VzCbXC3mypBpeiDPzD4oGZiOKCuzFC
85dAPVH9hJ+MJny+wJZA84vL5NJRG9OqtZ2FMvzHG/cHFxi7mtKxUqnkmU9X0cVD
qX/1lh36iueC8bWw+Pk1MYXIrvtJEeJ6nuxrE9iuSrJmRtWJfXMsnH2eSUhXcbqo
u3i4NUv4lKnhQQoxUh21PRSna2PvU778xMc4qHiT3+xDZxq+yx7wdcuI1DzRBxcS
mpAyhbDh9pfuVSnn0DegdA1CeoyuYfsXrdH2//MaPkLukDhuBE4UHbYTq7A9QOU9
JQ+F3w8Ivu5gYieI+1h5elVfyYw5cYFuVnVUi3VwbuTCaHtIv7h9BK06S6gAGdhT
HbxU9V6qVoyc9Lj03e8q84NEQv2lDQzsyX2kV9cZdB4EBkAJVYTdRJR75zgNlma/
9eoUa78s0OKIZepvNz8zjqMxyQNB6CqqGuIGsZx0Ps2QBkUp/5y9yQf3ApayLTSA
Di1qvWMZyHz1BysRZwmog4N4u34zUBMuU3FEUi/P1HTuT7AuyreWJJUYPQAFrk3L
9whF5ydE8bjSsdA35+06D4P9fySTlV0C9RnNRLwyNR7ju8Dc/hlqPyPPPL5iVsMq
6mkDfyFSajsTyDzlE8Y6Ixfx0RMQ1Rqma9JXzqpK2dRrZc8fWFA/jpjFSnix+ngA
dSq9vAGGFyCvD9c5Sw+nBa+T8dre+fXLZbo+frKdEbwetlIvh/5KVFwn/Hnb/9Yz
aJiTEOvonYqrwnQkIy5RGCXbfRYIps2CKr+ZtyvkOTQZctYyQdK0fpQhtT4IDEps
AXC5tDLPdeY1xenUVg0PACeDmFREj70psYbm9moMuWCr4zy0w7jMlNmgrIjYVJFo
miZSVFxK/DO054n9U2gO6MQqpySEPLy9S4O0h44c5SI0HBdejSdLusQYa4Z7ScFH
NkF2zoKhDlYOW6W60d7jH4GQaqxFaK51mt8CEMTlCNt/nWOjo+T+SgeZCRLsPF+k
oFWnb+gGw4MN2xZPlLzMsMgMq3M3tnFq7vb+J1VVioTAlSoOPHDQ2nNQ2SCjAymp
JvDvKKZ7BozIRQP78NVpshLxPdCh24TnW0MrII3w55Cz8OzfgROXxCjbv4J8BF/4
rrcWrVz3O0BtpHzgOTYMmFyT8LkarVvNqDKLwosZh2EStRxsbuwh82NjWiQ58jMl
ly6jqRH49STI6StD3QTArfM4KWBaHk5c1M73WYqpf/J7GcTl8qPnXmzxJI6YKG+w
csRQFJ2c/Vrd94Tayzx6MKRQaLEL1RT1hFGQvpXgez17PG2wPM5oCfsCTV2eeiTz
GDCu4wPbkPPaop8vtkNS08dXyy2iTH7jPK1ixYF81CZhtZvhBo2r7lAS2aiDQss1
7y4Ga4AyNyAxc8CwE1ltRIAR1hFdqladTHYKXxlKNOkSVdNB2YsXSt+1JWHmO3cd
2jr0x24NFfi+AV43zbo3taGePpdSjbujyPOPSm5SM0Y2mXBTsb70KLk4zR5+vDsk
fAKgb+MNorGqxy6WeK2cCz0rCnIXcvQhyuXWT5L3Rx9eq6ztHgCXzaCUxsQMnPDk
yCHZfWe1QJuQNmfKK+YQ+IMTqrCTfZxKVpbhK5huQxv+uQXgmRiAFmbX3OT5ZVbn
NWvHCWnzif6XdR9hchOX9S2WLgDcZRW1OCwW0TWuva8dcT0AFxRiJboZDrMZ8BDB
3tj81yWtBtuEZcFtCeUhQ1m9CT8n9qw3qt0pKzcxH2+HCMJnrlVUdyVOCLSkAzJU
3BCz2oEiOB3xyna58Ap/WPSCC9X9dBL2VAmzBUvoILk4BrRq9GMGUKJTdyo5oJ3j
Y7g5NnNA8CkpZ1kmQgVIMlfkhWtxRstk/njwXoZsTU3+TR2yLxZ0x3tw3NLo4Opf
p47EeEipB6JD75YXyhmQzS4DOyTzdH3VLXDQ+kM9epUfu9HJcRHFEvxhFdbA1YPE
zaFNzwruXgtorZyvkErpeAPqzOhU6XPOMz5SEsDJU5kvB7Evk9Kozy6FphRiDnP5
VgtQyNHIFB6IBUrLgCCLEhHDZMYErZbS4+gGSUOUSrHFg0jDB752UtN4tDgOADs0
8nu9EG2QQF3D2i3jNBAXo2/40FPOupbSmDaq+m3nSjlQKB22D6rUNXc5xb/oV9ak
AdeUcfnTCmOAa+MNh5GrfmbVo2PjPJnyf/+O1X/C+nASoC1JLrcYIbTyCy20aaKT
AH2sUtQsNGZypJxFnyn7tvkmXaDDFABhylKJzhJQCAASKJde9RVud0CnPEEC9V5j
h1/0LHB7fZeO+jUeNfVEFDRuny2Zjy+SwZcY0jfG57fis5Li/kuHBUrkQ7v6Vyxy
fyVSQbPTjYdU5b7jg0xYrlhJlpt+tVX2wXAmJwedj7yTDqQhIO9d5a6nhYPbFgdq
UDYKLr5ZAY/OY3KK9cXLkH7NFIRQNZrdrPrsyPHzEtJbW8h3KgV6oOMhWtqpFuE3
IZ1lObnPaPlD8QzF9dNekxduznjTRbJAIq5un4yIl03jLDsK4GlCotT42pDUqwjk
buwjnZ9VbHjvY2XWMtDMIJXmqMEEmypGQYTEQAos2OVXP000Bkr1TzwSmj2Vz2r9
/G2PL/WHarOs91xuxTFhJlzl7vJ9alEobd9UD1YAio5N+luAIDkhY+pWpm+PTv2+
VQ0+AsF8ZQMP3T9Sqd5MOXmI0A4YShVyfyU7+gqd8qHXqH1HKS0Wg2BvgNmaQu8Z
aI3Oq1cqAgRJoS/ysKlYTVg7CYatFj2+Ssv//uuglE9D3pHcBR9q2ZC0aPLqHHVw
o3wCh7hzZvYDS6WE5HQ2yw7Nj9ti7yCSS963WHMFIrMPuJB5SLFNDoU7cesk9Dyh
97inFn1AXoa5m6ulfEwl6fnC7FnC5IRB/d/iEdi0pLZ/NGnIyQtrx25ii7aPG3XD
tDfTWRcSKbcQyYH+T2GzsvtczDgJ1CTS6z8sms1ZVioV74HIhY8e+LJJH2mNcGo8
uhfgCH2ln6e+WqwA+dt6Dr6LLYyOdPVRGsqAJVL5LvAFS35Eq+vr/FNcOtfXkUol
zV9T9xaEOhlg+2GaMi+PcF/ajtYrnWDwzvn00dwGvW9JNLJVGoCq9KJQCzIBu4L9
oRmHpLZN9OGrjd0Oc2WvBxoXJXKDRER86NOiZEeXl3CDgCTUg9iBEYcZhZ6/UEuQ
dWDXBooc06h3AUkSchUkGvcdKOUDD8z/94q0fwSlsPDWdiwElAWrH0htHFYWQryQ
70n27sbOvqeg8AVvOyGUzUXKQ+K/uA08PSv6ukDkfj5cILmT8dpcuPpwdpcVqAkV
Zh2n7GxE0uHuv5SZYVD6Immn0SGzS0AE4vyrzJOqYE5gkiJEKHGrBxefCdf0kcY9
0gPY+DP1QcsWf43MgY8EJvYrPeug2yKaRms1wSocF4sjdo+6OwXevi00AEll/vOj
9n5LteQTeIsCvHBsW3F3fWYZtG5Yt5p9lk7Mk3v6GOwAKe9szn44HLeLM2/IbcK/
R1VpEg6SX5ofnXOLOkkDH+tBrQY7krWTX1Vpy121BOUMDyfrOaz9njU/lHGIg6ny
ri8wJoJWt1YyCHpV69hcMabwM0TbaW7A39hO5EQd1aCkLE0YLI+BXZQflVlRwiHX
XjiqFBH8pLh0UJJa8hKI9z2K0pwwqRetIRjWP7avwKRqXX2OnJCGAEh+zylED4Q3
KjRzQ5RW4vUmgr/ZkzofOwweHFexF3OmQpi0pKeg/cM6ui9VsCjZ8zGJvnNXAo1g
en48LkGOekC04aEeidOtJ9kFtYQjtqsT/s1vndax1QZa8KuhPcvRkv7u6IKMXU0J
3yajDSlOAZ/srM47BmG2rqgAZsifglAqUff/mXAqW1Iv/nvGb3D+d8rbjywYcEl2
FR3OQ2fEKbQtxPo+SAnUFxv0BjeKEIcZkSm31Q71veubd+9U1J3CkXd2NQmhzlWG
CXotH9C8ccn7beNEzA49K+tH20OF7LwHm/U4IPrgDtRDVpPiU/TZo8vVBR5hP2kj
GuIbj8LluiUZc/DeSeLr/SDhV9fz3PAzHXRs6YN2JUMYzxc6zezgWVNFQ6bogwLe
tHiPSztxF1Lef5T4hwb6Mplp8PBZh/inQKDrbTEviFIJAu38uq1w2nLmDqPK52X1
/HxSAFRNjM230tE8Ba+BJhAdYZnr4Z1Be+TVXnDvqvbOdUnrvT9JFoVG0cBkHN6H
RFdKdTLmNmTqwgTC4d3YMAZIAWaB1icJiarwhSGcUsZaLK71wY3ZFS+FRdzPjbwp
LkzjrN+HXXFFG7I23Y8G2kAVymmifNCr7XTJN/HYIh7A9H3pZtOaCH+GEPF3gSEA
b5174Bgr/QAqSr/nV8nBvEevDkv6P0osPbkp8r5G68gPrna6CaoZDCesvXQY11u7
TLi1elOSyI+8TRFdcoHh0QLBXSS6DaSRFQf1vjGZDkDMZu/i0QLd5dpg9bR3kQnq
8frz62XQ4XDL6ztJPq2z+D0dUZ5DQ30lWth9zWtOuhagi4j0uwrir2dY9bXzBRsN
OwiWWxKSFO5xZ6JQVFIkOjhy+QdkAoCyZVhvFz96gs7HubtKGBsC27JLcjf6+HtA
dlZiG+Ub+tw7rHu8YdaSgAsX8lfo/EitpsZDLsO2sArQObzZus4aYoxcrPU/Wwck
oQAJ29Ebsd8RARR8dovYfXxBLaDCA//hxt5/5ebdYV6pSepnQEy8ULINzOMTZDSn
eN12/de+6r00OYJYoHqRO3sxKfd10dNCMyiir/3I4b0eERAM6OVp7EpS2ZaWbMs9
ErK05H1Tfk6awgILaxNafIGlcsY6R6KIcGfJtltsqgVgrGQebKfoT1vdK1MRIYZh
HVAMChfwLJkuE0I3jlWKNvOlg8UESJEt8MmNMSqlAGdaJcGngzqxYtiYSqP5WXj+
mQ2LZitj/Tt5W4G4B3agLoTPluR3rKiOGSyoEvDBkewctUQFNxM391J913ReCRUk
bVdAbutJOpJmdwwtHfDr8DHbachA01FHdF+H0pL2OXs0ftN7jlscfihUaUuC4acW
pwQDJqxsV203t6vDnq3ma2k81MXt/cx+Dd7kW1F3G5ODbjXp82l+l25FjTotQLez
P8oOOf67syPlvFNOKKDKdDvqQsdN31nf6I5DynMy2wFeGX6jkQ/x5klW2DkdNQco
4YWUjN6IDSwlonVaMXQYw/2dpTA/YmYjYfIpozNk5YJCJx1Sv1NZBZP+lb3U5mgt
BctmVOi6vd0rxmrpOaK17O4/gHRqYAoEx81iNmnwbcJajn+wfvJsWshNKsai0jCN
VaeeccsuYkDoNuCKrdbQ7ubehKV9cbFlP0f2s6GlwZGUrInXPnlpkUYLQGHzWKcH
sSbHGEi1LkmX0SVTGIT0A3pkqoeoT/N2x+ofqH9NX4QKsmN3QVrUDCA/QVM5GAhl
beaAfvXDqQdo+YN/cLtErny2J8FVF9tD0SOycA3u34PEfo4tH5Il4E2VoImrEgS0
f5f7kkcTzZD1WGacCuQa7LU6imGKTXwfJD9LZx+ZgpvIuT/ZHw+nLPh58Jbg5frw
6Z2QffA/wVtBC/rT+zR3HPk4Si5T+KOMn2AWHJ8cCdf85aa3xSDPHr0VUs/62ctG
g7SxP/mQzekhaYYVaDWnHU2EHnkKZzjB/nexSEMx6iAXFJYPpCrA7mQqQpCJ/RQT
ntqpi4recvmGp0K7h9/T73Bs2EEj5nvl7CoDBI4nVKUwIfUAKyXKa7Guzgi+fu4w
xL3PAKK3k0z34NK5bEppUZwx82jKfpV59e/wr81ydBMap3mDTd1h9Eu4+OsnozTZ
yYffxJE7ODz1z/pofCUWRfD9WGulVidna0J7kWzewgBy1fVnQ/h0on5MQDREEEl1
skg7lSn5KunSYLgVCP4JzVYhkTNlv4iYb8k//Xuj6pF0gncLjHyU9539wQefCeHC
ykpBKNccZuJnI6dW4bZo0Hp7HgDq6KrkW61O54V0RfcqLBsYhBUWorvmXICHTizB
nqr4Qd6QTxhhnFJZESb20wBzNzDVhYrUfFTKQPK7dVJQp3KiemXsEaDGGsSjspb8
XCzZPAlLzr0yKBdK3+57iERRf/R4Zc+jIx7spASDthxZD4A2PsTNGUvGXVidW1N4
Vcf4l47Z3oyUcj4lB14Wnu7Z9AEsgUW6cjdLqLAjXvG7udUwlnfONjKsIom6Ci9R
f75JjMIzmJDSFcFuwehX0oRSR4JKEq7ir0xH9qBatyuGh6ShioVRkK4xBC1wXmRM
mRkMrMdHHyB+1FePBeZiAyZMTzOV/J6SV1oSHIzASr8rqC8i/fcuYIYM571FHYgV
zEYAzjHb9/XhzAF3tPEoOJgnvI+KNCxY2tTiNtZeAJFUUGeDBvr3VZJZq80MzlMv
LaqsXn5o2wUM0njKN88zeR1SIp9YPb1s1V0NFwBSs+aSYIF80IID4uwNxovoE/2N
KVfdTdOoRtUEfuER4fuDuls57e3VXhghW+vv2aixtHhk+trenb1PzNi8b7ckaAB5
reMH/5rZNuQd/wpv14R1+tILiTTLhbf0/M42GS66siia+Qc5JbkKxnkmAC+elyA5
yCxBRfwtv+ciGZyZ+0sB+3awNT6AndfibzG0JGKdFPCQ3vSbCI3hy+SKDW43JFzs
ARbU3MU9Cjqz97bcDTpZdsdsIKq9XU1KUMo0w1wn2SQ61ESWV8cN0VBhZa4NMTX5
W+CUnclcs9Z+w4yxC8TkO5evDxYZVorgl7uhJUNGwVAPGqyH1zXjPDl9+hG7D2Va
/fz3LO566EWgGRAwrIIohT0IPFT8XjqnypPGCLHt3pCmIZ2ImVIcv4adyHPIsxOM
YmH/xXdqdqb0DfRvBw0SWIR1NHgdM/0VbbzWrazy4lyt21ltTliJ9PQpzLpB7Q7G
166x9UIHBZT8tBDVtJqO57/8ZXxDn4fF3jGkMhxRLVMUQgNvRuZA9z4LXY6U56eJ
b+pcupWFZncEmG3SK0haPnM82k+oaLspO3zUCNQT5FhpqdJXBzbqci+n+MtFNOHu
FeD/xqs/Sg/tyV8n/ek6HGJmdwR8Ci8utW9wdrkFRA4nTt3VdAsR2oIDXfE0jKfT
fMifhZicoR4Nldbmdn1F+faphPAwBdBxt4qm0Mwns5/J6+HbOPIIIc5ngSGbiA1L
ix1HeFxrI9+FrbMcP1yx86KZpQAbdtvo5pVIQ4uvCYYuhu+8J88S8zMk3NLjjKDd
QvlXd7xGswljB4b4d36KcR0VfB88YWOo7MWfwoqph4wb1aJN6rwDBRgHcfdjN6k7
lFS/T1DtuRLymLJk2IA5rIy7VUOYT0d435ZhkTH/cEcmxgNpkLN90k1qrdDs7JNC
HpK90uNa0U+ycIgD5bWWhWYKntrDvUUFQ924zudhwddv/2KB9JOOFAjk7XmjHaG3
z5RofNy0uQOgXHIEJXPyZAHxg5co6Kmu326Z4Q69DDHDolUdcRo6HXBEpqAUeZvu
COB7swYaeTZBxCTQPYUXBe8kRSVYWoJqgduMMVck9oyVcDFOdRYsImGIJ00CKWkP
T5xgJNCmaBCG8L4vwsriYYwscvSr60UMKsXaCR+s1xP4eeTJ3JCVgjsM6ZPe/3KM
CL/wNJS5ydfJPF8gnqcpxD2FB1Bcn78c8JR63+DxoQUHH8dapPaw4SXgyvaowtYK
e9ZPMN6CjIHQFxG2C/rcaninjZwrdFBWFH4CQeTeHj+N0zVk9avfL5mhtF30lwmV
kex4Kapt519RdpmDXlqdejlQRW7/y198tpMbvUFb5LU5CxBxzZlB+rdPufBJ42m1
xrb3TGRwwIb8tCQCN2hFSKxYUO/vBMvKio95483NuKTUvapiY0oO2LbqveM4+k65
Cvhe36PRbAgBVM5HMGlzWYKxNKqEwiDGY/B31H3oxUIhzJ1yjRQz0W9YrxrFuvh1
uBgbtvHvColZkKXSrQ8iYy9/UPUJxYcRE0MziH68S5Rz8Y1VLk3Wcu3DHszlOQIO
bwnR3XdyChjmADGlVzKJP90hmsW89lmsjB1sb1lpxOz/nReSjJswn7URKIfnEqkJ
5mcTF1Km6vj1uf/4FoGsjCDNAHc2J0n29Ev5CVujJeq2rqntuUJIMI/pqTPKxQr0
Bv+o+mtkU12GHslN66fQmreCJ9m4KExjPJFW/yec047XI9R7SpWCTD+5NvEvubSM
uy0BJ+CSX3M5n35nZvyszILRvr+BDDQqk0mtZoOGFK7go3QSYEtNbLgmeZ+PBlI0
P9pKZisRSavbcfLA9Tk51hI473VcEnY41wd/oTqrSeU9n/aQ86feYtzjM3s0uXio
nbUaeKu6lyT/vJaXQtePgscU9ZtyUoQdIzCeGeYT2/WzK7p8iA5yoWNA5UsnI3a9
rnFuOE0d/uMiVJ8zzkZlky2GMrpcvG5eRplFa1DhD4OcIUAHHNYK/qF3pshcIL4I
Bjt25yYWl0i17Z2hgP5NiBqjPlkujyD0Nzd8WbBUlKnjGA4XQQBXs375JxRNkCpq
t1/TEecwtOta7WWnTbTibVJblGvQw0h/2qAmMaBnvr2uyF+xB0jHEZIHaXGKDPyp
hQkc8ZLiXhsX5vwANWb7ttL7z/IE1Ay2cWVjPJoWW8xZCwIGu/ng8cYOpq++6q57
vwQsfwbh4eAWh5so2f4cVeK5t2QtvkD5xTZuI5dUNH2RSrN9255eVtaKiVnYBZzj
4z4Fef4ScPBue7jGvIG/0H7qP/JS7b7QPCktaFKw9flXNve2+musYSR3i6L2zwLy
wXM4gVfT+nrgPUJCdJ/ahAX4duALcyjADl2+miGL3c6MGc+9IARrsDsmXt+B5/8G
CTObAhBEsLpfylVg0AvD99cmSWR6rpcJnrKZqkg0k8nFeiCHi1aRzOJNBGcPCYTw
ReHZYr9pQdFOffONdhTwB79SMFczw8smOLq33OMPM/Z6s63XYdLnbWj4G1Fg3Zso
+Qg+n70LgENf5qAEdSFqsbp/dgzqC52Pw6r0ZEH9+EgVaC56SuReAaf3DpPYqmgz
sYtjSdFZNKy/ftJt4dRaku+FA8sFiBtefDHO6oijgLkef7axbwCPXfOYcRDC89xh
leE9/sqIE7ttZym6NFVg5SMowBwckrXXBHgrWlhYo661duwuPJCI2JoSccnfBmIU
nit+gd3nXWtKQPOANQDbPxLVMBZ+GDgUendnGmAx6mmi+0qEaCHyLiuQxa0EjuR8
n01kTIftJKaLSBnGOjsG67i9IC1rWuH3HVuBnnRmYkQs0lcoeBXvtLlaV+dxHMQ2
L5Fx7dFoyZkyWSFm1BjY0S101tO7ub6qcpflsrN7BrqtdFRVpwuizSJEKebemNrT
qSKL05Ea0ekRokdhSapSehR5djY/HtJEodFAe1WbTN3erXPmWo8DYo0ebzVHtPcU
C14wyZATPIbKs/TQv9Q4Gd4Os8iBLphm5G+xlC3hxBtpVrKo5H33UJiNkz0L0eKn
whXfxE0bdXcS1fWIIkUpKmUxD8u1TOD8FO43q2wkIj4vWbxj5eOfC1S4UM/r4gtS
Ag9iG4kJIbBgvGRzoU/ejlpIDGHrOnEl7PpdYfvlJ1a8N3hBl5rbYDjVV9PcNIyl
W+Y/uOJdIyfITni0oB2KjQSY7NEqDffVUAAd2ijRd0S1kdMrJs/C52dM6dG/N92U
NiYfWu4pfSEymvFjuENSVUu3tZKWt2giaOLaEKLn4x2QAitwX38pieJj43wa8S0b
XAC1uMadLe8bmrl3G6/Y7cPDURA7lsRW4kxTKUvxoFWZX6zdn+ozivp33rh51uZH
mJcAzK40mB+UugRSSlel+sqYhxmokuBdNVgD5s3JoxCG4f/3QPQZIRBkA6uZB0g4
A9GaBxfrP9m+S5fSNmrkDOXYHo5xmGtdqk9Z6MuxSq/k87AeiJovqJWcpb630Gzu
2GGXNkB+oAv2etGLJHmO+8+1vbxKMUXbdMVJ8XAZcoV5aox0TQ8Sgy/mpeWd6NgK
oaxUGjsljObsl05fjiBesZbAorYRK4gUReVrM++eMp7hF5RuD6LQZilbbpNT/zgt
t0msuDGhedJNGh28JXPMs+CsNpk0md1QX/KLvLpFBAFU0gBesml6Sg1O9qYpJc+z
gc7tm+HNk4lYA7Oiizow6w==
`protect END_PROTECTED
