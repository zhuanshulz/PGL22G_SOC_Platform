`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNvhqf+I54IMctEop7Jmk4P8OH2vMV1GUrnYGz2rh8WhgrZcaeahPybaMlR75iLP
n75y+iYwYCp0BNfjkHNOk8F9tph7sMJJO99gD1XAxmyLyKie7JpCdzgmO5YY53wB
U8tJaYUWIzTQA+rOWHuBJi0OzJ65DExiTta99Zcu9gAPlHsaL2jQ6F3+DgAnEP0P
nKjvHaFFhw2k+l6piDS4FLpkA3OdaJhAkpnWr2/o0f4m2TrY9GXsg9BSpccvkMIJ
WcCVCEdj/QE1FXZP4z3PajImctGaPnEYtTvk+kE4VyedbBxE0jsAMch3Kxf2RS4c
Kb2S0sHX80NQ2RdwoYAgcysdSEQVCOd1dyK/fO2gD9SU4i53MxQWkdh9jdY46TcE
u/5VVrNd5wVHm20WZhHbqbT+tM2E6oqal5nsV947jevzbBXtU7gPKGHeO+YBvT49
e1mXEP+u7r7a/8A7p/hBY4sAspojl70+o73cSWvMzYhHIBwOYVBt/ysOM8yIPkT0
Kxocga8+d/VULg28hNKUDcZxPmOI938IwpozAx1mmBM+FleRZ4xKDu4dymNMFrrT
0e+PlmTVQqBr055Zphp+qbMfw4stZK3WJhv+OrsNaUazp3Ai8fAYcPvOOBAibTxG
ISuSvWJFxYFzE66yaHNkngRdYAlm6vPWBh9RacDyeHVXyIY48Nv6ERszYWDpvrIW
x3zbnq+Q1wgY1yM60jxrHr++uyjMvC74VSVcplqWdzk=
`protect END_PROTECTED
