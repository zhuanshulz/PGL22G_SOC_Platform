`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnmX7Kufru8wT8y1hNWq/931hl24ZHq/wMP5s9M83UcqjgiHrmDAqN2rnkG778XG
kvsnbPrtMwKTlnjX4WAye5rs7W6VZc2NrkgA6JhZvghLfDEWZTYv0Y7spY9QdW6s
9poM8TMTvT1zJAYQ8kWy5PyzUhGQl3G3bEabDgn/H/FSSineEt/01w1lP2e4qz01
grhtq+mklTtpXfAkxq+5YCG0lTzFZXjtOl9FgmbXYsptzoVV0BqT+tEr2cKQlmkK
giu6hF2GXXoE9DzO0U4VJ6XCkik7o/0ZTN5n45rEwLWFJilGm6QYEtAuX7byBjBr
YN43wrTwaEFM40rMzf2CwexP87orxCqtZ0c5Rg8Z7mXIfxccoxU7u5+p1k1aJ3PN
OPNtt+WjVeIyVbZoHYnc1gdNOORFwnbMRKo+o6EJ5knmbxkhBKve9tfJ5RT24cHR
rtKEOSwBKk30vSi+kF3q72UP2esMoCeowvXutt6izf8BtUYrBjU64/MWVlVBON+M
dM8FWiJgtv+RqaPh0GWZOt7SUjrsC0KrtrcflrprS1hjMBHLupOGAUp6FfzCsQ8d
Xp9QTW21806aCzyRKcfLuvPYrUQlRwJ3U5Shsngisvzp3QOdLFHpjriLbwjF1VRh
tpeFHOIqsTOBhi5mwkMU0R1xEVm4Nv3P8EzbVHSW0+FOZqZCuTYtMAETYktSKhm2
SvPKQktInY08jLgh4egRSB0pqR7BP/C/0iEOSoJBkLdoQ9L/mRCTGzNvlNwozu8o
3Zd7tdZWHnrKmRgCcO5VcuTgA9CVf3GyZNyGZTxeb5NOKXj9dV6oYTSNyTSyhhSO
Ef7v0Rqu0K8jOtiD4XCJWki8RkfHvtHxKrhLA4cqTXKa6NqFez+hQpcPLuS5DOJh
P1JOE68fzo3zFIJ6lWu4ww==
`protect END_PROTECTED
