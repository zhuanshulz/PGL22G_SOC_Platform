`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EEABq16kYCfNoeiSx8x3a1fqWToPVG7CDNld2W1cSCdH9zjQpY5mxbogp29KWAli
g6FqIV/BKUQnA5+ddPV1ut1+UEisW0/hrI4mYLOEe0IvVhttD7D8gZsX0m71raCd
RHTxP6UrpETlosOHn8bGB03tEr312p+Wm83ma2McSvPekUbO2jY2FDtRvw6hCiNn
UGPS7Myof2hhXdgDqqE/PEwI3IlxxJTU2FivuxHgA3CPluDJD1g9/3qWS7fer01q
2+w+ElmxBahMyGxh5/ogvQYxxkV6HXfLQyoN6LDFtc+Q+PS1k0q6IbZrwAqjYeZ4
hTiRFRlgSKHduqJBVENCDhgwjWaCNjqUfUgbxoGIxSzkSq8roCJRtTbIT1jd3dB7
yNBxr2PeXmPKJbuNCs32FyfZ0bTlKZ8Zbhl41YW2zhjpaQ//XBFQP1UI6M/rAd3I
FpjvCk3c86gB2ng82CdZqsWFncdBVrNhwLPWvG47ardoz0JAenw0qxYV5/p7pdFM
OP4/V9rUSPDkbdIi6Xd1DEjFCjnINt16lgs9hJYKj2ktzeUyU0GAbwOX3Oc2U0ZX
mZkc7UaXrnUu/eg+OGQLPUOCOnjuLEupkY8Oz3mMzvaU1c/ku4wm3LzkgxyS3E2P
osqB7M74hkdpgYu/H2dhKUJctGFCfvjMKDRRuDzbBbu+Sj943o5g7fNRS73Pcn8m
T3zEEiib/zCF/rIZzxiHse3wIhO4Axu0dx2lgmtJkjxzfWw5Wf8OJDBOrbFzRX9A
hwtPPAVOcgJmiU3y/LdYfDgG1WcN9vLkzt45XRL/k3x0HN0sI1ge+Cqtmrv2EzcT
9mfo7jz6oSja5fY9ASQsdr87H7SljKSIPFv+9WLjhARDCMCpZ/MdJ8Qvm5gMMhl9
yNY7M+iSxc4Ksh7K+Zo9VQOvIqTm+dG0RWSFLnBhHIMAt8LZ95BSq+tG/DjGps+0
EU0XCFUdUcc94l/EuvVBX7dm91+I2FF1H0ryPb44F/CkjM3AATYngCcmDLgnk5f9
9FPZW7KCza5vBBBUAFs3YHRLZl5MisOYbABfgoQm3x5iF+6z6wfvR+DGqIfsdNJ/
UMFEuJdWh+yVAqja/rEjNBM/Gid61MX/nbib5ZhO0BRepY47fR1LsRGdXYBqQP5+
lCfUQgSCB2o5vwwGglsTiIpEbnPhTfmlH/yioa5eYEUaNvDcH4w/Ss5s6/E3V8Iw
jl90KmwXlKTqW97CZef5HS97CuwLXzoQSM6IVSaRyMLy1Rv0Lq8cKbv6IZkxCNEc
8Jn2n0izy25IRhW/YXpqaaIQiwbXZdTyO5rMeYUN/JdelZsbw5abesdd5MJZQ82Z
pUJa/72Wsgqq5xK7lrPDP360gpVgdyW/2Idh8/FZGaCkbqLt4c62BlS7aV6S5VaR
5kV8qgKtXdeDCrW7UWlr32IF6BJ1R4wuH1z52WyQkpFTeSHoE49Sg2W73k/9WjX7
B/uscRMC1KKkFO6Zx5ZR6jWIs7pRZtMCLx+bXyyWVSE3KkaNv6/Q6JftyS27ZTIQ
DZcUaf7CFLB4lFv+5kHM9aPrV8fMKSFPFGAzHS1oOj7L5ANFcXD+m43PkTIAxFPK
EQp7B97TEOEFseH7VUmUZ5Q5ZtnRINpXPRkqEf0rZFBCXKxXSFvTlEtqq4LmLgS2
G51KfOfNencFt3+3Fcnm5yAImEhVqfcKNdCvrjv4HU0GHW52/EOFKSr9zP3HwPWu
vPwxXiL1OH8S+FFBAZ9A8ufXAj1qP9gP8CF0p0S33kQ4kzaMxzoLs7mWiqr3UKOB
SDOAR8xA+iAdikt0EJdZOvlDdxaTzSuoxfMd5jlchg96Kkjk8yJ1EO/e/6q40CH3
mTTMfnTwJx0+cvHh7cDv8iLg0HBAKSXIEKyBTDJ6uuPjxB9c8Dt9n2sx1tgyEK1j
I8tDFvTA5Aoe0k1wcAo5PK36zTIfO5GS7uho2syFd7NwqlyCFfxLGXnf6mu30Id1
WXhXGf6ibORQsIFr6MzzcuFsG6o4yisVzijTv7gBSd/Mwuo4OYDIK84gtuavEmGI
wMWAQOwnjjmBGLYY1PbfJ5Q8QsLuOUBeGZNVUV61wXPMW1BS21Ikiw4xwAHySwdv
bzcvi6MBVhZnE8hB+14TFdZW1f3WGkisPTojoO5BA0GE/4CxqXndizJKupoGDDU8
etWZ2lXob8xlhiIIt47ObEfDphgueWoi0Aem9LuZqvsHbc9Z9HJZFD2lXY4Z1IgW
QVrq7QaEN1JvoW9aDjRutzucdEn3ON3dO2LGC2nfZPtaspg7CJSJrErK6I6B1lKV
O5R7PlaTgTUUJPUrQO0EuevuSF95Qq66msAvxk1++KAyIbDGtrc7P5hkzrPMDSHC
gtdQw+Gu8IzY1JiEFUfWse1hR4zCwNY91tOnXn7ssnRC0cnElElx1vzr2W4OeTdR
m9x38nPe+vryg9k8HixvihUe/LWg/U3+/QAbySnIGNY9FOfh0ElS1vzV2FKKb3sb
ZmkC0qP64mHisEyV2fGWR1UIRetVGwz2v62nkJ764YfAAgziyrIKPW/zytWbFVVW
YmLAogfRnu0hhVpTLwzoO6eqg21yfv38ZQriiYrwB3xVQzlGJTFxe6WkHx+L16au
OvrhlypfcyMlf1UtfsPTxw8LrIuaNu4Jbtj9ROjUTUmQb27ewjwz4G+SKGeLkecp
RQ0sBlVE59JhGfkNXw91WbPGHsfZRrwCa5Z7VBNKVppnTHpw7Tn81O2UZi2eM54O
GaWifFUZ44H5s/0bsc4gji3U6P4IPE4wu9CSDWggLqS3fXtoxXXu5I/sTxqYFhAf
hXG9k2lRvcU2buI7L5IEvs69P7dscKuizs2sHRXKM7xIJ75QdM8Q7hujcoiYw7ad
NihGYCyPGv4iC4sPvHDA68AkZdSSCLotihPEBqZsA3fgLBHQSSORMQ/OxEQbym3v
dEwz0f+pVbaDwbqWQz4KcjML7VVmSMdxxWbvTWp+2dhHaE5nHnQtTrpRgTFNWMf+
iFr84E5vHDCaxVeBm18X6a11rM58+XvwoZ4WGZEFxENGO+I6CqmF3eo3Mpk1nIgK
4HhzjTf0k5uxMSAjOwJAi+ub40XRDTch6LoivoOJqtynjAmZTTYnRQcnoldkSZEV
fz+kc91R9vsn4bMCZy4Ez+6M+t4Cm6jwKZOO0UhQAHmaMvFwtM1NOXI0W3dEm+oN
b0MtZ6XYywyTa8KtgNFZoO2T/gNjwNAlR6Q1RuaQ4Dm/rh9gPWg7kXwfP3XsW+mw
rq+Ky2OrtIvPCn6yFwHs+gBsU5kJ9celQw7VMuEokFfJ4DHY7wvallA66hEBiy7L
3/C/trVUeN0zvHMAOiYCe9fH04kabvusV6w5KiKixnzJWr0oG5LlW+bgnn6BzQWE
MoiUNt+dNVd0jXkNEGUKFh1lqovU7+rBmpzAC1Jr3IzLyTKM+8O8gvz64smDH1iK
+hkxsH2CbtESEWEy8gZIRY/tpPgk9Cv8nB7Gba1qTpSlnsWOZxcCE49BA6FaVfLD
lm+3Jpxx3e2gPVkWSQgsHncEB2nNtHldqelYTWpasndfoCLE/LM7+zjeKmzvC50R
AmIs0fGOFtoSNJYM3JAbHYPLjOvVbeWVamRZZqUDln+HQ0k4rjetrDsCSSEcTV6Q
IaEr262S0BHR4R65KKZT49+hTKPSRAatqB3jSuYwbEFV24+8BMayivYs67GGG+2o
Wf4a0kCJZTAOf+I7Z61QyjyElpQc/2kI1Od3qKbOdwyRMLNGb2rtY1bODpeU8VQ1
wS9BpfMlKJvBpI+0rJ0anlYBsYjJ2ycJ2uWtY96q8vuJpemKnsL+dBkd62fabGXI
SOsEmvZF3l2rj1utXzrTN4RU0PGy0FzJWFvn6ONMEPoffome8NORLdj9tQyBuiyW
OHRTqP7Mh4HR0FiRArXQBdTSzngmmS8+DoIgNo+dfcbtZ92QgboPbx7/i6WRIql/
POsTKKq3rGNHYXTpRbJVsYzb4yn231ZBvKN0euy/hfyPnYTH4P3WmBNvbPLINFDv
SS71OpQILPGzgukj2l3ubE4as+GFbOk6KT/K2dVCSsYTYhYRSyJIqws1Gbt4cTzw
ZNdM27pHo4Sm24DCfVMp+IOmgYXOIHDk7/INtttrCBngQ4MOck+FAYn+Md1W1ASw
j5ayMuXfB8YvFxNILBHd1p165mYFDONGKxME4D3uQB9LecI+rh0a0SYWuwJnPbli
aCT/joUKNVhkrbz2Xqi5RSVDnijiag63doYZax39/MbwtxZvQ7UnlKMM0UQlk2iN
tBDIBFGuYEMJ9crz/qy5VesqOW2/CAGRZhgx7cFcwtlWb7z6M5RsdYViPyY5Ccvq
LUC/B80mX3FI9fCJ6b8wVPkEGthc5YFKQJxj/O3l+Zl49oSL9EHJ0e2AL8pZnEXS
TWppcBuYC2VH7NwT8IASqooU9ZulWRvct1FjFEhhlAcQLnzenUVPMRlNz348U3zW
z6KZnFZrqsU8gyVEL3lUPuU4Zi91I7k+SWA8Hkc54Fnb0r+/ChZufvZWN8nlTWm7
Z3z8YlkRQqfPMxbAfyxMK9Qc/2C+0yp6mzLVy+0sxTZ8RhKsV/H6nlkw9dGIKSJG
ZAbBQglU0igwSPdYGJykZP+ztH0EW3YIE84tNdvp/hLlqsZ1IPSgxvaw41Osk4cO
0OIKGEH9v1Ml9uUxw/mphTXawFoyvq7oELvs/xfxWpFwVJpIJ74QuoXprjD2InFX
qmQIwJasWT/ikgqA09OxBLgnkpEPUIqbORGML6h96Ft4dqAcZAFhnC7W4i2Ysynb
RqPSkAFsNeVR9hi0iIAYJ9hDLc5R71dIIq/1bINCWZN17tOCjDhFJSWu5YUT6N35
8sRK92EajCrb97LEODhcqDVA36/ansjWhBpxvlg/9Fcv8tknmOA5sa9oqRKkmvif
DKTHgS/CaoY7oru7mFocECnExWyDcC4+Xhj+sq2x/RoeuG477OgTEED8tixmcx94
GzaXLW04DMVVvgs+a7rXic3AfqVt+v5fIWkGdkAHNjhm/Q89FFTJjpjtei/MDOBm
oCMVs0xTN5z/+8f8sEio69zyrCkZ9C3YB6jD8usm5f9UwQ0K+zVlsPlMviYTjjuT
Xk1vLzVKr6m507vqZ4od0+StuO5jend5bHjmE5CbT11d23ZX6WopCrIsAvTn2oTU
wDiQqrEO77A+tIPTGeM3xASCyFr/AxxPHj4We4YPkX7V7/rIVueQhmuJwzKTns8a
yfAGx0OOnMFWZAR8CP530YoPLEaaw7Bk5h0rrGONTBEH6Fyjf7i24n7DhWq+DVqV
+J5gmsi6HWZbk0JrWw1FjYORd5AXn7xHR6dEW1FpnW2zleYJfSU77dfACupumRDw
C98oa25EQRay5/7xEziFRZpbq7/7AE2Oajo1E3YNPdhAfBG58+Y6frXidcYTbcEd
lIQ8GwfjYudA+XYm/NvLhGPrGta3i/XDr0sSYotmdfdx6MthEjBmQyHvztwq5wkl
2Yh5nUtG4NL6XMCu0JqNiULy+U80KhraF4ojqlLUMkC+kMwg/0hQRek4X8yIMq0n
fLt0WlItD0IZp+B7PoKbH23QszD8yk7lbmMcGtXCFYEK0dEPnaGFacAyj3L62CDU
lLEkeNEQ23fG6ymt+vuJwqXn56DAxfOC4nHS74wiO0GdMq+Z8LbqT70I1lV+j06g
XERL8IHe1WHPo2MuxH9ffk4KIxQpxX1aSObxtxgnZErfsF3IP9Lb+gNSOl6FNqhe
BtPx9lH/PExoenbz95oU7WcGaiFuuWL970KJBcdTp+207gO1vs6XOUe4BQBfaDb3
WAfhDTGUm0rxQa5GrNzCZCLGAi4Luw23gkXlE0cL7BRI0UPenawqqwq8cN9AsElu
lhVbBg8YxJka4wh1O3FkuPkJd/3kxBRR8eJMgfEYfs3fgopPH1fpK9zjpj/1lmvG
gEM7iuar3MyEsYL+eblJu8vQnbgj/ixVnwZM5ZVowHEWYxgKW6ddA0Jicsk0+qYc
t6k2Ne0XzqKeUC64PgqfR9EE0DoGm85dg0YklNYucfXdsS+7ZHBdVtgjD5z0etVx
GFKVSvU10TX+vvUkRyj7jxZhRZht/47OSDuzr3j4sRBnfQOcSxTxB7fJYZrT64K8
Y6PCUZ5wJUyXcYmeVv9d6pb8MUuZ8EirtJxWAAxYIkr6W2whFSxc8cuNLtdMiLua
X2JaXMXPh/IpvS07X/bW2bV0dRS835RMfZvGYVr7bVX6CKGTtzVYkF0RjTUoQoP6
gAgEjvd64hvYSNRfAPIU7pi83A0f5OkRM+FHSG9wiafOdagoWmi2vUdREvqgxsgX
lQVZ9EJWfQnlWlaYIO8gjjUd1Z0RbBcaWruL5CChc1D57AaO1y8wwB8rtij+tY/y
Bj+bLLIvr1KGuAfUBUWWmKNG+Kcx6pGFZIaWF681DDq0i38uFTxwR3f+f9ZnFKsk
u8iVnDU167BMeeULekKlwrNfk1XjWnRsmz+GnH+ZuI9LPG969g9uBTIBGFGuLTsr
a+HuQ4Au6bEq222zPkYR81M7Jdu4jLVh7vKFWGDgpXJ/EIfwhpoxhcG5PYzzsa42
IFnxqmnUHgZ4/RFUh7RKqvkpCCgGNFlXmla5HC8q1BQe47H8egFM8EAqPZtHgMMV
RFTPyAK7Zy/+Re1382wxoVjRQLIXDCfEhXrpokYJf9ntp9T6N0DZ0pUM9l4dJuKy
/8/UsxJq6F452iFbDKv+8u9noZlVxRt4wbhDoCd6TffkjU/zEr+9xPLIYrXeOdFE
pzEjyDZ+mNJJemGfgSELquE1cH026k1znXURAA0zayTu+X4egdznD/6UIixahR6C
3ZBKdVt48yBERdSoqzKFHYSfktcjsksEj1bwEi9inawn2AJ8dmd0O2pTc7hbV/vC
2OfltTrHKQMDs6cG7rhdcWzaH1oFhD8+RyuQ+yLpNccTnAtGv5StDyS9pw+g8M72
qfHoqVR3YxSp8BjiZqB/2dmYJoNU4a7haYp2B4oTyC25m3QjqvH5kDlo2WRB72L7
U63/izsFpevQxWuK9crhmHcMFdjBh/ihUg9Xcr/GqJLbAWClTUAwZu18DAngHTzZ
QdSr26kBJFJ5xld18vzmz4rtdVo4hOp4MsaBeDokfhosQw2QJrfHpU4dqb2h/0Tl
AEXR5Q5A3uPdmLNSXkig+VyHFK5ddBXEIbHMBKvm8kope9z2RdLFN5u+cYIr0Nov
pqz/HO8zZ7sqLfxvGDLCTFAdZ2ztO2YrdJN1VinPc/A5rHUGOnAtxvu7IJa1e22Y
3m0vYbG48TpVUgo3o3fuibfxyIF+DQKC+dkLW9tw/m7XJvsaCE58J4z+IF+IqoJn
Rflap9nuC9CFJqIe9NC3uj+/8OIfb4NJe8546pdCNqI4qxJda999z6SlQf4IP0Zg
226pfbNFZoN1NYmwH4tqQMgBzzy63hchixYhbqnwrBKiGKrplJSPIn6pylIjK5bG
RJ2yf+MtY8z0LzHAZ9USUV9aI3RGSMEJhSZo/BIsnFH0DZ+JYRexcYP/DUnUm9PM
Aa8G6/QcPFHU2u8FhET315nwHCFZoLrW2ihimThfxTXyFwbns9QpbIh959zSqNm6
5sh7hGLxAuHQW9DKfv3AMxYsXq7fpOEM5Vz/ysciqIDSwdwSinEHo6k42hVmJtCF
LN4jyMLEWJF35Mz7+TFrSJqFVOCsyMEu9eKSqLwcTuCmHFkGC9XQbe1+s/AM0V2J
RokpGh6rteMSmSVsfARf4qkBlh0Fj0Xz+dUi7A02jGY7p//kfCRW9KQEZBRFjNX1
vlux+xBuTfjlUgo6rhMcT+mVdzGPVJLyCBqCvBqUN83P+iQpYxYw/PftJpuCMEW/
I9ha62MlKVBD5YuSG+ft6DmoGty6XdB7NNe7+D937izy6q3Mqafe2+URtWjzgBjK
h6V7aet3bLV7I5vR+D8LPBK8CnedTb8SqTTFgB1Pkf0a478r3YjqTfyvYJsPHxvX
6CY+kpaATiH3R/hlpTtq9IF+mKYYQugTx+S3+VYqq04UZ5gzGTiRWNQVfwQJpTV+
3yAdpspROTs852rbI8uCCnPZ17/Dy8mctAoTWOxPk8UWXPorEg2SYpmx6s1XhQXc
gY+nJ7/Xy8zH4IUdTrreMBdFPzXDU98SQqfHNlfHyuVwTac8c4GsK6o4EWexGHOO
DDYzKqYNiLWb4EdJZCOxFfrum0yIfgE40+SFky3JFrO3UvUX8SB/X9wzfOHB43Ci
VKFNzsOxd47vyUgk0j4pN4kK4wMFR+eMt52dKK5u41dTrv1ZGcRLKdej454UEGMz
EzwnYXRNUYx99+nvilasMg06iqq0B/02SKBN1hFXFh79EF3D0YWhzlL1y70YYzEl
F2CpMVvgetRnQKnJICU2ML97mOb6j+4JhghGGFJeGbFoRA3ilBUt00bPPYnpaNNd
a9Cb0tRtuosrEuByQ8oIZcOVwXkZ5lhjOJtz5Kq6rs3AKb1kPJJRULZFqU+Vg1eK
7OWwXDuJBQei7WlMpUyUtq6IKJBEH5dRjFo0rTxPdNzX2kzohZIGYwUCQdcVnif1
2onDFKQpAiql1+qNUaJRuTjYWJmqwLNBmaO3+Ap7I59AUdidjg6B0oo5+5y4GcGL
39aStP7jO+CGDnCL043vjAwI4PYPLu6Mv70xbdC70UL6G6+XAz/4Q4OdsuH2G593
AG9EmJ1Dt4JNxGqVPcWgeDa59ewkBwXyH1+ejYyA2QmGxHbbpkXBIo0XRsOLE5Cg
v6KcbHQFVGG6dhqI5gtvV6MQKkCMCYr7WWHQNTRSgKCOFh8zJliEWbLJ3KOxVirJ
mJ5e+xLOSsY2ZltmvtiOyXK6zI7rZkVMv6N52z2hzfMG7GltElglcDLyw9xDr1rw
DT9QALqPUHCfaSEMNPrOkxsmS6oli6iPnx00W2Dd7a/CNZiYP0l4CRUrIIasvlvF
qjXV4A9tPcV0RWc/lWrreSAURpbm7pVmyT35/X1eDBmCIvheTkd2WUdkX4XiNuZE
Gj8tmSPguYZ14FLFt/0B/9eOuLlav1jgx5YwIJVVjqbrM/1Oms5jk8b7LF/UkQGV
+SKTUSTF7sETMU4hm+ibPElbJded3sULFbIEpk0gVIiDNOH+aoP1Wr/IQVU8BfCX
Pku/nn4sLhhx3RU/ebrlZI/hrTlxElspGD//Su6aMIfbVQP4JOENi0PZ6oliMWIb
1l05s+uGIKCVJ5wu02yXJX9WIzUf3VuqMJKuVdMZASKDzO2tYjXeXvKrBY52MeUC
/s8oEFyUi40aPxUK1ZJXxDv9Pp5qG22R3+T0jc3Ynljz7GUnUB7gD28M+GddxfkR
ClymUn0OjXMTP9ohbjaUGRUSe8yq+del29Fqq3cNN0bv6UV0Rtdaodpxpa0ojiVW
U5tYqoA5MTbzXD2uvcSvBXiEQXZHGIJHsj4JXZyKptQ0rUCSHnH6oHwWmJ37OHZr
e3apP1TrYaxqBxi5GyAJU+jOzEcdsIYA3TL7HbJdK9WX/LrNJzgYLcDabDLAfGXk
hHM6Wvx/FNglwMyqhsATx1TXJkasfHBlu4gp0NfMooIGRnBtkuokxJQWnEwZHqzy
WSFL6yKnoWz2RFM5oNhU32TdNxKb0DZ6DXIU6bVYn0sjpyJIA/7w+W7DyNJYfyCQ
Tw3r7hSp+ADimGnMkfSoRDnzFU+YBr5P1C1Tv2DbcfYa0nW8PYfrIjsll16PE0W+
LAnMbl1EEtznsUEMUOiA9/dH4OMi7kUkn0VNQxTgC/CYWqCkOjSPN2B5MxABu8QS
OOwvHSzjLDkzZeziwD2jFesyzg/oV7seTsdlsMKuFxe2eZF8lLmw5+5DtA2BDFgH
AU2nqsaGe0cDjGZnNf6kFTWmauolQ6YgasXnvz7R2R2UJEXShFPMcClyi7Mq9lmT
yVuDI91O7tAglSLddCgnl4KvqDIoJCZQhBkJwKgsftEn56v5Az3y1mPJ8dwT4hZu
eV4AfZ57jt1WxxfYWWScGl7eCh8520mxuQgdAd3xN+UzLuN6Fo79uDioBLu/W6Tr
uVPe8Q/VHFjmIL+0Lir9z/9+TGLemb1U1937h6DvNmIYd9HqY7VwpClpvvGEi7kt
L1YBpGiEpV0UaLBMgO1U5Rc6nk9F05UeimyZoq4I5ch1myCShwDQXL0rXhLkRPXC
qxxub5dtM9OIU2y74wcNIZwwkpz+txNI9Ts0duG77S7+bdw4ebaeAX4FsaIPdkII
Njqe9eWin7XGpSfAd6RvgE4eh+lo3PQEZ1R3UJH44DNwc1z6W1isquHSiYM+5jfy
JUjBJrnFqp8I/UB2PUUFLo+QkZbhDxC81VPyDYiTR3pOhQy3I3ZrTSXyFxuHrx2V
PEeX2PSvE2PnVCKWR653UYBTRm7a1IjlDe5Fsjbhbz9+0EANkt0Hqg7tWLcz5N9u
R6cYEOXUu48oETk8BhzWzJ9zPbbBYfOgHIqRNVbXUtRulTdO3Qgphb6iEE+rsdy9
bIBRpB9EVAGgyKTV0/FEyR66Wz/jWyaUYHaqFGihp6GkzqYUwu/iG7sbEGmdbp+h
4t7DJcI8S0F+COPcw1ecN5yzT2+6EuX2JIDjBGKHWzAbGzvAktVvcuZAW6zkue3n
FzFW02Qsa8A7RbhkoweKLBOU3CyyunqEXEI8V/0qCUdFHPu1EGHPhLf3DoN779hW
W1Z7AROZ8hpMNZME8QBB753CsVVy56qxAkRpJJSBYYLjPNqcf2S6U1Tkk2O1Jt40
MawRrLK/jF8RwjRT9lj5J6zBm281nSOIKZvKnXEyQmM6Ao38jYtdQRAiQ6qFfebR
OGFtAwaVDsw0N2ZIYAyUWmPlsoTmwnBHJ4D1blSFh7NhvO5b2eP2jHKOVj68SIIp
6OkiLQ/pOn10NMIpGljaOAvdHp2LIJUBetVkQKbzvfdXBEiWz3j0mVmS+/H/U1+g
FFfpfnvLxq1TnjLt0tLbx3Ep0CDa2LaCnN6xH/DBYHgDBu6vGY2UgjSePbzM9ope
kxjNjM/gbRYVm+7FN988bx0coT6HWxM7LjXTstxTliJpaA8821TLVgynVNjwAOg0
zFQBpd+vgLhY5veQW4DunPFzlyytCHW7hrxQ5WwAzWDWkVN3VaWtpPxVLO88pjKk
pfNI9NlSj+xiE1AUpzxV6/RYeHNYx2Cu5tBFBKKH/dJf33vlXKBlZ49LHYpg0IBW
dU2fiSgyL3z4JaUYbY6INGWYKTFn3yMdPX2HCJuvWO+JJ3iUePiiAlobl86VEivU
lE3o+dD5wDt2bZ/ZZuG7OiReBaYR3x6xmE07IEkWfnh/ks7fBkx5VXBkL6I56NYj
4D417hqlKLkco4TaMAa8E11fzutQQQvqz+y0kqAQASezsgOviQqhRuUVhmGawR0Y
nD5SoGVYJ7IYIaQJoqqLtJBEycsifGn/G5jVQCjrl5/9DAGUhaeGd2rCqCHbH5OJ
gsf8nUNPv83oLeqoJUnYyXbi4YsQNzpk5K2kykczWdSROFTd5uDzFdCTr40HunxI
6QAAt09eh6cJUDqivk24dONessJK2f+nRRGVX+T6oC6NUPhRXob11WZDbiKHxi8J
FM9AXbNkvrC1w5zjlQUUMUo2NA8NTrJgtr/UN4Zx9t3rramgHY99Gbto5i3SKlV4
XPY3cOlam13k1JD6bMhNPIAaWqSEVow9hek3v9N5ah+GvKXih6m2TrlInZ+A4T9V
jmP0qjFYsPZTfQnl4I1iztvkg9J6I6OflbgGyORR6f8U2fVcLk6rvZxhzK368z3Q
YxwarJ6xDVPMx+WEzjnukTzwFf91A+eBW5CG438QFJfv0lbMiodGtLDt5x7jNJdL
geXfIEHccnAsOsQML8QHDAZ4+pjFThtDvTDSJ8InH3njciqCDwdfU5AVNaRnneFs
U1Lf+KblZzmiNozS7GkVo9DWelIHlGm1Tu5S/698SuDH10AcdtKtAMeMwxskDOIn
lWYGDoJlaVyn5lNyHcmR1xf5cCHKF6iN1hjKs4b/IWiG5A+MizpU81xOftFsZWfE
Mor5d+b63UtjVj8sG7FLRT7ZH5z1DqeG1Yq8FNRY9bunpLnuxfm6r7NFn1K70EmZ
pmTQIMxa/LfFIWoksJ04GSKvlGSlPO/VvOw/1L984jIYuTnW4KX1QjPYzQZ8WN3A
6BhRt2hyTn541wurFNVHKZzcwYq84nHlpVJpaxfZTcAL5DQZWj6sBoMscLFbte1/
4tVIrLI7DbLuGzJ2PqaZuJ3+rjX95BxrteSmzqEQn/xRtDe/o7G6ZBFew89ExBjl
seHdlQW1fY7N23g/XnSrC2D+FKiqYQyEG9VIDF1MmXgK7b+d/5/0c7p+j028zzZj
T7MbrSDP2/nIsqhDqCtnsQ==
`protect END_PROTECTED
