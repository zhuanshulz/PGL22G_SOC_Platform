`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j0ICsVWVAuwbWUTARRzYCE+J2l1SqE9Yuo1uLSlTnx6lBnkF17joGL305b0GP1pD
FerX09Sw3XP6DgzsjYopF1YPMcp8kuftW7Scx3q+XEAZwd7Hot+y9Vg/K6vI+uo1
qvb/jY0XlmSwUZfzpwry3CovflS4WT0waFwfSZlVvqilNAesrktV8VSwXDih1EE3
btw5VpjvNYlUeQYipznnEv735Z3VPxJFRPqAZzE3hT2IbJL1dhclcUACcq7/hiln
L2CQhBoI648loQfMRzmbEXsJmXAiOWLJOOjqh6SlKqj2Z6I4XYmblp8VLJQmbAe9
7d3uoEEa5xPzACXOr5DnsJNQOmnFV06bAfyKHKpmX9BsszxoVMww56pf2kNUoK8R
KRDWR3vwRp55vPCKoGdKBw==
`protect END_PROTECTED
