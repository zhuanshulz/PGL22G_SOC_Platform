`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvFSfnrwnCeN67Xo+lNInFnMXAtiI4JYGv3O1SCWeD4Pnd+6gBPYCt4aVRFDGhco
Vw0Ew74zbsaj8ZustZhbGBFRZQsGpdw5MbW7ZMMUUNfjpCm+01rOCnD6YoQ9F6b0
AZBSgAQF2ETRqV/1J7UL8/GIUVxNr4BeaLc/R1C/jzK8tLz1GtFNA2KiCduJrhxn
iB9VbrOL/izACA1JF5HuujD3inJ1Ein+utM4JSRrdnPk9LAwTpiJQZGGjvyer0D2
gNsq3x91wws/WWIYWQitHHUgHc19QswlFYvbE9SiW+Pv5O3xVFJkDEwQRfF8n/K8
8VdB8X4uElDqJrmtz1VVjZVS6eCCN0Wv1NWJv2QGaV6ZG62TQtS3Zce1L+IGWuHP
7gtV6PbYsQF4Wq/QA27z6/AYorxEvEEBB/flQ+f5350=
`protect END_PROTECTED
