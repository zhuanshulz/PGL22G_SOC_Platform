`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJnCRKNdK90Tsop5fIxRq8Do7h8tZV6Gy71uDOkBfKczBO0OLeubuZSC5YihdEz/
/SVkLxNUQBCj0n2l8vIpVTlt1UlDvLxfrtN5Sgw5UNqx4O7Xfv0D3jxIsREa567n
kDuLudlyitI5k9e9LVmtei4TBK1TivZ77qZECT1ggBe7wDeYBuQDiEs1NP9Wrdjp
rxmlbYwDRqr7EmLHb9B7xOeL0/S0T1DEpA36OT/mJ2aAP+j74lmQ2yAFnKD0ORMV
AGrBCXZvZ2Z7mDjIeSPxsTIQIcuxMX3oL81Gv78//nLNGvNbynEtJstGhJbP9ylY
BDBXenfNFZ0/O9geS6Yn4Fv8iqvOHWd9d9DINBEoxemH8t1QAMC6F6jNP7iMHqkD
UKApHffQfwOvCf7H3uik82uEtRpiHO+cMyyGVQmjui4MDp2Fmgywu+gH+jnHxHpw
wAI8kbUnXKdGdM93vScCoGC6PsRN1lAiET24xKoayEX45ODOYz579mBhAemRugNt
JKvxR4zxi/sTEmSqq9bxTtkb4x+1t3LaMMX0bI5LyeTAsbrirJnSYZYBV84GMLUc
zoMFc6f/s5J+C5bNb5c4LDWbc6jMFVnhfaJYTVUL82SjkMNsOBCIyM0s33cXOh+Y
ukoS8w/U74uUbH2eB/TXikyamcZKaDd00+V35ymcik3IpFzknMPaZZcNdfUyp35T
bsPv8FvDQMXUvwPOKZ+ufoD0htJ4a7RErYB0sze5JURM3w19rpjX35u/Va+soXTq
SZieXaUpvco30pT8TLq962/8eqshMTwXVNe5U8NX3WHLgU4bckVyQOtPp4mDdD3F
AuqU+A5pgX0cqaa0Clwx0AkNaCsgIFTfSyMebZvYrPP805nj20toAY8qn1WssWsR
G2NDZcSwYIShr2q9ywlKSCFs27NyKzWQgh91ZQ64jhq/J/Kw63dF8CmM02fowsEh
wiwsxMnBRq0h/3fl5kKDykLtJkb136/g6Fv0ia9GWqmwk/2hJ4LKxKSPdtN30fk4
HJ3o3438Ms6QoxWk5lS10okVwN8WU/Uzhag8wE8LwIefSJ8z/mZXSPI4qWs/jK5F
NylG8Jde8Wg95RHQ2guwNSpoYvtPEDBLDfsHRa9jeHNnfYcJ4II+4o4ClfJ47Vjq
6bLoRIa3az6CSBJq7Yd/Cfma7ug5V5pzAzWba2eBjy1oKLbwfT4+gWdmDUE7WeXq
bz4bXUgT/3knqTlW8jqttA7ijxoBFlHsKxkl+Ek+JStm+l3KEW7lEzl/VP0ihjZ6
BkMEjorI/Tk70iIVhpOfbfFbmPQUbuFdzf+waVIsFx+jZm7sIkvKXPBswsZSminA
uhGjR4P6MfcmJxo2DKnYox+nFHEpX6ytsQtPXd9FPBLIWZq3KEClS5exZsabVT7w
usHWXocIW934pGbhpFtcSQlKUW9gK19zfYWfX27dxUYes/T6vhHi3ETb22HxIYVA
B4ussLccectGQkLAz4CT2IuAe5bNfHFG+yjvQ4NmpVcmmmyFH8UQoHOK+qBfUrkI
jzHeMdVox6otMdwVqso7iEAmZEWmII4m2DulA9z8yOL0PfNn1LCO56k8V07G0wqT
LWbrBzTxe7EagPdhYHloWWOnYmfrEBgNniHTVN+bK1xkVrL3YC84lTliI4VFtxC8
oJk2trBKpyYQgRZPhl5OApyp9YXD0VHKbLh3E2vtpm19ZwAXxBrRrLpIXxR4u4qQ
8ndETX5QVo8RX6GSwvCyCY3eQyJrrU6mBvauf6RzqnGXOP0WcWoZhfPIIW+3wd5E
DivdVQD38PmrBqBAPYIKxSnTNuhyii87CufQb0oRUrp9h2ae3c+3LWSa7+D7g9px
QEkrYZNi/WCvCuSaLe4GDFXhwfcooYDnQHc10npIjoqei4OK7km0aEXqYmI8fC6j
L6V4QSOTFxUh6i4VUb+65cHIesrC3CCGBKZAye2cw1eVOGFS42VzpT415Zi+Nwe9
Pku5Avf+czJsx8ST877/AdB2yicgbgHjvZVu9x67opinRbaHCMPIKDy9w8cTP+Bh
tOGAFhRO/FE/TBvkfMpO1jdi12rX9l4HQgQPOUx4irDUnv1jWCjQ9eWVNejLDnY/
v4gGrkbyAFWvoVb3nd41pjDmeM9hougLCLNu6gERgTzKYykw+2XQHMKGSkyiRqiH
WDqSy8jshtw45uX/VMUrAFOzaG+iC4jvF/mwAoGe9JPerVEBvPgrEi4RELBpQViW
WZeErXuzpPvWiTmUxeN5qEeiUT/or5J4Gkqvd3f+mYh2gsFxfexcVZNsuceDO5RX
AziY/YOs5BsfShnOOk1UWd6z52ESaJUnb49eNLOV7qqzQ3hZZNojUJyL4i+lo6Ls
zedMh48EnOo6epurNBzhAw==
`protect END_PROTECTED
