`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zu/RJ85su3I9T0DbCE9yxmO6qNmOsVlBISc3mLL3q5HKsSiu6stlYJF9gtDYmrs7
t1WZxuZWr3fG2kjH2iHCG1siAP9FORTc+19aImTAexFny3Jjl05hb774B91LxV41
9Ek+cnkvmybxWZbQXFr5/nmiSQY/zVAGqWbeFrDHFGoSx9FOjn0HiKRQQGkDKLR6
cwEXLqVS6k6GDMGRJ2XJxhoyjMfwQZTMWDBWJCj4doLmm1W23uQosbtXkfteFsfO
az6L29AMZz+Qei9XLDUGMUaxnhaGaTv12r267co/sHjkFNm28N+c5WP2qSQO7VkT
qc36sMjXlj1zsKKpyqXm3Ydkr5R6TWF+DPnLiE/qSEE=
`protect END_PROTECTED
