`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/3lgfBTkGlMd1u5ttnp66t0LQbHJoDFS38uRiHZ05d0fZH+fj2AkJEj1MtQGHZX
65OaYHlE+uf/2O+BlHoOyYyaVXT1WFy7BytO8YE5pjojEXFk+qXkmFU8a67d6G4Z
EH+YGOM+zvv6TGdXCzHoRnywkY4CtNtok8rsiNHg9z2fVMYNcyJ1hJmdehlty6iY
QeqaX9GGQkcUKRa9p+RQSHmA1UBw+vdnfI/e/A6nTI6toWqE1EUPv/SIJMMhsAxo
+Bkfl+iOKpu5mMb9eFGU9D54i/LpaJSBmpcpA+fmosqhuHvrZfCfIzLmf4LWmIm7
aRiNrk4Vr8mNLJ6Y/s0RrRtWEg58Gg4wdNAlYkV1v49x2+OeLcMeAPpfoNOLsSee
YiT0/6hogf/3PfQrOAMF22xKGKIiZTp1cra00xAHlHlbuMjvwf9R2thDqFt9J8Ko
NONx9j1HkNpYlH/9++xYoP+dKJ82o+9nCpTUahZ/penEIeKDFDe2PEsXLrWEiSPB
OXIIKtr0XDO92x9KcLa2aSs8tdjq753OBs0zqrC0FxqVDEro8IIFB9TlqyJdPztD
PGPdomv+55QwKMvbq1EHDwfP5dlOkx+Fax1kxWXBVxMQU2KjERlXYEZxARidZ2CT
SF/Lb/pikb0vdoG4r2BGehlb9gDhOE/JFfFE+a27SXXrhOZ1Ggza+NKHewSFmCtx
wO3cO3W8v02l+fRa+ir+xGAEh0uWOb3EV9Oj2+9PcgpDL34QVzAGBlbMuHpr9b+M
X2RxIMg+cWWQCk8siAR1YsqETWROti/MeZ5NwZhGR9ZVGQngsq8wPdQurF3g6x3y
NcvecdgjaQlUvuejtwQ87CGUbXOVYNLe4ZViXWi5yhbTFhBfU9HdE7djlOr5xmUb
6M8XcZTuMxi4KlqJOqqwSWRFuHkAacdcWNm/sWiUbUcUVhvUDkA/c2lWjndPoBBq
zp59kdRlm47esYqGzHbFYeaRpr7nh/aHisgG/3QbrQdrzZSo1RLZ42T9AVLe/xo4
EHlVjIpsIGQnIopnkt2p2O75vV7evUbaFqWwdJ7MxA6NngiXzhqqin5WNy/VWdYt
X6spINMYVap+hIn03lsKiYbzOXX6+coOnLiOr4k6OjaILQ2UAhNniGyffMyn6/Eq
hmi3Jkxs7kjwnpt5xUNqWaH5Hj1+JCSIPQi9OMqrkE/wp5P1Dk0bwEnO1kD153Lp
5tO44tR0rasktWXIXG3OT6ZIontY4j4FoOYLf+kHw6MHFCt1YyrCA6jZ5WMoDL73
YMiczpLJxyL8NuKDkHrMTSSVdrZKfGaAtsCCSQgUx82Fu0oG6W2AP/KxjW0OshPx
+ad8vVre1f86+xjJGcd2EF4LEk+zKMnpaLbI2DknoI5gLGV3yFrTCX4mf4P1SOSo
eDNZfAJV/+lybCqx1J2XX32O1wpKHnZ6jsWA6Am6YPUWRYwYKrUqITG1J5JDS562
N213QVGSyv0h43+SoRYR32xzsO1ysUv4oEWnYqudXKQtmTZbCtAdpmsVYebjvOuI
4di44e0s6Q2nvuOTKk/CErJIVJwLJJpmVfEvUe9sLOlHOexS3pN3DgiCVhjCrpJ2
l5bNdCgRWVk9DIjQj/1G831+OGySDhmCiZWWFSvFIchZG68wQw/z2Ju3Wv3Cf5HJ
IbPORokPjpdMufpwTpEfvFfD7rxhJYDuNtfTv311/idnHxP/kAN+R1FtfrA2+0K6
9nL/2vP6L8xCBHELrrNMjDoo8kYz2PGiBnfLQ0D7X7GKaAphEXsPfzsJpC5HY9SJ
zSihHlGT/MeV0Q2+qFLCIMTWvc0szshmtkrrLEa73ORA4aDXZT02hHBvd7kXwm7z
mEoarY6g30ZoFu1/nCYOUPJIi5j3GK9GXfgIOyNd7AxHKBey3fbpTAuwz7cBn+ci
ZjImwszxzuA8+eY9RtfDgs9+jJrCB/eUOr28nmr75gpLwy/6wVkW3cOlmc2sFyat
J+1Hen6+bWlH7a2QhMboxnp7zAQCA35hs1kKI1DslpNyofXT6CvTyyJgRIik5eZZ
97eWI/9uNtzFeYmDiEKR8Xb3INzI3osEP3gtuqugCV+8o6oPtkihZGBqM/ijPJEi
jQOIwNWVvlqjAEuV3DLiC9daW1TC2L0zUxPq4qUW2qb88lDk5Q96/lddeQrbzopp
swB6cslpgaEyA1GkyoSVFvBhRVNDR9bd09O7UacpwFiZWIhV74Zo4Zy5wHpPJIYU
rf5QNYdIRA0jDXo3uS+3Yao9VyLfMgLSvl/FHmoTvILx1E9mM+ZAgjW+RhJSWNQm
8eeQCR/2KPUcloshXsU/xluChcovYaP3YSgElY2I+Dco4Ll0w13wEI4R/6YE7QGp
207VOE9NDsQjtK7vslOE5GHAi9irur8U+ZwR4IXXrAVXNDJRYLn1bCAVw6lfWHOB
7akegs7XUPasRhcKeReVUxzaHkMYGs0NcPvTB+kDfIquZLWiyOcnUQBrZ9Cl6uUH
LIcjlUax/+N4FtCxnXRiLx9GPF+U753zETCngVcilwdkq2avsMf8nsZKIBIk+VwA
jwc0BuLIw1vJYszx7eV4PcVOmn0r9KTy7wk2Bd9JRWTDN+K1JHIddmNuBM3GRn1Y
2Ki9E0MzgkIsFyuMF6BIrGnP4gE1N28BPgsnavH+MrmEEWlAGXkai9DFM3skNiuq
Efli1OW9J4ZuI1hLH3eQqE+QJubwk65qKFdkjSp24tHoP/S6yuEed3D97EC2+1gm
R3tdlVXKfkstc7PWryLUoFp5sKfB89Xj3ZxeOitP2qaqdMa82S/IYQN0ky7CGP5e
q7r45QtlF3B/9GmHnY0ezARL+CSdUZxKhua41dPBEcOIDFNzsn2iHXBa0VzdR+B2
JjofhXnHrXJDz7VwawstuqVNEwufRx+iRGvHlGKHMOkdUAWeZMO3l4+0smlTXcPJ
uv82ULvPvGz3VqpziUbxahWIGYp5+E2q8gJItJgk5JJIGzEOMCM3cHKW3hGHg+D+
3Vnn9Fo4qQdL7vzv7OTqNIvqdpk1uReNA3sKzIzcYyfugxDKvSvJC04JeGDp2k96
TpXmXu36mJGcRgADFzLlXO+bLL0Kz/MNMJqFoUEe7Gh79kVbKFUZyRM4m4WxZkcy
VdA5my5glxtUzGSqI4XQ8IOyx2wdjbP5dngen/lU0nC7DiuLE6L+PSfzdG44DbUG
S5CjlF3SxKfLDasPVPlQSfDLTdKuLlDp3k2k03Emm1lqHd+TKVHPLkgssb+S+xZG
Dt0TNB3LO8rdd00Et6F5xglexER+zITWZq+yZ0i+Of/3nhNevX2uwXCCEPXdOgIF
cZWBc6MD7PdSHoGZRAbqYSWzqPuqn2HAldLdQERRJGs/S4hjVfXXTK6rFCtIAty2
VhbIXxvXl97SXfLTQdz5QQcf9fpdoraKPnJ+C+5l1nrFcGrzU5qIFefxG+uZQlvu
G1S8J/PGKw5OFwkLIfnZNF5iP5NAFA4pYhPjwN8bzRHZ+16RhmGUTn8YJ6hnN39O
YlmDzpti5VhxX6cIErAp1HjkRWon5pHezPPCj11jIkjM08GOfBqQnnkSTxrrOF3x
9icHvY4E8KG1No/7DBAqcXITNB6yXDPY7Cut4O+Q/eKtjyyuJhwgboYg7fM6jJre
ujfKtkHkBUqObUkQBMV6orBS1JOt7L7vpAFSmg46YvmYHRLkWdGuoGCSZLUfhrBL
PS2nNLHyEvX2ag3V94OtZu3pZwJxsiyxD3tT+aSwypECRPgyNJQ+Bg3OWo2Deerm
ZvhHzn3ocKZjzsNX70kFbj20FutcubrftJoxHDPKDaT0w5p9FLOMY4ltTr/mVtqu
MSYqfTS+uxymgpIDOVGkzu41hAGmgfPK6LrHB+MZJKRBqa2mqx6OIKNYE1dYvzmf
U4kTs2uKfjB/mAuFjjQz8FaP1dxZHbEkQ4H++5NTMc+/kWUVv8fwL0Ii63hMUft8
/7rGhIDKOeTAqVE1m0npWpuYufm+qx6a99Z85YSoPKvNiBZH7y/fkqEoeaH+Mffo
FwY31gs0SyMAf4lcasKjixTzMG1KNwWcDeH/8NNMjaursz5o3h3uJfheQ6N/O3Yr
YXYMJ3Wb1Qc9Dd8BsGtF8JULIukb6XK+z766++FsS5KBfye+aLlFoasgrFGjCtrM
yNuxp3KBV9g3gvnxr0ciT+ZAtGFWz8OrJLHaVmzviuUG+9/7Dh/0XZvzXPkqO1tC
dRcz6plqhEyRpnf9VZGSBwGpOH6xJkdMtprtwFRBnxNRDCGtXEqXcVCSrdI6JIy7
CbSgDVogIFbuJv8QOCILY1Yjj3xmRZ0GGG2nUsBFERHqGvRqoru+ZpwVni7oqsn+
n4IXVVqClGAfQEQYteYL3G4lr1m++Z9B+zuOU87gZQ970LAgVIMNOxwU1Y0O3ho9
Vvy04Yi8n8gROKLTyI38yf2MMIxjnDHNkKvd8Piugd0QbrqVCiNSU1AQ3THEKO00
tf0DYDd9Gny88g2+HFrVII17Yl5dr9NAuTQIvdX5S+Oq+0n1VVmx0Jbtb50e3RHH
BPX22fz+Aroa7UeiKqH+zYcCZcqYfLIgDCQf5yvmpjm2nXOlPWlU4Qoip6obVC/u
W3TBXnpOgiddinpDRD9xDiyaK4JiVaz3yGxXd3ongYf58ruhpWOuk7dV2izS+jux
L3zU6j2zSWw+u+o7DaJa0J7epuzdT5sd4ZtsDqHHlSadWm9Y0BzdC8CQFaR+zeuM
pSof6YBL+FJh1NWYD93y2dftr6CPMKSGkRqQZY++xGa+5daHE+7LfArFFBZSovmJ
cpyu1S+JVu8NKTIH9ZSsMCtg+a3JoJEVsiomKjlkTQPBc5HM86JdudlzgwYEJLX5
h7VNq59o8cMwbQPeg3W238anqbB5ezagbwttDxeWM872S6tCmvDb0wgoTZB5agjp
3VSFHSCojbFrsc4nWVIjjd5M6ygQ8VAPtuMAm4remtujtutvHpwkl3KhOfg3pkuk
vNg01plbqXhK+css2tfmnZzz7OZ8IJCeW2lWQghQHbPMhj9D+bUNmvAouc7vfwMB
8HeE1wLQxmA7Xjd3YHeISzLcVM3XQwqkmdpAObZiMlqlmScaet4J+hJKbls1+pKx
hYj1pvdY/wWjU+JFoIJFKm5C1HepDhLTXOItxEFtHlefBEOa0nkcL+me2VcviOen
CtMfYJ08O4OLAgZGnXZm6bdyZLvIjV+GcF5FyG0ACI/xFdXB47l9ZCIjXOhuUnm/
UWEenqxjVIaYZhc/mf9jw0Ul5dpqJPauGVDA612bsLVO2J7RmDWIaeNPlUA/FYIi
9PJ+bmjWmr9MXBmmphalwDDqwbruvV4Ykb30fXkAn+1cw5WsvKz4YItFCSXonm3V
Ia8eYlgedMfmRB3IVtXPX/h+yHPSbXSffUYCiy+0urF8RSSOnQI4Ekn/mJSfZ8jh
/ue58oraWHUaJ0NqdsjqraQHSnDM+cbPxOYaUFkVvhqQqbi9tlR7ePO3U/XTMvJM
hEUJ1U3O4KQXIQ86Ry86OyVpVvna/Yws/Z+mUkJN4IbYaLZYdK7WNfri3Gp4pqUf
EoEJMG9lhCu7I6pUZYpMtzou6NmzQw7culZoSww0IEVAQawP3lwH/erb/hc/bhAA
DHxGhEGQKIAWK+0DzrG3yj4Kta1W8oCw5yuHdqaaFwzAewoOIHgZJCs27k6CzyJF
2Sougqax6PmN7yts4xiENxU3mrGonupLu/WbaEF6aOaWzH2K6qdRNrX66e7JkhH+
2tw94MJqR5uYIyQXVG02jKUodBDfQPTFKwRlnxAqvRnBNgohIPqhPeRP9wJdIDwk
/ZchEwKc/gR6uXLGc8xy6BNTFcTc0dDOGgoBfJX1b8C/u5F2Q/XzjH9NXVy1rbMe
tkiHVajdKhQgnHcU+LdlODq9wmSFgQ8YuSqQPgShjYQzwpAeDqLHz5p4K0ZwZZsK
NVF05r35ZXfN6Qxy1I/9sCEm2ticDSpWbRdnoQTWH+Nq/+iF6ebwZr52wRIt8dHR
t38dz2mZx7DbtIvmjR+TQ30dnsEsWFV76kPyaZizBFDD9CEfLWkPxsHUGcK0ggCE
lKfQ++slqLKXOPIGy5nAkblshwMdFODlb82BRFjdru9Z41iMqxy10eUKrrfm9/do
S6kyhD+IVpxEeYMH528SfDGkDvVggRFkgHHZLUZdbd7hCkGwOmq0QPrpfvvlxefl
QzPA55m6P+NWJl0ClYIz8dVNXSZh5dHAMvTJCwZDwdOnp/3KyERjNxSyom2ow2F0
tM7f/i1t2i8MkS+G3QJKqSAy5p2uUYulSMh4XhLJ9Cyv1CY28cL4E/qrWnTZfVjW
p7t+cewMyUQWyHHK/IwabpCg7gcKTT4Axo3WQRbb1niNbvBdQ1rVfPiMSPk2o1BG
VUcOCTnYGNsr0DO4C1nQH012W37ukA04YKHljaiXX9w5K5pypoRt77R1uafeGZgQ
17qltPlM0aD2COKSr/RFLf5oOjZxzsE6DaASHDA/7ooQykJ5xkMM3UNmY+IPmMHE
RphUsf4opL29KaLJ6DeVOvrPeoUXPyh8vmpxc/wvf3yGkYF2vQY8hTd2FjpvJcrU
8IPaXx/F79vuTQpP9n0W1Avgg50mv72U/SxpHPs1vUxovtgvoafbL4/fN1B3zGFc
NlBb1q0p4tUsyxqaZhB4DDh7cINmLOOFOgoL7c5HHt9vLke9eI10hySFfWj20XG8
tkX5z1TEgkMbBm9lI1r3b8uuNKuzYjrio3iSMjR7z+qIh6IcrwsaRrCxcjTxDLUa
vBJ7rIcg3BWK4L6UZaQAyF+WAZ+MxOCcbYFyKZr0HPNn21EiPNyuiGH7RzqrUpnA
7ay3wQQt9bZDSD86yScwz9mIMg0p5bmtVEOIJlLLlLwG6Y8PHR/l2ccMpWay83iR
HeMMc99vPpCeZ9ZgqVN1kRmc1UVChUfRetnrjJgtknYnxnasBiIE70x5tbnXwPvy
Zeq+IEpo6Grh67xDOR0v0WXIPVX/hYJvlLIs6fWv5bOS4N8P74AhDCBtrOmlueHm
zhhc18Ok/aJSJGiPU6nvdKPWhD2JxVWPOLA/Bbo4fJ5g3q0iqSJztmopwZBANpP4
DUBlOYOR+AZLXdGy6xPPxy5p6gWpzheBS08YnvWQYqOfgJ+l8/jtSo0K3gbzMz6K
JtFceXqHFkZx9xR/N0c/ppDGBqXkoEZ5iAlz6r0M4xcpBoicOqYAjy1TFDUMg3+4
ABZ+t8hh7sOwoYcuM73D88tObncd+Mr9x7bo9NSOgH5UExvezj0GHv5AV8BSkg0n
ygYXqOHqBUvDRMHcniQwdI5IbNBkFnjc45QfE8mJ4Fz/JTSDiUNm/MhIVtD/AGbj
EnzPTO4uSp6e5WC0Co5r/BtPpaa8xuaesjc40ILyNONUM8vOHQEEaCCdvzBZCTSL
ajczZX0diAKWTRMQebdsBuiVvKehIeAO9dpP05jKVa7rfTzqIGIj1b/jT6QHltw/
+uO03LwvC/V7eUlF33XGF47hgHlQB3Kw3GiCe5KEAMK/0JflHt6Rw2I/oogBhXVu
9qnNtRMGY6Gz/MyQmAS4dq7qcE2QwRAmw4gcj52Q9eNXPQSKNr3oyWlnqq2RtSri
Y/ApdaEre/qxAZSmtNbyLly+oZKm1jJ2m9w0gsrZSM+3whjaQ3aTDpTyH/LZ2isM
YeYQRodnv6d7j+Fft+gEttQ0BB6ayyeBnkw9/FAWDPcj4+S8hBu8p1XmMPtswPXL
fAuW7Xo6oTsOTmY9X6niU3zWOcZK6NNbVmjqfmW9cYXJEol8sA5H80jrzmDzxtd3
sq1l5bG5GrpoDjgb4ZSCyuuOiHU+Nsi+cVTaw0zA7JOUTgW4/SdRXrVqRXYKutqF
km659bADWKLQuotRP+k1qgd7eaNDgRc41OSfs9CJZYH9ZVJLNn8iRG+z0enM0jxB
3oaF5c5WGPXZe6pmsfRJL/Vi+u6/j3ESajqMz9X0h2P7Lkz/ma4kTEHwISiWO3IK
4sGRFNcBIwShzQOOoPfn6tJnnY5php0HtwsuBsewmgQ7RtwhEyjtkAJnHTmZjenX
kxQKJ/jKY3bgmMQgB9HI5hGza03nOAt/x0GL7li7fz8as8WmhHW1Z/w/rRwIsHcP
xhCDVtQQTxikuOMKz3e7rtoyYJsR1U/tGLwEJVg16hcwRQ9jKAcPyMNT0o94cXWC
JVsycUP46Pfp7exFkgL/mHxnU0MQSK1MhDOFqD5IuTpmMU9fl/Olo+kp1fRza3z3
1HbBgNCzpetK1Su1x0IoD2G3/s5TMJd0LSa74izxulIHcvkW8wYQ/LH9sB1VHIER
0oZihrxcDzIRyn/ktkPqECC/g+8JikHktq8IPqqKoeimJSeUzqNuqk2H/9qkjQiu
ffvfkUIqdOoUD2o0m/ZIJ9/jeASJCTCk5VDL+SyS0ULO3ekLjVxbQRG5rpsydWvc
0XmQZh5OT5iLaBa86r/AM6mx1Raa3I5WyEDqbshOvSmmNznZrOEaptbfhSq09Vdr
Mvlm3Cb1cy/ZP1d7y3pAWMduT5QbZBW9nnSsbVTvtQOgss4wuxWmAO7Sm+OGXxwD
KYbOMYhs5LeEAqBdKTiaYfo6j8ERt5Vio1cbWUBUbkSROMGvJ6J5mEL5PoUnZ+Pl
ZzMLKnLehw3Mio1M+mP2UmG84TGS/uJjgBX7W7o3lMc8sVn4VEDgItzmTtZKYxhY
L3oUJwh2BJNSPCbQzJRDaG9V0O/jGxCUvYKuKh9ee0XL9qd/AV9Pay7NhraS1UJ2
Q/1i1Rp5sF3QT3T8cS6MH+xeMbgxqPBE5UbMMLIL/yhnFedp/Dz7FFq+MRSdA/+i
MIny4adqjamvIYP51ix97kgupg1RAs3bghT9AzAx1FtBQ50nFyRdqIi4EeK+NitJ
c5YYIxP7n3VUbFqSmu4rxsat1Xne2eWpXhPhFSPa4m5OOVYuh5gL87KchPuOYk9l
1NFlcTsil2ZBNyn5Eip1ZP0yDpunFQyxn661kd9A35grH6Spq/tFc0cZFTAjUckA
GzN7pIKxFpcnl7FMrv4TuJW7J7XK+lkBu8L247UPlAVaf7bJdpPYDXwn++q49uyv
jmhuaN1j4mHeZ+/4K+SQ8C6hIykoYiABHjigo/h8Sc+mJPuHGWHGbiBgv27+DFXd
+zfdH0Hq1p8mGQBfkeI+kfUBBvSrsWleFA5L3ghHfqTmkRk9m8eU7kpNqVtEG5oF
Nzq9KOJ4ks0Mw8mBCpks+fL0Zx6qtNCYuBKPj8RNCW8mnYh2xJSvdEFVW6LVygNF
R9QFT1tNXv3h5O3XSXr7ZonpfGgY5ZRLz+g6CD/EctgQkt/GREKm0IRTklvGk75y
nckgg+G6ooQgIhLTmEvH2Zln+/zotAmJNzMPc/Ms9OxrGejcpoxdbO7YA0FqTIEe
jXOletrJLjEGjfxtopgw6muIpJcxjnmwrQ/xv7LAGuMtIfNIDQnUV0SGhaQDwd4x
18xSjLp4OiJZDqbs/2GcI3FKKyvI1hCqBCtQXE3eWyA46q0MfrtDL/3071gbXdT+
G6FFZQS48DUlWn1UNphRF4IoJs3QI+TQpZDM62l1jS6lobZbylHwA5zrM8ZJ1Ms8
6SzNdsRitvMWzOIhYQx8CsdBT3xhdkLSG6TrFkhuvvKOUsn1/s6kXg/OJJsSyrIq
Y5eLilH045ULGiV+NPrBmWivvU2zVbpJQK2QUdXNGjwqIU32HU71ZhW8PNmb7f0+
42Cvj0fusNGvEMmK3O0MfreiZfb/ldO3uqjQ/qP07ssbv62kvKmOK5k3Q1Cyya1H
HyOR4HviyfS6xYetL2TiB3JUefxVWFx/LdpRr8MhTi4ALGgEVCAOHo901Xgiz8Fv
DXvkxfnEKgaqwQ0DgIXEOHgrTLr66Cw+vakL6gZrF2peW0gIIT8AfTNj0If660rg
1z/CVgQhfeaVgaRhdRZjLrgc6JzxTJKCLNdudkHioGQUem9dLcLt6/TMCz8NK5ZX
nUlKqc1W7T/SJ2IKKD5fjXFmSgGstZifT4lnBMueEBJ+iUrUoIhp0Z9cEGYd3ioO
D0z8Kk1h3/IOagO6a23k7nYD8FkgiXhDOVnOBRUOPhrpquiTZi0McdCgwDQzu+3W
aZ2m3VynIeAT8KR/OBRH+fBHEDqG+uSt3hmyPwff9lTu7ws1/5L8CW7YUlDOKuC+
uRKNxA1rIbplVRyDr7RCxxGN+qgVv5O//jk7NZHOpTwUAfiycrN7MoIeN1VqXtWT
HwwDtLtj/Zf7Fqr8IfTSxg0M2L2s9I2zKkSgY4z07VCxCDTPipDS2B5QnVy5tXgH
PDiMg4K/ZWmT9Kdh/zD5xcGhVLUQKtea8S4geoAHb/KBb+Zqq/UAZiikZHdn8wLR
SQasvSe3QQ2D+hlgBpQvC1Lpd3oV79gTsEIwwN6daD13C9Eel5gm5Vz8n0HVRMNt
0aN8rOXwUl92h0wyb8rjhDgai1qrqz1PhcbskoW00trOyO+Hov05+hpFAKYe3IhD
5IyR10JZV2vg1Yw0MniUn9zMyZmmvPVE+F2wLWK9U8uAd3OK+Yh0TcsY9SlKeEcz
2ZzHkd4EU2JKxK9W2nnpo1wowx7n4om/i/CFXqUrpP3rcv39ByeZcjnfVuwds3+K
NkadqyH3a9MvJ56ip4MG4w==
`protect END_PROTECTED
