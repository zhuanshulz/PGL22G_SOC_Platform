`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwz5NUvX1ZAKswQLwOFrA7qDwpg3S/WQQ01j9gdVGutCRwWv/LbKao3i6ndXysVp
/28twFvnmGna6rWY1gzysEzx6K/ixVBaVF7jwTWR+Al82HhR5zMq9WG3KTsl4fCN
Iz6CJM3jirSH+2JVVXPWQn6R9t7ymqj8wGaCdu8Jd3ujKCRq4wBB+MYOyhWoLZqW
rpnL3mfVs/CMHfcOYS7F6GndP2IUxNHfJNtKUN3wrWgnrLQdVU3xG6xbtIX7rO5c
KRz5l7ibu6HLAcer3tVbhXV79dUiZhwo0Vqv3x9+1YhnbSWz6YrXzhpVlSsgh9h8
ghsGO88sLW3SI9Ff1hnLgLzd7xgZ7xxgULzOXkVdjSKWWHSk0xNhu23SlmYEx2h7
L3C5wPiA5fEZwPgAXx3xcDDhHbCZpFP1TeNB9tGo2kAQ+G3d+w2zjUy9nlzSv0xG
EG4PMquhj+WNvpnK7DWF+k4F1/02DkiCVk6QGg6jiBycMsdJwV9zG2YUlVqjlpwL
1L1yBxp/wga4Qp5sflenTJWGzKGbjSzo3v/MDU/4kRk7SlcdhdBzyXGkVRX3ujfu
hd8AnZmpXRtLJHeSEvJAIu4xXWE143NUIRtrrzLlcyj8powCFQdS/B0mwA9TZPy5
kgv3gonqmZqpB+8P2jmLrFdKfVPcoORljt3zjZY4c+nTPMozm8Uj9V+quQtZSowU
MceMtQBj5DQpi/kK4kuvHqv7OXz2l4Xiy4Gzdyf5RC4UcUc+Ag3nkHIqsGiQO1TY
e+SvXFi0vuMgCMqKVuz40T4Qkt0k1Rs7KCt98VyWpAwqBK+iWI44+KTStb/jS5bk
RIaKf39uzbkvyThXIZFgJV1RqwGJcTK+tnZP+/NRWdHtP+HhY75QdUOokI58vCc1
E55hs5SyQYS9On8qJQqPD9rhPG/YLC31Mphn2cwmHW+7TNloGAeuBVZGisUoAC7V
`protect END_PROTECTED
