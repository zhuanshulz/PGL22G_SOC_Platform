`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dlhDMytRfEXTTJLha/fSxzr89BgwFEZ03T4J5rl9k8o43TA75eV8/SpV6+acS1zx
7Fpj5tHv1fE4lbis74Fh6WD9RFY5lgb/a7rKlesd5DFOQsQSzu4jStOAH7rslNLt
IZZ9qJP3tSvCFxdY5CLwt9SWaRtxe8Qkf5ci4Fp6qNqE9UNNar8PYHvbbjchpFcI
+Yo1P8zUh/ThEudyjnkHYUTHSE9hClWHMUHjoNHkE1hr01KzWRMovmH4e9XKMv3L
0wcYiiQnCLlGCDdYVcfuFLSRIv1s2DMQkZLERlTG01oUnCE3qrZ7YAblg9lGAwDl
cnhLJBFuYycufFD6fYpC1sBj0+W1Zz/OQt0rWtsdjmjrm4CeAE5Szd4pUSUvShZL
Sma6KAEJNGNKFwXC9QMibQ4uB+Z1hNFH70CWnkDcK3sG+uJTxMeFd2JbL9BJSIgl
Sd7d1JgSwx4nOVaw+q3oGtL39j4zUdAoZPZS4vwSkQKvlcMN6FAKR2CICrUHZtfR
Rk6kYkSP+bikHZzC6fHEEAgFpFLoAw36UOq13pmKme0DNFCotr9mPYy1qicT52HG
NCQ8Pw43IcEtEvIR8HeAWB0kOscKnBibvvf5ACiQu/m8Nz+6n5rCs5LV5fVaK5m2
yyUXipmBbzIjyq9mwvyZc+Bp1hwBEaRbFLwxCwKtv7HaREARem5m+KAIRzOa68Ii
YRLECknOtomQb0zqOQrVhZmol8N5QG+8zax2LY412+cJvw9ivKNOmyLCOu90I7W+
6IyNOQgD5ngw7OwsZB/ZDu1Km5b0UAVnUROYftVpQhLlVNy3kVpyroCAdxOC38zM
YQuIGzsXhHLK937o22l1AkPKfyJL/SEGjO+gcYNKpP3qBHfPZ2V/YfLO8f1JVwHa
FLZEC5ltuRmOwjMNkRhpTxsIwi/QQ3xSxcL/nglQ7n2Eql1vqDWNQzJa5OT7sCn9
5cA7m25Z/uF2LspeAD8XP5xvmD1vxXegTuJcf+QOvIXwVKAnGU3JIwNsSsmLwQbR
8iRpu75Nd3+3lR7iON/s4hMBmPVlC52xhOGX6PZLlusF6ZcbXjkLdzXl8nsD2LED
Zp1gfIU5x2ryGedJjvL2nYmaP1Q5s/N6e229NywQzIoXZZZ5+xAdPXXI5dCe6K5F
oBJuuy6Pcr1wSwYQ/iA7mF+0dM9p0JisZPt0IQKAtS94iJiTJZrAYHE4NVLgnW3+
mP7u+Y7Rf1vt537WfK4EaJ1w0201EFBM49dT9WwJCC0/m/lyoP4Zt19VsGN2imDQ
rNZISsN4hUv9cnSIw211W0LqVboIlK7vhLDPcZY0Obl+kR9OVjoNka5hYeQsZEMS
ONbp94s4uKyV7PzSP5mbl09h20prDcavI9Fvm/z/uc4Ux92kbUI4lLqHacuqCoVY
b7g/Tm01eGDyAjgvPRUhJHVZhNJdit+n5DIWoWZIuOKD66ypXXxL3Af67zdRp0R/
cgL94S0kuAyk3+VA/BziYZ0oQKC8MpS55E91OqnS/5QyKBuIFyLz1Bk9+f0Ee056
McmtF6BByuI79TG3MwlLkgZzKEhAzhZu0gY3lYmMcryxLZFCTvQOfMuzdMghM6X4
F0gZ96NQ2zud/y20rTU4gl7zDxQt7D1sIv82x56p7FzOZPPqvfk5Xl8ohPEKj2QI
Q5+SG4MY9wITNs3hvCi1T6Mj/h/CB/6ZjdGSYdp0x4hTlUZgUv6zVIPQubbAtN4a
guC09Y5hYuBwh65z6jHovzTHjNnYHXGeFJkGMP+/4uasbwB32r0f71d9ss6Pzy6O
D8nCS543NUGvFPlIUDJxkl3BMK+LOI4FqXH3iFTa0i3uj1d1bu0gZXuUvhS8t+Fx
IlApja4STyv7bDSWiv1IuORWTKSYPiIJZZ7CNHn7ppxgsItvXyU811tLNwkjl+Zw
+CY43N2pYWWWGAvxTheRBWuC7Z8FdH5Awu7DbavaR5ORsLZHC5rLzb2rYAUoHBUV
/LMg1szta6u+1H3jUmU4oYv7eNMhJS+b7CTkn4rveMgV9eI67hHG1POjCXNluSCq
l8k/7BiIzVHnS2h4tnv9J1a+TAtmoDMYQHxwETgTI4nCQ9AQzn3rC1FOYf9eRQm6
O7a0xGYAKRrhcgBW4r0XeH0cKCcSLMApYCTyJLcf1wd+ofTZNgdI1s7wEmycXktD
6egSM1OTWtjpZ2UVxHHf84bUDezGZiWuYfm3nXZpYKG7devnj8ffBAjXG4AinFap
AA8zoo6xk4Xx82knoQqh2XZRPMWZAZUkF6/unRyz3Dp2IIGGadg/NXIraqJMWlB5
wa2vU8UswLe5UOZKWN1cyN13dqdD+JCN9uqibQkyGE4EGaE3Jv+SnGFmA2spjA2s
gKoltyxYvnlaCPIg8lnOHQ==
`protect END_PROTECTED
