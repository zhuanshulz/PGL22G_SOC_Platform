`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cu0lgybbEiYKXrYDmMMGM4V8G8t3hduEf87XVftxAjlaRiwvsbzaCk069/NZ66uc
R7nneUONVblWJRIWBCgA+I7IS1UA+hVBhdc5+Qr2x+lZLWPyXx6Z0fvHY/QrAIjd
8uZNstLoS5wvpfsZjLv0ykL9AZHEhGZFN9yk5Rofn11oDWta2mP8wXXyDb/0RV2T
XvM/emPDgqdR0fOLScH2d3ZeNBlLb5mQ5lhyrB0l3IX1hJjrdwjthp/1bisiAAdq
l8djbVQTCJKYv4VBq5tRQQkSzqnnPJ4uYmVhCohfhodQoEXwCCTLqVvHz4W3ANGC
07NaPt1U5KZuituyW9yz+frl7YXexS9KFX9f50owFpbOrmWLZMYQO3Z9n/H/f76V
7NlYlZluR9C7tfIE9/5u6mzBAxbcTsNJFgz3IixYiEW4QcvCA++7S9RUquIymb0H
4diLnHtJXMWber+TwnNRzpw+u2Vl6VGs5ROYFJ0W9AwgkWOc316ANuTRL4bzvD4Q
0ShUcv2OhMMn5jLG/HcWGA9HySw191jVp/0jpyarND7AN21cpniMCAvJ6c2FFVEF
Nb6mavPybfr/8roSyC3GzO5t/zNQNFchwTkDss4D7kluWl2bwOhk01l/Hx8L/F4/
174j4GtXmpfjy+ooXM37J8ExF7XWgoeFhlGwv1DGI5YSI9Lj1hin4QiCcvvJfMaB
T3d7moev3Rd0mu5h/cAZnimpUTkHlNtIz4YaYd6y2oVe7H5hDiqMfHcYglVNBpSz
Zxw6io7SvxzhJ5Ec2Y8U0Zv9LSJpNfN/ZJLa6QgB47UMMd0IT2id5wxCaJBpr6TQ
HGnpI3EVQc4hQ7lzFrMZoKnBAyWDFV3mP452smxaz6dBqcppXFcB6iJjAPhdI2mx
4+rnZzfUi0d5/M87ZRJ+cH+L9hrzYu0HE6KMYq294i/K6DvUFuOqv+Ph5cjaRqkf
g2MLrQmjqrWy9ky3jpYEebUGXVoO72b66S0nyMI/ERjgWM7mntku6tGkXwqx0hA/
/EQvK+MC3IBgFawo+G3RGuKT3aI1GnVGKOiNancSlTbgc1iNdvj3ZDpd6wMbpTy2
4VX4BSQn/mIMdEvuRhpzj8BqhOFabybU5qts8AY3wy0UU8J84bgOGlM/u/wFFDA2
ljbNEJot1Hk8cUdS43XZnHoTQPqKrjowNy62jbphfT97QEPf/0MSgf+ngf/66klu
iSwL/SSMLceUysTm+SPo4zu2KvxK1RTZajdVTdNr0c2WLHkg//hfOAzC6o8KQaLW
BKHL4JrdhFKhMaDdFgZgOj60/yvWQRovM/XZneIbT3h2wAWq1vpLSunQFJWPq9ql
jePR0kfCs1s4qUc+DCbP4/rWb1ajyEbsyjlpy4NBCAm44RGrRg0rrjLqe/EMx+Sr
LRO/jK/Lz1ULWNS8AaX1FaN5uKEopoP7fQ1eVkUofOgcRCQUu505E9aPPnuwyGNO
J3kO6fKiJYdewvKQdDd4QzthxpeEwv4Q/gXLQNdE/VUH/vR5jNYLUtDWuAEaIiDJ
WsyCvdimdUGJAowyPMql6QnNraK+RR6b3MEfldaHszuq5ZlfRwxdVm6utwYVJkWh
DWPrDSJ40c00fYONP+5MgdFDzZcTo6TqAhZp+EV+npSnBoZXpmEGxxu0DSa5S0Mt
Pa/twnqj3jZOiN7kwvfRW3K7iLfNVmrOQjY6rVQvAJJo19+YhXmRn3neKVuKMaiS
XQ6gLyG425lBGBgsJTEiXOWMlnTQ1YqswekTKEIokblWp8k0zzYGZflQTdDlKvV0
J0yq5at53n9t+5DEmjVNM0QlWeC2xmWpcUKUAJ9KbyHIIfY+HKOQKE6gvWJkRY0m
AEIdVVvmGptK4MVkHwh90d+apZh4ENr8LJqjgzOvfbUcQxfltR9/KquWfRoEjrdX
XeCT7aCyFPwF+xf+3zcfEDY6bSedeLS2ehc7fBwgQaOenCchAz59nO+WtSqT/luO
s2hw5xgbfohJAiUZGZ7H9otlJgpc5iG6IBr5uXezzd5UL7i1zoK57mjorq6zYlc2
38U8tS2j5UrFl8JgPLJFsrLWlgiCJHNK9ZpMHD+bVur5HaJg7wDY9WKsb+oirQiF
AF8HEFtYZPfdILrnpy7nVuxTy2x5pCRIXuXG1e1IQJ60rtNZfNUUsSojeAyvqTtA
kzltQC4RNPS2OrhJO47tOksDKHzF+ZZ9sXFBzmxTIzGur8ZG00nXfhn0kk165eO3
DF5bgyKwJJLe8QTj9C+Im8OlyHh4pI1SwSqjJq0AVpH2655CkTmvB9u6ezoPcJqo
551CjuhcQ77O4JY4V28WYSNvIQB5VDBu3wk81PPtXCTvoSrISUEVJbp1XsRZj259
YryMneXuBo4pTBrwHa6MzT0oCiCjQsIqHSWQoHbyBlKiSfkYgXoQxgBC5yuZcTkI
w6C5vq1k5BImJLCshCS83iEr09g79/zQH3TDhisNIR3WFwZ3EzMiWEw1BiesgvMy
qhZ57tJME8RqWR1yB13EZkrqSaXBs5mkKsw6olcjtNep5yB3oT7UIPmU/mVI5ues
s+yF8UcgmCEU30ij2pnTPDo/dLL9vwZyg9Y7bC36mpcVu2ETrvhiAbtFskek0lOO
tpOI8CmMJ0W9tlUaiuaWqcYLQvwX8gWpcQSAU7kM6KABNRV7aoXr6GzZ0g6Ds7yR
`protect END_PROTECTED
