`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDUKvIb5xMzkGluRsZDnNv1T2t6UgpLhU3MAtixusn8gtMyREtp2tyCj/AYAubjl
/e6C8Q2ksgKYLGn228yg79KFyGO6KUAgkE1WRCSFjpq33DqVQ2VxKgfR7JfyvqlQ
M4j1hHthYrwVDQWHdUS3Dnn54fhFpZK/fgLFkfY+utKYRICDAJ3wYlsPGsjkXIk/
VvQBu2gt4/1TzvYjD0jUzK5k6vLMyKuhuyt1cVI42sThncYUfao4XsrlJkLtC27l
PHLMGUCHJzN+HGx5/IWUYszoExNONgBElcINW+NQtPgD4FFqSeAFyuJeC1chpEpo
SSEQTjxLG7BTnsDM+Rua2phb19erwr5viMu6Qg58a9RDwbsw1rooxjpT9bWvM7vE
NRjnFCjoEZMWSsPCcd+mLb1yjikfPTO3iQBoIbOO6Gnjc3132MoL4Vt6sLUE7ZnZ
v/mYHNbp+kM1VhhxAaYrX/B/JOkFw8sxSWj4D1HLswKsnHSkW+rHCxaEeQ98VrTk
SY5t11+ymz6uNo9HHfFdygRWFF6m6dE+lRX3nGQ9NTcglFS7sS7mhiD/97R5DOmA
jdhOICqht2cA/5OjweW/I7U9DBoFb6HjW2L0HnPTLCwCzLSXivMH0y9u185OfOeK
13flVDS2VP/tt8TzMIWN0ZwNWe10sxCbTj+FRlW9DwfgUlvHCyDspsgmgxuex+0p
zW+yh6UkWREYdSm/h747oICNJNrilrD3YbRvB/8G2TFnytFczHjERi5zmVTQBiWj
4Bsn9FUQPiFJjiEaQhpzc8TdMbOn0fEiS0/a1IrTmvUH0v2KJT7YZOstANnI/ImF
fQxX1hw2+0fDs+ADhRWbB+yMknZhCixvC06vd58hOnUmh0juqJNAxQxGxuJpnqLj
2Xw7AFDsX+zbFMq2LBStcB9JeX/F6udo8qzduwc53YgYsG/WPWyTvetli/UIkxne
ufM1Lf+M8PxLBXvuFt+3Uw==
`protect END_PROTECTED
