`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MiTeOA78grv2E/y87sSJ/6pL8SPKTwSVrA2EJTwrjUPOkbQWsSPdgHo+x3iLHF+y
Pi7Qcr5V8ihQ2xY1ze7o9m6+6pW4LCdZXioh51x0RDfCFmR1b5iWVirWr/h3vJB3
nITFxRk+uz7aXZteUCuL8b0Wy9ph6UVN9DIAv+ddszDtxOH61aus1N9qh8rzjzap
0gk5seZQAMdGh40Kbg/bm62M9Sn3hmukeFYFXvMlrZydcJL1HpIJh+8z/4Qp3hks
rO5PeQwmdA+4CgRWFadJRLTmzG/DYb0K3MVoxQs6NTeq7zdgFI+QButS6uEcjw4Z
JeGFG+nBZNhmvOiMDxKkHggAShzIF+UaxRQ9fpozS33gp9Lj70dfbZy+ELE2o4Oz
O0hT89TMGvs1wM4ImCnA9HHRmMwDdT+ujvXjQB5iUjfr7+3EHyuip/THADEyVs/X
Mu/BW65/EHM8bYdqm9Tm6wnFgRBv+R/Ros0god2G/f35INMgXSSaZ/bpXwSadFaz
DEH9a8AsqhUgX7ZMXA8a3jkp/87I92l7kPjWpdSvu8NSuHSS5jHTFWoSxet6ti0L
zABW9sKZkc3vy2G6T6lOeDbbXmp+mkvxzPaS5NZELQc1xVE44QJMNXnQ/+ODYXLo
Nq1IoEnVjtalIOGyThSbz0eYR4+PpZrBZiA7XAexiSLyRtHm5rSTflBxq/x2FQBQ
6wE8zYHmYBHWf0FG3fArk6ttj9xl/FXdJURwhAA9FzAvxB5UMVkr3YbQGMDYAotU
m+8VQAUArQSFB2W+Q12z50Hnq26SolNA2BWUadK7Zqri9nA2pee0X3fXVsgQ4msW
Pcz8VAlImXBlw0SUmJSM88TybukDN8+L3rtDAExr7RuHH9cNJFQuJzlOqTwLY/1F
ars+yXocXcCfPcPUkCkcmG6g2XvkSMWm4RiXYo4ttXv7GYahUbMy8P+Em2tHEF64
zOgL1pyFfcND2QtclnpBnNDPnVJxv23bufn7NRHB1tmflfZ4uQK2MHmhuFscSG6H
vMgEc1Da5qvcbbb3bW8/k7Jl2fP7v49vmTcbL2vspZ8MyMhpet0OmwkRcp7W7kNC
+VtVPsaE01QdWKB7UlO+DV+Jh2I8On1G/rqY9XceqsE=
`protect END_PROTECTED
