`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WdISZeMjrqthntj1sF9zp/W0DeQZOwvawe44z/nhbLYdHYhur4lTI8UO6Hx7oVi
ha6CsaiXH8Mv28uxgbKYf2aa6ay4RkllJ09Zq9yVJHSpCxXR8/BlSWayULFWcTPb
DB9DH9aQ+So6rRfxsRaMQl1aHcNnxveu05AujwQz+xnksyr6gWwySfgKdbT0pvXt
vGCO7fD1gpaalGnFxFf/S85kv8kKINNzUoGRIF4Kh0MCuDz00KNNCgq8pClg3e/i
b7WhRfyjUI1kIsDcQEq6NeNV1yF0FzJK5gym3HHa9FBNFDwdkEYyNHXNWpMnW/lj
YFDmkCpCNpWfPicQb7ha9jZAvN3azYIYO3g26NatpEWuJ1MHOQ3GAobNsNiV0SJH
BPQxZWRILbsHRANy3lpkSn3VpLapJWqwVbYnWfV37VLvFaktLx3miJKmbXNR/fS/
CZPlr08LaCzn3BPE3OhbZy3DX9Z2wtFup74lhBn9xtxCvp+1wzW/yHakXmxE+sPB
JnZDjMi3A1ZtdZ5xlFo+KxeYmULZjqbBv5aqljbvxfPNQH2xRNYOJ4PJIEd81tCc
y6oHFngYIyjkKF6b0Fy5bkv9uSQlIQMEKTBuWDucFPkvvib8ZW+IfS+nto6jvuyZ
VIc4s18d1TIbtAx2DovJbw/Wd0X/PnneCSNvnOaZobx+c7Ir0zXJ588PMbFdyvYl
4rTCdIMbd3N9nmkWq1LzeSxktOJ8s6RRmBwviUsDKxBwb5B0PqUPkP07Bo+PAM7t
5Ssz57I49w9na3/znyyOpFZ61VRzh/Aw5nHD+XKqK5we1WIE/AOyRKEnZ3WoTwZ7
eAdDgW1RtoetvgeqV680v4HazTlWrzt6SEFEVYHiJIqTLuwxovGpqWG4nmGDUONk
JfIqWHkkz1TtgKiFM88VFTV2LnNga06b05Ubu1idAhqRuJXA1iF31i53H4Y/vZlN
3i28UA3mtkpYz2lPqef4/LWK1W+hhsNRK2kZSwRzs7Zoc3trp4286YORDywO/8QK
H6qjOzM5mh4NLHpWDorMKTjazlP5KLeepe0pmmQEuC/auK5erQmbv8dbIjCXImnk
Bv6ARTuZRMMkF1p9mF3gfnYb/z/wpScFKFDzjFBM8wKr48AuQv/Zo6yu2cnPD90T
5c9zNztoPB+Stj+9Fy9kCri15vXqr/M1HREDtdFqEUJhAvwzV3RnyKJIHHg0TOvj
RbXpsRJ58PH8EHhiJEdms1LiNy/WJ7m/QbglcCk79Wr+NZ0ho053rHBjF/UJCX4C
jtrxfanyyR1vyyby+09inmu3NfNPMW/tPpO70SiBVlVrdiMRUg26MlW5H4W0Hjj7
hPqJ0fBALO+qxzda4lqzjc6oxrKYGmNuWcZKUJK+/LubEAaUUdiuRPuoDWUJ9AxD
84bzMQaZdz8lrpZfq0SF8z5RpMW+QpyMWEioPQDMDcw6/dwQJbim8iyi+KnzjLMK
Sb6cVYWvIUWLIUy6zC5qUISQWZuGv7pZ/gJNhAhsLkN306WKgEocUVmGLhAmmudR
he2cn1o7c7lVQB4TTfsU30zcH5hlwPJN5tHrRdgHKhhidw1wW01cgB3dgEiNoIsn
BYBasqPL88W0C5spXNdKgB5aeT+rGy//REwIAiZk5kuri25k+q4dRW5OFWUg0SZR
oJ+jlX18+WL8Lcnf2YrrxgEPvC1vrGhZtfceSjca+VT8UpIOUff0c/Wtc9BZT8RV
bryy5V3LWKPww/ASgorYbmy5ldGkwv/ZcE2pLKR09zQD5btPczLHgyxYJ/ew4ITd
h72jIWfjzaYYhx30bPSi8xOu+PkqoB0Mrx1mC9jkp22kvVB1tdYnJAPBEmOxeHkb
KLmw4H0P0jm+C7YiiLQbnMsBjNSBLiq8oqtSupr89HSiE/fppWavXNqqDLsP27eV
08bfPF4yLU+KuQlXzBb0DBYl8suwhVVGmCxJ7pWaYJSNXrCzXktFsdPrgY4Ch0Id
vsS749R5bCGylRH+vtqDJkRqUiCuBzR1pMtRNt6mLVfxrWXxY14wTLDxsrJLqYTm
je3mCG7b7foMn9+pqZ9IGYru7JgG1FkzQshDc3l7y51KpYelM1ts7GsDq8wHOHAx
UpYVNnq8/jZDnkfCmyy6q4/6RvEgpsRZbS4VItvV3OJkCa76JzQrr2aaiMq7b2dE
VMM7+PVLR+Zy0/bg1+eqBKUZc0fpJcN6aXFFkSCN32M28VjzUdD010m25IcQDn/r
q8cO/ezXnWBGpI5ICCK7tRNZkthnyLo///eLCci0E6I4Jzp1nGQkVKaZ+YmtZ9Zs
nVvvmaTcL8Hoz7kEZW0AwQahOHTJtdtOTgtH9NwQfMCqblpcCn20/YcgPPJ3mWDc
53iRFz7c48JVKSc5V4jKnofjilxSG545DohJsFPPx3Zoenvs8dB/zFlzvMlJmG6f
OeD9fbc/an7TXQHupS0nqM7UJDarmMtzOE96NXbyrhXyYYHo1fhk+ovWg2XfD+HN
LPWMdzLbkWPKOOLKvl8Ua+NaK/1tFKaKZLpPVwEHruoVqKPrGxzL03pBfTi2urc6
k9TkVT/G3VVKRwlDHnZUQRsirMbuZceMyUJMH413CdQkUiIEphlHLIV9U8y2SMz4
RKJRH4Tc5ikZpqtBI6zJ5FnTEuR6BMGqXzEOT1mVu30juU6AkeXjk+WI3zS8PCyt
v1yEHwJALntZjQGctL9FADBiv6//5gHKCkq7PcutliNAO388vPTkVMaem5QtLt1K
fRXq4BCRl7fWnM+aV48upE90d2jC9PZgElpjjEcKfsQyFYK1L6eyRwZMoczi54uM
IYAP7p6usBy3hMoLXKV51d2Xy2rvtp2UpbRq4NMSRpHQkAyBi+aC+5GIQ4v/vhI2
cILgBMHqfdwBypbWyepEDAfP/XcewtlmbMyjKet7xJYqZc9o5TB+cLc2YbqJ2d7/
7GDo6A+fUX9W8KJ+zUzxyYaa+5fK4BtlBGV7jhmY+jHDN7F3uV9pFwZrxXFur665
8GTmCuPtmR99ulUBZe8znEcB17Wb/ob4Qpu0wGedgqIgqco7w8OL9f3M5lTQCSNn
UOXO8WhdNWEG+gbPpu1fh3Te8SCKanOnfEX0kxrZXKIIm1m/26Jba0D18GrxfbwB
ScL/Qb0iBAeRMZI6Ok4NqfKTpgS8WtskvTbWnqitR1/dhe22eD7f3C3FhFNH4+JX
zjvT1oGEDmpgm4ZOBEyTR/NjoLq8RhZxgfFS+DrMDKuQMMp331OnbnuGN8jEIy4J
SjAkBm10/Ra9F6BFscjnTPbgFz06a+aLKcsfnXdG+f74+dZZA+mTeJ0BcYICsNvF
`protect END_PROTECTED
