`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiPGZpWEtqE6U7cbqbC+YCuTVZ64xwA3J9JVUh185iUCGXrSb+zlK4QfojuFHnSt
XGAEEvb7GkNn+Fc9Csdg8XMT+UXQnI/KMRwMRI/UKlVHpP1z3C1GbYCUmlCz1oV7
nm+WfAJgoUAe7/qgcOjXigohr8jeGFSovac+xyAGxbkLgo0l50dLLVk1z+M2rIFz
fK/PmZsxTnmds9KF5KnFuNpBU3nB9e2njcyUb8VguAk0TpF+/g6M1V154A2WlYut
j0q+t5la/SGHMoCnLS4xtvlEIPloBYOII2B6Gnzmbqkpqy4no4i4xl58532Nvb1A
pgHp/bHfwrrx4fJtEO0Ux7S6ol2RCXMGOBsK8j4cGifzyUYl2+E+adcdGTmHkhCb
gozZREnNQABKhZPZVBuN3hawIjHLsA7Q/t7GL6zFm1dYPGf83MuHTLgmrpBRTN8Q
CuArPWuIYcpeV4zzaoRh9tKaxF2iUywH5qF91Z5LSotHX0CMqWSVAt+n2VwzmB6h
lrsjoZ3inhCZ6EnM8qj3H4+DbXV+c7HLfypXFKXTpJXuX/YnXtRCiDn0GuOaYQRb
35gh/FWuwGzLJhxsK2g+U4hXUdicaDTZqnlMa8w0JMtBStZl5O1Wcn9TPMN88fFW
SFYu4l47jnZ4BKihNgwRJ3jsn98capYGXNfORiurP2UbwHnkgA4s+diuGyj3F4XV
WdkTQ6rAMqEzTUM15YN9q5xUehs3RlHMlLisXE6P6xG1tTZ37IX+OTcdVFCIRekt
SH01/mCh6EkbOUFQ4trFw8CFlm6gnff9yEjH1iYkMAn35/U6+5Q4nZMsGByqVmKW
j8PpbhgK/ETEGF1CW8CdW2cRQtqiBpbodQ0F2s7iNNqHkz1AQS9x8LvbcwXap1O5
Y9LOpWnZUVTKrfJzU1gc2OruaWpyXwetL8K6ixXUJc2RLUtqPDa7SZnQCbM9Oe8i
ZEWdgll8iynjVIX/z/Ty/8REaZxUl3d4SxjsIj2/cxy7mC+Tsi3mmtKAwQYMGVVE
f026w+LHgU8itnl6gD5Stl51ZUbLoYMRxNPkxw9je6LYd3vIwoV98xTykGWN5gn/
p9F6k2vFj515tTXaIRFuF3lRmh5BcszmMqYF/qG+HRW25CagHF2HrHXxiWCIO44I
ckNr3k9xpOCs+lCjZwaKr3RE3M4JKtoWkb986an9H7eggzl4zoT2kogZGHckUVU+
j3Urt/oLXPd1zGvMN8LZFHsqInY0mjlKyyivWtMg1XO0CPeYbyRU3Du2sYzgGs7j
vZd3Wt9TotwsFZoWnujz3zHFLIuESi9Lbt+ToUjRNXeLen6KFDM1i2UZKPvbrK+2
D6+q2oE5snITQvcUQADbxxjXsV/hHZTS/IMSzTzCZrI84atLMDK4IyY8NP/BdpV8
TvkH8SsQK+a+GDHseilUJQ7hQ0JnXNXabzaR9oly6cdqDHoTIQcnrgMBUCiMrR28
Kquh0L3DxFluPGgm973zDXuAoMG2d3bbdB9KA4RwJH3rf2vbnaP/TDX1eIDH3NIN
Ue9dIZYmb6+M1aHtW9nKsCqLmHBF0iiMkEQUg3gm7Kg2bhhSvxuMycX+I8WiPGLh
MaM+HEQKm3IOn0P2oocBL4BpwlK+JgQfDTuH3e5+aia0OJBYUz0VDAoRKJiqyQwr
cHdHSC+CGkffy/LFpp5eQuMOn13OgEVEHCAG1GJOtWukmLLcRaxFLxI7r5OTDiSn
gIHkVv/zUIzsEHDlrFyFIAyoAYnTairmh5ko3ww/Sy4tKG8KzvrPdZvorjjl6D6S
UOQFR8EMf4tdhE8uHlDmE/ERt+gfh3wqXZwwyprO50X9+dY8vekxmSfb8mq70h55
MBmfajiat5xjn/8iRAuMuNxtvOzJGdQTNvw7Y9gjzOg4kJQwaX4G2gv1HMx0oypK
GfzeI22CD/aTbP7UXDQcFnIfGf/faW9jCOgK6BJUrJ4Z998q7jWecN9Eux5GYUpc
`protect END_PROTECTED
