`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qwxnhHtCWeyPuIxN9BBjIun0CJw1XzqSq2XukqcXyGM+hYmAd45Xju3v1hiZrRIQ
+oWan1K9Y/ylhX6/7kZhT+aenIsHIKzi1iYt1HuUIttVbzOApbzEhJAhVh0v5hd9
5mmRrnTosj2eJ18CIlNjHbhV2pzClvSRnPK5+cdRYAXptx39SjN/3M9fONlcvFtE
kKZzOWMRwO+CRaaPV1txRu+ubG/SsY0fHTOm7VbjNf57UAIM2OfkKbIUWF86+q1k
JF9HNEfOhE5RPxAxkyYVa+eDT3jr9ej3obAAtvs65kHUYmA0FVd+U4wsJC2nhyBB
FXoSm/vXhgDd6VZHlIrIN1YbDX8ZkJ5cSKCYUE7jjk1bPLwFPB8mOKB7l9Hc90Ps
04QyT/wuGdLFBn/SZMXvP2s8DoK5Baa1bc6oz17yCxDJgjo2DhdCFU1tXCLBcNPt
aavJFX0TT/UqP+y6PIA9BsXSzlNJggu44SbeN0049pOxlt7C9hoxjnuJqqoB3dqk
0LppVDjwuvaXYtc9ow4/Gecj1Ak4dTE/NEXOPSjdTcxJgXfxEOfM3yXveC0gXZo7
2tkomwlJTHKbCG0i5s8Fdw==
`protect END_PROTECTED
