`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uNYjyX1LTuSxrqlQHuDHpumJEBranMx4Yfiy5FfrZDZEQKOPa18keTwjOsnAP0m
fKoyJz1xflOFHeRi/9EKNb7rVjJTjzDGJjWtHHME3mI5+Fedkh3nboZGwwyewzZv
q9Shfu2ZcHY2CbTbCo8FXJB6VoHpPGFw05mx7rsEj/AREwdwGb42F1h4pnv39Bse
2Qg8598nA+PvBMgwSP9XyrTu2WyIG6JXLv175I6+0vzvFhwhnB4rWNz64wCi7JZh
K/CuHH6c7HsSvlsZvuH5hMQFLB8Wfn5787OXmN1OYUHfJQxVQzaDcs3GqHoB3skQ
lRql4Q2x9H3Zz3WmK3ZqrmNdl57ALqZdkbmm8A9K3lRBppE28QOpVOPyR48X+AUN
xxA2EJWOgFHEAZCZ9CU5DWwtYwqk8vGCinrF4MGL+NC5lm3zvNYKZ+20pgkD2kmq
0IjpD2kvrAmcc3OwI51rkvOU1ouH/W+h2JR09GjgP6zElhzSwALJoLUGp08Q2Rgq
8hNtD0KQx8KOLqZwsmZS1w==
`protect END_PROTECTED
