`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xmeDrcAvmYt216UQLCR6tv8KsnsC7iAr5OKGZoDnv19hlL9azb0QkEI5YEM3AAxF
GKELNa8XYUB/nmO0sZTraEUzYFH02+lPvr2nL5HMtN6s0SXqLBykSdXedxaL8EjG
irY1Aezf6rLQZsITdiOHawvA6sWYw0P7d58EVjGDS9jEyvaf6PkUTXss/TCkN44u
5sGdLyBgrBZwGNZuVo+/E6jGlaXFcQhikIRxGiFw+1tc5b/f9ClWYPlZWLLQqG89
bHNetNpWyV5sa15jALouxUDMWGi+BnLgGFp/KO0cRIvfoVG7l8kVKOtiLaV9ZaaT
6DucDqwF9zAP8efNHqoVWV7PfwaEKl3q25LH1VOZf5auSUItbwlehrRP5CDchAU6
qirZ/uAXGt7DXQh+y5OLs1aaRc+tTK4rYW0TOhVMC+1G3rlKXpXEu+5lpWm86jjd
gRVLcDNjKMg9WpjGdb5TmPRd0EcK6Y3j76osz9+jsx3glQDuaPrckGoqq2QVeqSX
t09qrWAiFzbuNEyCdI9NXQkj8FLB0vXvSDroM+dFLA7iI2xUAVMffxssOsIuVdnI
BfBU/tOyTMa6XqbyhrfhdSDbdBEOytsfcRxpKohj4DSwf0zC4J+qLFbntW1h6Nni
udfyjXyFGUAbZwCPXQiwWtuUlX2qEmk5B2cuUoy1hFg5JNWy8zjAmOW6xTZC7c66
uUk1ifL+U1j74Zd4MMCw2TQB7SgL6Fsl+IQIu+LHb3ioo/S33f6rZWhy5WJPxg+s
uxCJDEdATS9aHv/oiPDql6Rn3uizsDcDjWtuPgEKQglKrPFemXdan3+jTJ3ruBf5
3/q6MM4sqGvg60fUxySuKZ/Gf7EmWN2ERLInfqfEFwjORUu2cseG3elRrSuBk0ZI
`protect END_PROTECTED
