`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzO2sn3apmcaApCQLHe4OmQVydvvPXUpJ6zg4Rwdcz8BGoE1n9GI4X8o9k0eoxWS
G54zeuQBSFZNG4MWLqXOgR5QEtow0ZgEqEP5TjlJ9vLevzY43i87q0UV/zYSyuH4
OYFUCP55P0+xOnEGtTQybY/3/JoKbO7Qw3onOOgRoXMj6dUo5ydTKuyzkqhzQ2JM
sumzydCsH7VU0nFuhg6zVvIs1wOq6mHxsuvMNUFemRlYUFGgN/QEmuzu2XeYelQn
fZapzP6mLqQjhSc2rSjwPFs7ao+iAtBvGtcT4G59MjWxoGgiPgvTThBOzp8r0lYB
nybMttUU8yFj+eJKxE+8Qwil7rhlzQhr1JbKaQ1P5YiipuaqFcHzTJlT2eZGaGgX
406FOSTmR/QY4SX9xB2aiXVv899l2APgKlOhD0oV3HLPulsB9+EEN0JP1sd6Qli1
rj6xTG7gGwTzTUjCnnuV0R9WGmbUbOrlQ9XgZvaQ9FaZNfwExU43ou/tY7UuudEg
9/2VKRPJIrcgaRAnLBx1TLzZUap1603KHc+zeou+pVJrfHRNfvIs90cT/BAgYa5S
C9qXd7Vna6qDPhOP9dhUEEdxfrKNI+dfnyBCC1bxmzHtWagRiTckPinBpWMB7TyV
+n+AwTjDZzpPWfT2GtUGH3QQ96kMG//YzRiIhvtKYh2vlRALMV+BhcSb056Lqc72
ZPWNOt+JN8TSdnF55liuT7gj5ZIQ7Gtamg7aFFP13DQL7tcL28btH5L2b3/XqlDX
AXSj/uYaTCfmdtGq0X+VAko0sWEMfD22oo3dPB9SavNw4UlrMiIEd9F8bkxE+qT1
hM/QjHPfDgvcKn7leEvtn2Bm/dHPm3mulgCN9B1YGSd1EWxu0stk4LvBIRihtNoM
EmDe8AstIvp3sc8AwwMMWJLpMzZlGM6SznXkagPjnYd2Jh13o1PncdBTATY3Qroj
nfIcyovWMh5DDWM82OrtRAO+AaO4Q7EDcF1FnPNlmSeuD74NoBBYvOlS8oNzOCtk
WXle+NqG9+gXNnlkMdxjaC17/ROtoI8Z0U+3tN9oU0wAVlgRc09lMKSb2ZyLFcuz
3Fir721Uje09IefTBs+jP+2IUUF46gcn6xEnR2HY7h++2JIJW8TLxuHyYqjzrCir
cCM3qG1cnDrNNhOG3h4850ZP1MpQFbc26RBl6hul4F17ICrI4fQ/6HhL04ovZjcQ
Lq9UWRzC8RK3u9Fm1xXVYN/TapCnpkRGjnh7RrY2VB2QNq0LL8ldLEiuzeZlvXBI
7IUbisGs8gIDIvoMI9I5MXUw3tDtjHcbmOWEs5lYX75tzuuPEOzSBjrXrWsmvllF
UieLcCxr4vkJhUpJ69M1N3B1AyukPRplaRs7QLBi07Uau4w8zAKQ4Bt/sYHzH6qB
/LlZGMCmzGmz2kRXuaWdbw8Zp3qAOPV71wx3+zMVLcX1UDYxCG6Sqq8t1aEOZGfD
u63IIj4Kp46fcG3EZj1YdZ50mC1dFrmh50g289zYhrUK7tcWS1UP6Wci0PGP/DJp
+XrtwSAn3grguy12FQzTDMoNC1pd7BZCWlmYuQ5NDvHGO3vh3MRGK+QeR19/6XmW
tTZocmEiDONVCmICd5iqv8t1g4tkauCmU+FvrYNOGEiPeSvuAJhR6EaGylkdS2Dv
gjeiiIRDEstFRyGUK/bMeQ9dDS9HzmUCW+eC1mwatONoBJ1/6Q8wQbQRzdrYSSZR
nVzj9cTCq5JdcyPKO97a7b4fx3jvpYhIqCPAdZffUD1gtrzKAVtEqgztOnwPt7Pw
y1M+9kzT2r25Z5ofYraSWSq0VuxfkEdkdIVA5uXPs0zkAIbJXXq5o1vYljZJBluu
wRiCkYsfXGpWB5EZoWHlyup4NAwyGdxXyHmQXIDzRwSLnwY6TlemKdBfQuH/slep
w3A31qnPvqT9qk5zofJu43BWdri4BSZIv6a9uEGD0Y8FWTKhKS+fWC439SlwCfi9
lxC986LV4BxAR98nSAdr6U2sHeH5u/zh2vymfVhhZG44Ge0aGpIpyo0QsYYGvcAC
StFQILIIlM/VWo0uteDIZKoU0vUbdAJc6YevD48C1oLR5ZMgf5ErUQwkbXeUcZz8
I0ynl6WzV5p2Z3wMba8p0RYJzW63VPTLL261atuCejpopSADvHXGp1lVDVg+pDu4
fYTZcRplv2XhmS7DqvTQ6mf6LYnmu9FsdlzTK98ZB3SAFjEe73+9ZuVJh8TjZGi7
ltfa/f9wiIdMO6V5ZQ/+G0faLvMwEV0+bmBsip20tJ1DfdmYNyUs4PDOX2FIkzmR
csiCjP5DMc2FN3fXzefqDImKqo9/ggTKnzYBplSUWOgu/pXK0Dj0atYqGjF5Xub3
A24Yl/qDmUDbNbafa3QU5EFAyOvJcxtFJEQBduRAjnts40T66jajqPNAEdlCKjYh
qqzsgDvYaV8ff5oQNyAFXpyIha1B1W4rO4rbgIv9V8GDM1ZgGcuUro3JsSEhDeIW
2J+y7Ab1QK0QurP/03S0QaAzfYx/TUr3MNmraMJ18MdER1K9h9XIGRhWZL9eQ+FH
e7R4gNXCE1SNxusMZJ+MkoQMQIZnY2wDBF6VtmIOyjodlJ5dqYWJ9a34j/Rgc66d
4L6omcnqmpTZwla+O9uknHJVTtxwIZpPipj2df6e8Z7JSDqiPJWPZQqBW6vl2v7w
V+mi0gbHTEIBz/+oK1XoOpI92ih/MBJBJAWoUerwMiVnEjXb5y8MDYL1OCTAeTBa
n6xs84wmKs6gVhNN5EhtMrAIQ/jbCYvdK3WNbqQEP24lnbCJOuVykJse8yPCzP6Y
l/XViK9U2hdjjp6jpfZ7rNRlodwN9c6KH8BKfUVfi6m+p+cuK6hkoznTx3dCAfx0
//JRqFYuAUFywX8uTgYn/4fsghFmRID932wcQKQBa+jIa9NPqqHmzPvy54e+DQjD
xp46fbMnPw1i1e8M+EpdC3CoaKqN07Uk7+eagW3TNq/GRGa7rCwgt07ZNYq542Nt
wZGdI4eh2otr9Pf5c5QDxkhSLS/E1Umup0IW81GesKNUO62CvFmpTcBT5EsfXv8u
rduKQE2q/vZ6z/jfz4JeFr6f70IY8Z7PJ6JM4+jk6x2AtJs8wk+2Osr8FmJgrthX
l8y5VsgLlicttmYH/rVl01NAZ/vWWTf/4k+DasBCQZkoAl8tQ8M7Bg3FZpnE4ICn
wek1lO88o7XUiE6Zz82xPE8K5uOsSLHY98is46v57O19jDgMDCQs4FDQ6j0xNmAT
QDzH3gzsSKxIvWk1VwbChzrP0ilipP1ZwTUfzdRhJDUMD9XhGsDGtN3//IqBE8XD
O1oIB8JAaEnsfp7Mpi6l8rmT8zqmNFsh8Zx9wDNqIjxT6bIcUORU+4cXaWOU4nQF
PxRYEnYXaj8e05Rm+6TWRRoainNVHZPdeJau9y+dTII89K7004zLwoTZ7UnOHNcf
E0J90awSrH3gpKF5yoQ4sc8xL52LddoZ6ThaQTKZwXkYhG6Or7QQp0cNk49UPRBW
NCi2Qvf09Q6vlHkgwUiDi0oh3k5cRg2pvd4v8ny5xgEgcyXVkiXxaudcYQufuxoR
QIe4oWdDFKavvAkdciG9X6z/4GtQrU8Bbh9nnWsymdUav3RK8n3iYEnKKFf/3A4i
MhpWgrAAzvAaImcUc2bB6Q1aKAtJ2t/TzuwXA8Ip1tCuIx7FeMeOyhoxRsU0wTvV
EVOwnkdsDGbvpJSAGQsISJfGzIzkzKMCloYHprcSuiBfUHzgo/iA8JeQpxJHoLWc
pCPnrlXjqFjhLX8y6W8ry3d4BaueeZB/OpX4wd6dvMD/mGWKY0z5Vkm2rotgPsW7
PBL2VsQQgfOurzx8lVGroZtqqE9SiQ3wOykv2LfY7fLTcjZQncxLcC87t9oFvOAl
eknCHAhnYrCK8w6J+Spmk0DJN3qUdbLJMNAE/JTTw4c=
`protect END_PROTECTED
