`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDjeBUy4SXW+0mK6KZ3XIzjH/vi/9iFEq9h0xdD3/9ospJw8M1uxy/P3e7KvSAO2
D0XQP1zGBkdZWWgJE59CRCgtmk+tiY18zzE6dLqtKEfShLfnfURDYOjwZnvGDM4+
r31a1z1VxAPivueEsROdp90imuGDJsgiWxwBGVt3h/tZJzg4VG3awzRlF8t8LyZM
OUAZxI5o7zPxIphoe1swj7FPKWEfcTJj0pf76OkZ9vF1LJvipcVicfsz5cVOIweX
/H+rkiAcLI/3dtAVNlBdpMdHXCU9gAjx6KFk/26/z2z2hmkvcqb8KAQiGvH6BNlD
zfLEfznyTV3N0DuEj1MWyFy27c2RoGV+nr50hqXmcZb6HVvlarCb7RBF+039Qe0J
7+881c2QsStanlp//sW2BJu2myPdKf50RMXx3gqoTycpDakSO7xAKDTGR6te7Rmj
2tZ0KV510sU7ySN0A7jyYkDwWZAu7nWrATDdTc5iuARW60/Hbq1TTn5desgDUoig
lPlGXLKLN636470v09PtCds20KTYSAqysi7fajatZVyiMYA50ejzMhyMYF4Jiiic
ueku8IpCY8WyVg6ASB++xxXQzwL3hD1fOjzjYGO+FS2PIO5ekkrVX5ec1RtOWqpV
+0C33WLW2EAWdzCCGQupgTfIa5LgFZfe5kWUZy/avG0CutYZnLCj4ZDQ7XTGTQjK
Bz8QGlYgK45G3JLtnfWp4Q==
`protect END_PROTECTED
