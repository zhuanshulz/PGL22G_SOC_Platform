`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H+pnFZsS61DvLeMqHyB4XWD1JSxMtj9WGrVzEgAjOlqAd5LwkYIwjV61eQD88Aax
vKsfgRuchabU6bOs4khQyzKZjY4+iVTAsV5j+YEkAat5RG37T9i+U+zfnuRz/noX
YnDx0tWZqkoQq0tkBi0X5L7chZiLGVvETX2cTRJCxFw76XUoBONObSQPjg/7gWak
YDl1/bEjZzhWSG0nVStVJCFZ7YX8CUM/DE8N5ljkoreJwvFN4CD2209XXbMaQXeZ
odNxsY6gCJ7WFvj/cPPy0McJFDwb9gqYeUpmGM+oMAO5p6n4vCXUJUL5qJXj8Q1r
LeV24bc/kehHWyEPq1wP10wYs6ZQrWa1dtjES+qj32W4Jlipl9+X/PQUVpDPB9ZN
1DT+EjkrFhMZguFctbCA3HsHx4uBiXlROo9vMavCSLx1eZftNWxV3VeiABAEKUvm
wLeZVES0Mg4lhDGMH5btzJonwa0hhCFJ1RqXvWm8ERNebK9Ph1CwxRFk0yZW8sKg
FJ6C9yHLFd1BYF5I0xVKkYFE294a3pSDBa6/7klnf5iYw7HpaMarZ3T/70Um0dLE
xWQer9rRc9ogNqFQ15pXrbOD5hD9J6bMFroUoLCrWrfU6R0LEBIWYAnwYniJRh4y
JoRs5mamyx9L6kgtCSG8y8AdzatdH9Ic9mIHV0TDWa3QemRwDajbWUh75te7N1GI
z9wyRyeqeSRw7tFXPbiq+ZvORQTYVoQ6m82Qu8Vw91Db2Ki4Yd7ykItYyrEJ/dVw
UtnG+rbhCX5NEI1xo4U+fsGVj7puZzKMmXokpzcu5kCwSqB158NTviS5pKfg1IWg
ZijujerBfbFElCg8iz+qqPRR3GC/vsPJ8+Rf0YK43t/0JPsPRKazWhUO3Josi2do
2Dnk5XZ0bRSqVwoL5+56aEKccZzHv3WcPTzhBkUY+idhaq2ViN6QKSTWwIoAOE2D
Bv6wP8NRjXTMaWUlo2yj+pRj6EjkCEnqtDOU6LJdExD028zvavz+jnhaiSiXGq3n
8pq7XRsLLKq1rOCba5Wou5h01c4VltIMM3Jcxumwz2MGgX6nsezjKFPheXeShN5p
IMica2/TT5tnOrPsVRTob9L1M/2hP+YmHuTtRfWx+xxCk4IId4i/y2dV9Xurs0o4
AZf7sl/cQozn3f545fs68+JKFH2ZD/fCFCoWnlT8xHgCJ/R3RSTuDOhSxCryti5D
2v+DRN8ZUSXEgrwYnegDot5RlYrpUiT5f3Wm+yJyK/par3zFD78LV/s1P696GO9M
9HvVGfDdgs5TX52evADJALt2tgC4b0J98a8aE7AfA+evvXr9DMqF4NKW7l7+bck4
Mwp19groe7+W/Cel438rO6nHrP1EiZNB4jvlRF1a+UTgsYvftqyOQgl/2BLkDjx8
pBCYrIlKkhKpqHU+UALum49Qyvd7xFmdJjfBQSFBYFntB68nLsPTEi7mem4YCHNh
kNsYix7bzeNGjfIBf1cy2ji7yGEuoSsrmgvtpmXkCS06TGd3UwVT/GNwrnzRcy73
LKc+61b6p7nYxcXfEMyE+UkOcCKInU3K3kHn1IDj/dR4gaESG2Wwv3+SNJNzGZmy
dftADEhI2VBO8kjnWXBMNUMu9pMv8Z5kwW8lgSAqlDYkRnLi0VMcCq9FkHtkylPv
4Ymb91h0VLo5S5VMFCcJ5I0MLj86fSFGxSIBT5V/SOg=
`protect END_PROTECTED
