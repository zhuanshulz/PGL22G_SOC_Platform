`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tv7DXOToGYmIhIUcKpcOCKAVO3TKIP5Y9D9ert50Oh1wCU3HKvlrVAOSdpcnLPBW
GyK3G2PWj9XbhJvDsv2QiBBcYBaS+GIvM/rLR22fVlciskjhHjLB8ZCpUXnhyarZ
gewZyID04Q/JOWiNrga2AVxGlMowdSZNpeyNBHKkiu3CLBHbe22KIFnB7vkvqrCy
ABGYpxwCYowCmH2GFyClrZ703UsTR7w+FCkxjmDTF8FhRmQHuNqXCS7f28VGSo8l
JaI7S8trDMfFShqohbbUbeX+uLaPLNvumVwaFjYCpYgphR0YsXDfG2Q2cm8ljeDb
RYBJp7ai8RWKo6wBNe/g81SzDwtT8PDt2AWvzxulRTje4SdDXo9+jW4MWA94s3am
YztLazivZXOzASDQc8apoebShgYP0kEHm6R8yFMcnd1PgniR6wy7I3KAlerdM/ZY
`protect END_PROTECTED
