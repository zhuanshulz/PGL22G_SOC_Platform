`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUb4Z5xJ1Ju5n1Jwz095U60fgqgV+mP/InW2gcjFo8PGq4LbQlVa5+kQ7lVVSupQ
a2ZYIVt+C7XJeArl8OZ1KXIBucMjpOepDKTuVNO0c2puiVBO5mLQnVddcb0/AX9S
2BRrZzWSHn+zJsB9isR0ZLKmI+M6KTggDNd5MDSp3OMG8Qv/ca6hz4Np4poTvW1G
YNG+Gx4r7Av0LC2bRjEIXVModkVuXWV7sKjkhpZfbKCej2nMJ6bvlJRCqi9s6mp/
E9EN35XLNl1hIGUTFZGalF0D99+o1seSSjslHsnqMh0zJuIS8C2d80KFLsQoUYly
iY1vSN6Bl+1oLjAfrQ+Lro09qjREB+rqghfWVT8hrxH00VIDXObvl5HWlEtl+nwL
bgnHGaDLyPKYmzkwdjCZYTZlhBqf4O/CIJErhHBqwuc7JpX2DpoWrsejE4bYQIGH
HyBFQiKIl/SN+H+tVJXzQg==
`protect END_PROTECTED
