`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZ30MSF5bvEsb+gbcVLBl6/2TD4fUeL0l6KsZzUJzc7DRLhm0L9RQ6x7ZKMBFnpx
iF0hnyiuPY5mylwwA9NzcnGGgeUBYDG8M9HmP3zHA8hH6w0ADwI1S0OqVlIoC/qx
peVUcoOpGP0yRoXHomZNNSHrySYxDmQDCAhwcwfG+5fEXR5mF2RT5XscFWnF2kur
RcjDjGS4JoIKdTxINVJa4MKp5Hh0Gc86IjZXU7V8jypjszt2gjVGwPfMe/qUKXc2
bAR/SeXw2EVwnupxJhrvobsthCFoYEzR7Sqgng+XhfAnd2jtf1n1JIrrzKCC9A5I
NRjHDTlqUHoHPFpPqCpWzDcl754SwIusR4cvfRG3CEet9pAltrTKJYH26vtccOlw
fU1iLv4+3uN0wqk0QOGjB0tfS4rQgQ2vwAhfwmpTyO7JbiM1ahAJ5+ETfQLuS51o
/d+3e1Le8UBPAOfsneTsZXKUW5FeU3IQIyyfBJSD5FnTqKZy2vasKdNdaL7L7xM7
mQy8qvkd0glpmyIyOqjHKjNg+LbfMMoD6IKe0PwuVANdp1QwQtFtrw1xSOy0Uqdy
rAZgkeE8PrmC88CYnumEn7T3mUfUoMG16n9Kh0tHj1Py2N3BCW+SYdF3XGkK6o8N
MeKiKVX1Vh85Thbv8IAqyIr7JrmgjIa2ZYlIfdXcD+qNYTK4VuGSvW0Xv7IfVJt9
VqcP6PEuahXrRjkQ+X1/IpgmOoMuFEs0Lvvueupc4rofvuhZ2JY5VhuEmN/H1YZO
J9jYuNE3RjQd9SV/J7tm3Mq3KU8LKEMMX9ZNCZK2HU2ZOyVFy3R6G0tVvPkN1W1t
CNadrRnOQExyN6odfAd9Xqg+E9P2ncLhv0893/UPc9lwwpXH71RpiZ7xRpJFFRBX
OAtcA6LuKEpQx/Snbtz8EbcKd2TymlLtRqxyT9XfaVMBe6H3X+qTPzgWwrES8xZx
akeNZ38HjBYpj8Axhdl8qkxgy15q+cBIktgnofXMpdUbZG9bXyZnfwXgQ0rUIaO9
mifNGUeTX80iSkpbzaYKmoYtKnG7wtIIScw2RU4+tG+GrOpfhrwH7uzuTOI1KN8g
u+atpMBMp+jlYTmZ48/C3hFj2gbM+9WqR0mp0Nghy3CLCQNmuJaXXa5qomiIphxm
vajgxfeobCvopdKVxPIUm2YlaK/SNKDCbNOF9oKp5s0KPGFf1nOkv017l7Wy4oMe
IfVSjXsUpVKeYDQp/gB9xVGM6vM0F1evb+wdOd1HV5uMHbn+GgWUKMVhq34BS9lY
p7sdnRwpColCXcxmtKsGSdllYrm3MzzfcaUR3c3ZaiZJbxsk1bBTU3K25omiwgHm
rOWvRX/5cHa9vUOFDwJpnhI7GEsyAZYRYheWKxivuTsgKJ8r0X7SYM6LktbFo3Oh
2kN+S6E+amsZds+eUbws0/8hThi8xlM8rLtxpPGUjYRYl7rESg2J2PlNm+izXLvv
DD8i9AgmRBzrT29cuWqjqzGH1JT7m3Ju4tLHA8cfZPbicHxXok0OXgIk7pamavwP
779BuSnbjvMiIVMOffM0aoW6xLlXw7sHOX77eUZTzKSYcvT+soNAkZ7BiPIUdwF3
iK+xsywiPtssU4ycQG85P0a8Z8HbEETZb94afjHXmkTlqcWdas+ubKtEE6EVZZw1
MXuiSSbOcBG1QdCTsQC+zYi3L8PMRhV4CpE2/4fUzmeGEFRT8bOz/P5Vy/aP+NhT
PuYnLn3G3DjtLjHFevfptnYUomCzMMx4EpLv9UotwdUZYrJ1Ne+pxuEBlAA/qXOr
K3blpQ9gZ4biVzFr2JWBcbaxgskzk2IEBTIGhOgSMTuvELwz/G1JABfEhXEOpUl4
g2SZrRoipDzb+hPKe32gViNdPqrZ7XFkQV/9h6HIw3PLPLEf03wbTz2vT/mf6Ajb
OGWkYL0hD1UhNmJHUAFzAjiL2OO481y2DR0YaVL1uZuFI4zgC6h24S4G+I7FwM1g
6Pv9uls9rLoMfGYjzO6Wl0Rluu5UPeKPqsEFAQqB585LfPCw8g9MiBoT8Hi2i+8P
zP8jA1ytLsY06Q8cXe/rJDfo8oZhiH4XWI/0PHeNC4iI6trgdJBi8vdT4gDV9D25
asAzTX9ug5+vPJmXYcbW+aoHhpi2std/ZmQTVoM3oFNVRfgVGn6BS66RLznfZ5UN
jpr5Pwqrrqn6ZtPvngIJXcMsy6mDxIHlQPHyMq1f/lXObe30AQS1d77WzeuAKElA
03hIjsDHHSxpipR02wKPSGsSGKtxOWvUdAmQOOzXEZJZuaJT0/iS2088v5C/Ahm8
rocOQM1a7yqEJJX48ruVQRNwCWgCGqWCX+xYfPXlPwXxKthZM2NqR/ZmNX874qyl
sdToJCsv0c/Vxo/NEfgQQzQPiMO6tM6I8Ib+oE+a9gqnovPDFLKpmetVHfEJmQ3E
+13rMmcPRCoKqwsNEKgrFoiqNKMLoP/BlC4Li3In45J5TMrtje5Mz6nVDcG8F0/h
0SZUY0w4ELEX1JD97HpqqRqVXgy2QPZisNajPhBm82XzXVXd/0mPRRtYeuDjQC/S
ARNEZjmIZWyaeBLTuGj+KYsj0eXJtwfljgnKLnHB00HGfB8X7uHy+t+AAzfaeRVd
aoLAyY9eAD+IGs9hLelinuSfZWJPD0E3R0P2Dad/fSCuUnuMk8zn/eJwEz3C4UbV
KBNVtJSMp9OsqSi8CSYbg/CDPOJuyRh0ey3K5yTiwSNCAmhGq3g+vjx5ntG2P8Fv
U4HB0DxUCFc8QqEpB81VpHbJYL3dPBcz2qoXxVMShVeIX4hojaO4WPPvlYI0IWX3
2L4HExhA5IKUfEr9a6gZu3cnT5YUXX5MS7gj+XYtYYwIWrlQ7ov78+JsYO5TzqWj
ziDnFEesV+3R1uY17Wv0z6b6vO/GeA9JM3+EEsKP2spYpYozBJ6tltXzD35aSotD
/M9mKtJavNGuzmpmLwWSGL6GWCT/IzwlN5yFAYbX04qdHfBiF61DfXWhdks1OJch
QppM+UcrVOccS40a8cq5ATPLwDXMtkJK4bW04+i6hRpnieJ16kRo3C0zJcr7ZMgz
NimsS8IgyRPW/wnkFBRnMA61is+/uPz5xNucUwfQTYsqUyhGNTTELGvH+ZUOIjal
bJiH+b3BC+u8j1ajHfyU4qFRnyIWoucBBdB5paJ0kFUGs/2SW7fAXDwqPt+Z89K1
OZqo2adP40nCECiDNf6XcMwBlnXqbWMyWn+TqW4yb7q+8MT/2AAEQlRBcSGDxQjT
CpjsqBl7CYzXSkha19dmm4U22Doj1fkOFj9Hk/5z7NNVuMkmm8LwD3DVvDmgtEC8
tDJ+MFMBzBMoWE5cGcVPfwDQ0CUBEk6sOMsVG6MggL5eV7oi2bayORKUkC6xvaM4
69Hknrq8ab6QqgcluoVjxT9xLqKm6/llHhg6N8oR4Llu/ZaY986bUdkOb/hDJ8ty
gRE4t/DeCvtiwYF0ONtg1UVEYL/q/P7kdfZzZfjUs/p3SY74wPvpd4onVuvJrpe0
GuC7yXI1NlDiRTfLtgvW7rvLILYIgSh7AZKeRBhFCWn+yFFzXMBvHRTvSllAHk36
Oxx3aYcgZb23YlK5E9oRrd1OKUQj9R1vR76DjNhisCRlEAUJri0RQaoaquhWHlmd
rdao2F5+rjoiAZL9lmj0uaorHsVIWTnKBcog6gPzaaE36zwJrNrRGPkcYgnTIprr
WdciKcK7uVWnWTcLFeIt819cOAgs6h1BtLbqFSQECGZx5GtuxiiOR9C1YWIsX18p
tESyqV3XYH/+Vn69NpQe5KIoiM9XlmqotOehqoEvgNFaE8igkDni0DjX4izl9oIy
6zES8uo54cKDHqaif9eWaRGCBbnjcYu5NT8wCSoMmhmZEpIZ/O5u8I10HaYT5IhZ
/E/5RqlqoJjkFisKpitVBUdADIeloIFgVIKwHX2SBMaitPCGQ9vil+uTuL4uS2NG
HRQovRaz4p0779ggxMGLFiQIz4IkKT7qj6VUwf1YQDmlNOqPMoLAgD7jIXYL+A9r
uxExiPK5zvXIPNQyYp00t04m+ke5SUfxvZ3HvzrDR4UDA1m8CQ9PH+AkUpo8YRz8
yrs/zXfo45Y4poT2xlN2S5gfO1HIN3PXWZeAIG75gs8dfBFClHx23TWIUHrqH0KS
YhsRokP1Aj8Gj+ctuhOk+ZfRnk+HlbiPV8eV0xc/eajNpRhh1D2OVgnaYQS9DPS2
p2uUk5sij2WsFvjFQY0N1D5O2diiww1HS63s/aXn/pu+cJM0gom325aaAaJM5kIu
GPX21TGh0TWUaWFg9rPoyhaHaGAOfOEoEDAzWgR4qIkXreJ1oBGAO9nToHdTe8vu
fcPMlgKIYNyb1VSLCvg18/wNuFsUbePcY7PX9J/gLRZKtqOVtPMsMjE2CrmqAX8D
4NbUdiH76dFjHPSCA3VqQ02LjLQBoMtx4lkTANDNwBU5BS/zThk7usFPFr9MCiWu
/cGJaS91eMj83n+4FwVxLAaBrlS+yy2STWZnFE4gsluhdcAO28iYvgoDGkeXuSJD
fThzlLWAI/qNDnFV8588WaLv6a5NjZJZ41oz5OwQrceVwoyJ/L16nUUjwlCC3h9z
lEhV1L78u5ENiDOf0lH4kjqWis337mtziNZXj0XOYWQnrsVYJkTNU/bSFnLXkZ4d
ZlxOI2/ICf0jwZ+e3sakZ7glpEm7bhJTmRF6BZEErBJmcv8V+vUPwp4AFjyGWmJi
BYkR6eN+IItBlVd9kWF0oAy16o2zpuDQr4NyKjm4qCHkp1KRvJHqqYHGb+f9ez15
4d+8tzlH1PwvMOHkq46GGolMfkl8bhnQpKNh+xG+QZlOofVcp2ix4L4CY7AOuJL3
YMd3obw2rKlJ+bQr37FUzkZtHEX8JqbEbS7O/ga1cMncvUidnqfam94jAB04JZ1W
XdHanog0QXYxnW+iZ2hpogpBjq84xnp78zIm7zzFwLqJAaKNLm8ta5QmaHVW7ZMO
8C2U+joogotlIi8cXqqMtNEOf8exlWrGjSkQGgcLG0cQJbSXY3ipCpCOw8JaYgDS
knVVf5wj4cKX60aED8NeysBSQsK5Hzw2byY+WNbTSdyMjB2i8NQTMeAQwDbffVyF
N2ght1H1gXp5AuDMSkXHEDbq1a8lwHGwyhS09IHGu2vRIgTENCL0hywjNUcqT77J
9N3aNkJc7uMoNJoZCT36JGm1TFBIgxhc9+p9eoCLJ0yLRYUjBajL5K8QoclUtL9i
dqKFmPhhh/4GSlWelu8CRWMTXKNhrD0c2nnH+KYr9kFi+N8q8HS6m5Kl19smINtg
yNxVucbnshbeztcXtzcEoCQEtNJmy1M0UwHLj8hH/6IhXcm2XGMFup0C3hAUT56D
l61FZ0WLtm2ElXpSQ9jqpBujiiz9eeNtIlTZg2Bgv/EJSN6Avi+jrDR4q7oc8mGE
6IrcVCbbyWAYzACsbKe/8hZjWZ15X3MMW8mSyKL1iVFUZIhh3X6yGttcBDIhCja4
5N5IVJoOjYm7Fz4IYfVvA6tjLUFUIjEQKgjm44MOHTzOyp/RwcSqfDZ355uJXZr0
Vv4RX61KOdWA+etHf7qUOCsP+wWSykfNlqjMUhMquLAq5xCD2cVoMe4a2BLu0Vsb
2txMpnyAbzI7wGLqmedw0qTearaXvRCFBmDema+veDClWwDE9RPbWDQO/H7COQQI
o5G5CbXYwM7QFv8PTsPQPV51kLC0OEU9Ve7ko7ZW2mEigs/hUbZ4IUq2YA44yOKI
Mw8UrUGlZLnMyYJYgbSt1d9sWFFRyYiN2WK4iUYFNd3FcwnB1I2Jn3gxXMOpwmds
EK02+jlb7u/duKDcKP0SbaTL1NQHSyNAkW32rkwFPORhONhjklfc70uxjBTmc3vX
xsy4qEb4HVljp1bEsfvWiGwscNDReYv+8TYDblrpk8Oj1Eeeom2MVB+ywwNsTAvV
t5jEwohAE8+vnevB8rFaG8FaJTqy6B1855irrRvwtZeaIjQbx6m//E+k3UcQ61WA
SnoGNzEWARR/3a02q1zENxstIfmnfCFYb5c6Q0zHDSiOF+AM+tPPFgGptoMFMZ0j
AaqFIfMAy2ujZb/jF9ZuicC+bvpPSvj0AmxB7W0w4bTvpC9kxn2e7nqALAUr9G4Z
HlENWGG3H519EVkiUfELeaOZDseoTxvD6iweRvT2sqBXzYcyhkRUq8hxKN3irLfi
gWZUrvACnsqcsSe+Iob6goph7qbHcoWejS1XHTQ1IgBQpci9zBJHYxIe3H1zfYoS
aPKcRLJu5pD0ebYeLYN/7x7WvoLmZ/F4z8VCLhGfBvJapJEP8K2vE2dUraHs/hpE
LVeXyMGzUGWOnStVrgJAgJHgz4R3r+mKeMkssRrohDhBTWLKzJXEWHNyspWDnZVj
UScSyWt+GdKOBjjJonkge/1e+8Grzb7cYaeDN3cH6SjXqDHE5+BkJji6iSXfmFqE
dcrJRra9C9+vxpEMOTSg6I09gHwXwnWwVSmrGcZ3Bol5jyC3Yt1UZLABrls7G2la
43K37UBJEQ29GrjD+AkSv7fd6Ur2llaHG2CW7yEnofGf8GQFCZj+LCHQV47/nL71
qENK3MAqKSoobgEJ4WOBsP03Noiqcg4pjtPKpOsHn2q86CUg52n343dHkIPqgz7B
72K84m/u71nFWRCId7RdY9n+Cxcc630Xbm2s9ZaCk9NMYnCWs/UXcKWoMy5KgFfp
WWqApEKoDnJri7UgzXAIfqLnKy370AJUeMO/rf2oskKk2lHjvmFiMrIhGi2ile5G
qcT65WCsaGcsqHHYOJWDKjBVEkPFG1du1EjYX3XUhIOaaW68oQU11J99G/VnThYT
QIkIfFa2Tlkpj/Rd0Xn4BV0DrfNvpntLFEo35KgcEMFw90VQnhQGR+c5YtKiPqwF
guSdtrv/jQyShb82HaQoNkiWvRl7gAg5jsamjQLMUczghVoP05RkM9iRbUtnIrYO
yRaqIX11YMzpcB3HqxJq/RFue/JJroOfrmyZgYJLtuVhUp4yc2eXb/11KGVqAtQC
HiTJiIpLkqjC2h4Hvgjexp4QEHo+hIuqkLp6pADeja0=
`protect END_PROTECTED
