`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4QxxBIFH4FTlsIs6tR8I/yVU8EsmLBjUJmsEW+XDMlRGmqqgKh4hf0NPE2b5Ops
F11UbmOM5rMogGbSgnDiwo6XBLKuVyP574tYgOLcSfbFp/In/t2pmiET2UR27y3Q
4cdsFd5NC4q5H2F0N2NSqo0A35MDg7u4ASGrxAFa0bPTjj1bhSsM+865W5/D8Cns
tnGCER6QSP8Q1wxRCHzGBO0jKqSfteweJG/893t2KQvHc+i3O03/bFECW5BQF17p
9wE3Ftx2zEiUWysGhIn9JqUpu9wqS1WS9pFIHKC6elCJeQbWflLGnrGqDSJWBx90
AOHcYXFgjgzjz0cYQaU2OVzcB82BJAktXaTbByZEdXFi+dOqw0xFPxk6F367XTKK
+Z1/gMQYMMtkXlBlkdZs9uRzOtJ6RjnsEC1EsC+qCkLI0aY3+tezj6tuTAlMpAgT
IAuTekQ1zjxTtEiYuesxw+/I5Y3L2c4QIhcKzeyNTKOS3ElW5EQ7WpxZgZS/Ljy/
PM11X2Y5iXHCi++OktumAN0zyzbmDBu3LRGB4xmEUzChT0+fA2fkuGLISVFwCBkW
HWGKrloLL2BKiZCU7Ks0L8R6LaEZyXt5Dz6zHRcU1ihvWhEjfhwvS87YhypEEgQW
A+CuXuPoLywll4DXPNCD1rqtD5dst810s/LvnlGEFbN5jnkskbJzJjjxGzv3Y6dq
pgK7XW/vjDcvE3WLwfIRZE6XU+nLJgkFvc58k/jpVFzh9xIEuSQYlkU5ZX37ciwE
vk4YG/2wxyMkU9qdkTIVHRWb6Sj6KFWu9moEFFGhF4hCBhLSWolraRVmeLVH2U60
Mk/WhTX4vQMzX0URYgFcZ2pG7+CAmf+iLiX8D+KJo55Cv1TV21Vx5lqyDsajD/6q
Tse2KR/7OJKriXq9LSX+my9EGv7K3p8I76e38n19odTBxBnrJe3crb5EvCby4UiZ
plkDY99RbcXunFfjjJOks60CxNCUQ56DSc9me2Qw3PY8DS7vEqnwzYnxLLyGfLDj
XsWmyPKNCSgv3A4p6dMEjdR9ET3aibXzu2Bzz1S68LrP3BlVytLVwpy/aOwBQQQ4
LQbexDW9U6Xpg0yWdvA82bLVrG73JozwIOEHWFUyxCflk5FeuqRIaUNGj3dP+eKJ
O7QRJ9D72xtQaGVCcVjOpjGla1XIoEsO0fUtD51jn5Cf2fYqi61d2KqmYsBAW9r5
FMa2gou/ciKy75NqRc/9ur4BKlkCZBiWzIdz1dCCu1KDGYDrJu91NYPUoDBUjMib
NCOHHgXjou+4MNI1IL+ed3UAj7NUQ8ZBv64SlW7VsmQIFTXivSFtjkmM2k92NNYU
+LKHmvQTz4JIRjcUMtlGr1UyonU02VehBQNYditFDKrh7hgtpCni7TX4JU6teuBI
2ZYe6LsLJq7Na23rTZQ/lMiRnXJfUhP+JwoIZd9gaD41kMDo3SveG08b15VWw4Iq
Xxnr7ciI5rtUtkz2668SaZtN9gMvLSW2is1Dq3ETz5OYN4uHJmEKptnifCoDbmoc
ZvFPedZd+Wh9JuEuUGkCZ6L8n2xfj+jeT7ogeSJvWpmQUX20/uqmuFUUMv8tFZwj
GohOJgHpKnab/hQlnxctlpDGLRof9xheu1omxUledqMKxHPOJEfipwOb8pho3JCZ
x5Ev9eO5vpPdKPM4YKRJPsWd1EU7JeoNtZxtbKRUos10U7sDTBAJ5OuioyEBlwrf
Dpy3r9A+q8SHqoZMx/PsaxLiHmxoNNIN+fcZU/4nQQ8V2QvvVkmdXb3PFnB7rYlS
TakRYiwgjk/QuHJvYAcaVg5v7Kd4MQlwLXw048+N7J3lo7khEJGuiQcDRTIt9RU7
NnPt+ktg6NnKvPJihLTcGN5FH5x9ydP4ROs4PIzK5do3XpyT+Ph1O/xzqRcnNmLi
ew45wC5PKo9NlgUFWHpJk+mpoW2v7mNiWkQO9qdUvao2zOeGMQE5UmzXmbGtCtWv
7NFZFUgcXP7x5WHAYJV1FdFLQ1zHDW8QDcNeBrRowqgiIy5AHrsHF37An4yJGpIP
D5+dhikh7OikiOqr+RZeKV04pllLY+IdEOEfGUtbDG6kn3sJ3crw+QiRQmGY79Hy
v50HajLzXW+ni3jZFNG1x3azVLsa7Xn6QbcFIWiBizjXRvAebFEyz0+ixVTE6Iar
MvAehLAd+v19TNvnwl79IZA0rrvGmfuu8mywmYuC2D1KxhHJPQmqJIsNbT4AsLms
YtXq4e4z+3YELniaeY6EB6ihZAhEpbzcd4uTFSToiaq8Ee0uDMV74EMkfg2up6dO
psa5qXFFRflUOlxq/fPTarDce0HO9e9n0q3Ca5XDU9oTdBZmQvm5pZoFRCzdiJL1
DVSv55Km7kUGOxGtOk2oNGyD7Uh+hwpxXznz8cdNIXP/hYsXbMMLhn79wzBBkggA
qcs19Yp7YlkXw1+iF0Y4sH9qejQ3FoNhdoTApwTc6F05AH+p2LNL9D+fGaXn07Sq
CUr+kbxORzQwjOprIX2StIi52Iz+zHFSp9BLuCawECA=
`protect END_PROTECTED
