`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGDo572LcbsWcswW1W2s8gJaoRqk1NN2NcV18fFCQIvOCuznO1W4gZAfILeLNZXk
JMJYZvgoJfU8gDQR1r+FFJPx/IRO9lG7BaCuo2Jzei82xXfDc2QLdZidrprj79+P
C4LGLtcDeddC6Zbxr9wxXsv9SevLuNa/m+bH3IXuEQI5t7dZGbs7bAc605hDzkzo
9tJH+INmJX8OdtpUzslHbg9hjvbqFMSoDltb70dZ8OEN91aJaz4YbMtHl9CEQLWb
ljwue2IucPIFTBDUJeU2HSvfScu4a8kidUKWqRzfNP0ywQgMrIuJpU2x0qHeEkSm
j80w0/R0Gf3PD02UeJmSYEl+UvLAzJ/YHDOv6N8utVmoXdjHCsRx5lOnGdB7Nu9J
VjMwW0ij5hnvFwWHCUCpMK0wpD2dxflrSdZxM0zNEpdLhhhpyYc/GRFoTCFhxGQI
KsggxuIJPbkRObmVqqFuGZq0ggjaPDG2EpaVALL0+xoDzfHk0KYZzVlOqG/7Hyab
TRpz5XcDrBnRc16J1l4Lcmh/3+NCU4TOiC8a8krQdKmPsqzP1/+tNZ8VeMkYL2IE
EiJPFvH8new/wDYNR6BOspoXu8gY0yrZRjrLeBzzUBs51mlD/Rk0Me/Y8a64jQ7f
L4qogryVA7spEUATbnMHk4C8gO3iCm2Qh6If8IOM4yx1/pGpRrLD6bM1PfInjKJv
sCYdwUrzt1x+7w4lHKI9ifsvftERXQfexW+/xy18iH/y7Y4Qsg0fK7qP7t4rVWha
gmeCNZTb12Fl+y81VzsuZyL1awLLQ7fvFcXw9Mpj9v9KHf6qrErClE/beMNorsf3
IstUZv6AZjhAIb9MPZvpueK1yVNb75pD10Ds7IAWGORcJX5PDY/sk7bya51gikM9
WJK2Eb08IBrp9pqPNEzq5uG4UmXFHNaFsX46G5cVd5xtsL6vRSh+Xp6Cdk6JOQ1p
z9m1jcB+OpwhSGKFA/BQUmsahB/5bZbeVY4w+Jh3jZEGbGQSfwXZggkLQNO2JuKi
4YqJDcDI2mFoIFWCzQs3iL27eYMK96Bp9oy+GJTWF4LiGkn+f1dI6s1jFWztZyob
EGMm3m4/VnwXzxxihb9+A4QWXsKup2DYbI+aG3G4MRXHz3HmmaKVRmzl7x3aZTy4
Bu687s1hJgEU6pXk+JsJE+/E0fXpzH4qtUtUb0PSkQ2HEk/65TGduDpCsqeOB1OD
XWDuvs37eyoz335ZiS//QxciCUKlogFs92VQzi2gKOlk4xKdRQoij2wRvruzNqyV
vLIxkoN9E01eOmm9k6UXqiG51ItIhbDp401PgVoSQL8rZN82vAmWpNjMPDYPZ7Cm
DMat1j+67/zZaDGA0OOzlpLV9suhrw1mxOc6E86NnxC/zBnwcrI3rK9w/XzFQlnc
BJ3uBgPlmEHuniXsfFoUyMButIume6mHcFplNU6/BZB1lTXxWNTUFjNEjgYM8Vod
K4TcmPPyOM7COXblGsOvNeYaavNohavURvYU3K7l1IXa2JWgJprqaGJrlq6FxCkY
FFCd94OTSVAP6e3QTBPnxXfFfx8LVJ0tvTviN2EOaewb6FqnzJZ1PLEbqDy+KHJ6
2HCaXtIi0Mf8e1aUE5DeC/xepmEG33eHPh72REqD26r3/BiWx9sUYRI5G5sq7Rta
Kf8FekOYJhhKhE0hUMNlI5po46brNMC129YGGjPfR7wy/gfKx5MGx+t0xsk1bKWA
8XaqY8qgYgkt0ajNLcbgSHO2UgsdtjiQWMhf6QijowNPd6WIN73OInx0xyQP3qX5
GaAK8qj/5hy5c/ID587CXA==
`protect END_PROTECTED
