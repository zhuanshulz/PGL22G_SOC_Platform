`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M1sbXWms41q7NP2YHlarW0N9Uj7ACqLwxUfqDZOmiJuboRBp1j/A6tqJabLh8Ffn
qCG8w5CELyXqv1+ozxiO/Ca4vcn6uHzqksemDQ9o15NdONpq1z1Cbu/TGujM2Ygm
E9ypTLo6q6cHbMAFxD9gbh9c0g46zB2itZoqlag0hzJWRmmy/yYvniFeumu7IeLK
qjiTU4DVWEAkS4iiCgmMr70prOZO7tEATSrsOqL1MNJ6jioSzNUKzw6qAehexwA0
xqhgBjFZ9EbrFgqx4KMRRaPZqgMQPt5GckkcCdKTo7kaXhEW1fQngcZgNssR2hS7
dW5xfs0aFrz3JuHePVodVc23JvAfYPycZ6u85KVyF/obSzlCE5WVufTGOyGo/zz9
Dg7wxNjUSlj1QkncEFIDhuvHMcIAeWJ61zxmnsxZD0M=
`protect END_PROTECTED
