`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9wesSpAn///mGNAz3duGg9D/kmMHN0DKWBUJH5IMM5S2DV0hZyGbuFAQgbRt/gMl
5pGRPS2uwh+9O8r/W8xQak31kUx+jc4dJ6G24KcfUQ1Hbe/ovsAnixvv+Q3NZsKO
IXlZUiwPdQgVza3A1+HZ/wcKxxlYbrC1NfTAGwoL7rZBu5x+WcCJZdgFdechTVEv
XUKNdgxZKIOajcE1+YkLrrLZi/FTuA52V5SbElJpqk1eFPzYtm9fIdmDsHhUHmqs
gRTeA8/lC7qnPFl1fCjFPT55HK+XEOxrcdwmgprc3BtMbQY0MgoT7i5PIoW/fA5h
32xZAyOHZlieLeLECD0Xv0MzhJPDUjZomqKPxjaG0PDYfZ5AE2lSEn9lVFELbJ+f
V+axyd8z1a5Z+BCVnOAhGCSUu/gnlD2BxdX72z9ZMH8pqOWXLnSbjtaXfbDHZgyp
6OfIyTKZsUELt31Po4LFwLC+cfUu8CWMb+IFTIVHmzAJp2R9dwKq8uUUCDa686Uv
H/3GEYvAJZx1irQPzXRf/WXBLfd60798gM88DXFVZ6v165lSYDwRABQhJE/MVtlB
PolM1uzcXYfQ9Y1pzz2weacLtQQHr8ZFmdKkcGGU1FpjGTo5ROVI6GAsm4iEWS1T
`protect END_PROTECTED
