`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uh0g/VemREUQukvATL9PJNopko9JAB6e7hsOy7Xa89gd9WvlLRpdLgr88wCfsrtm
sapPPr/pTRstHF0ckNCLLfvZaeEKzyiqCJmgA65R8KgFM+tFJGkvGIUm532TM7Rp
828NeqOYn29LTg0Ela5LjmcTr5NXFWtic/YDssl8U6c9Uomjzt7vJHWe5E8KyI10
MZfjEXVsq3if3JmusVZQSqtPG4g9MguPxWBmkCQK+WuvioV3EexpS92vjKjiaDf1
xXaA6slNP5npCvdnXH+HSOcNs1YTB5LK7SYI+HJWkDTWTM9++PjEjVv4kQCI+Dvo
8pnnpRvGpoJgBTKOzHRtru662P0776BwosXcP57BTWrmkhtpzD3X1yDspxbzyYJW
aGnTJatQ5ITtaW5HLq+zOiIzoie0vwG+Kj0KI8ERP4SVMg5cyA0SW51OAt2Dpu4+
ARkrzpuw4fQf1gP4UsA+PcmCN8f8PfwiODBUpT8wIQ6s4OVuYFA8UkVbeXVbOCVO
iH7q7uXXVDJVg8UCPAGeXFjUXHgvRIpCNHEvkSjlxA5AtbM7j0JqCXCDG39vTcR9
JVt2gKb4QjIbxdhpt03alw8fK+l21ZL+4XrfDCoSUwMdkKKXPHXPiIqpntE0zVKl
X9Lt86fyl5t8NmkztDiiigG5h5brkQgUkPevtaplAWLnNwl0mWVH5Kq46uL2xc8F
QguP9YcDo91S36yO0C9NU51PDioK5tRKP1lTwmIcYevBVnypB9XXVrze1yaHbyJp
24dsLDAhFvN8FBouDBQnkw==
`protect END_PROTECTED
