`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J32qoNy4ALT2auhT1Lvi0jYhH2k1hLnpVx72NKLAync7I5hkv+BzTiiBC7XvDFLq
32CpADwrCLkWTy4fyRgAUPyGX3ADnAMNkHk2+8x9jF8p5Uh0L85FpCYrZ3+2Mosq
4J9htscdKAzh8htDjrY0nxD6+MFkyPIS72irvJH4MLXj+IA7P30JmfiSxfjoU5sX
vhNF338SufjvPHgjayS3zLwLPhbBpJ80fHBYh0X45SDkWkNBU6P52RRlS4KqCaOf
cdaJmPPtKyhNe/Cici9Jm0GPjoe+kD6roTfHf53vNnHWE6cDvKwhYg2UIdqzk0hA
ZEC7Zx2TamMczUwjUePFJ4lFdTIcmlfUv0oud3iuaNnpwsihFOsGIxaCnIUJtG9c
KJEhliM1nlgg2W5OU/VuNg==
`protect END_PROTECTED
