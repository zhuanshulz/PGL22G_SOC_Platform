`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6l/jezwjnsu0v4KKUJBslPu8/C6xWfcTm47PCe/63Ao9u2xWme+W6W9CvW5P+DM
a8iOVo7nndMz3kkJvio+oweR+LrSTh3YKKcf1IcuqMsCp3tsTDqi+lj3rKI5iypu
DU6/cXSxX3cSzvVq9ji4g2oNDFA3NPnNuf6BL5UTPl+QXRcdYIJZ7A0P72Vz+DGE
CzOahbQok+dsDGrD1NgdLW2Gafdl/p251dZPxXOxfjFJq8K3pvp0EjUf+XEvbc5e
qm3Qtb9azdFKKnuuZWHYkF6Mm/EnIU1uJCX+pWo+puhQPoTFVTkCChqGvBu8xppX
GeuSGp/YacTwWSfIB4lPR5TShO5ebKt8W/ucI0kaJ22suWn3rivs4lBhw+XguEHs
r/abQJhJAWa3lHxdDXOPxVKfksvjWA4RDwxyl6g5q8z9JB7x0DveIeCJBy+mAqgH
beI33GKPJYILcHsPfSf1sHhqua4p1E31nIox119ZZXzt3RvH0Vhfh1JGThSzpqvE
oN8MwBaaV1eSZLHyFjsjAPC2ynN+zVzUQtRIln72XA23LheZdpH+sT0vmVX3FDN3
PU3+kaO0y08PqZuhP9LRskJQQxf32Mg/VRN30s8bh2gpGj+ZprpPY52ezGRCr1KS
oBDHua3EwEvBXkMLKKFksnyRicE6K/M+MgK5QuGlgWBwxyIOFSdMFFZpMHF7F8A6
3xxOhtMMu75Bjrq356umam7iPcLYq/P1E1IjYx+XM8TEMVAvHPZ6j52sJm4NZmyL
xQpbEiyJ4A2pGFJbh5YKTl42Q+fQvClbZDVEodacGTXqt8/V2NJ79mBuj+dJAC7l
eaPcKqTYZtT1NWnYdPcejHVm+S45MQtX/k2jMA/VX8M57ZkYFVKZz096ho0mY9ez
adhMsuPQ3FamIn86SfAjEgr2oF4d65iLLa5yk8cuGBpeuMjqwC50BcZX9Cu2OmdG
PjiMtubB6r60u/mKBWWegYBXJPdBtiAZNPu6yKCw9ytWCkD2K6YE/GKR/FD3HO5d
OVXo/mZuXSSpvFslGQQv2eNKcDLkiYTBYGxuxs6kZ0qMipmKcMbvUBHuRb52d2Lf
28AZEzNam3X5Fvd/hWATCjddRg3r87wWxT2sIqvMsu6Y53MQwj4h/sRQCwB7biMQ
qc2Y3gMCXc1ZjfToZ61Q/wOZnCLtE3VjhXYJDoW0tUfK3Rywl5Jc8+V54edHBr1Y
/G5Pxmz9za3h5f6nEWwUzfIhlfmZgv3uHaTJvaKRRqfAkap+pkR/FydFvPIkTXso
SHnMdKNdTn6kylKO3SIHSh3kUhjNuV5s8ASDQG3QiEnDMPHzSaOnMKcNHxP9wsU8
sDk2pSESD2F9RUmUhslMr5PYVTfYBxkz4O9ez499faZY2vdTt7xBs38MFfliiqCi
64/XghBhx5RyKxezdW9ooTDQi3iwt1FOhQLFIeN/UxUJIhzmwnm5N9z1wRGeAogE
AohEiB6LW6Ndi7n9WatCdOFI0n7DByKvq6oon3vCncIta3T6oKgT5NUfBjDfYk96
khqNGtU9ihkjdzYXE3f0r/b5UPj34ikD5d84TnjaM8rZnNQk/c9huZpN+kxUFwjD
7jYXc8Pa++APw1TgDAnJXVrqVnETLoYhyXO0ZbNm2JcDfmt0ppWUQxAupjAUBNGk
ZT5tZifCDogBrw/eVY8N8kBZHvxFj//TOam0gO7qdku3y6MXZhtbUdxnoWhmyptp
tzjEGMYkrUKF2YZ6dVbjJXYA+r0YIqk6h8X7SQkFD6j8m/dCF7EcH3pltkakyYpX
1KqqqygbdLA765W3IUQ4pLeECBr66yGoXsWSMgxcupWogFq6Kd31eoKWv3kPEJ2V
CN9ci8utXyhNOw9gCbVCVml3tFxEgml6nO126dI1LkwBtQjycmtqNw44XJ+svE+3
u6gzUamiHzTh6MqSj3WMWpbeXssvvA9REPOiuIsdE85uGY3LvcmBOEoTLvZubaGG
eNvnntv7a40EOD2XJYc2XXkn9mgnumiqYT10Uajj46NiuT0uh3xuyrIwFyRgc/4g
cWttWwB/PGpSJZtA/IsTNft17+G5puFFK3HkR6Zog148ok53S3dry83xjKxtLsQQ
JaLykLQacdXWSDYCtgXEmGj+WPS5iNJN5Zp5A86mjRrJEnyTH1qt+C+ptYHy5J6C
q8yOMuBdZrcP9bpaS96c5RBO85E6Rx5urzdASB9t3qyftG4uKBGnRcyC3STUNRys
oPybVDzFUcS2Yzq6R3LfhVOpxJ8nKUYKaqmxu1sPYw7FiDLnM341nDuEtafAe/a0
DF3y9H4Vb85t159EJR7N1mLErKXM3bdGY9rCMKpd6AoB2BMB8Ux8VpECaX8UYuQ7
`protect END_PROTECTED
