`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BeXj5SZZhO7eIHCuCgvUCGfoox5FVggc7WH+QXnVQfX5pHBAIfVB3ZmDHfv/qNtB
AoOxE4PN5fNdVmRGg02Sp26pT9SOGGb+Q7TQYEDhNx71KxRUSAi0590+cHFmXJED
6AdvMB+CQO/eZVNeoTM56Cl3hbVKPMUoibNQMY33VJmAC8D0YWeDro7N2Vi07smh
cxZVgZY7KXYjUZfLCWXagVQHRDCoCuYJJc25QEKtuj6J1zy/5Ymet+aHMaRc/vh/
AeHRqdETuilBv4b+f36pCF7PU9cos2aTabXe3FEgfGr8V0cg5rPfhRRvZ/DkVn4E
DmOqCPMvj/eTGflhOL1JWCTLcumOqdgNPm60niTJDNcnJ5bFfyqR8UMnwJFrSqyb
kVnkbShDI1S4/sAejKFfjr5GyY7rTxZwxZgs2IDnoE+zEIdRr3W3e1DmboYdYme8
w1Z0c+FiAJNYPCbXP+DE/krb5JvjTv0DxZNS7QVGbt1XG0K3Z5SFuKwzwahLUPXu
Iq410HLESC++aLczAjX8EW+nv84q37YiVXSl5MhZW2j+pNLl0PAsJsGYg+cUXaw6
e7uRqag58wN9gZ3KXu1ARgz0Xn0zQ9sodSPiCa+Xnp1FyS1avmDb8GMhkd6tP/AK
mfRzEN7martnDyeUhgeB64rqX+HkPnc6f5USlrQSuaU10beOkjlRWDA9Td3alcY1
RdkXRfoGwmVY7A/m+RYKcEaHI/ICCiHvsUmwmDpVrncmtG5moeJ2bmIdziJ6jAUH
hMhK0fjjJsfimAHFxWzxlcrayzEZMtdNc0g6zWn4p7265OOeLBmbHKGnrZG4mvot
6ffEZ60UPqech/op37biWEHKkmpjY/wXRgjT+BLO9yo=
`protect END_PROTECTED
