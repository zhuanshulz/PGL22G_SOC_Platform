`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I5DtGOvauuU0OiYVfXomGWhfdvnFLp84YUYBk/Rdqtoycru8c+NXoSPN2OPcaJdb
3fNUHtClZGiyEyJOci0skYEKbQOjivdfWgVT+Fe0M98EfgBp0Wcz7kLDvus0S/zY
fDrm5NiQs8ChXy1Qe6I9uYcad8JJhxSa//loHMJUTQ+60GcYqir0nXPyaL9n0dfN
ee1ntfVrzMp5HHl/hmRH+I1u6I7Wa8EgfPQtVrBtN6uGcEuBLZfoqHuSjZhJN/FB
z+yN6nMF2Vl/NJVe8pWKT5RzPRn5pMaomF4PJ7M2wT79XOPIDCVyLxyJklQKqSpe
2HkIsV0xKygkoBR8XwG73Erx3rd7Zslzi3A9/FSRmQkm4oGqmOkMC+aooqSTzja7
1a7G5wvVTY9MqK5s5RiwoLWtrYkzOFHSGXgyhK7EvxknEmTPAoL1p8GJskPt48ks
BJ8qUUqKBPMc7PShLFqa2c6QAzpzoUtFNPaKH5X6owg/DZLyzzZ2DVaJQ31uoS2A
hbHdMOTxBfEj8cSsBsi8UIwjmDfrGN8fWLw+AP+XGQg=
`protect END_PROTECTED
