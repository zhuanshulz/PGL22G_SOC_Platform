`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/gy55x7Sjv8s73Y6BuH4ENqKCeZWe1iSl0xRcs3QDdaByjNkU/fnZ5cS4YIIbNk
gC93N4bCSSK7PhmQ95WMjAEVQ3G3TJVsUvP/Egohfq2c9gnpSOmTdd9RNBAE+5QT
JNcSdz5FGv2Dn4UnO0dDTQVkuRIo1j6hfsyNUuD+iCkuziMwaxcowhrQatwkPkmk
zUHnt473ns0IK635L1pRQz2nG0OCu5ml5rkSogVOQA0aBZl80yyHLMQeD5YNEXdW
nO8BJOUgPB+VPV3tKTMXUL1rbkav9N+RvE2Ts2nAeryYkGjHnYrBnvKBdiRNUfqN
6GUazwVFfZGlDVzvabrCQ3cqgSh7d3yAvey9OBzqSYCuqG9jComZtiI+wfbe7/JF
YJVwV/lf5o1BbLiicancS0TM37ZTLOuKtOub2fwcW2k+p2UGylbp3vOjG7Bc8kpo
VtMHH/F8cdgn5mSm8AgKmgIw6iyVFqHwtYF5dFiQAIqiJvQ9vy7kyFfj4eBrI44D
gG1sAHjYDbsIeYizrPjeB6YHoDb0v4804kaJKjw9CarrKwoyETu3cW2hKdj1bCNI
Qo36qFjQqzZX7mACsig2bgKbRUJd4WH0Ab7TJxZXCJXJ9+R00K/JPKKhb4b6ZUN8
T0mKg5KPdXV7A9nU2FvFARXmHSox87aLV6zxZMZrRTzM2FWhLlTGgp2Jd43vYckc
I9nRknufZHn36wQlkWMleQ8DoRV1KDDAVxXx0Wzo0t8z1XHvA/ANyVnmqPy/ks9m
aoXUPT5alqaq3VIHnelU6/0vo/OxQdEgXqaIlN5GOAFFOY2D46kdiFyjm3kHPNjD
rUpmkpbZGEauet9+RwbyuV9u7boS3iXlx3OYCC/VYx+GewzPB+8pZxgIM+8QY1aS
qfvOpiQlo2aB++PNHRHQ1EEHNpv0wksB+hKTELuTN9wU2rVJZAPrnixJ81iButhZ
GqcU+sT17lW4zdSfv2XEjIKD/Ki9T0qnOB/O77RRXS41+ongUdXs9pvC157vTpTW
1MqNHYejwtDRB/Ad8E+efwkiogFRmH1yhHo3gyXCI4weKj0rzcHPDkczh25Aw3DM
JAxYOwqwbx4QYVILy83Yt3wU7Hzq69QI3aTUIhduP1ggogare8LcJGnNtsgF4aL2
U6GW8g7q3Cg8ctd+WVd7tdFFF3COcgiy5kXRN45IdWwfLiMhYWA5+J/ewRejULwQ
jvAi7xIi7iOtDK/0yjJW4R3kxgcLhwwbxDheVYSSKo2A8X4EDkaPk4cMciz32dyU
Pb2YgE+bu5PkS6xtt+pU/EvI2h6VYTlwDGz+LLIvckJ0ZDJnU12HRdIVqVJjuMIw
YxMK7HYYJM9WTkcxz0NHVYJAwXg9x7czVUULLxrskEJIrhC6eTFLLtRxM19RDw0D
y5O4gs+2ecaKicnLVXKG/NfawYIp20dL3Ociemp7K3FDvVyOWstglD070qXeWGDw
pghL58264g/jEEXG0N5uLaW0EMJquPaFOYn0W+iTIq47PlIPS5KsUIPt67dAoAwS
jv+JNSjKZEKuWsfeLV44oBMgB08KQXzNfjuJ5y42fcyPD5dekjiWuZPqbtVWei6Q
pHpb4pqJ1cg8OHqVBTPEm4LNiuKY9HxR+AQKcEBhhulZW5Uk+7tUglHmTkwJmpC6
EjxwsmCypj27aIKPR9aG66TQMrrN4KIQLKhfv7txh7MeAYK1TbVCL1/LZ+8BUApS
aYyi/a2Q59UTeDAdcxDL+IPtVaJa8OI563jiN/tBUvrzv6EM6Q0mnnFDx1iP7nIH
Mo4xBU6R7pQkEnbgQSu70xaqWwHJnd1M4JODeadi9mkWSVUMgSl8dD3z2iRtj91j
SgRPfjEbMkvM4ge5Ihg5V4nLXnjfeTbaQ+LI2q0UrQoe9YcnUwMHUXgS8MKC980S
rR+SduaryFBaxCtrND92veffu5mabKqxRyOmykR7Nu2Ohj7K6dfGSUckyfCUcLoy
bKG1aL9J3ByoYKgsbqYHVrKy/wCDTPghhojPj0H1BKKt8hKXY4EXymWtcCMysIuU
w6e3oFKCweFkVFxaEAJO4KvY94Ik+4SkL3bT6dwL6toDhTScjbdoRGvYoEFE7wbF
MfoDn0uRUFQCfYPo/12NSfC9B9v3u3uJYl9udMtW9Oct+2W9HnT6bS7iICd93+CH
BoRDQNBJxNjdTTWVXsgsBKyQpYVq3qslVN6FuAHmwxW8+UOY74DtwFTKxw26KXX9
NzpuVs1MS/jAazgQDHQkxZ/pc9ubiOTwSIZ8LXbICeTM3r7+AzmhbS3icL63yqMj
3H5dV6H5aujoOfpiLcv8nBlbKyg6NhyLAM7Hx6IKasxIohypx/9UcSH2S9TFzKlk
XgZINTvbqS8hAYokH3AV8qVA92JgMpmb5YYDceabZbN7JiPEJdgoxDZBv3WIJPWv
/T8eEUlmzAtv2Qo0Vp7WS8Enuu/D5PVtCvmk8XX4FLbiguJJbR4RMfAEIlNthSvI
FCKffLjNB3bjqMD3XHWE/jNlO0YDOzDnKaZLeARP1r2UMaFZAek2nDE+1IX9UkUy
9rHfw5oEMqwT/UuQgytG7oV/t+LzxA7sOuiLMF9QNs+vmQvNS20gANrqCzbrbkve
nkds6yPVlME6BYMZmZ9LNZZaZIozvI3BEweH6TBo5RRVLoWOKwO+M0k14AZ4udsM
LWVqHcIeWhlpsGGmh/CbQYSpkyGPOPvveZUx1ByIjZQb7/B/pzvq9YvZL8ngfsZl
coqpuaScib/V+7yJ7SHVJn8KkC9T+yNqsvsE0MBrZlTmyand/o5twlJQpIX+T9nX
Re+mRacWB3Gi4W6KQHjOcIEBRtz782HE6sb3mLiqSiZauUa2u5Ev8Yq3/BeR3fZn
IlgrSkp3wNpFs48wSw4zMPknmRcIOI8RYsTD6eSGGZ8fTfNLAjhcdkywAZ6u4VEf
xezjxqqBK+PNsgu3Mmu8rtJ11fRoNPJIeAfh/pnIIRfi5I+zxHlhyj1PGwJ0nwpr
MYtSOckXnCiQmal9YnCrGeq6I59txabp+k0726Fih44qKH9DLwESqlOU8P4d+gIc
h4hFI7yEIEi+Q/gG5rFgksVMORCAjzE3CepLeju9+Cqd382ugeZGuQiyj/lwktSw
x1a8X2EQXzxL9wsErOFhn6s0DdZNKDk8Bmt+nLkPRO65r7X/FyJhJXirGN94+D1m
fu/jFK9246EtqtvRnA8j+HbX9p3zu+0LDM7Gx3X62ILQR2ZCWJmvxNxbZRdXU5JR
BuhKC4hZlg21fgK3qVjp7N5QgFxkrgrNgDrtlku46bOmzruo7WRDYN5+XeaHn5pk
POR+PwT0Eo/YUEHGHOwBlRFSH75IXK5aFwup5939Hk0dnf+Fjxo3jkTGsJkoOyCe
tpE4rSIGyuzvG37CkHVHFLYcfcek1MSf8lmmarzwzPwfN6qGFiTv7nFAR70NjDdk
sJ1mi+5O5wOgk09J8DOtHwl7LH5c33JoE3YNu3TKWmylmVr6DiNluLh/6x2pOR+E
B9TYHJWuDd3E6ZxXuKhWwX8zqqsX0s4MeJVRrqUF+0qNwiH11gdN4S6nHEMPRA7v
et5N2Ytl09gJp7XmJqfeK5aYrH2SCQ5+BilAUvHBmkeN7FfNaa+p5IUZjZVbdJMd
S3FRhooS3i4gQ+mn2Lf+ALM57Yo+ah6cySlyB8b8bwZEA2KSh358EpyGl0kzX6hS
OEr9SjVNynRkXPXjvPbI9XYyzU+FQCWJuujndQStNNhGC8Auy9SdcwXEF4cxg4yG
zRuDvEpHfkGPV8rY+VdN5M2jZsxKb9E2O9fyKwajwN62h+XfGpElE+Kk255GZFCN
LhLR5veWnR72juU0OfAkCOpAnoCGG/Ehnam1aygm3t2DQeeabSngZjie1hUY/yOE
wuhNyr5slr0KEOlSW4orLjVJBkYBS+KFqHAgU4GmrONB/8QwX17/fqmEn7rloke0
iNCG7CW/trIo1KhGcKT/re8VEdx2TWyiFJsKTM46iM7fD9s6W3YlcJ8SA5MDwqFT
h7NXge9MCgKm76R9muzGDspL7ovN63DhvuaiPC3UCtuyvXMasgOMHHIGSKGHtnAj
tuh4b2cYhpS3REEsitgjz0knO5MkvuAE8yOdS1N3bi5XaRN7sgwz8lfAlCwDOf7e
pMOeqBb9dbgnkkbyJ5U4YgSOIfCj4rTDLqRaLte8JAZandRMQK/n7NCI5x7Ziunn
hFk2zFa/ESw0MlDFQVQgsgpqHbWPfWlV243c1vXsfgFMX1vs/ML84lGkKyKHE6T9
V2wfE3CAB6nQIsL/E9CJOQC1eYJtCmulyX65iP69GC3yNQ1E3owaS0SGMfyOrXBR
haLQAb+CnDlikfjD1cf1LjgnZ5Pci8ptJGp1E+PTN+Xaj37JSieiK9GuGuP2Kji8
biq8V4PgAw31WY3r/lSnKGrt8+IPb1gOUP40eX7EmIIDtrvqRxp1MRjTjqLOuBMH
FJY/IpH5kzfjxCmRI1P2P4baOgH26bPqxMaUnk6kRRJbuBVvowdToapPzBS0vuKl
pfIgQVPq/n6Q/G0BwQ3PtIR59vOwzRN+/Mewm4IoqN+MuYMM5I3iAkbWvACWKCcN
XSHWKEScKiGyPw61vMZk2HrhOsxcRQGqdOTv3Kuf4m61/Wdo3ZZiU1vuOEkDkfYc
iv0gviOTs0haCdZGQuzKI9GTOlG6RPYXRtgGsCB1tFJ620t+PQ7GF06TR7nKIg1g
yiZ20NQhr3ImMmxqMrgL8v5eCI/i6QY1pTnJxdV8oc92fqoYECatRFOiOHhKXECK
8eYb+VGtMAIIIXcMCTaUngfclX9r0n8JjbGxNwAu6ftY7yEsrMacVPLqtbEQcPb1
dak0p6MnVhXacrAFuxBYw8LmjCn1y94EATLGeJZ/kfUaC+zXUefH5i/FeiI10uis
R4vW+mGLjdWzMYanV0qp1uOPslQ2bdH7mPOh9oiZiexTo7UP3hPfQrbEYj4LribK
L+alNBMxyy5H4VlyFy1FGBpJhvY+axEB3DtYiIFaSvU+KgzF/g65UmYZ0ythlUfr
GUjGQaimhM+hAAcuE0kjrRtS8kA6id5ofBVDM3EgRxSjvlftUGhel6COJGP4EOSm
ZoECYWp6Q7xwcrRLz5pCxyGVx75qOLeaP77sRTwUrC9WonOs8ho+PTPB6Rd9V/NY
Xi8eHNWLOqlqPRjvMlzWhXXh8iqiLd0xvnhiXsmhtzhCihlamHrUOnVJSxLk5Dk2
9vd2mJNEoqMDx0DBTWRjInCBvOY/9RLDSYCjGAxtYDx4Fg6caKCuZMBlV5VrQM6w
mNZ6ZnGwdxfyCVYxCRFnYJAzdGNirHSZTqkeAcwe/05Ta1EgaSWKhYRbBicNZa1I
9FopeTKhRwMCUOSa2/suF540kw8H7+Xyivo5yyrS4P2Kq0s4cuP7WwbcH8yU/0Fw
dPVJCq+PZQb9zJTgfc94moVxKEHd9t9IahjGwxsHoIHDLxpm4AzXtJEx+wLdQ4Il
xu1RzKuqJHXibi2BPhfTFQNHAJnHM6OdfY3VvcLq9M3KpvoHdBcHwf/rud51qyIS
VeU84RBL+XsNbMa0NLy1imX0LCYH1wTJ5zoDbfH23tBt4GVzoKIZKBFYvtAnfU9Z
6c6Fhpek7WJtQuzVTsNFm2IH2H/1fK7KWegAO7gZu2LcTvZzWleg6XZ3aYVBI0fF
OG4Ic48vdzaC+lGPkghoqfB7BM0KFTQI0sdxRR6Hdnb/f3qqzdzVpsSu/n7c/8cA
1kqsoP9HOoRsuzj0xCwu2MXns39bLUDnzpL5Lpn+PDDCWlQwMhFm2aGhxJBi5oB8
8lGCjTXfuRNj31FgnuROQQpsDykzLFwFGqF+kl4rkdQAzxgcCDSCr49EDkpgOcmq
c5R22opQaRvfb5u88ljTyNJfNkaYqG2sHYtlepuOH3VqsTNjGgioErdM4EXNfKcf
cufsDBdopxeRRBEvPVbl86PH/fuTpMrmK65tzJ7AHEqbXOBnJyqh4MjsmxwahpS+
1gHCAT061urPtpBjKLEcLumHMlNzb/rJyia2YN/i+GMUVU2/KN+4diS8/vDfRRAh
qpphNxK4Q1cVpSSfxyg4uX8n0xah88PY5cXxZLkMwnPBvlRHXmrqRowdeYghA9Oo
/xVeSKVnhqBmqOgaCCeMV7vg99vwAR1pOQKOYpGz9rdXjhV7RWxjvjQ5YninK/cb
msTj2EU4gkbTe+zPW3mk+TyM6c1z8X/OzC1p3gqZupZhh9KstwqEbTgrzIBvNH9C
Rx1Mo+oZc/0ClN+H/hAw+b05ydmztpvWCfb9EooDDEbE9I1q/fhzIjGHXwwppC87
lyftrn8titSTAOhDx2DApI31F85xa+XX4/C+AnHmWSB/lUiA5gFlwUoOkZ0eq+Ql
YIIWqNGwQLUbElqbZ1sKaA6DdspMcwJFV22NgWEAqRVk+Tr/GPk0lsZxTEAaIXsn
+9Lklvo3RSSfuWLSwHHqysq3PnPKBwpF2GS9e9s2Rv7DIS7Kwz1uIKdT+UcCQGMI
TjE8SmciPL0SedfiWttJJxiKsnsJpawVtlmIfka1fyCu5UL3kasGz0hVQYYMyQLc
0hcG1BGM/M05IacItxqO5IKSZO6tOvaYE7h3UnqUMNHYUt7e/sRPAF27SeXnjbHD
b+xN3F1b7hfu8WiNsv18fPbtKpvqarT+ujM0PkUv1GmvJfwCpKpTiv5jfQXKxVg7
B1/jqzS8ZC3d3pPS4XPZXV5oRkRogAGvQuM/o60GMfy1dgN+upWONsPOnvKU5CRX
z330HTrJV7r260O2BU/8OvD6IMV1Mk9ixjjcBFBhLPm25DZ/nmDOqqwy4K8mwX9J
HKojfRHLyG7teZKpie4xPpHA3Slp/4b1OOoj928dNnWFxNxBN1Tv7SPVI5bUl6rc
dAEKYuBUyj7ukr52CzHJrZnoypWnTc9Cu+ehY1qJcIVVq9f0SwkspE6XG96flj5x
qvs1hFumawDpIWXXTuE7iuPIJyTJeIedCOcZob5Wh/t9R4NUcfWiHdp1IE7L5N4H
4Ka+pdCG0R3TMhnlCUHTn0Wv55Q/IVkeYrimyXXRiOPzxYLeFfD7aolyCC3d4oxV
i4CXGoc+0bbcoE6iHIvK28Dy0ugMO1qWzZkbowouIYq3MRYTXW+05z2YUq4Xzp/X
R5Qkf02+Wc2g4JFrSr8rvGyu+GOLqRlKRaVjb8yopCWunxX+ekL1hzQdvKNakumr
DsmkpI7JaPTioT+BHjqlQlVaP5Up5Xvla806Z+zV2rWBbecdxnpcy2E7G8CXm5Ha
1TAD21KTUa2BFMjR4rJwDK8On/u9jc2O8YMesRjwWjAFQJrTXjwvwfCyujlIrxaY
SrewX7N7YPuCQD53Z5xpr8SAifXZPKd+UGOl6onL2LS9rj7jTdBk9hS6GbiG6ebt
vuVWWpf28b7GrHEKog3N2BfmAqC/wqc51eUEsHsLHYLFjltHAfJ0qKpxSObO+2Bw
aqaiyCEZGnwnvNyQ58puQDLiEe/Ui/tm5VKOqKrRRnJIsVfhDS4oszCTW+Z+MPMu
UNhF1kZ/l81CsqAHy+yvSQHMeej88Ve+hcxjuTcbfMv61j9tHWZyOoSumq9ELS/K
m818MVA/F31hqb4BBIuDpbR2Qqo5QnY9jIEeFaDhp5Ez7NVy908owSXfU4Y4pqfP
2oTte2qBIzy4YPaA8sz+Up6Hq1ZwjI7C1Ny8SykqARjVntduNscRdHvptMMLhItt
vJsOwke5xjpa27VxDvDC+2W8MxJ7knDwJDFqKCp1MA8rvLquSCYPRLRarJeQmKJa
tXtecbm79kbJ+0/0WeZt87OE94La1UH8pxWxZeOdrW8SYJ9puXPELl7MPpUmb1S3
SRwT6Qr6h0W4Ey1dLthfKQl2rC6Gh6Lr0OOWJNOjGMy1wV3P7PZAQkj+o6Ep/R3V
goNNwqYTvHu5nus+y3ThRuONzL8nLCKDlEqbD0yOf5UQMZxYRZORkxCiLxP+jtKI
gZm8V5E4Gb8d0hjpnQaOvIRZy3QKrAC2EgGVSNmVgQmq0Y6aBPwGPbQ2HhXvAYip
v8LjJo9NKdS0E5nwTjOX4RzrEcNZ9I1Z4+38AgA/zGrkro+05IBCcPHbI5NIMhK5
EDVzulAmykAibZ7gb7i+54pXuH38pqyDyqWPYZH4BBSuHwh9/KQNoMEJxA+gvoT4
hidlEjLruR49f0i3TU1BCjtyP11qxBtP0VlX9I2og271cFqJ2eHKMyBk+SgJ/Tsd
zCH5IwyDMyUnxTUOktSmB0Uda/xzcEIakbB07GPnnCzG83uFbz9ktRwCQU5UX2z0
zCwf8g/qyZsMYG+IZZ1v7inpcK6FRfgA81lZNTjX0AC59RQZ44Fm1RV/Xtc0ZvrM
Lvh9VSU0fcbgxSem3dlPwDH4qUS34FYKPdH6jl5mScvA6FqQ+fBwpNgjmJ1R0dnE
KORAMLTK57FqOcmLv5zExR2AZm0hK6jk2PlMo9Bi1gJ+/P/eGN1ptezveutkebq0
H049xv8tjJoNiPCFKq7XlLVy0O/La7axdSEpR6dVr57c+LkBxzkTH731+2hPt4Az
yuIUMt5lVPk8bmc0esaOINt5zctwPm2+p1dixSMtSPTbwDofVyAMUPfEQ/ums40F
iafipIX7qmqc7vS/TnISUXcnqJ8BZmr6BZO99rkvIzTH6oN9fGMa2in+NJ7ASv6U
bwfYalGDGkutLXj2UwQVSOuLOXBe2FFIcF8ZXVqfP4f3lH2fUU3STuB+b/aZe7rw
lyddgPsFlSWstHixTjBovHBJlLTg9OQqap6l1CsyxxYAmCKlnxXlu5wuOxfSUyyn
Tt2JdWHefNbjBZZHVDEk2CCD/a7tLvB1alWrKCifWXmn4oZQlvAt6sgHGRDGS3Eq
+s9Ngtzqxu3WFEBW6Uxa+Hlgmp8QTTW7xs0WWrmka3KjagNSjv6CYaIHej5tvJKH
0aePLrFn+gSoGW5FpFVZ6Z0DC0ROOs2xWRqIeoOTYTaqBB0B35iCqU3yWwcg854S
ik8YFDyPAmyiIg0osSvmxtVzqEIrZUjwQsOrH1/5R7RRAEwC559GrvcZ9ivGL2Hw
5B9O5N8y45xitvetjt6MpJPjG27obMIUypmtmyVftMhjLEwZAf7uiNYJjG3UNEE2
+8i5XFuYm8XMpgFj8lmsd6gWfPOhhvskPfblnl9dEjcH6c6ahwZ/F07AQ+LSt8w8
UHFuqIOD+c6CVHQ2pu08CqOwtUR2tQmhi2nQSvkPsDjN5ZCJXERc2MfVUpbH/Yh5
MO0dotgMa1LVZir4N9ZudJ/8q9PYmXLLQj8K28y1yAGPL0ZtVGLfqPxBFSQl4sk/
b0zvYEZWQPBjvAc7MINFjBxuvaVawAK45SwogkXVOAPiZiO7ja2ruhxMdwEuHJR/
7JpbV2ihOhXxy01+CFhizoqzKhmDdGNbuBEgtzzSQw/TTnyBL1MKD2dCxWvLpsXy
LbCexqp7plGHcaqRmPFIv0v1S2ZWHkxdW00a/NstFtdd7daBZV8loB5tk+EcTnsc
KkaOv20NqcFcCeLCs01u3DFcL4SwpslkNZCX6Ot+nzhjUOj2xW0Jda4KclTuVupf
nKdbRNicLbT3ODtHmBiQOmAxBl93ETiGcUXzGpJyKxBOv+QZYVwCjXsMn9iRMBYS
HNt9o5WMAO87Sptku/2ZrMAY37+OnRGzVnYC3RELQ2Oxdp5d7nR5JJ4DMPqZu4sz
TkbrhOeHPdBkdzX01UiL1KB3FQGMZtL6cdQa4Icexyowas7N6dyeCvaJ/Iy5moRn
Ct8QIN1lLDeoBHIhcp8TBunSmce+cONFlKli15WaWRM9i0tMunu4DuRoXFHla/gJ
P8rBBK9GEAKvbbCmMBj71x9CMq+p+VMEzU9ZHSuSOtXmxUNfwn86hY1CW3l883ui
PQuW9F4cSsKtHnJp+PbNyHmMnX183+pJlUOISyRh7kkiqNjTIP6aPoHXR5Zy40h6
uMMfQgUHhw27l7VjuAhENpQplmM9aovVcONlfr9pJ/KxRpQmbc4vZKL9h+V5XuxB
tvxQW/CjeoZVLL885ZcsI3uUAx0B4mJLCjLKFXZtLOAWn0jOT9MxAGCsmylkRBNv
X09SwJUh4P4sNuquOyY2j/JBYGEm8YPK3a+63psLL+jCItxM5ezYpeKGb5wXWEKE
CIYevqh+5S64T4WK5lAr0/LKLVAT32IMqipt0GxYow116gyfci0+pm1scWFDMHbD
XP1T9He4Y+hUkuHstepx519ndrWLhFpQL15Yq134i5IVratkSpYnBUQPccPo+ZWv
YivmR4BYefHlU0mS+cqyUoOuhk9OJ8Gqw/N7HmSB9N6RR/wqXOOUYqduURJeR9NB
9O6b+JvNCN0Vfe2JBWT9tn02fiX7urx3L4nMdEUH5u6eXk+Wd08xD8DuGu5ffNZy
qz3Cg2P35vemaxhgLezo4/IFoHKjMnciO0UkoZe6ByUQE4FJBRuQ87wB/hJDFJH/
Ud5mL/3POAai+ZVGZZe6Dq/uDfIso3ddUSLFVJBB2792CCgQszx6RjhKIzoOfBM2
F1z0fOACNkXDu6llKkOe6fWv1VbMSM9R32o6Dk290ECIjpxJtGmkwBz40crFR9bQ
cc5Tw4hcjcOKan9yTfkPh5lXmsilwCBKeE5L5GfKc2CV/vIZBhTdgDMnzqer4BfT
3gAwe3PXCwN6kID0o+g0a/8xL3qJGYu8tIbZO65/3w0lWj38mI+muxPNNM49rbwI
a0UKtHH0rNq3Ad3IDmWZSXLLa+J4RcRpUvISuv8QR6IzzGFJy0W/UgH8mzoMrkIC
zme784ue9JM/t6kUdAfntwW26Yl7zEi4A9+ruIPE8qbxw2PoEIHBnwiHrPj2LR4y
J238oapzzyT7AQMv1fgFCLYBBvER9Yd/n7LFAb1tbbgKrHW5Ii2QJrF5+PXfEhrD
Hh0EQss0L22d6G5s7yUqf9CjOAJ87Nfz52U/6Na2W/996w0Syq+FHg2ROKxm8RhW
n+8ZqW8gEL6aTllHCAaUeyXJmCorRX8tZYF4mO5naPAtJ+R1bVUQ+K8BhOyuk9rr
v6L31OtBfaSt6TTRlSHDLD+otOdWR8UhpueoiP0QQ7zLt8h9ihNwyGEaslWV+fzB
qurW0niZF2VWWIJRH9OnpN9wWQooCwMmOt15sKI5TEnl2b7ka/S5n5NrptysQn4K
/GBALfV0hO7BMKKnYzcfibS89pEQyIt38X5NFg3dHnIonD1svMZUVtqMSY1zynoA
JRwC6DGOUjTXaO07jvbQcNP+vZIBxgsduKxP5l1HOC+tgXiT+HIBfsFjjpeBdQaq
RqSajRAYfmer6OmaVRE59YGpBpJ2GTdQTElG+Irzvzf8xUkFVLUpjZ/wXkZ2t39N
sAOyoGFyB/LRKMRMYjAtkKf9VLJq1gM9GTIclOLKsvQybwUye0sGw5jTg9wdT+Gx
uitwf59Z1q7LkIDr3vSOh5hSTPkOzJ2btbEaR+yrTxMIajawz+Ey4cPYSCF/IOgq
cKQyX1ppakvCbKMfCOdOgEq6s5RtwG5pyhByFaBJGrC+cnS03hRWVJkMvxViFQ5p
OIrp7qsdDYHL2hqiA9TUWKGWN8jq9XFMJUOm3k1onIRf+foN6jyY+G1+Q1w6g9Nq
9Cn3V0WpX5T0EF5D94FmoZxZ2WMj3q8JPu8XyuzAQ2kwDtJpBExj9TUVS2ILVMyu
UlYYbVyJUTmIVvE8vjDBHk08fRGO2VKMFhznnsLsTB+eaUWInEHCggHUc1EjY9ZB
vdZM9gM/2lgRazjfkoQedQahc1vuFtZqH7gONdV2Ao2b2HA9TLjc9XKL1zEAd6PH
Qxeu/sKPRxi0iy9btvkgEsEcGhJBdIkEzdixyh5h2m/TfGKROMdyhGTMqXz5UHO+
SUd9eCxSzfghF5XOm+8FGuj5KT/vpfIhLGR1yDltELYRcmgrZdTMb609xdkVZvlb
j4yj4FJulXj2djaIKPfhmYkKqwkznDb/uBf2lpzdyG0uVqa2fvaOwCb9/EbPidxi
Xx9v9ArBq/5XOpVUI5TxMr8H/H7PPG5WxKAErVV/dBA22qoCCH0UcC8eQtjEctyp
GOTrX3yf8eHYa32aOoeEgqpiGh3VjsmIlwhgzqPI/K+VngIKamj20sYzsN23S90z
ZjHPTBUKLYEoFNWzpgwARcoLmwFnwOzHEugQGjJ3tNFuzY2O1kDkyo5PVR/GZ6zb
+tDAO0PriyrGfksRrzKhrNoxne6Sa8iQtnTvsH4mzt9X7TNk4fEPsLWnQF8u2Fge
2Tiudqwf9B+oi8oPDJoyfWBny4+cxheD/DFgI3Wjr++VlqQMKpCJeNRDMMfXxzaI
zYngkc3O2hM+j9A1m1+tmCxnGlQ2x4w5fVKH206lWR2neAu8vtma8clKB/TpXczM
MDCq7lHzNQ9hQiMrzGDwlHcLa+JsY1iM/4OOpsyAJ2QS4cplFm5kZUmLSC21HXMk
YHhmHkQENjNHHUE23Ugw2JErHtXwdHzw/2YrO8Lo8CL3k07HafOQ9mLQM2gV5swm
MOPqCc1oW4YaRTiIcedZOpwYEgNYalUU7f4Hy9K3suzgSX8ZzF0/bfIbfW4RZLXX
Hnv9nGHTgfQM2YW48kz/9+JdPHTQ7B5h4xMxL9oFV7QBey5oGR/ANvE6u9AKKS0o
u5I0n+Ym+CKDitebLGFxdt5y8h55IzRu+5DQ93Q+GNVOz+jF08Hdd2/tf222XHDY
LXwwSleomQo7wb/3BzdlPIqDV7/9hwQofBBA6hmzAPyIrix+kQm3JfsfR3JiWS4M
DzIwpjn0d8T+KXbeDyr4UxImBEGchUyDEnVPfcOFyKlZlFyIRs8g9F9Nt14plsxo
JUgI1yRASqW7A2DKjF4k/IcHqBEzDYfKxgoBwTCVJ7S7ZGlaAN5IBP04nKKAMjOl
cxOCyr73ad1f4dhXq/DgoBHr8ltyuSybWSNhOQCYJnPPpiHzCXHEWpZ0VaZkLrXi
ZWnR/bSvZblHZ8DkkLkDqFgrRw//jdRxQtYJvEY8no+GgXA9GIG1f0f0uLJAkaFf
L35uGiiyyBHBnZJF83qREw91w3vpYPaZuBqE322z5N0uvKiQ/cnYYASEuxtEld0M
W+46mEcCHWMeUuXvvPSYLac3yqE51+Efe32wHFoHJuIVIUef3NWBLdUrx4W5zIzW
sNpc6EHc+b2QQFiuyeF+cx0Oa9HApXaLr15cqdoDqLP4gc9bYWPWc5azYgOC622K
Jx8D11FLIpQv3JmC1zH412EK8qTxR+sNrzeRovEl1Ikh7Z5ov4bHnapShw5RNJgu
vWu2YvoEs9acB45j5uiVjuIDMMIeJo5ye8nIMPPCyTqTk9hQcK9tD/EWuSg7hJwJ
PpRjCFLJImaUKV5tVDz5uegCWSeh6QPI2I34kE5uAgYYDMdm4aZUasUGnb8Jx9k5
QeMFvjRAefsMmbVKOYVTt0aYct9pl+8gzPUPQVINfHo+IXoCZ/aC9wJ+hiZ/0uO7
FAWONuQKw/jZ/fD0yP5WmOBMTxWdCLcOkXFwDvgKzbjHtQx4almnK5XzIvQgTPr1
WVVbYT6zvBX7psnzfj4IjG6w3OaVZu8ICixAP2yeINfnvfWR4BbsIaL9MOMo5qC6
33uM7RKgCAaSPnWa1kyCDj8zeKv3jfTR3S6meEhmgVkF+c2IaBmirgyg3dEM8OMG
OvVuHqjz/JyA6xtQSMhstpXvPZO/vBL0Qts/6mQ48J14gAqa/VBqxKd/lHG5XCuw
EApJVtNhm5qReaNXhOmBN+ZeVU+i06DSNaW3CPPk0V+GoJL/7nmBHTduLtGUif+X
f5k8NVFk5YNt9JLgO5AgmdvJU7e1bBWVWXoYbJjkQvIAMs0C8BOSPaMHaCEQ+0dB
wC1oYjeHafKk5q8xFidWc78nZjPEIui1WnQWfVKHs0vZBR0UxfqbF1gbgdLcunT0
FAxDz+jf2b8ApE4wI5OS76frCIq3yTwKXC4Wd72APfhW5ylI2K9epcwDSSXuRIKM
0WO1ndc58F128V0iXt/gJihiNQPw2Aypd9jqHSRTPlxGM+6jUFakjKUOGcwO7IMv
15YhawzdRoyxwFbR7b1zue14555R2O21MPewT/+YY195aiz9PFZivBqm0NOYeo27
XJI/wQ0qa4mHBD6rSieCRZuwZPZsAyW9frejqsV4r4htVqf0vSsvNnmjwDr9Buli
FzjYXWC8CONtVnMU3cpjvGoE0CV3bEFSstB6OhR6uowUdF+1bh5uxp6ZbbuaKWL5
HljN/HzV50eOw2KPaI8rwq1dhpu6MzEQp56VtVZAw6ogeeySxKiB/ev1YGF5DZOw
w8ppLYO4T4SnJxktxCtic8xgpatZ8XQEaf3vC1zu5epZC2w5/vWe4YeDhtOZq4NQ
/ZFHiyIoIMS23VpBm8vuZmPmAw+soQG4s4lwxpNyNpFDExUFj7p/N8ubJYvnye4a
OGPsPWti/3uaAfubEFHLLiMzxhuomYo3ojWCZmkyD2YPlm5a09Uvp19f79sawhjT
2+zOszaly4J0l6/iEv9udl3+JzkxIvGCHIRwxThnq2mu31NqoglEocfowyDWv8V1
Xkks3s6y6nQcmmXKuR7EqkELWsmt8Np0kLK6XlxD1CXpsoU2pYIOSS9K3cYaC7rR
y/W6SUijeTqEKc7qMf1QEjvoQqStdBB8MooHbuNFDRVO54JyDzRA0wdNKi+VBVkB
dgd+tMdatqkRaA5OU2sqkTJpo+H5Mhabqr5E334NfJXDzUgxaawo9UQRixcszsQh
6q+LjCOg2BXZ9Q/HW42auK6eRO05uEhTcfEKRdQaIVqvmhsQ/ArChSt1QeMYJUzO
R5F+6Tp1/8CQRnoqOLnK99/r4ZDAkG/esanCZTqIg+3vJroeqz2+YQd8twPplOTj
xM13iByjXg5tFXZdWACO0DoAuds2IamyZGHtmsVSnyRbwiw3mtURmf/kraI3V/7v
R1+hrHxDjQdulcftLk40wLDMRhOrbEvchpMMtTZN198v757BNxP0JJSVcvmDDEso
Eag2fATdQAoVzftKmsyZUNvGUk0VJ+ZApktXK1YHA7w13zZTVTqZYBjMv40IEvVk
5sA7stU5ysbxl9kzayfUo0JXcFKKsgJMAiI3b0MpqLFxG06PyV8Cbewrw21b+xHW
yDaUdeQX5hg2cRNJL+2YOuQopZOVLtz3h1siY3xusCbbCznjASCu7VxtDkG9/Fra
PxlFG80x5XHDFXRGUnF2gos3qiSmo5ALRwoRIvRiun8/yNI6TpBeGpgg64x7GaSU
RAjE81CijeXSc908YBihTXXtEeoVftfYgtCO5adrgWLYfW3ZWsZBl02cy/d9HMED
6HepjYvjAP88USW64dkolzpLvkXyjc4UDc3hUd7xBSB2bGVB36ebrBPKh6U5s6TH
q9t+pmR8v9FhUv+8pmIjaI/JrUg1NX4IIs+kM3WRVyQCRrQXv7a2yvuH4LUkE0M6
dyRvO9eupjiTAns2yJ2XRzrxTLPaPG9mIy5ce/TmebF2qVckLjzwQ+zsCQgGZwA0
N+94G0QPpPLlqQEb2RVajqYMcz4/u2U0/vLIaQ7lIOiUyDvN2uETfyFhtF9UCJjK
C1j7T5LQWWrTzGXriaRsbNRS2znKV9gT/ZfBoitcY7MjQ7QE4/3NnU/qxihiZgbT
iwR2O/zM84zeFHLlVgjgnJjzpzToH7yvWe+ISDQ5EQtlFu6+h+AI+NqymMeFMVkV
/bLhVuyYbzYrslcPN+GBpewR+CvFtmUKIXb3LLojJFVcm1AFHA84/cWNnnOfUBDK
MnF3bdOUGbAnuZliH3AQPKw6/BDLd7ZEjaFGFDlBRXxEoxKFRGlO7zssoa8WcK9O
p8uuJ5L/SeyiXoDizXq0JxlYIRsadgvDGu9nPrUAMlTN6TMlfbtMFlbDxwBuR9MU
eXX+4HLrThATyB1iZRT8jqEk7W+n7RQLDK1TlW+l2KCNi6rh5KOkEh2hPz/mS7Tr
JgJgCbIUEXGAI5Kwc4vrDPYo/S7GCVFp/aP2ihVH2EpaLL9Fnz5sPO9TAMlWSkD0
K/hj0XQ0GaME05X07TfANVJwaA2EsmdvI7kmkXc+9exoQaIOlwYhepDGnBTyBHlQ
4icPhrRyL7O+eRfdLhV1waR7w4BTk3eQk/V1ouSnjWlnA4IvmxVwotE5STgbhPoP
Gq2VzxtlWOFofFuL/tEi8nIecNY56mzfwyryFI870bxdV+PiVfqnD0Ax+nx/e0pD
1ljxs6hfsEENNC1MzPxhVbYaOLQV7QdQXnGobKMp86Bxs7rbhmnhjOztaXNgCKm8
wns1uUlu/sxM9T222FgJjL+55KnDWRVPCy3HGeA3IsRNbJEeKz/8O2KwvhBf9PhB
aIZVd1Ubj3eRgS9PgvJE7zzR+8NmacvsoPTDLyrAzQZNxIyRw/pljXf1ndTb5IF9
5n2q25ULGujXQfg8YVLpTqCy0BjJipK01T32WIg1MkhHx2OKMOgTw09H+kUfVAFi
e6SE7Pw/FVb63tJOl553qDjsITvZEJH7WfvRXzZM4wnvlVpPIGr/sK4eHLQHqMp7
u1CHNzRKcwSPkdOzL2+JzOlJV/+p70zPUU5oQpoA3RHORUGOaw3mvHBcexk3vSTc
6d9m9OcowwTaHVNsS2gmLYIcbzbGm1LhzJQVh/cnqt60Cp3w7S4KJF6wtonX4iwp
JphjLNlpWaqFn9bV2v7JIZHKPr/0qJdr4NSfst13fZ1AUdtvCzRgG+5/COk6h/U8
apPaNZWD58xj9/7R26PFdVnechlbebImXI0vFNfaP4p8JJh0sOuH0F+2HTgEtMSG
3HNLkAA4yOMJQOaSASc0bYYAwT7tIqijM/dLBUpoVYoAue3jTQusAR6un06shfzN
MYmrIpvTv+ANE6xsDCeBuNJb3fD5A6kXMn9KNFu/QDp1H6tz+TdM2UUP9BkotkdQ
yulszEirq4dPdMs7Gmk/3UBIxc//oJIMvRW79/Eme/Du35KEsRLn40Xj8mVGdtSB
u+Cc1modqWsFdV+QR+SPxFfSgVwmw44MVE3y1p+SNwbKiAwGNNEVrWJGJ9gsSEol
BG/q3iEEzUOcNTbVx9ExG2L0Ci+sZJpEhc0SuJlf0Lw34nj+PDpI+lqdmvZtMCOp
gSwXa+BE8ZcmBnGRExzdk4KdRW6PgRTTxjlUB4o+4VENTv9QKGjw94MlsDfCIpdx
rjKjBGlmx2I91gH+aCSAwrRYEeli9oa37xJ3XKnBpBUWD7nMML3A3+7GzFhgOlCS
yVZjqx5QflbRpwrZIFHh5rLnXaPIOM4tfMphpiGcRBZ3k0OvPcocvw/hlIv5xvNA
pY7nmOw7VDjW1Az94BL3leEovr8d+K1U+Odqf8y6+Vfa3M8glSrRo4f/jPudrrDH
XfielpgRPDnYMkw9xCambemtXuumq3wqegR8DYq5Dg37aRXC8lI+BKKsdkRawqOy
YajwCswg1imYPsX4SMdP0P34H8rNtfXof+uiQYdD+iLl5BSMf21KkYMfsA0W/Kg4
mMgglUW579X2kNL5uoxSuZbui66h7iPTubl8UiNM7WNO28P9hwckXj2YwSyjPumM
KF/h73GEhojR7LQ0r9jphvUzpkxCo8oBatxHX052aCTDPeWeosoKqpPHRIfzSd4P
98y8e2ylFSlH/vZx+oOQJ5NiXkFa0/3eHOrK04E3p5CcVu4Oi7Kir11mb58kGJ96
7p36RPTBRtc7gWjooFWpgbxAvatgxfxieRU9cE5HK5Prp5yr3Pk3yuh8Flsf79Tz
GybkaEtL2S3K7AKtpBcThThy9zppdk85C1OA4iFsLKY8+mAzUkyfvg1hlRWUtWCJ
QYMD9Rh+A9Nst7QEja/dutSl8Dj+l5qFJD/Z8lu+MeLx97YbPZzKz0Ko8Jz8sFzg
QzVLCzhHGXImYPySzUrVda1ryfO2Fo/sKFePVesYr/Pbdn+zyI+ZB2RwpSYAPMXu
46th7E3w8k63vYTii2YDlby22ppx+kwj76Q4e1oJ0x98aOi10gdFLSVPz7WY50rO
/7KFFcM76Zty5Q+Qn3Z2s+nyj1I06CrZnxsrZrCIst7Pcsap/rEXxmQByYtG1V22
Xo63qtUunqJqMGOiAXBi4vc5QEh1sutc2MiuOHIPgpVV3un0wQxKnfaH6/ivzUf+
lH33ghIpyc+NvNpVlyF0jEqfsWk21BgBc9B/tN9OiTQhjDEph1aOUsOKVeUXfBps
MZxTDuP2wzDlcdmrzLKc84suDgCFLq7EJV747HlN6U9zc17yO/1s3FqBAlE4v0NR
7otc96gYQ7NFz0BLyCK8mapFWwOZezziYzFZfyhIrg5XPA3gSaJWo2JnjiBOkSFM
xlW5VZKnAPmNYt8iIggJiDXonsiuSk0UAx4cbOBVfHpEjmvleEIbJY1Wo1A0RK7w
SSL3JKDXBUWdrpdZrS3az4zRBh49Gt2H12222/HFOBpAiv3NW/Ass0jCZlgp3vuZ
OgJpj/Y0G7N+V/UPmpfe/0cYsouUq5VcwiJ/QnCfS+nuugIpVHBGT2mBsbWJqeN0
uyJWdyoqMOsm8IHwcZvJk8ChO2+rXAW38DrT91ZPItNqWRdvgpzUt7NZPTvoHz9A
cuKT4/a+lpCOusWnWqefbu8hzI1BycHKy18u4eyn2l2VzqrpWd1UTFTqc+h2AXhX
Oz/qwPWNzXqjUD/0h6sd/IPgM1aSMEI3sXx6RIzvOLLHVtFlKneBZaLAeX3z8Ftz
GDhTteFeSBRUbR8mHq0ogiBwkymJGEcPby137GTXADnUklYUvE62UJOxXEn66iL1
JH00I0lFK1h6tPkz8jaNxVsmYrKGwtUh2yF5KLYEF7eJmOegIMfVNGBV58LA81fB
fY1xImo7v+Xy8wfkqqOGr9orsorJq2UxOf2zz8PwLgteEeRsZv99QhPvbFtmXhjc
itENLfiU1CBF/lx2Fzlmig4iIdrY3YDXQB7XrUN+TuTP1hdJwoDl03gXK9EjAiYY
0pjC5VVJ4YLjRKvuD7WDlB/8gv6rzPFhIB73sIlt2vX4VjU0gX5j/0/1Eoe8zzQ+
HazrKhWq48ZFnHhBSsWzXGr1BGAfhUmWmG2U+l1IDvsOtBvdwnHGMcpGoP6KN+IV
CB/hgGSKOiKrby5artIbMBKFJ+a4yhQe7vEyxO+thkDm42hWjWSxa3Cvy1HG3Y4R
B4tLtTxZu26bXBcW8rHYgdGzZirk5NiVyThvyge9GplAmZlEtnPrAcT02udLbkVW
cOvXo5Z/t5sOuXKstqGHSiXM43+hyoW0rJ8pwclD7sm37iYMoMDPb7lzeZuubmZS
S8r5uF4nolNOG997hqjKIOA1hV4YZnFn3VlJPK4CGiWff+DUe+m4xDWnx/MSQ8py
cbt+pBjnA5D4EOm9kv4rumLMDZJBnDGMOa/aSrjdc0IAuANaQJ0XRCOSpKFveepP
zIeQVTZuJt3bghaafUks1XIFgqHglDi/aDHEhjE0gGxNVGZzCVk2JUPC3SNRld3r
w6EOHSPPGrqsGJnLIj32yp+/F3Xe2k/aeqIx+P1Vww+h5IM9QiPDvcMc7IZvosSe
Ep1/5sTC6s66gAsPDjE4+P2oLxPUNjCAz8RovKnMapAeMQSTZfXWVniStQFevJYT
Ot9mPLNkfLUyAvEDEU+9d48K3kK9mlP9DpogbvHF0jJBo7IKjASq90vRexJ7+SlM
0M/6PFO7qKBMCoqiahBT9GLVlXL0GzTrgcM183eBWU/CNzfFa2ZNnS1ufpai1VcZ
9Jod2KcWPrqnfzuh4XAeWk18ffOeviPyOnpg+cd+999oLiEAAMiHZOcd3sAsGo2T
qpC7U50qiKWJ9zxjgM5e0qsTUfSHF00YUM8vfiFaLo/Rp4QI+BwPeq+eV+Jov0jH
waoG4kb7mV4QJHhoHo+DJKt+lp/0miGWNCYSiXKfUISS1oahsY0jokC6ypZ5HSWa
22MAaRNw89O/RjFcHqOihXYol3NPe3lPsjGGzl0YetJUUUKDYfBcnFyfwI1UBBFh
8gBx6xjvDXmPFb9ydvysrfnLUifBkRW6mbE3vpaqRGifqZidADNAyV/6TvCte43a
FrIMQSbTzoabwCiMUhecsKwzjQD41CDRh3vaEAegM0WBSLnLihOT8p2wlf1hd15C
eYx8oEW/vtz/tw01qDu3b8E6uOZqhJmwMPgO6LZ2PLAgn96Nf0AoAwtBxjgnPYDr
HChIlHuO8uYPGaDdk5QFEDXqKPBWNGKQDTCOS0dSGXfDFAAmI2xwfpuHWy1gLQXS
S/EO1UFT4yIqj18lFLYXWi1d7GzghSJa7uikC++Ry0suQw/1eALlJwx5G9G4X1lU
R0gSe7qXI79H6n2bIwJBr/WXKlCdn4Xp09/JsM281eX756Ap27mlsWb9yNUPLRue
TVmjvmTrpJv0KF9Mjd3bxPRcr9QE1fa1JVGJ4jntdiMH5nUNWd9sBwcjX7AM35HZ
2PWCrIB+fQc72ZAmGj33YdJNKwBKwqIVNT7R27PcYnFER4wbj1fEqwtj/J6LdVN5
EyBYN32HKeK5dbh0HiD4Sv5PMKAg6mfI17Ul4jHru0I=
`protect END_PROTECTED
