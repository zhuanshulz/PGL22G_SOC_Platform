`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOJew62lkcT1i8P74OqGDoEIJ6bqHCD9wAqTvhLm+7V12EomfYrk+SKxPMEn8jWn
0TbPLHIJ1Kef6BXzhttNJ8lOx4guefK4+eqbFwI8kXoSjnGTOWa8ZE0Mo2fNATuy
mGABHDfEk1WGYbAMZWQ8fj2T15zUFCo280fkp07FRIGDyjkCK50xHShWzxPwkG6u
MEolwBNIeEpqAwr2dy7ijMqdwWHVuvpxa7e/z55WVpFFYGLwWLOE2+FgaG6fohk5
1PoQiRxnC6N4Fx6Gm4KLAoWEBzXdmic4nEm1ag657yLXLC2GjBLgxQfyv73ri8UG
sh7Nyh3yZBNAsu/PQJcpxZd+feoVs4Xo49KNTSh/q4JYF5Xv0quhWJLM9zUjUAZ4
HQaHRmMWlotDEHXwLpayD0L0hSb+U8xh+vTf1YRAJiVCD+YI0tuEx85dP9rb/JBn
XocXxZeX37V8l2TvBClgCON/GKfKEbH8aMRlLHuNCy6XcAihZFmP2trCVcxq9xQT
jKxqjVAfzUpDOfR3T3DaxotCTpGTWsPZ7o1d5PxVY98OhP6/QahAWmVMKj3OOGYs
+C0Cpeqys/wn045kuo379BJUwjLjKBP3fno+tl6EfWH+NsIe/6k7cG4uspeSk537
A5B4SdPQRpOMQF31KAXrJ5h63nPGwTzDFXUR0iwLmKL/7iEn6JgHC20odSHmeEii
8WRSSVS0WeDkIVHZ0hz4pdmuMwl8QxVJ1SK9JVfT7SBbUNTzm4UT+zIARs39dUNw
UBMBTHb8E+JsxSV1Ec4GoHZll55wLNR/aJkmotAKu9pbeIpR25VliHcVMGJZbAMI
fyedf5tzK7mnCJ7VCY/7F8exeQERRIRH34bfYuTeyLy4x9OmmawAomxEM7zygbED
XmC9Pn0cFVpfsGumvQ52pYABAiDYHfHL9C2wo73GDZU9ZwlDgfFcrot4ILdWUAOP
sKwXWtF//b31BaUaGU0uoAm7ZnTJI8SHgzaHcfYfuHv3DURj+/QehWMC15FIDDGw
PPJq3bU2gvi9T7Whj2SdIdaZPbOwuje1ynDcMpnAGt048XWHWMyOGoQYAc2SYANV
gPEOSbOv1f1ol9itv+m9+JrGdMg/uaNIJO4oHYVWFGQ0RA0ypt3F/ccP7wkfW1WB
x95RAFCPJiVh/FoKTahnV9rxMV/Rkcvz4uzYgrntywwCDN60XBRFlmZlxn6H8cXA
REMSUDOMCapapLn1G8JXweNxYbnR62w8JaVggWxspCcLbOn7Qntc2fjkjzvY9rFH
PpoKPWSAZIAM/OvIusCsA4rt5V9fN9s/M4fWNLVRfFSO33D51FPT25tYAx+d4XhY
J0N3onyYFkHgwu3O2HFZyFgL6uive+EQcmN44IF3r9ie+3wNbP9kqz/qr3/qvlPJ
W65e5Hf/BxSPtbpeFYqD72rHjNTy+SFGdOAc4WQiP/w6pdbXduZZvdrlG6MOF6/9
pMm1yIz181tp2TEtM9/c4d4MdViHCvwxiPw5graR/tDaLTSSXGuEwFAN3sUPMDKU
5z4WnLknqsC+x+mVTbnte8Z3NuaDFzMUm5f6aNz+rBUmMyRmMe6Yc94y8Y1nv8Gd
6xh7aZbMH3DLPScT6IIVrsojfBZeZCWOASP1Ym2P0ccDwedL5QTQyPFRQhwHqzU4
i/wanLG6k1nLYlSxIGx/NZZMzHkdN4U0xPMi9CGh/zDeOHftftkwAqh8k/vD+COm
BbZwn9VvK5Iilb8bBfroQKJ/BUIsx2IrKkA5jM2sbuR5VQqhhkPOEtUqYLUBatOx
v0C5nxEwpi5dhuof7hCULMCAoEwRnWQaGqqvS1WHBWTzd1qxrB4fRbSvjLocEuI5
VX+Rt2cLz/too2ZEsJP+93SoFKOjsMPwH8zo91veQx/UsOKes5xaErlTw3Do5s70
JpK3iVOj8E+MhmFick7JML3CCYCFsIF++zkHGlT2XUnGsHxwfw7Ehp2+m5j4gFOn
pxJErkWxmoeNxswlo2dEQxLm0+xvpTTAa4Oosg222yaCMxYJnJqlRphjWxXWA+Ps
jfLUgP4gtooP7mo7QkVBw4oPloBpC6iJult2XQg/4Rr+zpNjDJtAWbpUekrPDcBw
E0YW6qVirEYZmdOwhqX3R8ISVROWzxiWnRUQJ/B0tsHLpQ9X/1okrJROFtGKYgJv
SYXnmX+AL2JHPAr/8efNrL277IHwAxNtg0VXbxIQnvA4BO8z55N12TK7hBZK81hp
IZnYkthzD+GWUYN5xCqGWELRnkZdYEblJTHoB3TJECfO7scdA2I9Ain4kqOp8xar
x88j77qGO/huF1IAcs2DquPVmUtJh4Imoysug3Skj+izmWYS+cS/rCpQARe1qrTa
9ilwIdRKznXIos/AHXz+UHyFtfLA7TpqWXaUwH7//D9ui4Jo2LNjF0R6xVGQDg3t
aajqkG/xyBeny8+BTuErq9l9Q6EG8xyk8nlkd6z4Wbea4ToTs+tpmAtSvCVYwDao
GCuskyaERImg6ENXjVInXGWCTcqejwfaNNwZa0TRCb3df/VvOf3owUqYhCz6rRau
ETcOALBbblhBMg54jWJr1ABHKjkMU4xbxuSa1flerCH+pAUyybtw6MpDryhPrZi9
9FldGDbtviMEoa5AjnQrgZht3GsrOdp4oRJ7BI+vls39uySY/Y2CcFrG5EVCfySL
j97RIWoykK4YrpzvKgzwAMMa56pW1p0jGyFSZA93e5p8DL7HI391x6w321USIyVU
bdIL/HqfSQwy4K0AZNZa4i7eGSbSwDr5Y66+UKRSShsrgR1MSkta3Vd8SkxWUffz
O1Sn0A3A6SFFE335J2VNnY6ePuDZNV8qLYxcA/Bjpeb5dM5lsqSbHi9RZgrv7+6J
8EILeJd3n/flwSfiBMpi3O442jvPDNqhg1W6+je3bR6eGVS3I04nvI9anu4iSAp4
lBiCosSDcIZ80ynKnAQDNRD+WkGrBb9FAzcdTXLHS556X25qgT+SKt6iDAl85R1M
YKeXqhAUT/DjxbRGYcakHnj9NQi+oG+kABtOph7THR7w+kOTtEUWt7WO2vmXuhbF
yyLX2JnKL/FeVoKN8idrNN6eZNk2g8f2G8U+/FGb4FdXpBigjwmo6JK8tBzMZsFp
WOzeygprrx02svvWrquMVLrVQWLgQgMKfdOIGyTto7oGk8Mndp/JiJWf4Bokpyde
D2tL7Edfn1ZoFlSpL+/dZrgXUiRppLUs/olDb7WCWgUPZtEIERG+dqgxkX9EsyJ3
HxIY8YCXaGrRJvyus1poj93k7pP5hbGYCCAqWMfOquDNPtL15Ma8kvBy8yKBtg7T
swYO1K6Yh27u8dqSfmEpDUFqugpIlF5leKpv/k+dT8v2g1u3Bfv2ldDq6QgtNZNg
U2zu96+GYAR5rlAd1CHZbgGlGJb0jzY61oP6CVqT/2yewS+tzWQGuBx2GEROaWmv
sI5lIt01Vg6nId+we3XTl6YcMI5Nad7ClDYlLuK/aqjPcyoNzIQ77R+ELmXlIjYE
zTbsE/VfWefbdFKLz4fdcsYWKMv4eNNhgAJk8s4pD4dw6kDkTFJMFzlGizlM80Jx
hbdLllOMeMj8kHJT8nG+0XB50YDE5ADrOwqsniTeQ+UFD+ZCvN+/NkancNpyaXf9
sIGzykK3bE/XHtnWBDgJ1VGbEbQhG35vzkR9FVGWm1vKAZFTI7IKcRbkOlRwKvnD
4wKKgSeozPZFZfu+FLq2EpjJj6IzDykRssDgb29wNMBUb0osL11eAwdqYNEHPDA/
d29vZmwLj5fVq4QDOuEjqAV+Al0IbqD8AkQD9ney71ejShphDjLwpv7csFCeqWoe
HRfSlmm8i83LqqoTC85Iy5vUXeaPdPB1sDUcppTy9Lzr8NNp9Ae82fE5SvVHMQCo
L5lvyOObgQRE8r4MsxvxcQ==
`protect END_PROTECTED
