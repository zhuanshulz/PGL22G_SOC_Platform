`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E1zAgLPZt8/wkxEigKdKfLFBoHVhSQPpzOutggUX5qvGnsk+ij10rlvtqQeH+ZNs
h23aoH4/dAc8Suw48t7ItU+HawbTJTE7qHYxeAlRAAmj+etW9mqSZmjwxiqtafJF
iBQ2uo/4BRlTQrOCebaYbewW+MriYBWVKxkapYxzLr+d8rdIpy1Yb6B+gF/kDzNp
uBfb3TPjApccEsogxZ4lS0wtV+/sSkumdTVVnjnE3MSYr4BbUFScdgU6Xsr9XMhO
4mfuRlE/SQcG+6yrTByW+6TZmnbbPUzinO6cSB0KYx5am6NNF3QF3zzuAlaRRhJx
5Q8OU4mOz46kGDbsXa2rF5UMsiohhIh5XHpwCs3CX31vt5bgRzJJ5Z+lcsrb0VtF
WGz4Z3QTDxtUMxv7AvBvEUL2UnaChargh8NzxBCZOyniomMmYKAzal95nNkm9jw0
iS9c7Hm4ahrJx4dI+5Ee4l5917PO67wQAhZLLQAs/mjqDxRAb8g8JnMDHG/b32LS
c9Xin0Cfziy0dTScB+AcMNtfW22IKYA2OZYPWOqgYTG7iewWBl5bvCk1BInip2+f
BTb45PTsGraSAG7epjCN5uILywoNzXlwrj8JpwHGfaZq0Qxr8mroOBctaISDAVhE
hoHTSnIQLMWTKlmahsLee7uP4scWHW+qG2jlrywEo9vUnRY4XegVt0ZNPF7UnUSc
RHii1KDkJhJej/0RxFccgX5pSXi3Z7wYVujWj+N+/HLeBUv7UkOzMZHCE3xsEuDs
K5i0kZ36ybc0kBhfuAWuOy++Hy0nFFPHJ9+uKvUNzs8Y0yjbNidiEYTNu7sUL40k
FqTNjfMsDP33S6Xs5Vmo49vgLIPtYoaJ+Na7zIRBAIHu1Meqh5nJ7VAu4wMcRGlU
gJHggiBQeTIYRKXZx4/0gM1QzSX3lJGGQAMbizbS76r+ce6VYkX1U5YunhG5fqk+
BJNn6SNwbg6YDKQuCpkpDghyiHtEMyIUVSYXEk7w6h+G9HaKkKkgWR/nnf3Fjj16
3yIYp94cAn0zw4ge45Mjzuni9zd2XzqM2L443rks6RjwJag/cK+0ldkZ9Ud6YFxD
8w3Z3Sx4jQuE7g852WMRceLE+QSwDsQPpXTgfMCtPKoJgeTlfpNVahaZ9DLs1SEB
Wo1blr+4f4bQ1bkTowQfSJIBiQNwRk8S6j7+OimrE3W1z+KqG75Z1KzH2UPYqaOv
Od3bGDCkkcj/ITaBxcWfdy//UPJKGmQsvRCHgMCzGkOfR+YJKGjzEAblNdHWCDrR
IG+FrDWVB/PJgivww3Bp1d0FUAum3QxfW+ub72Ddwqs87KUuzWXYgp4li0Iauphr
qCvpicdr7nhnw/jMd6eSS+9w5bMhRT3/pONfOVHjtuNPv7nBwNfyJAUMsCPLsDj8
7PAidbjvjkstAT4Q9YWMReb0wKxdk1VMcaez6smCWiK/zKNJKwhTTnZvFJotKrbb
w5ABTuZ2Y0QScerxYLomy0L165GEdMVeCp9jgUIJKboTnzpMUPcM4d4rU1VOh9tV
CLxVg8YIREl26MlM3Q7/k8k1cA35uVkuP1Xi2wGnYoDL8AxKpX0aDpyGffz0KOm+
Hjpk9hThFdstnVlxwd/asMpFYpCvr6yj0uU8HOjydRtRn6SBC2TWAdw8CDFFjkDj
3BdNgNTnRp2Fgwc09PDSrFwzKiIBP4oF/IWsG6FymDuByAPzfJRlhlO+plCzqVEg
pD+yEhZThw6H8GsAxogpChaSDmKr0EiS/2yZ7ZJZ6wV8iF/kn0D4yDs83Fn2yJMB
4B2bVKBSuKkF7Yv+OvwrwU/UatB2cxCtodUtvFHq3GfojS4xxp1upzMKQJfFxMfr
Cwaa0iQbqa+NjLs9HGvllU5nb0aJFzVmjdoJ1nc0XSNVNT2y8OQ/3OFhWGWcug3w
gWE5EgxudwycXBr3kEEhWsiistHE1r0EIgDZoSr9c+cyWW16d/V9mFwFYXY+rDLl
e+U44U4Ws/krmPWn/S7oe1YGs8zZIfHHG+o0zLGwWHDy+qJjlZaAdex5oP2X4gIe
mkRxIBMfOcq9KD5u8hZJZqjHYofA4UaSEYOVKG8IxYY=
`protect END_PROTECTED
