`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iUsNLPGMwPeKUmre16SYUf516fvx/NWSO2VS1gzFG+qfLppnqG3sNanmufQgPRIC
fY5oNnxuwJgRvdhIQjvOXs+RupUKLl+Eif7H63kYVYd93a9ZlW/Xp2SU6CyGJ7ns
nruFynEnP1+aTao5jynHc59M0a4EiAZKtww1cPiAxUir6qBcr9tsRgFTGHWtZs6R
DcnoxZ6GZJhs3l+3kM72dhlG73Dt5Dvxj37tuTpfim3AzQ2iOhZrm4zUyj1ftM2b
CECxDS9z6EJVc25rACluH8gGKrsncCURTNMKaHeN0AHcdZY2eND97kR2ucKMsGII
Z4oY09/Cml2wxcK6YArI8kiPfHqPmS5RdZ1oxi5gAcpYqhxBPqW9eh84x5X2c+n0
68JTzHweJpIjk1uvM3tnAMZvacQfY9pnWzHA+AfbTeO3Ye4b07CSAiQNlk+tPO3H
D4JmG/Ii1eWS4//P8QYfk/7ti+efC0v7dDlwNCe7c+M9SMkSpzPi8/J72bgWER0b
qTCRlZltj9E1eamL0XiZxAyoIiDAV0Iel1QB5wXfARgVwPuzLb+cn9TmL20TSfwK
68pzqKOhpPeKQq0EKez9T/t4/XCZ16/Xn78rSHJY4GwoGbJSSGgeIzMLUvTEfSor
+GXZ1ujkuk7RaWJQtN2O5ANZvA5Y3SoXMr8AIky1GUdCUlYgo3ONJi36wPV0q8mM
jy15l8A4NpO6UvYzKnD/5K8P9ushhTHOLcEoPpbIu+Jn1iA93kyE5pCqhrqfb2j2
iVzoaBuNPmaFpfOts3l9HmGL/s8I9ZnHcLfthzgqlgbodlocPz7lm9PztczgU2qd
hq79+2SSKz7D5S6mHS6yQNhljSznV4mgnOsE/vVVhli/2GG33HwcHt8OLahDfiUk
jFTp9tiYdjYym4xDBKwKNFPGdNbxU/6XC2OkRcwlGRo8UxMCiSI9mJSfGzuJxu7H
vuiiRJdrRnPit4bznY71hF5g26LP52vacIOtZTUGA4LykErYtn7GqUA5abkSmpsw
NGiG3Xsiqng+86UcjFFhuFuzPj6h7LiSx4/h3nPBunjv9GZMwDHDQ+ZbGYC4gEdx
WAHIqW+jcfm5kY5ZgJ5R4kRkSyYRNNpMEKnRxbZX4cDkKj4ZBztBOobLwwEWv1ye
E7QeY1z09c7iBQEAMUIZ6aZbMctwaV/HXg+ixt+7FTAROTzkpETQLQqbOgNFHJ9j
AXzvh3kHvEpW6J+2lZEgfU1erm/iZof32XN9Stzjnusn/SP5hFgEIxlmxrXv3neI
YV+x8eEfJUmHmmekMzfCFDb9Da/9I9NGbc0kvfZyagw885sDdmpnYR8w6RJoMb9/
1v593xNTbfOhPg82Hs+zt29PyoOxT5ueJNrzCttpebO9P5v8z67DXCyINB6ULgyf
MWsTOs/+T2bVcjNGIINi+FbqzDUiUaWlqYr9F2zSNuhdxpkePg5eneTHH2kw2x3s
2d+ijGaQHaC6fPqtvFBiqIZdkauMCGkrFQfZafEKQFqY0unL728mIMM6c8JdN+cL
/xHwuoaU4qTxyBSzGXUTTPw8pGcCy22Hm4/WOZ7Brfnr8Vro0NwPHi7ZLtuVpW4f
Ql07dlj+Z0ptgyZ1dBv5mfWx7ZQ7J8vFBkbpxxDnZ3UL6GnAoB2G5SPqnSrxhmRu
ZpmXEL2Ih1+LagoWGvKHE2v9QOK3Mgt3aNnKnWTaKyCcjUjgUE0fsTyZr4A9oYBt
gfkpLtinZWxVhe5/Obv/nrfhrUgDaT6x9GcAThorMBHKWfk2VhcC9OgR6riG8LYt
OAZwT0TIJcjgX3bLC4m/57R3m9Aw1TAJszYvzu6RsCmOaxFtzn5ORCQTvDL1RORM
gbFH/QbfEtGra9ZQICoYGg==
`protect END_PROTECTED
