`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fPlHU2QHyv6Z48s59eUx+AgMpMAtc4kIe+EkJz1cxo7fgdszW7YxT890Um/kK0W1
67yeE7dYGN2FuQBUg9j9gh76bnDFd/oQDrI74fO6rLTv5wxgTvSI8wW30x9JNnF2
8zMuWPtgtntBAUQZNJn7Pmy8GheuLt6niBPG9nx+OHbFKZZAlsP38hJHetLXuU8b
As5pZ/RyUmDpwVhW2QWa5hGbOLwUrKsRN7Xv8w58QN6/7Gq2cnIt2I8X0g2njzHI
HUQjX589Jn7NPtVZPegUHSBQiBdqY8wY8GbOuxrabXnq59QSJsX7nTkLaS4mq98D
XW4pGnBc9YNixLx7Rg4R1Q33/A+V/X1a/KDNdyZKDqRVMZIhyhu93zc72AX0T7wl
6vDNonZ0UyMojrU9Sk7As8DSvDIfIsqlqLQoqvbzLOUcjjX3tMCIZkG8bxSNoYdF
5PvUuB7eEO7cZVtnFxWscuaGTSGA3PLKYm3WYhHFyCHZ8EcypHou2ByQD+TftXBU
2V916aDKCNyGvNfu2EtNm3ZctadpEjP/+gJ2LL+mlA5oB0SI+nWphYec5Nj0QN/6
/gZq9GB5YGwPFQ+Wq58VjlBS2xXcwKknaDJ1l1EGpukbkuh/hM4JLKWulTYDRar+
`protect END_PROTECTED
