`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/GInKJ5UHBG+XlbwpwDGm6+hFeuMKhz0s0YS+9xnBLfsIN+8836cbOBNH3fIwClR
ApmV/ZvolLpTaUF+2re7xO8/7YIfQtR+p8zx5TlcLG7g1dYEzxQ3WIjW2+h0dQtb
Ggw2Jhi3pzV5RcIcOgO5zTuKxn5Xv+aWU1eXdNXrKYQ0MFPUzqcd5tiTwQnKt2rZ
ZbajkgGSLN3Devq+jeBG+sJm8NU8hMonhLuEQPZEYgKOHyYMEf+QPOS3L1i11w7g
54EtMQZB3UsDSNP3DH+N0PRLcsf2GEFgci94RZS/XtHuX8hXVJj5q8eY0NuBLfVb
TcY0oyycHUP4gny8ig8CeSiPXh5vEV1w10BtfOWqhWlSYdXCbPPitbVSPsPhF5qe
cP6pjgsfp+BQmR4p6j8D+m5i37ZWyvoYaRKMZObD9VlX8drPxdhvQYt1wJyg2ZBv
Mb86FYkZ8Yq/iVXizzC19Q2hhRSqMumUoJrm6DYbOz7QvvnCmC94NiOrP6kroDEk
K0k64q+qJplSEMvU5N/UmyfjXX88bqknnfzhbIjDih5BnhYcDM0KpTUgBBlTacPA
69QkmuwwpiAlFosH8luWHvkfO6KzX81vvI+fadCyCS+UHJ5pG+8UizUd54j9guj2
pwHQh0wRChYAWfS2C3eyMn1iW/RrRC1Fcu3V8ZpGOIEDee34vrk+I6U+WjBN9c9O
sQ8lZC73wpBt+FaVAWBrpe92aTSZ/n8E0qt3BzcmuPYIDh0uFiIHYXRBLCrVpr7s
4IgZts4pOyr7NsEtyxYMSZVYpI1Wh+vXlYk1dZFAM4KUBZThwuN5Hi/bLf3wl231
V87W5bVDWSKsNDNeORzdmFIcOqJfHsCOjrKFhR/x+9yfyxk8B15ThYBfIIbhUq4G
RVJ4xNkbC+Ud4ORShpgAqVi6ks6HvgCFirOsQgihhuhNW900cPCB5m2asA71L7Lh
AGoEcsnYgIFJr29ez6wQ16XxbBCL9bk4lB7MqMW2N9GF6bocHNVJDWZmMJJ2LXKm
W9BnalJ6LeXkpPtNnQTtLA3ROcT89KTYlSt1YiM8ceipssIBs9WcRbCRohDmampQ
2KbUZSmMAA0ezNwAkv53fv2pCLPfFoR2lWJI38uvOPr09FNdwKKvXliPHPZRZqzS
pZZ7Pyd+CEODkuMkYdUl+77HeHNx2E73d/COgx2KSuFkWxYtXqhiIX2wL+TwRWo7
6QDx8umYcy38Ort9x+iKpTxDhG0an2dDv17NOHHOjC5yYshEBAZR5INi0BVCwbxW
815uh/phnF2qoOsv+ohKS7lG8cYRXLYzuwLQxto8u8sJNz6AYw71lWJ9Zr1N2hKN
zoyV9ffa8QTOZTdvBqP/lvPQ9afrBHlDfEk8Gwrv716Y7a0bLseEeBrI4CbljP+N
MKNfXzicX6UQ2HiSmoj6DIzrXsPBPV66hnR5QLeCUPB7Kh4zDJnAtYcjgOznkJwN
gAyypZowQ7UzsHq/ZXKTemP/yhyf8U3JcnWbPfD4quAK4kc43pASxusYtnLfsPmD
k9ivLQ7jKt41Jala9Wd3U0QsD4oAB7tlOdgBpEOqF87mVmLkOabneRiu33O4FX6A
YX6pIwXUbTjhI8cFB7VVbUe8netOPHagpXNTchEnWDmHD75cm+mD6rei6g887P2A
TqNmKEzVT7frKw32iaQk+NiI1yH1TCIDLzSyCbyO/9eEVUj18XwrSmoDRU8Wrkdw
jKueDrfBOms0LPc8F1DQcvUzLHAcl5KZpyJMkcDJcUIKsCk9xawCTcmrMzk1WvFC
ZjfRkYWR0TrAVH7AfGGqJxllr6Cu47NW4vg0jC8/XvtZ7RGhKHUBrykhcnKUIF/X
18QwensBkIeUOfLyjvOkrcfp6c+wYfkeacO88DTZIY6FhuZ1GRRNVkyFp8FMIM8Z
qmp5JY88Ofg3BU1Y83PyA7QzRPIeeBq4ITOz5IozwvuoMRBASZlHqxONwZDM5Fqe
vv1ZjKzou1YhYdq+ObABSGf0HCRRKpekQa/ktm7Eo/hv7SU2pz8EXUvht7dRL5Op
+QZVfY4ZMazH5aFpsSgVGl46udAok4HqZfPjbSAWpFDnVmLHBI0TPqDe4YU+ZUuS
nNGYqlITuEoE9b1AKUhhQ4vKVQkXm9akn+uInMNnE2vOegakw/9Vs3KqsEMBFr5h
kGxWOYyloVMz1EpnPugDQstW+OCsQlEhoFpK5R7ODlK9r2TXXD0r+Gelm/4IisM+
8GeroHjTfvFRxuyWROYpeLbXkYlgGJ369sV2y5OqTRZFu9062XPMOEIpbA7c45Y3
AeZBqdj5Hp1kQSjwm3W0YSWYskqoWBTmBg/YIPqK0RDyvxsFAyx40D5N6qZlBCPB
vMbbwMl5ZTQ4nFTiz5j0RCgngA1Bg8KPEORPgL0B0JX1aFP5edbRh5t6N4iFBHGN
l3GkgYMjfXH0gEw0AlDNbNwyZMbMOY7QI4UuwICT+M2AI3yXqRfahP2hmFDRc5L2
j06cicqfwSj7kuv7gN3K8eInuwIwaTvJGCEo+W4TfPNGLnFut+gsWidOU/8AnHX9
KTjUGCjW5KTOJMAXncwn3GU1+f+3sZqxqTmXe03LYbrE8R7tVtw2NyYjQOXAwQZO
w4ctcgkYF/zhf8rYeccb4lWqTApNfymGsNqCRdXabF1yTZYun2SgjYMYyKJh4FlA
V2GZ7VjfvihknRklcFG0Gw7zyF4o+vuGXvnoTwgGQnFyMvISwhElSJfkQnTzN+it
F4pPgHazdQZr85Wzrd6/vQVjRHAHX0XRGmlmwMCvWH0zsNZ7ad1Ise9Xg3asGLth
BnFlXFPPfDgeCgPTcSxBuMdOgPmZBJNFRbsYgO5JLf6TjxeX1373tSsI9US/XGOb
77ipM4KLPmqvkRLS6T4RvIvUrK5yvpPmMLL9coZF07VD0v/ZTcOEZVyPnIysK57F
YsBDjlNgClmuNEQhvdEUW8BQYOMu5tzbsF8VOMK4jouunzBl2QEy4lrGhSqRmtPm
J42mcmxP3MGzqy0kCLunJkrxzLDG0nGMl6iqw820Mdw0K6NvP2iehGW/fNT5B4iR
y3vVDBi94siQcnljUYwpgQjAnCiGGtvDydWW+kRGkZrJuqOIeBVLaIFUZEtifz9C
TUznk4VEVE9Uzaw5T7hSfzg2CSgMVK/uFvMw9LgS+39Mv5kUhc2+hUulBXfeT3/z
3Rf/EsdtVbxq39i1JJC0mYW1IVO1sbuMkGaJPt0hxv5RF6gFzPLGKxVfxYS9aKJ1
t3Hj9pZnvPFr7pBxd8tfH9EcF2vLaptiEAvCxUf2V5SQ1IjD+8wTzXiDTgHqZy4D
ZnHLpmb3u6CWQ5/9Xe5ETJlvbWJvaR7SJ594xN7dhQoN4IcaiXIlXsFAtM5JmV89
61+9D/3aQ3bJj3DHdnv25cR6A9H5BXh3xwlV/jRlVz6XycEpdRpnSZexVBDxl+ID
Pbi/kk+qIIskGYopxPdX6iGfr4POmlHg7gaLTJzYN3YaB+uZDXelAFhzJ2No/Df7
OSlCkRF5vBQzzpiKJJR1SR8J+D3l0SVl9bORolsvUj7MCci6/158naAxno2n1E1C
UMNkGergyXo9OmtAtA8AEA1ch2bcStx168vkEfsanY1bN60LgIjm/TJF6b+TWRw2
JGMAN9zD+byyYG0WkS0XUuLDexRqYXaOxZTTYSye7NyMsV5oyE+7XAMS1n2+KEXB
kEz2c9rpTzMlIFOSUfn00+8IiFi3yELJPgHi+P05G3B4ZtVI5sZVJ994Voo1W0qx
FiuOrSg8icnb3bR71pB6oP/u62aEOTuhl9dRsohEwOdQ8+vetZLAlaakUEl9I0Kv
hNBdOaEMZATQFOLjOtWmkhkFgg0u09SnS/3KPqvNtEzJ6uQCbm33r+e7Q/rV3n2B
H3Lt0GOWWbe6TDCQKyizrL5x0hSoqMGZnXLGzxoYN9hYyY92M3krgtTYJvyZoRDd
mWcs4Vhna3nXhTZEqcnVqn9qNQ7mV2maOoT+pVoRmKY3n1WW7A3UlKPK3rFHPR6Z
CgVSm9TOCu680rNVyUtFjpckcBbZxVCQXm/y4LmoM7gubAwbJwUWZTSU2VBuQIbo
L7HjIc8Q7FSV/rMm4CrQ/ZEECZIhW/TX8rXP3BPsjPX6tfsBsUqEDKhd2RwMQ7gk
8BJ8+ebmqa98iOkbghnzIAEco4nYjtP8dNq18+XKl9CHZlpIFrlJ8tkHeWHerqSK
D9RrdbbLRx8evB2+V+7Zj0oRGkhwQLa1sP0/nmb1UiGU2SnGhajBdbKliAH9yupP
iKHBkMmsxCtEZXua5XrolVpWvQqR0yJHO36dtaW8kEE+uv+gjXFxSWGtEXlarnVX
YO9nEdbOA6ouw9rhGSaVsYev8FfJwhPq0ctf1br9gRTccORETmfqq7k/Qul/lyXP
9xqAFB+NzJ/nCb7V9XmY39lF9hPaBUrWasSq1ry2P7cV/l+Ta2EAuRaOTNxdEAA1
+4Qs8yBlocYTmp5BtRsT3dwXc2bnIM4itZRC9idXjN7dhJCNgoVeDNJTaHlWs90J
S8IPJ1bwJVhHjEgSKHKBJjtKxZBU0/1KLKhtYM3DCKj1kB8rULKV7nzSK67d4qVd
tM9h7OTsBbK41DUh/owV9w8USUvKXMnh2OwhmNFQHpnBf1Du0VkHzyFy/wM+qAez
Q7FqjyNt58AhDdoCF3+h6DSkvBM84G9na4FQF01LWECXzZzq7r0Szo+xuXVp7PEY
2OpT3IGXxSLO/CKgfF6Jpl1TB90Quv02hZ7cxGtRQ5jbfdV0rUiIWj8nRNf3Uhod
L2RUkXIh6vuWT/JqAL8Eecwhb6VsAJ3RVQAoMxkqychh/HKWYt4CBHv1LGWorrJT
vPv98Cu613+kvEayPXxBao7Y2lplpPe/SH1/eD3PNIKC0XULZLjS6iivmd3h+c2b
MXoWwLXhfr4ow+1wZ/+A51NrWWCeo+No+T9QM44v1NRO+IsmnaUM6AVc1GKWt/H9
8tZfsRE5RIPNFRQfV0OE1A9w3E7VKdSgKtp/Wc6gKA8Ad93yWAvbXcoM8GL/MYkB
wYG5/jDSYCF5AXLZPyCrV3r2/mJoKT+M0RyCqsh+8wKBKhm1C1oyRRcBVsaRk1ET
WoliDEKgF2toyv/I7Ft5tCGeBczbCumpknLQt6wgZKOa+25qgkQN65HG4A6HvvhX
9S5YnASBJvjKdXA/lmybT2tP+dHTAkSK916z4qQfOZQohei0DkUgYy9Jt2CZoquN
WoBfW4dmtiXh9Xxlf5UxaYwnWNVFUPdWmeVOvEHkzWDUjJAubiP1SRZFARMaNILK
rJrBd5SXNaPSREaPhvkeS9kcU8IQ466EtP03gKFYn+RJ7jCKcpCdSOZrI3NZxjfG
LvrsU+FKfefhynNZb4y7IdXtx4SbfWuDh4rRcBq5qH2Rwns7ktaxrAMaNZh1jnY3
7KXrYfBdfqv6AKnC4FSEdC0CziCTGO4pZtFDmnDRJR5qV/YZBN1NFi4oCkEOTyS9
6pcs1KCdvPBrYfI/uLdyajzwxtx+V3P8hOmCa45qYK+P4t5kumPT1WlYv5bNrHmV
tdQiqb1BDmPHFVKiNIIsPEsOiWMRXJKiXPbprwTPsXYwLLuqGMOxlKMEgUNEhALL
9YQqB/4VeHmQELt3rM0Zf4uUa4x1rtHJHsSHK29ne5Wf+LMQbM6oQ3CLIjgm3Gp9
AQwsN/Jc2SywhoPn63+2qU5mSHOFhij1ba2Hq584+Vkql9azGkleE9+Sg4AToiKN
rWUOjFWw9zROKff8solbC5oy6vD3CHHN1vAVE7EYau+T/Frn6LN08PSiEZ4KGmW8
NaNlmGebjSisVuyTO7Zc7OWo6UE00GKRV4kCOtSU4bgn+NbObNUtbzDSqunA7Qqh
VjSQAg6kVUH9Rbz18sS6/m8vn5+DDmjlh6VmDQs8EtEoO1wjSdyrgUlQNs3sSxgL
3IfJKdW/KUCp91ryJovhurw3bDJXpdNO6imVp32Oqv0MOK6vL89Z9Lxaem1bvNvB
YFkZqBlsIcGLGsGtw71Gb3RZj2IkL8M8zgw2u5W7wtrRIhhxQgYE5V9THeOGeI0h
ZKNrvblhZcFHWqwLpv9VSm523qgrmhair6C6tIbjKnhWz3ozeHkR6+p0ujmmKECo
prDTh/LLKwhhMFQaXAw5t/19Hi3PFFNxaD3fbbZi4QaNTRGh6XGYkl6hxjz2VMMm
A6kLhlPYFO6D+s5Yj5TVz6WvG6D3ToWhK1ympbh8NBeEYiQqPcwt3ApkKNBbExkf
aayz42blMuQnbdQMMTfy7adSWeXTZRSLa3F53ujuUihJng1DQc49JVAO0SFyrF3O
t7Dv9L+inwgpz7nj4MysCnThT6odkOy2nq2OvGxAeVJfwbQn5NaDqVJ/0szGwmrn
ciXSfMt0u7QA5jSsZFzySqrio8xSy2y7Ko++Yqq69YXyLswX4CvA5D6ONjAtr95+
Gc7ZNZcpq1/VyFDgp/w4XcRUDSXuh6QRA82CZWRldnGiZqTRxU4KKYnZgtwK7ceY
76E7XfgLl385Tk7HHLIA0u/ale5b/Ijo/3MWrCx6oQ10S49HlFX8mexGRWnj7f1U
pF9t1hZetkTBSeA5gEq4zeRUSeV47tio2wYydzRuf9DM6XC4NrADsaQC6suZheiV
geohnLgPxIdRKzGq+3R0L8cKndTXbzNOUc+s1rocZEoRkj1VbSjwmMQblD9vJFCX
IucwFyMGHIMHKfOQ4IGV5ogC1o9nO7C15rU1a0KAhBInwIBVuII49Kq8jNZ8im0c
eUqzNHTQwD2MK0Onbx+G93ka1X/t7OnEft77uKLwYv6sAgMCftS+axgB7/tSvce/
N65zfQaryAUoiAzYd3GfQbaUNzQBm0QB+Fhvl4ooNKjbEhc3hMBxFPsd9iMPa3Bf
rImfVzlDuOOR8MZ/sYVmFG5mT3UAo2bsi/MIHe1yQjIKsDy7Tr6dTZTeCSzInHVQ
fuFOwc8MUbAIJIWZF2LUECvtfTjWdu8p8qJn7LNkRZ6nI8rNBmL7cwbKBQB8BwI5
jsHP2bQaGp0cFhnMukZmKfCafXqwcbfCtgn0uwRav9YHWkRSYzEgDsGJEpsKpI/C
8WAI2HNE3cgRxpYVXds03jGEHQlfHPPVKJSHZmiBWzKy0382tqJOFGahUznahbve
Tr1RPwRvQ3aEZkFEpGYJd3pQVUwqKUbtxmZSV1BHODOWJ9CsBleAtMOxNdHlSu8W
l/dxwZFYkPRzjYVLr4OlpgxCbI5itEAZW6Tm/MsjoOdMAkADj0ddQqF1Fu/m931d
F3jUECJRfg+yPlWe91qpHqNy7l5m7vYBZjIN56QJyngHfHtjZmEd8fiyQwjhtBJ0
mRlVVNCLmgDAyr8PDNekTMyTJaM9OzEZhE+2UGHa81wmHjenwBhd8Q3siibGKqU6
hBlgQpLCXjm+FMIoUBXmZ/t+L7r5LSktj6gcSGHMbmMr3TiAuCapc7yXHU1vEX6u
Z1LUQsE3ISqTcFxGVqWdvhMUTTz0Mpd8HoSGm7YxMjXRfnf00NAHmnrv4yYjHC/H
/QTi7My6x+Dk1NSH3ILhzu8IQYZrGu8uwf2Is+nR9nADrFQ0xFIY9l1YlB0emyiF
P1Vs9mfvR/lVVUduigq7mqzzcsZDEW5a+t+h2BaRMdDVX4Crkd7f4SQ3VHNaa598
pnqK6GAj7+QXDYt9y7Rivvv3Uj2kGoefnQGYfwIpmA2XSSj2zX2MqlrDPO5d/+4p
9wBLH5jAW2DXj4n3wsC1GW0muav8J8lHG377zHPd5Dw2Mh8xz4I73DRjDxo7rUud
N5KgZFzbPWDaUa1KZBzMblFuDagZPbMnGl3fAxI6iHgjSpLnDXD2w5mpxQN2kbxL
6rXHt1yYkzQNXDmuibIZMA1AGqph/hlPm0/uwD2A7IgMCnuaxlv19blYtphtV/4+
neDDKnsITqI92kDvjKcV/OI2OckRlkm3hNfj8mq3O4MttKH6c54pVCsxbAjeme4e
9jfXWb4t1kBrivLrrQr0zkd9GnnLYeMvdC5VuMm0eMOyLwJh83Mp51BL9gXTv3iq
hE2UJlRvRlLxHqeEX5SveJvivHGWI7deWSrvPAOJhiUWsjQuB95++Xom0ljoWviM
UJsHAJDcD5S54XHVQ8ZRPRp3UX+TurGHfyaR0xzBpOyrcI5SDvhvX1HioQvLGFXR
IMA7wEF0n42p4cFxdZ7b0dpMD2KqnmNMPgSG7srVixkLGutENQlsp6FurmIuUOG0
b0mOjXs3oWNwQjrXHbTXz5RoMbVyP0qN2psJnzZivFqeUn6w3eEFRomqI6wvs31q
Z8PeprTwR+/aVQJRqhj1y14JYkRz/ZCTrR0xMpzCCRLwjBZsAqhsVw5eBGwCfqS/
xt5B2lsSspzd4ZTJ8p4Htij1918Jq0J9u8UDLDQhN2JgRA6w7N9Vzf9Gt9Jk2goU
yQib44hdi7zzUfMvTFjZ9bMs8+gXeg7WFer7Qaad1UYKmx4iNxQfCDZ8HKKj4GYe
EHns4/w2dPgLV3Z+lbm8MXQp+D9bdM7dH7AdIfY+qLTLAHDVqxKqz5yHUQoKKoKL
sTJVX2usgkpP5i2LnEPUd2wdmRsF2ItVYKVSoZhyqVktZQ9OB3YcpHJJ2fwez4Ky
kp4ShDIxlfMhH4DmUS7+h2PpPog3EBQqw2WlBNCzlxC710ztfPh+anH1cxE0Xod+
OGAuP31s8OJumRSH6qtfXW0GNj+VNwUkdi6DcLu5uOFD9aColNCeENPcfCF1nGFL
CfZXdPoxQ6P5h7ZEnuAibQ6h37WnMcZN6zj37nDFx+nujrpNvCoZ/sjqcQnpFFyP
2a5bjyCeAUx2L5eODP/F/rbEF+i+FMFTUTKRJsK25o98MkE171bZ5mWM/KqqLor4
4rolIolmyXR+aeDrDqt9fyq/+c1MZccOJ8ZB2A5WqAZzv9WWnvNYLEihyVsOVU4S
FZNhojzd/5Zi8Box56YqkZZT7JfsYvDBjON2OxktaMM8FON+73PYCL1DlPC6/i0j
9WJUSyllwQW5KradePcj2DFyEhqlzQRShKLT9MTb+NochKL7NpkC8rFyzoHLKHkY
ZoFodsClOLfPybKUy+Tq/U++iFP5wMwiADoxWn4hBuu3AcjReXvtJ4kC4kyNxYOe
EinVv7trgo+lGkhtC47LGe9rGoDNmk0PEwneCKtx6XgvCqdLjbpeNdE9U7QmqbTi
BXzSGzSEF7/LcQzQkKIiVHfjhWG+rqrf0yzcBLNcxj2tv1uVMZMDf2Ft7iXCt7Pe
uvE6o16QMWRtetK2Z6kvlwU8SO0pmjUMibT1irhNjVdm4wvz06+jn1z9xehfOyeD
4cTZ2LDSMunu54NKul9LqYOUbKBjV9gmn1F//CkJNxsJmsE13DKSOggbvT56lHpM
m7F1UtP5k5Rai3p6VsbNrOaDyoyQPO1bixn6zVKM6aevo1tHTP+LBy5fygHHITH/
QjaZqP5ECMCjIt27da4lwcvvUDkhCUpEZtMjVc7mjZNloF6min+2REnZibHaM1r6
7RBVGeZPJfmsHjs+PGSwr22LiRCzl2gs+Y0JZl0JCbSowHcLnQMhPYNaiaO3AzDN
Kl9DkPt8FBoVgTle08jre9aKvkVfiZlmJAbZ3mGf78H7GvBw/iP3BGyk4tq+Irge
4hGC3h/RmJKyO+zY8KUvE1cf4XTjCD/QlG11q9Y0OYpxkLIKSjtNapA2qvppvHPe
YUVd1BqZBtOaNqFn25nk8k7h4M7PdY3LKo/+5NgPkVt9jXO8ljPYw7V0CxmYhs2z
gmzP8FVtwZo+jfH2oGkF78mrkRFgK1aX7dFBN7bQKwCT4NLYTg8eDj7pYksOHuJ3
/ZvHw8gw4S/1BdJ77JTMg5UFoxI+SX9PVUzGId6d4qLN+P+9tFY5n0hYIp8LGwJq
KVd8OEox9c2Ac3mfuYwgwkSeYjTADQc+r1Jca2RtAphAxWmib0lGnOhNEDGlynZ5
A81xENbG/lrvp8O1yu0QKUgvu6uQkX7XWGoZEWdJ4pokgiSQWvG/btUXCVckaFNH
+OaGvAgMAeWoL9K/ckWvfz+Z4lpGbxY8io14q+x00UHCIW7jWwfWbUIzLTsyaPaq
mTTT5VU6LRkQM/h+5w082uE1woWBb6AKN7TqrGx+On77V0QQLRfrvXNZcIwxx+3W
0TMC5IFJA07ZuT6dAbw0sJhIsV1YTG6PIDwwFXPEpuGTrTuGXK0iM9+vCc9fnzV2
luaV2mrkwS6A1PimCFZ3n3AVT5y7radFM8+p+vpzhy91l8Es57mlEOt9iXL9ZaIv
mLtaLbIQR8PH6SEryHqhpnm2lg/qr7z+i4YMG7VkYKBr1hFUTVYgM1TCOPsYI2KL
pxoA25fOhQJml2Fau4C8wPk5Reffh5OTNaD2nGdI0pyCeeDhYrNlRKloJVJDVu1i
koH+opbPKlXuW23lO25gX4wh4ApqzV0VDLyRJD2RiRo3mKGOoZ/Anbi7nuLb5CZF
6muCrpcllj43V24caeXtZB0gt5F+CE2IJi7FuJ8Y2cCLFFnA4HohHP7/AQ94vVa3
0EKJc4kMfXIRr3fKD/74a02kEeBCOMKRQvu8slVC3wbv4w+81+bRoOs3ufTgAaak
dl+4Kikx10z0MzcBCw6gaiSUJqzm4ztsF5mU0hJ3VDwn9dVjaGxGQGBv8q9l0DDE
Amth7LzX7V4QbDWZA+Ad5KPH4gWu8SwRaQMd3ut+hfbZv5u8NX0kFw1tVfIQLLhZ
i1/mMvdB8Mp5cJQ4Rd7mtsr1N2r6RTKX95FWxjyKM+4UOQDLCanG1lvDFJL59ASB
ReaJXujn0zzlxTPyBBZI5EmfzIwjvdAteEP0AfKIHgCy0wEgmKPSpCE07uHWAbdQ
iJ0YYd0pwQe5+viyNoQQrYm8oE9rq+Y3LbveEdIRlYB2bB8AeXWZ7/oU+vxPLU7K
FW0BKWa4qWwIfNrt/gpdb1KGpTxqZKwrbUNFuOMkIGebEhldtb2WC4S0FhaGVSHy
2eOp4ut2ktfqmTe8gVb12OU9Bm9jtNDEr1s/9Q3vts89h7kDVIXjcW6CGB4ussRI
VxNmwW+hWHsCbCKaN/C8onucsaGnQjcU/YYIP7KXAcEYhQ1Wut6RCsdg+JRk2wyD
w9euMQeP8o7ZhV4qxnKBAkrG/Qv6A0Wfqi/8qfY0IJL69googQJ57Ifyzxwmf6Bd
zJm9OztuVYm+JeyrTlzY8L/cGgYl1JRutaoZcnJ6a3V9UxMURjbCA163D6s2Q+Wl
/I8u5h/g6yZABEDk3E5zGaxsnvISySl74DyyzP/r/H68jkQridLFyKKtDBfXg9B5
LOLOWl0vNmg8jFlaQnYF3seEvvA3k0O6k/HhXKGMFiQMXJTtk+3U+dolnkL0QZnn
AwRFgJQZ2gUhOmkvtBd8alKR5QtlJ3fbqrg31CQuB9qIYoAhSqMbXgWoivSxsmVQ
mnBWuVakK4D7tD5zgiVG7iBHl3oFHjYu8u1U3C34yPHWnvJU19T8dmtK16G05zxO
3BNzgPcRLWEDGozMsrIfLGTp3TzURdnyGCPkzaGjBmpr4vdQiEsXcl0DNkEseh2V
0EToyGNrzzzRQFULHSkM/H90wpi+Otf6ml+12Gd7E8XWdhr2LI5z0f8dhEhcTlOo
kXcmbDg7g5QW9p4poqwAWI8ouyFFYq4Sy9uUlZHKUvaCPMbN6oTHVdnwlbnevfaG
9lWSElLK/VW+E4p2qpPOpVzhdkshBU7wYHCLVmQH5BwGAZZlZceE2g8LT+dDvKMo
kfq1A/80yc7S37MmH1B53aaHkoVheURBur/gvB6MfvCEftQtBlBfikgL4u5igQ6l
YePbypPyKV5fB6SOuTTylUzOIiHFJaNcRrzVyjemNjeRsXxKA/wmMFpjnwi3viho
a3g04fsM72QrgtOVx6MfI5UEI8mBYn5JT8ZOvK8WmnSlEFJA8WetqHJTBvmv43Yv
1Of3f0dG8px/RpPRQGrsjs41BO2gLeOEDDNqGrr9dw7qYgpF+98h1UpM5GTqQXtV
IgYs8yqiGOBgSFcTuJv2t33vbIxJ4QE324EAoI+lqYV3ftL9VtW6jm7wJY8J10T4
/4BAV+0U3ak/kFqSzueELoanC2zCQnY/dM45K2H/bchz/lz1kxjbNp5jgRzwyqS7
1ZxHnqpvVL/Yv7LLVps9YhKCj2Ocds1qoR5jBQ3l2Wsqfini1hqTLa1YfFxOszr8
K8ZkIodiVrozrTHvtIwphKWz5L3XoAT+RwRDnbVvMk9bw5UK6SdRrWKZXPE06ahH
qwnw+/BcTr6KCXhqcbaGZOnuHadQfz+UdevmYE4vmDR4J93P9SjC33uyFoMd/Ri7
1Al5dUKe+6O4zjvylEztHxcSHCMODCpZIPq8a1M4S+wVfrNXHsXMt5u021s7y+3k
Ta8ANP2zYg2fCuHizIGI5yfj4jMq0JPMG+egNhBIfQZNPnxnovgkKR9bcuyR1ZXG
C6p1fo67wqqxCvUJakymbiU0/sGzoJI5JGhvTs2GoHDGBabzHYTqECyLrNr+MOGZ
mJF2BSs5yoLr/7RUxUj9B3KIk9yUOfPib8JP7BpFOWVYjWsbmAJtZokeNXa9pDFx
x0DuOAsGIHuclCcpKR402oKRnWTewQZ2V47CKmwzxKMw78KXAicEtAv5bX4ZQR/a
YSzKxq/xwHAqCC4yqMgQuJK9BnVz+cNqVUYG2JHmTAbrL68OY648BQrGuIRhNz8/
LaRz+jqVEEuPROeEDrOVJmCwA3BRb/hyx7yiE8yynICiDP+1rAl8WqRlPHJIG8Cu
1pAfn7+KUe00lPoBGnrK0vPuiUjnabNKNzQeTiLWHTraw9MOGNASiZhaxor4Z3MJ
edDNAgqTWm3fwbSzckXTVVsqJjcJQnrzDXJrIiOMql1C5WZ+ixQ2A1aae2yi/YLe
aLNSGpMhbNcIz4SP5REJLEq+d7e7bpIFCEIAhyX83LcTbnK1rZzRJZdiviagTQbb
ux8jJ9msuTb1zGxhNjH5f7TYtapqjdKn4T4hiCmhVp9Ws0zZmw850/CaRAAtPcBm
Ly7veTRXFtwhLfxxx2lw8SAmGVUB1Pbme4JtZ+rWL4CaQqR0xbsTNVfhJp5wdqfx
ioNBNSTMzRVgpdU+u2qVoLLzb4DTUWqZjJJd5iwDj8SXNZhbPJNoOpGAMb9nearu
WSHUqwNKCWENX5n+3FZv09CQcO5Mmc2M6FA/h3lp0glSIFiOfXWSVDuTiPy9K9ap
cve++hrlefnPaOFePyHMlfD/RnozN7U8JkNNPMgGNuImlx0ufQLt+FlPg1fp+klY
B0mFtH2X2Z5NIagipE3tIkTXgNwgssVeWLwjvuUT3AGGWhAyq7Rka/1SlVldsNLS
dAvPbZyfQ0eayXYcBa4kZ17pfVVplvZY5EKG9FxEz6IcovIDlFC6DWaqtaHHPMP1
INqbUUvOVLSedWcaVS73KxeoZs//kwIkjsH0jUBy6vc8G8I0i4uX4kHJe6DQrtSi
zy+EfFLnt/0VeLaP/SY2wDlpmh+FhqgWO5me5AoTXfYvdpW9Cfh80dfh8ahIwmAk
MmuN5E2qelbLcm7kHY+shHbdhdD+7YXJLWoW5+GikDj6rV/8jeSNhBMnBdPmecB2
XymZnqsbvt20nhOzdUkhEEfymm7fJ/SEmayd/oZrIMsUv8rpXkVY0PFqwTGiOJd/
olS9LAk8SFekEUDfK6FciRJKgXD7uUBMK0UJbD9zYrV217U/x6VCAmHWb8LQBIy8
Sp5gXW9oDFkCRCw7e/xi7rldpQGwqK1DxTY6a4B55ynFmhpcmCjiJXxbaITmp0I6
cZHxMh8vgI3YiA9GIYjVBXqANg5Gf/1FRuIEfcPMdiwBnbUyYtSpNJ2Dwfff6Zu0
kBTViuKYb5K6gRSZpP+zHKiY2YXMOvfW/n+hv81NmTIzhvIC7Qv53oWehYy2Jagt
3Prcp2x5uF/FxYrBK5vuagMhdMkwE/rEkrTIb718LaQSU7umvuRGFnkUcaWWbAaK
sNBy5hIiEXzG7QYH2lnbhyrZSTFH3TmPg3XJ/PeUVL3lu7JRNb3jerENcFsVBPVf
/cy0TiVhChQkLQH49+RkCHjNBTL/nM9NU8d9ljY+koknvxAs8lOqigDcg2E+EBB+
F+vXl3eNemdkSmUDIM9aLyM8VdIfe+eCvgGFy5motzgd1ZLfvQiXimrCMo7fg/wt
EndpkF/lhpAxNM6G1w97tx+sm7XexaunshDUGcrabkHPu2B07FRcFbWA1Ba086wV
zPVJ0TQBxsaa80uai+iqgt0m4sWZ23W8O4klALu0pEbE+857Xwq/fz7CWKwHpJkd
Vf/wpxYR12TyHai3dWc7KZVI/cU/XDU93vXtv7GijXcQt1gc19iUHtypTwn5bTdC
gsBuRY0mA8NTE+VqmeSDAN8qJDze2aCpAePSmZQSDPLoYatM/EOl321yTslK/KK7
80g/qvJ0CnzihtwYjyxyYlglYt+dluc+js6MEOmEKBz/O8H7KbdAc61z9y9jihvl
e6r/ymLMLJUZxM5cvSrFxAhHmdTC3s912QwmoxNBHFQNV96FDgu863QmP6D10lE0
fSazQHswDgMKETLJ5d9/GG/CsatAotEUbOTbIN+GU7IPQ7l9fEZSlT41QId0mc1x
NJaW1biOWj2cY0g0Z4A50FIQQ7j+0diS2Gynei24smuINeWcWxhxkoosCeb1Fg3Y
4tDHFmq75/PV8SQ0rkmFjHz/GHKAWGFKtWQkRa9Q2YcuyFvISF9mRRKXuShp1lEm
pDutuStkJIlBooY3lVjrkXXQtuBcS4dVcaZSqn7bk3ZCdWl8Qj4i7wL7JMAXuQYr
bNGRDEWDNQAaG1H7rBVWv5FB3vjwCUNhaGW7O1gtEj2HfXFhx2VBFMEyajFRPlyi
NPeXAKJBGYK/sJ6391XZV/5OCaXWfj6lFjx3mANn0mCCbmJDkvct6eCRp3Le9LRu
00IkgJd1qlYF3GxrFB3i9AP3cQ44x0RET8bhCzbYGgTaIEbbO6ddNjBdHnjU2jd3
JVsULW6DjnpHt6QjajVbsUROhKJ+zgxXGUhbD16kX4w6XT15zTCfgvREAuTcGsdC
P4t7NC8KD6VSKBYdYNQ66h61mO1tRPA5P5f+JqHZ3J4qX451OLOQLEa4aYFZY410
u9rmdjjf3BwC/2Yjy0vb462Qh9IQzME6HOXREuCuMS7YCFYGfQenqz4N40I/xHju
tOLmiJHzk8Ym70ttkQ1bDsl6WcKqNQGt+XQa6tpKEnOi0zfmz4KfII9Nn6dHXvnX
SQ8XSCfRPUCCd0Hv9RJw7m5aIfR2uKIjAQG+UJUuiP88KE4tMVvfUduQZBIJeDoV
8/3118sjOM68Fk5rIM2d23iaF7FoAXCoR+REmv7tH6ypCdeNV//XjABZ4PlQLsCh
7kAWaDLs+gvwbNXmJlb6DZYfVprEEiARzWh/CuRIDvb/TdnbYxJpiPAOZ2KtrURf
fYBBbl/Ak8z0UT2D3xR/saQ6mdcjVoIzUwpAoKtPtiT8tHvkaMTCUK9BkeoxxyQt
hKTUfRCPF8xenIr3f0Qfw3/o0ti5Z+at1n5B/B7XNi3Z3YuKnDzNhlEJiHZ5HH/C
3HiKjHG56VUQAwTCghp2VUktSjzzVp4p1bv/vfDYm+CeXToibYdbh6MJtDM5eiTS
Q3+sOfBs8M/2DP6ffREATA7JPYXcUtWRX6va6tJmhJOcWdpQi3HamYO2fMwMp7uG
dzidjcrn3w8X/j1+ln0nHbdwxIRhhpEHNU9ohuiQ2jkUJPV3+wk2j4I4X1w+8gGl
mafbUB0tvuVzIBriVGp8xi18F0FOdT0w4bTH3dr6FAmC+lTlAtSnAT8vAX+4ESqZ
xGfoWjONfKOVlgD+2r/dArGGR/bW3pRrU/cQoX+XhQebfSVIat+429m9QE6H5iuN
OWBb8py+YXaOy05vDGCKLn+XV2ohPoSe2YpQYkhbFdFm7uOQMOGAP118X6o0R2cx
IWU/bGRXzDFfb5ldubejjrDOE03kS0/RM8Az5lPW666nYhbaIQCQH5bPdZ+uZQ7c
fnKHpWEFdruiQVF4bA/Vc6+saJGN+8RfRgdICa/wApdUyJcJQsdCAlh3j8AlrOm9
SJnSLcMfmIoCVuMbWbkImzHVK2AHWDxRFgwVNulVJU02mYElpfwrEAu2NZK3eNIF
vBsRIGYSpBwYj65sIkcsAjcu4W+bo+HpWKWXUqkgeuVTtv49LHI6eAzkC7IDisXj
cQpwow/FONl4WHeZy2PaOTaRPLu7dwsN0ikvZvtKynqD5MIEPMXvp79EpZf70tdj
RiX3EQUoN+5k5kWrG25vbpQhTmCk1Md64889dtwyhhKbrcmo1aoTPMcRKJEIsh5Y
Zw1djAAS7ZWO5EcpGElPqscO6FZ1ZzuuPjDSokk9FoWkCRpLn9UMC1VkbyBtER2W
SveDR2Ew4L3wxDAZuNCUaK3lAV/GVSV+XgZd6dti4RQK3IfgT+OPXgxJjUhvHSUG
31CKGGfJRI9yZROhaZQGqzqH6Hudql7lQ4j0W508YD8iltHYogy5SbNI/CtjYtve
kECRaQLVYcP//E2BdSxFr21DVDv268QdBTvfP9R4ltIKfc5wBQ+tFPkY840ZKdJw
oavVvbTDEW1W1nkerGALCMu8W25GTTyNe54KJrdCyc4pemrDFeReBDITl+1Laeot
JTcK7cacsIKZ60gsoZebpgfIHe9CwXzXT/GDpztgxaPbOYfo4mYUHQAIrY2KgxE2
MHMJVheSf/8hdVMaiEdkFWKclMMGHOuLEYnF6LI4Zt4eQYl2/Y1LaNXGe8dg3089
IfNvoUn1KZuPcmSmMyNsSl+Nd++17gu/PAd5AO9Fcsoxd9GNTUl8+pE5KO3sF2LD
34YHEsIl3Ick6KPuzXZlDO3XRWYwQaokXep5X+5W9zV+RARG/ogBkYT29anzewrw
QnOkdjh4lV7MCcTeS4Rlab2+ez0abo3QFtFarVYiE4V+V5RO+zIyypgBQwsdP3jV
bYRRneaiUgOqrVj9+un/stLZR6RvAr64uG+LpnyWSylUdJZCFeivrDCTNNvTz1OD
Y+nDnk2IYPeGrq1shcesipsO++OVDxgk7Yl+tgdxl/di1nXv1QF405Z0X1s/9ure
Z7YtW7qgvzhLO+v5S4NFPvhJUJRCAnU9l9M08zPljsv7xQOsesUgDiS8oGWTxc5D
8Re1n1CMv/2jrw4ydE5U8XMvY+1ZF+KagU6lt7Wuw4+Y9LAST9ueqLuGAVNRGV1C
3M6xLAzY/oYECIYcfi3CpK6qfAVTYXmrdvwoViUniB5AnkH7nVxb6xQoWAgLXypi
MHLWIypaPssGPC6jImE2ubD7c4cdpTEmfDN3BzSSdyCwx9QAKMH7tIXSNSYJBZxU
oJ9BmbkMuQGNJeW5nREMGugy4e8pAAabqa669JrhBWD+9u4hYAOBLQTefHNEYC96
bYVtumtA6oPF0sRQeRtJfIN82KosVmCDDaJOlQOv9NJb6wfHmG9b78lPUU6c/CK7
U0VYhKIaFyLvLSn32A/9PWaKiawhggXeKj51ETe05AhX3EoF7qARUxgKlqahK2Dk
pGJkmw+v2297VVKeO7U4QG/VJSvfJmfk5ruzLZFqvWCSmjMPuZqad1wj81j9i5LP
7JNshJ+4fvi0G0L4Lig6OJnqfImYHg9vrEztUGIROhRwJEXYTat77ULX+5eU3CvL
UFfmDfNz4cMdWwGeFRi2U31xAw5jMntFCj5+oMvpyEBDavTJxYhlMqyplhIHSzGe
/lfhQt/CSxu4QfDnNsxEx1+48u6iZ5Lm6w1oHmYhlGei8Qw6lmP5rz8EoEFBeTpX
lilMDfkj9FAV9zZDjVGf9nDKNjr25HNAAeViRfE12jhX2LQ8BSpzK3Yo6WT9/8pM
BveV9UvTQSTP0+sXyL+FqH/vp4QyEVet8f3DLpZVMzB5rpiPPxg++qpsl9ioLNky
GJLDo+ZdXOZsQ/fZmuTSx8A96QzhuOLwwjK+dvc9m0fy1DRV4LXokw6Wxv58ZYMz
Jzwa0CkjnpOI7Nf1V7g8gukJeMaBXkiI+9ZR1A7CVhvk0ymlWpOH5VgVQ6aSLGuO
34m73ynPDsjzio9kYMy3dyF5SDT1gjDkIYKNzTgDdRxn9bHZiatupqylqQHqlP7h
PiGbO6UPYEtqzW1vz/2Zf2J5CNd2UsPVJbQIAyy9AS3ngtH5amNvsaKWhC9Ae+k2
o8DXoNb787wWmDsJzvZDMCSlKV1DFVnQH9GQj3GKeWXh5FuJpsUkGR/oU9lXAA31
heRggcS0jXII+B+v7CaOnwvCMr3ZOKAPZOdc+hw9UWquVBedyAPmkhu7HFx6nUaN
xLOrnCd75TYipYhYYcCz5Fbyp6sOjFIGfQMvak1qgTcTQGck2aXjpxHzVzY3FhNN
vyVV1Req/U0Z7L3KpBdY8XOhIp7jYNaifVd/N+21K9s/ddLMUYj5dXYgJ0WO5U04
2Vn+J0LJDzPpklPPKruyxbi2fciLT7EY4KMpblwd+0P01bquTwVowwoc1+CKWZwQ
vKeOnHY7zlmtxZF/IYSgycsYvVDiIymax6/1SkncGaJakiHQMpzXeNTHr0XjfCvJ
ZJGgFcIkldEhOwKxpwV9sfCgPcrD+J+59zIm6JIjx7pA/J8TxcpJLI7f+UU8R+Fm
EbjvgRIea4VtVdj30/HxyUr34z1rGMOT1Iq4WoB3PjC9pfiSeqsnalfq6C49Ol/V
ke6XPM8nbff04Bg8esvb6fDjaBT2hie5zz7bV70SHXwKhGLoQvq2WRojyOeDay8k
4pwvuR6h4sac/7Pe9lt+vy1n1ffH2DEyK3IEgXYtksiYIKO0uyr4FjoAqrc1NSiW
4OlUZiWH+X1ythy3FYghLO2MMWQyafxVtTGAu1YvTRe6QvR6d+16i9mrwv5l9qnk
eA1+OKtwMxidLfDHsuPOokjlvMHyL7/7D7GoSLb1CLPQWeaCYejoF6khX55PW56p
zVqRPJvAR3bfXLbxYWfRDZvGZzR/gMF90Jpcd9zWfD4yomcqcwfZoCBtI0FCr8di
Cypf/gfUaBA8qb/0toWtGJVnYaGiVU4G1DNfVNQUEHq+BWRCr0/LF3iYOMcYrdka
6KmXPQJRcq4i1ZKpop7f6M4vs/+fR3ouOVCLd7WJLMfYQLz1udWGvhRVeEhSsskS
c4S34awHuLcZvuohbIGsEM21JnFIytR2cjZUxpbYGdsdEZoUOx0Gm5/O3fa+NhvY
w5MbAsbEUjMorOVe2PhO3atpGvetWMwH/+jNYXlZ3RlNd1j17mwREPMvtX+KVVv8
D16GSx420MucVQvHNZ3I9goPQgIWUmrRAYM5gAMDgwqLrzXxoWGZYHSRBnsboFwJ
s1NQDWpwY26HIArMH9kaDCsbbbp9XOfQVSJ+NPC2DP859Xiter4IXx1l/jMFHTeV
hCUXYaIZAv1R3LfE10BwUg4Dfbwli7J+1Nni+JwxeWf/iXqEYaIlFix8SuF1rsAC
2Nz83cAZkqrSWrkGfh4KFt6PYA5DEzz+LaQoGK7HeFg1WHGEvUvXVpGtYVZmp3QG
J/WfMXtmcQiKM04rIPzVOuT+GYYHZHrNZHyJjKTwgCXwmLfDy8OUTxgHZRe6Swgm
fZv2quLIhEhAkahA2hwR62OE1vBpH8lWDdCrYN02Ma2D7r1sMdYDORWUiHwm9r0Z
4h+R7s7vTA3bvegzxajTB5yO2rCKrBZY7aTVE5NGFTrVgYnL8CrFRQuDaLUbWIN+
A+w+nSv9JL8fdu2yyV61RKXWM/DjONgWLmNdGnccqctQJvG7+Br3IzeDhU5Yio9Z
nFpDEAvrSxy6zc4q0eYo/azzQ9OmGiq3jWd1pAFNuXAeQgylO33aws/qpItVMczO
BVQdBTflzJuxoFys9j1XlSqbim0raeG5djYGEqtHvVbjfsJzjkExQ/TiaJy0LYZQ
oDNqaeYh/gcmkxKy797K9eMq9k815KZexFzYKyaVS3++G1VIPwOZGUjlOXUdsfWC
5Gct49T6mXcfxEYnbqbsyVUoCkGe6mnrOiiUhpe38pdMyc5Dv9ChvRlOgu8iVBzC
pvmK1wcxW645hvMqCzqQwVFGWo7Rc6dh1L/dcQ+kD+34A8AdMifKhNsxnHBiQ7RK
ACaIXuPTowrCgKeyaveSomsO4vN3QvybS+gGDM01QzeCjgFJKFAr6cQlIQ7xzgc8
PEhXsc/UBr4l4lq50NTCYrsx1Yklj0D0KlW5J37HXv2C9EcZjmEfy+twwMvuKk61
885Nl8+8A+KK3XN2FcNnyMWUmHMqDxhEs+rx6Ie7dSSvYpq+W7vdw3mUXX9ReXBw
x2JkWl7XZx3bchkMJNlcvDzHfhdgYMDIPSy1I1Dw/atCItcSxIQO+0lmhWO+hS5t
dmHNuMbsR60jRazYBMHzK41V5RH8brWa0tQ4jF1W4SF4PpSUzXfe5SxDJv02+bmV
TDH/Z4JCiGmSsVbhPfXukQJD5qeaPxbz5AEDJKBQShXBb5a/WYcVcMGlp5JPICGj
QMsV2O2PVY3PaPHXt3NURkqhBhqejOmiv8ng4FgTtWOQqB+8vKNkFu2mp1TulF5O
i++yOoHpzBn+TwApEgKBexJK2O/VUIDRGFrtTW2bOOpW5NaDbYKw0f2gpTWwVcY0
fOGcYtZ2Xkt4DLlVLfM3pj8Xvn2F22Ns06tO32TG9G1Jl27iQMCXcieaxQl77A//
nfErBsGyoXIim/MIAikK8DN3K+a5vEB/A4JIL/7FrReHDvh2yVJvLnXRTGx7CZIr
PJj1h+oOtSak2A02w9QtErdhNtUzd+nYCWr8nrK431vtp0AjZynK73cNpn3RELca
C+Bjcj+jOPm0fnmV9ZbjyNyeEK06SvOQgA1eltOe6bLIpJeIhFA32Ul0cwuewgzG
KduhLc35iudgI2+qcVmIGGRoasCFGjIQcpMow2j5jfiT3SGid/xix+zHUOItkPO3
l7xHUphWLugH7D6VRQRohi6vwMTgu9vbNxf1DinmvdIua9fA++WohJ9W2BWlOGnk
85hjHOTYA2kxzf2N0d7dSQXDmVR9Kystk0pa6OBDVY5DFcyRztX/+rSM2BfRr48P
U1aF9NlNzQyjbdW2H5TJItjfndeGubboWgxOqc0yANdclIaaJapquc+iiT2kVgMZ
ZRxpxGEz7YZLK717pMx+wTHqf2aQTVumy56ooO/Fy2Ex7rK1b9+MbhTpT9eOmcEr
jh8uJVaq2ws5BYzZj2g6Q4t9SkMmUAFF5MtxWuIswkw9eVnSZeegtFUdXJ4ljsCT
a0EC0Bak/q78ql0Tq8lGTCItmmgZ7iyGWWfLz/FaXc0+z59xHuNLXCBbXWHJX8We
hZyyzbrWuFwUSEYP84szJxZGrJyzX14btHDuTiFX4raQrKqRq2f0FSQbhE1+O5Zu
y6AxgDm85Ss6Igci0SRx2R3xiamMaaqeYWn7hET4KvKQDPNod9KsKpRYdTBt7LFk
m24QCgjHFQ4Yj23QHT2gYB6+sRFhAbSAbwt8h5yNn0HGRgsLvuG584slUOHzmfKe
f7wF6CJX+EmgcF6qky2KC+0ZSGUIuDS6N1awC4rDSFktYsLcZ00STATMRIX9L5Dj
4M7rM8d43uyk5sSNIZ1NBl4rCnkxS0MrWdaWzI95wj7wJJXkrM7lZZlqw+V7JFjx
yy55EMF0JQ6GRVczhjvT53h6uyJss3WpFH7ViOgBYCinVWnkCbY3y7IbQtL0YoF5
x/D81yMsY9G5J66z6Rh1sK3cQsPNmLpNeOMDi3uwvKXuysQvDGSLzmJv3ygfBmQR
uv6vfncKe21HLewOAMUpjMvqqXM5Ww3bAb+0usIdTnamzd1e95P7ObDecpKG9mO3
BKofVw7sbMjsnvk7A2bk7NkoXCLE1OleNXWzQ2akeTN4Ixw/6mFdUY15obH+YL8b
TrxBIo5k0oA8D0DfSaxkjk8S1GflwlzWTgCNj/60etoCCqSQaVBlkumpK2hMCsxN
KAZUr4XA1EpBc5KBdI0ykCwTjHppQ4X0yrWJR+ZXl+4j8JrFtLIZx2CHjK9IjqLA
PRR/2Hxx/UG43DlcM1FMq2EnUoMHZdaUR9WOnR2vfiHeATKm3zGI/Aw7iWDqMbdT
X85S6LdEVW7Bd1PYZmyqtpDizyXgkXE5022M6Iu+q/kjKptXlBrQExZpofKnF2FZ
BjkETxvM6iP5VylGH13/4qwD7LUrKvzinmOVqVCaJB9YtpC3irl3nSHBhdOZLDSP
32Vsd3bhwHRvJgi+A+mWXbZgBFQFh+lZAMGQV3hIG/swJhMLP5L0iM9KgWhNubLq
hWGZAGgKT8w1Tm+QnXgDT6dCNXzdEMjP1SL69WuAcePV/LqdBE/Rgs0n5//loLXC
VBpTZefHruWbtj0OlUUrj1J7AJ7IsBKdDds8UP09vZc=
`protect END_PROTECTED
