`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2I7gyC50XTCsTOnfHRd7y8tz4ZX6p0ou6mycuVYxJ9gLPvwCcBLWtkGb9NmHH4zN
uWGB/UMsfU6SqrHLmRePKvbmW01rxuXyhtvi4RORDw7YhCm2Pfb8gn+qy2Vztpdw
Ontej0qJyCGUmcyCfnzvtdBXD3AzVsb6uRC6JpKZWaHNiUI752VZehi+BMGwFd9h
exyZJllJSh+KFuFE6D06Q7+honEFQcnXgiAZ4WkgOXM8IQYexpcjGhpUi+1RR0bm
lTXpw4xGzEf1vWNL+jPAkz1s982T1uDUPeEu8Sp21xEppWApDyayT2WHdJ+wUYkY
SIsQ5KBn/uFq+0eaEXWPj/Qyb7Cx7DURtUDAF9aVU5Z3W2Z49u3YZbcrWjoBR/Mg
FxZY/+JO8rkQe2dbxSVN92fXasw2ctYp5yHEG11nJsr8m8VKHCffoTNU2RtJyc3N
wiOG2Rgti1PvLhjkwGF5W7y1S9NDn9xvznkNEnXl15Qmzb4l2yPTGimT0npfxi/Z
LH212P6DluMWlhh5tYLRfhTeEt2TD695mGxD6xXCIOamjBN8mmlu2UqT4TDTSwiQ
qrdUpszbJlVUUkNBGFnuwZyWtE6zaMM0uL/ZvEsQNvdBAIN6Q/R9Ab15ty0qsepq
EIbm+X46HUYIvHqFuI4D6zPeJfsY4L+oXDAa70mv0UB5LE2LU+qUezMrNixJYypw
OOv6Nnd1K9qMuMt7jsdFJUOpwGG9vVJfSeuj9NknqaKiuXP96fJcPUH5AC6H40uC
AG15ZZAr3lQ23w3//345MxzFsTfko6zI5En21nYc0yocpAp8DIyG1qf/Q3LplEfY
IZ9cu+Yicze6k768PfeURBDkkqWZrBbV1rVevYUHKslJ1XiEElFHJ6aUlDhl0oSi
356if7313jh7Uw8xD7ex3lGeU/4xq6yi9O4ErEApkUk6hdehFSo4tIo9lMiTJClG
AgZLjcLcwJmtng0kN1PP/oW+ZMlvAMMAmJP+Nqu8VHiacDIEft4x3wzAEVu6Kz8X
SHC78jDvAykIqcfquSVZvFM48F2yRv7PPib4HSM4gOlF1iegaFTkxy+P226+6gZ4
bFihC0fAb2FCH+95gHT0C1xZYKfH+3PRNxP2aRzn//r9jOp3Xf4nHd1v4TElTVSD
Y1m1yVnWE3mE0tm/2eMrEJqI6rCoX7YDDT1x3JyvJ/TCHcWSEsZ8VfuiP7ZcpicG
CGgN1qHl+69XksIo3lo+YBrBfNWPsY9eCEGSRp79b0UxHOYUQPUZDrm04PxYHk/P
L2XxHkvWcUAUONyCzKuIO4xkkq5FS3fOt9bKSQG7d7JGhA8yiHxhvVHU4bnMG0pW
1GT61xWxA8phMkgvdABgEXDAkk+K659YAEMAqOJihyvjLSxgUYYjzpb9wW8O0bz9
mXOriJBeBHh85YwTp4MDxOz4d7DgOUPBeDX67HsI0bgbxZvGynqihPJXbp7fxpSs
CGlCIL4j8kgFhA37CxVC4PYPsYAILj9a8UmQIV5YlFUkkDv8ZTQk/JQDrEtHdKLN
OVYbVGqwxfSd8TRq7up0T/dq8F13rGz8DalzJodWkhl8E5unMzHfmlcwffePc+8G
Rnbpb67HR2qBhQr0RqciLEfXaZjNZMIhAz3rnUBde95tfl7xqdtbk8fuFLP1dujP
fdYZdZt3sE1od3AQIghDMJhB9bdv4+5gbM+a9VQZFBAD+6Xgudkgt4CYCVXRlvVv
UTgnsaPW9UpSaX5wXvd/SH0CZuy8gmFQ2BpM+pVV/e95aITOT4J8nV90mBVLCiSi
3t6cugcLiByjZhiAlg1H9RYkh3BIBDxy+rtZfhaXmfl5zKA/0QDNgwJb5zMmpQPo
UUOIoP3Rct2tBjnJLTTBb09xiDbVVNyM3kQrIxNxuXl8h1anBgTHnZfZS/ZBk36T
7NbhXXOwe8aYzEsRi9H29wdJORyKBgiRnWbNOirJ7bExCeCOBXIhrKwT2qqnvwmf
rOPJV+lEtYTtN/M1J6sQv/chAsMJ+b1bkL2bWs4P30SzKkwr3GOc1Ka5z9qE3YQP
whk+NQeZp4wQi6/j1tyxkhz71udQKwT8IDcV4cox1HYedUfgKjHMO8V36dBvrRMB
6Hnb5GCIRjYgot5kRcMB+5o4Q67I0TIIO0oVy0IL1UZt8Mb8CDv0J4K5bEhT+8ep
wKjt5c4NL2zGKwCb+XWpyCsw6FHYaBms3dLOSFTuYHETBrFDYjYaMJ8+VwFMJB1t
eh/vAleCnfzy+dsYOFbhap84GvjGFCgBFHNHmiax6+qY1sUt1St6USY43hnJ//ZW
F5q5xGNtZJxI3tC9CSG5wmD0PWut46AZacb0nfGaPYmPQIBkm3oteeJDTxM/oXMM
CbUh8XX61tOaC6KdmT9vRzYEkQOJ1LUweXHrPM5N0Ge927HyD9FFr5K6ipQR7UXO
ylFujDTvP2AvtPxbcsJl/ABfHoGuWkhPLXMGe++5I8WefGZUwKoVk4Qdau2gZGLl
Z5E1CvgM7/ZaBJ7UUjMaoGx97+m1oxqzzSFweeYuaAJdjTSb228P215J1IZKb1eO
lcKzVu4h+ZXMlL1LitauOPQbh1vu1VrpA4IIVLHZWcA3/c40zhqBNJCajyRYRXtw
gsaP+56qfkP3WN/v5kl8qb4G9+oMSfqT8xHnhUDmMU7+m0BTfvm5j//Ml9oq7g/4
tfHPUVyLrwud5E9k/z9vxFEBJt0Mb4D1hyVWK1WQKJF1L86gCRSp6lY1V68QwsMx
ocQUM+fIHE6MZM+v6BJaK4v5XdmtY7Bfx0MPwBy6morNfMjZk1XWSuuEpxLgeHiM
Rd6YWf5SNnK6AU9UN8qJwwsZ2QNx6uKZwNoAO6bXXsbeoI1iJ/S2m2E0u52Drtis
T7p/V72edP7M/P/Ipu30U0/eIWBVeIQngHMqpQj0NWs4YrbeGYJ6iOIYTVOJe+PX
hRVVeefldIVos+c1hjw2QN0X3k9OHb64ltRlCZQU82tOfACGnvI9Tl4HkBObC1cW
PrGc/VBsbP1Sj3VasLnxOCYKvzwvyUWErDv69f1xP7JdmScmrq/v3ufWUg4Gxj21
7eB+rnURKqIldQyONovwpQzDfRYE9jLqeN4rXI0z9ryJHax3d1x70pV+8jq93Ek6
rSAic8O7RqXVatMoBo0vaesbsl+7BaGBvP4A+z6zW2w8JtSdH3xJ5W8Dmg8b8v4+
w4zblYdvlCxogSM7T3bb+bWieT3H2NnsvjUO8i7UGlGX9hYDk3ZTpo0kUs217yIN
5gDQhyEcMv0gsdbnkGurmkYR4VIHmzyumoNLFTB44BI6uQBiQGi8sFVZWqqESOl3
XffdgVuN2ko8hwYg5mbXvomJju6Z5WbkUVmPD2Hp2JhATb0L6vIp7OJk43qHEWv2
ORlKxFWTbe85fmdveMxYY2uViTb/TcncsgPSD0tIgs/8KTZxwkY2I0GcXGfOTP1L
Q4JUiFwRLJUfOdyOHaSMO5xXreFaHBfUCVpIh2pOPTUlHjmOH1CrM4lm5nhUDGgU
xJQlfo4xSoRG7B9T9n7H6SlZtu7J/R8VIXDgIETEiIEA/0vccz6qL8DSCTsvD2Tm
R0PzH9FcZOQHwVm4Pf+IdfCKNwta65eD2IZBe7SS4LvyfdSM/N+QZ/xkCdpxVZ7A
18dgp8kN1K4KgpWYWV/uaNktoMLCRTaZFzOfisbbh0WhkHRpTbN3ll54oMrUCMWy
BZXBXde6nQOwW0HYmdmAsfLHx5J3oy1RtwCZ/hUEVrlx0MkhS+wXLViWH3xG1qA6
AytQXMoqawva9zb28gKimSIZDLUuQ6mRnf0d74ozhs0gd6fVl5yXVgAPlyZ6E4mH
3j4qYAJrwF/eKsokwUG6ndM665/icDTdlnEslUZnpsbMjExZTVt+jZO4j+mqfGVB
cUY9DwiGq4wJ3gaLULU4uKAFrdEzzdowQ17+uA3D++U0ATPZVMX6/V7ZuOmh9Pvc
ZNpDin9y+Iffwmi+tztVaAdPpl6WFMeng0q8RhwIEML63UEKbKnUJ4qIgzLZcjK8
luvunTynSiCcdEt5S3NggTAa95pSjNJOOPZjgLEAzrHNG124rWQ2PQGSLj3Taz/8
vlFSAOgsNs7Kt+icvkpgrTLp20Ln2DTF0Fzr+I+W3qPtB256KEZv8b8dwT828VON
lR9UcH9Qv9m3qEz3cqghEaYwSnzi2myfzrjDcIzz0suhna2afcx1et/2E29RCtQb
7fxZaRKfwUG2d1ImxVgFvTVQ9kHeMAUxr9RaAF93mHKPm+Ex3n81a+1y8tSkLRsT
Jtt2LSnSMH03JdFy2CqR44fs3Z/51jtuQp05TAfDBhsoDh0WM5/REyWIexUN8UE0
o7NI4potIm3tIErFP3opgttENCujYjc6YyE1lkaONGfhwWLC7vkfHLZuKwhw6WhR
WSBgpnw/lt7p3PoggkpleZD3UZoPGwJ/2TTXTr0rHhlXhiwpxzdDgQ+PKJgZ5OxG
oHPoyibV23PAPv4c1YvmOzkrbclIxIWmsLcm9KRsBqswcb5iAxJTDm5nBPfkMzzQ
0GisKrP3ncN7eNFqpM/sWRhSCXQHchAHSNbMepdwjtbjGR0n3rkFh9ol7EHqAf1i
MEaSsGHL552wP2qgtPQSPYSRwmx7YYyDf2SMcFFCKw81i12MVbh9izuyTgA97Z0G
phztP7UAnyqh2CAFBD6SBXOBbmJWdMmYuSsyCNmEZuVxnN0DiZ829iadHvgCbmW/
YGoAYl14DhD5H/GDvJk50X65o37PKNfsBm0HNsnXqxLuIGkH55zBFT+iuONuLEgr
QG/zDwU7dzuxS/DEubGZy0EVn7Jj2rH+EcwVO9jlTKKmfSpjaR8Pqj+vloB7Q43f
6D89BgDkW2Ka3U3n9GhXDZubna/BHkeYFFNQ6n8CN1NPu5aEzfZZaIUI9JVZ0KPb
T8akBaTfe6hY2RX2e32Jo9mdGoJHio4z3BIe0ZX8clJj3wOe/Nzs1HnkUqVH3qew
nUa8nnhNdMVyTH5arAjZ1/J4xEobE7QquJEXXN4SQ6xb3nGYrB9XRWUbDgizx6qK
hVBsrsIcmiwbcCFfdTw4phH2NbJTOzkb2q5MjPAiAq/BzKfovbbJ4EYVeXoLF43N
NNZYIZ3CEoSxf0XZTCfAmINooL1zR0KSp0kYgW6sLhHmXzyxYJkjZcexJ2/NNqKC
H8vELyrNn7VC0Psp2x8NpGdhJ32YxW0cYTiDLcVY9taIHFBF1TB5MGGYlsreoDHk
0ujkZFGYLS3RIIrIzlkITcW0DkG/moARn/962BoGGlFy4TYPT6atCo+GLW24T+9C
R2cQ7UBvp3esO7oPsPoxqXk2ySEs6DroEy5ihsRqNm4UgJhcwQmtpokL7YdGvC4y
bdLt8iGaMyZC0Vw2RFHZMZnzP5jMWjDCjJnc0Qw9FicBT5/lVglulB9APqbNogzO
IX4GgbYYZ3+To8oottEhiR1UL3yLo1b1eU2NUcc6aEnOefIIIee+yBsmznautU1S
kTUzQV2I6JbnmLgted7DEn5dgsMESMmtWGnDT5on3htgLsqsbERud2UAiwiX5Gp9
HWTb5MZm9GlId6JKZ3i9L9gWZr1sPIPilR7lxaEtehPspuxLFn4NqtQK6zQdG8n/
XrjbXw73JmrTZEiZ+RKQsdOwp/eD2ukM5kFiAMx0a1Qwwh1EJ5/Ca7npaSaoF3dt
/W0A7n8sN30loZO5Lr+XR5nWE4qp0uviJvgfGQmoVWV9zkP83ye89PNXNDJAekPt
qtEP329dfDNjeFERElNHtszDUqdIDtxW1o2yw7QDG0cIkbytydL5xmt3bCUzD46y
GwtCX1wWSIurCYo626DzTWGWE5nbxqxAIRLOkfdf/Zp+k3qgMUYJI5KkzfXqfp+W
/8GUSRoNsrD5tSvwd01QbsKcjYLLjoXoFBaDn+pja3p9+YrP5LbqELHAW9EYSQ+5
DqpVrrCluSl0SWqIUhnHiGJVSaGVKVgWACJoXocY4PTycWVAi8zUlEyXqbINdCyg
nH0GXiEvZwwYhitobUSf1xvJlOEXgpqEIAil4/p28o/xjCziSF55EzRtHSKhWSfP
zF+49vFu5n8D9rIUg/CtFvSUS8e9htlQjbCAldrd7BpUSbr1G2Vgnk0xZDH/yLaE
RgbrozsIhpr5Hn596X3s3FGMZp4YdrumeeTInR/Hj6ei0m9jDBpaN4ecodjDP2DP
PUpT3iYJJ3hpTbwTXEn8ahlYej0s+uIi/JyBdlm6eNN/CI7JqKKq1YiV3JC22XS8
ACJm1WppQ0tU8JxZgw+rimxFbUF2N87m2qzvjh/lEfURiQ1GXQCc22C050vg4+rr
yz5iNjTFfB03BUvnNXIhObobQhPaxtqkL8naWtdT+IH+O+/DeRtl2GQ7ynVBY3s1
SXmvLEGSuSIqomNHVVcPvD8G78/Yab3USOlksnhGUli/oPQkxPyAWNic87H28JYf
U3YpzF1HsmeZhg0ArQ8ALhC9d9OYbY+rz6KVXSxqpB1R/5vGrekhrddhBZ6QnHE8
JROiES08tF5dEj0PgFDpenLeTvhB3SY68K8cdFdW3qowYYP9CzIa+TFpWqI90Glg
ud1Z5Kb3Ii63j9w/JyCNXZGwt/rPMHwcFUq5nVtOkkALmskN7IEtaOiBfs4q1Clr
1fXgpi4dWF3w39LjfOId/GRQJmrsCDz7K72dHoD4b75P+D1vNPArFaTkwgFCh05W
q+AsKHFRaBoHIMpM55258PPsalKAqZlUuIksARHHeCvjzmexUBYW5McQ9jl9qB7t
wRTdGsmFnIZL6QXEaV/Tw4KQCr3cKaI5afqrUeEGGxis7JdBDMxqaqj+jqaaUGR3
+rxHDT9Nx3mVCXYWUC6T0hOoFg5pTU9Qxo+jus2Il2Xp8dKEBAyaHMYFYqr1JGG2
Bh8apB7Mw/xZ7cXEj2jcUnPS1GDQB/pW+upt+BibDnbuFqAlzQOQWKXhS0SPYlp7
Uht4pbKgO+cHt65UvQgnfAelITEN/PO4f17hcNnFJZA2PfpuZv49cZ5ZEPpJ3qn4
q6oNvhoOojreicaUjtzgpXA7WaPakUKs1tiy7zTFu1EHCa/+gO/5Xtg//BvwxcM9
IkKu+rTn3E+S61re9kldhCuCoePHkvIOZpJncdI81Qu0yAOy7bo6I7tyvkPQVljt
W9VsJ6ODmL4gt0A3pTi7jDlLtNA11pFizb7XYMxQ6bOjnEJoZAIogZkzpkojEarz
xae9m1G+YR9AonKrirCcGw8ABnV4nfrFlnrkpaqbMtLsTYwXXwT9rmmSm7UVbGxN
grWSPyykFKX9gfvruUCshZSP2+QB1Xq3iZJgKcYbdJrJyIUY569KopNlR1yh7yCu
NX4KOOMxG5PexO+F2rsLBKJja061qCENgYHpJVWOarBpS5oUowcCp1wuXDqDj9Ik
MfujLqdhVoWA2O4oS5obYOxt3f6OjM8R1FFG3wKZUlK8XsliRkVdZv5sGUGE9cn7
V+sEtkKIO6PxiVF9pdMgZ54xrGR99KqwjdJTAnRHwThldKRqubX7qfzoEVywqx9H
xb6/wo6LIP4lwJkLV+/QO5Xb4LlWpJyvnJWURucFAIVcRgOAD8D28lK4KZ570IwP
Cg3d0scsARexKydNRsnIriZwUsWPrO/HUiYl0TSfY+kGRsYnjDz5vIKeL3ZPpX6F
HPmew8uAWCK3jt1JsngPCj1bXCmWeMYDN33RJ1nfljdxAtWs8G2sN+ZNY20sLIKl
J/SPKcvu/snDOYq2EF+1cNEfLXfzueQl/ysoYjxRldKyUNbx1FxDHujV7u8TS4XF
sJjsd+dGZ2eD/lRQ5ADDGZ/ww8IsKFRXR17K8IkyUmVh0Do3Lcr32DbpPqWjqHCj
ZsZte5UGuAJyKU3Y/2Qq9ztiHMxbeYpshxiqMVWC6/xY9/HYi48+0xJUDY0PZLWz
2RA/M8az+uzc1UbprufYw9dyd9TmpmdrjeXRzJZik+QauVkySm4lTfyh1btd/cRj
54CMeuv9voYaiMRvpjZZMLD3QBnVchf0Cf4dQ6YecavuwpRHzTmIklJ9KAnPL7dB
Jv2m6lQBZrkIgYVQeGorVvql8AMNTsLdLAtj4fZki37fyPFl+ve8xSqcurqS1WGr
CQLxlrnWy1rFqGTfQH+/0CBA6G5BwZraCtcdUqp0fIDYbSO8zlghZ03YzULBARtM
znHBKk4ifKXVdX5ttf6lx2RXVgpUhZ3xZaFmIjcNj3pdFUqr5ekB3p1Ot5Y2w8Hi
gVtnn+Ncho8lDFN74RxyPS4h8rTXdnfKqSGGnUJFx0c2N14tNS3C9+X+LRVAAPjO
0nx8zyLGM1TK5M6Rb4O5Z4oAX3DVhurNm7APPdpLFCFhfyOGfBM07s7oMg7U3l7V
gmYeYEDcNNti9X6uUf+AHbCw17mCWPaB/sBzde2ioKVJSVzqibg0TT0jEXxluLSJ
/RNOsvQVjR0rC+EyAcSkVMzt/EL6ZL2YGSiiLpX+p8y1mLATv17+9AB7jWcBZX0F
sODUpzwXzsGLJTwCIMGaK8BBKcxBcEYDXP+JdiL3L+c2aqkWnvU9nWDqlwtxWPad
+CAvhRgA5rdCuuit7+bSJUGM2C6Dc868KWgQYeLpUWJPEkoAT/SzjsE/FptcifZb
3kb0bVh2KiFmOy5jfe+omgx9SjjLOgTfqowm+n1qspP99xHWDmoA75sigTeG9RdK
XpB/a7WdVs9JzG0rwlysNG1ISBbyFL+zxnI7bem+0J1qLysHdgX72buX0HYtnZ9n
zMaLpOuHOwgALRUSxZgvcvdF9fblSjjD3qAlGtx+8aHxH/ifVXvC0x53W70I4G1K
u+ZmeB6A9XhnS89j6694W/qRBszp/kFpZE3tZapGj1AzG9fx0s0mrVORTjNQoncH
8g6TmSzc4sFWuCAEpvK1ZV8u0J2YIZxXEH+eOqmHIzACVmJFCymM+y6jtLjD7HPo
ZQv3x/l17LHuhsbgPGSqrg24Av9LvEWAfXDAGE6TbT8pBFiwn2VU0f4dvXY48pGI
Q7Umv5FuxotDC3lQsgolz9ol6rn4YlPnb/70X/ljVix7jibAjWit8MoMl4c6DQmw
Iw8LL6/dcSxvQcriYaFk/blTDcGtmBipyEHTrbilgcQEt8Y7eCmesa5LJpFBdJ5B
6EnHZdiZKV82Mq0UGI/08TVgL5TnGTITMkU9VgRbp6RIWJLcUdHfh71RhZ9/MAgV
ClWJ98Xrxhy4SV1No8+Qho4B0fynYmadgptRD0Ec5j/vvN8TLe9enEWlTXCI8g/B
Oacm2dH41F5Op32RPr3zTdX69Rg7oU3wmlBllPJ6LUUPC6zhqyT9PJypKbSHjESY
FigGFjQFElV2ClUIFwM2Tl2PytLtvuBl3CkGR4lacqjbH8N59CLBLO7HyNueJRdS
AfWbODV4IqFwYVBEwKfL31stlWuViTEuEM3RxM5qKy/QOAY2tG7CALo3AYRQuunz
48KgQE8C9rOvmB7W/l15ioBvC2ua+CiEmA+yi0CFBMjonU9xwif8EUkAvrfyv1vt
fdCdMzdiPtOd0P9+kFFur5YNwE5auTFOPxGmgIVBwYEtb2O1SMWg0ws1psKX/UeI
BRur7OEw6gbSQm+HkeaS2Uz6bjcGXXe1sxpUONqgp7jEdkoxlXNQJrIX5bPDy6bq
4cAaDw2p5iQBbLIL9yRNfSON09DOlFulTvnwM8Mq1pRHbR4Xq08SY9WRp2IA/ynH
+R3Xu+UiYvTKrdbYVKebQelRSuMiPL5xMf57fjcz3AefLOFgbTV7z2Hw7uRUAdC+
FGbKbyl72vwXTZ9BZrvL/Exb1wyLK6EXfWO0ehiWaRK5g1dZn81FOMAKnAmoVca4
INY4ccbpYFvnaRQ1A3rX3leRgZ80Lxp7tm6nuzJBmZfVMAIFIlnmoci+u3L3l590
/vsmUs3jhGF47xFxC9hPZmTz1005e4mbNEfo/Pe0bFZ8UUjYFnN5D3sTE7Jh+TM2
lrQzhNa3fQjDw5awk1XHpbjhiGS3IDZUY9rcYL9ihpTLke8qflgUtEe5WX59lH8l
uxnwV2VYV+AYCPfp3tJsb1P/QCWTrvE2os0M80PrDWx4K62KyJ1KyP3Sqi/l1rqp
fKZuvMCybgvtWPexYePHks8z0J5a2VlTzoV6PO4WomX0TdihenG8anP6x4RYCqJn
K2tr96Op6Yavyxk8i/RYQcrenkayZPSH2zVgOPCZrvS2UIWP9jSbQWHtzVcZE44C
zV1CsJFyCJ3SpyUnU0OY5gmHQAwWmwn0Y3DFAXTZVWRUGe/o3+h2T/bl/qK9NwUV
gWq8Ujxh1OT8igoUZUnhjvTMLlMK1Yl0eBKhWwltIXyOrCv032nPMxyJ5lXE4qOB
HSPll1gyPW+LUJovhaY/0w7ri9iy4WbTlwAgZfa5YWVb7ARGjZhecQyPD66XbZm9
5LlETNKHpCZL5WN221jLQ/5QMjnC5p75mg1juo9ccTU7D3Nnn9ymjSS3rESYeduL
ZdiuIhMON/2P+Q11DIses3LpkGk5FwIrJHJlpPA0S0CtyCWpew/eIAIsc+ZzMOqS
1Qh4JX3t2xwT2liyRSsI3ZReFzm/4aod/ooKfX0QJSqEEPqBVG4I19/dPxo8UXu7
J7+4+K7GIwMnUcyuzrtqjXLiMmV9lI/2E9h1Yd2XgT1owHy4MQ/PPwXBaRvYJyAo
bzyHAws5s1DeUOp1XiaCqiPzok809ExrOz9EwXCypPsYBgZ+nVWTch8x7qw3S/37
iJf85VjUUe7cx3rgilwS4biegfBphZP5wsfOPByBgOBFNPw0Ik73v9fJStK+BnH3
A1DE357qbimoMUOv/uBvIynmfKuDt/Z+DIY5ULFA6N+xPvGHhe+08QVmufw9pUbY
FaFdrmyw2X+ykipJ0CKEMHi6SJqGKFSPPFy/aqOZOKMa2fD+ocwmxNWzSpj5D535
ENEFJeJOnvSgFGi+XdWtbScadlMHKF5K6j4DpOj+PM1mMJ/Dyf4dnnaHOMOHv7NC
3oiV/M5h2/qezRQaGMuB+lsQZ0evaGPCvZX1tPEA8DO0fyFIygHDdIUCz0vgGq3K
X4BX9KqvEhuqfGmPQ6getBFB3kdQywEpUvTCEM8fU/h4xJvM71qi0BIOLEzu/TG5
wY5WMwZzTO466mRPuw3m0EqqDkw7DMHJ3QExgpZyA5gzXg6xuBTW2EGt2q3BGFdv
uuNoImV906k84z5xsjkQNr8yMHSGdJsPzcbE16kj3Q7/kl9XzkQV7JcdYRdqkOjG
XH7OBfhYbwDVoiA/KIKsS1X1nNomIBZCj0jCGQCboJkEi63tssDH8S3OlqbDb0Kk
/4oYcZjlLcp+7JHOBq3KXRE2vprnEKEX5FP15NLRm88qwjHF5SAElem7eUVYw94h
h0dltbEoEZkfvES83+r9cn4j5PjuCTxxzqBuPaYlC1aPYV7LNZeIkuZ+V1k/ii/0
bF45oHrmoUbm+lT3Ctn3LS5j/njrPUsNBLFF6asSHNPmR3HQYN4beo1MFpt0lYhp
cjt/m1gKU/Z1tLEs82HJqkEfEpp2UhforTrTW3LL/1pLUFJxOsOJ6r95HFoXAv1f
V7LIgNRFCNO6URuBsrzleSzWJaQ3y16rlXLbWSl9ichRV4xtVfOJGduXmpzlY+nL
ES604vYQGnd765DNtsjHgPN5hystbQPX78TAhnfyWRu/ZPS93pgcWnYrKtOAZIfd
r+sTCq1XO4uzG2JE/DyjYdYjj24ABPXq3V15oCkcDiixLpC/rsWU59LOqVK2OHEm
F5pV7UJkT5boeOB3V12EI3lXryqlb5Jtxnaoq7Q4taVC4CPh2r5e0NkfgxPkiCGB
obRrSDj4tQt5mDhBP7UBcRYyXP6aUoC0ep+lnYfLge4zQM4Kw83lVC4XAcfEHTAB
wYRBa9KoXUtwtUrVNjE7svQa6I+aM1uV2DuX+O7q15wNHYc3c6GrtbaBccsnjxlX
zwdQKxU5ns3556GUXNmINACMbF3uL9mx5VMu1daeih/UdBk+KjLTn1lyUMGhUNPs
cawe+UKYOoi6CaqDouMi9aGJ/sT7EIlaxyP99mhDUqv9xW+lLVy8OxjxGET4u/30
A/HwI4W7nG33J0L+kNOfWLoKF+Rjlq6xfJjbKq3SbnAWHc8Uk/DBAYaVXp2ytylI
HsZ0W9itYlqA9FQsmpRrh8NhbYHvRIKo+0Uz93MvQFuFvpHG2vptZI2U55LnCgp7
bXgmzAWejjKTGbrbFfeoj1R+8D5yTe6ebkqtVP+OpbFC+93llfH49eUwcDMCnTmC
kbFIHXbx22vx9cEgjV39elLNYw8sIktND15ZJquS30Gnrr+u2e/YuAIH4Yn2BiI6
njH2Ll52gPJSEddCGwO9iFb7gRUOf/TabgegY4V851YbXbFDdF299KCQ/skg8QBN
I9AFLYr0GDDgtMNMR0nbgBgkWYxd5xHKDSjyEKctCn0/UaGw0SzjSYbHKXBwNGHX
4SxcIwYT9vpG6pyqHbgeEH/ZvC3h1blRIreAO+jYJWMOeGJv+UzdKqTEqSctoO2Q
CvBnVlHgZGVMIp1B/fKN0Q/RZIpK7guG2j/ILxgH4TEw6HqIZK6OIuOdeYUBn02r
hbP7xeVSvXLDBt+Ad3wro0pFwF5HHa6mqrcJjLmy+SrtEcXMRT7v+grcmc/fbXFJ
v4AlXCf5ZAn0pziYzCUIeKMZRIQ9WjIrTdzH95WzsWzc2lmoMLqxb/YMEl1V/dru
Ti3+N/6LIgzRbue8RPNM7Z/piHRTLAg4mtHHaVR1CYsrRddY1DXFNNa2fTCeEG/8
gbzvXCTn2mC4+BzJyJO/7MCeLvYfPH9+ZeBUC0piiN1xB7sdyLrKadYBtb/S2jJp
PiJQby/B6b2hFl37fLRgiQbQCFKw/9Y+z2KH91eipMjVUbsp/4V0OF9BXBRsEtwT
GyEoxczbOJstU7BNr8kwEPIlxUmjtjE/Sn6Q67MJ9eOXp/ICHMwMg5eX7mIKpvYV
FoosUlbwEaBufnl36LrupJPcFfwKAtsx3HwRgpXlKaJYRPm1bKkHAT42EgSlgYdC
/KaAuwCqztHUdBFucsQP2+GIV/ctYAUQgDiUBtzZ3HkIOpkoXHQyQVKoGrpyD7VB
73cpDsN4CrtFCNKK5n4O2vIYxiCwlI9N2e4ZTf3qK70PQB1jhGBEhHrfhZfZpBiM
6Re004mYhakRxMIbAox3uSi/lplbsTqmy5ctjcN+uXoDQBbDhkmQlsIggFC88xG1
C5XYaVcY4GdSC+l/4z8JGSBwUTxK9qg/htgd0NMsgWiJXK5C9Vw+achUZXrFwQdL
dKqadr8g2SnaR7RNryjG2WTnzsng6ipUPUHT0CcYF8zAYPNx3Q36JlqyK6/40COr
VQWt/87vt6Z3ar4SwqWWFl2UNSishv/ty4p7ERh3HiPTwu0mQ6kY18yBv4NQ56wi
6Bf0eAp5vKTdv/wJsMyAljNdP2ihWHK68fEOMq7iQ2HEAE/iySxXsBTMvxvp0HmR
N+8NIOttOMynWgeybPqlEnNkjO7FiFTee79mOTy1MITr9+6Nz8j8oOzDH8cmgxWb
5ZzbCOYZd2qEf6HQwei7wmDESvD7dR4qe5wEm0wfsSOB+Sx4txFhc9vivLF9mgdM
Iaqw29hsvlkhdzVEgr0iXpOPc7KSSF8WttvdhN+bJupEmtxSFXQ+o3ebYyptmXk+
i7v1IP0q0D3g4ZMdSr4IvqlC8Hs6sTvquk5sDQdggExTDL+gfSJe73m3lsEJoAhb
dUQaGeqxlKxDyPu5t5gRCCJsMptXSVQ+gzPNopb/LyUdYTkV4YT8esGDnHEKYCbD
g/OYgrMxzr3wt9XiVKRjuRl7LjHi5Nl5VyA89w8T3GxKHpbiUgbgL/4KsURFy/Mf
9Rw3j0A4C6VCU1rXdU5gfiT17vjuzMkh4CYswzniFlvgG7Raf0uxBCK7Bkr+Qorj
U96R0lZAaPPHrqo7rZGe30RtPzKmz+785ArNodXsA+oMMtD1GnNKh6gHpNKZ4QG8
kMK3VKlf67bn4lu4hZlI4v8/JVM1ridFHTE/Rs38GUe0Us6++yrq59ibbWDrTlxY
uXu6BbFvib/tPnTvWLPxktL8e7YEuBsSvrUVFq6eB9saN+TR/ryKepGcGJ74NQfD
AsK30Ayx+jrdG8m9Vy/52wlJRne8nfok5SiPzLHbWecVW3DGOBkam0AbMF9jVDq1
7cTiJOjS7l23JOetbRNcrT7MC4RsUZS6jEjO0f3hKl6TajXefBMXeIDKBB1mFKQB
8TXXjXvzsfkhzJwhHwXzpIs61tlKu6PBZ9aNsHTQUcGHEQX64yxeQhI5QzORuJBt
EMybJ8lQpPxCldSj9zYct4HgGa3iPYLqaTVwNVc8lh4CciFLGUofMfmNWTZ6ezkU
kVBDpXB+ls3P9aSCBguO1JGdy+c2A6OISO3jtA6M8EY/MPZorEDRbCG+7exAx4MV
CWbovjuC1F+AJppIS539+4luzj8mBwkApWbtjCZXetqbLT+KJdQZVTWO2I7UUFiV
87kVyWXC/+bsQ0OeXGShbu8k9U/tLr4dL2frzQOX1Cb8rJuJIhdWfIkqWr7H3uiY
LSE6H+LK5IVaRXyV+M1g1hiHvBWrd18JxEtCUVjgk+UurulIGY9V39TL2uGsM7YT
Tip9DAStAOa+yYl23ZUseXewG0SKJo2GguqbnR3H7tBCvONmVpmTZsmccDLgRGp8
NRkR446ddaXETqdarg36EmR0ULjXIG7KFRnxPS08wbEww5RdFK5ZtcZHr707XIFk
dgGDw1M0q8AnrKlTGnxsBpESK3aKjqrQephkKWd0GFn9utNxKsvSKCERsAO8WR2f
6yZvtlp81EdcRev9zD57a9WmDsc/FXFJkOsP7sQ2f3eJ+D2sdznX6FkacxS4BFot
mSC7H16ZeArUCZznWR8VdSuvkD51/517qmU1AiElJOqLY/1KZgstNJxyNgc5NyJe
d6I7tEgiaHnxVUI1Jiccr2hGu+xyZkUVFMASq+zsAIEB8+qM6cPdKxxI27oDAya0
RIxNZStuMLrNpkZAluaYjvRJPWrq+FZOT3RNneVmx/hdjm2c4zugEh+dmDIOlMEv
2LC9yKtl4wwjyDVXi/zBtbgxnHSzMQatoPo+iDdfIMGT2la0BIZPp3jAWEr11Tw7
Oqx+aUQuke5tQRS+AQdNCVQObKv8I1Ebm3dfs2FQCKe6ven2iIsAnP+aJU1EIpz/
uF0Dc8NfN0p+flhPj7a1k8yjlZkvfTtu/+38G1P0ugYw2DQuZ0J3WPm9Nqg05K1l
TDe3l4pTzskCSZ1G1jGHVWS92tMSNGaRtLU7vncQ8hhk+LUVPn0W158+gxdtLStU
lzHh/kGbVLzJVS8HvMGd5pxZzMJrdcwiV56cv+PbaQfRE7l6FGLp64qJ8b76hvrs
cwvXQ1jvZfka3qoxM77ct2gWpS2N36Lfi3NgmXo9RDlU4m/EjJLDARA3VPKj7tGi
mufvPkOv1mc14WqwNNEtan476oD0Y2xtZkNRxS1CJpJXAf8h+/Fp4a980SdEyhTO
esO2uohNELz3JqDDaJePpGX6KJ0+Mg7UkE3qByM9u/l31P+Qra5LFGc4DVSx0KZF
/JAY3KxFLRAD5vMcZnVwoBdPtSGgPgfi3lRf9dRRDHfAE1je0pX3hkV5oKuqiImN
eVtCZ5ES6F8D8sgynyJkXeQLYCoFrwRewOxVxMMDZOt8NcmF9TpU4/pd5v2LyYo+
4L193L+u3qLN9mcU6kNtZ0cml4f8H6LgDE93ZEvu5Yr95zH3cEV2EiHnFod+0Z+N
k2rq26KWP+/Qsie7EFnhcZEAxbkOELR5RS0V7FgbzPwvJkkdNF/GgxUBQ8cWZfnt
WkwwMJIxBOcaJbObHLXYODtlS3UqEXc2q97i4lDfQjc5Ai0mRN3UuJup3XzmBuUg
3/LVLNlr6Uq7wb4zzlRugxgbnLyzBewl/snW6gJToz4eSRsJ3FyWGZJdx0aoEZKQ
9oAivUP2ydwdro6e/eHk7Kkc0vzEjdafmvuG73hP0QbM2VEDN/lNw+BvXQ/hs+Ji
J2HJM2P7XriqOutl+GG/KA/m9BAbe5J+VbmMsE3pSyUDvowO1McvFHoyjHoj1zPc
XX0pqpI2NDqmp2Yi/xknXhi/86jHn1egKiRoMqKQPRAEIsk4WFsbB8MWcRDTFIpr
mrRgLf+oLsHFfodiBKGHSWCTFMlq8QnCT6RW0u+5CCeC3SO3wJkp4+WPzmdZdcg3
oEW1RzD7bIpfCadugAgH3G/pzIS1f7WxrMXOF3HjQh6TMaEBVVnC888D1ISBiCfa
wkz/wNH3MRrTp6rU2uttjDGbemv+LIN4wYLQw/ENvppLgcgEB1DwIFOFdKNRWJ8r
q05IsBJ/hDoYM0neT3crpYa20snTo8XP2T7fqr8OoDieeMFVmE+DotmOi+qgKQGF
U9nk25BnnMwv+G2G+11+5rFKgeZrUEv7+Eva1R3qor/nKciZJFw/kek49pU3wUT+
LfaJwJkRqT42lje86g77MsJzgbA/yThXlJjnxIamXm84vo8X04XN8feosBGETmC8
3hIUnGfkuIg7x/UblDDKPyGvnRWOCAssler1pwJgMIXFNMv0QLXBDe6ddRxYdb7O
cFyCSzOpUJdok5zsRRedNiNs8aveN7ht9BKHcuSL9ubbndCtzdIkG/Ns+H8N+f4P
ZPKGC4r5vBAElEtIu1wPY0HbEQ09dLYzh4f90YsV+B9w0rTm1qazvNggcQcOt625
Hed6ouTtN2jC6SDf24HULmD8PEsG9eDzrYWc9mxdaJFXrMnofh9Lp+MdCWzlp7sK
iIyXuVst70qda8htPmesEP4baA0qHum7L5q79ydTtli7abkznL6q5/FoE7mz2xfW
uyddwEmWWmKnWbyn313XjNAjSVSv2154K7++UiwHi65qWSulXUKXGWS7SR6htuUC
JCklG7wRfbm/9NvnelTBvBfhb542GT2s87eCURpi7duxuAio0mFEDX5nv0a5jGvY
mZOvzTM9ygdkBWwWGgnro2e6wKyCax7B3iO7sU5QP5RIPZ/Ez5NWTsnFPUqWk+wB
8BzNVCkAUBHqe85WEG0N5gcA8XBUWo9+aGLsQ/XC84PPouieFyZjZxG2MewWvIUP
D8MJ2bqYDIZpB2aaA8bP79Y1lUFTpmy/vO+JZMrm4QD1xeZ/Gz5nleN8MChT+h5N
6xUapZ9Cfbf8WiStd5xis5RHOHZyjQQgw4pBrw5wCPixUmVbvINIPLhkeZXY4rz5
RiB7bk4pJO72UcUshbEFHYRcPNROazX0UyqNbeGLlkG4N5M8u+ZgiXHvW7cCGLo2
im094VHUf7B0rPJy9xfaUvdlCjAI/JK1qcs30CS2c4EZcX28o0ckdvUaIKeTsomE
ycMivJAmhHUIeMS6X2AtFatK50bI0i7JKGF++mA8rgUP4wVPyhizD8XYBE1T3D/6
VnIYaJ70Jy8frbXYMbXr72nxRmzCF4LGrd4d77bTlRkRHukfyefBIR4POjOK+E1K
BuvDaiy0MYyCV9XjQdAcc8p1lJR4V+0tcozW+95LsFHzZP8XVc5TGvHy1YaMHD6z
dDtAdyXOL7+KdoyN9+X1kAj2zDBizymv6kF01GzAnzwKpkBXQY8Joe9iYvlskXaS
pnIA9iLZh+v3fWodUwcYudbKgE3WJqByQ2+n2p9lGJ4Pi9705TkIOVBIJLfBohqT
dg13l9E/viIDcIBlF+n7Wz8ZU2YVld+/4gxb4Wq9NxIOON1beUFFPA60n+G2oHYm
9o+NC2YzaIgGOBwBhJIETQmM+BNnBi+3t4nbv01xfooSNhBUka9iQY7zB+88bSXu
DJNH0tJ9A9xWQgsgNrZX8s1Ydbd6X7lY7f99TXGmFDpIXyhJvXSOT7gMssDjB9+e
v0HLesRU16rJKfP/gQaIY/qNfK2yqHvpWNhj3LKbCn8g+2yUP1GKtGatTMuu+7tU
i3LkoyJI12+Gtn/Fd+it3YFoQQ6sTDiT8RNcsdRG8g/T2q9dwAZGoGdRLF7EgKf4
iy4gPWI9BiuEa0zBTXSeDrOoFll90P9Ruv6YHEYrS2YUI/KnkaIAfV5H/wuSf26n
no7FvS9aLPn+0XGVEMWeY3hfTEwoCTy6amf/iNvsGpGyKPXKTU0XDddlS2o+jC6x
gozyN87F7QqFg7XJY+6JRZS7Qk8S45eUNnPt3vVENkM6hkPHd8Lw/PcpAzmK7pXE
QuEo2H9TzTimHSRHW8x3HLICa9ODKj7ywjTor2P5hbEVQRUKuaCZsWW/8QF7MWlb
79gPg4mjRiUSiu30lPf70mcRHLzLehzatkK2g/kf7AxxYz0s8PsOAjIh3Cd+nOIC
9NBClkkEM21+1mU6fCk5qCeJiQjJ+xodNRCKhCW4c98FW1xWCYnBSyHFuJmRRzTG
UmQUSzo27dKfcmWJ9Tu1bdbSTbZwXkLoRIgINKmNf1arh84r57m9jHSm5HiyxG+h
NaFNrG/l0RsabX75WeV1sU7CREeK8iKBMzw/88P1927RAlxRQX7/0V8J3ftzXznm
NAjKY29cGvcEMorytfiBJAzopjBztqGiqDL23Cp8s3fzUGCXPrHnRT3BiFyeTXwB
JAP0GPkk4MairdXA4j20e+LbMx/zGcrNo+DSeA5nehIjNnphDOaW1p0TM9HsYrzO
TUUSZD2OP4XmCVllXYTDJZSNpa7HolRWGq0o5RYkL+hP7LMbIprlutcvk6L6t9ZB
cWDpaP6YJsS044CCXV7/paPadK5/4XVtGaxVDvgi259gbVl4qJb++lwm+8NzGEmn
KH41yxW92Xc5fw6ZUhVXcZmNGCyJ2m95GVKtT9x1kCZE0N4w70KfHOjQxPJAzT3z
4a/GHm2wXdug8RI3kPGmx3tIaw5M9IIEAugTLKXS/Wga458QZd4kMTdVdFLlHMcP
52Ypxoendp+4MbaeiHLGO6J+lHfgMaE4/v1UpYcQ2qpwC14Gb64As1imRW67x7oq
ei4h1UkS4lZGLF4B+V6dO6a7zvdROL2xyiF9dXhii3lbv25gcMi6/KnSEyNg6F32
BVS5j5g6Ypveq98zf5oJsTD2apT71SvQaIMi7fVIUdF3J0iVEz77KVH436/zQofn
DIXebgmEU59macByMR+qFGyViBonlgPYVfKzVjJpL1okOGdUWSim6Z91yBMLc+jj
ZVh0GOtO3KGS1cBO0Bwrf6NIvf/xGZpTA2njbq//gE61O+uMj9ZDGRR0ltencl9E
oaGgdEJ9z6qE6bdVhJibBcxJZHaWwRcstp56hW33vjpk8JNjjc3r0K1NM5brqaIj
ZPF/Mi7jfrgyelo3GGMu5fOi9EPNVcqy7pYxneHro2nVmhcXCRK0AGQDQJfroOtu
a9JiFpRrbi/ubGxZwXIeV2SJrZb5/syxQ0MlcQO8s4VrSB3sg3IooNQNBKz5BpL5
Trq5ezCYUiOoi4daQWDcScIp6WiWFuQPc+Fg6/wWYV+LGvgw5cGqyu5iQ313A8H3
HMh8HlHP01HXJA4vq4YK+bLDuDZYtlPAhhg3Go/wDJfLiwdKkjyvR0V6ylocv9WS
hYvZseFj3bWZSdh2UbcWmDGNw2rYUh9RHlVfdiBH9/rclh3hRenhCKzhufDXySYa
O3WaZV81ibl6wWqzLwOENH/gSso7VnX5y2DuTxybIlhxK7r2F1f42rg4Kifi5Blv
J1QlUJ9eNRBfE+E89TBfSkSMieWv9+Y5M2erim/clTgWz8cjh3oQdotmkoIS4+RC
eO8o7ciD80OiSSO6ggIrtTQx//dh0C2rb6WauVLR3jNHiVSq0l1BL6galOg0WIEZ
PN4+wt54AaWoej+d07UGv/W2NXXzVJe0XVkdraVmUxt2Wn1e9L1Y+/sxbJTUWg0m
sF0OIa0ZdihL19H+Hs9H9s44yVNZGSckWwemlVHwq6KE/3E/w5pktXwqor7I5fLS
KKN6fsaX4xIPNvmpClKE5/DfGbgZUtviTp8/s7MPFXXTG7LNKd5dUdA7PVs3btY8
02ggP1/9r0/7xuiXiZjh4yD4DNQI4yO2WxnTL3NphgrcaYwy3WP6xZdyh6Z1ZigN
pge6/IB/vYfmaGub/FsbPyDwQTyYnXvOR/j1XdtnhPqhUNOmilEm4ovqiEoEM4ik
h0fyORCtC0Wf+FF1mAkEy0UghtofkDB4WnMK9z6lerfU3pDiJT6WcYWKwLFuFFeW
PtRelLpjyidx2H4v6P+NMQJSlDdiqG1DcnCGO6rJ7xumHYGo0mUPvYi6n9/LYpDb
f9wZnHV4L4pG2oyfZ5v61mLGHnxAnJW9V5Qk8+hGgpw8kYUIFwdYfCAvwnNxDIsn
mSdmlaCg1HOQG75tlgEeVi5lEKxEE1H8RZ2JYo8HSuYV3rN7fHEvMpDc/YhNmr23
5gJWmvtE6wzfkxfC7T0Fg7etqQef68j2nGqvqVampkCc+m8hbo/7OEPJTkVzPQpT
y586z+mQu8AEhqom4RkLyywQLM7jdzEdThVm76iOlFOgUdgrEDKMbnQAw/DGtebU
y6pPR7wXpLpSqwRnUu58+uZ1FlUEpoxSDj0oCxfQqy+QCc+XdRN50rfZR0dRrPnS
yFs0RZ1BmU6wt/9W5cvxDyAktkqP2RLLqsEQ8Zq1asODcnYc8qIzmXaxN5tslzCQ
FHAonCbmGs60cjAJK1GdAcsYBkTSA639w56lToiL0znu38/D5kGsacMrrm2VXMn+
UjeOAq2jcjTXLo2pvKHU/9UWYEC91SHoDLxP7Ssjap3KCg+EX2RGj2RaeWLG+Coe
ywh+qBJcJGCVMtwF5OF8JeA9aIhmGa4ceCqazIWJi7VcPPXbRkE8Wj6NWwKXxA6T
Qx5gMzdCRWt77sL0bUAssXc5OkZ761cz5744O+aOp2chh9oH6ejhWIJ3xUGY2KXE
FU59jM6HQ+JeE6QTq0+Nny9B5xhrOAy8HSLSYLAtkk32LyVq2PX2Itjy+5IvzE6z
7AFa29lU604Ircwo+nu3PSDss75pu5ftFaB1QZDRo4hd0+gWctUu0KQboKIiwL1R
X1qO8TGAk0uMSdMYSysz2AnnODidk+5WomA5xIlXHmLNYWO+Gj9+hSOY4hwxQZ/2
8RaE79gdVPlK+kJMAwDOS/zFSsZHAiYgqF3t0+8LbpkMMO1Ol4Yig8soo43wKxnL
+XmhsJkkyD79V5SeJ1YjyhTUY2x5ceTP6InhRQabSwpttMyosM50Qcfo3l3flkUx
5L8nnz9+rg2jiqvJ72OTsn1tYg9q4NEHA3gU6bwPoy4Bsni5+ZMFaIvl/IChRY+w
Ve8SN75BI1vhlZSCEp2eWMf2Zmn2tEfNRdh45MOJekvx1QRPggyaMLFTq94dijJD
YroaUNWQoo6wYJVwD26DharkLMM8QgRZEG8/vAYhKYcNjfbUsAfYhptkuUYZLZx0
W6Hqu9SOqyqzf0CvEPEAoSNZp34S0lo4Z5uzzb/OOMsvcFPXaSLoluKwoyulYZvY
LOU7WRJeu+86Dn0NMWmNLYOY2GBDhv1DGH48Aq/p9GXMHQ+86SN1EYX0gak/N+Jc
JnKts6wERQKPtuD10izP9wL7KknxN5B1gRB2YNM8RIekapUCOuzEkAdZGan3SBUj
ITgzAXXE084iFN7wR8P+13IuBOzDthgGwBidg8MbfMEkgUxuhqhF78ouh/tCNES8
WHiJATbmwmGRsS+URjdThhhITc6+rSSeIP9xLNwdAgQciThe438uBwGv8U7dOjqr
pDeJbjLx/2uGxadhXotmbWNLMrOuGZpbco+RVz9bos0mVkSbYxFGuS6bA4yCx3qD
MCSZWLFaMEsIxfww3zlHHYGWFHqidXPMn9maz9cCKf4mC+7g+MioMHUc3CMnBq5t
DtdnD2lytc6XCPlUlqZqhKSaXcqPxnIF/KHFZqL8vbVjauq3D0ZP1rdPLJffr7Pt
zi8YCY8xQO2aD+BmMHfguP2nZR49uNrb8qCAKA+yZuflazz9g6nr8xLXIkQz7smp
ssV2Qsf3Ja/UTvyYRgCn7scQ4YnWLyThvUVTS9wABq46000sFROGeLaPACTkmeSO
nh0ZHR+Nlk8b1SwJUiWAmnDGLQVCwxOVgQwLC5rJM1dSPj9MZB6uU+/5yvl8bHq0
8Ci+8hQRPkQBpGarLt96LW6z2RBN712cAoaLvhW69wcuNc/fKvB55vXni2rXExFO
jwH2puHqw9fhlJ43HsgXlZluagZq8qHbmhzUGoaQFqA0P30Hjq1OoSkJUZ0vw2kx
IPBGcxMGr8l/q1Fk18Z9yID2yVRaG1ii3fGB8EOUyQHYXrpp62cCJwhmnXeBrq+s
WfYgQK0t47KQaCuYplrBSJ0giEShW4HIC/otAezS7suTpoGnuobxnQhi6kf6LZsq
XxM73mFngj8sKB20SQKAuWxhdaBRQYIj87sisrKkWUmHnYhLnGFGDVFmiY5RT8pE
syinKI/SRDM3ThycZIdBwNCc6puw9YcQZhnBRZZyGJvnG2kNrGHXnY8v2RaBrd4q
aai8hdqS426XrJYQF/vuY8Pre3pBGFPr3dA6drgOcKnnOHH7P4R8awwsJiXTX2I0
vDfZCOviRAdJBOwnbMdDIzEz+FLiqpEiLb0j7uR58UNejJSDrYyyVUwd2Ry9jkNh
Qkp1ubJCjEssKeBDasvc4dUgjebkBUZwCe+oXTO44f+0CwE+f5RtsCnXusv1hyCx
bTK2CYajmujKG5kjiR83MEDE7hgFdYKf8o7iUVdoOJJ4l8YB6eF6U9c1Jxmq8FI6
FP89v7FGpoLKOjvDlzJDeB8a+OxkyBMlOu6FXWlnd9irUcsswFWVYoMhWOsoHIBk
Z05MYJG2w6+mCte0eFKKyhzl8rEhEKV/Ly+gn94UBiM0UbLlgbeKl3ycT8QwYBAb
bdVzaji6dOhsZ+EG6ySGyzmtSvQBvQzDgfhRF9x5hNF6JozuRro3K8IhVgYY7sIJ
AsqfWaI+SaUxX78gwdp/+TAhuLngE62dLw4kJNtRJGi22sJmOVYhtDi6aH8utcUt
RS9wHW/9LnJLLyw9oF9HqITgbwjdC2SpdXYeN7dbsngHBsNWDJP+jgojNWNstfMZ
XjwL04Bwf0jPbLRnHpIRjIjRAaSK7Tdq7/Wp0vazQ55czM/WLXuQGEb+jD3Hkl0y
XTX5UXDpAUb35TSEqJaSm9BgNPSXAQk/+kXFUz+i0ygz0iobl8WKF58WkxrHXalC
fi+TQAMN6+Dzv6slu+KGNMmL0W5o4NtsqGlUaQ+oWjUwOPa4zzgqqKLHJtNbCQP8
CNlz59YdZIlocH3avWSWkN2gXoqrXzTrFXKxTw5012TV9sKUmZg1R6nOuJH3LCM8
7KcCfTNdlwFsawkZD0xTW8fGhwbT6FTEUki3f7YE+lXj06ln5cvFWxNk3VRSWn42
z8rBscsn9+/vXm7+H9YJEHVnlSiVmbx4VwGflDGzbP0lNkTEBero7ASxAVWWYilj
EZCre/6NwuhLQRQx9pG2fgsng6B+z2TQr72RhiZWHa7VVN9JSJHlGZRBmOEUS4lI
cTHppIyUxU7EbluPzYAqpQAkXWCQ25/7ZjTZwFzx9i2fFZaOY8yfm4YCig0sxm+5
LkCVYwtXvpO3/fOpTY9aLwVWSSg8kp4MIGK9QRZscRe9vlVnIGbYltZ61K3Jrunm
h4K3OPqmVQj7LypXDBsBs/mnh+zvACrwhslviUOOmeTZhV7FMaIUSxP3Hq8HG42g
JL5fk8JBoz4HiWup4K/XBHj/xnPiC8hFClDrWvC41RPm42fZxJSi3knCsOzuatSp
OOL9ENLH1BmdOiW9wpSJHCkNfzQZR2pVHmdx2XlNInMc01a/RbOuM94B+NQz65jH
8NntNg+sCObCC5FI6mcr3AgQjs8BjOGxXf31zL4h+Y+ueAmtug++SpWMeWqhDvPO
Ih2P100UBdKP75fqD0mHOyk6FnCZYP24/Dcxss6F5DEIXokrBPfyxkRH5h0xg74A
yFwjFYUqWnBhlZTE5tsox7labsMpaLXT2popUimtyq1vf6PHUElwm82qheOx0njz
dC1PaRnNzhPvgB/1181qJI2BLVZaLL2sMjB+DPaCAfz78RDtDH0386rxRwn/AZH5
jTSUhSYyPdd+es+JqDKDUFXcpDyCt1L4QkazPLbB1IOScExIlOOpUaOuhwazhxxj
0yRLe3NpOznrGHx+5dF1XvLb154hle89GD6SI5ZDglF7LP2jlqnRRqkV/l82/NI4
Y1/wKhEYMnmkQGQ+uua5O565PL0v0zZYP9MmMGrlpmVO09R64x69PJZGJvnb6tLs
M0Sm5sxkEqIjNtZIbQ9qf6O350PZUlbvTv25EbSeOdrCIwhCSQZSvrGFQrOhoGxv
DvsrMTv88P+56FuXZh8E8ngLiewll4aOOCoTX5fvfsZNtz4+B7mdVZ7g8PWfuFDn
Z1WUrXOAnVnhKqr2k+GN3kqZ8yhVjDjxqyVr9XlFY4YSjVv/ut1pXpw8WMYAwB5P
A8vc5B9nhEZ8WVot850aHu6ktQ/Kk5o/5tGxPQx737DRJbtIpwG5uQPNATmkB4jg
SmBvaBBNZOI4BZwbVK7nDFZYyyGgHuoz2ast6n1v86UJ2EZGndMV48Zer9LBpnK2
gc8UkTngH4GwfofhSX3ka0Qvm27ErN7tHpVXHQcsYW4td1hQIiYWky29TArt4+rk
AUxnnjG3ZFYjLYebrEl+rc4amASqpr/E2+Aujsjzj1AeJbZqEjsNSRcAAunToUhh
7BM2r/TlpUQh2l2wHm3+8t6jdt5F+AJYIWPNmIr2/LbMQzRD6DvPO7O0bV1Ea2vY
6rvbaP6nGRZrYATW6VjIotwQ2cWeiP/Nhh7HzHXiDQ42jRfcpC93X404Moy8IIdJ
ow5ZREHvFyuG5RTNm9/A9Co3gdvdTfwI8MehCGI9dd2nHsK/fTML9vk35Ludv7pC
ILF49hoj340in30X9oCqnEOn0Noe4mTJmhhRm6aZYb4aYvT41eWPF1Up0j+JyV0p
jc6tY7c20FHqae7mLEBYDotpvjYV+dfvjsFaW0DWQUbmEXzSR0TRuFHqRlopNzsi
xbIz+nNk5DvRqjFoy2p9GWRxj614+mdKmUeKBqjqPP103rjxjgN4DWeeioILGNC4
m9e1AaAoUU3zXiB/o1y+hy4HUSEWVajWXEHXntATdWnKsvfcQ+mSMtbLJG8EevmL
nGPZPzqDEyWFuX7x9wJoQ0taSK2k6A9QPPbS4Nw2qftbTmCYojBLqF0pRFVaQ/O0
`protect END_PROTECTED
