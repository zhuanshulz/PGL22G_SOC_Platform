`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7+OjfKt2l3j4OgjyWZz5muaFvcxKW94BcCpo6cvgoQ9aTS0x73n//po0MuLZC+G
XTPoTNn6zAjvBnzs7L9INOsjOy2jpzTOq5q/kTtPaHL7Jwssbz6UP+zB1d1hA5kL
F/0CwQ2dl4iQ2cGRQPVYaS+OZLiD8fp3CrO6uTPXSDuFvFgxXMaoszbT3PmLOKSG
AdThYF1tOSRKlH+6uJq1ESmgdU3L2S3OS1gEzSpBxNXA7qrO5DLJlMIoO/0K3Nzf
lvi/AqHIv6iijbueQxKQpE0PAuCSknq6NPM6V02+J5896r2ITdZv8y4RR1NT5cqz
EhEhp66mirysOjAxAcIB3IwzP4oW3vqnWXX0WL6mif49DjJJW9CbK5ryByWzMRhM
VFgDjsXd6bNDD+25kPigVozFE77x4sQWNrzI/eT0c/RIda+sB9KPN1Vq4RjhIPWr
F0o5V3YTDbfDXUtijC38Z19vQdf1NkhP/ANbcOCz2o1yIBwoPKj0kaamP9GdNpon
yqoTtMD/t/TPp9DBEHWat2OeVQAiOUs9/tosshZMT3ViVVuyqzLJcOwvtW77GZay
itpvNm9iYD9Aa8PkbL9dsFeKvH08wtf50JE6PsFDL8QeMX5Xq6+x2Bf0s7Gc4csy
XZw2a7ELhvYwKleK/p21jbJMVjL3/+6PrAi+Ly17VeBYQwR37pFwPbSZKwMgFhfE
POEbpkuVTAJObIhOF0+nh8SeCnFRVxWWQ4V3PwCGYj9pcSXzFiIQk9iNc0yxuFRJ
4eUnvUTejj3sUFG5/H9llTzTNSdGIJ1eezby261o4L8Zuz1cJil5m1tflcGV5QH3
tJpghiyfRP4k7al8wwq+CMZRFGEQN+KuOCrcrfo0tBp73+/hNfKNglVEc0Kq2IvF
BWBCumdzwx39+zB076djpkRUMdAC7h+xvKNru33L8fGCcs1xS9w52akjfVqoHGpS
NGyNyPLdOt4B6p67KGuoY/xtwJatZ5AUEEY8amO0sJOagxYnFHVHUlBm69DqKhLc
0bOK0Ult+ktRACaWFCFd94FL5hFW4V83Kh6Q6dfu0I5w6687JImuzju8TpdkMUmv
T7VVSefhCDJFOBkFj9IHOJh+xQEIYlP0czeyLQT+JD7eLH7nD7/e1PXnphKu9twc
TZQ7Mk0feh45aD7qGzE5mVMkbiLk97hV3Mnkh2U8DLnmadUNUw/46QChlfW0zFx1
wTki+pCHT/TRm6w5LcpA9kKmXbfDfF6sbH8Km+HEYdPCX5IvC0T8qEChq/wz2dhi
X9Zj7XqG81A5qlJNzK8u9n1smgcUyIIg5sLpSsqkcgHIMAZqyzJb+pMH8p19DUET
ZrlTJBBEu3o9QaClJhB3+l9MH18KFQEtRGiz4KiPSWD1Q9xVtkAY88LA/oa+9TKs
wn5PXvAbP8E0EP6hvYuVASzktaA5JBQDIO0mQ6pO0NMn1uq+crGzKMNqDFJbHiWF
etjgn78GsMsmfAQsEnu7YdNHqAS5pQFK2fXMbLVUVsknTQKK+B2o1OFcV3GDd6r8
tySEGhDw3bgY8aq2ho8ZeTVbW8FgOv1OrVgfK9LzXLb4qFTH9aI2u6qIsd4V+lag
Lxxm+FQP0r02pIyauhDFHVhRpx/i3P/p8/ANXqdoz8ChZRQijpuwD2ect6+SPlm0
kLJxqyjq9t8Kaxmpte9OL5Xv/6xHiFO3zuvQ2QfVBNtrLmKyyfISdVbj5LwOrxC6
vBdykDNb6Ac5/rR1ZdQsN+17QX0iF6aoWHBNCg18JgNicL76mCw3MS+mZwTaCnLX
E29EVvILQJ7Ti2ZfffVszqiFOhty9+M0jQlmQGmc3UZSNq6ZLf+R+lxymlY4Yhjg
JnqT2RQgFpSNcd5RXhLeVT2SMK++GKvuTFsknIvXeh3bLb6qufFzthvOEDl8OUQB
JcfMEUYlKoZt/DrbjVhggKZu5KQN6POxbO2bbYglym0qK9LrApt8cwPLWjggraBv
Qtg9T6xBH9YSpu6guzWsXaurnUc/HlKhkKyB3rnOj2KzRz0FX7taZsyECdp52KpG
B1HVqNF85LPbNRchxD0up0whO4+MD+w/+ErtAD9RI1X9sCjF6D1iwoY1Ba3KdiLZ
Px9UVuCAK/opuZtp0ged/XqkWCUxAqIISnnCeVYMsC2pf6g4FthZfwv5dF9IXVf1
Qmd8F2x0g1OZ/5JlWuklSbciFCLoNA7Q79lawG+YBmiZ9COBB9NBZakKeP7nUrxx
5CR3KNOR/xUxOYC0MNkjiDB3gtwn68Id554pOxXM2E8EKaXfgqPtvw2N9uDHqpCM
5Ez8yJmuB754+WcmLhrUdclbSe35V4gHe0DkWnreoMN+UvCRDow/j7huy2BjaLOf
Gh3je0e355lAyPQTFuylMyM8goc3Jla5xXOVOu+RTO4SONkECtGn56HzqzUUtJRq
cyMxmKN9ooRuPwI7EASLqM4N7g7+Gd5uJ7sLhzmOO7QXD0JPaFj1dcDGrmxf+AT8
XEt5CdcWceRm3w1MwzNTf598JMNYJwVmZq+09sa9dfcj5Z6lXpQlrW5HOHFrNReG
wjC6M4BCYTyFvah2BOGamkogXspDnz/MM6UIYE/wHYuuIDCfUwgzdezCGuGvS5aZ
g1/sOrDWYCB5EpkdRCB9LRu/8k0Zjde6VdBZ63d8HiUlFC8IPqNiYw4TJm9JnyVi
QMnBjuDRhAtU/PLAV2p6nBMcTmWqsqUYk4rwhqnnkrAophfwVQ+oUZ0IK4B0/xwR
u71WB38fh3fmRNkTJHhqQGOKtLP9pWum20yFmCSNrws2Eg8B2XRBv0n+UPNYFT3x
8qa+ZXPSsnE2QeCN8gbw0roaC2FFv2Q9OFeFgTHTo9RhZMDRjn5zVswTaQWx96FV
5KzkIw7AnnOz2snQYfrs26bn6SRyC5AIWEoUpU5pSzyPPD4g7kO0+fs9eez2VppW
NjENdJvordmQBtNcN77RuWALgsFXrQVhaRH042/cZTsFftGSSqCPd5TyXHuw46Pw
QQBzQUS+piFzpPmgGXbAfPzACGrCftsWwApmhS+YH+MlKdKSLQqgQkjSqa7ic1jS
9Ik5EeovaB39XIoEdsQlJzUUF+WiRijtb+1qHgJU4ZjWRutrTIOEPlS8p5CKzBhB
tf/hAGq8MLhGk+LE9HaXtRZuFTUNQbsnbsOTxsoSooqmbHtprfXo7ZF4StcwCBrz
jN0WOCvkWU4vWiW2a72nAd9xvUcAAyXDzzMvZWcDEHqYgsoSCtvZzC4OiSJTR+YT
wx4+gPrd3uHcE/WPunoeKwVJvk5scRLCLSSegOtuUbaruT3BvXt3QHpF7r86wCVw
dtjxD5mPH32mSUfca+NItVb4phZPm7DXbvL4Ud/F2Kpnn+FpXJURCx8scjZ3s2zn
iBnIyJnXtnBFvaZ8DWgIKdxB6c8Igw/vtOVO80qwB1vQXO/n2pZvvO3+4wRDMjQF
D5LyG+DMLfVWoeT+RoDVAMcJfCplxMk5gWLErlPlpVNYANEgjpZ+mdgpcMprEGMQ
OhpR8E2efTNvS0k4bT4/4H8rlsBDvq1B6ViH+xrKWxefWS75uNbDRZEPzozJcA6q
lMsEP1PtsPcImrKhN2oxrZd+/Bf+yGECDrvJFX/nztmpNs1NEDn+J0xISxCB0GSu
2Ndb6TGbAC5udf8Eho8P0RkVqNBkPFi5a9Bu6YSHLDkITljDPmzrtg4JeeXKZWds
rn+oGedUA2ULjw62qHXr5D7eRZSxeIabfecX3F7WrNudpz+EmEutICK3wCiYvOsP
d8T1pHc3wDJmbkupMyJC9f54es2w3eDW7RRe5n0hZs3iJL7xJvHVR6oTfov21a4Q
ntETJDGT3Y7gROjlauxaHQ6zueiRPpHmsiIYQaYYbCVi8m81JfzhixvtphUPFI4k
P2HVTTholC6fS29rrRFi1cww8UfdCQSf2RdAfXBuAzmnRJNn6IyIJxt2xXykiw40
bRocbQi8v/0WOUbTR24IMgRQ78nguoZwiZ5HyAcg6X6Nm3NIfcgLIClcTMfSL0t+
gNilhUQAeIjThgBkSisB6StdsuZSzznSO5ijnxMLhljpM3cnJ9i31mTaDElZXu3U
sbZKYUX2t6k1JTNlxnRPYxJXkvSZMMQ07PsmunAToIwA02VVratrP4r9BOwENrSf
SDgAvwt2iXpsMQEVjV7qkSssAHW+xO/Mki8qVqGmV76b/gkP9OZ5y8JLxFRCQV4X
EzJU1gYmomxrqcm4lMfy8h3mZ6t81QlvL9wP7Xvr/15gNjoY17w4qBi4xPtZshvj
qKANxU3d8vbgjLvU0fI42+9v7yeu4CBkZOoe7UPqG9H4PHRAKU4OMziwWRjsWdly
sLEe/Rchco37/BOoUc6eqMVD1LOTj58BZoGyEYzjp4JTbWH7Av3uNxj6V3HUXD7B
Z46SRSJyUGwKiX76VZRbgcKHvpvoDhyXhywisDESVWljCWnYoYkw5xYawkW/HBOq
8UnFbwDXhKV62X8OI/3mKQ808/1MtJGp0wNHzjHywhbfkWzJjzYchc3GmnJfVyeJ
eIsw6yRkpaTboH8ctpYoGzRdfd+GFbns4WeFiJOyTpdpI0sqUNzDbif/ygzFX6o2
8UUiXf9VTShsYzzenSb10zYcum660EIhq0qzA4u0rMA0YOD9INdiPu/QjnaSAtmJ
DPk5VduyI/oyw0hQ4SE8VMEv+2GY7IFe9ciTgs0MC8MLW9GQvkud6eMf1mKXWSDo
NgjBlsKw050jZPW0NiM5iWZQOlFua0sx8fxRcBja2i7PPt3Fzex8kqRCKMd67uIb
3AkAlwuSeuc4mnITWP8+K0TcFzyZv3wz6vy+qvmiL6e2XGaCniR0/j8f1xQcObiP
jmtt/JyMkFebaz2DdlPy6Hk7XvcqDi5KFERevaywnplniTHfX+Lsj9SqTf46L09h
Hisr7U3xUsrNYaTf2iNuL7/7U5xjDpWd35Mwovr1UcyzeCNQSDuGN6u6ssjfKr0d
CZOuq9emVvJVH2nuGU3v32UZBKCqLuJGEXk4y4wurmnVzbM6zarZLmggPym9GBTR
N7x6aKtaHUTU9Z59zAxOIdqN8Ymn5WsuDlzYveuywW/9YQiW/Zj7QmdTd4kBUiC0
VeQBUvv7f6tP6iIfr5CInewX2zXsmjUIYGs11+UwzFj+Q3dS9SaCnBGxAioaH9MW
npRujSsHpmVFCqVg3ltIXosVaWoTfJiAHfUWqAOVHkaAtNo62Xika/8ADB7HgnaR
aXUlL2FmG3ZPzUplFvPivpSTB6BPGdHrMSUwSZ3NaCd1fP7A0HMaiGiJSnrsLKi7
J9N5sdfVl13QXvV4YgYZPkUdCCpQ/kxFWji4CKsewEEWc76iWehciFAweZmp9LUR
3oXE1PiqcYlV8wZWuDpigv2jrcMQB0x4ZU6byAhOwpnSW+qLrEh41KJ31yGKGlRx
6/4GFAG8PPfGIbDol2w2KZp26dY7SJ0aF7BtHJO5OAcNBAVhEWmuiZpg7yDz11Yk
q14VaFiQfu2mK8ahXjIygVV+xkuZK4R6k5B2jY55iHTFfycDD5V4RVR5BzVZCiPe
X9YDh7Mh6rJQwCoRJmwjN2qIYa8+tkQWAPxnncGypG3/KqpxEUxpzY+EsGinhYEY
GWhg17bDpdZ3zMWVaCu8/wa23N20aY0X8SC0+xiZF+ryZyzch3jlFMqL1wz6TeZN
Wdl9cClXHpZrjvjZus6sgs/RtUFBmHgKt2sIAghvcsZneTV3n4G3i+HABWf3IHwb
mgESNQKSew4sUYp7Be/ptO7+2v4sleQ6EzbcwuhUnTxuESDMnQoce06PvkYBaHxD
2YSlsDxbem4f3o99fiBIbE57ygEde3NcP72jxGxRVThs/SFAMakoR3/rDZaMn5J5
r6o5ykyjCZMtuD/YwHyFwDnfqD010S8rMEyMe+ojuZ8G68ku5nUMwiX9NfiSmRCp
dPr0D8Zbi511XZSNrSY88vSqEab6bhJNA+X4KocJ9Z76640ubpnx2dfuZTqGu9xq
lp7K7R7YqGvRCmx2G7Bbhtvcdhy1jZ/pyfJX21LSNz+esfknmMQnyCoTOh+1qYWt
E93QlvmlevkjaqBtsKhwMQ7NLmQXo65zm5G+soYpALqsBm8PQpTryOIClFtx/ZeO
5dsXdqCIfbsckDt3PXSAVksyV/ocZ3hJbvO+6XhfP5fgUzNvw1sYKXuwxbs/2xVO
Et+BLIcCOAc5IVkIXBac8fTXkfbRJv7+Gruq2S38loUWyftrbDvC/Dpar8UXpx/C
wulSbUSHLUzEabblt2Pw1KK++qDjfd2uJr/hpTSzPMxz/Okw8bSHpqZfAIQEEyJU
y4g9rsuaaXDPCEh9MbKzLiCwNhDLI8meAV4IKTGslcT5ehHoNa17RBfK3vM4mvy6
+uHShqHeY0iVzkRpu/BMnTUi1BVoe4Ali+dOkVc3U3Dpf5LM4h5XM8xfSJp9lMfz
0lXm0/LMBikbho+a9LrjLKrSFn2buWi1RzLw2gcadhjXJM99D8aSBriflCHUHEZ3
YG4ssAlDzOvr6PHUmpPZ9qv9wqk3J6AUoOgv9EKAcscatALDPEMN9jDOq0XvWK3H
i7Ggx4vBBsHLNzjLrpVEEcBEnmzbCJk12YDizO/GTO5fSG5W6tvDn4fqnJfMJRjh
9rgBK+OI+phFSnB5v4KpzH732iSmXjTUOCIeKcLn2O8oAU48XnlCO09IyOuxzxo9
nVaPlEHwgutEOEeYZU9BtJ6Ez35gqw1NQB2ij67qmAgqM4MmWe34ndC3prV9+W6N
ZJ72KTGyjwI4GI93G+du2lWSirhLZGp0itx0t7LNQaokOGSr1bB7imi+slT4sW/N
mOqC2OPqtyIpGtl1/Sf7LvSmqdbgUwIL2gELoNHYFKskNgiHHQnyIldiNt1/YTqU
dsoJEqZamcbqGciT8BC8p9gyhPo9wtKQb7z8JpGOpMzKsfPLCMK8ucYnQvNU8g4e
+aRvzckiDcPLU8OqQOzrd9nBlAb2KU4lW4KyDwXP7L3sErIfYiw1SGxVAV8HkXo1
S8A/uIsjmxtdqltrqxqI4oZPMFwOWO+b0ic7dbLmUucxh0mrhOUVTd6smucLksiH
H16aXfwcEHkka9MhnQQfqLgueEkKMQeCGcbcjl06QplGNZmqjVbYxJc2PbMHpfrP
YLCcMhxsYIKfVQRD+yafyNKImcaLLm+cyyuTTx8CuHUgFqKsRU2AqerBtNDPJIol
x6DCSzSuQkwWJnlwcKlSV8etemyFd9qxYGpqSdTWsvlUkUHKHdZkorlcvuiqZcx1
GVIzAo750M/Pp8uAdCceAw+jODQfutZFlDhwRADGU8NolyfwtDpInF8qPK4RDAk4
AU6qMRmWbsOzH3qszTyAVdAUvSA/3nwfTHnYO0/8MAuxYs0HCynRlhGsQ+4Mr2iL
cQUmoPaxp8e6APjgC0XwGTwuL9TvITfwar2oA2F0MLGnkGP1yTjrSQS1BeSPMn6o
Ax5yI4ZQYQnJVvS4i5LkFjw1vlAwqJa9+t/lLg7iuLIRID5qWOnxYxShakpo577M
8xg3iuY700ZS2NjHcYlfy9f23HbWrJvnaiHCxXH/AJmIjfnQeAW3PJ8Kd8y6Mg5X
avRM40qb2/mOyPZnp5v71geSCimcuLIfVbdcyyD0dWJKvl1wtsKsL/wBlR1k836J
rr+0ctSNxjBdlSWYhpCXv4EC9XlDkH6I3KkO3ADVVbRxNnm6+3vnHF3V0EnUvHY0
Ki0wCSw5xjGTJBnkx027+7wN8YFAmbjoZhbWNlBQBJelzrRWebsOz0AzV6PDJVBp
ZVXL+smPiNk0Ohp0E/82XT7X9fyAPpfxflImodNat8L4ck0Yx0j3UwwxnU+43zl/
FRYOjP/0whgTYmPF/ouKP5GzyLinJzndqJKmvIvajVm27tbdrrl4Nn/zjdFdcqMQ
9JQEmqyvCELaDWJ38nwTf22tu0uM7LKAPrsoNmupR8FLEjwyVZM1aWph5J8L4dto
cHcUqPNkGOJPagIpBdsoXkSZXstdcujKTMBSc9ht8I8jSPu7POHP7BnERZownp34
/01bZb6Cf/BMW8CaWnBg8klkzIY874/6F9kBCs2OeNxWZ7YyS6+2YTQw/Dwa6NVs
tsvFoNsMdIsh4JCten7dtHgdvg/pbHoW5z/zd4rK5pI8skcBTNBT4iR1ZX/xDHVX
2cWu/ceIVkK8ufftiO0Q3ZACu9NyVPWxr0OfelEkZ1sXISIPJqKoY0/B6KmYQOpC
WmeB6tTmqsaVHE8Su6j2MsZ1LhJ5h3fhDbeD901sRmPYJAh8qrGXpeQeoKKHDYHj
daiyqHW+mNd9Jbni9tSlLQOmxVAWLRVkgkFJVYU3pDTEm9gvIkvCdFRPefCEQpUw
EWDAGs36g1SlNJ7lhV3Dtj8EpXj4r0OkFWEx1EmwwatI58iO8xYPN2p7eWfJwQsx
IYrupYpvLD8jAQ8WaWc9bzrgofQbseapJu2BfBG55kSRuuikklJxuJo3IJo9ZnF9
aaKOp+MSrolEoleqyGngzzYnDW8enLvJr+fS+eAeO8UT1I2jwGdBAb4WuornnhQo
oMT2tmCFdwBtdoIuOeUAwwmUT0Zv6tnn5QGPChLf5pC7D/0Sg6f4+Oe/TpLfS+iH
t94sE7RGrs6FSCdqn5DEVIbntVZjV7j9+9ZRS9JfUbUcJWpJtRD92V8H7e8I+81F
iDpe3IuqXQ9ZNqBE5DzqN3ZKlDiphVHSh6Qkr2WNU5KS031ED87TlM8fTNwgm+hP
ES04RgPgFKizETIhNCqGgrCs/pdf5rP2G71auhJwcdbYGfCN9+d66VPRBeaIJyWO
iLhJxDxn/H80xAxvn5ma5M9N9eMonkMNPDIoUltfBMcZRo/LriemfOiMqUOaXyQk
47K2yTx6HOJ4sCgRIRVF7LJgOeeqdw93BvmE2hDsNm4ipnWnNqUu8ezKCR4WQtFs
66xDh+tvMZCyOc4fUyf9kfu8ewa3szame95TWtmdiSJKmLuRGMKqrQQsjM0BnsUK
xLxgNjcvSKrHqwMxrm3tFP1CKaF+Oi+NMeNhG31yGxJX2Xbbv+PSWNQxXgyQHXNP
BMiM7QBXwn9VjRUb4D8WPvWyy+wOEfyOGIQ3c0neD54Cat8yQI89yrvc6adxF1BJ
Rv0mhDQype/mQkfhR+AOsR1e/MtYw55Idt9Fj4GTSP+YuangbsCMhu/svkx/+bCb
TkOJ87ZP3uQ7XjVqudscTXDw2wrks/v99XwXWKb9pL0gj3tpNQj93e5n/SGCUGND
44trBLAF8kNWy3PmPLMEd9E1wMdpS/4y85CZDsdU7m6/wKuyEJhXwKOj3X7ua5C/
oG77vMaobILc+hAmJDRBNVOTieTzGTNtvoYr6KZtf6lfj/L53RRD+KKx3kzpNlPo
x8xlBVqPgKGgfKsMjUo0075gOknh0tRZXaBFLDQ5voX4fHFm9fNJvd9u6+Pgs/TQ
7Bd1q7BrdIAkEQYbO4ehswQ4suxohPjPfRVPUcV8ICr4/bN77GptTZbGNQCijoXr
+ggjP7Mnsd0/y29PUIJwultKkbX7cL/Y0C9Z+TPipOH15iYaJPJlrGMjnMyhIzQ6
JCsSWTnuXlHcdkDf7EFAIzdyIQSPuPKeh9UsAeohKMV3muBIOJhdAEfDTxHEjDig
iPZ5hEAE/nfUupcaV4nXQQyJw6K5TQIQLqdy/rAyNNg2DkrMl6tfS2ziqqjTnDtH
83S8+gMctfDzk4Cc2UMRnvlZtFoaMlscMTeF5QwmLIUALoSyo/Hg23hAnaMOD+z3
ACHmddeGliegNEfrN8rAU5Tn9ghpgMQqQ+BSfZDi47qzN7bvViyzRuGgiNyNUgBB
OfjP7lXlOHRfWZ/e+TbrIOOl3hHvJ+3fjyWCcvk1MD8IGQrfscnSDW4d93XkAS1k
zA/5Nj8FGgmvkUzqyUSVzkBwYApGu13XUK0W3HI2NiJM42IdT7GKL49bJhUQGsxx
dijB6LlXZamfi9v0meH4izh3qp5ODWtya8HCejjWGla6OkO9X6cCc2FtRU/ymSNE
/re1uTiZkQ3Py31SMKaaYx/vuMPK7RNfscPlvxXVDS7GM68JH+ePwfysTsjGYA3+
MSU8F+I4dWixUpkxxJKZOTrI6varYIGPbGGEtwrMUHG0E/vZLvNzDXzaYflaQyh5
F3fi+I7U6VrGI1FacpXagxWmjk9dVUNu6wDVTG37GFH/f4WbzLNtXI3IZOoanqYr
6rAV/fGTYITMhIfk2wZ9EkK4hjhHLK8PJDuYhWWk1rNSObOFiqR8TMNNEkQRNsDl
0HcKlGEYeLlARcxSmjiD+iB8/4kHqJsJs+E637m0WxbHBQ0+xEthDFpMxW5d3BQt
4wDveXLhG2ohOqYBszAzyKtIi30I/qx6Bp2mVZiRoZ2ibGA56VBacWmy189JV5u/
fzXbQGLqz7cI89wxQukPQ0XGV93pln71v6f9w5elCRGJXpzArmyT/oJgbzLrYMyU
qsuuKoxxvPnD1/t3j4gH8dH+PSL/z7fsj4IoR7x9R5jPqSc5PF1ApMgniR95RWgD
37SdvlNfZ4HC+MI1mK6mC6s4syfvTF7xsT/O3vzAnB5up4xwjKoOlt4GGe+VS4Mp
KixDEPYluBo18R2wZhZwJ3f/HwAsJhADZdQ5oL87gGOec7KVzVOcE9rwPuUh14et
JY5AGMUfCMRVMmc5TAYWMxkWz/w8wmti21U926UwDb4BIxLfUXxWZXjIHykIXoQV
7XeGTrErn5UpiyYXiKes3yW7/nxPLtaUcY1EfJM98YWocCEnhMaEBni9B4fFQQ/l
oeuKEIlWpqFrZEB7Uvx0D9QwdNqWPcNNS/eK+maGVBjDTUKeSVJTkODFStCmZNl7
KbGhMzLoch1zqF9yuFTmOygVnpbFGSPlHKgubyFxjd4mrchDzp3+a79GTvnO6fyD
4ky+O8aAE9HYOlneiayRHw==
`protect END_PROTECTED
