`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFGgtiH7JxvQ/xiLNFZSOJjSY2n1osFKSkmZMlfjVRkiIgRtAnEx3Cq6JquIQLhS
Z9vXK5mnXYjhK8vj7l8JwyX3mGCrDGjXM50uQ/P6oFHRe5wsEMq258loiTMCgZE8
vQ+HNxVX5m/5d+TcSxiI4pwEzuwzycGtEbtYVHobuLS/lYQWwp/pEOmQa15mw75J
msI8ZLZR+9Fg+H2+rzvuQ8aru163dCQPwiterk3q5heYzQFBHL3Z2AEDM0lOoZDh
c2DVjRj+G4oSjWOZ70WgOUhWB5kbJIvnx5azVSocVMKOvz2zT/CzMUdcafVnuo5v
N3CVjVTlnoLbm6kXmrAMYKADsRe3rdVDuq3Spaz6BD+mfn3TPs9aJjjdc66CvCGE
KsOblLb8/X10Q+qjkQfG2V+4/rTwrNNx22sW/mgAV1mdyWfepLxTtISgovRUlRV4
M+GQtH3zHCN3TjhXG9yYyrzh3mKP+YOVkeJ/Q1z1U86K/mTaRWExXUePcGKt8OCt
tQGbZUNdSuplv0XNaVokLec6Vl5pxe000O7vSTFC68AsLpPthDANvMRlFYnI7N7A
8S6O3keJsXj8ABK/HkWtGCkEHlBj+EVQutI5RnPYiqlfJpAWcoME6esSDS4BK6Ow
w9RTSCJf/TVx6cRNHVR0g7egYI1jTre/Fm1XvDzw2Vpn0ZOshwCqRX7vfbcsp18j
QLTosgA3VGF6S3Koxhzs1cy1x+S6HVYOg3Ntb7dEEXPDvU85Y4XiU6glVU4f6QQP
elrd/6hetlBP4pV4BR+kku7ABgHnTRywlkwypyfTDmptBqxD0IZn3KvdRNT920uP
alhH5RdwXvpXrXLXCnYam8vtDall/Primf2Gjl5Yg73jPB/ah0GwQHTUmjj/DKiD
JbJbFKKg7RFNvQDVs1D8GXGx/iEIakqgKGcDPbDPYNETl753R0vFBZvhc7+s1Chd
hwB0jz16nYbTObpjNBkb2oAg3u2pUvRKiN8HZ01+9b6P5eOYTw/LaWCaFUyXhq3K
M+oMCDe/KVX68YCPDaZcB0tHM5Fg5UqOk4Ym6b76rYU1Q42Noa5Q4MjBlkmGukO6
WpT99+wqcYXEca4sJp0UitFp5JehlCb8vpnt+VoVFMPbbXD60819UizDaENNARQb
8a1MFX47Qa7khtqCbEftcxLWRV4QtPRhtLQfD19AZouqxqwjkjtaUiMYkXE5r2E6
GdIyeS+PxfKWmoavoNnDwpGWEzbQpFj0Qhdh41QUof4qtRqRjik8z3BsrGuVlEJt
SD06Wc26xDSSWtd2XEORj9MP9CHGv429T+QOsQ/Z6rNEk7AcPppTNOQhY4GocCMA
FuHO9P0htlfR9WDGmfHCAMPYOWBOK11uCuz5nKnza8hj6ZFzDhSVIGrHgj5HuQob
OVo0ua8Bix+hlgntG9XvufH+O7lUxU6luGz/amBOoF6kVZ7rZYi8N/vSNB1CUuB4
dMKqFx/vKgxmk7nmoyYh0ICwrFlvOY/9ZgeCqy88ZmwTPbanR5zY8Uugudc15ei8
1bjHN4/BZKq2dyvRcEMop8N9CL8QxoqdkMangmw3dmzTRSXQ0dhiinyPRjM/cwU1
NJo5rouRkcSR2SwGSB14e7LOh3N2D06dF+l1qj6uMu8zV2wxVD90RnP++f6dD29d
DfMjxDz6TxuUKHIRjvwvM0Tqc7feIQVNfIMBftnS+hfF5tYY8VbsHDFE0gHLY+iK
fX8PEn0o+cvbEDrmfl+MnloKP7SmJV80ttrORVFMthwgr9gHWib2T+JspJ7Sk6Zr
A5Mctepsb/BNnn/uQ8sJ8z5L9jKi8K6AUoxdVj0jaqYXRNxyspgNhb08teHz78UU
5GDB9Ggc+RuVGbfxb5Kt4I3gz87UUa6nYCwnA3u/v8+Zwm02FpMj7xRmLfZ7bzDh
CwQOOb2QkXukNLKZaUQeUaw1UJHWC1JbLIOwwVP0dKob0wIJ9N8BNYxU3VP8hicv
23GevJFf6wgJPNhCG1fTfp7h8oyh1kCUL9nUU9zx8oiw4huprwUfqoVPm78Ljh69
BFqUNEpCgvqVJ396FMz8sLrHwD9fjjZFvPQOViRk4KgZU7aX22D6IWJ+2dhqQbro
nW35dAwqOg9Pi7KYUcuQwdU4Zmo/RbZ4oa9yxa8dv3+/g9+PwuwzRoQIZXtkTQNt
oD9GZmR/+rnz46rrlB5957fnNfOG3ZLggu7p57YKP+EeHAS7VdPelgUYfD+rkH+u
D/h3OFjfTa5I08p8VxLPaHUSqTdEMJO7rtXs9TAu+rP77mDpRYT2f0vxED93q87N
euBU+N3P2F/ktLU9lmUZL/GBv1ADV0qlppWhvp7wcW8//HBpDyxYUBECDTzqRGiH
fIsI21vWBxEc01jUTtD8rnPdmgHtEfTQRdMifolfstdRdCo52+uTXcEvY/jaI7Mg
PMCFku5dfuHK3e69OxNBavPxQYcwrhzSxMEvr19iBlGzrYzBJ8JZ7Z8P4TwX8J5S
Ap+B7/yyrcPXK0Q44RvbgP3ZvUzXbJqCFgYlPi3aecfoi27MSqhdhQsrpE5u/512
eW5lf8hefuao40E/LqsfTphTVXasLh3+hfZYDzBfUlX/VI/hmZWMdOyC+LytZ8yh
`protect END_PROTECTED
