`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ACiME7pu284WyV/DXwg/ptX/uhMs4PgYVpfLMym8r3FNAaqXdcFLk6iZUBqFFPED
3U9AOl7huKrIbApPJtIXGlJkc3D2uD3XXtIZh1hmh7vLt74kvX8VoAknHNs/LhJ6
7X6QtNOxoaRUXo67IGQxQeg1zDmR0sLo9eL6hwyvhfr21Ykz3PR4mtity93fakY1
oJp9BA18YiMvnr+99X8wkT7oG/HAP7BMG9b7tkDa0AyeZ40UEgnE4Uyv+bnqBQvr
ei1h0zp517P2Mm1FA1SA/5jMYNOMvQ4mE74GAGqXjpk7B4ONi4kKOrRbSTZ9dc42
01QuSHEnMNtjuUefQh2NigAVhm4vUp4oaj5dRJtFv0fkrnxiUvT16FpVIh4GNKJK
SFrxitV3uizIt1AWgGiUP5toRraT4Yu+DaDlnGIcGmXDqw201eokPyQqhxecgUh8
1z2RHFtfTESfsjX8KBPnf5jachH6w/JaSXE8UGBc+cWSiJkFtL0ULzkUOZTefEuz
XgHhQib7UhZ89aYP8GmdYhZCsLNjuvGSwApTvPPz0mPgtv7RSI6qPpnTO5oX3tEF
91s9wXD04KACJRvp2P2tSTYvXOK/WHt5M+5N3l4MJoTbNhz8OjL9VJ6rnQPdBX8R
ivHIZ3nQT0sHzbqWRy32YE8SFTVpwBQx2F6ZLAD/dqicQG+n/fMjRJUJZ6n2KSzP
`protect END_PROTECTED
