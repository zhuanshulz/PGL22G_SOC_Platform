`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k431VL5URvrgqQioF7X0vyQghLqxLSWpGCY8sYWlW0IThvBYsz4jpzVCF9boZSug
bFJ61lNZJpHudKOibtr5ezMBNoZy4ORQI89OGwSNMpxVrIMYTKWU4PRDIgxj/sGS
+W0/xGnHECkDbYMvdNykMUB2hiKUKqNOOFwSTrYa60tATejd0BAqB9+uEW4f/tDP
U2A1u4v5i5/o9BOuZnfCOK8K8OXF1N0QpWc6eBaywssMCgchs1yLBBbC/l6nofQD
MAULlDIalY/w7Dg1hfTe1dTVcesnJtBck2YfYQSw93IvR54BnCtMtlfw6ADWV6ZF
oH0/YS4/LNDuslkqC5qT57r03Sis3xtRx2+lCJ1JNqJLUax0GauD4mZq4jopCgmJ
L1P/NUmQ/7yf355kBBt38ZkVh7JMlgDoOKsp7lbpO1YB25R1t9YAlTWnzttYQhfj
f5lCjqzX1sN6wSzdWc2f+ipzPmchvneVFPPgBSgj7v2jhU5Z9xcInEWOlNLm+fJl
J9jxL7AvfrzERWf5NosjPpQAPovgFY/ygdO0tWHXiCN0JIV9UJ0oW0d5PxTcozqQ
Of6iInB7+I1RX4eKtlON4fi75Xqbk4TJSAi9mY91YIdsmGtEau8heu0zdxOp989H
gabGhu1sXtqGTzTdbVljG/j7+S87xytNkT2S5ww15v+jILtyiS0nWmDS+LT/zMBe
T3ycqo76aYWNRHqcanSn3R1auXHVZtinRGIS3H5ivJkjydlgmzyTutQn0+s42VTI
7O/00Rj0nT4c4+q931gqE09I/re3Xce7KmeWR0BWXDNwxdROapGpGB8oLbUwcSI+
wgABfh4qhEHDHKaHX8Lp6Gesm9fda973WkcU/wwOnxlOAKwYao2edfxlQ3gsmi+m
45Bvm0X5LCO+gkWIWYyJw8AWFXfcabof+ebQKl9lx212o4AU3/WFxXsUJ8BsxxBM
WncKBXFL6/jE3XiNvQCkIXg2grnyIPOYkbCewpJjNIY0o8tNigT/ZSh1MjNQwAp2
oKncVqfdhsMgJmeQ503Avswvky2nFM9rRcpzGMMlNFYHb3BNntm6XNXvff13HILh
IyzYo8iyjl+4tzCI94Cc1Q4BuE8Z6dW0VOk1NXcWpar7Ezk6pvDtAJKYWsZvsKQu
SMkB1aoemSz76rJRTcAdUyKmLatrutrwwJMz2A6wv/79VP5FksTZNxGvy/cupvs+
2M7ZTJayosgPkCZ6+Dotw3kqT2FneLLgCXTdtsRo2RTeK7faFvLW6KoS4HJFKKmm
ge9v8Gil/f5wynSAueHum10QVvoYJb9ZW5/7ZE9CLDYyz3syspg5XSayB5Tkhwfx
nQRWINymScWQrwryBvBo9Eb/eGAnfXbWOE8BpIlpoLxbLG3YngwlCFzjJeqHimDD
hbl9ep3V4ado8Oj3IdW/qLVUE5WFmnXfMkNwT0xXGZ5H00uOlVsfgI4KhAi9HN1n
XqJ1z4NYDvGCN0FaBnAD4Q6lkrd+S/jo2Ms37Nzp57pSbhHtAbmogb6Ae+qqguim
6GmZKVlSpeuGHiXEYjRelOxhWAEou4Cvu1Zpcsi2XfGQG1nGaz9kQY2oI8yCNuIa
uo6hiDtdvYYqomNz0VZC7sjyIh35510Ku3W0pFilj1UBwtaB/3mHRM+BNf5OMU9B
cvXdczo4LC1NX/QjUomXAaZIzWK4bbANW0ebjoTDeJTz+6hLLYnvbn++UT+DraIm
ovRHEqCqhX72tUJlJk/VPjzwjn+N2UDib58ShWRSf0TPLW2Yg+Mmwrsc1qKXE7mu
/GGQE0tXnnsoN9OGmeKIdCeAb5sxBGWZjSnuuCxe7uVReRAsRSoYf+IIZo3Kgnby
Axl6f51BI8S/ztZ+tQkujYDTamOWGIe9VZuMtNao/3vxEm+/9ID1/VDWBWm47llA
LjXWLVkCSBkNPgX8oWO70UYnNHy6dlOae9WiTQiGbktlHT9Xh2wsWkRif2Qut2Yz
Uw73IL2tlctdx2Jv0SQf00KcvEiGTR1hPpFNIAXGVn+OlI4x1VwfqofUQIwMXRxh
Qi4o3hnvvbMWn3v7KKg5jwJkprftqXnBby8awH5h8u6CE/P7Uyy1iU//MxWu6543
UbGUvOijwnzHhc48VsVCVOm9okNbu5G43DQIuwx04PVwGy9QjuU9HdZn1hlzW+KS
/Wb4TFqsxmkVUrKJ0Tw8sjBHHZmptm5UbiIjUlaHloKj4kOWdnHq9xpdnZMCmO2d
tIJXghKRnmFfPTxsV2laMMQPA0fLer9+lCPOwQxHErwkvmr1UdmznRq8AWB5IiEH
fhzT2oxs8Y06iDycq6PFt9a4ou/E/4y3g8rBoEL17oYziE3nQqh8uRCXhiqxMnVY
3I+6LUFSEGVP0UJK2rvHHwdbUCPVVTfDqYK8SJSZLqU/7HxMFJHfPC76bIQVrPqa
na1b3PCp8DpbHjEj1vPN2dPep4nWqUleLX0jAAb1tKbmUqEl/2xp/WGBJLJkj2SF
0xpnNKzHlPxvV1RWwFDEUgq2/4Zk9g15ONysyHGoJBnIUpq4tg7/LIvSeQjX+kTH
wTgiFKHGmXM00/6tvkSgmwPsH1Ho3rEW8IfowzZQmicj+sentR37kohCDSYupk7J
NKLavROenqpwuHA7pZbGtdNpcMuUNrGDCYHedddRRj0VxvDCh3HgAK0bbf8Y25np
8oQHEIkvdSmjLx2ebTECAHbvUMIC5u00V7mgDRryJxpBDAjQ7TcMwK42mHW62hpU
kENoHkmsLRGJKtFLoOdMgCtnHNzxniLCWAtF+C4AOOrdE/PIllXAKZXpMXVHehTe
zX/sfFLR9aL2jTQVJZZs7n2+ggfGdn3jFvoaIhpguQV8XawMqP4u+OwyzFecVLOl
VpYHNdVN6EwL6cUbUaxTZijTiKoWIoG6ybsDhfOE6ProBuP4suNW2CJrYVS0YXY/
JWNwr3N24Mrf09SB4Y6vZgOTXWM5ipw7dcYGBTDOPXwk+YWM/YUbImJW6wDzdjrD
Rxu+ARGmXUL6nus0oTosQ6qN9Ly36TQ9eyc4Q1SJwuWoEAOmmp572RJdH/YR9UG9
11pjoEk7Z7Yf/PS22avZVoEgORrAFJCijrHbRbgnp46cg/leKbWOSXFanrDWgcd3
YwjtcCHT4bbyP0v2Nl3eUgpMvAKShMFb6cqoqmlAlwHsd93cQa+vtVviNt+F7dsC
2zmiUuxyPXJdAjHaYlSsBxwPDj0MRPYCmaa/ZNxntqBuybms60+tuNFNqdI0wkT0
L74eBWweAK+MsIpard04SK7M/M4gJmdInGRnMtCDJO/HOPxGkjcMZkCrFSg4s7Pp
UiOUIIK9nYXp+Ic3bJHMIfJhGYPA/V8rEvya99BZJGZXEa8PrUbt3bzcrYM4/A/H
sYa8e/Sb5U4zFuvkg96if1rJK+fwnvb2mlKLFgkLzFl5y9FsxcSNMnFZitv0wOCS
JcYjK+GoeYkknYb9uuTGDP/h1tEvR2g4bty+yEJnfXSF9XI6sNL2Fvy5o2QkJeU6
YhEKF1+Cyfytle+xg0K1OttZrppca3+KEdZk8EZu8uQXVkglpaCISQC94Cq1EqQd
KVjA0F6TbnIYEcuA6/kx0mVeroJp98RiOPcBe6pe2jBt/+YTCqymkOh2ulprAduy
OFUaTcYjgReCvBECR2m3JwvCIbcLvXsKpelebIcHY6E854Mm6+NVXc0Sd0/Tre1l
D798Xv5Z1KMp+TptiSbDMUeiR/1ojx0DmRds44PbLKHTqpbXJHO2E7jWffgT8Ap6
MNpwtCUfU85bHs98q3mjiYPzR8Sfu/cfi4b/VpOb6rCHl+rBgu9le6dsMXh6ZySs
L3OcDQRFY8lgwNUsqpCWob+i7h7mw0Mg1xUUFKZZYvE5LT9WD6q14g93rOH5Jm62
Z5FxGxj4s2ylsfxrmD7NoJw89rfts7oBrIr8TPWQEzKjLckKpKuudk6vrT/TLnKz
G0tyQWeK4v4uDAjz5D6JDdXiHl+vjfQGZlIexyzyFQJU1htPCxHsqJFSWLdnxfyj
vEdKr1jfXwOSalJe/Wgp/j/TBHaTVzmCtCVDGbybbW6afWLzeamAoXVYlvh7OY7J
61/8dMlVviQpqWH2KISqUbQPJTm5DrPNGrVLUFAcO1XpbwzdEAwneg6RSQV42pm4
eeslS1y05vI2H/gHo7EHmOZ7E2o+pRf6Gx1i570CD86z3WuPQjUJkq6rgPK2T0U4
zKMoWSZ8FSpLHc26GpQbd0ZDdAfzmQGx+WTM4H3mW05kyoKJ70un3y7yWdlFAQ8V
HYPCeaQDjNuvZ26CTGb1cO6M7KHJwYRT9gId6ntjbsk=
`protect END_PROTECTED
