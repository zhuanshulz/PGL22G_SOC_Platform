`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnxJ0PbCBnQ3+9c0YDcTnS97weQos+eQAJae+YLqogncJJ9u8/k6D5PpUxZ9oPqy
ldInhMTbv2V2DF4bEIMLpSPMrecuOXfWx9EmaIsOfnCCH5z6KmOR7BtwbgLQlB7Q
O5NlV7lWQ/r89VpmSNrlQedGSShTbss936INAaZKQlinfkIFRaGk+69xKsM8fB82
oC9qDbJ4wm1h6AcZBm/zLcFUwARrhs7yigHpChg0st+cqL2CPD3eos8s+RjwmHJ8
vbiLj7pv/O5Ll8vmAbw0rKFxNwS62NPoTvNZbu3412t2DNfk8ZrTdaLLGmaPMj2U
ckYHRiJiQRCdukBCgAHmRdT7uhed6NiYIIn3d/dOwsjs99FeykxKRG2bmnx5E8GW
uqo61BN/jV05Qzv0VtGAalcgEAsMg1W1oFYa/XzUmL27ue128TVaxX4pMVR+Msi9
jWP+SacFpoE6nd27QIi0iR3Xu6XWCD5eKkPXGCbJmpdkIuE23cxlSSFi+/3rjL+d
tZv+mc1GNRoYjl1OjE0ltg==
`protect END_PROTECTED
