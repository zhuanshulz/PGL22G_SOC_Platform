`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KmiSbJ8vB79eJ8st2eBsP7AClYFObpc1+j0jcPdbs8ZA7g5Y9tc4b8GL9LtP6Koh
QikpMdjGdgepilF7jJEfBYNADdMTqK05twHc9o+239HE+7xwGH+SRXmdONePpNhy
5/VNAffrtBU+NZMyPwexFdXd5rjZ0EjekvUqosohq6EmZepjq8e+7X3R0AV+BXiN
Pqus3vkTFyNaIcNyKOlwiOni2+UDAi8Nrhz56kX7NhISlx2ObiHoCwbH1pzFc8G9
Dj3g00JwXNlM8FhJexrnXLzVov9PKQB9SWiHYNsmNNv+nH1q6/VhBVgsTM/j8qhW
dkY6tsrlHrJDLwAQnlWhpXGWqZQ13nxiX++NmXtxXw/nhTdFe5MzTunHM9x0gkK/
Fps5F49FRZOdRBxSxxpFm9waIW+0TT4xFTcdTyTW73Ih9puxJ7jH0HtEYCMlINw0
Niv5KGs6plNTQwaTvxLBp/aviB52OCdIRGWhq/i7o8TcJLJkMFdyO7lbYLbOEH/E
Q9L2VAu19/oGZMgYlU917gBFIHaqYOiMDsL7NacAO6O+Ag/+oy8h79Rbmr4FB4XX
QcXVUBz12juYcNefg3sM8BBnat2f9jKfKnGxRQJbwzJ1WpecgHoDAQU+eGEl4SdZ
+9g+/owa+5cYrc1fP7I7B9lbejeK4G9fvMoqAP/pneWNZMA7SFvcegR8j4xRTXmg
d1FCGfFa4GBOEkbvn8K0I5kbtnXtsD379tQkb4M3KU8q0FcN8RogMfS9ZD0i2RwE
af+4/ZMthYZXBtFUSdiEiROMFpDignDwlWjC3sYA5yqKP2ai7kb80NU/GJT3Vg54
QZdH3ffFJ3h6x1kKHRDasJzbM7uATeSrnHw9SxdRxySmBH/EjX96KRU2d3Y6B1Bl
PsPjKz2+wM6jVH7CjKh5mZl/k8k6+BYD58B4UJYcWBkG0sINQYmJ59/DL30up6RJ
1eMvI+DLTEHjDK+i6mWbmbePXblxf6namlwYJjhCpO7I67VxRqwdXzsA4b+kXNz7
jvaCNdpSnB2Hy2eSpnuODJ9YzG2VW8M6UpYTjgqeQbXUTzDX9+nFcHFrFM84J5w8
0B17BT/Equ7CrqNgxk92+71E3rfqBLvWstr6iqeD6y1xokgss5pzLVL2speBoBfY
Uyk4UHKQOwSx+kcfh6ymE8r4Z793/D6WWu1DEAdiAitP6vJFjFMOyslYOpTDUJxk
x6y32dubd4UhGHTyFVULfSsSrq3TMs+zqmHXRuTKGnL0hkbDFQmxQiRYwX4IqZor
4rwmzD52r3DQFeXg5ckqcmhh88x86XVWQQlElAVxtQh56dTB7U13PxJR+K6xUrnz
tLW9/murXpXtCToH596y8Kc2B0JLU3g+9F2HQeD/2VRwFEx4liB1xrDN7IeSpNtl
XzuCcIqu+IHfzZV/lsvQhDGbl5OH11UsM02ue8EO/9ROBHtNwxAHyEwUsg16xn58
aD6QkA+Dc2URNEzmpghY/STbGjKsRNd0NA0r2FnUPIhhAEsGVj6bKUKfAoIyz/cO
/QxuDd8S4j8kw35zOxsBwgajSb8Pp63Yjyw5y4LKKZtzz7qMsAzW3m0kN3eLjnjw
03Xt+70sTvDq1J/Vw1b61T21AFCb1ptft5ew6DOP2B5ABf63/jv0lET3uyFK+4ui
ZdmNwu1xpk24Qzrp0B4EraX7T/MHJktDNHINvFkB01sYaPGU9libxplloPR16bD4
bM6UwlQJzakj65AWZ3thi/y9XjjlthkNGAFbtTL1AEY2o0MF/Pzcsg2aNU/tyVVA
If2/2mHQO4KgKt1NlHGzsqYpGpnTNcQ4PPNBHkjzYRbHhap9BqwuaMVCyjqcEAA0
PnWE8rsYM2Ahe3piJ/vzjZP5UOlFXuSfGgebWFkpjA7IYsv646XSlDUkjkAa2Xlj
exiNLLXuTlWHmARCA5PKlBZbC8Hd93aHiPKxygtaoRX2VE7KgpX2vWP8ptpPdjB4
z/G5gBUomgN5RPhKxRa2BvNjvypJF4nUL/iPNF8eCgU+l0K8NE/x5KCeFThAdHqu
MNUYiUeTApCy1ZFmU0BJTXtIyq6d4EQo1UyPsLo7jHuQ6pfhkxi2eq8YNFzCmNmJ
nvlBCJK8ARqeu0xw/QLuJe7E6uA3gV1oRQSWyFRUphQq3KA9OMGdHC2d8/nXTsYw
vgqvInfrBdeD6DFpGHcYp4qbSVfV9opj8EK0QyW1p5jXQ2E8za1grsMps/eNsQxs
FwECKXCtmyAvdtAaHPc92QijE8P2OvR9JgTj0lD7i4yr6egpV4GvLjoY/ZehZXjd
Fb24CsOcSg/4lvi6b5E/NMzaGPaSyHZ3Ob4iaVSJWMF7hSnbarWDJa6Tmzmv+9r3
RSV6Lg6KgNLmtwZrWRQBdsUD8QIx3acN3B3XjUWYmynm/Ifviq/g6Ge1mDLX3jgL
iBvDkzZOHLAaFHtxZPFf+vLjVzl2Aai1DyeRGD0pcaHwBu9wLSQaZk45/wRwu0rV
AaUIcdUrdlXUZphWq+YdcJlJC1FRbYgGRPk/aBcrewQeZEE/qD9IpDi3uFi+uCum
9T0RKZ0rdI/PPEnCJWvdLCqrsc/pMSxpIsA/TJCkayKNjXl8uQuk5ipRAn+nPWiF
nG+WNvkCb0eQs/4nATO2jSrUEm5SypFcalWgK4Jn0f5MPTRaA/xYcObtfOzrqawU
l/sXlkVnYNcoCbOM06+FEhpi2XOFmRI0Bjgs6ucgihj3+CvJ+l0JkWarZ8i4PUXX
rhXHHah/z4Jbw+s0wC80+8q/FOVOqP12/1Ib3ewGBAv7NUVYOfqvc9bGdJjWYmXA
3vjffqKeCKAE4jJ8km++XPaDczELao1W0oZKH/GO7osr1J1fWjDWGKwewKEji1hn
aNcNGrTwE0lo7FQyvwtV8BAJ4Tn8q53eq0bLlXSLElzf128yib4NfMBPh+UCeYz0
tbV7xRCZl2YoadThD2Wj+KnzqAztiTI7h2tBtwS4h2fEDjNzBx3WAfcSQYyUzsxs
Oriv71kE4hgqbG15e64Ne357r9tBHCPFJgFGpgoJYKPNpVFfJREDFdUddIK1cq44
moB+fcWuIc7vhe6qADwf82BgKjRuTckVmmyUY7nJfdihXuhUeDtUT6vu3ZtYZ5S2
bEJ/YvV8cWySOjyDJ9p/AFYtION+phDkdtvxm8bqg7eeDF6lk2ZkmeRrbCfsA55k
/8sEc6NznX0VPJxG8CT+BpRY8iQgLq7/qFOryKmKQ0EfhYO0PNplPLOrydRhEVIR
HEm/j9RwEfgn0MzMg6Ap2fCx1OFMKT5cN3mvcMxWXA5dopar4pJp2F02xBVzMe3o
VVKNGAbUNKWwE/QYZ8q7siuPtPayD/xW7GHOMGMv0+gX1GVs2LA72+OXUtJ96gjq
ROluIcOLI+/ZI7dL304jotzCeP5niuLckZ7F3eSg2C2VJ592L1tACDfnEeUfJprE
ZLggsEKyG/36CSvPBv6DE4vocGb0YV3IfjHb8AxPnQUP8bthE/C1qCP58MgzysYC
Q6PRh+Ehr1sGf2PSZIGAf5k8x0yPHoYhRE8rtts1RmUs3zq5d+G5uc0JwMDri8mb
qGVSU8A/UM/HuTDywtpFkccD64TjZhr0IEcbJkcRnU8W3C56uFFaQQXZcOykGkEv
FgI8fuldlMWk5291xG58tOgT2V0Nsjrq/Q7xhOR1GK5hNncNcrUBKxwRQ/FBKHKH
LXQMinbIHTNCDMIrzGvAx/RbmTjHEMEA9JsQqBshr4y5m009mwFqj9CACswxpzaC
ZSvQxFT+GBS+adUiYikMLhPiOb1tDyc+9rNR1p26c6MXsSlcCtW7T9ZecaReKjUN
q6bSTVKy8m3tqoUilWwT9uKE2HK7aHASNYAyNpmwXP6F8A5WVCRgiiqMjLgMnjKz
0lfwOvhQHQEigkdooJWS3C0Fbaw+y3egkVqA5AFwmvHFAMeoCzuQcz0Sb2m81x77
bixdi15m/+MwAqVcE5DhRAwN5RmwRsdobjJJRX5hLwgAtvj7R+FjclBP/VLz9PCm
RWhysf+qbnARs71DrNDbvgBBp3xQu2KuQJl61dTO/4K34PPB3fc5k7ArsVDIJoUV
78Z2Xoz9RKCfqHO+azUTVO6vGK74CthKn8QKytpn5GRhOiPUup6SVSTOQLgHfaOz
EqYq4hSBFGmJW9/eMMKLiGVTrcgmg6LMp2USWS1uIQmt6f8FD5Ub+F1nPxTC2rHm
8walo4Kh1FuKfDXlXcJaWbqntEd4mTaSGrrjcboklTQOlCrQoc+b1tP9oBxc3cAw
Hbe0hxE1Pup8MC5+sA42HkfrPAUdENWguBicQk+cQV4gxeixxF0LWK/BH4fkDLBd
bmcqUgJjoL23nKP8zonBaITXcEgT8zCk1nAfUdynkzpCDSEI1vG3msNeCZQWB9Oh
lfJuMND2HiF3ftJde66Oc4/Y5qUV4vimRijIBSkZnCNz7P3U/szsY+nxJGJ7xvHl
y1WDZWDOhi/xUjFDp/+NgLSoO5X4UxOFIWO6FrvfzaKIA/trmxGIoYOnlyiZ9h8c
6iJK+f5jVpjS52BJD/9pNamtwkkrH0WMhq/KokWx3T8K2VzjpR+QDo4sjM+eKp1w
bgRqJi/QA4s8j3/1dBbKwm1/BAFNna8ugC9P54qhvZfZrCfXkI6FlU5VfowmL0Ut
R2R1D+RBuHzy6d8VX1TrLYvIG4PiPtTXCNRw1cEute1IpzMfT+YF5lMksJ7f/HGN
Zi9wTb6CAP2CPW/+YYr8x3Sz8eQtHdmXyLOlfdfBujsc/9mvLQjnyWhIlDXFLxwg
X1/mE8PX5SLrz9V1V+hZlVRyGemaams/vVTLYaFaKgK+8Qb6qWnCs1SmI0hvSQ3F
ONLID3x2ZNwBQsI7bW0DSaRhbndHAtPJswG8uFiMEN+mdGQBEMVQ3wJ72ClL0soQ
/KBFjVP4lRtXv5AWnYm50FYKjx1GSQjcrYfsj18nBXAiRvOUBxiLFY8nwUlAN3pp
VwMF8GVFgvmIj6jq/VYNYpDCzt7fWInXK+u7o2tzRLA=
`protect END_PROTECTED
