`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZ/F1OkWVvwv1irA1H7MH2ujEoldOmqOubCN8bcYB5Upgi1L73UW9TB4kIoDYL29
cnJXazwc2cs5kHyT0jTlmwUjzooqird8frB9+YDav2DeluWQxoHnaUpJeNh3cyHr
hyFkLjO0pS2aJeLF/o0V8cAuCG6VH64cfiXfzirHotiQDGLdzg/OdgYh5yJebfJ0
qjt1YOk+h3AttXnXEx+X76aEDPme4qPsZr6m29nNljUhlOXea05Ix7SrH0HKOORl
M3hzq2IFhKm4gLEZeNvYeNM4dzsnrWHqjWdMdtDl8qiJtcSrx5Z+doVY2l90cRLZ
Tdr92DdTdN/tm8QWaW6Ho8LYtUy0CHRl38/TtPrUXweRYKAZ6xS26qaHFkx2FK1y
B+m/JfQ42EXeKMZO/5W1yhizD5xaJM+c07IJG2uAZWfD184cix7N2sjxG2xsgCYb
EKJZlMg65fX7e2r/ERLs9VE4l1duq4HbdnHy21F06AYemrkXxSZ2OZkyepg7849d
d6hgTDOch2Jqqk+ga/gYXNej6XGuLsSVwN/52MrR1tdr6E3UkGSYovymp7lfBfi9
yYMX1ZK8PcLxk93iRQgBX/Sacy4ajQ5Q+ETvWt+z89KZ4WCSESpaHoKnKU/2tYiJ
CRtM+FbYk9Y0ZaN/7W7djH9MaihVWQI185bcbQaMP/BvCX0/8bqQj7NYdNDZ7Iqm
hCwddbCcvuuAEelCeumLZE9QZU588Tw9BZfR7f0RWC0MMFWlRHRWQjYs9UMswO63
5Nmtn7K/hCiRvREM5qrfwV9b21g7f57mspwpZbkYS5jQiyPzrwHcB1/T6WoTVZTV
a6J1UKTCHNVZi2b6KwEa0BqG/BS0p667OHETBWv8Rhw0eeW2ssvjlPaovLudgl3b
qDP7G6sqXfS9v4onGokbFez7FqgSw4flMGSpb/+py0oDktPK7Epc6/VUfgAgsK6A
Ld60RDhwtAsah/giJUdwyCud8VjSIIU6KyBi9fH5zgbhpB3svtdDQyZgKSgUWTgG
HK/nWS9JQNEaLhzg/KRcHE/+venMLWwhYbIx5Vlb7I5R+zieWOfC2ecy7KtKiNge
`protect END_PROTECTED
