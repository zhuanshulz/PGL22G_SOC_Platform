`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8lbAgcnBGojoJfnHfJzgCR0SjmVNRVMWG4STOz5EXFa0D3YxkGj6BcjHyA3/HlHE
8O3IoxJshDT/M/2hO1TUJwJFO0Tviud5LR5B9As29Q4DqUvlCsM5J/wh1XtoqajE
nzcTG57yRMU2RQ53N0O1k3nuFd+tRl0zpK6hRz/m5TElYHvzvafDg1bI/mLSzpiA
6hLFC1ZO8FT21EhQTVI07ba6QKCnixVagJ7PRkYgavumbRUSBpKXsjeNfjsPKIno
4cF10XQlFpJSisQOOI/p/bc2fWW7JjstljMY2V2qtuRRWD466DwD1jXotBLUTPyj
QEUb9PNu9dnffqpctYGiqdMSjRmh2TT3aTwiIyXMdsXWNsL5Gd3uyyyilShsum9c
3U54ephI4cm9a0Pq7weYSkJCXY1RBOSmycI7Vh2D1NS9POfpy3jxJ7FkBXO56ivl
NiUUxK574urQhxE+M29/L1e3on3iSEAVts2U/8Zq2LkmyqwwuaH48uEU0UAJyBgh
jgnvfWuWj3uxvE5zkd6I2Dy6nwHkP7K4gB2mKdf7ZKflYe5gMBypLBb0NafbmTLv
rHp9p5TQ1rbZjBIhaMA490eoi+PCx8OgpJ3GHhWFDO8Cl9L8nqbN+5150P+gEvQs
fJ5ndeZVMvsX03yr5WdXftO8zjfCE/7/jZ2niLGelranfq53isu8QqnAM9KyuFsy
uOW/eJGbe8i40nWXdRVPRRlenS2MdF+lvmKLRhBfUAtuCgPOIwm/kQjtDqRTJ5Nc
aKTtG1OjCv4F0xbQfq1LmBXxVdhOMZzHhpMRuNRd4vcM44cH8/Og7EYHDWxOIAaL
54im1W/aeTD/qCexY6xKMR0Rm5gGIGz7B+npnWpONnN5jnTXnMRwijLFfSQrgjvW
LKLv/373966MP1kSjfNdBx0yoSu4k5Cjoks0iPZaukK5NhIBqjByTBA2qSjZGmZt
e715TnR7vgh+towKKZ4du8F6/kk+PpwsqI6z9FSs8tgHlRJ8DNkBQqHZTrP5dfUl
bTbC81ol34QH3cLnHlmIGAOVLwV1ru/qEOedrKKfrDbxHoaQsS6s17RvKaxfNuyW
8qqopB5fIaSXM6mQnuIp03Y5OjFVCup0zvuZI6XwtqY6z25v7nBgLCGMFgw0tROw
j9DKdt8hUjOQMdaLJj1z9JIXj6rSOcXsB/glWM1FZHQ1MsJCqJ/EerFTdK8onuIN
gwjd7jtineBLI5X4I16G+zCXK47lJYVk21NCuOBlsOntlTAsfExudcJapU1nkE4q
UT12mxuZrWNuVKD6+GzJrERlNjOUsMPt10NhbQHKxB+JCcSi5Gp6xA0vQS7biE3B
a3nHgEw4vnHDT3WDQyrGS8IOtBD5pwFZZhSLJgaEmwzj6Rv4WVicqg6zKdDATeB/
kNvIk/tWQtS9vlrPRzRbZD8BLcz9DTn9LpRo9jgSjJyySyujt5vKdITAB7pN4SsO
w+eYfSqAIGJ5T3J8fyYiIJEiX+LkNb58RUZtkteuNABGziHsleyrLKaGPfY/5Ad+
6pJngYd81aPaMhJIl0PD3pKxYyWyZ/4JmYJcpSZKW8ky9ao4AyBvRe8XtK4YyUtl
wLkhLEkUmqQAaPrsaTV8G2iNGIyFztv04OYPNEcJuYM=
`protect END_PROTECTED
