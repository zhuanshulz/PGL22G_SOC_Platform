`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJP33/m1HgM6QhovEGi8RVuTfKlzEq2gZZC/IFb2qe9+9e7+HAgL6rcGcvEccM3T
Nksm8Hs8uxojaD5Mf8BKiVgi4YaQalQ63VbQolraZHmzO21puKSgfug3OwcnLzjc
YhGbuP7lntGJIWpQu9GVDtCubxPE9LsngJBJvXTcPbtnHt33Iu3iU08/f3LYf+eJ
LNOXHYCZLAvUPBq25d+Nrrm26Idz4ZCy4mLjdPBxu+eZMkv+JqTdSs7fbperVAKU
iUuCU8Nj5EjKBOM82ac4uf+/NW9FVwPx0E/H1ZD8uy6kzPaIHZsV/6eRKhdWBfIO
JnKfn+RDw63bCjE64Pil76L6jbbg6Bqp3wd1Uw6xor66PubVKew73DVJrBBN21IJ
4YYvdeXStj4h55n0w0KC9zfne4BpWFY+jtI39v6Zwkx5TGQ3q0Rt76Fu3vM3T7Km
V+Wk2IWQLAhzVZfTUybN57zun9IvPLZm0lAZpP5UUDBGRIiG+VyOWsWF17HIxVmF
G++Lq/yFg8nz6ipB8PDLOoVhHcqPbpWV7bSYO+gvoMCDjiVUmBXjnMpw+mrHFRMT
2VFZfoeSOx14n5Jxs5foqkwIvrZpxHXCHAC9xX+fXSPz9UV936WmAicLXaOvQDHE
DmojrbDXD+7Io7t1g0rNzOKRjp9xBYYjMD5AO17n9MAnf7V1Ceb2zO4IEKqamTE6
6tzbQ5nRvtEFWgRSV2KMhLfAIwn/UVPBP7OP6FhZjK7P/QbQt59Gebcs0e7OS2/m
esc1z5To78J1IxSsIccBB9F/5vAJ/6pS7xo9Aa4DIclP9ulX1526Kbx3gEWackWy
MKkx95A6KL3UiLqzT0YHHiN1jeIx5hBnCOnQlA3kaQ1OUuTmP+pu8oJG9+HMWFsq
8p6OZxZkqpLNqfSI893au72F9ZUBW9ekeupeA2ESsIoVI2QNBzlhS9h6kL8lDuFD
7uNGwXqNReiBNtl8nnvuV2DzVOnhhIDxSb3CVLWOMH/O9RQuelbmKkWKnRx2d1hD
RI+lNdM4ex7Vlsjg8c7+RsK7tADwCDX2mmhx1/M84M8LB0CwGq4MTV91vS9MRQky
tdAXay91ZBlCZ+iC8kHv/LLKcwWexl+kFyX16FOR/shD6vHRDsZk3jTYMtk/ZvfB
3Hb6yOS44XLd2hbrKnSDW2d0seV7NftyWjQxMWGajYQ=
`protect END_PROTECTED
