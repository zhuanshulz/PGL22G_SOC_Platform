`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YDw5W19JcPg929eQrbWsqdDQ4b4cU5j8d+TJb/Ssj1JXdm42tFqDtzlxbw88926s
/56QzEGkSJM+CiYPK5qnFVNF/hAxNVEYTrSyVmGcNmDs1XkJ8orbwXdNUVoFU0Xh
TuM/xotYqKOIhdBTXwoWa07qrh7qewvxzQhPU/QmjyOvIsGmjsX1a+IGLikJLCaY
ZyV9Kb1iER3iWqDsJPfsAFNqsQ9KNUQr32/r+YwL2fuqLKrJtxEnf5193Y1E4tEy
DBMrjzjO6w4HI+gWbCOIp9g7prY6oOivbHil5oHoB0650XKHc7x8qAicH8nulexK
flSt0NTcKW8D7iWhb9Xv3ySMWtPylPSxFNmcYzaxrfq+3drSnWY5AnJlDOpMC8na
HzcbFWFNkJdLgZ35B/GRmhC6QNup0UXjFDBLHx49zG62I90y1Yw6t2mmXXIiRqdN
jgjXtlgPuLKuiKUPSFGIUgJ5fCZq1XbxPEuxgRZgY3FTJxISTIiU7T+bshrhDv3+
hcQ3YQjMyXlzHYu5/EU64J3gzxklPE0Q4clDBOkPHM4RMy7U2FQbrWjVBNJ8KiDa
J12pNb4rcBprY4eG17VIpwV072ImwuP4l5t+VBWJy0IyiNCqqVbseR9nJvptODX2
Y2TK/zTZDXaUDOOTf7Z50DEnzAFcWPi4CjfEB/N+v8edlIsmT/hvdgdSH/6nycCW
1/RSLKVps2ojqeFB/TiP+k96CY6aPZcbuPqq4JMSc0L7QiHGCmFU7IsGlp8tAfYk
QIVR+Fo92HKk2ujz7PI0aIo0I47SpNEW+d1WQqsESOvRImHRjLPk5UhZpEh5t3AI
4DNkMWrPU9qWITaBgTRS3bKjkGXs86LIw+xzFvKZMxj8LyuscHGT53iTYhucC3BU
c7nBQCzFbNPLOysDrUIJF/k46YMSF/x8ZQibBhFl60O8RhfLfXLqzbwTsP48Mwt/
BW37FrHWDZUTeqnHnrk2yEDRF5YjJis9PMZ5U3gYXOnTvDceR080v04njifNgZim
pN133M/RExB7pwaNH+PXPGid4s/BVNYx1Sc+weCIXrQmGtSbXhy7rBn8rzbdGjBO
Z6CG+qE/RIpY3Mwq+APUksSXSBv9Ayv1V0rqt+3eUFkaywZiX0ZgZCjby99DL+R2
`protect END_PROTECTED
