`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgXnTIQ4j3gHEeBeIvE5f32886Zayit8nTl02TTCYFQNKT/QyHHcXM/0OFq3FN8r
cKeKXGNJjY/cHLgOd1+sEBPJLcRi4rWRRqC0tR86Q8Q2diyp5dcYjWtIlwGwPoaL
cBHV64R5eFuME06vWjA+aeLrsX55OyuCuTcYIHfm0b6jwQS/8VdYoeOxHtDSUuCk
ThcJZoYvPRwpXgdKWVqRWUGona3YZgXawVbf5G+RrwfoPpkxrh1YW4HfYCdtqeJa
i5tOsELnNPt4dW8qGLUMBM+1UURxClJfY4Xxr0HHX9D/yQFSL+HVsTL+IsNAb7pp
VtMHZfXQDSO7lmcKh/qq2WyCbh/UKMfjwo5vw+DmgoMNT6EM3INQ2ndpF4PimTEQ
qDUbhoFKAwQhbuFVUZ1C8GPhM4VKOIJeYRTGZJTtqa97kOQhWHVU3NWAknuT8L7q
ouLog/vVA/WIPOHDIkEY5NoojdyyiUGl5HfnuUwiw/bVRhLI0vQHsFJrNUq/qdT7
omOkPPchaTXmVy2n+8O14VUSZbcACUoikG13oS/raOYUoD8pO6dwX1XndbrNvIwS
HNVxxVdQTII07ouxBUUglaWRSdykHfVBWIeTejbwCj8O5v73vm5tJF+nHVILFub2
fbq1zQFMuP3Z+SFuTnzS0K4fdYyfmH6VaAdNNSuZXExBBLn5yVRFSxTScQ5xiQfr
kK0gxOX581UW+bbqofoOBQMvQbvrsrCcHPPpRAgTZkJBmmpRNGJz1Hs0fvPOvsF7
LZ6n08KYzl5WdRmYwSKUacw4s5/hxwUehc6/QO9by+PdRFRa0EdgkzugT/FX5yiK
fA9VYTGBwhIFuq6vkH++0PjLaKAcSkicfajoI6rr9ZtyRBQbViYpHohgiXrVGolX
PMaVodawlNcvi3+9QQ2y7k6h2jPlrPIiE/lANe+JhXP0zY3x67GszZJoCNFWDpBW
AqcHizSQXTSpoWwNrMpvkwkGE30encwxhvY6L0taMkhHXSwcZ3vYEDfM/EBQaCAM
KhzuDr99k8oyag/KJVlPSUeiPtePEmrHjgmzF/UJnRMnB1VQxg11hWh4aSbqZ7Nx
Rl28SHEww7WKg9vIo26Hc1UqZ8ukOTZzKC2SBAPHtTs2tFOYSucHNIlRChOuyvIC
Pg2UUHnIRfxgjMRS2PFq+Y9TvTrtO7Xe2bRj8MEKMJHcxLiZqkSMPHOGvOf66tMr
y06aD1xg46zQ+A2hnH0dm/WBFlHyWVG09DmWMR51BNIGZa/je2eexV/+LKvNJuBZ
7mtDoXGgoaF8UNk6Wu+TP2WubHr7m6MIag86Y6fUl49G9OiO5TX0tU+rrLtAg8LA
wsud343A2g+7s/qZd/KEdCU3eCoNptJWyuSFaH9XDAblUJQmASksOUVdCL8EZtaZ
C/P0SUF2PDSaLxAROikmMFXSjb+y5NSUZMGIKXHC8RoWtXHRvgAXiy6nFEOQp0Fh
64R8rvWiorFczcjIhNrk2iHJFN6XRxko5FMF3WYURGkJG/RNlCTwJRV6US0B505E
u30EBFOqhzNrIrYJjI4H/Ev1GtQrDVZCdGIY5yLRz/naQK0UJQ5ObwQStS36XV7J
NmmQXjOOpAnD30choovhTP4SF+wab0DAFEAq5RmVuyzQ881E9yf68jocWYsLxHuX
UEFWD9cAb2jVFtstmsWHk4utjwkY1bgTRlp0YrhSSpCiFSRjH/2Etxgj1vI+kyOu
JmtmjmgyiGNCCKXTt5iCE1Ki5Bs+A3aIQSw7xb1Rizscs1BVNtGFOCoWF+0O0+2n
LaGcQLSvEa+dZNsCMQyJ9oalVf78NLPzmR9OijayRSV1TmrqYrOKlqx1yZXZEC9i
y8SyWiNMObPR3OR6/yApHYPxkQL5cYeKv2Q4lUKZ2704iphpSKhZk59sqGVoNr2e
lMdSjfXaLc4wwoQcBuyh8H/ncLeKI5vMTv/ViFmFbPT4XBpXZvHhZ/e+0pHnd8eM
AnR2pxn765ik0QKJT8XCGw5vA1CgJTot0q/CLxmch1EFew/6xhiMhnSBhF9L5akj
UYhL2v2KK07bEh3n1dLZC4tv/81ImaWZNrvmO7Y4orkAulwio8ii95K7uxn19V7E
bSezer1gvdtAL+nYM7QmaloyxMWPJsLRdmbv3CHa01PlJ8aYoK895UPl3Xouevko
1cEmKFKx7X3MdWF+asH40FY83VzdRm9DXgHSPHlRIk5xT8x3gJzIti3I9//F635j
h6WC333sH9eBx/qyaTY7Aa7X4TIGUuUvEz+5v3m9aFWbXB2SClOPH1AUxebEOAyO
ELJdaiXlqBdoEPYAma7MI/kKD07iaSe1BEVL0KAxAKjtXhRO31TBb9pShS4t6P6q
pOXpyyKe6TVmwSjBXsGuHuvC+7yaYMHbIgmCAjhFz+dooiABTHpBHF0wiE27MXAM
vlbv65TVgFMfTY/XXG5Losz7tSUje7E6OSkX+yW0VSiTlD+kCqu0wsWoc2V93y0S
C6z84erZ8kcOIi/R2PaJ7qcwKikOm+I/6Ty9x+T83dD/pSXKrQsFBE2XZkDJfLdM
IITeMEy1roeVzbll+V2fpWG4dHSags203sLwNCB7QezPxNgWoZM74ymzDbIQPc1H
zDslQLmUQf5ajqNWjyvvP4v09Pe0/3inCv1+A9VNirA0fT8gRmQ9BDpeGRC3yYXE
QowR8OuzZrnSS4XAj8TcMCZGU6/DGBLoYU+F/xgnJ4ZyPv9MWHhPhiKwEE2nhi43
y2NWWz9gkH9PScXDVPxq6cI9LcebeGhRx9W4TNK+Ef0qiYRHmsUUcxBVqt5UAkgt
B5sUFVf4vTJTabYHOX0c8EiqR7Ux0oPF7t5gUncDjIILxnSN1B5amEvn8aBK6cGA
XVbEciu9B1kHo/zWYX9QWVj5X61uOlS4AjLsrTZ6DEKgDNWrbqPFRui8ueMwJf74
s5GiXaTztqm9yaSYoPuVmeiqtfDoO/OTvYZGQKlTbS2VgnnDHH2cmZpsvEXxirTq
9uBqHN0tuyVdTeTdNi/qye3fFyEL9WERHMaH0xkXm45j+tNY1PChWAFJrlt7uJMH
320i4WvfeYk+zwd+sAd9WiEnp9ufCoEwaDEbuJh2fWCUj0tdfKYuyGCcL/sG43rS
5STTLU3FtdU9bL4548jsRCIB+0/jeUIWIgAzVtLIZx6HoMIyb4I7g8kQHOPzhzF/
bHe6bOc/dQaG9LCblYyHUxYFL5K7uKyfV11k9IqXe27Puz9yQ6uorihTfuQ5kVFo
WLJMSkyYBm/aeTisnJVSWWqgcBOKDFJ7brGXbOszSBBDMHl1xWQnTXc9G2mih5EM
eMjjB+9R3WKYUvy1ajKRsld40njYfcNzIbOJd9ALfOTc4XfylT5Hkd259lgQqhME
usiq3Xno7BEbgXdVUNLU6usbw4Jo8FcFQz2/MAFAighl3A6qf3KfdRFKpvkfGXha
Y0MvF3D4j37pSMGSUwtwnKBRUiKBveLbnTDrXpe2d2IcbELv6dBWCoyCQk4ijS+s
ei5/ukHxpltXyBdzLDERRVBd0PVT+yFvaVU6UWYbKdPCcn/Iaiczu/U/iiNgzf/9
TCevV+grQ+Slo/M0EvwBiefDV4snDtsSZ3iwEB7qR/OuxzKlU/UT2JgWIJmA4np1
1Q2qQDgCdsk3IcouONHswl0fOnzX49Hz4i79u1+lrFvKT2QGUSws2hJBdrhd83rf
9xs+WW22rejQpJr3cEy79dVMszUwUlyuwV44tZhXmKWS/KQpJv8xFKTmSB3EcZS+
xjDvz/QLyKo8vIEZR/SY9gMc3g+mNkMjpFuoAC/LuKsfD18lHdLA5JM+BtVCutGq
wtrO5Oxv93/MveO7lTD/xzGKqb4YJbqCMXQbvWJiW3XRQh8lsuYuVKQz69wvIn2R
D6CiQKrqAP+U0Rg2yySgs0HEqABrAWucvPWlFNhoQMQkfI/EcGsVAN3db7vu49Bt
HfMnecPV9vK4dQxiulrVq3zsCHKVk1/g8TZ7/5uC4vb8l3QFhFwLqURTIpma6ykE
mPXyI4W4gPVU4K4NBFIdH6UyzCS+WC7KlPGVDIdPkpCqbbh5mTbjIrYitxHX8+T1
KFomcbcGxkC1QO2QkKw+9qUvZ1tlYiwldVJGFrghOlj6mBajjk5rSSFMbd6tcjHx
Cs+7ZRaGWOFGdxBNN2DOm5dpJm7eitrTjves73uf5I0D6crO44j3/5EKKMq6thhi
jNUN1H2E0h35wFX8ddXfeHj4c5miaYGP+B7UBhJsY/eHexS4fmNyhMuIWtb153fV
Hvcdt/nMN32BEZJed/7hYZd1QjUkxlOYIl9v2HaZSDxLBq85SSDxQufTgc4ihFnk
eW8wZ3cQ7i3OoSXoUfKqKtsTM2YWGUslJkw/nJKNZQzXcMzRdmFUncYuT8RkZz2p
R84ZpAnEvjAK0uET2jICWYAMb834BXWqr5M+26Hfej9Z/j/UOXj6iisICrNlwglh
tDeiLdLorvA+41dCnsQeSAGS7nRfiEA9nfKzcDVCeILgB4iTn8xPohVKjiMl3cE0
N3vJ9lILSCmH5m5l1bIX48ua6iNnMlH88eKniVarlf5SQ4sKAW4nIvTIUNA2vlGW
Dj3/W/tEBV6kMiffJiyj2B0jmlEmFKo1wqNRjWThei6XRaRmUxBwGca6vzMADhOQ
c61mi/ddnI/JCuoLtHiZbhlu073EJY4vuJgN/eWzS1l8B4Ycqvw2PzCUSZDXBuoQ
eA+Smi0eEmUDht444QuK9V01q8jY4f/OPukIyahk4B+bfxk4q3tK4Hk7tl65Wi/V
C/KPA9Jwc02f7cpLt2hMdeOiQJQ1sjC//sr6D87mTZ50MkYETrH7ZVOjzUlG3tK1
4svhdN+UjAyFUpT5mnCuNWZ/P/sZh0SL+FQEVR1beARehe/g0UK/8NNUFUL+qXyq
JZGHJXqwWa0NSGBc5Z3QyavxF139j5LBFMomcI7LFY1IYXXUH5i34pC3ykY0mNGZ
vFZKcqE4cmi9MFQHKuGyxt0OmrBlJEM0bZhRed3vfhe62p/mjW/qcS/HKY+qfbc3
MrlnLozd5NwBayt92M5b2/UwOaUyjxLuYHcSgLuVDkJ2MHoAt4PbqYgt67sD91rK
JbRfjEoqFP2Ro3jz7eRvO8Kg5SQeIP5TToWaNc7M0XJm2PTTXwqaC1NR6+nPdX80
IPtfsIC46s6/IWCMZXMXhBVIHVAAzjTfuoSn+Rhcoaa4zfvmcHPzzgiXULBpxQ0m
dhWu60d9yb/qkb8I3Eum4n+0l4bWnuFdQ5J7FcDlrqFv5kLFwtIX7zwWjtR8vGKB
2Tp1/QWx3mjByC6OTOE+Jqy6xj5EPnVym8CI/sGsOangi8p0wPObx87o1TvOrH3J
LA81olYdWmTbvSuukDZk530klwzrN1r7zlAApYGW3Hje2MZGZqoE5EoplCvV6/+k
OeAZjcxGXgBQkRoJRec15PwN3rvWT5zQ2tnmTpugm0nvX/TS5pMk5stn+2Gjgks5
Cn9gJMubKiBD/GHk0N4NccuMQfZ0jhDV15hHPe1CRAWUf6QBkkz4jl6LEZRupxdC
OUrQlbpaRwWfrtHpFOUFWS1jPFGAtL84meda2Tc/8unQ8GtGyGrq+UCkPRLlxVIB
HHfyb0QjqmKkg/SM/tRP8X5p0o0b5Uz/5mygn4NFDteG1yqx+hK+aj54i6VkuEyF
W4dd0wawxVseB1UX0OlptuTbbpG9+Tj0q4Qd+ebikkK7B5j7+4yiwzNXCooM/nZk
p0wtoj18WlRaZYmebdw9h8CsywkK0K7glv7jap+8ufrjhkQqPOY+lO5asrp27SBa
liNN6c2eREDkVym/eMNlp5GHsvebTwJ5jp7G/MWRro4MDUhYVf7g1VTE+nzaZKDr
UTfCJyd/EueUGmNmiN6Ttp5gJf1TcGm13Dl92Cqm7q50Ywud2FOb0g+MCzSTh8aW
Hu4obFCP74kUI0y05aV0OQSSehkJj4IBjHXGrWFjlbwx/TRITdxmot1uQ3Y8Z13j
+WJT0x1hF227L0IlLKWbirOG/Rl1J6eWid1nBndafBKj/fNtip0+vloWHBFtChyJ
bnUN7kQtWFON+ahuc9GuPdu1D2tg2ebNJGCVOEHxLxC7zqjk6CiFGnKnCNw0X6qR
KOUn1ac/+oCa5f7DAYd/ujTCuzBsnUPvwWAcPmKj8VYKZWSlGQ9iXlC4b4Hmabgl
JG6JAHzWHck3LSB+T5SB5xOX9LcFBezfzQUJN7Sa5EWgJpsDng7wPUHm1DNWigTQ
WY08Z4xFfYEOlpwAj0RPKmDfejVeeoQU2z6Uzw5TBcaIknDER6bg6xqfiUUCgLAI
/yZwJQ6+lf0yN+oxKWmfArBnenSQoPMJqjuKEYLYT1C9aAs8tsa8OxUhRaHqF0/8
iI0nGrq4athWAxK2UNzOpg3NZkys+gZdp34Nk0QgdKxF2yWPGxJ0nDRHvZwsJ4Xt
aC5up8AgGYqYVk5h8Mw/CWtxCXgkcDsbBTc5MXO62lsegGBYI9q+EKBVY7BDNJ+l
oG0vH8f80/GOHOzHGhTXh+fWuJ/oa3i31oJaURbA4iLgR1nxRTK177xWKMU8IQzz
HWoQ+exNy6AdtAikPs+h/c/yp1QYN4ZmLqVyz6vV7y/RVi+y6uWhAdrvRt0rhCou
zwWAj1E5A4OwQUeoNwDF1hLaWe2lYeNUOJiuzEyPl+nv+C35MgRWeXNOjMgbT0ur
lG0hzrohO8E/5t040BP0MaKgIiNEbiOkDFwUcqC7iICKXxXDUycIcYOqa9ugKmM/
96giBRsk2VrY3DYfl46gC7gNjjYzkxTeF8ZHSmEXJm4xwe+dR/8+XhuD7wjg6MHF
FY0/ptAFMX2ZNt3o8ZDb15onJZPAI+TTr9sBWswZrzV/VbsGOuq7OVHh3h3Q6mHr
xOb1ngefp8zDPMiK49EaZetR1Up9M1FcKZ5j6jfRWSnEJyW+w31QsrRur73/ueRk
rnudmW/x0HGNcphdVIZOYwrWRHp7yLLIirv22R9WVJO4HQgnhbx9wcfX8QAvynqM
RXhtmu8rHhyR+N7hYDUAIp/2d1iXCgz7sX+tE2hvn0kvpqK/nlhQykSPe26uqFxd
SIs/gUAJSqzRake51mzCTJMeEk3rnpvQXU8Z0CUwyy6HKdvzpDzda9jaISDMWNHT
1ZTD5xcrNs6DlkPQbpJn2ojgbjcNovU6wdkI/nipxgqQTCtj4FCC/e36vEZH1mg2
CVOHuTk00CqknxvCf2+a6qQiSjpj1iRCTmZN7pnCjQ6vWvlzQjqyXbtqfpGgNnWU
EPSRtaiauGuF+JvBlcyzAGgHhVsSluG7b26Quj5svmWyIXFuWIvXkMBMl18OMQgY
+MerDpF5AID9ddHuqoMtKOiXW82+kdBLkf7R516618p4R68LnyHGmsl79VU7p0T+
xP9MlVb7pIjZSOYbb4GhaVvnlEqxOJXHDpUgg8DrnJ1aLx1jMn76q2UBEl09ioVm
o+nlQz4DxM16AHgUOkYWC7DcUCnPHInKWku5ycJKmpxBzxHbh3XDTf5NsuYZIwh2
GlLZC9SvgPCkG4TWsh8vcoicsf+Akm0kA0oSZ0zsx/8Eber5n8kbzYgCRyOSXTcw
aRmBHvBIz88d0CeC6NUi+wL9KYVAwx1zDraRDYz5aJSaLD14cYebhzK9WLOBRfuV
oRqoT+YRJWmqJAuYSPn6OW4afwdIn5ffHN42oQTUtiElmAjVwL4fucqqK+HT0My2
aUJlhE0JuW4hJ7qSe6F+Ip9vAliMaLo6MgWRWZdVssWSJJsJxkynCVzPiuojf+qQ
u9J9qcu0EY7Vgo0ooQQ4+cRiG5PkJex7+I6uf6sIlxSqN00gVUGbgWdKwqaXIkxl
5XOZOTX6INhQdn52GDP7vXkijqY/xHKdIestvoyBjsL0Ep580Uo8mKgTbVhCf3DO
7uczTrJMobxHE/9hYHPy7BRbpnl1wro6+nbn/z8Qpb72Tae3LQ4Kwucz0RUR5Njr
juD0eqOrQpriXsuU0soMew7iBhR9OJtbCK2FCiZRxHj3ezSFWuxtn4SGSFwQ3I2h
Bs8HCD/RoojTsjzXBPl5PwTbNKLAFwuWv9PW1LfPKBE866Bw6KBWrGLmDptdZhiq
KjywJjGRcX/isoLGnDzNCN/4ieZIug1v4zMvzSKrurFfdHEr12x5AJNSOzaD3hHm
7fP7HSNm79/ylCebwgG57hrh3zg2S3v76Q8jSxEoFH0sYaTojo4sK2ffODyhmXvb
MsSbMhBQ0X58uTbzpAOmT2NL27cxBxjvC/57TrltbX29jVnrp5AtkVcYRzdbBlm5
HJq6NooQuhufvepUMBbV2RnujUGueaVuTh4XH1v4IZuLX7tzfv1qRneWJJ5BMqjM
f716tyv+nSZHK6sp9IB8pGwgYbxqYf7DADihb925E/tuTYvxa3FmnJKoXSMONhKl
75WcTxEWKwBzQPqG61WqBh94+2MUaQp7m6p82XwOjRHjQS+eGlX1GbcQiiMYrMjk
gTURfFO5UFaD9LyruE70N1kWF9ToJXBcx66knL2HAfuDyGg0toogSFqcHysWRdP0
r3JXI0ds6eKqYeMkIHPzxLZHsUapc94Po0lT9D/wfEi8WVhwN3LqUCNV3sY7wK6w
KdXLEh28uuyYouz9yXuaqdkBhU9YcKC9F52w9KGR7+A+0v8ksD9DphacBi1gcDM3
Shbjtea6GmyPwNekVi/8lxdG2k0X+aCpoqYAYY67RHGFxa6aH8xNjpFsqD7oeVe4
DPVa1zgY0c5TuKnZxO6GG2RU7/nMBOA8syQu2LynerLPpzo+5kioGr4gzblT9fPM
KfuArx3y15OItbRJnPl0NLsKrJyzWmYhmLXOnfFXirNzbWkOeBQAQjkE7lJhfaU1
ncRP9NHGMce8lR4xWZ+dVQR1tL8WnIoD6ATFcbUgGmUrZY3IN4YvSPJ2Lb4gcIk3
P0s158iRxq/ug6fqyMkpSiW0d/lRTPx2MurHiiAsxopvWRDekaBSWKH01Azf43Iw
jqVpc0kH66jEY207FzcLsu+dmN/dvkrDokcvmfUAfb5McnDCsjuh2jC8hPfMso5Z
7yxdyRXWfRVEkp3kie6s6PrY2Y9TR+ymonAksBM+57CPJ4nC4dtr2QhN+Ig/sVrs
qwDPeqzE1AGdHyggoLQbBnu6giDV4zAnA4VPygf5KPqWczwqRA6CgO517gvLV1OT
mpEfIiIPxVp9z/alx9aOqz6ChZexsoj6wKb4AwP+8WblC6RqlFMzDkdbnqp7WlwQ
+/nL/quJO2A8ZsCdlqK+uyAyX/TPDkDBxrJ14AhrTPDSAcBUvLyut3cb0F6mWUSk
9GLGr4xBIpAAEXQS1dvJSo43AQtkfJXAZ2QCc/LAR77o24E4qd1k/XlXrZHn0Imc
x5Xh3GAiQv+RbTGuQXssXv+agX3RJIO3BWX3mseVfH9vBIyJpytMg09/NwfGxcmY
yjNXY6V924sO8yXw8HOGFzFuP5gmE6NSIq0gg7TGYHMhC1o9hmMxP7h0yAnum3xD
LMbVTOqmVtwgEaqgzF9U0M/YqJDO2kyhIOr9No+Vxx1Z9srPwj4QUNvriHngRTWP
FHOvCphjQs+ZPA3WlD4lB5a0MeXNJrS16pTJeCqk1wSFaAPNkcpvlHg09hlnjnmF
6sFg8ipY/7gUFKp/3o5Qk3eUDojgyj/k/bofHWu80v6IsaVnoj6Yr0/bCURYbrdV
2w/sbFtBrIAJn0CCr0KnEnoj/LV5UtfFU5IwNf4lPVQoJrw1muubd+LfgTKGlos2
2PcMLnziA9yol5E6khTFK3PbQrbXD0kJgtlMbI8dqqQynatDS9vcwlkGEPbJg6CW
RgUxTO+ILsddMW/5L8QRx5jbXPMCbXnU5NFaNRQ/8Ek8e5OjojQ/Gw3zpnQfrY2I
NVgIm6haEh0uJLa/hB6QP3Kuy2uJRZd9FeeLsHkQxso53NJW02UCfamhmz/oQS/O
4m6kOw4jLtQ6L3iJkTqNMB/EQTudLHUHNLnZItpOgC1jLfHgzhy7LJEVqqrrDUDy
k6gYQvN5/Wg12xN4pL6uCsMXzxDQQd/NfJB+iRP93gw5tLAHYS/vFpSd7Uo2+ifN
QtkF68/tLB9eI0pSa9YTokpgyf/pKfEJtzN/j6hC8VqlpewpjJZ4o/MJ9RaOXvhN
uiRaAFhOAS6jsCtJefras4XPJkvqTw3c5qd4cftpRlMLWsspHsk7uHH61u8CFDs1
5Hy/bl9hvf2BbldAs7BmKgQtjoh8+BWZSQA27bazSnqk0r1C1InJEdAm/ZQWUazU
6GTCFDL71qYSHv3FJHqiyyrE0fEXV5cijYf8TmEe4xmHMIk/dIxBa0kxMfBQHlz4
tjz/1o9oNbQG4echvVqzOO4AHFh3fMQ7iAXiPw8RAlvOxWV0+up8ixfAEwxbR7TL
Zu1Dix0kSCzPBVUphhlg/zrj+ym6xVg7BRBPFsupLSiKkGWF1rx0QHH2HCWntJSs
Gd2LogRYb5vpGFJIJ1zfuucbVBXYd67W9E4higGPhMFMM6ngAgPA3tfNb6cPXtcY
7vqljvvePCtghR6mjzwiwBCLD9p2SBECp7tDAQIB/nqcFW7x+z3svgx+GLg1w9au
TbWZhjfdRVIB54tpKQwbYg3SfRHmlNr7p41ezMNN+OyBHst+cCfAwpzu37rNjYO9
QYJRyJsUT1uQys8h9x/IboGDeLQwL2keXRMTb++RksVSTYer1+59wD3adrZ5MFpr
XsPQE97GMvdMKKwfoNdc39N+twszLTE9GtwlaPza1Qvws19NCJoD6fZ8Wy1H+R+F
z8UteSb6hbLKtTD2l95cHbPlz2xdfhcofsitiXqCwYlb71WcRX454b2dR9lbwVic
g7DKWsFWokF488iccGKciJYSr+rYrTR2zOIHOFRwmGk9w1x/kpgJorb8yvcS7G0e
Om2yloQKWsiLLpYitvxMqEF4ZuBbcvDhuxdCKGytataQj0Fh63/8EQ78lrCiUW13
KV2oA+HmILkqDRcD3ji755foTfDcZ789e49HpG3hc16kp8owz222yRcbERgHY58d
Hx4Vp6cTduhpZci+0QNdxj6/nXKddiXk+u+TtjtUexPKf3Q4DA5Z93Hlys3lWTwn
1OJnT7FQVYqU9FpfAUqEQM7Y9zaQLd+KSYEXur/Wu1n1t/ELiGfm2sJYzaICLzzl
iDjMt61aG1hUsculj6dDgA7HESbE/MOd4gnmNVt/r/XDyRn5al+X2Pjtwyqp2xUq
9PgZZNMO4dZvbQT6ymuRU2UoiQGCuH8qIc7B1s0LMeoFCKBZ/xq9Hc8L8JS502K+
ksvthwDCQCFZ/xdV6QOL0yWbgxyLveze9Iityk1rgHDUDM+2bgvBjIVVNpHIrNmA
727zUk78H1j74MPuiep+pM5ktmn/bfUGrHhFscVLXopeFxgFBrNirk+Fqr/XWtaD
iSUEdOkMWDgJZLywgSeZA9S0WGD4cMsgoV4LJ//7mV7OMR+Xt6NRPW0AmNXXtyVk
JBixoh+EY7ktmGePoT1+FltprXYLrVNRH3X2flDK2PNGrUMGzGWFCGvO8MeIx0Ec
qICyfJgY+yd6yAklUNBgBjKUx+Cb9/D8qDHcJyTNTd7YH59zCejX7Tn27page68m
YTuTkLnt3VAjWk+LVMiJ/5F/xmPekYaSW/RpuilTpd+mflMOLZjPONJrvO+qU8yc
siHK05MkZoBuv1wPEv+J4G5MKp9C7OELp1d2FZlE3J8Jw/1J5n/KtY6LtJuLaI09
36r4gjTeiumLR2Ioi8xqqSBS4d0AUkV0IE9I33NSu95xoucCH8smsjAoh2fw1Oxy
OzlEa1Ae4DIhFeR2uO2+XNHi/+BNHm1xgUhDKF//qbtyffy3RzJhO5Q4NxFcrrJm
NOY7y476lphBIcJdpL9Im8zd6GQOqEjZBAs0HF5bEbJ5TmhHGScGrD3WfFkFRsRI
WGPKmADXG3E5dmx4EQSCWXQVwb78DzMW7Z/XMCbjEofqsLZOti4YpYVPGHYRWUcD
qxYsp+c6VqQ4x3tFcX+ZGlkUQJEGLu4S3qoPaz5mMUzvsNFrL1CU02VCL1Jc7YxK
CtSciped1YMg9ujU3psWDeTHHa/SW9/ye3Ju0K+t38vFPppMzY5cD39gaBwSJG7U
07oxPAOWW2uaAPXn3yW8fB7L4MDsVXDEnYP4LPpaXouqJ1A+SOGCWp7vszBMLu+B
aXkiQs96N0K8c0VamE5bHpiAgDaY3nGjL5l2gQpZ3vMfLEqbVbU1zMqS8BhC4Lz8
RCanMuqrUgPsOyfGM0z9npaFoV/xCOJOQQSHmGXqT5uTS/ZyHt82CDG0lmKV+KqY
8k1/goJDpFY3VbkYhqIC3wx1yifysR4kLDaQufYFXMpJOLgnYA61Qsiol9EdB4v9
w6fuY2uhaU0M+PwbICGb0pRl87IbAUgPRH9xojNl7e1M3wlN93H9O12wjWT4pKzY
YntdePdApzE1ZBPatvG11qXMJawSqxgm6fXcyuozQ5eRU3wbcB4N8lB/5kbrpVTk
4di5il3Hw5vrfbsBeeGOhP/nVOSh/WP3WZtZ62g6U2fdWJ7dpC5FJxGN/ABvfr7y
JUlfow3ErQ2HDTFRiMTdTaOLBIE/PLZAWNZMFN8QcZUc7DjXzSVZxBLBd9VAfQ1d
K68yWqix/dF9shO6xG5PYqYgFrtoiXsZ5mx9sF77u1BYIwYfK/Tngnqmtr9tZUc4
6kBy8ycHyqEbZVlG4uo/rUpvXzI3xhCTTLJgBQ3SP2r+BUwSWdaevwFXojtau6hD
JzJOr0cU79Ls6EAzVB5FECwG92YC4EBKy95gPyI/6kGM743ew/7812kMdoMOgEiq
thQtCOYvazuWKkzpNR4tZBqCFtaPnIJqPkrqbF6A11OOXcLxm9KP9X69Da5IxTot
z6z4VrvI5eN1JRMzT02T/GUO4K1QqLgxRpFsb/HE6G++qS+FAX+eWyl6/ly5pwLp
Ilc7W8TnFa5+izSbLT0eDI/g748sciBB9VYlfzgukH97WxTqiOypNVpBJJ6S1m4x
PdzC5nM78YR26+i283tKsq5BSMZ+z6fN7DPNtrazRe15Qh/+jp1rvU6zeO+pt61j
17Fr7vb5SLGNmbLIsDlz2KkhcD8FfnAszogh7Hbw4mCEVSalw1IEJ5H69je2NPOq
Jltn3xxCw1Ul1cpGUV5z0hB2HvNxAUbZJVL8k59Q1pWgxTzC583VSUkKlRUbfp4Z
HXgIoRi+p7pVq7PsLADhDFu2dqJS96voKZJXmtLs6H0IBC6bAdwRJ+GHDIAgIRI1
SOJjeUq3gA4fBT9/b/QkDZ/k45OJd1Y1fdaswZq+lUQehQjJiLsTs7yJTFJlLTwm
smghXmdhggFwj2SvHxAQZ2Vkx1BZVyKQ8JL7yMe46wM8LiLvmmiK890wE1p1VAyX
B9UJK3LC46w7dEfzZLMXy6t34ht3sPGwocVrTLZZa2BU8H93rDgJoMiwRqJ/KbWn
De4cjUve34+XH0+fvZR+CjXWVWpLQZxpSdDPzAhQXwZIHZj+f3kvEYWdIUfOmUSL
I/gJvOtCP6se9+i9oqlB8URHiXQWmwOfqXBRtMyH3DIfwZ8y6uhKWLWSONdDku+1
7u6xOPswN+uVAO+8rVzCVwpIq8Ip1hhk4N9QCwcAXjXz5oW0PHvqm13Tv6NpcYax
FwrEYOGUyLDFuYwqIr+UpKnf9f35EfzGiJNPoNzch0n2LhZtdtsGmIC+zzVMTUhk
CcSPFBrlhOFPwq6yjQXomSmf5VAVkJtBVm+r9qNEnz83o48wZn2OghAfIbF89y2N
QtHvmW/uGoePW6MQ3TLp+BOqSpFxup2Qx3KQNEYcJ34SuhmEq71APskOEWx4NOJz
lB/o12mLMb6iAB40ihtME8BFoDSoBDo6kdRYftji8L8Y8jEPCvNpuf9OlaqRTqks
eY2JWiOr0ym/a0Cimt5kVDeHuBjyCn5UpiN09iI61NQzC3OlnV4h96rukEgZUXj/
tdjYN9QdaaXGra0KS9ieR53AxWl3jCvT3syxPX0IleHsT+TRXZtCOm/3oV6h86AR
8Xt0xnkI/u3efF/1hFkdRZBrzn6KsHHNBTSSgllKZf5Z98E60Cw9KyeeMsnXAqOp
1bzyf8/GXc2wkZWhoX6DDJgu0DoTISDuE/2i6woGobypIoObecEo8RRO80e0o/EP
n7DHuaL53eKee0YI1Ezfpyd3nHHlIsZEH4Znf8ySs5PC8S8lk3oq4RibrdCMwq18
1/O5faMOHDLq+bsAxjJ1WtB9nyHl+VTl5iefSSnBqIcF9quR5L1P5JtYIk8sq8kv
yojoI87Q/snjiaC5zsrZGiVxxesj0u7vYIzHW6gBSCal4ojieVZUG8O8FJN7CdI8
/zjTAWHOv3rEjUUMtGd99nyI848CBDsiujq3HVJ91TZjSGKvdCPlNdx4Ae47xbea
Bbo1dgqlwTvf8TBfar+mNHYFyylwR5bgIkHxAtL++SWI6D36Hz2xUi5hRytNlsfv
LeFpluCCGdrGkZphT8HX+Ep9UwtMCsjueLREU02RkvYJnr7OdMVfkcF1hJ3cOaGR
YoGhN9BhgRk5HUPRqDq9CADM6hh3hLZvMm3L0FJz5QwlgmgtQMI5+I+VacrXsGhE
UWJrIyr4xUV5lV9DOx3Uwfk7cdtPEDCfE0ykdD8RddLhI6KM8IrOzqkyxlUwNW49
k7a4fdAa1dRpIwc0srKPCg9/tC6vIe52+D9Vnpgi8yj838R87iVKZzZYdtr3RNc8
9w+Fne06KhLKTcU4lPcKjIkChuErCB876RgCHJ1uljZVeHBtyrt8P/iBr/pEYoUz
lydeN9usJq5SLFr9CH7Ncbjfcq/GVrOb5D5IW+khX+HFCirstIxs4DNljDeDF6uD
2PK2VPleDWG0il5t5eEcVE2YAh9vqapUWGN6PZVR42CbQs6NG7qs80Am26zU9Tcp
wtLENFifX05fcC2IbvHjb2VK480l/GUtBRhLGAGr6y2Fte7EiTnLlmhAku9Z3lFF
vDnriPcvC+QuoS13uuBwPKBE2hpgA4UydGHhopH3UvbzLN/QVtqdBWoo/kaeN/L5
XNyLQulpAamhFguafanX6K2Ra1VbQnKbmIKy9jiIUazYQ7RnpvfJxDYJU5Ygf/qb
OP9mqkTrFsthMC0OqCNkqqgoA0/xRmzAAP6XP25SZ9kqnhn/9Le3Q1Kd9dII6Yy8
Py3i1qL2RqcOz2xe+T2V0cdju3emTlkrv/ag5qgvvCN+cYBv5qQ+iZZSTAx4tsA9
RjI/QYTsluBhZRc+ywVCf/NOaBppOw/ACF37dSKlpVw1lQnJNa1UWxnIwmESVSfS
TJ64z925vIgpFeSk5+bUxMltAeVpj28XEbGbwuqHcmzu3s6ZPIv2H8L3w9yRVoeA
Eihuhk2bjYVaG9L8XpwFZDCnK7TWQG9DgWqVCdUP55pLKb+DCVpONnjNwtQ4VhgE
DMVBucvWboemZq90O0toFHzFO15nhC0I6Z4pM+oFCWDJISecaMLxY9OKZlXzI1uH
kvUEfKmY8jLkPSuzxJ7z/oKzZVwI93RAL6FNxDe2m6A3duK5LS58KITXODejs8sd
sA395b31ZWJ3YMFc6iEhokifgHrOCA/j9+C8tA4nSHdaZJ8dCoSv3RpJ2nROZWsP
GxJB1gjZExMBSa+C5g38GKBdvubDmVme46/he8XnMas95B2eFFadIUf6pcXnt99B
7EJfAVMUiTJhTGMPF1vE5xPcznlkdhZ4shaEhAgD9dWwRre/eMIec/F0L5Ul961F
SB4HnIb+fmADMjBRyepL3xi+bAYktX+YMHGBZKp4d807j1wk9MpVka15a1YOV+Zr
Z9pu8cvZ2fNUyNrSPHLIfbI7xDyfHwwZCV5tiNtBT3qawI1AU9NKZTfNqIToJPft
A377PbUkDRt9JsSH/TTwQvP/tIq3XFsYdFDqlWQ3MxPdJVQiPoCEYO+Wk64MsZio
pPFxFQlBDSjGPBApq2A1FBNpVcKBALtmVd3yri9lKSrmGWVYkIdwjxcIhJegGGnW
tqTxg0D38/8jlnoo3F2fLHIcmgtf44QBN2tLJixyuw4Y9M7KfEu0NyJ9vRtNAfHN
KjKcvIZDJ0iRTIoOBtQNo0ZuCvGEu8MmsheBX4/fRq3dE4s4LLS9rPJaq6vtYO4L
adiLIvBKi2H/IXVwoX06sTex8OXz8UdSOBu38u36KtsLwZGdPBvQvtlIeiHV9xkx
7s82kvBd7EoNegUOjZ8GlWKtvqdzEFyvhaGPJksdwZH68TbGiagfKCYDL5KiScAa
NBLqKBUnQ5TLNZRa5n7aHTxuw6AXebQQKc+fqfMb4B89IS2x3PVjoJARIhbYaCuh
fMG0QO3YMP+UkQ7BNbTX6GSHWYj8XqMtnEeMsxrYlZELtKix4W5qBHX006xTbS4u
TjVwtGlzeUHjYj5RlQm3eZ0KdO79vv6zTV/DM6ievT/DgA+woRgI8CsIoEPhAxbv
5VJSsFBvCzNK7IwqIx6mGa+9Cs22ZUWFclDajH4gT5TYRJJkl1tK7EomlATX6C+Y
jgqb1xH3DpYrNILVd/oL64ZO2tN4erVB2tNZMpsDynzWQqaKid1zC/o2SZWW3BWT
NqFa7nv2usI2wFTLW8C63GAfU9Ic/kSmWFMeTUwoIh4OWaIrKIGn9OUvzs16eOto
f4fcaH/VblP3ciNmQ9sVAsJ7fSuQeaPxcUbKbo/flrMbMmlcJaRD/2akc3ZaDd38
BPLAMXXhSTfvF0JLrodBZUF6JiGEqXRHMyRk3OzCnmT0z2dmpfTyhbrcUJIjbotr
JpEossxRDNVGrdXu+TQ9LqMB71h4lgx9+n7N7QWriPD6AXgf3YdGQMKu/YjNx5i4
qX20HU2SkUIuMtEYuAn4YoabSD9yf0Bgp9X4NIHd7rqlhLgc/aKbaZnmgH4x5FTI
DkK+A8eygwfRU3eCvz2uM+D97xox2nQbCQckDdmA0PUkJWc2tDMeIJXk7hudvF1o
YB9zJrmaEIFhyfz2ncEBh/NeASxRtyMg8RGwUPkJRe1sm3MlkKx6NmMZjSV+qQKB
zpXLCdXNeru85dJzgwtXVEQvYZrhA34YnYYA8eNkcW1AvpLmF/j5YcoZSVlxWav9
nusWUiZ0Her4e69OFiul+j9Tlx5HTdX4afVkrTOsGLjXQSgeHLBi5SHg4/QuDNU2
gTt3TXHaejxeK7EUr0djhBJD5Uhw3We3iVqt5fl5LiAX+1PqpOZHaI+9pu5JQCCZ
0Qxw1ZpNjWI67z2NmEaXHTQ8g+zTE2GbKtVJvA5c/AObUxuIy/Bjc0kjxmTugJ9d
aXtTyR0LiVhk6chqZrwT2dNshBJB2KlFgAytIqka09KW7hqTElQ3mgp200TuUGIj
TlAhG6bx+BdZKQ/k/GfANb1pM5Wkq0MNJSkjdMAIfM4q+pY58OlOPGHNajysV7PG
o2pzjTpQaBuRWu7qTe36NO7JrE8RxkUbeE7YTbTYnOiE6iFC2BMsiXqhWVBin43q
Z9DPbIFNmv2R+v6iGjQIr7ks/OTs2F/HW8htsm3mP4r5ynD0zMZc8SG8KT+SDgX5
y0DWAH8L96bGnHDppeZOPb1Ulg7LFNOERa65qrAHuM4MxOjHSOevU4VPHsT8aqVX
PghHM6SZ1kQ0UNdUEK3bIv+NVD4NSirKLBTNABYK5fiJKBP59yYfBpeMDwJOnAi5
L+zA4PJxZzlRl1U5sknD3Oc3LZnHIYwC2xz8hA3hmg+52ltTr2NvO5N026LXs0zj
0MpgKFPVDHIfHSCzkcV8xRdjEy42Wgv6UwbMhe4vJUUKHE81hZTeOtMlO6YMAcV/
xWJ4Pk965+SV/hliVt3DTeVxXUBAwMoz9voBXKF+hTOyhjuBmaefBAL9uWtfJmIE
29MACLV5yvvBEg6RZ1MPhVzFHpdUJAoYfrlS+otuOx5EhYDaqkIw9Ti6RM0j2nYj
zhYN3R6DDtiwMp1NLPEMiMCnNZKfeRdR3XQaRBl8oiO7clT2an4hATDpH0Bowc4A
ekSt79MLjBZsO7KSJMrnTV1YbqrMxLJ0vIdQOhuOgHmnPUzzr3meEe9BjRiZmw/8
OnuQr35LQJ+rzvCPlfIFHdK8P5WztKY4qFSQLVeoejvHTbRqDIG11HYyqrs5Ywwt
jv6wtMZPW4F5TKDDQ3lrM978/0ldxNhxs5BfS2MoDT8SgGaFu/w7RpJvtC0BU72x
hw8ck0xu+ddkFHT25IWIzk0yuI1xssdm/7FRCYrAAveoN5p+9r82F7IOXXK+Ap1V
uCiAzuaRqLv7S8mRTo8a0xTdRU1un07Cw1GYNxUmjvGxutCBzx2pbFElVx/H6Yds
C6LL4rIZkM96mGSvAadz4Nv/+MLb9j9FlKmF66b7NaVk1VBdPuRS2WlIWVTbghch
fF5hTMfP8aqU+3+C2OOFmiwcjtaXRA971LefVNIwfueOBXUKm0ObVvK62N/r662f
uC2F2kd5AYw23t2SGhFhRnJ6zJXDp0QMOLZ5Xjuv2cN0j7MFuC7+DPedo05wGwiW
iAe8976Oen19QQmcqdQMYZqGrnowCn3h8Es/Gkwe7T5yg7WXQAkiwe9zSKgCyM2+
Qw9xotLSl9WPjP4Iul7l1YKkHtoOkhyg0iP0LRnFvX7P8tGd7rNhsuJWtS0F5Wz3
HFWpIo833fCwBS9JvK7Hwb3+xITpvWO3nEcX6PasN3nE4nZbK91u5q5/zYsUF1Gt
0OHuP+AyzQtL4fE38f7YahUX1cd2NNLnRVvcqueGOdCit55CU1wOfh1rW3FT/sdS
eQZTN13gXRyE2IE71SyRazeCDC5HIbibOJtG1Ba8qVgPeh2DrLlYuSx/rAhIcipX
VyPLpWKXtPO8OA/rPdicKCRV0mFjrHuJU+/TVeoODClSlQnqr1r0DG5w2BScDKKs
Xmj6e/EQ9uV9XNvsu8wG6d8kSc8dFpvucm6cAOZU8hxaRDwb+gqKtTOkwQ5zxwuV
ZMTQtCYInD2cRDsGHw9kTtoGX61jmWppVj8vP/lpV8lmwTb0N9D+8tg+trT9z+Ak
btvl95o+IKP1MlUyxTdMqqC2XYefg9VMSUyt2trTeJWBuDDoDs13k/8P/CLaMpbq
UtqEj2uSHd4BeXUDxwPUlrF33GgMKtJrpxLPX0MZBxrlxean3hk6XAb0zFk12ugQ
Jzzelxsiiw08lQlCegQj2YUjI3Dp/ypohelB0Qm8bqRbhsiYhGwOeda+J6NAOxqy
MjhradEEGKZDY9qe7ISyojKRbXN4952n+7ojBZPfBJD4hDYV7Gaqaut4SxmjLqAT
9hhv9EtV+rViYc6yzkVZg0FhkG0mYI2wqWLA8EsfvwuBYxC0zRzGv5HPWemZnRP5
ILi0J9rOW7qs7Q+Jhnt1n4Iu8sVNtPWvbr9e+EFC1neAdMKQ8fR5kbCCjuolg7iU
jQSVmaUXJroAhDp/5XNrl9mhvif4hcnBn4UGmXpHievfEIBJEuIQyjXrXglcnDeL
91Nm3XgC2kK1lkIXTfh5alsbkMLvE2yH0jpeA0PGbgKu983WUzKOMyijXURk9Agw
guWvfanH4kdUQbECu98wD3VkrpSwJh4FHdr2gIk+4IxJ/E9ws0EOX0bmK6e3y4/N
Al3qSJl8ShFYPcoKCqOXdBB8aaLBfzCqxo7T+7tUP+OyEXAoxt4Pnqkg7YWZaOZ5
W9V/5TSR41BpuZA5JpSucTVr6lEWHnv8PRlGptZCukcbXaMF3DTV8qPCtWRgY1En
TywQeXgjWd+QD300W9t609MljCHGCFKcH2OZixCt1a6/ie6xsqrIEjKrn7sAHMIK
QIJNx5/sBhRFLaeQ88n0WcAypzYIPLU0AP3N04ZEQUtMAO/TISDTaE5Dbw5sNKX/
mwubuXX2GNrCNtpXxZ6ua4oIMmaqZVBBfGRVoGKNSg8sQDgz/XiZH3KfdKGn9gzV
4aPgsi2wzNfw1KtRhdCxkfCtdohpqbxutnVnF514s26JMPFWG4b7/+RPJgCL3NRQ
NoP91doQG129iNJD44XDYPEqB0jl9QYIhw9AkepgRnqFlWLThdffPuaAlOUs8J2A
l846VVgTw9M86uVnAF4UO/b7NZ3pXNb/PeEfxcYRyBl7J/RsR3saQBbF9D1xQMp+
lnLbVya3zmxFC4vMdPxKceUy1xbaRm5uZXmXKuZ6hT6Dw6L5X0W3zAiBtD9NenlA
X3SQKpTx5h2J2aCVJQEdW8/7c+kn1kLpJyIjB7CxacFWuJQdJk+h09gVuESSjynE
hKpE4aIn4jJS0U3LiKY+NJwCrvcnjonxs31uU7jg6MsdW9Qe4+0suWy0xbmU1YHh
eFvSPzVdUmqhs9BSVZjbWE471VbZn+J6xVZYQ+EC9+oNEouSlRlsAqyTlgM4O7AW
NbYehohWjN/HscTRpu/XUGZPuGgtu6kJLewH1BYeEr40BLh2CM4loHvRnhfUo9pR
6dQSbS1SIGrXj4qYJDtk72nT6cuAndusMNfECZngyVzi2xDRcVDw6Nh5FCiQoCeU
7ZoioAOxxL6CdmLyTFpvh8ii/2W4trmL5sEoE4uTZ6FbuvQcb3I1Je2n8/My893n
9OIuJ4jzJop0Uh7cAvWgQFZ2gYeYa4KnbOTam0wfWhTIScCRB4kQs5R1OelR19Ax
TsRCNu8pfU7wWUTsKRYwkx5k7qSthdZ98VwCy2oxPxqvBAVGOW+qOsQHcfoo6BwB
grkudJH2Y8XYggARgssAIULa19vQ9tnZ2bmFb4EatFgdIpTJ0b3BjhvAHP04dhmV
IVMdbP4xaQpbhg/m2wBsmG3l/InSV+1GHNqzAPLQi7kn+oEPMEjeeVHmxpclTyQs
J+nKnR7qKjQ9wAkRrjpZk9Mk9t+f5ZzbPh62Wm00IaflMkHXA78pYebbcS3UAspc
kVs5bLZjKSXWFWMmKROduCPapGrSxxpeqWDJvXV0cmQ/a2SYXK8iLwTzkRmMiwCP
7DGhR15y8/j19WNJo+unFI2x2y9m4pQkFFh8328hNreXGLO02nXYp1VIfzjfRaCw
+Pf4x6TCgS5rAPvBnextjXVqjLdR2/u9w5Rg0mPax9ZF6+HgkkNU4360ZSUrcn3E
7zd/Yf+SDuUQlxHKu7jRvzLJiyyOAbJvCk0tnhKDuJ6l/9Jzjk0JDkIXWwmjj6Fc
3PEt+49NYcHBYJmKvUyTHYPaWEpZKMw/VPRGhmx4CNx2YWW1ZxJTnEm+4Rz56f/M
HgqslzJ4uHD5vXd0iZTIibmxobUOhv0phVxg9g1LzM43QbhVT5CC46mY3WGxhlwr
QHxPMbzYzdUscU33MeIxKZba4psDVx0wcrXFg3BWoCK05FSHpMfLN6SbwRWR6kYI
//+A80sSNnu5lJ/5f/+kWLGBDicyOfTDkoiszFP611e4IAjYb1wwC8aqJHRQ2BY5
kv7rEeDvacVgA5gc78/BvuI7QmJkC2ZrOLSwvylMnmYlqc0vQmKiPc5ZNaByVXG/
JSPTXcNM6JnybNba7qhQPgnWX6zrrTeW6GNYGHKDWZ7DsEehQgJ+4DVNpEGgZadt
bZsqTLQYFB6oPhEbvnwB9bHyM9dHLOJW4eLLEsKz1da5DSpzmLg5qcXDSstu2yX+
QPjHvRiiBqFLGUllgt7TOk8Gq4ehQ2cjAbEPtXRpeEt/8SALpF8uIVuQPxw2uiip
kRE77lduDSptaP4+z1razphM+9bCUqtQ+wzsRjAFmJfncyBj8CQGLm9Q0AajnF/Y
yAoTzptP4I8kusuwM4owgg2C4eFnOLX39aRto74y3qrI81pRstOyQT8XOmkkYA/b
jYMv1BXZ+0/0YktlpORxLtzzusByiLNpvNCyH4V0DxSmJdsXkfVO26J6EfWbhTmZ
33fQjxXWH+T7HNkogYUsU9kihTUcWvlOpMddVspchXMBH6bOXITCi6kwuxXV+4sP
ne7y0QZlwj8kCXNj7EeCF0MoAWmgo27I9PaEYWkkh/jy5oX7yo7mI6CrtqTG4fM1
i2F1joZ/ev871TEhfN5AE9a7G1SiI+FLHFCkZANIfl96H6tokSS7dH7BvbCbB3JV
Ii2IWo6rfN9bgq5OyDB8y0ROE1oI6TiUaTUhsmOEfh6gtwunXtAXlDzgiCjqMHGY
4LFTrWKVz2rtt93W8JsoejRsd7hZwnHU99b1LPYb1sukxriTEe0UtMra+uft4yYv
JXU/0HgbanHmLbcbejaX+YRDWxLt/lNQEv0P19IN/IWoAzabf5d1q/AFea0D2dAz
rAXYXDBYMdwv3t+OyU41VPqKWmScUYU0/BAgQCDz76UteYwmIQNfak6DlZXgSmOs
7MEoDaq+LktMMjX1etfcus3JGuT1gjPtWe6LVCglTIahhJMRx3fthnIUcQozQHFb
5Ckmf83VwTr+VKb9qXIjTL6CuzZm+50i9zs/samNJsLyR+ho+z3jJdfqgdhlgRhP
sr4PtQ27L4nxt07Q5Q3mpteZaHe9wNaruf4LfenCYMn5T80m7DU22E/o6s8bvhtg
ucCyOGE922aOndF8+/JGt0nkft2Ep+Kqio3lSiJdTB0NQQFRfPFSByxX6pL3/Cit
1upgZfXFMzzuIM/gp+JjQ/J86MjaqrseQ7p8qpmWWN9mhUMCBkD1K0wReNZ7iBaV
s/TY7dUzDliZyI0gu6PDiMSZdGcg/waWbwPvpSzIbFXaSdeJdm6cF93YrCAJUZ7t
ftcIMU3vXvhSIKsT9bGqISUrpAaiJRtghmospU5miYjNwGNGoMbnIvBlvube8dX8
FDVdgbsxXFwZSjTCyz9D9Q9x6KpCEQ8ZOnoyCJ5jPEOvtWGtRoY62Plb6Kxxs6xa
bwY9XC0b2du8Azabm7CwoLjKVggiD/d1fzk3X0OCYvISPHUfHmPNc3CBIfYKPUH0
Iot2LX57XL7wqPzuDYwZT52d82vnsFMccQQHP8mHwdftzWh9QxNq/Rh87g6z6tWo
4vPs25eIM7/1PZb+5cQUPvQpfburVKgtXMVjTXQ0vT1Vn52Bzvv/T79Por4NT+pj
dP20w/BznQIKzj7CygUNRCKt/RSY7g403lbNm4mnjz3gBnwXakjUuo7vBY7SzIDB
+19O6eOwFtTInwzZ9of240K+ejyi26Gh6e3s/QZFdYJxkJ5G2rtpMDa9wFvAkSW/
LNJEi67OcaqNLZjUeM24OEURM+Iu5ZL49gK28uHOIweT8QUlbzCynIxWvH6GSC1R
kJ09MmJtQT15Bh3HEGHIK5t/uQYGeLwX/0Qm0pAgfCS/+SJTAxY/gxJhBnJM42rV
gPCOX9ocyYwY98qTWxGDljSD012tKcMzXY3UxayljYN97567hJs8+LpaLMmYC7PV
I4KCnvc5hzUxF6dbwkYCT6ocCq6OnGHtKyMWWyWwcuPEYCPicYeg3QC847qNutBz
zEeT0qgU+Soe8MeeVbdJ6vY9yCcxe29ppGi2G3o24rk9Dj6F1HaU72lvcLJWjw6R
UL+VIEv45c2Nh1VSOlo17MLLcqNjQI3ysvAOm6Rxf0AcEQ8OlxEFAJOrKdo65goU
RWpjL/9dBfne6GuWmA4lBJta4a/dm31wHhEsUDaPBOxccLRLze3BjvD/VGT7CxP8
9lsBxRgROhfVmGkOwHRfIaNCA7iS/qFBOQ7XcoHjiR9IZ1lFNeXyyhrEmFJY6hQc
smMjRGajESMEknjRfrrUNCU8cAUl2a7ms1LlcHqT1ADEjMMEE43b0H8fZwfYE6O5
IRx5s119vsXpFKbykBYYZpXuMnz3d8vNyczbs6ytngT2syzeDeJcMCoTpf2qzJtx
rr2N0ZQIjDji53k6e/a/yaNG4D2Y178mL+HFXMvyrxs0w6A+pp0lPcValjs2b/P7
9mBrl3VsrItRmlu4+ag9EsZwDQKu5FvHKsGX0nSkUOYlo/x/TFT4JDvso8H0EPYE
LzQJI040F1CMqxBycom8giOtRMNjyMZbIFfq9rgRj+3sEmwYJoY1tlX4ChUEln3g
71c3OktzgSyTpOd7UyZHtityvqT90xug0VwFrqcAr9AEXE1iw74e0jiEh0GowUmd
2C1cy9tX9rLkFDm690OIkqE8q3LqJnp9cUVO1LzL7DyoC0jvKIa1i3a1VI7BZi9n
DFktxjrM0HffYK0jQ4OKl+NNjpprkXVI13nJsStRh1vh/UPaPsHhDoHqnQNTNYIp
VjLkOpUzrCxy2gboitOM9Nj96/6Gd1EHkpXjzMhHmLEymIToDPAML7EunrfBHlrD
YEQiWPOoZjoH4LsY7VIMO3wS+CB0xR6m9nyDoiSD1aZk+QzN/+iPiFzBVXAyUGEN
GJ5gTNW4r5jJnkFXc2ClH1Ad2p7d/MsbNzAzWarWim2DdKJl+Ou4vI+CAfbdFQL/
j140cnqJ1JR9pa6jwmZkzr0/wReq/J646R63gaVu3WWygPGlAfd4a3+gkkCPkWYc
cc6EKwQE+0OqNVhyEM+fT9VedAB3257UJ3/gcPYr3BN0kB/pnZJOj0cdyQMjPv65
B+5w6cSmy2Pv+4NKwjPc9VLMtYZ3buf0XQbm9OQ7BW1075MDx9CuQJ0yAFFn0QJ0
DrgBZJvYiIo5UlrJPpER5v319tB5/TZ7LhUuBlQ4NVq98TgQbDc/oyT8QGKERSal
wNUb/BmA4a41lBaPRENZ1w9jMgpMd9+FwAuyr1prOo/2/WnEmgBrkkfAVVu1p5we
YxeJoOX4PyE3H3J6GwrjG0lERQWH6tNncVvvZNcgAmLuq7SHgdCTlmwVEzZa8cYD
mPokpP/VxMYVG3FN3dvnsw2UeQ659Rp+CxY5adWVIC2I3ybvE2Unno3O2pvSdROr
xAksfh2zlL90Y42enIrU71ctF5tV9aGkqd3BWR3a7HFSUcmOey34x+k8tF8KhXaL
AxmtRvHdbaF+SGMuyO3M0wejLFrZmhYfy4FrBp8JJinhiPBsRag2UNWxKCaNPEuf
cmQRLKGMoG/dvVPkN+7IEZFoW7sBKCnfge+19TzgqyrJF7NsEOlQ1e8i2eXrOK8u
6bzBEk6ypGsSl1S7TpZfyzjIO1DfjuWBNidfo0URuJRoJhRZQVJzU8gCsEvF1eU1
eCrjr+enVZkKqVJIrxZ1zOAmaeHgywaplJFqDPXpAIkg9tj6bZQxh1Gz9+me9DUQ
lnj1hHFTQSqUTz1mV+3Rh+JbXKSleXG6DmSPuIwwGFsE/E9s9quGbqQ5rl4cBlVJ
kuU/sPU0Eg2FEfzqZLHAopJZUlrm67+DeKtrjAwvpiUIXZkLVGuCGkVEbNb8KVGt
iptTBOTgS0L9Mb0x0JQ7GaeAL9/aoEfBvyoRv1du92HEZOxUpWB0s/XMeeImEmI8
oWbk+0Q/W/O0mRuh+ibs9jl/ViwRTn6zunVVz0YBqZ8lO39ejguCrosT+MYoINKE
4M15cbVvHizrP5W/RCDYAeW9wYmHvkK/DFI/PMtMsSWIzRb1Fcw4Fqs0DjZFmMwm
Zhd6BdUqvR4w2TF703wq0bTewbsgbiqvCtQYgoKm2C56TmbNDCR6BPl9MCJqqqDn
AbAiiE40SlDgldAl+VcfPrwa/5rfLgnqg/kpZt8HBYk9+7KgCAnB1PGx8xJ29iXS
JMZ8ppoGPX3MWMQ4SfRxw94qbLRrtuekdLjldz/+95W/uNBlcvisNr9O/YxYydhc
yC3qk8gHNYBMh5TUV/4Lg7JlaOWFzhQ7giPS7INdGub61MtFDF88qCI17Uqa6YlK
iFrhk9+69hvShAaz3k27F/Ojsyp4jEjl+0eCkjlBzpMScsGfBQqkNzShMdaLnyyD
u+cwWjlCDsGWc/80KcPJFax40H10gDeNNDaqpn1Bb8p6Ms/Pr/Q7buQIhGDY5uBe
EtUcwCfOwyydEMFcA7B+bODXQYuOx8Q4qIXxRiAwIunkRUdCdl6CA7wM6e+6TNdQ
Vh1WuSrz+7kWrPy1w4MksuCqdGBW5I0e3ix/+EeouzTGB+r+ZZNGUb+7JMkJEhqi
2W1MlVxs3UyilcjuTC4o+ecsIexZGlVFY0h0IeeIeLEJxq+eIqE4M45S/U3dHJQD
iwaQWmhcORgn9QzNIV3qtM0mNRTrWUxCLXWUZilrmRZTLOTHtydLU1p8Y/F9QTFE
H43eEEQQqddkzzfNZ9eP9EtUx6BxhI9Gg7y4hvf6uvNSoneOg/6kv2o1T28Ho83I
qjQ7puDMeX2MmKGikxvlVAMrIxOszDohb0dAeFAXX3lVziDhMyb1DdhYlq146sbj
w7kWlcDcVbDQvO3IfQL1rRN1ZfUt8InM7U+bz9vj5xNMvdKDR2lEk9ZCSIYOAQOK
1kT78NKdNDbJ3eeT5PCMoyx7IdeInxokUjl8fSvTCm1cvCZdlHMdMYUPiOkXJozn
w0KLT8ANxqvJgVPV8D7+TwZcE6mxvO8tGybPiKSdOArq4MBbaEhBgTdX3N7cDN9Y
q0QPgf4ryMtCtn2u8POIN0mrttGsYBv6qmZOQMzSmnw679Bn1/+6wQth862N9qRe
a5vwOD4lqq5hhJHcn+c1hkMPg431zc+un2SxK8F6paYaPEtOfzGVjKUg6KhrlSbK
2aEHOYRgPWpj0sgAspR34DMk6rZcW8p+pKsX1ch9sm7WG72RmC4RAIXJwyEse6Xp
/jpmwGeinrfx7AZE3LvcfL/D0F5oKiRayBCEQ8+v/IinAFisYg9AmO09bjaGfer1
68Uqjp5NiuXZXoyk4QmrcipQ3H1TPqcPct1lHrO8txSL6dahziM+gAXQOeeylB4N
EP62v7b2GqufedbcCZUiJyXGtbIVyhEtH0XTqxzo2Tn+dLVkSfY4zBbMWEH1lduU
s0+VwuIJbKldTbBPUdyFk68IBWcn5g0w776Vl5wSClw13dqz9LWXGRHconFwkX+2
WFks62/lg6ExX3vZ87lLF8r+U3NyJSRQAb5R161HmHf3c95LkjR+SjRfPavWhpzq
Owh+MyXBKcy4F1/0ceZTqho7oqEbw9LwuwpZzfysY93umoK5KLgP5gLCIYSReo5n
JowPnpBl+hqgF1dUqFRSZYP1UokjchVrZPCF6E/56XSCmYKv3c70ZWh49tdriOKc
p+BOmmTulR/WK6S9zbFxD87DRQNIIg6WCvpXJPntpcrDNRgjIDD4ohr47DlZv2/l
s+V94+u1NgmKvAXrgKDPDiuUde/dLcEy7SBrDvtsYMR8nYSYVHIhkBZTPef/K5JG
tGM9qUhjtMRFZILXgjIr9uA81HmeVHWtwAg1x96yKnJlAL3TKJCnrvOhZ6W7Mpf3
sSBxaxc16jiITtBeglcfn/YVcQUssZz/ik52dtdXt8+g5E3Lvk/hymUjYmPEToQZ
3WM/uLFHxWhzV6dNUSVuOZcpNP7fe6G7hpJbAhUzTQSjQ7oKIUCCaNlcXMAfWTCD
KxjPuzsBJRGkuvTSXv2y1QJOvn8exuobQ2NVnY6h1wZCBmog7TmpO6yZiNwmn5GF
Gk6CT1gsl4WQbsMnd2uwKdbEpIDhlqSmmlvOtK7g6yZSvCms5GWfvMVniRUqUx+R
6kVtxvPXY4SJ1aM1RA+kq0itoSH9oVjl7htdMdbZUDFrJa1N+4fnHjR2JNzu75e2
5VqYJ/J3b4kuU8f7YBqe7kxxSRTkUYi6FB/pqjDU1Vx6bwT7XhDZ6DjhVqQQVggc
uVkQzDrug6F1X8eH1yZCCVj65L17eJBFI/IFqo9o4tgGF3TYh4ntSH5umlXuh6pV
tk7QLDl9aJa+ht4exEYiDfT6QTh6kCQbvBYYq+W4nnI/CMIRIuInbv9YctIIVizm
He1zYdeIuxR+ruKEAjiG5UM5ZqhZ7WTqbnuZrK0Vv1iUPebG0LtycSEbo89xZ+rg
Rq8ygFPaCjSu8JBRcR7SNAONksM4MV/54+06DDoKzo79sf4yky0MrWInNO70Xjsw
TFMxCVQd8E9hyuuFy6zFYRlxPU/SN2nneh3bn2885CSezTopFQzIBq1SzC7UoP+D
KJCxonrxZQ57eg0I6WAO/rIzxdYaG2lxhudeCOIEXyccdXLXQorPqLAc+NjT0sfi
cdqOI7/QyMOXs04CyFaeAz9zEqtq9CW830am384YFVFRdQg5mFxmYf+29w1GdGLC
+b/pToGCkmPrs3v4P+k+h2In95lb8ZmBfNhtapdtxwmF70Z65583SY9LZsjMQ1Cb
eg2mNgqeLtyqNMFhkT5n0w1oX1jk0+DOIcujLqGGQeL06STXCs3V6RKUsOK58dfh
PZzpjvW3k285NWIsigZBNjEHKdcvhF0TE72ZeJRrpiwJ/fG8i3w5mNOBukalLVtX
f3WsC6ArU1OakMZoRUJekcLnpZ4lCctw700NxbQkqsTq8L/sZBAzdZ3iD/4HXAv0
ByUao2CW7Pf6J2kT5gkg8pCJxM51t564ClAHTHkkP3Mv0EyBJZ5/g1W2Tg439+rU
208J+4pacsebuv5YFjfpk0EqZLysPoPCTFqtPApUU7cl4yNRWQXIxFdfDReQM1Gf
QWnCAXyfmJh/rX98vYSLseaPA5sBWpMC/GBbiVWef0TLvWJdTAA/+/vrwBgQalOF
1zrr1Cj4xhI91pB7uHlpbzzfDyJt4gjd+85NIBTbyubC3pDKbB8m3xMvJo6M8pas
cIpEoIQcyUKxf0n8AW6s9uzS2ZyM2cJQlomcAAByhLkNhAGwL6nEmCMAEIJGx57L
V3G5kuE2drZdORwije0vP5m6YK4zvTnqZ5skjsz6rz8xO/Q19Iau8Ixf/ZnicuPS
gq6WzsMp/5v7I/9AxBWGKNaT6yO0U4Mh8TAlf0IFs71bUYTAsDmkY8VJVdB0IjBF
RlK8u73guZvdXKYiXcxz7ZlRokcEP3KMIjRQJkgxkUH0pTj7OiGKyBXFO7mva50z
9s8KO8hGf49oevskMilJUaX6diOrY6OZHe8zryiIgM1dHDIOEKDZjSSy5BfskCGf
deqkZBU8FnLbpBGOaXfrGiTqlWZ7VVg2/oQg0oNSRmfL2jsHZtyy2fp19JguZJ+6
E7J9s2Tdslgieem4jRkwF+hvHQ6G/JznQ2wgzbc3Tnd1CP/QCsYERy7CVWop2GML
kiVXE/xk48rcwbi8NINgANrusDbF9tabLdXJjfuBoSdKxGDPQFl0kW2zD5AOSfrI
wVRuRE4F8Zh3B0rQUBB1GVXwQgL85rEsu2quCiAKGpfNPy8iJGl1Cf2WimB2qP5U
jw1PnXgRlA82sumHd25JSZ0DiH+OqDcMl9yeC+ihVxkrFBOpSYSaKNmkpNsNGpau
1sdcNySM0lGOV/DUO6B7dvwdfD5O/pdrsudvBIWg6nqRLFr6iciLeqjXI98IA5wu
bVyGJhoPH+rnigT60D+xUEXohsHnhapCpxX/XKSo3z9JPkSo8898MBKdPtL4m92B
dkCvMaG2dM45FAuw/dsfBKJQwLdidDVgTnh1RNgh/AlbVWt7VeYutq57k7IP/twN
42GJhaPJZczaIr2spvHjDgcbec6KcMcmFYRo0lTzdjm20riRcktC/fKQsLwXkvrO
TN1oICXO1l1+8Q4gpbNn5D3xBGAPOsvscXF2ydlB56/GW9t/LzBh4Nhd1IhcTNUQ
2Q/FfxsqQcqqxfsls+jAF0duEG7pJVghzgeA5aq1ImoBfxUZ0rU76t0Ima8DvhFr
kJ/m6weXXRKrv7OndkjpC1NI0uoow0NeGpGU88uOMziMNDHTfOiWTQ+DIG//zZux
jpzNAvcr8j1bbbDf1Eja6Qf1QL0tt88CqNWZEJOKm8efu1DWUNuD6mHy+QltG5hC
jFKCghcRb3KX1pg/SkezkkygdZyTACVkXYZJEH31eNfv7AIDs2SbwC5DxiS+TGhI
158NK/6V30prPbZeCuU5HLTeWXDubQlbpa3RLn/jh8mfoay/DjHkfKv/uU06Z6qM
cR594dTo/ZmreJtDWVV8GkRBp6JoeGic9ac4oHfCzqP22b/T/B6YNDkX2orzK3G7
6ybgcaQYFr0Zj9q0zYrvRnIN1U9N5EkH29xS3zuRXzBmq549V6keMFmzuAKj4gsa
//eJ6hShFzU09r77osTIhczqQH2qIHMbw9V5IiiqGH0qGNcOGwlj4BC0fVUCn23j
RSOMZGAog4c4rw6P+K3zaSYlzIWoBxj60QpsaJeiuro28daSY7D44ahP+YZ6P1em
XRPiXKrqbyoc8+rirLY60NsuSvNBumvlmfYdhbtV/UurLrLpU4+/hf5i7USQA6M6
170yE5mqsPJc2W340ZeE7H3Q+8CTWB8Q9LnvZr3MRw+5oxkDgMvMpxKnbIWdX3SV
mJMebhRrukwGpow6FKqZFyXWaSqXj9moaibBnLTIs3ams4F5vOG2DXacSX91EQ8G
E8I+oeSCsfWp/4YUHb0SOidC2We25z5YADi4sG+XhswvBOzVE+Vxv/QDGt7B0Gu6
Kchp2XucsVOiZ9gNQFSe7Yg+Sji3DFvVC+mEWHVqD60tlyVUZLS5PyPfZMO/AIzr
2pL/SC1Jfk12Fs+Sb+9hZeNOcrYzJynpvOGfTPLEsgUujInSVL2Tinl7+fhWiJD+
jkHAAQcQBIzD3xh8P6qIDDA0pPjdiSAglfetI5KAbkA/Z51NSvTWiDCAi8uFpXE6
Z98Un/IjqfHD8m5wYuGZhGA5xPfOl7McVnQAn55qGRqDb6oLZ+EhlSHmdgPAOk8A
ZBRUKK7NBpgd+P/U3BWQCCErXWCx+smqgBihD3B+1g0nAJdOq5RqaImpQBYI7o49
6vDw5QLr3383uaoyas1y05hmYCdB2G40oCkDEEnUhaB+iq91KjeSRXvKrjY+3zSz
hgq+KgjvjROJiwAl3LnxgSQ25Y5Uc323WSe2ACN/F20l604g4AnkE4Pv5ic95rhL
n/41qOFHSYyjnt9K9MWYl9xpTDfKUKlzLj9o/TU8br5VF5UUU4B1x2EhfqfST2Pq
+GLyoGAc+gU73DyGQYXjyicH3oR9md6cw0P/FpXg8Oame71DD4qBiQtb3qbD2Jkl
Lh/EPN05haDBJ7cX8M3As0IBtdc48Uo8ky0K1tFS77OsT6Jwe0fZsSV3hnNS9exr
g7aVJLjK/aTSO8T5R5zzZydmw93zOYc48za2VUWUvtD+7z9zRQSV2Sx2E1jU1G6s
dS3itF0csgl76McvwFt/1vuehTaJJIEdQWZHeS3f+ximoXpJMorKKbf+cNzzQY9z
SQkDfD+/PKLqB/hXVcaJhATqid3q6kUr99JfkwTkw7LXiBQwH0/lDdAkf/EImAFQ
oxZK9YfxHrBF6SRB5G0+74HntA8LXnBqvLyz/5OXbu25vP5ItEYl9vNvMwdph+Qb
UgAGh1viCiZBnMafxeUgn8R0DKOxBg61YOzhI8tNWT2BoSas9Uc4CCKtBvXUS/Zv
zO7+fQ5ACV0HR8MBO8y9NA5PuNOPz2H2l8raDbFb/k2r3RQcDogJoo7NrXKDGplb
/nppho0ohZlvQiM9+l0mCm8v6DNgFY/VobHzpbyRPocnMG2p6/IBhpbmMP1DTbdt
+qQ3IPIcWLoZFGwR53btFciEZvhtNhAxMlblgKIE7gRbytPhgaB0TPzuL65eQ9/v
SQhdIDvm7F9uylOKb8n0kXn86TA8S+e2xNiMOV5/4pOwe9vf/PFr22gGh1SsnDzL
StVdzAi6vMez9LQTreQ+2ZpXWzL04idFcWH814oJnAa7Ja2SkCtlni3gTWHbbUqw
drek8aGpiy1t8BwH/OalQcbDKWTgXZLlPXN8T7B0NC68U5s/o0GBq7MIMnlsroU8
5P8S9zKwfbRKrAg49iSiMmBznbZHJ82iCB8k6gHJdOBvnDXSSqhzAMD1r58RCf8h
AkmVFU6IGOvLZlxImYwyxZy1JyaDt3SqxSeuPnQFbfdCYDvC3VGaQT/5/iMe7VB3
ErgsE45EtOjziSsDmwQDJMUrZPSVoFcJu6ohkkQMJcDvxll/CWDb77BlpJfbTB+X
8WxE6eRec3xi6+k01/htXf+nEZgK86gZlDiyq/I/vv6wq1/7+j6kSO0y6lxxddd1
dPlskPgD6v2S4XZ0ECzk0Qk9XvUhS7hN+/Rxeai/Luz+aWMZFk4iL4a3iQTImoQD
+OhDP47UWCbucExZiF0VwKNnPC1nYXaWNyzjVPTlZUOulSeuxnilfnzQJdgeHmC+
vZ1eEM5RWEjB5hHYKO/M6T6lA0eYLSUA5z6RY1hQiwTTk1oC7kQGkEQ+iHZsPCga
bdaaanZ0VdHkNnNOPKz5GLzFC3EER7uFrFBAeHQSu35EfvsypKdJqvK8V1PlGXms
yobvOWDZPuoJTSrkQMnQKcJ9HXWNiO5UhG91QMNg2VwJtoiXYWx77PRKkJhqYkVb
KX+M6Qid9OeB3switGvpcspXOLLfJKYDrMj5FRIuqpd5rhZsW66xtVOzlBO7x3f3
oX7bU7wE2wvZzGAroROjUw5kTHyhu/CgusFGPU1JEZizEM308OiGrRKikWd96CV0
g4XEIXap30Ctee3bNoxA63aNP4o7dZUKro+/rPP35tnY5c3v8bGtCDXNFvOCUtnI
IXRJvVUks8qd5nvS5Ofjupel6j3qXQ3HbsS9I2eqyHT9dSPQiPP0XRVxujsLC/P3
oAlOid2VY7iV4eRFqNk3dWjlszY/ReiO/wb6QNodk0laFC9QdJYNoJXTpN4Fc5Mk
UYCc1u922AXlJ7W4GZVs/d1MRwAMNkwovSKvc9/2JvMh0Jw6gSQKi18mdaHDsa38
NtM9J64hv/Jx/qolhVihWB7NPCy6qu3iVPJ8/CmD2kaPSxNi/sLvLygsXd3SXW47
t5Dt9vjqLG9Hq4TvPVIaaOAO5325J6a0r584duZbuPP5AwGvrfK0aUmtmPwsTjaN
KluIlfPHP6GMC4gG3vjCm9XRlUqE1mjQKAykso+Ftjknvx7TkArmQVYJKVV4UJSR
Fr4uJM+I6RqCIa3iUrjGIkqDSTK7vyd9YaE3NVysR10EXq9m6WLn6/6ExqeAjHza
60LTaQbcr3VTQRZ4bH06QRzZGQbtoZALj5EjDVJ4xogHzf52gg0CUvA5t3nI8bih
dr6h6fkDz1qWSsLdlC7x11lcgQ8SX8krK10AO6dO8J1bG0MilZb/auBGvpwowW/N
4gWAN0vUpuCaKTpw0/0c4SlQY83kacNnll07ngihtYYkN0twjSPpj/tRVjl2W4/0
zWKIqzmQHmvigIYoEEUInPpx1tpNy3HfFK1PbMFAHZx9/A/jbLN+Qk3rAj18vw0p
j8O2XTIGGP8OdvoLQVuk9CMZFyGWbEuR5sgEbuEJ4kYyaIbu1pHKk/ntgPgqH7cT
cpLLvEK6FWPW2Ja/U5NidnrDlMY9suszzwAEt/11O6isjwLnx4YfKg0dX+SxLoyd
y67kVxNlGQnDqT7DfPpoMX/DgqnrOp3Uy4GGJOulXdB9YAzxgPdErgawui0edcd2
nzCpKpgCNTjzTbKlqqWJsFe7tVha9gYQgQ6meRCPDr6nu38kqubio4UPb4dsI4Jk
c02R1YOnqgWD/t6wvOuUIU/fj0O6qVNvgq/u2EazG4V3MOvET2cSD6SZ9otqPhvj
E1hzdBPaP8iv+q/ZNr7G/V3FYorUl61ttTs4oJOD9e7KIzAgH7AIo0LgkCzfYMwk
Ev6rlApwABpmA0XSykmKIwqpAa525tCEedozFTf05rVkI8yrWGcanfj9f8pHxC2p
8F6wvIAw0nSDZvgVhARM30PS6q28JWq8RMDlIjUHLEzJ2v7vKglA8Ox3KWwQ0dHj
Iruv7FtgAwebc9qs9BJ6wHPPTq5R+JQJtmteIC9VRPKxwmTMEocqFGvNq8VBX8OG
gKIKTDSt6di9GxL4dMwu2LMFdwNdRUlNVctTvDXgC2dJypNld0RhNUSrPaecDQzJ
hTn0Px8CI9nmUmoTOpz0wN2lagD1WB4Y3f3HOEFof1j3Zi1XDE5a10dMvFkf+D0s
WtgV7cBCVt681r5HY0sL65rR9jpD40Ocml0Tg+NACCDZHNqK303IgfKYbc/QcEk8
ffBU2o546bOJNmeRePnkOgw3Bc3fQPyKdyYCvndzlVYfZoXw2u1C2LGiEChUFeY3
XFdESLpSJvfX1n27YN6d8NvbPUEMzEuH0CKZV5tC1RCSCySvYYHPfdOgPeqeSRoK
Ai2D8u05+IGHlMfNUrWE4wQ8bGcOgQ91EOkoLZtY6eobqoNFq18i9qFD2o0dPi0I
ZdVQFT8x3ZYQxEV3S3djAS3DY2HBmmc/HKXeaq3Udu2i3GvzwjcPfYPChu7mbJOX
tQvGkic39GSWtKfxP0Rwv2/ABj7U3aRKVg9t7GFrWWWwYyP94rJrPBsbYFuhqpSa
5RiF/Pts5fLV/lFjRfB7Mor4fM5B2itrtCvnqYcMfi/RTbdMdOKdfJ/dhD0fQbc0
kFyZjo699XgAQY6kyJg35GYAMWmph+4m6iV42j7oeybdQY9EkddJpNZKDHgyM+TM
a8WoYfrppGAd6B1Ub7sJBk7fT/t1wuEjXcHgq1Udlzn689y9PT/ITle25PAS/azR
r5y32tIVe+/ulMAkt/u8KzIW47gHMbZLZqTyG/ztiPGEUOh6qqXnhbYLImU1Z6z6
VAarbPU04RgpzNuMN30XTUxJoDHCpYoWCYalRvYHcG6L74j1lgudKcfinoQr7wgt
L0c5ey0GID0MbQ5Z1IK81OwayAOIjZPkdhcycPmi5XKIX1apZWnNjxog9JIJYH8T
MU8/HI+ImSqOVElQoyHiRgQ59Bh3pjzydKjdAipqSZSGzwbzKd9/tQDXZlYdH8B+
hW2fyjW8Kz4oLXozXp0SBCOsuU5iPwYEetAC47fHqRPKFS+v+hJSTEF4kOqLSvWH
pm9ypTdAG4k0SuhArU7MwsHnQ/+B25xHn6ZC/duWin9IMfuRkLrppAxNNYYd0YUv
qzKThE3CF47comBWvVP1hU/wYArJVEJK5fjf3hLbAOOFj4skpmsSmMtZVoziiBhv
cKNsphra56dlCBKxJb6S1ySjXu4SXJFy+StPWZaL7c4T80qv/FpzvALcC8t3k4Lf
NgMXEBVdkeNPDfJAJeYiQ1NteKOnK0pnx9E8RxIqS86D2BMFelOmMcHS+gE7seRJ
CSTpRKf1OSzR0upfUaK+b4A8YrlylHm05wUd8zde3PO8aObElDceiHBMJ7TpXgeT
3MEWpGtFQZo3JVLPqsrVhoV3m0kYJQRiBHYYceUFvKJoI0j6IVdmWCpowkb29e89
fEZM+JAqy3wZ8Xx5Bpteb76daNL7nU8ZZWeBuxwWhieaiRUe2qrF6YH5kq9+2wDR
bsY0fKE81gZ3jiEc4gM3RF4sitGxZ71IV4gbz7EVusPCN3XFEBZEk3mUE3ZyplWg
IKLcsaOVqL1P77k5WoYTvUpVwNzTIWJF9RzDEnZtFaGeuLQ/LtMHuRqYPNvTSo81
/5JJoJRSUwoaAtd+XvM02tBaI51cg+an0k8TDMfJyZhomyYUddWZ65a27pZuba0I
3ghcS8N/iBWGk4vv8AFETPNUI5wDaCDT4BML72o8wDzC47hDEoQX4sXyplqVzeVT
YABgMsXHjCFWG9vg4ZTX6zeM/XO/RVTFLvAvPElS1pUQa+uQAQ0it1Q1NlJAQYjL
AP0h8AkZDm5IsuV4oFs1qhHqSDtssTznbKPAvR33su0QCpA2k3alIA1KMdKdBwwX
I6NaoBDRTcYMXxQ8t9d4B3ngpDX7HdiV3sD+0aO0eC2JzRkoJ3U3lFIxjNUOpFv3
jVmVx49X58nF8pVBkNGdyFoMd4mHNDpTO+SRzLSPUXGgumEg2wWtw2ATVWEhfYYx
Ap1EhatNM3AvJx7whU1u5bKQu2bOo9T5YhKHX+tazZ93T6v1OGKgeH70MG2AEMUB
kfe5G2lKIJiquVnFQLL4qvsy0ykQETeQKZg+GQiHpvoHQ6b8ewCRYUmwTPsFWqUF
gyEK1lgynyDXCu6yU67EjIgWpg6XvkckNLbtJ4gkbtF4CjcvizvF3gHw8GE1zAmc
3fw8xmwccO5qxQVtF78FupgdBl5HnYw5nIPzPpHvhy3D6KTsDIwvACfPEfdflso2
irbNpjUwJqt85rLCmKvAsuKS8/AyFkMTCfSHceRX0WwMB+gqOnrI4ga10kOp1FOY
STE9a3sOoK6vpM8rZLP+UeQLT7FIuHOPj2J/avZvOtz6rbwlDdimtKcdTlDDoim0
zdiQggRgvt8B+cucNM6b3/+EM491+UFMfF0mSbeWVTpXqOrL+9ZweScLrEAoE18S
hwVfZtxoM2NK+Bvj24u8UUvtraFS3dBXkU9tMNBZkDC6vQttuaXlnCarLdIprsvo
2Lflik/qQEwtEMrbwVVp3ib4SfV5dprsZs+CANaZ7vVNygKG9cXJN+taMlaCD2ZI
JWUijUqtuQmMxUKXBUkj7TQvPh3lGzINAaFKuXcqMzk+hgv+qpnxFSe3OJuk77vI
rhG6syAXofeI1xJy/vndCC2UiZ1h1bAld1xDssxXin3CcYv6WMRnLHLOTQeLx/zU
IPJEvTDJ8hc7HpteDl5fIIdf165FD635fUwgyFfJeqCqmq9KfFUy4mpaucCswEhx
ggWfb4/wJhUbtnp82jcuyVx0lF5fgeVxmZ1+OSYc0nTH2ZNFzkg6/f/FuQUMh+zp
g8jhyIFe4JbcOuKi5It4wemDNQ4lmqdsENtuvPT7Yb/FXsoazwjj9XNzePOxi1u4
ChGE+9PrujXNfeZcReSB0YuSSbMNz6pIQlHu8wPXfd2UXeG+4y9WbrvoPY+Wj4QA
/l0tCbKfK7mD47NWnjEx70IT9OxILGNOtWRyOUdWewk6yD38ZaC8v+KLk4xkwL+n
O9Fivz3u42nHwmTryWufZ3A9pI7g6Imuke1n/zOj6PJjUO0aJYoDkfxB8oM41z1X
los8idXlZIqoY4bItXZrSgQxMg8MQHVVHQbO+MQVsU057PAmHzVK8n5TbsWU3ELN
e2gKNx6GgPbPfGF1q4EIdEchz8sWSI9Dx8aaxot1PY0KZ1p10UM/5q+OkteYaB8U
RDhEiOj+4oR0isZG64NWaV2cpiSdx9rz2EIn/wvw7SwJAFxdSXIvfg9qAuYhvquM
1Jvsm7exTqeJNkO4IO4exKFu10ou31IZ2DZk4wfFy1K+y9cgH3VfPS/8+83ZQ/ZQ
2Epgwk8XlqLoOljV/rvLhO1fqjWpYQt/mee5kZPBCjsLt/Uyl0v+pGXjn5IIO7Bt
zpeqJvZonOqTffg1IDYxfbdzvBVkQX01QkYmaXezj2tEz7fhYV7soSJP/JbDExnJ
tDvBPd1ZlEMjM9y8d2OLTuQVLNw5iV8num55N9px8WtFwfLcF8uHxxfboFk94cBL
zCSjQmtP03DwyKAA3SlfyzSAzFlROnT0W7JircwNN3Bee8WqcC6UYq9Z1GvDANlJ
pYsUaVS/uyBcyby9h0uZPoIMiZspssDM1lgUCIsO0AglVNYa5qkuJte04J54rgr+
GqOGW1mrK3ibYIIox1hGOMHqyX9gdOWSdBe95OhYz9zpuVekWsWl+qo6hAGnX7U4
ou9CZnqKpT7y/11SbOnpZZyCB/J3L8wDcd/GWdeso7b7nF1yIwePjvefJxQamaD5
DXPriOHdfSP73ZVgwwX1Avb7etf/qteCMbYZekUVD35gpyFc/uR4f1JJBybcTt5m
kUbjvDHEDwEoAZ6g14Q5af7hUr4/OaNA+rFQzNMFZbpha8BWtrJg4xrKnzmfDUnP
OD0186B2AroTqk0UMkdVDldW8hP7Q3/G9ybd4EyhRkrYmqySPWFOn3Nubc+Ikp7s
L6sEW/JNrOR3iSJ+OkbT/eSQ5TJpOGQBKMn39flqGya60bNbT1jCl5i6Y1ESactX
YKw1vGIzW52+immJlnwX7mWPFJwYuvifT/BgJKCStkJjcrQ2TyOvitY3AsAUuKEh
jWUkpZaaPR9QUEFF1W1KDPWQXchvqgzhT+ctXOdfnVEUO5vH2HiPDyedEsSbPwpI
eY+3j1K6qIUfvytC7fwXM/cJHbhFjblDC1duWq98+2tRKZMf32hVHetDpqrEat2e
ak7xkQ5wk+7K+qWXSTb8AaAevNCUpz3qN2A/23XQZViUcgJpLMghpVw4+KZs62L7
93s3WsbW51xUIon7YuBYA3d9IVoC0yUHOIlsri7zqWp1ChIocatcSHVH3K0c1Xxq
bLJUAuCQMQEpzW0M73c0gu2rvNhrV82oCRUblUVUUOTXG7x0QhC4mpEgABAHSJH+
AoB1prvece0GrTaUa3ESUsiPehX6Wg+QFaBCjtAoYgXMqM75sjGf3me1qpEO1WLj
rkhaUchJ7un5UDZPXxZy5HrjjW+pN00zTlruO0D3zrk5PMpzlgyrUCZ6JlxMKx9N
Lj3Cn+Wnwvg7yAY7CCNSFpIHE3aAYAh4hM0Km1eTq5OBZeQ0ivlhLYJ3THFk9bl7
gyfsS7U4Vzvb1AraH4oQnkhp9MVMAnAf+kkGJXbb4CVt1r3wv3JidfB/pGSAB5rV
KnxsglWPHwK8AXq7mTkstnDjkue7fYkJvWNV83bE3F8eF5MWD670nsx6o79yXvW9
+qeXAT9CMQhh4XgAlHBGsmvTo1zEo5ntQm7wT43i0GuPm52HxG3XJiEiNGDr7jnX
l7yAGczRkDOs70+dFDmXkAnAClpaf79VJmPINBq0lVPD23691dN3rm8zTJY0vVLS
qXS9kfPioh4j2QyZPJcBBmEBdip9dg7N8J3JQxzL9V72APRXuauvNu0v2Il41O4J
05vRBsYh/fwaNZ9XhZ9XC/CnY//MsF6g/FMzALqwY9RyT18AvGpmo46oROdsD1Kh
E65bLC9ekCdV4TEzv3aLJI/e7W++7YIXzPagZpnIAUn7S+6iTSvXRsAS37s5PGhA
72fe09yKiT+B+l5cUJ/FkBgYTtbwCatrmYuXfstnedQTBfLdotDZC6B7fEDkuwEy
7RR398iPToywJsEEuodNZAzXPAF7IDNTWui/O0uaWstc9qKJsK29zJHLTmfuu6xb
jXKywr42fhKQOxph1oAFJRPwtneyqBg+PLw/usnBkmt35/T0S1Okc1qYccUIpwVo
D/ycf3L+HGpwXZcmX7Un+un+vWMPhgOz7CY5nfKPmuzIZ4lRRdsno/hzWjQB+5Vm
FU5vxYPgxWYienKZpCOYcTfk1j2MnvgHPqFkKdnxdSnqwFqMi5f0UWXTtgs0ChAh
dsWQ8JUsCo/dQXpIO5mT3/3d+4ZpRWAOoulozl4jU6UHeAUhrAd3ZYRa+1prgAP6
04wbOEgtfpSIjmy9IRSj7YkJgvrMWd5Hg+kE7pQElJP7UGTsnc2QiNi/tGEnKy24
vSLIoB68aQcY1zDl3zC6A7UNwoCXJJlA9CCzPb3UOh54+ILZdzeAPwHJgIN3fpvo
u8DyN3ev2LRojDVbq7btR17r0MXfAXdVj9bPlBpmIZkdaBzkWKwTa68A7BHpXplP
nilbarhisb/ExJEE9hqfDiQbGESrlAuzmcuvBa/cLpeXs/uFbYXYkeALi8Wcv0hM
RswxFatcfqIGTa1Z0NoFLInkHI+WRINec4K7Xq2nQld0JOmWUH62CyCKlHi3bwxQ
c9oTk8VppcmhlGeno1E7yJqWKGSy+T6UPt9itSY/Md+QY/i/nSD/dzyuPmg0FgmI
QeBwXIc7sVKFyOapZ0F4b/KiDdtzTHQakvcc8TstMrBv+b6fOs9OlBz0aeE8bNDv
LwsD5ddtl+zVA97sTect0JJ6X9SQVlaL+UIaHvsZhE6pYMsSixfO5Wi0uv/RQjO7
qx/CmyKKIry5g4Lj1hAiqnUQ7l4nFKHs7HDJVbXOK3bB1KtQF1TXk+cFcou7ozPe
OIF5yiV1upE+xab6mVxAJjQM/NzncdpeQV/e0DFk5FZJuYE8owwoojKgpac6dlv4
7RQh9XLlQZqdQDtXDI0bMEh3Frq/VfhRVUzEyVvDUTDBOZjXzO3u5anuKCsXEnJU
QcDahT/TSNF8ioJ/WEXlhT9xHZgm6tgnUK8zz5o57CDdWmtIBz1fk5RMT5p13ozn
/8PHAMuFU5snk3PdgPJnsp0+9OUxxsoF4dQVsp7kPjRlh+qO8U+NvM1vAU8SPE9+
a8PUaxY+8xcoe5U3wrCS4wsi90Z91Ofs1PC9nf2W/vt2xW5IdpdOMykkt9+iIjiG
bbkyTk8waecow5lEss0w/gRUe9RktOkG9lqHHwMU9DfiNQ8XylDZM8M8IgUd7Plx
4GnZxubtmEx9KLLz1H9TSWFfdwQ6smMh1RpXbCySHOygR0arcJLF/xIXi3wR9AKC
Di8LtQnQiNQ4HfN6Th8Bc4+bXQM6GDDM7MOjxtpv/lSZV3x5khvc35YELwFHRdbl
mqz082hyqKkGrFuW8bkNLtIuj6IhD1oQMt5eDsB1zbgOtk5t3Nj4eWGpr8VGH9Hi
K2w97pTam8uldZ2ZYnwblknaVI+BDN6xd8dCixwKgbtRMXKCzC4trXROVRQh2ABq
gU2IS0I0ZZmTgj+ORTg5w59+vT2WF9hqzLPod+4S9ch+91CXqj8THFsPmwAMnLYj
jhZZkNyQCFnfXdf9i8WrtH3y3Vp/ZRv+y/tMFOsr45vK+gRFdvrqOH4fv0+D6M6u
YIATxY1CWCLsQoiDLuQwzpZg2jFg4k+1pbe6Q1LdNmvTvhLExt0/b1VQ0orOhAmN
sNmQQSWTUBJ4aXnPUczQkZdxbJ1bbjzc8N7Lb1duPjL2veqk2ASvZpR4ijY8mXJx
na1EX4y51wNJezvZmpkUEhC/jUP51q9moD3Bj5qwtE46SuPD5PJGFvw1bdmDJk0F
uVc1zxsTYn9jW7EEPgnjbllAD6fcoM96/elPWjEKheogptcCoPfP7hdcLh7/JNJS
wdkoZCWdB8rhsRWX4H/Moahd8dpOeuotqMSF7PbIyuTNi9aicQHv5rDW3ZWDSqp6
nOPFKwOnGUhMhIajxyNs7fXn4sSBl6+b9+1gAm84XTKnNL6Ui2r8lQ1OBYS+4b0h
m+ldwnB4YGhVL0y7H0d4c/zBEVtSKRp/yWQzPqjpfAWuoRcZCTpbzV/Da5CFpJVp
0T/KbI5BCgj/WxqUoXleItl4J6mLFUDRkpLXUqKsYTdIeUiwRCT2VWwbzVArT7Kw
lUqA7hQsykG3+igNANlk4xdLP1yIrKxGI3KPCzqg6WzFUlF2hwuqIndWrVDU/JAe
MicBd+neKa9DJ8I/Vw4NQ2Riu53YMs55P4e5zll6fIhTcczEmlNYQkRnLt1/sybn
dKdCHskkP+u8RtoZc/RfTLKp+DuO98GuJP/OdRszt8BAZnX+yyJa8AxF33lHInah
Go+y8mTJCtqB5MXdWNYMxSTCJ6PNO+3tzIUkU8YjHqXtvxhNWbErtfnR2qejyy7i
Uc8nbi3l0jTc/yEUMzT319wU2U7W2mfQ0So8j3hfPK0VLy/olBf1neSFbJQ/YbAA
FZ8KpMBpED/qg3M95z8xOcIwR947hWYKEnZOqgD+Z94B/KLgd32rbAswJKrrCRO8
HojASl1D/rMKSYWI3LuV/WfJNWVGUxFPRFwZ8zHystyQThSVvYLrVTjgKrXfg9fx
+IqT5Of7oYN0gC9LUDHpdidEBSq1i4GVJrpjg3vfNRJYcQg42+VaA/vTKJhxuPUs
xCAg//oW4/yiF3r76x2ndf5fsqOywFRq9FtPJKrIsDw4xoherzKnQCFYPFnZLnrK
2JqMCbx5jZ69stxCqyz1vSbiXCAi+Phqdti1FnGHlJPFkRkmtryb3TBcThsk6nAP
WQDd0iuIvwx7CekV3TTwxTZFn3DnKwtzTWCP9n12o+Ypv8ofhyN1OGSCuKeXE7re
Q7omE+Ke4ElXnqoBQCgsvxkljD28cj9fkaIh3E0djevmU2MM49+IljY0L584SSiA
4VjenraMdR8uTmWVkN2dVd7thkbwBbxdYGXjQI5hwgbDNRSzaKhbghwahwGKoOq2
BNXb8qrXx4P/1Q6o8YfCMrtI6pfbaDxim6ZD1VE8ntTUzBTsYyYlwUQ9uGDQjwM9
hTep/YlOoqebnFVxDlrC20Cz1VvzmvpYH3HVfWyCmTsSLnmx6kN0KKkd9yYZA0Gm
jGnEKtPwvmqNsYg8oNyyZ53NuA3R7OS+sGV8udmhqgrmLtUesbsq59V0ttUNMWYb
0K9+fF4AKgiFwUCK6fhp+WYoAQFIXYVp+nRE8t3SHbMwDnQGmAX7LQs/lpTiizPs
Mh23eaiBb5MTgEjFCXLNj1EzyGsG+PFxHLo3NAgRj/uccHwYxaAwXscASI3GkKIk
Grg10YzBwcsWlgUZBU5on84svkEE5EhN/PbIFB0N2Oaxp8tocJfjERf2Od1hDgmc
Oh/o1cnu5ofZ401mYQ8YMBDASxrNEWdHacLh2YuD1KxwWNGMdvwEDrjQqqJ7sKGe
0kBkOnuAHfQ+j5vb3LBIDRvXq1la+B1nfHTvJ7iatfMVvBHLZrEVcGXeaKUAW7wO
+60WvVQhdyFl4cP173rERolaAEzLIgpz+R776VJ0WfhtH0qBm4mJRLDvOok3XjA0
CWX9S9mCiPRxlMRMHmjUpS8SfxBWuctMqg7ocU+C6JQEWTPZgduBIrYQvq9KdjbN
uak8YCO3Ba54omgyPbJKACLqE9vSB1RYn4ZasOmV0yCkDOKNuaduaV+55zDP7cOS
Ol2wb9v5eUiVsZwhzPVz+7UTCXCer0/Lu6MEu87yc7Ck/CKfX5xYE/O4b/YQgdND
AlXhrQeUBf/apK1HrOZFdmq9YU9Ys6asermlyRTVDLTCh3owCJMnY9zqyh2OaT6/
Fp3+DP7PwyasuO2/ViLBs3RHk7mUwTyOQHlwt/wVn7H+KPP+OXSQVKke3gmnQ3vd
U7yh37W9RYKEfXe4B6tTrMqq7mYkkFJ5wPrHlGeg4CUNN9I+K3XSOg+xAmZzJ4a+
EqAZWHaEDROM4uQJa+sleyLApLesIsPwqqIO6IzqyfBVDZDsuN4QU7cr7SeNo3I3
xzkoNfn1LWr7TUPbutBovB9XGJ2EQ/ZX71zoMgF5O766qSFPHJ/Ri7Pfwc6XNehu
iQeYPLHWkIFMSybfDjCwV2xvIGq/UPu8PnyyMbCfbKE4EAKPwiq2OwV+Rn+a2ini
ugC/Hcei2JdVekQ0CEAGezv1gPlBMyzn16NuUfMvlwpWJUbOGdRHtqcWvskx8OhJ
cPaJ1R+TuE2rRg29MV8YXQ1p1Tsika5hnWSbTm8XTLaYj0TXrpvX4X1qehDEi850
GNz+TijEio7/a5Gn6MvxpsbZdOaAzagLnvRxUnOfEc3I27JG9AbV6tKqziFmo1Bp
nwnYIUh75Gt/f7AaUtla9KWVfVa1i1D9UG11u+Kr3E6ypGKUd4piqutR/n8JRcNo
XnI73WYRlYkGCb4LgV23pC5MnkdyV5veN2zwHYKq0fpUpKfx4YGIYXIiOd1Hjkzq
tb3rScDv+GK1/rYjmQ6k4sbiNqkU/jcOJusr0wc61NiXV59Wqe1HzctldU1X9bln
1gpr3MvnwJfPKbz7IANd/wlnhHna4s+ZyeMKRIWzUWblu6HmqhTUdGSzKte6WwIX
8MLqnk8vWedxDHAT5JpQQOkl5Eab7PMerh6G2nw7PP/4yIDmSd0kWX2XUinhn2u1
DEx+yDJPPpEngnw6stIONf7JI+MS9/+v+SQST6Yc26rmSJxjGh+bwuY+8fBUOYCr
eYWVOuUMuzb+eir09bRg/iZPxgL9r7ytzatnKw2TQdWpdxegCYl9c/wzFUvmnz5X
gW6ic6zL8hSCqkIQ6FqX/eKITN32ybCXoynTPROrTumkHqxpREAFi3Cy+HvpnAo+
Qnhr1rXGNi6RqwIZqGsEJPqOhtxqZVyTQXNEIwNtgiHNNhb11DKHI3O60sjg1B6k
leHeaXkVQSOAfCDPsg8E5YLfuTSmpSyMvcHMqa7zTzh/M5f/W4a8R2jrOal5SObq
Om1Rcck6ATTsFjC+avndZD0NE7jNn+5HMKR3HLWor6X1xM3DWO4u+ZeXi796xNsS
noXFK0vUmG5d1A0ZkCvddXThvKOUlj6HRpFuULJ3XYyJJdVFiqkJOZMJwQTAt1hV
nILl9ZfPxPFR2j6sJmm1Y9yZKhzgJBaa4UwSyStypqg1zElBpeEKuwi53yRRPZuO
+ehTc/3MJI3+T7ynjPZn8x+5TsF5GwX5uVYfEP8ZkhXjQc1rbnaqox0I0mmmz7YT
RFTGROBDnpur8gI/RTHIGfjQTMmcAYhfJNmQCY38i/RFSkurHCXv1fTf/UsB4Jzr
r2ygxZdMR2I17zbviCwgZJMEYVP0sbPcOK+gQ+JrcdsuPaiFIwYxDxR2cF4QnI6s
rKZBMDr4TrGcCktkaonRffwx0mYuEgG2Lo7vjsm5DjwfvPhdMBu/f6T4Ze7VAopu
absVtTV6xdSGJWOZv85hxvljU4iEQ2mEd8JXnpeObNDOj4//iSVftprT5POIdWik
whuF4u+IpGwXOLqBpaF5ilEUC3xqmGxEP31PNM4DJnZTBGTLNJ/QzoDYtjE5NDWA
QgDok2OzcEuyx+FnrnSwt7S9MQtuB846NC22fVI1YwMcbiULpPzmzbIDoNoJXOje
hCVYsaO/j3yjEiwNgeYN9o8pAmvrrdtv9vIDnxihpbAhHtc3jkzeKKHd11aPetyw
yGB7s5UGcVzP5CPny+cfJncFTyyXiUtAeVIxEi3BuofREz396LzCe30CfUgpZEOU
a01OLeQD/vfDVhSUiIehR19Ij/DGQn5wcfcKLl7eHdSoAb6F/xOjgwtdWLpR5mpe
VbpzwYwt790s9KkApihARDVY4Z8/54t0uBxiMjX5n8txCWXCTaj9TDYQBMg5zfyJ
VKp5tMCuIXy+oX+qrEFEfL1lE+fchb8FGE7RQIVDXsy86NQOer1vNYhqz94qovRe
gZJOHK0w1XieWTg942gtEvRaM2yE3LuBlN/ThnL+YGspNbQ7yQLI7xxqkyYiJoPW
phtLiLXMWYb70oVSTHxak510atf/pL9t/6I3K1FeUXIG+GySDOXwWnIZty84RpHK
HqGOxeZvIVhN4opPAVb79g8cFR0nHRDht0QdhUyI9OnurS4Itq8R/anaOdSfsK7d
2NAYStCCwVEGYBxc+kqZbhMM6xeqrCMxVwgnJB7v9/tilTWOzP1cJxdAiqN7YsRM
rmP7nwFfrC9GUFMce2g3FoCzITU19KjslHZv8YwTJDc4O2H70NxHLDv2LHttU4QG
tvS9Bjkfw3Z8iDybnahfz6anyhhPPlBuEg4iUBwacGCuP4kA12uLRtObgax19T2Q
L7M0R+C8Fyvb46lmApr7onl3bxCvRuWKgezUtDqA95EhlmwzEVzAdq3fADu7gyA+
PPLp3OoRej5Cua8qUHjKW0YndTK7lNeBB6ExcYcDMgpUhbx3cBtlBHZYl2N11qve
cTpbERMuVV+nrVnAh37+Nt9/ZIl/rc4LhQUwW4ldBamWdckwfVit5SrR2ZWPmmQq
thYKvfyPZ0W+dvBAtNRh7JXJI3UFdfkkJOBiVyXXaD/zrj6Mh/D0nS40b2vuA4Zo
90XUFlgnY99iACEWJJcxAxLle4WeiRqoMl+38bi+JeaFOxyz3JGKSN7jJkf7EbUj
92da7IubJ82xwmhsF8/9aqRrfU8KK6tq8BczN4BasVrpAdFVhL4xY9PIHlXy7dmT
eC7H/MtJleJD/XF+w0rkEYXypTXIYRgjlMheMy8WOZ7lpDxKHZyxbQj0hoNpVwQc
tyAtOYKVroQCwvVZyIhT+0+dQZo3HO5Up2ZK2decvugy5+r9BJO50+0PqF64UAJN
CTPEIDTvOf2fCdKxtdC5j/S9nV5hzX36Q6/LhNSNcbvuGdAS8xhUuK/u6jqG21k2
NJ4gH5pry8ZVqRe3uxvULl2GqcQfFEZICGm7jFFAKBpZwQOoqd2Si+ocyHMO/vVU
up/boH6IvtJuWkkLT9+8Yi/DlIpoWs5O8szk2z9KX+T7nHP7TAQLd/o3goG34WJC
qh2JNFCi4xZDNHeCHf8LSCjQHtsl99WS1VXWBmM6EM81oKakA2eDvX/U7jnsP9MC
msdbPDDjxLvgWjwjz1cSkt7Ya80FDFytwWAOJt9Prx63PxKESYK5UTJqj/G4NMzm
CVfPsky2MfVMY/1YcRNIdzFSMpyDSfNSnOJRFwS0YOTSORNswTSwvHvmnedM9feW
5HB6abDShA52Ur1rzBh69YnuIvGbXK6+KKTx5Y0eP5wXLc4l/TveQ1sFHqyqqMS1
TNsWmafwGHOY+BwfPqBXm6gsj9nWXa/Ra/e0qLZdnbl/HBMJ9tIV2zow1wkkTORe
CBbx4CwgTI+euVK1xpmonsYiTLg3IAccEAvqPpwzMnibn+wbLJ9DX8tXHrrh8CA/
LRoo3nr8KlzyxeM5AuRuv7Oo1IszrQO3Za+OiZCRebzxBsPXCBdW6SSbAv2O+sua
Lf9U1VlabuBjjqNU5vatT3C/vrnGIalhmF/DqHCYa01176ZaAbDcJaAr2qDoNJtp
ahM8ddOLjz4b2B6VJ6rXHhffaAUSa3CqewKwSa/RgC8JYfQI62Lc7U39DPX8NADx
73Hk+UTbdrKJteR9qiHuafrlNfy/9YCbjXCF4Qbdeo0FMmTxgMUeasV9duBqIXvt
MPbPnIgLPA6SFNHZo1UhvgSaEAENJha0wacHSECcJO8tVX2u1eijtwIu6cophZmx
vMyHBNOa+hPdw1cShPNQcW4dogd+MrhydQU8SyVrhEAc/IW5EI7I3BZJuZzAYZP0
b2nQDPM4QMGOcwbPQQGah6VkocXYmxJ42BdyTZ03iKT7dr/wikyb8ipNZQfGbRze
MEqbeh3DhnlTW2S9c5ACndQjwYMtiIiT/67Nm/PO/04Agpel5Z6XP/H384+M2DN/
zvsLC6zmx4tWqBtC6IuxANja+7mDvbmjuBll4wZotil/RDRFXhU98jpGeD1puIWz
U0x/rR+J5At4zTdS7cnJJSkT5ItZx+YXIkVo1hVDoZ+SIlPKaiCE4/bSJ/02lOeW
N4uljYXmhSmGIIYKligOWv9ebvfVG2w/L6yHng+WDzBdNV8Sx18pfEJ8It3HRz47
0HFUZ4QkAjbMdhrYCCGnkXbSS3wWd9fTejW7CHxf5CBctNK6T+XlEXUE7oXkRkJA
VRyBHvnGYxuhF6+DOxNzXuXcV5+1BGi3FxaRSyqdrKAVmlNvqAiWHcX6ZSN/iC8W
5EKVyCSVSObE3N9HgbbYt5ePZV1QW1OwXx57U9NnJaJpzXldYXfz4yz95kt7a3o+
58nbAhW8HBnSJAKaLknLUKUQVsslUAv8E/0Jkp1hbdtd3o4uxnKOoLyH9/dowZTp
GSZRMYcmGJewjd4exxe+7nmMJknbSlBL5+RQsNyIWg6QpLh+GO8+8T2ikYuczY/7
OJLzQqqS5Y/awQ3KUhiBBjbq6fkulR+iRnVFaUX2GxQ/m8VA9fMbtSwQYV9OI+Tx
LGlh4i5gWUSzmCAf9bYbNGWWqt0l9RBBeV6maOv3s1DUedmkpVi0boE9yHmZsill
zTt/z/m3AMh5XnmPHWxcmDu5m7r7T/BBEfJp5Nfjg4+5ChgfTG11MpRdX8kVZG9j
rJ/yGL04HIugMhoP7wTWvBWxiQ4eAS8jBe7lFHXgRxEXH3ffh1iezmB+6zFWJde3
Vh1bcHisPC373pXjg0BwVw35qqzqjyfntDj7y3GxmkNrI9Om7I1iPUwojdC9F9xU
GTeTXdMnxONFF9pWNJ+qsErUiGCUrLi79oKf9EegdRStk1X2dsDQNfL0MLWzvgkd
QAdFejiz0XtrCEv7CZ8fog7OELsbYROJ2ipL64xKuEaoKLBOqC9RokNQC3dPzXC1
Gx/GgABAQxu07sT/vQ82rV1TPEngQCKNMJk3Tw+ZHG9H7GFa8mejuXTy2kORQi4d
R0aTUvslrboPS+yacxQvzfMjwRdh4dd2yP53rajP3mBKnqviF7pk7w7WOXYuk+Vk
/+mZcrMNX47IlAkF6oMRRxo/SzUIy8auR3oIGyt/mujssnSqPgW1+PCiwIal24I9
XuEDw0vumP1o+pVVtxUeZVbUi4QAem6J31WH/nhza6lpa8srKZSOKDRda2/66clQ
J4PQapZVKy9npXJrel13r/6A06qpuUw8rdi5aI5PXrPg/LgHh6U7ZobKYKYxbyBZ
7TWVQSL49EcgvUjazyl/mhOI5cNnW1KbRJH1bA2BPcKl95Sth0bA0ppNxJv6hb5w
rf1KlqGz5N3YtO/+xGpfU9sJ081P5lZTy7XP1Pw1VC8nA8NBjgD2R0wSnLrlCB5W
eWo7M9fNDxdi+Frr6GuAP+XfbUPG7bR+vkmXd5Q7sZQJtqgY29txjqjv/bSYw2j0
mL+o+TWrvcIjl2kwH4WKoIA9wUrSyrNICSKHgZaFOpU55BWRZy5d1aZi0RKQJZ0x
r2rQrRq90kr7XhCRKX+M8wQ5Jbgzy7PiUTCQgCPxjXxO84hhFmbF+iUp/K6BTkzQ
3naPx6iLZvSN4rKCzHMLzDqFVbWNTkYEVwRC1D7IpRXFWxvTbVDZiDXqIRDbXmvQ
3VVqVsDBuPHCmuBlYfs3c5OF/z5BaCFgxsusrSvR1tCOMAqNqDD7DAFOPZP+7aqI
5SNjTPexQOPwj65HwtKM8fiWz9oCG8b6QuyCv2CTFnqiyFURSGyh2e7y/zxZFrNW
ADihuRvxf3eYFrUMzT7DlJcAJaOs8UZRX/qRo93AjS4FPHvISe63pml1n1n+yDR1
m7XyyC7bEW8s7AgOeduRFKDII93ef3l3MDnAebQpzxIV3vQ8U+hrCQSe6DiT0UEW
hfuYw2ijORyKAsWebRgOdZG5bUYafOFplUOqNQcypo6UzOKE2O5wds1ogp+I0oXP
soSj6OFMq1h8PNWHciO6JySoMKtD3i0G2iRruNjuxyRlh03qTYGXs8xlMtyFGQKC
rapBc/gO8W8N3YgPH2QMylC/n0SXwkcjFOi7Gwe0g/s2icq71KEahrAznoUPFr/n
ARn5Wz3o/WmFWwsXeH7WWQ8GD2bMzPDo4SZ0M7T3iIRbdgIWfXUwXmGiszF2hhDQ
L5q+l8XmXTEJvow+5IpCYuFKPmQfCqTaEwCB4/hElQ1tsx2zKTW+KF5arwIKaH/+
y/+eBKGs1LMfVYWsPak5HCUqAh3idOHMFSiJTXQuCBpFJS+D7+BRYjaq+fsXhvCO
XmI7baUckvSz66PkQucUtUAuACJ5beBXCpMU0MwRrBOugeLeXkbycorEbIH2avgr
JiLgaJP4Y8RXUQbInHVzmpAfacDaxK2BByGYFjERoJgROnEtEmhAirZuL4GPOxsQ
sSwwkt7LNlbbil6tZGqy8u+68FORYlKwER8HRWcOUpEkb1FAqFPmOE/BKO7bHDLP
z4AvwzQEDjs0IaLnhYQOI+Hb8Auf98fkC2Y/aKNifKObkpTGhYVaIF+U+Rb4dUAT
+TI8Wn1j3IxbQ5lrh7xya/MTr7LpJIfPF3QwrPW04D1vWGesfsRhUPr+qScttLQY
WFXBTDOaEWBQ8RKseqaejv1FPtPDDlQc5BtzwqkPfDkAU186plJySfrsoR7vbVqW
M0d9nmtYy3L0Q8e4pDI8HvhKhbWGQjTNsTjLrx87jWIuyRdQJG1cFAAdrpG//k3l
50axV7dqh2ZnQgnziGNavrsj7WceD8ShquguLVGEfbRRl/CGRuFsnGXHrDBV0UZQ
s49C5j4lgj9FbK/E6oCFbDuAW4qPGTO1XApUInZDCAr5pkvH4vQ7i8NJE+bCXeor
GlP3GaC/10VwAouahLu5VDnUwoWUWum9QZ4YkELwAXigqq+62Xj/SbihUnJvRJVJ
ZtOAjWDtj0+l0vfXTQFJsDObdfiRUrV176mYsjxM1RDI3qwwQsSMV4KqrkVX5OfO
5yjfOdo7i5ty8mAaCVULkV+eBs1qliGau3Kwr3sczka5Vx17C4UQKNKNuobOURPW
WxAKoOcXo2FlFKVCeq/kyBEVYMOVWu921aB/95kz9mvQMm6pstXMnK2QJa2SERAB
Ef+hw/7ejbKavKdh9pj7xATOdnr8vlf2FOjlKOe8g6T09BOlr5Swb9VKeeSUP+QB
+dNJE9LhNO6x4bCegvKz14Gu8CJQDHcrU7UzRUsKgvyX0LP+HzYtYqvS9/uuNI4+
sXQ2tHIb3reAp86lBluRyHbVswZ+wrlouAq6zG4BucoqlcbzT4JwTH+dmhxLvjYY
xsE/f3pQ+Qe/veLSN2MXRJJSbRi5jZkqg1nod+h95f6xvRTJauky1C+DkiVXif45
kDpYjceh36KV5kfVgCk0Dk7PhydVC6IppNECJw7jc3yq9gH+0dNzzkfY+kNziJyW
4If2Sx2w/1flKfpUuLCteS71qLx+u+q0n2qwZo/IA4VgSNCd4Oiun5Sq15Z6yjIE
qYMwMGJ8PXbPhygjdhXv1mil6ItSvns/Vp4eHEHW2FadD18zwgPHEhmByZbkZ8Zf
QdaFM63Rpx1HNQwdxDRNgQJBlj4IsLMr4z9ukLpELaXUjtgb82vFlP3gNKqddJcq
gAzHfiwEmEA5tTRhAu8M2ZoNbrEjRBK5uSQVJ3BOq2kNCl6R7Sb7s/yEWUEeMLRB
HARgQD2RXOCIkkC5nQptRCmjSOlAsQK34w0vPzF7nbiSeF5pwy4FaRDHwe2jSalN
4RqTUO4jxSjiS/yj2quqVANpgFuDWwTbMz+Oq9X47ORQnIaaqJiSsgjuu/YDpKYn
EQy7SzIF1/FqDpgCF/uQw4OjrU2L6fxv6SOhmv5q6DR17Iw2AujP/1aNoj7HcyK3
Ulw3UYe3cKw/I4DBSx44Ypck8n27Hpd5MH3fkvulCF8CuQh12Jt9amI+5byTvyLh
yVL5fO62ChDhQRMppaiQ2jRC0PlDNYnsl0z+dgtaBwty8OYELznieJuft1ZfHbLK
kt/9lZOwUUMbjD7I3kp7lduTgoZk86exi1Jd8E1kNeXWQiaq0zDEnva9ry1pNolG
dD41MccdYy/sTDfNOomH3pKzEL2R5We69osztKbwSg7cIKt5x7buZvpL210LIyO1
CniMdQcgKbQFTptnfJDO+71dbmS60Y2L74ejnE2BcuFe8CUydpm9ay1KO049WdsY
5QyorD5rKnFse0XeItfYg0pnsvoOuGNZ/+LJFEYhtN03PXiLz1PV2FmE+YAl14ti
s//bAL4pTcyM94164VLoKd4t7LHc8Fwo3/r6J/5fJLJolTw1ODbgXzBexrAyd4cg
XPv5KvWkcOnEnb3/N2erppmo//h2NbC+OhqEy6Lu3RWB0M1FE69zrgGeSPUb8lU0
l/SMgTTz0I7t3484/J9YvLvQ8O3geD//1kXyjNyLYMqtlLVtjyxJIUDleroZhiF4
3jE/bw0J9fvaHzLGsm5zQXmbAWw7unV0DTFQuraHTZz0OREbe7YVJxcGVtxpP6sB
O/OXlmzsXbKz3aKxSuHVXWcYKRcegEIzdH7ox+jHywMxXxhMrLJ+lIrhiHuvLy73
vCp8KaaivaszlMnm67wDs3I4ygQL6kY9aPhacbMAfZf4YFnf8TwfCHarU5Kpb2Cx
0DSWt4s1KbKmR4wJMEJsA22PxqF62sOE8sCRPhz1DJLl0GMWSuj81wM9c5GS1W6V
tTt5qiylBV5Gl0jXhjTeMJi66Tas4O0QLWyUMbK7jjyl7v83l284qMxJXGx9q1RJ
dw/lcv4XWDZj++lOYiQcaOuaZDUR2EIcdo3UQTB8E15PV7fLONgTPriubEEsovBt
vqlz+bSf/RdFuk9zM1gHDO+ZelDyEaQtepXR2j8Afw1MQeCqiAiaV33va5bn7OQt
0oZyXbgjRX3d3HtZHzLd2R1TqweTy7epfTYHSJmxjzFywbDvrIqaVdpYnv8l24Za
S/QHkh61GvnRNl0gP4t2auFe8886rWl/rhl7FG7rOlpaxNoGJ2eYQeXfKFL1nJOd
gRnHzXvmCiqSLlCAqC01vE42MAKev/SmzAg6RNd1/2vGgtygSPgC1q6P5UInBivq
A7dMefEJgaEJ+0R+HoNB3/nhQGjB9/fqdGExmMSIa71BjHYVXsTNhm3i1m8NrZ1L
c2DFcaE5In0cDIDu31Jxh7uDo07yvOUqWpd8DtIgXChNMU7FvThsoW45AeduyVF0
xLNAHuvJL/EM05l2pVItg0eF+f3QxkOajY4iKWTRW0VF0DiyNMmGYJujs8EmbQXR
8ksLWZjmQQYFnugKSsgZPDiEi4nfTyhMSjbtKarH1bDn9yQQUuE8WF3aYE6e/3Xg
ePBjDz0DuuY3MBni9Ovsz8sB2HuM+al1GBJICN0bC5ru9Z1por+denTKWv0og664
2zkM0fFfmVcCYzkhCixE0QxGhQcsyl+0Jgpqn+Myfc7pDzmX+LRkvmOoMlsjaGjR
iOb4GVdBw9ggdYdUOVVkXPYW2h/9zQJ5+eAtVUVTMlkGtKKxj5nptmXDCSXGLExE
6C7EF3v4JExjcrIQRAkJWAwIXp7mbdbMRPhVJ/HHouYhCWe+pZtqyoEM68TT0MSW
ApLBGTAzOq1vjIb2Y33Bc27wE1z0qf54lur44M7vdVgmW2dxReFBJq7/E2p9jzat
iPs0YLxSmEBnuuR96m3Z90Tki0wnoyKej+gry5SmD4uUTyG1kR2S6PyS5PiDIUs3
Jb5ZfwM9op8PXjVZ3BKTpd2h34KztvE3EusiDaKeLAnu5XRwFxxNOKRpLe5a8NLu
5rujjJj1uomtKaXRK7LCX/8zhbXsY8NUHRpiWEIKPUTqe1Q2WYBvW9Zzp7rqzmu9
62l9KlDzKwQGwTJ5TyvCYvlWCsm0G4WJUlh1CBkKb+p5WXAt7zU6aYPpVDEhP95w
vZiBnPbQSKjQt4fJmLCPUHioV6qyHvKVemVClVPZ/WbJg7Ug5NAv56+BdSyKcazB
9PSr76q4sK1eQDL00SglRgA/k4VcrJEFDDa6A6vx4BUyZ/m9WDUDxQ8kiLtbFFIb
2b2CwH1OkRmx5zRBrRQJkEmb0Ifi19qzT3kGsTM2BxcWj+JWeiGMvLWbSU7Z95sh
vdbL5aGRkLLJ38eahs7Y7ocmFL8lunYJQDhX89rFulSu23C2jm3Q5mFAlQnuiX49
xZYl9ABPJiOwTfd2eY1l/YZd/yqe/UYNqb8rl2Bj0bAoIL7xB69UIECMFIpbLc6x
sLDqK3Tv8TqCXL4vFLwQIRz2W0Twr3UR+767CcldP6onxjuF7gTuaM6Os5qdISx7
uAf187SCfEILzry7YF7kSTkbZzEOf9n+57i8T3oUKwPGQPuWYC4xX1uVbSWoGaPC
1c1S4YjSOdTm5PF/bXrKSkNeerbRpGk9qmH8wNbghqg8+CRbecAIWYHSh+0d7+9y
dIjIt6w9yGmrKe4CF7+QgxmLqnt7Nhg/egWvItgTYzGwdtvYhO+tqt6M7A72n6eB
Rtrl+DSiQFJkP+QWylKueZGlnpoZtK8XyRKKuHVbunb7fzfbDB1AXR/OtENPc+qk
V9SJRZK1sFDuzEx/a2vnBvkkwosBlgUe1oXuhSm8XN8pLpeUfFhjhfXRyH7jcFHC
8bYWtbIHkZcDn2YInkZxzWFaY/93NMH2Un5tLxCa4wzIWeVIkD5FXqJSV+2Bvt8Q
0+sV0CouPX/EFjSEfSM6kn4xTEOSRVqrJwdnHhC/kfZZb8+JyrQZFVfAd04ivDop
ez8+IssoBSod3snL5MYxq3iOaw8c6ZdLM+bwAYQsZ5pAOvZO3wYhtst7rmPxtnAi
VAQbs17VKO93Szy3eRUcYFA+HuNQXjuQaFBALq/epkNJjH445wHhUwb+UDe1G9qz
rNMnqJyu3o6J794jntki2xGo0bILWv4MMQYjmmZpf5HaZ/7/EcU5BD+2IMLe4NYq
WFD9L9QczrCwmFWVHryo3H3LjwLAhgGeM/F9M2Lok8HCetmSfXBzf7zDBeu3hrv/
l+XRMhsTEOgFvoJwVIxoX36ApXXu/5Hq8EshRDBLKVYvIW7pqS50tLLulg7n94R+
oOFfFRVu4k7M0AanYBK5NRabv5ussU8yOIAnmkjAN4ts3Z20jkNoVmSGwa3hqqBf
ilk7+tlyf2BcYTyQP9oOduuZqXnPFFoxw4r7DAkhkhwG2ql/rMHapUmH4MT/fSc6
o5fdpmtxYJT0RzICMNWnVMmHyDo7baAeoZwjk1aqh0V8zsRc1rLvWoacYhi8Oxg1
9v21QvZ/v4x6haIHYu6C5L1kY7cLCNkncXhmykhofu8mA2UzsAB5FbCo/CIVYkJp
i9ljJ3+VtyNVshVbh6IRUpCMxfwArfY7YWQL5DMg+UO/aPF0MoVEU62rnoqLFjTn
ENWLWQua2oXxkI3Z1eCOlu4dpJ44oA/Lxls2LwL7yp40+gRyA8OHcQpjyU7b6/ff
y+PmAGYwaakRJB4SUTbQkkE/mQ0j3ENE7drU1njZbtEetstbfPDKO88cID6yOJMi
Od96HNHEJL3Hpac73nlUYBHOnw01iUhgiY1pi66t64Mo7wR2dR0MwYLjvgrf0ZNc
R1UUQCDh6dvAmfNHaoGs8g4eeJDqcChXiUTsRpZDH6bAUjvgWnKV0a9baKe6XfIG
/ao6QXuQvsA5L0a/GYEtelUwgqsePvXKUU+OR6Rz791H81Byg1TPtAuUXm4nC8pc
21TDEWV0aAS4AXwzabx2dBoohc46QANwrGM9l1DA7y5EQtBL92gVG/d3JH+gcc83
kDAsQtFuNWdPyr8WjNmfc0srOArheppJoCEFg9FUrXgsDvmD87juOw6UvvYO+P7y
4qYQj9TwWHBXV82j+Yj/brUgEsvxA+uaaTFHGWxW7nHbwpetvK+XeEWqsL4YWvxy
TadRvYv20gCM8UAyWRqYbkWX2waVNy6SZyFnKZE7VIn1L841G7Zu8YnUDKMHQOGt
InZyaiKVrkr9HAhN98Pwx+VIw1KwCE/8tzAvLMgH76AuZs/OuKu7iLny+P5/mjyl
QcC5Eqr4qYh71aY6h9xrtXJ4vduDDYms9g9KmchvQ36Rl+hPWaKszliU0aOGYeHE
UNbMC6N4O7ojLqriDjKwjcgjnmXTpGffq3quoBMOJzJZGpWXXRUJKS0hg4GbOnWw
QeVT523EVXM7Rc3b9hbEHpsFtlLWr+Ql69yRwNY0DpnaYUr5rlAGEjkTrP7zf6Ou
+9gLasZoU1oM7gs+r0Rg4+23gKWPvrPesWr75if14lfQOYeEzMK5pqjA9k988TmO
v2Yx+ev5u/ZI2vRZq7KaKICJ0Y/QjnmglBAnUpVL00d2IdYaGQw4OiuoMYsEqj1p
Uda9rQZULWOIpb8XHLzC/Ehsj3EfYXMUsmsq1rF2gwNxLi8ZTLZlNRZt7xCBPtwl
NgY83y7b/v8hMfp8k4/aNAk7EAFPiBoZZFaG/ova7H0lyxEtbHazhlMeyPOFV15Z
M4sMeBq0DCX8G7rNlF/PPiWknskU/KMLsZyRusvG+X6MmFUmd5Fyu08gDxJEeQ/U
IalMfZ3DnZQIyAsSbmI1GO4GZbm2t/8xJwH7p+2CiUFf6MYVqZZp7azH4AXPfRHr
mfAmba3TYYsVrIqtE84xBYQCTPx9yflXLOeHprYO0BAa85y5o+tvtMDVBvpzXrXw
Bkj21hHsikGnnNBxhbnvxU0JC0CsGRifQrZbkERZcsS49I9SZ4KNvCPn3JQ+rc72
fpeZTxS9wYyEGpRHpb0Qlf76KcDvZCSL+V1QVPYrehYisxt9tRPa06brPCR9cz0V
LBl2kq6xGTdcuXx8H8On8Sb1ltFxmtmwD2bb181TYc1annn6Kw7FnygJfaACgehI
JKVAKBKC0YBPdCMRho8ioX/LjlxV/LO5Npn01G6YxrO86OWNwS0G6Y4gLyggLSZI
FhUlOFKIwaDmabgnRzIhUsMNRxosljfQ+ESgg9ZL+oTFq31S/96ocFixRzB9SXv7
+KutW9n9RW1iYizfwsJ4ii3o0I8reylzei50f0h1YLOeyDiEUDqZYhu4OKLyjIN8
whu2SqHat+2tzVv/QXYoQMVCY23OV42N1PH++SeWNSfWmsGa1hmhRi/XaP932pMC
5bM/Fk0T3kZq+Hr27rI4px20stQh1cvm/U/t216doMMXNAO7QEOtlFZIfwxHw0pM
JHktgmmn8Ov6g22A2kfjp5lfNU6CF2IgEnMmwLpLWeqOeypezNaeuhcxFcZlaFyg
0OH8xYwInkX2EKKr4lVAPTnU2s9sHU0WrOqqD2SvMVJ1QoVTsK5I9NIpNklL7Fmt
VtUidLUuvhTgYmU1ezcjQjfjn8MpN6+O5uLHsRh2ZAEc20/eNeB2II8wuQZfQuto
twAeEB0F+MQMv4rSynSO+mVrmS725wb/aD6fI9Nf7OXrchhWgIKXnwvlf110UCkx
oHKVzptBPq7S/7hagGSnUkTSfqFOSM92KoExBzzoec2jRkn4dstrGnID3lhn1wer
rMItfeAhSrYeiWDrWQEnIi2VzWAyXXP2l3L1/L9zYqex6/NSzMHYgMjz1UVMHURv
dFNzgVXqpPvgJJuh5OixHsh4TAXToqjjUAgKgYO9UGM6uEZGrxZcfJHAt+gFyOGr
6V+/vH7VIcXQnh6ZZ9P//hXFxrtO2mjLNtvjPQejWfcFDklqoodlNkegf4M5iw22
Kyz+6btI1jWTUF72ChgQ/IlXZu7U5fzMqUIRqe+BKkAWucAYCw5aT4a+C7bTggq0
zGrPKXwtyLWnjGRR1jUdcbTIQFFzDHtJNheU/fxUqrBf4eVL5IBWP6YAASQM7+NQ
JDzZ0U10VvhqIf+49N9yNzvtAVRbO3f6rjn+YuIMmpBEvo/IRl7g5NjcsEuY5bCw
GS9dX151Bjf7rfVd2srwy17avj5GNF+mZzkfi6jKeER4jk7DJpRlKdhTshI2E8EO
Hi7fLUUga/RrfhqXUZAf5ErJYK8DOnlCl2NjnIxckPLSVtudh7UTCCI2acmWTwze
4eTI7bJzmadfnX3zwI8xUEmLC6/uV/Bc4Y8sLEJZ9jsZQ1/EOEx1OxwYoyAMdH7l
FDBuazA5Uy8ETiVOGkTX45HRu/1WhezAxzwsmIox2Fz7/TVV3EyTs31FtbaU9/Ji
xGeSKs/Oyaoyqbivm8B1CBfbXttMxrfuFhPXnBpIt4MoZXdAqxmd2yZaDlq9aiIL
52/x5qnGJDU5hSFr5/q5ub6scZVhXi6yrj6mTisXrOYeD7FMh3+7SKqsANg8Zpiv
I2QWdRUpstwREYUQykhtmBiE7GT5jHqIMKb5NpLhKTDXu4zw5oBMYO60z+jHf9X2
TcTU2xjo6Ks/X88KE5H85uIgBdppDepCEVYTByLFKf1g8SgV8SqdA7rgp0WAZGhV
Y3PTUyHrdJJLpCRXgyAJVd1p0OXvyuFO0u/VSjBuArrqIzHDhx7WnwQpijrbjwRY
psUAxUduYqVbZdOC+kiKCLq2icuHjEK2GvQeA93GrauarU7SnsOmM76vHi0A0BpW
BAP3BUUnMF7R9k03IM6hEF/RZ1pbDH9NH6cz8bp/hsLqpQWqN63VU9M01L3MWcSX
H6R+Nebk+s5DbDP0dKcJp4XvYgcHDD0JmNkUJ1t0GDXVjSifxJ1QKgRcUb6Nswvh
+zO+CqQlmsSGpKB/N8u8HH9cLw56l2MAJc6t7yPqWqIJQ5/1exEB35M+yVZEP6Yl
4Y3/oExe2+Gm+fGXWP3IudUYR5+O47diMwu8Kbek4woZLJIce0XHoiy3l/CSz8Zx
+hMYA+n/YZJ2MgzYUM5+sQSkjP6CR0HzcSng8dWcBv92PIgw/ZsHYptLx1Xa34Fx
6AUjPFOi7c0KDpkI8SHx8ns7FkJ4ZV149JbcbY1wCC4+hbUVkjtq9afR0t251UBY
B4PEI1GMWRk2uv0vO8jWNDz91jcg1OmwBrNXHfgOtvBLkNdPbiiCPqHinx6CYQfz
LleDtgdE7P34U5QlSjXd6XwzuboVrwI6Qu8IuahM00FdlPuhPWOiqvlQO9YUsw5J
eQISbdoYcyci1WAiDWg2Q8VBwOUM32QGs8lWnQFt4IMi5hQlv1fUA+2t2Tg6PE35
hXqGkjR8WJ4Mf8oLFPqKoSpsflmIa16tFo5b85t5lNM+SAkEFmn5KkjUPuSt5b1A
0bH+kgYzbPNmnEZYsWif8EDl33LOees/uFk4s776B1dEWYbtkC5UNgcQtNABIqCM
YOroCddSAYfziNS8fEjT54ZnRVrEBqJOcM2CrPVXk5+1x21l3R3iblm93/ouQz5d
uovzmlYH5yTyRkESgfoHCOEPJbD03G1gbe/6azrLetZEA2n+xIs0Zf68r0qGQvZB
j2sQ4N1SV8kHkBnpJPm6+wW599DsnWGgV1Nq9L1ZUwo33SeW2d1NxkTigy96MPgk
r0m1hZ5Qx6J7Q/EidQ4MVUyW+m77ceTiBEsOYeDjiKJGeoXwsiTx4msl4KIEl6r+
2WDR6L9rIP46JSa2pNRSGgBtyhNB5QgcMv2lbuadbbiFtFWrqTXZjtKf4yDL8wuj
Bn7yHtJ+0YCiBUqjADydj5khBnpiTGm16OLNEXG3DtguVCPg0TAo84pjyzJsJYha
Nv1lHj80sCIzqH9sKzrGSUDOxcETIgIGLI1dHlqDMD8FREfUDIIRV07ftohIxE5X
u9jipQ4Rihwx/P2a1ClWFjk8eO4I2yxImKnfHPOcPW3dZni8Zfy8xtSwLqZEtCua
+1IgE6bEEwImKIplJw/Y5Jp3qRanBKITn8tCkgvEFFQwtftSBK7rMtOt4WhHwMY2
9RK7bPaozOf3EC11zn18Op6TNeKoox374ZIWe/SyqQ2kozUPiPoSknDtV4/PRMW0
TDKFa4eu3XaYkbDJ9XdzzOblsoBlG8H9SYxhTwhggLAH4Vv9c0B+5GkxjZlcLXbb
5MopJD1gkGI9BqiicG6i9AgLtUma5BEt/JsA/RQItL5nGvSNYLcYKmA8HymQT7JR
8h4/kNdl4lBw1fPhNoXf/9YhCSlps1s/fg1ZJ5G1YMsSIc0/UrUuyS7DoNkKPJsP
64fMolBZr/rTef6oGBj9BFseY7B7ga25b4P/LW8fQQa6+1cFn/tAErc3IqxqAX1Y
wlMeG0/1y1WLWubZ8JpnZWlGaXhPFGWC2qa0P/OIuCnNo0ZoxAQJMpjs8MBx7R1K
DV5T8whpk3sDZGbnfxfNi2Evvxdi0Yalhc2Bfr5hcTqdTIIDodCnpCfU+tg0dULV
80ATKglTYstbpzTNLOBY3z8HJIcWhP/bE1McJ39w73avkk1dAbcyb6JSHFILhGAW
1u/MS3+/fQkMEtu/JK9xjrNr9S3tbzn1v8dCpoKwCGDQ2GhV6yKdhsC8xG6wIUEh
KSmpu4w75YLywFS7xCqgQVbnL5tuEmaqYt/nJvkQ6ZVLbhh+YO3qsR0MSj1AQXOD
w4V17+lWKgUexvkXhIfYABD1kUKcil5uhUdKkdzWzY92O9/mIT8Xth3LGyD/ahVD
f+FiSz887UlpoHyOlOKdqTqmEc4hVrI9zRGtWHoqVI6cqljvZXvL7MD3U/eAVLOX
JAZmkRgDQa1ZiMSxwWvWOHJzheAIlj2GF60KXIS1Z6mVzWWb4TMWSkEI5D2S4D2P
T7TB3IlpS8fvbhW/mSFVRAts0FeFh/d9EQm8bL5nxuGLgH6dOW8JjyTyUb3zLr2l
YPXaEhnHp1vjRJcOve3aePePtrSP8j5OCyvAxXu/0BzGoxW008G79PzE/QGvautS
nOiZq8MA3ooy65Te54crztZPPqRz10m8VyfcOi09CKRuiUsEx7k/KP+UwMNIfhBI
weJ6QnXFKV8JNloZjoV8kNUKkl4aDnshDQN/ru/1w6cfcNldEyMmrtlIJFJWvfup
94MhBzrOEbsdjzr9MNQsQWa+zByv6LOjl9oEZbpKbmtCX+Pnqp6z5m0Kp1yOvBWt
zU1CQhPt8NJoyuy0oR1SayZ2/zwdukD/WTkEDcG27UjVJd8wbzOaj+11kltMtCOX
x+gZnuxbT77LL5EuNwQs6ZYEu9QsR7C+5+wBskUzwnHmsXRcfDZq9o8Xjov0Dbd6
C9bD5aQeRIETmvtjAcIMFOM4efpwFgjYo/5dDsiWxJHjGkd7LBXdunU28BFyTDrP
rlSdyEwj68VtFFHBdkQdZk6ETeFRFaoS5XXh0pmW4q3+c5NgLQnKD4LJlVvsunHP
9SFqQ0vnSa3Iw5LsVM4MQESYytJFISIs8H3IPaIQfVpCNuVd/1K8vQgmpLeT2hvG
lu5B6QhXhCnJrQSSHzLNAgRwlZv1yIpSFTGTdlmqKswCNV6vEr4h9EcRC1zfdkSM
TpU4L3pYYu3XEBLISO0amdLNLo/M4Nu1UihOC9p5dqxI1XG9Cfc2Sr7L4lv0rt2W
hiMrtGywma+BrBVfZ751K5X8/gmbg8Mc2Hw3N+HoN6dXRNEIFDDHaCrjPSBBTW6F
V+B8IcrO3PleIFRohwN/vnjgtkCl3K0KW2O6HYt0N85BTHggqQ+0RnRphkgL4mQI
hfIldja4+QaBigNpPaPLUJ81wfI33K5jnR349u+B7AdrUZBHctcLgV9oBENlf+pm
susFTgELiQu+ekG11PTEJ217R+oi0c3pZvqdrbYpub8m3JryetxWkJt4WPzPJGPi
mtLrS2Xyi3zAfoFKkw/MSz3rRq4Oxgc0iEq9+0W0FUACPWubj/fbWgxOV2sEyD6R
eRoUX0c9QuLVutOn7U3iIbiXkbYDisUqsipnC0n6xUefJiX9kp2LmgbF2nu2bANW
Q27c5vplMj/RUPtNTY0Ib1Utj15KK/aZbLTG6Z84YSFdnxpbXTZ0GWnMp11/WC3+
NxPfL0F6+QP3FvKiQVpYb6NTwQ4fLfVekQAM+z5vocqyWA2T0EbNsa2Vpqae1DIu
fnFyD6xnQ272coyQkVQztSlxk5KbeiiCcxVIqpN/21AANgfgR/VeSQdyr0CDdr+Z
2UKyzoUTg10iez26Z3U42amj7pUxEkY5lBwt3lVw4wmUOGLm/5QuFuUEkcIC8U/L
zdsb5LTZrGZql6B4yzV43mM+GkFFxUd6Sd8xI4eEldvRrg8zyXTOWZbB7Hqo9SHC
ZD7WARIjMqbcXt02k0LBwjlvEfauYyk0j/iPtMnmRTy9SKqdoi2CWPyKm9rCOA1w
QS4oXUkTci0ItWWX8hqAExWtqwrvMnB2k+yIwE0nMsw3N4fgHAMqcMt07P4oyYyh
zVnzkdJ+7bSyKf+OvO6wvR3RmUbyv9ZtF42uHzmcVnoDSq9Ry2dq31pPn+hHWmTj
HZBCoSLzripj0BmzrxODBGitDe1vHNvg7qgdWt9A5V6SJEijffWm+bs37heTqPV0
wBV5/RRKf1nH9bIGBfA5hXih/y76bRR5l6pwdhMQRCKZqcvKlDUrdp4CY4j9c92z
XwtPmP1u40fClExmyHooAbuFrtqRFK7oFGbyI4QUXMneXv9rtJgl2PVza+rl79xi
/b4mS3kVC1qoJy4zXugSHrQNw70KUHxBEVs03WGzOqJ/Ms83CmhnnBunlfkqO1N8
Lrx9Hv4bGymHsF3zamB88jy3Oxba6jCxx7uHlA1MdXu55+o4KxBdPZm+0hEyHvK2
zGKVG6eC7efZ2nFRaCg3qOP9zB83O3jkSjMu18h0S7FNK+uwYeImwiiNtzBa4Fyj
DNSnqmaSfeUeHSUyHRouZUqvlKCPrJ6BwzG0Is81Vi4Z92QOVCE4kBy+LSw8PhUB
WiPKHNGUIdmsMWCG4oS1fLq3jvXxEZx3sosjkSLrSWjA/Mou81uqEr9SJc+9b3cg
d4fOFxkl1nkmGT4mqcoenP+lAS3C//GG2348Ip6K2n9gEcUzb0iI3hjBDxJ19x8m
3Q3FYx16ev7016vUfewOWH8S1gvYsQ4kVH2gNZr8oOMSI1NMqLi+4t18dhCeii31
/fEU3HU6jqT3A6T2oZDE11GTYdLdPNIdRGfUbxljkrg0HO0+caOdkJ0tou8OTZcS
dMSsQSMdiR3cpzbPMt2QJ3/ZpJijCq4zdlJG93t+Ou2WRUAkpjKthC7foaveC24l
p66xJwy7R6CgQXCxj1Yd4NVGjfvmDWjHDQq5fToLKU8wxHWE/s+nsGSTgKq7X/1R
vIYeAwrM6HEKcf4Fc8woIivQfXWYVhOHtSg5pfqr/jpSZcSZ+lkUIz91UBl65xu2
X43S8G2ynh+S1eS/T/lByOGBwV9bPOv/QoTuYlw4TgY4MezeSLzKuBJSFTb+ojRl
XFocnQfplFBBMWQyS816g2IvWJB2Jc1qxQN3VyEnyBple9q3vTP4fdvAalnJq3ZE
invnFcn6+0DGi3PwnODWmQTNEgFQZ18LzKurbNocteFrj34C2IGBvKp0ES8kCgDj
juRcA9pCNegW6vHA1waOP7tHv9ebtOvScCzvfVyA8CuOIJNeyg/+fV42mkWcjiKD
fHixD++/CwSqhTZrnw2dEyo54skarW9i71SNM7L1j2Ks0msXiYWL5dZCS3X6JWBY
of2suQxnWvGAwcNmfP3nezdy8uKdxO3mK+RUgkWlE9h4Kcu1q+WKk0tXH5ii4s+/
7whRcd+AzYHOA/Pcfv0Ublj7/KbqtKNKb1cg7SC36BXcuXE2O0hx857z1Y1ES//N
p2XlRkYUrZ3ITPhPg2Z6YdVUJ+CjGlPMMJhUFvqR0967Uks55norzTyHarmSO/9V
tEdfWMIXXflt+WdQaRkMOR0IAZVg1weJE3Yzm86tNOYAKjUktQXejDTrMT7yTr5P
lGCo8PPoz/DHCWPdhMEF7b3XlnMDMP9NopKFqik3Z2hERpJqj33QAl1wJ6rJO1vK
NE8DvDy6a38Ac5My4cbUk3uEmJeynL+2diifTUyLXW9bdkuu3qkyRtdTaTpy+T7z
ZKeU5sEZYYS1nxkJNBG39t5mn7zy0yUUhLZJ4mlSkSlUBJZpmBo0XgyoTrrZGWPF
QNab63SQjCnaMe+O05c9pv8XZScwkS+42CrQYYj5h6G3VzFOGGv3gnfWonQVyPXe
eKo3e4DtNRmH5iGkLkqQfmKFsfg0RVJi9pSxdsyCDcqRjds+0PZ6REHtLdgfxbXK
5lelJrbvseYxZGocfK6T8/myoYrLoLmGylVrNmfwfIschSABh8WpKQ8Vn+bawahb
i1zcLD+LyYjtobZix1nn0G1aTg/Jboa0t/qhJujdNWRbk7BXrSSVmqvQMNWHyiyo
HXZMsDpJh/dMsGjLUvRJqtOacGoMZEpmbLyHUplnC/OA8pOkm6j9ZlXMv1K/ZJHg
cLTNz9UxgE5MgTYKM2yKSe9LMS1SYS2Mtb6AP2RTDxCQud0ae4hqNAbBB9pjPqZd
5g8UfYwlGqYaA7OUKrCelZtZW6xCZ4pEQ9bIWEnhP8CCLvUer3ag3L9vL9UhNR/8
vGM4f5u1U+tcArLE8an9vlNJcAf1T9KwVdkfJsA0FcmDJD/OA9olIU1E2L9uw0Gk
PIelrOv379OZRlL0f70ESJCkpq6rs6ZlNmDQoi0xL1XweJoGkyq/B4v6eLyus61f
NUDTAaQhrAbNSDNCWr5Z+hzejG1Cb9bUX0w40wZ2sUixd9g5TjB8y0FIqa1eniPZ
HbxGkCBn2kxBn9uXT++THHrLcz39EuseanFYdzEtFpHxzb2INn8xK/EnbCBSblZq
u5uUNh5HKRsY1gBssCXqeJnClFmMzA5OXFUla1WPEiNs0AQKbDvu0jf8OZedsdsq
mac9NUxhVzrqdV9wyRh2aQfVI35AxWDoH23OQImtV8RODbdLc5lMI13RRdxbcTF+
9RURxZZ5yoZMLJk+N3D0CtMDIo9/C4SGqGEJ2TkspYROLIQGIAOh3bx8FIFg7Kz7
wSPLpQZVMqMtzj0OEXh0uy6fX+sskm6lJvJcusSuqa0gmjUZbcMy4K4STMobi3X8
hIfdbdgOJ4RMVDy0Ipeqfz+NBfVqVnwGjDh4u5F4M7LT6XqQKo8w60Q2AWhmo3o5
uYHZAm6vAQ0wA0OrRcB0WRWBJg4joIP99zc0go2xPv2HE29at4V9M5A4A/B+g5sg
v4awwN/O2o2sXFALNo6Zahn0EstWI4tijZ7V6l1fDwsqNI4Uw4ukOh5zqrQoCwPm
bPj8QeUi5OpYNtF8n71sDgWg79udtyOXjlXPitd92iD3lIVKL3YSCLY6scILe1uE
F0LmS2mreSKtNZEnGRqVIMx5ZZcOqXVSHttrdTLnUfACn0gszNDUUevxvIns2WHA
qUYRWdC/LbKYCODETTndesaOR1hiEBRcTJXznqGhhjocvnZDBYLAe+dbF91X7585
mWlB3cfXIqg73m3BQPtYZIkuE71vYenBsVpQw3Z+iorI/sHc8tFPFEoNwl6340iC
I8QLB3h7ldFh64Jf3uLw7hnO+iCgSe0S71E+NAHE2uLg7AhYTT8NKEadUGvVO3mE
U+X5DiWoOaIdnBL+9cq9z96kdozpXYxfXZkzPOKHlx6fymWJwwPx3sLFdqoIGf7V
bQcOUJXM++EWxl9pa8UwAaQXdrEJXeJVKqpuIralzm8X+2Bb/I00l+KrH/QwG0mj
lKNTZgdzwsXQtmMrRAqov/WLZVgYmdPjCWmCNkHUd6R5ZiSaTk0RT7R20ZQCQVRV
Ja7hJsYdJhQmL9sXbAriesnrm6yb9QpGAMCaW46Mw5hP4K7VJNBiEVMxvTysJq2+
y/RiUPn/RGopktfaAZQgslIcNkEfeTOfRcIeMhjlk556THYgGfglaouYxSgX+dpi
RQeFj+K/ECArcuWWL/25rvfumMOCQ+gvY3MPc2nM6jJD2GviFNS3ug1vZVs+dLWa
vUfDOnaOd2u7AqPEImFeQ999iKhUvRv8kdNbL0FRBixxrb3kb41PIJl2zgr5cplR
zueQiRF0qm6cAu6ubRCqQsjTO0PJ9g0X2MWjNmqDTzEKGlA0/ze9DEuujLhc2wi8
vaVUZKriCm1XjIgZ7TK7t0flivlLUuFZLzh3fYTaaka/TZYgY/6aFT/Clo4iDy06
rH83yH1i9HLOMnzBtMEXGRhYJua2H29n/7uxu/Mmf+/amTjQCOaFWW7FzihfdCas
dOGrcjrw/HegJLx5xXZs7OmYnmdmxYLW23ujkgIgzlR+bohVKTom1mzL3DN6GkI2
AGpwpdM0tX0PghSGg9fWdbmJouRbjLGvpsl0eSoFBZOIqT6r5tdJOzrLnDV/diMM
fb+6V8uSfi3xsgU3q6tsrU8oIYbPhqLXZ+MNTMjXLznNZDm56SMQJb2cWFx+CsKw
sejgWCJK4Ln/gCFMmoYoi/wce3IWrKvYi1VEbQ6lODrntvI1JKPnD6ZptrXliphL
Z7l/YBNWoWg/DLmS6VE3lbL/YuvX6Vuqf8+DooDrDZrg0ikZvMcBHm5tXpQ1j5ge
pcJVlbpJDqBk8EY4z7cTkbb0w/n3TlBaW4DI+cgRgzzt0+qjpcpli6glUoDyuKdf
NzELqspHoc1Dp3sHK8gGt0YJBNkf/aRge++zglGwkClsXbezgq6CIjWa3ddaTK+Q
MODZeygGwNmYsBKWCRJMbEKCuz8PT+L9+yjQWZLYhY8vVaRpqMDLQbkVlA0nunuj
IjF07nHROvI2TBhvn4Seg1HYey5amPFx7uWfTK3fs8sU5ffyIJAZCp1uqweStwMO
JOUJh9VS2Ha94qEtJjAWyi4jCCeewS3CDWdy2DIR12oKIOs8AGCquZoDpivXwSLN
T7FWx7jM5ZUO6PkajGU15Jbh8RiRFmh0W6bHjcF+34ug5yJWMlLtK2XWqnQW5hbz
y0D8lHxNfQjn3scL9vSDxPpMEqO+3rLdXyTjJWgu/vZyUqz4mIWEl2rKzQWBXN+P
Qn474+7e18HChy3sEyPPoEN0FVJEukkjVUBHmnHkBfbtEvaEYP/s/GteC3gjL45z
slwjxxUKHhY9qxG/DwtlY1odiN6tkLmvZfG1oroZgk2UGFr43kFHKRU0Y8ncdlkc
uR9VK1pHhYPIf/5QruNdiRoZ5P4jXUSBDpl6IpYZ5Xhvt1Q05NCwMBNEmz7ytb2k
Su6Bqbs/uVoNCwxHW7O+U1MoNh/FTr57kftbw9HhyQFeixfS9f84KDhvC609DYDU
C/MMO4yVjoJCWs9qQjRZhpBwpnbFwrtyk9Q2ndJtfoCTJnPCPLejyC62tRV3cQHA
d9wRYU6/pmiy0H2ixxCcSuNldj1LlkZt2r6e1NWeVXBEf/DcuTw5fvKgXVUMff4d
mnx3pLhWht+MtkZMZAq2I0EP3Mw/73GS3H9yXY+nxx58742c2VDRHEK9W6TKz2zt
nC7FEjshtvx9Lorl7MRHXxt4Kfp0gAozqxSsyfNifo9s+RY++p9HDeiQKy+l8E28
9dFBrCGCmimmBHu6xbZZjxjY0sdmfCvYpoefv/btAcXu3RUERg6g8f0tF2ZoUsu/
5QoCv3MvTSgBs63CKq7XKEtEHoXXMkRW3NdXTcALs1kSmHedit5ttp95oMvLz0J8
RSOGtKIGjOWVpyyz/SmAsMlNP+eBVqzpthqvJJJerFf3K7YWZsPwBZsn4y6df0Ag
sjVlbUt1cYDJA2G0eZT7CvqaGOe/cBp2F49SF7CSNoVKM5YbvZASM1g2kUE7B2i4
gXNRNYanxvgtQ2BN60gJDEULO7Me3+qBE0zy2chSrj6HDU7fvw5ptb7LEI2eZS3C
XKSFrTehuYUQnEw3joOXQDYNvf2DqqCULuAsMFqYRUhPT5Kyq4U1TbVN30627M1M
JoItXQMmm3IQ75r5RpUJ6Z3nqHkmUZzsqMYHOIpRFFA9Mcxa9YqKnMzyg8hDQKkK
iKaf5w01XJZbMFISWt2XWUsTtXydjITx456xgO3Zu/1GicbCyhGv+PFX4elV5sQf
BsMAkaQZzFgXXOpT1SW8mK0F8A/9R08htOS0knnQk+N9Iv78M96rDC9pXqgq5QGt
jb7zqBpieWzWJWEKFVj1I6fjEcfsSmnANt0fwGwf6J6IUsopEOU5pGmgZB8fCZdx
s5Le3fYuMGZcrolp3UuUtD67wEMXfzMFg8EisN5COTR5DROJSoCX5+qrIDieA5Mr
xPxRdmRuZ6zed1JDWfl7f/ARHxeFicgfHOhpC5NnKSVDB+D5TVj2DNoztrl67uaN
pi+ES7fNR7U8mQdp4mG5EhxCEbgnqtMn1ani8KdEoCGLf2yLTYkfyvdjTJb3Fvpv
0yxJw5qwlv6TeFejB/kb4sheesdlzJUe3t4TsOCr55mhRX7Wal7zwDvd5C09GW+O
JVhEYux6CkCQoClHVBrA0Q6rzzggBctOW/DFCuFljM6TGLz36Vf31M3ZHHQN7qGt
DVNfdTP5M96Ftow3BQaI95K2iuGwGHvzxohOxZGkJwe+tfbr0AO9r6+Er4pkLZsr
b7Wd+ukJaW3ZaCytXCxttsaQ6+PU4C99gRzWesdClEasVTkbubezQ+1WYwQsWBA3
IMGNMrQ+wxrAYa6XIrlQCiVp83z8zFwHcqK02G2spWo25rnsfLpVVqgEf6DMuAYS
1yQB/mtvhYmhOo9DVfKTFCeFR9Kde7Sk0IZhQeoZefSmi5vjifwN2xvYWV1n4Ps5
sxdnaGGm8KHpuUwaY8jW5cG25/1QEAasLyZvuXp4suZV9FFVQtSGeB6Oe2N7WnHZ
+3tBW98+KaIF1sZ+EuN8KeuI+71Fl2PidX/fxjfYRMbcyPlEja1h89P+TNuLQCOo
0iBej+9i+UOtHqan1y5KO1I8ZmnBy9fgxBwWBPEPSuWhmPWKGHygZ+KXWO0kmAx9
3ATDUlFOOKznRHcW2rPunB+YHaGIPOQaUXjrtMHNis5PRQgtQ68tTL9+ayfzSwxX
JTCXY0EkMtA+0zYWzaMbIXlY/WRvgU5gJvMJfXMzi/kHHeaWS47BOZMPUnpAbwEJ
zq5icPAfJHNjsIjBxX3Xx0eMQ9aBiIQhxKaHZjdPl4kDN6F+9MZ/G3vuKHeeAvDT
vOdbjd3Ji58WNYyjgTX4cpAPlUeEVP/U0hmfvNr3HGGNe68hKnpc3I1Emvc1Y2tA
o4rm0h5o4oMO2s7oogZxaMjuYVFzUBY5xw98e2Lz59/JqDMGaHYQUMPIrYPeBsft
wogljugBsLfcn88MuT+nwxtpZCbESgie1I5vp/61ZmyPe2n2NSVDfPx1lhXrtZxL
veJRIa7TJLbzTY6Z9TCrLv+XXrpCnQJl9pbtykWEkh+f/2mA0DqvHVGHLOAiBhhD
xX/R9e2JVHVhK/bJBRBLmorYJDCYq85ZYrgBpRj0YQzhlKQ2xge8DdP+thtsva+c
rsIocvGDW/i2ATlAIfgFbZcrNGnLuw5spcfuiVZdoi/UL0z7WgbtBcxbjlZ+eaMt
YPCssvkNqvTFyqFm4pXfxpdRRC5RtnH9kkpS8jSGAZjNh0+AvuUGIllyYfFjAmGz
FoQs9Sz0Zjq2diO7/axVUwzc9PvfocaPB+d77JX4d+91UmJdHaKYWTSgjAwjIChN
2cJQl2BrK74sITOQmKqH08PdxFotNgdSUigCLdNjFyzM081Jv8iIXQ2YPW33jvTV
irbaxriOh+AbfIJYR+xQGUOqHCiGVgowWA2k4iG745Gggql5Pj4LpcAZ8H1Wv+TV
IQ5pA2um0ZNbvzpYu4hVGvpsJj16lf06/mQC5ZGPyaUOWnaBD/C3kHMfi+iYg3NP
OEAdx9mgU6bwvbb/83WvDWr7Jj+pvyVogbIHzOi3UKtottJ1/KVAZ9FMDK0EU+vn
DFBv87YxRs1zUZ1zy+v82ADbFExN6eHvZC39dZmdugYnxPFcDeh2C3Wbg+iKwJ60
N9Di84xb9ik8ybLkr9OfgYuSQQMCBNvBS9ceDTN4qmFt3ghdhJV18TqxzP01w+OT
a+6zjXqzbJNJCNooeSSTeXqR/nmvVAwCk7pQHS+9kKr/y60WDT5CA93ffbt4CCvC
fsa66cMPkQh+vmIQv1fWzslcPMtgeWzoMBRslrX8VSexexJN6Ls5IEzQtmBeX7Hh
GVTEPpRcwHWTKPCF5y/mcdcoFqhlcuBuYH3Ok2eShqQPUG2mu5kCs502aeQj0N3+
1Ob8xAoPbrtpvkFcyR21PSWGqFLvwRu/7yeNP1CDXNozyr3q1ePZFw0igF9JXqeq
hhoXA8PQmdnfXK6lbuW3LEibXH7HOQxH3uP+PX4XTs1OhfWJuMRjKJKbkL+PqmVn
fKUbxYm3x6KnZsNVCImdmHO6cLOK/y5GyWrkVCZ+NLbAPQPn31fy3E9F0SmS7SsC
ZZZBjvcL7ix0O9yvMVJ0B4npfpEWGHHeJMK+xIdTZ5Csm+rfAli+GURQW4fKzk4p
sxGTpInXpB0h0pgRGtwzM3kp6ygfm3I2MwII8EONQ6InH6EFh9rBN5fRKqvPTZhF
nT0I8L1PW7bmwlynY/W8loJGiHQVdwUVSU2XF+CdzqeOVj1AjbFO3aBVV7vW+2rV
zF/XCWZcvhV2DX7IQwFCVb1rF/ySu+T3Qc6Tfv8fff6ehAynCQPhw8BD+c827mHr
hm+g84bYfxr5chV/JzyTzHyZODEd7/bJOQ6HCuA4UsSJdwBPWrg+E2v7kSqWuSOf
P2GDvTcJiAShMcuq00Pd3WUpMotqAsN7Uo3QOB/e5qIn0PLWOS4MqDqNofubE+cz
hnrWy2cdK7k+XqpMRbJ7aBa43qFKNNFY8jah2RrsXTbxHfD3n+GH+Be0ruP1eJU4
P+itQUY6B0DCLC/NCQFogO59BEWOO9IkbYB5hXEQFfn2eAAa7xDtUbdfyBZiuQAS
P/1zjdA1H+ygzZ2fK4VjRAmA8GhcyMyxmBjCWOkOA0SD6GkwJ6AgZIejgw6bUiFE
lkCp3NjQYSln8LcVvuBfUGcy9yIViYfFvDuiztMjP9MgYN8krzNIsXgSF/vgejV1
lV0zSzX2gpzTNIgbFzrTTTZLnztO5wB3ild8AO9jCPINfzAWIHgV2JaumQ+X3sZ1
9ahlTcVd+aTqmBLsnLFeZUpydWAxt6LAR5RlO3BsTyJqKTZJZnCo7upcLF6Yc4A6
VJrLNIrxRaLaxMpBnKvmovpBXV4woVRKbSoGk2ry7xXCEUne5N+gJb94hkTjEoL7
3ZcUISjTTXJMiTOtV5wHhwxEHNg+oXNEXXnF0deD5jY91BHt/gCyu6sswsssAp5i
wwL0rQUQcmYn9MTWsubyjtP0hb1qNJZfg0GZViVG8T9u3h9r2wpTutUC3cqlBWUg
U6MGmu/SYtkHm9eR8X+t4M1TOox4PEIwQynF9i3BeNSK4Znjf/Ko7ikijBKMFFI/
QWkMjhXjkYoI1p6GxsI8YPP3rGlQMjznsdO/wPmbxIEYnL6i6waBmbYxcDt9F4sU
hLkUZkxFniv7JqHcBfYjRUSjGfv9L7xphan3PlqxPKYkSheUKy04tIywvqjca58k
mfo9yhzESrCey3HPOsHLZXQPxOL4WkmWAAXs0vIdPo9loYyInd/kgKGO0G5qeSW7
r1S9bPtQa8qvPSaaA7swdgy5TKjFRyuFx8RrP+MmnRMqweH3o4fSny+EvhJTWrjW
FNvE2oLLdeAuPF/tgHzz194kXFh7w8kfP9KU82LOQS5Ts85u39G/Tw7Fko/taTDm
wQFxYe5SLeGg/kE/zYTq8wDaFaN15Q+qVtVmYFR/iGSIFAj6TFn9TmTskTUXLF13
HG9+PQMMrR0ojZ0sM1ojI+idA68LO7WBiX9jsuJf68hPQXmXCTk+WourxL7apeix
K7KHO0c+80098Db1ft3TU0RIPAxhrsf51WjqxhzP/o7SE4AypZ9zpkF3R0wudsTt
yUJ3MwWKITb4E0voE9RKBJt/mGpWKEnkJfRuKT1Zyh2bkZzVbUsT8Pkwx8Pqx+gi
l2rDpY9xv3tQj63/kHkKJQ/N3g/3nKCxnkf2/g1hNKW1nR8VhiMHB5O1gHUi5Vzv
uRESsPpHeUBtbL+fbRCuaoeKlchC65nxDcZajsHgkywhfZTSVbfxhWtRcmfZHVMr
jXE1cFgjz0+arhmcsIs7brmR3GE4pZqymT0UXeXc1EWqlwfptn/GilwGYeWwDhE8
ddGHkDLfIR3IcjHiQXIqs+/O6audN3thLSjRDJ6WAoqtksQJqn/tR+RB0jKTWJI9
EypvGPsE7AgfL2/rG8EBuJ6ec9S+KaPuFJnsLUvmnZ+vx0K9sYvwHDtxfBzXdZMy
DC+c88r+k5nr8bG2FEKp9y1or/xowhrqSSApMCzu7MgeTYdRBn9w9mGruK8KvcdK
hOwOKk7aA0sT9e6VZssxJceFqshRcwpR5dh3YbKSXwujrqN++/DJmyzvMc4h+Bcr
boFq9VqebZvv0kOrhTYX/zJhcXhcuk7kr3BIB6bgGBXT9JmMZJ+tt2e9V3Mmfbzu
GjYcE8/RzeAObgPTT9iEsDZT/EkvpaVfBEFmMqsahwuDXjO/Ez5rAhqsyUZrj0/G
5STX88rZBak/JOcMAXmlnlgoiuxa9pQuQCB/wAwfkW912am5w4Aj585QbpFHoERI
XKhlhCEn/k11/ecPfCiYwngnlZ+PyCc2VfnCl60s5EWpGejmd0ukCUY0jqzEjwXo
b2GqyFYsqgN86tnB/x0fvMeQg0i8Nm7Rp5o46W73rE99RrcuJepdFSMGIVJEKNUf
zfc3g0ci4/eooCAHWBxRNpHGjldLD64xv4e1CvVH2ZoNsS9MXYb6pSSUJFrdrYTB
VpbhYIn1hlZWA10oYl0mfuJ6psrk0oiBzhlKqJRxofN7cfPq2SEwADilIKLQ6vK/
wxCv25opUfSRsU2ps4J9NiLhDvs9ttyscvHcCC3V8Td83FzAtkBPGJPRSH2Grj2B
3FCaIiFjjwbKSPRYLQeNULACJljoQPebLmLT8tdJM692JsWroa7RkYhVke5znWII
3KyAl+tDKyESsIJixc/UBhFQ/98jj2vpE3n7dcMlhAbqdcxQstJlXbcsXF0eJEHB
jBq7WuVAEIsKFJx/eTnyHjtz9cUwG+LWA8XeRqZNr1/ZS9EmeMZTO7fLXw1hNAZ8
JhIQUyHhf89ZsfNn163g94PL6VHFFDMstZIHj0jgAla8nz1PAcegZiCCfCs8hw5/
qoC7/P9ur6W5Mr71GlUbw5tcKqJvOh3//3vagRDklkfbnpM32pSxl56a7wr1bbX6
phQ8fFsOrAZLbcYTpDPkMy2jy/+MpUw0GBl/MxOIQ8x8pjkHN8VZrV4NmZIuQGdL
d+RgiqMnpj0GBx/3tMiviJpAOeNC5N0s62j2IGQGXsdcTgd2VhT1B/kSyTTcY5Ho
4mREagu3S5rWCdX0fobVcknlCujIwQiHgbdW545WzGQ61hmG8jjyQkd0xKyMLicF
HmYh9WogBE4lt5t6Mv9qce9WQgMQd9zypI7DgF6KHLJDQvzRQnNYwLn2eLxL9Mw0
Bp32MdxyPWNY+aY4qe3MFq9/hnSr4izU7gs4QgXJT9PoGRakgGDRtNJXj8HT66U+
mhxQuln2XuUwx6BEajQXdrcgTdF8kSzTMqUAzf5F7H24tlF8N0ZvlD/VH9XrTxMN
OQ/9MiWhLAmTjniV7r/FpV95x9ZHoOb3QVxOWspbsiN5dS4dN2CyGteJAEhPQqJ5
Am2hTLt3FClOOuy1S8qQEolHskihXVkIlnVq1cbRY8HNSZcYGfPVBGJWx/jUi6Cp
bY8wSvUfCfaIc5cKynL3FnC+Pc7rHhkyfPkay6Zl2CgPMW+iZamGRHh0t/2ixPtL
S00S2evUHq1ERiL9yRRbJ21OOJV/UjygApV2c/n4MDOOG0UtHrYPWeoAWC2J9NSS
biS09oAU/F/8MU6mowLuVf1gjz+ECuZMQviOovX2chpusFqRjwjck173bkgc5zQZ
6+5MU7Dds6EhunnpwXYldbYNpx8gi24VRso3lz96FDgfzwK7ckzrciGsUjQOLnV4
7LbZkAl3jqZEjrng8a/FcEMGV/zxDRraOFNR8h82qtQsc4Rzllo+YuuhM1yEaslm
I0dpawns12XDk/QgPgWQuOoI22tRDRT9XjrzfVopkQ5TG2S0AiN5cU5C4HY8J2pn
uVxUOx0vdweGVFF9SX+D2m22BrcYtR/uX3zaha68hNreRSxwS/HmoZ/1LDMHBPH/
HmpmZUtbrAarpyqIbZ8aDVB7Tp//lKirp/nUXCWtRjyJ7zhVFlKoqin8nCiSzl9C
c7u2/F9g9l1hpuXA1WyFHWofWsn7NNMVqyu1uoqwGFoZYJXzZuroKf/w7fXC0kT+
rLR7R6A5jqP3PADqcVDjdFOE0DWsZCDK6JDsH/ObrK3fRHQS5k8wqlJ6B0GwcTZu
AuUrHU0EkVylJaVtpudEPeL7GS4CqQfsPvscbQijA+k2pSql4Fk89btJesiijw7i
Ouh8UPYBRcm25y796BGfPUBhxKGS6VJtCMiL+c4D0EIthSuEOuZ2jLrNNVRjCA8L
4z5YaI6vBC3f9SoJQFMRBUohz4bh1PS0N73wjdw5WQkGOYEMRg4AVIO4XMWXmcFe
LDPCucqw9yZ3wAeWlAcDMr/D9f6CN08tYR4jWHUvoYBEunjhVifdLUzQlQxYSA+P
XGLbYPGB6oS4uWicMsdahpdyvH0CPMoPGKUc82MBHSx/bTY8AR/ePkssn0efaEqK
uZM1xyyBilnJrYFy2sa7loT+Tnv+JQw5nvOraTqskO+uvZ/Rmm/sI/kiS4lPnMCX
IU6iAu+IbatJ5sX058STaO5AMDcgJxM83rLqXkeXjwGIdUQSTrd/fGkeid0cC0rm
Xk9nDPs5dsP/efazWmRXKjfrklIrU3H1pI1c2yiXo5e3XB5084K8H5K2DgwPjvQs
bHGZaKWZvCNsljR9JWR8YA2tgUDTLYPL2aFLmY+ndVvr0Y22GZoNEuYSxGpSSzaE
FqhzZGsgEM7e06ncG301Oj90nMcvtiRrxCGIrvA8gQ1bO1CltVLvROpGkQueJ6iC
92nxuCfC7j36snH6l62aWOZO+p+ZCzkn8CZlMPEOuwoX2zzVIPdOmjnXMpAjuPa2
oXvbH7iyDMmsrCLFqLtI5XCI4gjTLXZ/tlpi0VQa6TXLoDVl4zQccndzLNPT6wT9
OUOCRF2KjySIvd3xfr6QPwS92uBnFU5jorsDUaKigvOVbv1HkcIrZpFDEr2e9ktV
tm700/ZD03xPaAWFdNai25t2tvWGhobhUeH4+BZJeX2n9fbw7a3adTuHKM5AILQN
JQffiuUtCVmS/by5R5uuWMBMrr0rtwVTS8LKseUwJBA1c0q5lGWtUtSA2nXzKI3S
17fFvZ3k221POk4gyH8J0jfvlK5zPQXEJ1sX631IRG0G6tYRx14jIvVMY8pDwDT/
MN9TbwwANy5u+wEBcTpjQqBLnqaXLnTFA+doqETc6EshdWHaPxt4O57NGOoPEtlY
T+lnVgRB7Gfui7SjMyPkQzUTbKMYqrV+lNwQJ/Mkval2kPf5JvTWLCwDy8S9sZ/i
800moRyy5c7mb9yZeu5k6Y1EgAfRZeDjFdNMPBkZfiPqaM8un81kEwM1mgs7H/NH
1FBANDCFjFCvZizgYFgVvVpx8wxdLrDKwDbdagIUCpTXaZS+kUvtJzBHhQ7D00Ap
tJr0dYKiBFpvLZ/ZnMtItdLy9IfDHtf/CXlm6Uoqaz9sTcTrOkRJGlM0qi22hbC1
FHb6SJ4kAmcNGYdJLUgjFmYww4/m1RgragHmR4AZDrowY1ibMtWnkfHWqcKV8hBQ
lNROD5mGxIfUupRZRWuHvD+6PY5u8+SzMAIQlu9dI1MSjrgf7PgaZdhrjYr1MAgU
q3yInR/oYjolc2jx9kcyqnm5jnKJSdLJPTgrlnF4yuP9G+6hQm60wQKS4s2RJGXE
27DYGpbcPjKk1htw74Mp0Zpz6+Kudggs4ZA/XFuOdHz7qFaXkVEEbP71YU0T1wEt
AYxrMPCIdF9nDr+1EjSbTAKmuaG5YpUjYN4UW/cNQzE1WcLocakS7zYmyYzYSoAR
O8fK/EASgDQe2QlKV3QQVlmnBPk3GZSSPjNHtFhDVxriUmoka+wEet1Sid6gUzNq
OWuxhjLJEJhy4/ZaL760GyMIHyBuCfs1uG5YuU5zznQXeeqth+HAnB3k32vWuQlh
uWLPkPizNOg/0azBIiiNDG3cdc746ImJr1MqL2PZI5l4cDqi0p0HfxbCMyW8nE2L
ErurWAgBCmG7Ns/S9s95++zIK5KSCpoMoyUrAj2a6eYih5HNhUjJZ0KKsBB7nGHe
KDQVzgLDdVg0sTu0Mh8ZKhl7YvIfw2dKl9y/TgbkoNCRsGS3gX5km+iNGMHGTaK7
UoZm1yltcyBEuMKQNgvZZiMts3AKAoOrwePmkFi84/IcmaqaIM121VKWldxBIAHR
54CuAAF1rQHPtVg563t9zTwnEPOmV79goCiWm1aELws4lXRnsralQFgzXjHy108e
KeDzenEQFrgEtUxyuwoZnbH0aLW00edWvbKeko4+sdd8Bt3ho9wecZ0ZBXO3xb/Y
J1OdPuAwvacLxesB/JghBfiFbL9sd9J0F6HfU6Ne+Jq+XQYz3ja4HLwEEAJ5wr/5
93b1fJpT9GCgNlzqVEB1M1aNT64Rx3TEVE+LpFFIEDM7ka//FCN1Rwmc0wayjmfy
5o/QsdFVgFsXkA/1X9/pN+vHQQC/ABGLd1JUNfUPIDUsFEwD61KNvLvGbEJSRJur
2n3+4Ctrwrt94xhZIUAOVEl4yMDBPIcguk6013adzE5JX1LgyXHw++xFbTBfO3Rg
aUvX1OyC87fVpnmmY2HtM9lYQfSP8nxZO+BwDZx+DzfV7cM8bHC0Tb5xCnkwx1Hs
S+VN0WQ0Dog58dnbhtcUI/ySEUU8yEzSzVSGUgGdUYo0SBS4JBSqtGKDZysCodtv
nKXQ+v0Mj4zIMJSJDi6vMgADyauAWb3ywljAyU01+7xqRDBDjepCXd7Ad8T8d3df
99JTO0lhNwFKOlPC0UA/MN7Vpn06xPeAirAqM0+VNv+kdKz0roTfE4DGrQJNJLUP
vEaLNGq59s97CRFLbE3NP2aUgiejpWm4dpLfwH1w5ARz85jt5LG/trmrPZNgs9KA
XQWTBdPLqmfgYPcUMxvl8wvsvyMgm3/rebzQeXbxNvIYP9l8hdLDw2Q4kuXojt24
oPxzdZ34HREls4e6x9uiHxfN8aY5Wkapkl0ErApEknViuSn6/WAn6nZA2+7zqLm6
EFXwbGtl9BbOVGI2KToHkMgjRNQnZRMvpNdAnGw7xyfIlOuzamCorTaGaJt7GCNA
3CLXVUBZzRRu4KQTi4dLRX8ku+eYab7y3TyVmCo3tIHwlSu22cvaRr5tobXRl1el
Ha/Oshv6ZoZc4PubOZON7c6w/WuQFA+/lOYf6hu30bteFDG+ht2UHepDIXI8+Urk
sYGNMGtpPKDJse53kYip2J3RSZaq8WrN8VVqMx1d4yzhckBmNELy6Q7zELIqKS9f
bqo/fjCAIiuS7Ssyg3Bbwk5jtp151zQGr6AXZNt3oSH7MlnhRQAQsPRGj8zPHBNI
R3oYpiuJ8ozoKgEM6p2tWOmFj1Usf4ZG/5wpTBZkInHBIw+LRud6tinGG/4r2O6v
I0gUqIcda/A31nLMOYBGw/uThvmQeMNpY4EJjMJnYPNc+1KEEF54XnD14swzsx3u
SvES5RY5+KLoA5j7xTFYLRd3VpJ2mVtFY6Dj7qf4Q2RsUmy0/5dlgTHF2JDhJglM
rb0y24vPhN86yQg6uj+CtJXlll84wgqlBr7p8YG7ihOdB2HI6D8KD9SbJIU5asoQ
4TWSVDP89xba0PO1fkWLv0h1jfnYFNWDWMpyuCS5WN/oX0i1JJmmqE434wh1O+/c
pzPkPR234Pc1f3KzhO/H7BTuSZj0npigQbksxXGEta9wi+kEOmFg1XcNBYtgXAIA
8NEjoLdhrCco0ibpl9aLhEhFCfuWRoMgfaNwnXLNJ2B8liFMnObPlt3FWyjpWSib
pfbee5nNT16M6u5d+zsNr9SIwQjrzsFZArtCP+Lk6PJiUdDg8I+74ReWKPiBZrCP
tmtbaDGETIr2Q6Bwb0qS7xfbA3Nb40eA9qJ98u32uVmFVxE49K7ZNCY7qSxDcuzs
uDYvZvyWhLoVJg91D3B5aHbPdZkpiKHDvk/yk4m9acgcPdXU7VrrK0doUwPL+rkm
BUvgPSQiHhCgF1UK6wmt69cLilq4jD97NP5Qu9Wh+NVpQTv+ZN+SrrtibNNF/bhk
WEhG6tMNuc+UQLGbyjOQf57mBLr/EzpT1/cdsxyR9Nzn7bYQbVKu3/2zg2Kj7125
4qwjNvjBy8BmYy3PKfxfXnwzRnTh5cjx61/clHTag9DLyAi1IpkmLvRYXdIkhZKw
ixsVWWp6SD1rB9IXyTjzhDuqqZ333DoRiqtxQYy7KD4Dn8WJpiuR6As0FMze4qQM
zw1bjo8YxFiRpoS+wCSn11NmOhXf23VSuy3PI9J+Ln8TA/cb8Q3wPStltpP05Ips
din5lOC5YyBOJiHdHQBd8HT3+7KQNgxv5PN7AlnBHyoLhKfwIfrG+RTxFDLAZlpN
cpV57tGFJXkormiuCfxjLU3Y5ZrlaEahlx+wsky5J43HV94xR2Sf8dhmKmswFjSR
DyhYpxUNDuzHdM5/+6hHIYfRNVoaLd8mTV12/Hdm29416gfLB9Mwf48h93kHNJFN
ezceJNVgKPyjPR59VXs76YUTl8TEHpwRrNDraLPMU71xyfn/QWoQaJhptK3M9mcA
qRp+iMVXhIjm8exdRBY6VgDDirRaS3FD18Hxdb2mcwdLjtdx+S8zFhZjDzcloAW0
eFSp9MIDbXSPA+REcfitI+3Qt+UEt2cx/0vqfMQEbkNaSJxN0CWhRE6iIcwZOmrr
PhI+95DSLm9n01Mg2uUzGz9swJv1XS/GZprMWQOembVkd8Kjy6c2/tx2jOt0JEwB
mgdm3IIEYuT4mPt9D6COLa3Mw7bgLkWUe8u6B0PkC45Hgjl507IuNAl1GYS3rI0Q
fcVtoIgAOi5GIDaBiyQRzFY5tBRxhlDCEDnz4bcLGFxG6I1tID0EJxGBM7BZpXU1
auqquIUqIg86zL4keDKNWUah2EWsk7u3UO2vSxYWoClZ7Aq59a+MVJu2ImVoP+WV
e176kKhGWSZ2MK3nHWDh7Xxf4z9R0MQYetA8fx3otqUAFs0YsUWYszXFrNH4+B/9
AIT/gLDBAEjCPAxMHzC0sf0QaEkxFpNj9JhJ+WJoWh4YsTAzxwQXnBkASnDGz2kL
QLOn1rqIQxgxq8krCIaXkBucaHTGennQ291FyRUUHmKfITHuACDHK9ZJxdpBBGKF
7B1KnH08t81304yBDxaZRjLXOclUgv9BDHPLrZdM4Lgy7JSLHYdtluic9m3RlGIf
K7rr7pAjARedrCMLT9E90GCgr1aV8zAeCtCDTMEEu80DVKFFF6JzZOH/hS3Y0TNt
KQwmNZL9kmpZ9xe3o9CeEtZR9fR3yQu4WwYNSiHGrtDgP8N73oZ7c7sPC92AfWFk
klawojOU7ekarZRmF6YHWiyQaUFkT+4tq6w6WKhdQnKEbr+cH7r8Xt/vbRF3Wr53
UZLl5FFEsqpSqdXq0Xyv1/KV71OCAU8exasAUxJwAcRXgg5qBTF3WGFyq9a9rTeh
FSClHAUF/3+T9AOq9/zIuw6c0PkaSkvpP4i8NAwGwqbMk5jzOuzr4zNzIlh2ikdU
X2lQw5TktIgne6oqVu+M+g0D5wxdX90UYkulkAm/mWKOa06nBwcYqfqYf0lNgqG0
6eaMr4vqPw0lllpfUKTOTc2SqwwOIP8EKn1I3YxNfF5GwG8tpPFrCf/PQMzFnYiJ
cisdXp5HuHb8cDzdqszjQlpIoVrOA80HJdxsUYhOPFw/fQYUdyhH2nw6G4jU1IRg
DZ6ysGXSdKl070Ay3vL80hC5VspQWKMt/HgihqFNwvoEJTb9Qu0tuZugR0vQrncT
lJdKdxhQ0RvrGEWLk4bUEzf/JH+wnf0jL8cFd7DVkAKx2BhbXVoYsJ/KfgUJn0UW
1y9xTLuKEH+22/9A3WDM5x6Xi11MOPf/zFEvZID3lufwM1VUqYnTKpfjxIU8FAp+
dg7SeP/P4gRuSGbPuLcHBWdkFDPtLx1InCTfOo2d4hMb2aEuYZAPCvHpoLrzvv8M
FOyxv4CViuA3kvh93U1r8WTgKkcOYNUJJPsDt771aTwSxjZha6hPwLxD40pgV0h1
fTWdekTbfjOoNYxEBpSnYyQfijLHczLv+SsuDR8dblUTPKhyuIS5gkH2u8j9erRY
EmfHKoPfAYoQQl19u5VB0exSnQ6nvACLjHabhE8wxxO+HU5xZOEnF3V2STU8Ft3J
s5UtgyuVDnelMY9H86IFMWstR9VrobFJzb4gJvRKpHMj3P1JaDcFg599hdGUldhB
yi7aFL944WseLkeUDuS2ph2PnbdAPe0nW8xMuJVhOy8V7vQjfEnB+et3V2Po7C1i
9iC6Fl5l+CQDrBUnFLYdHlAFnWW8aFcoW2tTqzN6nvsSvbKfeNzGZJFT2uuTR7uO
rULn8WqYkqmJrUCZoEH9QQMmfMXx9tnI7busxde8vytqXqPuhG6aCb2Kmbl+uK5D
p3DAvGgbomRDOaNDtjcWrh0RHU4gToWBAIA31ugV1RnuJIFzB8Mf6f5XNlBaIyLW
iOUGNV8z/ci02WpapAeRFTqXBYC9ITOfyqOtHEsiuY1YUYMprLh2jwRSeHbjtkw8
BZT/xlC9TEorRCBLdAwN+H9SkD02FdykVUYmVLDdlZuCJA9Dsh1fSF2/Jw+YzhQi
G0dtaqDjELytWANarX200ROo5JrRMoMyhlN1CLHrbh06RIefyWNmJL8PbdV2bevO
Comfj6IQN/pEJgNfTL6pwgzWdElJaOaPUaMVbe+2Ld6hkGqRYYBoB94VXwM2y0+2
/R/LTANR1FZ8JDO7xZjp9oUOC0iwrj9/6RFqqMJYCvaxFlphuR7vphWHyhcWxxYk
c7UzpeArChjHGj/nZpVuXie9tclMy4E7I+LboeDvdsEvZc1+fB5NJypMqXDhM3AV
t1ik+cSZsChgCfCAJjSDownoeXGMg1Fh9op1PkYp3TmZxq9ZQF0HVpYRN8PCX07d
3V/LoTTLe49HMxFVT1+N7RIXZYYMQD+fZC+/ZCKDN6PsLcxZYHnDReyy/TDco8EN
jlM5Vi7qZ1oeyKxEnaShBs1NZK68/ItTUl9IxICyyxSB816EvCj8vtODOS2FAyDX
1wjW98oWBu7mmCnTvi+gJRAVkkVZIG74UeGE8QqALtrH8VnpnQMuYuN43uHGP8lx
y2LECJZSJ5MisCVScomymbpe2bzYS4Hm34QjXIAQLaGe0ndRIsYa1ivVxGXSE9j4
Mjj6RXmm3uyL7wTg3XV38t01xsZ3dzKUW/3wyjEppsBxFtyKka64Vc3MUCQrCKJ0
jKpkc9J7WgcRD5QC3hE6BUdUjKpk6qTdBsgUrogN/kg4ck7YsvX5eA0IOr66EGWq
yGOgUxluZGz5F7rH6htgYTzomAd5LV+LXMqBZvoM2bgbcBVIsLV1HSOxpNSJjADD
XqmDLBeDB1rd0YqeM5foVYlgSBx16mODU0sxC0HSNs+V/m+WAM7Xfziipq4yGkN9
gYoKoHsMFZhLLiNhcRbQjPt1AKlC4INJm2weEN5FbDPgpe/w4Jn0QMWOWuUo0iou
h4axiDhJsT1hrQ8b7SFnr3x9h+NtCE7HTu5CPC5E+GStrDNo8aSD2JkClar9vXi9
qi0x2dQHOEMkbz/rcCbZQWsKnKrLZu72oI2axfylZeR0jVCaVZ3luIoxePu6BWiD
SWUxgJWwjFiDlDLzt0ze7J8dx2rfI5Rie5zKQ6AsgeQH620LGfUpf75cAnS7ySz8
vKmFVOMNVAAlBJK5H9oClbREk4gHmUyv9JFWR6yfx++PgO+4OXFFREowt2mVSs+j
q5w6MBWhKrHi+NX3SFi3ypWrKwdf2tRe/ciQ37AlNjVayof8V3hZKUDKqF7/VVjk
uzPrjCxrepkW1DF76NDVk/Q0fJkSMDe9t+upZ7kqjkbe6fmqKYIVPkre8DkaEoa9
9B1B7q9PAT2ZqgHmVMAtAY+dZjZsVDOnSoCexXCZBcMzAQSmAqJ40sLF3AbcvSUw
ncxFDiLeoz5fY5OJlF/dww2CyTjFK5A8MZO3nSZTf0DgE9rRViQsSW1/7ssTGDxW
hRyKXJGo5HeffA3oiGi/Gjs1MwVAWJL6MuJmNBI5/BumIjZpY0n5M+TTEd6CVNv4
6Q7Eg46U1r1ip5zYdGckbCrIGtyr5VHIE3F9bUuE2KEHtymvtXP7/yYwmMJ0a3+G
3stViGSIDsVFzm7MB5Ac06zG7RSia87H9xLXkeBvEUCGIzggHK3f8GUEY4IC5mH+
QktmJqM0winTeroNu5YZXIo6JaBu7sJruluL/9XFda4pvMJ5H7O/f1MZKf3KcB9c
Ffnfinux5bhFdwr5f34xhiCVVFS0Dt8ApIj967c+Xyn59jX8SVJR6doiBSan8Z9Y
gd5qAJDRhNGlcnRFQ6GZWm7VaRk1EV9JaT0qZVXYVQ2dRrP+7PuTGi+wpOgQJSht
mOB2tXAGVXEIkcHURvtn422x30OKpJP9GAkMGWpi9+z1tJS4WEsTkrcLSZhKaEtp
BIwIpEnliprA5dITWPwB+SJUgTB+BcfhJk0SFoWd/vCJ0TmluXxzA5WMm3+DCOCG
4At0Om5bc3nQ+Vy6xmz3wY5zBxJuTl/aAngNyOPaGv7wokZ/7K6CQroFWtIrUovh
HIQBR5/wD1kUs88z33FCYjWmljq1Q4NpXikWIB/FpxEW2GRO2Nx60B2ub9vxj05q
y3+n8llhgwDecXQWhmdVMBF1TSidrMqlx2wI31XbCK8vF+gEcczJd2N3IXMMu1Me
/c3QZ9+uSL6wOmS+4MROjFwDb5r9V9Rn9+nTe1m1BLWEIGiZw+SBJlZ8MieNuVJM
89FuJ7LBNIQtA/ly14Pr1zfrpjA4ATREBbDUziIkDSCvfGSnwEbWa/JuDVPfNckd
a+GmM7Y2jNmwUup9Rjxah6Bzr8/CAfZgYJN1xZszVWCg5I92az6Suux8LTfzf7Cf
Z+vs0rhrh/dvKKLM/oNxmTQnq5Pg9je1cadsAyl30cQcT2ciU+pjdYuKcAHqfZOn
tICLRCwnEEJPoT7KprK1A6un4fos1sCL6NOFwDBO/WcGF87powDi8C+o34oSlhCz
teq72x8ZMNrSgi8BInDsdw3v/bxFDgSjhLEPMbs6FW8dd4O+K6f8NCAPYygLHk1P
mW7TDjbDQsjMcuBIyxDxyk86kxdCzWbdqXmxk/x5GccQUWViAu9dVCBd9RrXAwu6
Vop9PgBcffUdkD5sXVCzr9eguyKnj/DSRk5pte1E4yYiYX0n9Q5VOd3dxY+mXSi3
ZuZO03oDd+PcYHArEs/Qzi+d/vBs/JRj3jDIK5JK6iQLL0xX0Ip1He2hhH49p+Eo
ZN2PF9IBdNMd//ymFaEqnYsfU5IgEmKBAEDJyBReb7xJzyttBil2AP6T/lpwvy3n
XA+6SpR9QXik+VJa/88kM4kbzRSDFQv34WTx3TYIwRruyT7QfFO764W1czNc7s1T
J45aHDfUXQAQdk3iXKnbLftOtslZ+X9Bwe09wPboOqKHaaUGRjNQ5hSwO8ZI+GKS
MVZQPgl3PnJxJxT74XbfmLE4/9SP0x0POGTcVkE9RnRu3iEH1AqRoUYyegJB7G7x
9kwT9J+gwFU9nZR4sD5Jd6BpOJEMiVQTnXPD7b9lMxZETbagrV2naWA8WsRdxSrR
YnociwtEEb/+R2vbDn7fERl8tDhIZ51heZDdH+yL0FFG+8vRuAjivUmMnnrNKFZX
elm9a26UXeaNouH7De9PinwpmBviqIpEFHA/Bw3iEJ7rKWe3DDh8RhzR0iRyKljv
84Mo2aPhbnbcV168zT/DOpDqOBOSKhhu7BKqUdoGf58Jc34n5Mv0d4dSXujO5rL0
P3T37cRUpsUT+tRwHneyIn1/sjEd8wKeYX7bhNJ/1kn9I6CQ9UXAE2Q3zFj24rJQ
qrxE3b+PkKET2kYrbYc+OhNBJoMH6hGCY3THNdI8+ghc+0kkE0yzbG3ulz2kYQ0o
Q3eIbo4gyYglmvnEGK3YVNjEWwQXngJcuHINDVMunbs//JKSQV28N8FmcP3DWBao
/8VQsq9++2iiYmUir9MVAcOOao2OMNxDlOaep41yw03zI/zsdDOhegTsqzFPvP3x
ZvyIMdWpMN7/xyuZn0Sqr7eexvQS0tTklH5UnDIfKWVIYZjuf8OpQY10MNCaA3Th
UfcuWAJsi4M9tiwBCe5itdu34GGpZLBbVfqQfjiCze7A6yLjgZvGEVJuS5O9yQr+
7Y1tYtFZfDQN9dTLT+sOriunLWTHO3D1T3XlvlYmEbgpzLCe0dgWDn0HRciwSjPU
nz5j37rGSYqTqsuiI7wCIxjPVH72e8m4YDfKEoEW+ZH05t6bS/wmhV5+368KCzTv
amF0J9t51YrLLgyWHTMDB+mLvh9LFJw4xUijG1WFEEs4M6dazEWwpp3464ao8EAD
wQEocqsrysCO9B0pAdoLK4850kpzShf/9xCSXhpfvn7PMKCtzGt3AQ/iUWbNKGoC
3duXVuUs3dJAESDYqi8YNAFabRXbjS+cIvc8uOJJrUyQkBqAsXz0OJ7dXFEBMsO4
20s8RxLYKHQ6fL34kXEElEDRWYWdZJiwKYFp9yxkHchbDtJDH0NMMdn55yV+su5F
RT/aous20FBdmU7ug6ZHW26lEKnWq4oOYDkbRvF6N5pRDtl9kq+fqUImm7NoaGnf
OhGvTZ1VCoPoX/cBrSD/qL1TKT4sxT/D0k9rwi1g56UP4mCvDML7tq5Bw5j816xR
EQeRV979Cqe+FCpHOCtzoVxOGbMbypK7CDzthFAj7pgmKrqt8fzpiKtfZ4d77QTT
0Wp8hgbwGkVkIlyFeTq8yipdxCOks/SmEne6KXv/xPjVezS8IuW5vdCyQZBapVHB
E5pjVd0qFgMCkKWuw7ZzPmicPqZweZJ+9arpEUZxltgMF+Qg6CKThwDTbEHJgqyA
UGtf8CNHi1pjbwJadVNJRAhUE0TZs6SIX4NVDkqzPDZo/m8e71MOKlvNg5XpwukO
L4Pw6rBT6JhWPJ87nDbXhkxk9zWQvZ8iEa9bEPmO0SKY25zlxoO3nEICRX5UR7vy
EFTX2Ztp6952N4WyqFenxw2KNMyikgFbh7jy5HSSNZMI547+GwdUTgfT/O7ktuXm
iFeIL66ljdIy6bK3ANyoTm1oP2h9wMCcUiE00qdFVnXmJH+MLfaYjABmHV5B7pFm
Wn7yN40Ubs92RGQWg66IyhuUyMcr+1s0Djs4KFebASI79zEozcT0hJdkeBLk8GXy
0XTH/MS7fiuuJdU/pOl7MZGyyX6oiQ6XEyQM3SoqSdwZpAAX0P9hrJxuzbJvfHv0
KnK7wvaLF9K7YG09x5ZWx3IvTViVV6VtpAJQVKKn7hCujXhMjXIRcXwgUZIDCzUC
Bo2ZNH5K/APS/r17V9iQMGBLv+iB0UnylZewHFoJ3RNIsbIxGXjL+pWu5OgdY3cp
z9DWP69qcSc0zuLYW3O0rz3HvlAow3hCPU5xS00sfW7iCr7x4A0wCBLtXRBjj2AH
6MNlViZAAwRpQHIed9qIETM71PjIcWilEzwfnPPI9KW6z2dh/RSBQ0E0LhVbMYIK
tde395uaDHvye84vQOL5H4jsjlDexrno1umA4O/+eqgnpLzIkYekmxB5q21z7n37
ui2ZjYjNUz8qbuv71PydPfksTurAFU68pMhZtRXJLgSgUtOb1/UTpkQw/qE1qrUO
1I2ISWBldaOptWj+7tHMMfpYKnBEJaY7kVDaagozSegKZM2X2aTBXDtElv3Nzy+s
O2O9sigFQubO6AuPpHKV9bIl6+DEJLNvK5tpCtHkuSI6HnaSbrhjJxZYq245/DlI
ebYa5GqEWzvxxiRXYaSdXlcRtoeF7xodjF9kQdl1d4QUldRbLBrdKiW5Q4yutM4z
js1IvCN3aTAr3TuT6jfrU9gOBmsMpVFbdJ1d0K0s14KvFKs6MUiP2dsX9RokSh8N
mdaLXijnmI7uP93HmR0w1qluBAZMvoXkyHimqJXstqV91J9wWICK7wylkuIHHirp
SdyvIwedqL2YxfZaMLtpTxq21XixQ9Mw4lybaODHJSYey018bgmLZT7wx6SWC428
eMx8kXKLHgLgarlhHsHqx31ZKce9JYSn/hG5/xZEFkb6TCsWiWdl6S2UQzomy+Sp
m16fWChtZjn535Shyj0YrJYavibwPMWYIdWRgAWzBKnj1yl0B4B6g/zO7xTX4mlO
yLGneiD/uLp6Eios4W/qjDIIQ+add2dI/AKKpR/rABPXIahzXUKLp2uWFlAiJwgL
zAXwdFs9CO34+9djQonRs5kBJoFio+uXAGxF3o2i+uY7bAhZ+WnpWklBm2SH6+FM
BDNV5ITniNFIsojtCeLgc+Cgq9X06eXmT5bXQVYonTjfTfiZMjmMGvEs2L6HkWti
eaLGc862DIcLiZ1XmnhubBdwC8osrE3+G0PRj60j6Gz2p651am+LaBY6ZEjATuT1
A6nfCAxrV9Bs9eoAL4TVcLpIIyjlMDAR12SjKE+chCL2Fu7O25dJdtp5UGsEL236
8EOv+LeTIWeIi9/0X7NYze26CwUFA1TKziFcTaJ2fYVzd+2PlKlEoyyMxIh50dWX
tN2uIJerFvDAEs5UwfoUr6a9IOtUlbezugjobHXGxvtu8F/5xCtAZLbFakguQCpc
c63XCjATZYBQIXkHnlgHT+tMQFD3JOBNtPONNk3ob55e6BEz8CdimoY49jKbB01e
2zm3WjnHlD+TDD4Qt30Vx3jrg2KNCipUGq3nVN6aTkrlXwuV13GREjlXbqGG96R8
W2rhx5S+5RHYyPknJJSQFzShboR1eEhbkTQkNRa23dS1vsnYo8sxyXHiWUu0T8gE
6erPaQPJSQn7qpnt00eGd//8/uhT24TsIibLS0bvm5UCVhP+FT5E9hq8RcMX6lra
piaY5lDmeuciXiYu1fbuFC/sFV74qmonrZZFy9vzU9kEWLsJbeUFzreH50DJ9knF
H9S6JjfVk9FwUzRyz7On+3HLEpmWOx1haaYuEkknj6aVET5m3U9FuPPKr/IkozMy
uprHFQT6bq92JISr3qEoFOfXOPVuw7enXHcU8tAGHe0ZxiD1LEP1n7wiaukLS4+m
EXUkE52G4DKQSqtzbvVE2Kg6c9xqNDcPjoMv9YOybzKmrdhtLmCfRN334ylABkUe
KcYSiXDmvwbVTBM3a3XNc1NjC/RG5coSDtAv3wlPVsWTAa88QZT7MLDVaylajaDQ
0dqEMAIGdDlYliGhJCg/2v3m6RMecc/1cmLzXJ2SN1+G2WnyUuG1pxMroaRKQHjr
JL3rxCWARQ6XtpIRUxz3nt8a0fFQ4keWCb04DGsyrfyXGQ3S0hslIQ4T67xf2t0m
27IPlMuEjLZqo+5ZtaE0t3QpLa98orJ3ch04mX0DpaKxPV71ZKNBRSmx9xkm6xXW
1nOkjwNuuKCBsOtP6S0AiFEdQK23hxBAL46RO1Ya2TtER+ooIF+TPPvZPka9de/X
XfMTkNx1LD7ov5z24JO2ZSsWL9OdO/XrF6L+xa6qZma9CU7B/IkJZEfr0QjLTlxe
mC2SeyNFZOvTHxKdbpfWGLfWE4idz5UFoXMiINi7olvPRVPzkZgOC0jEosk4uaNC
RSuSxekz3nrC89/MXBWmCtHRnEOBVzWqlMC3MYiFWhYRfW1vy9ANv0+Ta0AXFBxV
6lD1XOCC8dmpKzsMyCRJrzo2cqGXQBUF6SdOVY5DnJNT1esZcaokZa0srq4VTcgl
4nCqRTpJI/K8ixmkB0RI1Jf3Dn8ZOzxRAaRRtVPM8b+epvr4hSK/IBusjN99cNKP
oolCApiDkYTee1iScNZ9LMDdxF3C1GCpbJssDHFTVrSQodo8ac10l+BB2NQp7hIV
pZ2dDvyqw2a47mkFvWlBPyzpHbbTNimkhp8Iaf3jAk3t6WAxcGqIv9hKqHPBlaM7
SopP6egppHuAhlQeIgUIJTDzCzMlUAhS2uw0kP51Q2zEKNxB9+dm72JNjxiQyaij
zB1EAgSQ12EQQN/q5USU/oQ2OHn+XkI/ldknJh+IUKTLp2Et7FNBzqk0ur/Z2SZh
VlbcAsIz5kpDzREJn7/PvvV6h7hMmepNV7PnnMawANuEwFEleP/JQBFOLN8hEMbE
RJqLclvAd2Amzfd0MUrhUm801y77pZKZcCC5vL0RMgy5/JQJFurgWkLN0z36GRU7
Noo8EqOHnmdO1IGZApTPh6k1uZnCTOQEmyyj/1jaYxz551gg0Lxir5gHqBk6W7Vc
RefIiGSBLHYGY0TFtwzf49JlOlJhDfFYr81+4gk0MtwE7DpLPLKfdAZxLQRNlu30
Qnh19NCCnNmUwGJLxiPVchIs2M5fNdOB++oKHF/3+YevHzhh+63+8cQDKPWdRRTu
G8CcwFR/P9xCsEv9mNW/HuVf7Tf1SNzaBZBisPYLYxuldFnO3xJHITm0xHQO1FRg
EfunY41oXS5/Bq4xR4ZBm6eTRp/8XHi5xkaW9teTGmzspktt8LjnfJl392qLuac8
HTNwJjum3uDODsq1frhe0dwSq5NgUB71wKXVtIPCPaUDUqUHWX7NtmPihKTOgQN3
IfZ6OPB5DyAauYLx/V7k+Xkf5ZFNZ5jrQ0u9CentJDLeb3jXQ1fH82KZ462E3tkw
AFKGMigoxO+rRTGrmdOdkkAAg7DYDPtLCGnwMdwTPVBDWoeiBCU43cims619CgA1
OAAnl//XHViPd9LRxAcD5EURA3cw03KAGguEGPgOesCbZ1eVeoKpoBFOicwl4wqN
XbpKlyaybQr1i37+n1N4ajcXsldSmCbz7XIW9Y6g02+/bt2V34fy1fauhkB4JZ+z
PxVtzc0E3IskVTJ0mYhF+BAHsCao3URW6Tun1uNbd4pIBPkP5LEtxxvhhgPWckhh
eq05hWmfhLOxrNeHT5CN8xEcH8KfcKM03g2dYWBdAbVqu1Iw4RvFRVK48F+HdxMR
7Yonke75gh0/xqfhzuF8taTFuKvfLe31RWpxlqZweT8gTBdsOrZNnijVrkG4OEM+
srRhLdP4a8sM2qvAJZ/UeqOfZxfRj/nUkgEn+ROwrN2XlAUhZCY/EIZSv7nce0IW
3PjHxAdLsKp4R+jMQAOzerYJ02IZi7ZVV0M79qHSWB/bQFwruEcWcm4rpv8BZJgJ
+WQ3zQGyZTv8elEkt88QdOagB1XYqRfP64PWdB3BZ5LGGayWUnBt+VnFMbjEJN40
KbdpaWKRdtek5PrD+t45VB3jbK/fRriujBsLnw248okSSUeymnSUoiaDqYHGe9hm
hoLkooWann1a9lj7iXZEqIQQ1scRLrPjHbBZnbqVkwBVaiiwB0bo6DT606I4ZM3f
ZEuJncWdKAq9+ahXeucFDHPjQO+6Xvma4ISo7ncuor0jfbHrjmq+V+26/O+bmTC7
k5tJCuO3cWEJtRwEDhcnZaKMYxwfxMmbxoQmqZFoLErE7L+ypjR6XeCEczHL4BCu
2QLtNc+e0I967HIWuXxzFlInLRJ69ljicJZTEqkZcFnfIvXAhZy6iqZah5ulX/0Z
zQp5rrpGo5DpN1jpJ9FPN44PgWhSOFy0rsN2AbCreyPgxlECuhNixgLbr+5m7mKm
H007EY54ogtrhieNJw8PSws5OhU6bLSRZQXHVdw26Z57hpA3ozJhf+LC0oeMtlmR
8jBLzFSRunbii1ufK4TBu83hCZ8CGlMmTqnYo5lapDa0Iwm0hFHbp6Rx4MOd7G3u
KuK1w6g5bKnEIxZS9zp3X85DqtOVyrZ2DcIAzYjerA2x26KFJTuLnIitLS2LCZcY
JB4pOiN91BkYn+JhEzXE7Q0475+iCt1rxQKTTJfyXMAXokPFuesRdx0WPX7p08n9
9oZnTSRqt2b1eeIwZGMDJj7O8qbul5na82bt0UYxLOD//zfEriQMVJ3c0FGClMu7
0hmqoHIalMwe0Ehdkg5pbDVMpSGCbeJis0FndzfCaqUogtivpF1W8rWtIp+Az/EC
14qGCzF5Rdw8Z1Q+4InMY0blFjcusD7nyBOR/iJfjJHFbWc0Dvhn+Re9kfRx1FRq
R3cowrvehFCaT+HuIfd7alPXOk0CThEt1njPplYWUlODIsxlY2r5eglmpN14TKDA
FJr1UftmnAm6AzBKfOwdsZkdjz50+wdXTAjXbCM4Jowm67q5/0APs4920mdO9RDM
/uANFnMvRGydxGA/Bzp1Qq0VKgdmEsUEj2KsIkFCo3TwbyGcQgwA3z/Y3qmnIMFa
e/+N4h7uTwGBP3Ac7dWNauXqT+fZsQndkNmf1eDEO/cE6J9eG7b1OPFHGwPwqcog
NjynLWs+sJxC/mlMfE3EestDwTC2U1eL57x/x2VzPAE1+YfdxicKRg6VeGKARraE
XTK4vYlBDyoQ2NsLsqNq/qBKYBCUBCrSttbxo23FW7PDYFEXIlJWtYmEvG6UV9t+
g2vnJdt3/c5ZGUN8UjrxN5YeYu/kiIqgHloobvM5rxq6/mjbvAqR7UVGTO2SzAXE
VdnwCG5xYESytWd4sQqNNqydMHMOFSgLs1QS79zIuR9y5IVYOowyi2xUibj8Kiwq
+XFxaEAc5wmA5+hDP2dFpNedBKgCLJDC/PEQwv25udBaF16C1/wD9m7ayKg4slQ+
qbfy1DjchPhPzmFJee4aOxWmF+SJVWpblXR62oBkwbM5Q4hmgYSC8MJsPdUevAKc
OB+BfL9in1X+w4B0iQO+eKw/Xqv9VO+9bE9yhHtgmQVBEzn9q+yMs7wedvkzEQJE
aNO+4eGWx6wpqeYi8HYS+cpVGZjxfKmmSXI4FO4QVKpys7zbCTaGaqA4Xl2KlnVF
7lgYKy4LLiMChzKps/XIA5GIpSptbwX7TNU7UJ/yOmOnVOPZ8ZUBHyfNEQskJbvm
Jhh4sKBGKrIY1snBmumxYymgOQKFvn5+v/+2l9/JSTnXLluN7IGVNTDoXnKZxqYd
Qhor6JBP061ovOg3/G45UBMcyUKbH6L1YeFHSDm03J08GjqXkwk8ZVpeaoEhFqHg
TqCIC5E5e/BNx9hWjvL24m1lXrTD4Uk9pUGNRrfId7wkhDNPBPeaJBbyYqthmG8p
J4u70mxCFPAfoVn+unXWfQGXyvrrpLbtFm0iyKP2I1h0IgaW87lUzgGB6AN4VFKu
24GbxwzTaaqh4qWFqQqvgNm/VZY1kTFI8yOYkbfvcLWY0kuKq0JlZw+lE1u2U7/U
daXdTDFEq7cUvkwXPIhZ/d9RI5m6Er9Bw2IVSY4zZMjXUccots7UZIueA6NHSteQ
2obGCnB4bLe/nQb4N1xyqHd6fPkl899cmizrYfOizrXO2/g/WN1q0E4kHJxFF/k5
IwFCtu+/tyiF0SGvjmXOLfI7c1LoxKte19rs1ZPgmP7ZM3qoVwsaIvB5F9ArcXg7
P2knWcrGkSBJvEisXjrDAutFIv1hR5g8V/leTt5508kT6oWLXah4xOo5mA6cAr2V
JS9L42y8FZdeyNuClQ6I3zQA6/nA8HK9pzo8ejTc3oZf1vEvyvTGdlvUd6BEP7PB
B8o5iDyWwX0f23TP3Z0EuwN7B4IQOosdCP9DnOUaKChdnjTzxaQxfjNecN+7bbEW
LjnbJKRiaoza4wlr8r5whnme3FpesTEzwAw3NrX+wqdZ1togeidS4Qx2ykoyI97l
c8Y+5AIzO9uUnu5V/7Jw3kiUe/NuIhI2M7nGjhyRrpYgAJU6VTbbZl4Cv4KLO2nf
v8mxi7jmXsrIgLUqsZpZNWP8tIj/jsQh6+/h8EUVPpx7fmXwAUMGT1ZRfZ2JQ+Jd
Po8r67VHwq3L+m/ESSBOg6DK6zPqf+YshiKmdqQvcNvu4bSxHsH0/VAUuiEe1VKM
S44pTzJe5bxOqofQGnFqkwwIWfuyVQj5BPUlXtKbgRDDL38rdV/Ba9LFR7aSITm3
L7AwHPRNRHGVjTarT3R8vcV7zKzI7AW176PDOWErhZdr8VxdNp2Ac/s6YYFPN2SL
9BUaqB0W4EaRXdgZ+zaJLCFi6z4w1aQT6WyL4Mw86VXv//0YPZBMWSeJOjs6OhSI
SOGg1hxYQTyW0c1giaenSvNQpTGVjobw2cgX7yFH0asPoQ/NK7BNxYlOly1XGgmI
8jEvGaRifp29OChOXR0b6EDxDJW9uJ8xSGU65G5+YMoxkns2pUMl1AOmrowUk0qe
LtUXaY+4MiIDRtTh+FgB66RmBHtZNBeZZKr/Nlsw7Z78n2pmVT6Kmd0ESPjtxOu7
kvcurvkQq9gOPEwaTGOPlrha8RHnUMjuGi0g1BvnAWH9yTTTP9cKKRVNzpE8DVlb
/aBV46jmIdFEhxkSvIM+BQwl5zgYURfYYV7rB9yv6pRbZn1miL8sNiTCId0ytRp1
22obgUOeSjpb0Wd47kpA66XuYnXVz5esGuTGpfjEOVPVC7YvTbXFktjuDDYWPOHM
r2TPHx35vNKIOJbQVTe7ktxt2yTXSx9NoutjYeUMwBCEgL5YPnLimEycgZTwtywK
unUccGv9thVql3yZo/rzI8c3OoBjKa8hc2n2Jn2LF1/D7soIkJpMuCe2kTxLzsB2
U5WvQDvWA9G1290HK2vsishDqdtuTZTey11drW4qyWSruJfz7HOacUnm7DZ2k8IL
QbIxD70rkREE7rfKTmGSUHxnYBrhRwzmXahrrZw3+QYj99dM/k2JPrngXZwwNM9I
ia/s047cfeVgkLTOvi+0RPjsjjf0vtZZ15+WJG8//9ZVcriR5ZEHbFy/LMuzBoBD
7RPH0RoIOewYZIl032G5meHRwi4vcQmqMWJnXCov+uhAEwaRgbB9AfYIFSlV4AGf
1JXiaHUwBQ3Xr7mZBNrnUAcg8l9hG2GoBxXRaZmPyv1HZAYW7sFtWvJaAKfHI3/Y
6CoKtwn8KMZ7o7hFWe5x8vSVKdsqF2fEt7wzbSBUgz2xxFa5nsSTZzBzDxNGb+4G
04SE3wzRgvqE+D+8Nw0MhVfKz6BdKaBEM3gKGdL6Xv9K9fq+ZfcVwg9Tu/JzZfko
vlpwNFh1Q6Pr7JaEZoSGn9BoqMteE9DPy3WcDiecOdwn0gbHX7/zItiB9jjwUDYW
us6bZvfJeXycsPfTmls+S539vCD5Hh4k1EHpJsSXi+dHugQ791yHpIDvfp5fMYnf
Dfn9MCrExGuBlib9sqHGUpA3YHSkToRhAaHoBf4zwEEt5qWzRlH5USjVVetapnm3
vdcrNmPakkksxFVd8zkO6oruKZaKKYfYYb0duu1J4AimjZUreR0BojbSp+Ct8t1k
4X7fm8hExrfERQJmEH9P/7LSlcaz6RoEsLxM7SvY3i0JLTKmuLhIu3Jrn3b8BN7+
HfqIAacd0FZKscVz33D0qWJS7xiLvZVoryWu2/KySz9At3/uQqbNhHDekE31V9CW
AEPCI1/mpNkB9m3Xu9nvuQIxXgQebjicWXp2j9nZ8r3CuKCN4Zp/NuE+I1oohg9W
8CqhnheAv71HIAHd/pyXBWVDmS8El1PicTrVmuK4oGQvnruCOEIjwk5WZ4mRhzMZ
6aAw2jDVQYyBXMjQ5NcHBsG11SW8GS2Q/qWXiZupGxXKiAmF5mKn5QbYFB6kAbCS
a3b7d9fmStrn3Qo3mvgf/MHeXteLBfc0MAYRd28I7EejitaCakzY1e5fcIom+lRU
TmLFvVRFaXdvGhC7q3DjTLvF7oMkMSMS/rE9UmkZRqowEr1EH2ZVe7qH1BDl0skI
asLJ0RL560jzAVmkh/BwPFaLovZHOw1Tfs3x//XjVV9xdjMzn8dTfaHIOu96wD0d
ZMY+cZqW89E/JsgghJ9fij2aCwXPSGYFHfKAdjE3jPN4xYtOstgATwJ13Znf16Gc
bM3dBJNQUBp8ESSr0xDF45tCCNgcFSVNomDSwx2bLU3vRtcvknFfHIZcx5g0MKKB
sjbwdroMcXEzhfyA/j/ImSJTCnek7wPROCtRcjl2O2dsIgFEcsIaX/IjKIIUG2Oh
nNn69irMC/ObRYkPhTMdZh8RJcveYRk6QX39ZQXKObTtUlr1v7+1+wh+L3IA7jsf
Y5BFjkY2dGEAAayi/SubKvTS10LJ/qCbcLHzifBDlEkjkZ3XerrZOX0P82Ummpsh
XnTu4egf0VN3WnaNpzUi5mvW8wMo35BZBIateuQV84hd/NLlfS5CiZfLxD9EJT3o
sTQJAgIc6I4tIieIi0mz8ACfMxveYVbymW4o0NTrvK8IuL2A39lATd/e4DpRjk1Z
MmaMDIzxMsd4MGEzM5dfFXuUyR7T1e14nhVzJBtxirCwpDuZjjonz+fvXtK3fHek
KSxN6qEMeZ3V/U3H1ZwHg2ZQ2CF4Hox1BMuAf0rQaY3i26ywtWdlWX2LoW86nBdT
ig0cUFFI+AZqr4GLNzH6bikaw1ppZxN/97M7Cee/FJBp0vUw/8la1drQMF5YZAgU
/aJSRj0WSOknhRDswQL4K3w0kT0gSJ1SWguP2VRBVzFnHWpGTNwKp79HNhfX+rRE
z5lQ47JCHCydV/ai5eOkR8deC8ugtPupBAECThBYZ0RJF/6gc7IaD51OxTimqQo0
dQ0bq2MBplV8uNuZe+o818QzkhwoLQ2+liV9j1q//0oQt1JDog8nJ1+N+1SVK/Sm
LehYwDV+W8g9wC+FM7esrQpAv9wQMPqwH3KBnqvQKXl6vr1+4BcNO5kOXDIPMPKf
iHtMYcDYcnvEuYCGrcSMtM4NnXKonJjxrJ7BTz4mgh3ZSkb9btku8v5Pryx7rcDN
zN82qnkSKpQdCJ5771dXIswgg5sPNQqawLIL7YE/xF5BhHdi+g0Xuq130x4shka7
Pc/mejRCSOkF8cGJBJ5wjVBshakB3wvo5QAqIParydrmWxH4A0PgQ5P0gN+Sk7fB
U6YGtx5pRRJ1w/SSu4G2/rEAbczr/QJPUbsRnxRGPCNiDGZZPYFT5dGztYFCOTDC
IuVUwiBSEuBWYgO/REGScKQGITM3BgZC0as9aQwCg7379Vc75Lyfk72S9oAqKAsR
aMzuKFYpYaAn1GIXH/Fir56n/w3djnu9b/VwVz/tsAV8RbPDxxAt5r+4sEoNF/MX
8GTO+mxMmHiQ5ep2YguAEgVc3d4DYjYUe4T7W6Qt8qHSTiQzs7p5O4NKeDRhhsUW
mzj2TqHCoMOp/so+zBhL4QWq8PXRuBJG2FoAioBqI8OYj0yXfxdEHLn0DUZAAHpC
qvNepPVr8Bv449F0Kja+cVHfYQdwYVbDW2bL+QFugrBGhzi15iDaScRXVHscT4hX
cJqRd3Ztap2VBMdgq9QbHLwJ1+3q1ou5xKV54QGjFwKanJtDRD5bd69khDNpjuTT
H+ufWwyUaC1OOo4I55zFbvhjinqECZkUwgmJ5yslew90njosLE2rlpRquQMbG/b/
fi0aTo6Br8TjuYoiMGQWJ9IWcBrzux88ESm+juc5bx+FcSMorRL7//C9xkplxu3i
irSMXmkE6n/Fbg7mtVazUoZhdaeHvwuIXG/dRyparDq7fCk9XgrrBzphmsIS/BDe
/MVZV97HM3eRWO4kQm94MRFYqHNZCwXQZf1dAd1grNGqTS67UK6YomayfDrQPl9z
aialrdiNVpHy7nrhtZgvn8OQF2Ikny9cSV0Jm0+kOUaMvaYmQs6NlsFz1baQ2aOB
CfROdWBqyrGwZ30xjEv7K0OsOCPRVuNpDfyzLAOaqRuO3u1NDF+0GfRJzZ/zaR8t
Mn/jweSYC9C81nQxharuuOQ/gv2HteFjn51OhIdK5thV8VBQrp9FK2TzGwsX+pvC
mnWF8y6ey4RQNKHO8bnI+nFaovLSZqGEPUMsE9fBlAc+1Sy29Om9rElQzyYUx3Mj
VgeeNxO0igJQUEdXm6X+VrwjC0XTGCJ2yKJqZaJyetU5iGcGjI+VI0OplaiMM10/
TcVtcQNnFTVUcQBz/sugZZHAuS5j9hfrYpDAafNUcgYeeqI1HIV1OcDZuL0OMeod
2wVSEGyKyuxGsWTAjdR5rcTp4APR0CYty6h6GV0eiTMlmTg+bJl43iz090MOC1Sf
Wnc2XvrovfrBMpkK+TFBZmjkCn4i8m2vl5WRw3sAG/6qk1AxE8W1iZnqECQvARV5
asdpvsGEsb/cYBEYlRBQYBqjtO3ExzlwFAsqgpRxBvHhcwst5ALvvFVyAsTWeLGd
a+faLOBT+JotP0Nqdhrz1C+OR0iuVNaYgXYzHzTR3uK8stOuz72n3NtdKfnrAL7v
tBpfhFMZ5qEiRLNmFePIgHL2maRiPrTR6eCbleU46b3M949VZobglHteqwzYegRE
3bBRUEt8+k6vufAr+vnu/osu+LxFhzkWqEtXtfQe9TeQtWQ+Eu+96zW6kzAAo5Ok
gxarfCLovdavGBDGF+/iFEUR7NBXDtpV1KdcsSVSCCfviFzUlq9OrhHaoOnsA/b0
eT/uuOCJUn2+3/qHokxgAyi5gRrP9ilSabIt/ekoSnso5NjlrdOyB5z/ref2Ycqr
OUMHM3aNC8i3fQl2FteIxDrKxmM0H7D+QiumcHyoGRc2ahU3Q6WMWre5M1fsX29U
tGj+K3wTR9f1SE9SvufLVxlKGAYBW+b5uKcwdWrA3r/Sbw08AyvIX6YEugO4ljWI
npLk2dj1Gzk8eRE7PhYSdjEFP/iU9lAR72d0PT781r6bOXhST1RkQRkvg4wnNiuh
d7DpXic9b5hJAb7sBe4EnTlq5U51+QwEKoSVdCinnLj2C45xepg5E4elQc/dmrLs
Y8n3N0pBMuvOcqW/oz/+onCcIVLMnYv94PjmnP2GKGcMO92HtV9sBwPKmobnCw1k
x7LYETtk0yjmXgzyu3wy3x6XqvpUE7NIy6atunKN7E4TQkbWDQKt+ut1vx7nua6u
/knImDMKWKskx/st0V//f0/xw0OzxJD0A+zYObvG+qbWn//8cl5wLbwmv699R231
okTTWMtARM1FJUlXQ3w/SDjnWqW5f/Rp/YIb1bUooHedEli771bL2ZerJxzQ1H/+
q4UIM8MRuD9UeC3b7RHBfPryhsv/Mzuomdzapsmnb6XHAy0fRp6VPPAkukUSvmkv
pSJI3RNe6cJh3KZHhgUtB/Uc0QFEZteMq2QnwuPhXx9H8VrMGa4ey6SagysT6c16
kAVL2Vzhq5AbnctUkeuGSSuMi899eU8s3fU6ssBP/hr1ktDhy20UAG5/Nwjggj9p
n5dtzN6Rgt1NR5VJzYG3HMMj+5cjm3vC/sXuQAkrtA0ovTC6UYt5UPO3dFCsMqu0
GXe8nxNC7SSc6uRXI6uPdrKKU8Pa/yfkhgSnlrrAjXAn5S3E3VMwTaHeVbmIXWVr
lC4D/KqVQNaeb0DGjPsN3IPMHSEQCZ15+U8dD3EH3iXjYZ2O2obih3kxj+3KDkhS
uEm7MRCUaXPWxHovhqynXZcnsTSUTik2lk62vbIaG8ljjd6fpjFyCgK47Sxr4KhP
iFJw9yw13uUPkY+JRiS/xHNBqy3N14x8xpZVNXKUcwXWM2skkkZLOD3oX2lhmsqD
CGpC7eBpJOHUuFyZHghD3R53xm1rklK/vbAcP5BCnfUAnLghxA/3Nkw3alulU5PS
CvM+hafb24jfGnCGFXgQupLI688lsWAZRBWoqSNqHRWLf2CtCGW1OO5Jf5/96T2w
1HRhYMywPph62L37OyZjJMOhY0v5gC9KI3h6jjyUPGJkPqI4AsYvzavngr2R460s
rSYuNA/tEjhPC4h6BbjupMziUUibMHUAzsT+gnbtxOlPumzH3Qj4MiWgbcbtRmzu
lIx7zeyu5SxcNnesCL300jdFhQzdJYjD8/L/P1tNBLltseYot0ZVhtksYxP8JvQ2
E0Dxhb07GyeYOgteJ9pW7UDUW+QtZFC8SB4+Nr7mivD6QCK+7xEgCcQ0iPYVijfq
ozDtjBbYbqSGwWWIG6rqxR7s1zLaTUidXpkFoGIIJIp5GUR97LyPOtutkkTRgRgp
b3xfOa6qckl9zvgcIdI/HMNwU+/6e+YXZUx4Sg43DqPlhAA99hDDzbhrfGbayhzD
Qmz2fN1RLejEnNYnn/M7e2umpVDfsnqAEXGTSFSvQEWzty8zCRxAy7AKyfHmVaTt
KqbGXoHjKUQ+8S3gcD5XnHzDh54LrFYE8GQWmrnqlnUdJY4YYJM4qRpNEgQPcpDo
aupTdk5tWa77emYW0s56h+OSifhXHMWKL2d0lJwZ82POMLpSuFDgjjuhjw3nVHeM
PUCVj3kF217fSskQhchFZOVj64Dyb8xQhanSILWOXMNPRJNRgt/TC3G6z3Gn9Fzx
/FDs8hlwwbXeY8tH6izgBM3mQMIGTKWDE24hakgTx6kdS2yNiWBODBwW6lGPngDX
az3P3aRnQ5m5j2g/apI1ph/xGoGMtc9BMfj2/OU1udAos1qUq7o6H9swurMQgste
zuNGstWAZ0L92JN/aahVzlA+xFq/Yq95wut5LJ/MglrN1VP9GbdpBtoUzCYgn0ga
s0RtJHnE92kaKOQRZMbtjq3nHEwyVMB/PPXBvPydSlBg1Jp91onbuDopub/+6zWA
pu1gwJBktSALtucUgXRfr13T6U/SCreXXBgrxOPzEfZGAEkryDwy8gTpB0fXEIw3
ipiYLF+BQlkvGbx/n63DCZ5J8QkkuqqDXyEG9SfO8rHkb3yjV8MRIPlSpx6wyhq8
M3R1jbW7LSZbd4ATanyKH9x/05+wAHGcPrjT1NIorwirwzctxLwM5bIFmjB+/GdP
xehDAfrDXVpUxEqFXSr/0OTivud/hhSgFQoOjtnRPU6gdqkGpbmygrlestdVZcy4
mHt56aTMZ8KCUhaQyeiU7+cJ11BqXLUERohqavYj5Ia1EVVe9noSDPXfOHo+e1lb
Qxb4OlFbfpjoq3BedEPdThsV9JB9VDUgQ8xmShS5vS6WorNum9xlKx6skWfr1PSC
K6V/u0OkxVkib3fssGEWeLRLpG+TbFeSYoUTih1BcgoHocKqvpCxzXHg7bQQHU86
T6Xr/ifD10IsXjVfoo+pl4iSORsxHlmzuqpJaB2t9qG0uaLVIU+IyKuugI/TiRzP
0Aav0lJtkWG0ZVgkle5tFPKpGnXK2IO+GHFzf+EIDRtIVIuJOa4oBtG1/lz35u9U
rq7U03Joyd/xLDQxKOrRNcoEEy24IwwYMgM5o+V5JNOR01irYacA5DBjWw1MaH1D
8hUV5aiWCq3EiUGmndFzkR7sYKyK1sEB2AfgWfkYDuboZrWg1SYuVIHiuIiMRvXV
zESiENz35gm7yB+78tVScbQItnkAUZTWGjytNBS4e3pWkD7IGqzbGtf71C/uvG3b
hRKIClSOBTSr0MWHJ1T193ZU1Z7iwil5yu3jNtWfOItY9g5e+z7JANglTftuksPK
aIP30THY1sldbvd5zAZM5w4gyda+xcwh28OMH9m7Euxgvpw1BuJGZ3vD+N7izR9z
qyV2KPbB2hZlan+1luCT/c6DZSU40IBXdbbttEP3VdXe+HRWj81jYDUmotcMKQL4
8ERW9eoZ0fukxd807ZwU8ohSdS9uptJo7UH8MOOEj55VRB+QHx5fpTgyZC35MJB7
4jmzDcp8tx6PaqlDf3GLu6WQ3czYXqkqa2Bb+WbRWdzinkKTllV8ymx6SqD/bqdW
71irRwHu83glGcJsjAbtqIihL6qrdJFKnZzSpE/43rNY/FxqSj7CVi/2c1V8vO2v
o/5vmMUDbwX/EfPwGRhZ6jumUjkQbao7hT3TyuPkU+bbJOX17rUBDuD1wS7LYFz2
MhAN1D9e70E9vNzxXJtm5UxqbAYX6Gg4sge4BA7QaX5tGeB2pRkMB9nNwtShRXZT
UFaeZvwLWnyPFa8upvIMokfIBs6y2g1SNUyZVDGGrOvy/LIco/teR59AIxsDZ083
nZz2IGYCrnSosrKdIj+I++CoEK6OIJKPBQ/Fr3HyalOMgALkcU57yD5k/l6WEkSO
BlMF6cndgqtMx4ixSYc1K0UhPIBJGmH9OA19Drv0naFdYiWpD0JqHOdrnPq+tDxz
UrTKtYpCL2wuDuVe23/0I6RI0ViE65iFoQNHy5kE844lsjLlnCyfOGPQGIYcJSCl
n7PelfyjnKmmPEzNmJJ5JfHrgaHq/eVMxFAWjvGttk6lEVGLKNbPMbhdqcd8L0ZD
8kzonknVc0lPtCnC9zZOQg6pRHyTSnA4i81OSZIngcVFF4/Mr054/HGlsw+r4Aem
V1+fKPNzJRjH+hDq0udciN458sBac8kNaRzPL7fS9m/Dk28F2GR7LBW+DjMSHeci
+9ESfewUkpjOgIcymQLVcurlqKU21FQs/EgzMgCiOwpHi2r6pUiHefgqnTx5/HRA
SWejPFTQC60UZWKQUAsu2N4J4uwWpQBH2zbzUm48RVHRO+sNShpE0EX/9BssedfZ
YTPLNFsUvib3OgcTcIqhCB05K8TjrAd2moz28+1HVmGpey/ZvUEwk8LaJnjLJUcz
Kar3Y+X9xkHIGGwbkeYtHr6hEv9kp1TilqK57VDvhwfD+bUvo4COS28ExeXo9W9e
Py5w2O4edPEau7Gq9TpLgxtPFKbkWDJBatrNuiw+cXU85KJapLhfvTrX6Dvr/vRW
ud8iIElnbGYi9z7Z+/s9e7Qt6cqCOY/cZ+1l7Rmvm2wxHid7wJNSfcWmXKW+Kbvq
uqkkj+pK3LeLSJCXZ+pUPd74E/2oU8TcjOPgyf22FVywGtuaEoN4aZel8eOLd5G5
0ZPN/cbyuP1Vdc6hgQwBNc+i0wEqXju43tGdfEaHjeg9PGlumgIwCWzvfMTCmB5Z
6OYRKqfLkbrxk8l+0iyoK/2FOLp8UukoFXSuMiLpMni9nRuC/dL67O/L1uGsxVwH
Kpg1a5GVt/ADoVBnxJ7Tbv/JUCaxteBXiRVzF4C7Ehs6SVFPdF6NYAUcRK4RUTIA
UtPk+fbjJFpJXhWjdj/04X+exuOwIEdhaMkTmy8nnm1wTVugPWjEqIPnAwlO3HLi
8cJEGZsulmLcfbAKrpbJEyC3QJQ5B/1NEilN7HppM4JnBbM67lOZ/1W0SxccrkVr
98790sWJaPjaCDaQVsSK87G0bRBPL10OlahWYfrvs3wgtsnGNIKZnhqSYKr7a1Br
KAeBMISE5W/YwlbCZVBU4HYzqB82QHQuwm4bRymV/VF77KHjiTUX6ZVskTaJqLBc
d+dqeZn2AIBwHXkcJ2nYe9yI3AD5b2VFvL9b79G6v9tCx3UUfAJD0YWtk0xEtuJ/
ypl3bW5lt0gOw4AwZekBd07LnAu/BYh6hSYGSRhBjuvRqvwQKt3ngaMy/eT9zOaT
TgCSpGWGRQ+JkRu55YEBl38o9hNruXnaZBS4nU1c5c45/Fd8SyOxaEXgzAYSAsGy
PeBBzyBdU8OxHYlzPaQ5nM0qjQ73678mhND9Is/0JQdJgcHl9+67BGda6kWI4rW3
lg8NdEv4WqDGaTc3h5bmL7fYW5g1Uu+KlFiF11RSkSwxqg4Ms9DRiyr9qxoN+foV
vatFcNv1uOsDlUxELRoDIvZlBGS/BiPw2dtsrZ2fs1qK6mvCFjmFbcJZD1wi1gVl
EThWIXMLTELKPPvGHMCyZQbaViqAbcrMEMOtsVLaHOO2VlFTh2mqwRDnMUULZwby
DjYAvK3IuR8ieyvvnoxtsoYkl990Vo/fv5eO25nrOchNdNTad6LE0R/hwg/w6T0X
/8C14xS+npp55WgizKYAvolvzVPNWrgNXwdafPSfWXznpf1g3s+AXp4EwD2woSat
TV0YcBKawUgx8sq21H1gWHCgZVqjKJmMX+Q+ph79yK/ejGH6wqSPviU0VPN8bG3p
iHtkLE+5l8zXebUeLaXdGusWzMtWWyB1bpN8Z/MpXYDzzTGp/o5TJogWC8p1rJo4
wWlM+F0PG/Ur0DAXm3rLFsKYXVM+1cf1ndWZsEFbbYHdIqLmUiMQk9UvdegGVphB
aziKWychQKXD5vSuMmxmFaB/LiYqjCiE1FpGCc4Bk6Vt2Xn1LF3ShC+d44hZE5Eq
W0ROLi0dqaJ0nBVEz7m6jGW0uZ9VFwqj54o0d0PCZm8y0zQPXGlBSmovtUqN+FsR
XZvNxtUYcMXhDLYxRCrk02RBz90ig6L5AZhMH4OvNfd92FuS4l37tF/0ZrxuhRdB
+SZolQxprTyyWxCjxXFWN9PCkRz8Ex8W0UvJ6/cytnW5aMdAz9xe/VB9PWfTWTLZ
PH6nWTIjdhPEgAaRreKG3VCbz+oYKdJ/guLbkhOhlmt9K10+6GQ8K/gxrekBsu3i
P6+Xlnaw1G+HCot51yQ4VsPbZWdRqBDjquV2bMKGjqpCVAIwBkFhhU+ZPYkAu+uN
nuIx72IMHRrSeZD6Fw2UTGgHrnFPTAWTppJov3OmTD64ncovmlb9Ds2xDcK8+L2M
rN7rfE+kbfNbCCJBFG/RX00FGrj96Let0MBEIMNjiQMm/Z8HLdJXX9szi2CNCyEi
zLB5upxWimMFbJ6jHagtFkBfD+FIv4EadMDQ4XCSzU4XC6vtG4IZ5dUHkQpFit31
SPa4aI+lSLNW/RXSYpjERVcmu67CxnsJq7IyT5jw6tqxArMxcrbt9Tpze+twuiic
a1HpAqjueZLXew98aUeLXiPKQ/sP3dngGJeLDqFQOIoTVmDh17V5ZsQIRfUcBgR+
PAxIdrWAW2EdOFtQyRXfFsJLB62V99/qmySxa/L60WBqhBLbOnxveqDHpvOMRQsc
MulDQvG2Nwz0XiOqw/ToH20y54C8g8gkvGjoNjYrpYPkmnFdBPhm9z34CRTG5W2o
AmGLCKpx8xIJkwkh0Gr93Y/r631+9DOx+uZ4Vz+YaxMbF6SccIKhbYDIogIOPKEY
e/y5+2dDmxd+qii7s0WuvDthtXkNIjO1+TvM3r50WQf+w4DWe4tsQGtXNe3SCnK4
ovKgFFWYBqmaHc7yjhYS0aoPt0LqmkajyUUvjJlji2nlhhr19mwT2Y5QxRMMcWOy
tAqDBQcPbnrV2AylJAXzgLHlKpCAFbFLU7ZAw7fOJwjTve2r4104BiPI3lRg5CF2
VYUsy7RdMHBZdMfHhpT0BKKvOd3plRqXDm2orIDvtNgQKu3AD/IcbFPpqy0vCnhc
JL1RCfTF0h6e0uZyS98r5Y/4TuG9NQYbnloy9Pj59Cq0DCaWtD0MncgI3KRydxA+
s9tb2PdlG2zV+TUTx8jA0AocHcyy1hD7SVPHj5EjKLlKgaTvbsw9shGsU2hVVF+I
/5Lz4Zau281SP8WehZ2lDaBxk+LbiGbYQDu9WZPQAl4psgfJdU36f5A2njgcqX3D
vRvddLuEKY9dgGwX7tSfxfcGNKJUKQoRMlvLo1GD8wRRLiyHYd3NyQD1au43sKSD
ixi+LejC0imVXrDhJvbq5ZazVHg/K+Q/Diie2jEZMH+zRe6KxPxeKFvOer1mRrSM
jZKTo2VNSSowcila1aqnENeUljzxkbrgjjfKykKoTDojUNL1KRsYCgrkK9g3ZkxP
AAPqEdX6q0cqyh0KOmwvqXkVVRHCAUUHMbQk/BzxFxfRso6U7SFNv/ErZmDKdYct
NmifYw/6yRKk5KxdKNV98KBlTxsmhjRCa0qqdQs1oCOLDD7lpIwpirjmSNLSvfjH
rS0mRkuiaMrauMdaOIytAjUlwI9K1ugLPDgmi7A5gRXuOB1LP03hRH1q7OQKD2Oo
+DRpieaCZ9lucBfBrSHNiIU9nmiAJlWb4ZSquerGHoJTtkm+2hw3+yws9UR9zR+R
WXApsWoexv1zbn3MsbXGnWqpsrGTt5TmfGZsdgRISgxGM2MJSVj+K/OA8QRE4g39
CVNOICHwwZTS9hRPk+cGw/WBXiDvQnxxW1KicSNfqOCG59i3QueXd8UZkxsi3Ege
wU3A2k5+0xWmV5NS96eMiG1HXiyOVes+XiapB/VuUgd8agUqUdU3GlN0dKxcA08b
0FJD2pjipTUnqQPnWbISbTg744mn6PlqY4NspMu7mtvccJuN20gdi6e7aU1bEMr7
1LIsfda5D1BH0QwmSDzu/un8SMYbZf6F0F6GElRVykzfkieQILGy3ir2JpclS4s/
2AbVKBdIXfnaS0r1eG7rGDMWkT/NEXxohYG0KH/oX3htSW3ocwG3Ss6nGIXfmQXB
hDt6Wqu9HHkeEZb+F6eDNP+5G2iiniImHIa/LEtTgYvoSOlK/DBDbHKiMUwx8Q/z
AkvqLeCqws18WNA+1vz2Srk1InXZ45arIzPEH2jSN5ayfAJGRwOeEIRFmXvvpPwZ
19tQu0XFmmDDQuweFLEj82myRHZkDBYYRTatbczpd0dBXfoLbcTj/d0Ps6wXtoLb
/H3ackkq1DFwcEeyBNErfOOdhtRUg/iuSEZyLDhiDi+OVO6/pWQhv4qAYIRkzHUy
afOi7urRWBLVYyGhXvNEy8yx/CACdjGFw+4WsIbEvPLUYFzXepDwoM8Wc6xy+/IR
aluzJf8z20lk10P7f0Q77zK7jwW8nUbAcJ5arQVtVth6qGjbkCCKD6APXAjefyv1
yGsv0B/99VnNAo/m1VCEiIEzP9TiN/4owxI14fK5+vDv+gUWWCp4UbIvV19q5J6g
fMQ/PTvqZJtgd66l/9KJ7e2J9SOct1OozORfjWTJMVf9Tzq5zmTnZWrmUGjuvPEB
KKKtcp1kWu8Ip35EeQTinUNizeA2hzI7tEZINwVNMth9xnv5T3SjrIUgCp+ewjky
X00LDqgLgnJ8Hdeo2hFXR1cmoGAJGqsUsfGwKwihR/3KxnI3epH46eYNho/DaGGp
VGrzDPSy7B6xHSiMA8ZBt5wHebacrp7DuNhrUyiXJ9bfQPtQeA4OGlYmp5UyHxZ7
eRqqwZO1UY85+e8cCtZYC34Cvr6+3xni/EZ5D+x7aOAgJb3y0nKBKAw9dJ5XSXPb
r6hv//9Zv6UusYVUduf4923V/ARQit7WgLXzlu2hbwcQieNSPXUkMiAMtvRbH5Sn
mPcMn/4yt2HuogIgxAbIANp9T7p4YPV/xsNVCRnYxc/sy0A2XDCS+WiHVlUm+ikA
1mNdxtm7SczPANiIvhNY6NHsc/Vqe9qAeDT1A/dGVqfYxe+wVyoBJhgkwm3zDm6Q
2APR0tyOj4orbwoUf/5MQ5k6qrB69imnTo3DDx2y4juhLzuG4D4TUeuhM2N/8lB1
+jwrq/EtVfblikg/GLNnGXnqRaaToHy2a1YfUyUM11XjkrivBxO1dM7RNiU13deV
T8xPM1rcFNOjqkCogbT4IErggG/brjZuVc2idaVdMAhh11KfcHyztKHXBmcjl7YE
hKjCNTVzV2sy66+2slapnDfUOowBxVf14lwNsM6BYeaqONy0atpgOjmqb/RUtJdw
NtvkUg8KVxtqZ2YfcqhswYSefToLbstATywgfxkunyEnL/ROEILQGgCttkLMMc0N
ErOxliXZ4JgmAEbimNKxf9s6wHricsdBeu4/zSgrflu2UlBcijIy88qenDkQyKJ0
J9smm0S4IJ7x1wSMNyCB9A6k5M/RmcIDhcxgU77uqGMUIvBTwAZ8cOXcXDUDYYBm
HYRHQdN/9N8spRdaduSGeHmfFNvHSEGgCOXctPO89KghS24dUMy457T0fyxMETgl
pZLs8ED7iEbcgx4bP8z3bnBMKo4fZREWe48Q6elFm4lA6d243U1CiK4KBLSjzgfl
vSj7DAzeZgZOGEhX0RsBzZtuxhHln/Z1jfEFPakvvDavQuAxbTxYbi6Xrbr8Vy3z
IQYQEa2RgHT6txrQOIyCxbCRl6B7c2DKOCbcQk/RQtvjYD8lsyh/zznhH1++GEe+
tG8cv39PDJxoDlv26NbL8SzeWN1vjsVzT6q/VNsBJjJJ9mCQJIARntNyzmWqEVdK
kPwmpqjNwV8cvKL6FzpprLlVyjBwihNB+HdMDvYcx+2FjiIZYg/XauKOtBQBrJLz
ZCcgq05uSQ73DN/k2BV8vn+4UFRNPMxqLTSAiyqgjRdz4MRtFxhfT8WH3hTdHpbV
H5ACnqZhZ2wyM6RrMiFIe6wqtBqyyqEEWvJ2EaWSPYUKI7OoJWhe8bXrUPPzIXfW
Qv7hVOTrP+JBE4Vb7aqtUrRqFeA/NK51oH/4xZjrgKQMo8iYWk0gkXDR6aUyQXG2
QjbFdny4kd6hs0d/K+RFfVYLtZcJWKgeHGhvv0ydjeCWWnmOC74Czv2tr9w9JFZx
7sb6UQTO/pdc2hMsTUvaJ5mGet74cGG5W3RiP+ItCIInqSN2PQrbefTyqQxPomZk
7jOY+0LipyHQoLFV6cKfqkLO6I07poGz31DHVZfCkSb9+Z2pNnbpebG5qvXJtm4x
zVWN4Ol/xVc5uQxW2JilR9tbhwE/aEifdSQmC0UhhWfhPtis4Ec++7dCtaO8uR9f
26CmI3rSWpVm1bCxAAycJWw9oQ1q5AKgaIsJ8ZhpjW6U47bf20szaNdwZNLncTBA
2fydfzBY79vk1KKpYc75OCmSTdVv9WNeTS0bcEtkjfPgJ16Tl7DGNZZmNE8CN29F
qLkJNDzqPC+AKZXgVrDzmyICnL+WC6Vge8I//R2hnpyuU9sV21MU0dZNSQx5jl8b
q3hjNPRwhd8s8lLNBvhxmsKucoiRFfd8IbYEfBMaKaCTPcRl4uZlH5ELDskGsCDB
g3jDhMHhl9mjStAIrFWam9Oro9ek5h6TDBB7Z+1IkcKwRz++jtjwGhUMT8DP8HN/
x+zcmqWlnT6JrHJQR1v/gDftp7m/oT+/PXzgG9ERUcYcOD19PljnDlRG+sVSzSf4
kTDdaVPuY59JXumD3McqIs7Z6SkKD2twHBo4qRqDm/PehSQzkhHM9kW4L/899FPf
NsQc1Pw2F8rF95F0PDRj58dev29QLf5/YYMhqHdQjtnBre4QLo0mRY+HIRh3fJmM
sQODAEJYhksX8uwlpa0p0H+ZuxYWzzENT2+5kvLDiP8M8PQdJNlXVT1Le/CjztaZ
9UPpjDGbtFbIZ/TpDM/ZcF3IWotVLpVdIHGgpeBZEs8K5QANAnLnwmuWtoOh18JY
b7GbR8QxIkZF9buZ89R6zvj33pYl+x8AfHHyrDz2dthYNPYCObyeUdq5ayFxTXSS
kW8clbrunQZ82IoDJTYIyURpSal7EpFP7I7ORN0RapgobQhXUPM6gNFkUtNqVhaI
28yCKERttCLayXsWonnPbbACEUQ9TvZzy4EoWYG/TBmJuic6hA7Ww0fd6A5xh4SA
DExKX5pWXTzsmxQ8q07g78BHH5vfb8KHKiNMSC/C0+nEjbezJ4Xvm1/vv4ud4Czd
2gVKn9eDb1sSYE3+vg6bJSf4phAB8+tO1UqT7IC1+sKAaXDjl55FCKIFWfpj/YoD
q/tDx0XuyEPf1eykjMhkV2RMAHBr4HACeLQORGY7+gIdlP3J6xkk6wbIl38iTcvi
NLzlE+9UUWFdJdNV9QayTk3wEUnwFfspZuYN0ZFGf6uwxHTbnmJoaMkrRzMWaMhd
NQjA2zht93drgAn2uagDz9TJ4K0SRIuEfdKR9d6iS93WPK6083yGHHO/bERLbedC
swQvXxApXH+MuhSEI9hHTQs87ULNMvsJRdp+tAfy3wy7//RuRBKnpFw1PqZ3I99I
1FyozTiHfpfsLSpaFvmktuGp9H6xFO4kytQFgaFi4DrzNFmXOOb5PMbrZpo1h6s1
sLF4nivuOP2CZ58U6EffMMZjXvyYfT0MlpspOTBSW/LPKQg0TB6ipJpEENI0lSjk
jUemqEpIi3FNABsNMdox9lFMSjflLHG+TmlzM9OuiewOSVeiOFw+jv2gq5Eyswqy
qLC5/8aMxSPbErgsvY2czAPJphONbNt1tc+M618VbSn/aJIw4AUtAwIFq4jkHDEC
2y4jN0o9ZzjEC2oyAzSzjSXHs40o1Gg4qZGXSA+J08MHixU338uetF4HsQ0AApEQ
6QRkYUxOCboTHAXCtVn3XqWMTVOv34obMv/y9b+UWOmy9lVAYE7pND2Be8jbE4qR
n60dk7ooYMVEv/G57f8DMVxmZ+zFaJhmlfdvjYeu3taDbo2tP/+XJDVTdwJPpnjg
rgBgDZj4Pxf7RDLvqO2jLD8XoJHOodTWHW7jbZ0qcLnG9M995G7t6s/mt+NNUC8R
3r4Kciv+nAPHdJ4t5uZ0e+3uyq/6ujMlDMt6DPdjYz9S4YnEaRbfj+VDkejr/CId
UAwiiHiU0QX5jM0KZtlpcNM24zJ1+r28esRT9+2f2TTsPG3wc6LqQD1IMwOhvpDq
6OnYwcrioIIo5RfU46HOarTUBXZdc2XfvNBr54zO6lztING807Ifv20eHjpa5XQB
aa4O+nIeZQkumhvrScI4JQXnUhyx5D9mhbXQwPtXp0BFQHO3OaCRezJTFuXgJS0n
Aq5DWZOjBw/oMRJUM0Fxo0DDkwFEknrxbLjrpaAMLDOx2JCfDlC8GdxsHf+orJC2
jqsAZttKIQHQlaSdUq0uFCTJN430b0LsBobeTftp0qcROtmsVRmCu/0eBqHt65uF
BcuaPNhpD8r8jQr69m1In0zuqkUuS+hG4O6NF2uR7ZBc4MCNot15ceuVq/FVX//C
lmPYpGpN4KJ9YomjtaWb618qtxxK0aEA2KK3LWU8WRAyiDNRTdD85HuUPbyo+oG3
ILn00qiXldR8rEIBZYn0n/oTfDTckCvMUjdEpWxnB19zZTYPZBT56XZVXip3xQD0
/+D5FgIPwyWpSP0vzLEPNYBsTH+CzILrSBWrxw2r1GAektLBQpddWbqnE+bVHkAn
j07OS2qL+AUquHbH6Zi3c9HecjRruyhuU9NuziSfYo0QKGcDzhbj32vVZMBrMCW6
yx46pffZvI1unnsIJ6e1J4aYE/aUkzEcBFNjKFEQRLWY0ldlguEYMBHS6rszemaT
sg5o0I3cd031eKIee/r8ZOrJOTcRAmc70T0RKyKaesJFY9tQpjN8Q+M0WDuBApVl
JWmt8PNMsztjoITUTa2aYE98Zo8u6SiL27iK0gpmy7B/MAM79VisMtBi7CV1i0YY
SLvkBL9yh/JBRNnHmSu1JB5dMP+KS0CM6a+I19lZTjSuhr1zXwIYs6BVz3yTwaoA
yN8UimFUTnaHuHLEZus4Ppl6A9mITO6Jz2i7JibBP4X8I5uOyRds1BuIhKFfTI00
pQgRtpmPshtCkdRX5RneliTQhFn4Net1uCmksrgIE0F8sDNFOByptFdHEptdfkaa
eaBY2wTS/CAznrLniJpVeBMimhYWlrWJsyhvnq8iTwzaNP5+rWkppIE09gO8otV6
SPJb44HhNsuu/i3vHLoaXgJ1kb3SNDyvW5rayvFpDz/yIBSaiR2nd/5turnXy3bO
KasIW030WPCCNmN5zXe2x5R9QKwNW2GKRgeSo5PTjaNQyke0ihUw+FXRXhR+4V/p
MO1nvLUe8PmQLeh60so5sZGjqwRSIPIS/8HuCAvMI/SuCTti2YqR/3LJr+e0vklM
FBQJ+HJ72wMBLCoUs7epc8LFefc6sRgYQWiA0WiVWBxPsIBe7uY5AzwcWxJNxAwX
rLjqtVf5B6yGiF8Az2kBjlrHpkmvgK3CLvgwfCEvSHJ8dVUNUGVm3DEMlnKI4AX4
zOHpWoswOIZxskR4PWsLI7kv/wKe0exd1lOUS7/SXT5DUrFupd8x8+vomP1szt8j
htSWwWW/AVCiwnbV+8Vxh0pZQEsIeutEBvXw8uKr+wE+O7Z5KTcGHb9oswP0q1JU
+cVEuUSXwWXXMgeE7SGvulVu7VzE/5b82GNG+Qw7KQlyfXBlJe5q3ih7ptViTfy1
SFv+tXhuNuJdfXiNEb2zYt9ahLmMF52H2I4Vkr0/6R0nemqB8WUGThqepK+Xsjwq
B9c/M3hNHzoeNaDVAoFHTDXKu/QRs7svFktUfbEi6PfyIjrAa9CD9S55+lpaAE2z
t7bqaksKPSzzaAkVFP4KfMhr+X57q4W7+Xhh5oeb6+NUAwDl6CTa1mfd1gPJ9ZR0
nunw1qOc5VJgoPV2AJZV0b5P/QR7zJmQHvdZkiTFPxzkk7VlNBCC6byREMxROo2B
PW/THNe5r69thQwGkUBVN7aSp4DH6mZLAVDcJ1c1DfkDCeN10jgsQeoB8YA2FP7P
cqoINBwIrYBR1n6UU6SEFX52XOKuFnUeb9EPn8XfeCRTUgYa8TutQUEjICemJFYQ
Egy7GmrZ37uzPzTgGhmKJLb0+KaGTxEJXOxQy9WqA89lUysm6ZgKBSNyp+JYa2MC
qR1cLpimVbsyKW1y4kMZK3rKwnA5ha6oWDDR+Fb0XT3leYVmtX6u01mMIg0Qo0k8
BPOROWStnydx4sVOWo82nKes2SDH9mULZjVHqqDp1ngMYwy7isMyhBEh56TT0s0z
M6qVgCos7Tu7AnNDHUFrOYxuTA6/5XnW/xc44rLupoFdAhFsiH4YjSNr5Dj9McIF
VvilW8hExZjdXD76z67Da7T06oUaTbwdTFx9fO1lp4GtqipNAJrbXbENCjoLxxVZ
1yGuvPxLievy90ePd34NdjTmK/UvyD67PV6wVLNyUi8aDQqx/Mg/x0FsE2p8fArK
Eh4n0LhqxP+ww/aOxxfRwQ6hpVZJEU9EzEuDLtPyg+12gVXxAz73hY3nO9EutrPU
/fqDhVeaCJGVvkB9ljayTzip+6cFJCn4vFFbwsqkkyFo/VpDTSPewX1wrzT6qpWH
Irks3f6bo3tuJLvnEA84M4oZjlOndJaYJQ601S0qM6GbBCvZZf+ThU1yEjAYWrFZ
+cOmhgrLiyZnU+di3YBT2wUZk8dSc1vzM3tiDNBQMRK97X8nw/ot0ltWqeknTjBR
Y382Qd5TvJRQlOTpUSQyTaC1CDvTM4j+2GbtNhnh2ty1FJNy0KkWYYLWMRKvIUoa
8h+lguGH95CkqtT1TiSC9p0nQcHbdL54pnO00EvZLfK/Q2Ap3QrT8jCBgCTaceSk
CMjf4C40WV/3UwquO4dEoapeKA9L1NAwAVsbw2bVADsJ/wpXfOX3o7U69robqD+G
qEepr3oEJLwei3NEWQrs13rTvJ9Jeodd6ezMtQ8da+xnLgMStVRj7e4AAYhe0IkA
VEqFI4j6wnZTfxokc8Pb6VMqfcbUZT9+3yxarIwyVUOYMbs9xhUbZVnGMZOXpx3L
DSUGZ11LR61QoL03j+f/06qS34yjovDI6qMjLpr/bJG3syIk2f0Tve2Jt88S/j5w
3pTitU6RbayvOd5lKnK5dIvJcz+xl8/Otd6eaG1B98jWH6svIC0gF+4N8HqJ6YRu
EHhGjJP6oSJpZ0WennOo7p/Kbw4EqY2vRKulwRZAAI2yBfXVqGE3IFqS8ZuOIG+Y
p3PH3wZ6UYB/JvHSKfLVsbjlH+OPs8wOqy7Kcxem4fBoItOeEPs/fiGJHst7ImuW
YrnSBqkLrSNkrSwoSNOBBdP5jHC+qvKZ+L5EG/2OThRjar0CfVZ8UtcVZwqZLdRY
b+zg11B++DHY7MnAyviqGhf19Qn4hBy9U4gj70VwrVpzY/kK7XROM0PDSPr1zPMy
yas7w9zxaj44xri/y2Y5zMX5cPXMYJcBpGy4HSWKnyAN0i8wTyD1/Q9Imo4mS2gI
WDl8OjE+NgoknH6/wofPDYseS4Nukck2gkinWt8Nbe4ezMppHefpWonhcTBr10a2
rXrabFDcRoC/4h37633APyS1bmu+Zo8bni5NwWVE/7n9Ah+LyqZcsNDVb1QGz/3O
ZlwXzbOncXk5AEvhIUrMUrrh/Cjdzwx5aq2cosrNAckqzGhr/IX7WiiFWEvOcU2/
RcEzx0u2D+IZDSNfE+d094wzvwTO5Z19INUIQgbmMMpSBDP0/3BlEwNSIbP4BLd8
0l5PZHoojGY4l9s0pgS32WJ3Sbcp46g5teWy39n4aIE2ptoYzpRkzG4pkifTunkT
BYcvr2d3RkdEct1Z+Ef/+/ydlMzPOsBftyVGZUEpoRUxEtSFjdXJCoXnmuM/QNSv
G2bA0vqpYnEqURw1FSlQbQVGFG7pOkxGUmAot7/a7TxucwGvDu0QJ0XTlW35SKQl
dKCdYmD9kTaVGvRUhNIUL19Gta2rtYXhAlvwz9RyWSwA/IrsJELehs69S2xsbHpJ
ges8svSesJqfRwUP2XA8gvR/rXw910zAZ+jv6qwL49njN74Tn57lpod8x1++QEFB
7ZpNISdQx5OFYJlF/2EDM+C1pGV5Gg5rjiDCFuyiMLoflJ/9MEMjqRDbSbE3paws
J84Ni8oUUuwOMT/ug6kvk2/YyuKGaYoltewdBiatXCVCzWFikeD6QJTCOjsJ1RP1
o37dy4xE3qtLdyaX8KO0cavZOfgfB5rAAgOwXXpJqPfU4R5GD0Tb/57S24ypan4z
M/f3O2GR+Z4yZaDKPygybf2V+S8735whZXOH9um92D+v+fSeRXOHCwg9ADudqdLz
pxbHpRATnQTsnYYG/OJKTUmMzXVCr/aLBEr1KXlSyqhHLzUxwZBUqPST/GuFa0Jx
WuCI4nWoNH6rqBonFZhgPprvKTiLlWHUpH49GKkiwEn8oOZSumntOs2BvrLC+yyV
Nv19bd+/Nha2HNmFnlVK0Ti02slSkjF/2ytezuZ9jNk+q2+68q+VGhTlobr/vpch
UO6GT47P6hGSkF5r4NH9mhWqVTZM0jpJ7IZENT/Am/ts0wzfWRAXvb+jSgvQsYrm
KKLVC29zE7jV2VSaLVxkgAJIMIGX6Zz+a6xN44SYhAeCNZCMVOzDdgaJlIOYvhZZ
R34HMa943KTRGH7Hh4TyBN3iFfLOgumxQk9JPs1GDrXKVsbH3uIERM1Wb+BJ95s+
uFWtGuMMFkM00rMWc9ea1tllT1HxovCcup5ejuIFsxjrtEZFgHd2QoplnV5VyGdF
Z2BUcfPXyPWpZ6caP5yvkjyId7WmD7NIoAFJXpHaUeHTiEiHNjLYq/r4ojKTcckL
qEKwHzlEe23JgBjUV6GQlX4t+bXkCiMVzjTwkSsLzILZfygnjSrLoVaTsQxriQMy
2DSa1as7UNstWM/dKYl8iKx7xZvIcK0ddWRq4qWUxKo6+WA45RFVrnPRtfXBogI4
UPIwiqSh5U0q6TMCvMt5IccTGBcpCQfsZOWFe5X2QHpjwWcy+Jh9JQ6t5kA1sZnD
QikbgOvLfuevTX+Dxvwa+0Z0LNhWvE5w3gWKTVTox9ejHxnWuQy6eoy2VH7V/r11
Cm2bhsPQo1c6y+FSZL3hlZZpJCKe0o+Y0emaYoQ2kNvHIomsDqSK6klCIZ6YDENL
J4NBn9akrBEwTEhBJ8kE4CmVHcEcVTXTwGX6OJSwhH4lnVk6dQ69Yn/8yUKedn2F
q0gwR9Bj2pfCJ1fvWUggCaU5aVhKM5hbnq4xTrCamZOy4tbdvhrlYgE7ARPYxOrc
s9ou3xxajDglAu+2yybMx3FwqWnRSk3Sxc4CqmhglRnEGrtYCep6D0l5XNc6BhTS
bp+Oj8YRDoTHgHuGHi9qwW7BXfNLh2++VbcRv8pd51F+SHLxI/WXdA7jZ2SK3Zsz
j5vgF61YALhtdJln3VCbHPqMHrClu2fvgv6VJqB7qbNqD4BZJxH5ZgtLxKIYosb1
tamwrthI7UBsei6b4JUQ/kQvh87aUfeKyCYZlL2IrKMV1CKuLn0fvI5aTQetJodI
OD10wQH0eSX9VIzhdvCFo+qTDfWxKnX16/ygZtgfAoXxyNKiJb/DHxZmDJlab8ME
g+UDab+wjHc8d1ETIQetZmn358h/pogBLalOu5NnA9TXeW4h1+WG+z+he+9R5Vxn
p72Ht7SwNcTvRiI3Hf7MsacE19UxmJW5g3ut8BuMiSwIp9uz/ucxhYc8Nai+IUCp
FIYGspNaGpk9PShTMm2iT8yxpRQJLGF8yVfWmFNbPN6Pn6YnyS5o9/cPF3nkf2Hh
m5udzovlbOQNaTU6IxM9bKvg0+r/LdbeAfpkKW8JGnmhPkjG+MKdXpOLXoPvaIZO
byIrwGVYp0vtuXpxKsZVH9whFENj8wJriX+4yzwTaoE7u1CdiXHGPBlfb0Wb7y/X
izcfwijQN3AwdC9a7gq9ByCusj0D6X7XbiXAJC94pQs1mIm97/SudL78oK3l0V97
U6Pzt9Sw9aCa0qE47rNPF7MgV+aZ4pAE64zfmdsrnCBKgUVLfoOtY6hFJRIZqUD+
KI3AjRyzRKcJ8EwPkUUGYup0gLPEAFTCjQ9dIiRrkGWd7W0G8y+5Extm5IPVuk3/
A7BJ4MeK6UytsgLxsQd1BOYXO2piA46tZsf47sE+hnjDiwLvpldETlVS2WZBJ+47
ce9AMhfzh/nH9Cfsdst89KDzd/IW7s9ssNK1YpmJcOpIfzS4DamCUerz2DTik39A
l4Fkl/a1agBFDeqmHsDhve/mcASxmD8p5FuXjyruqXv7Hn6ujmwa8uS8zo7Wa32d
POiOJ4UR+FSNv4NxdOg61r2BgV2swFBFuKa8/sJVAWLgSLlLh1bGzBrAhnM+wTAW
DS8cWxGF0QKVXhiew3vOODfsXt2gEq7tKneVbVennd82NA4/qkX843/3h/4pmCCU
U/FP/CkFG4J/seFTDLern8w+xXOvzMm3MrSevNVvKUEw6jp+j1UypP4UJKPpo3Rt
4yIRdXLZQvs40a8Mla1uA+pKqMuBXm0mRiB97Cf62tP6f2Geu4+keZjLVvHZwOdt
ndPTGcSfMJ+d3KXuGaZeF2L+JMN3GQGwZnsfwf02SKHX2dGcfIm8CfVVm/NsRkRv
VebO70AjvntVa9xtmXmocB35qnGxRC1FegRzOkE2Ijd/Nks/V/qM6XfEsda4a41V
VkGX839D4FehrGYXc2czOxrBn+K29UlW6wdehilvT3LIPT37LwhRBuUCeZb3PL68
+C0DzvTuF9tyMKeCoNUujD2uOVhl4xOtqqjZCvVSmDyFyI/89I8rQz16zTQ/l1Nz
cvoph6rHDdngtJI4464/6kiNIrkrFKwSmGgUWYhgWZwLt/gENxdXy/jJfM6i/c6U
zI8mru2Ks5P289O21RjOAe6jRKgVXDfucw+CYCK6KGFfCS9c0SYsUjTyD+ZSVyXs
JERqfVR7fY7Htc4q0F/PDFcthgFcgJFzgtKlhAJk8FlAiNNtc/Y59rS00v3wqJd9
dy8De8jw//Uw/iTyyKnFDN5N3oVYvA/A8AqFiioAyiRDK1193eKMfcytkpA85FL2
67J0ZKu9Hgsr5mo43hXUZJ6k3TLo5T5wj5lv/HCHlMSrptlgazbjrdrbA0ltUYJ6
SB6kK46PI4vKjXJBejwldzDx/aaXRlE0Z0V3J1XtwYekl4L4XwtzCaGcmCIR20z2
VXJzNTM69acMhSg2wbwOMrLPx5B5YEGhi5a7b8gRSgqQj+SAT8Es0ULh0i6/ap7U
UOZSFwk+j2W6tEKgDAv5WLWO89NijVTv8HbGt/7Et45q84OAs48YqO9wSr4HbWbW
Zev/PT4iIAGr8OXktkszqUkrOaAqtZJKOOVatTzFjyvLY5qXo9ETNa4zTY5PFOuz
L4cdc6S7tN6Ur7ajkeovGK5hpusJntS9yiES4cXwY9uvSqdp9xBJGSsAMurNg5Tc
E81R9ciCTKlIgIGGRxbcGGYA95w3+j3FscMiEsV8BZeqtjp3n5UnYc+o/W36plB3
EMsojA0NBG8qnQUELUy5QN2WalRhDlhHR0aVzmK2uwsAJyJ7hjo8kMkci596xAgd
D4Kc8yGphG22Qhth1qppBGnuI7tajeutYpDCozZsk3UttWI6r/EcIu0aCmawTzYn
wXcP6jKRuz+cer5REr5h/tuEMaY6f/Q43iFPGbSedVIwBOKaCag1gOChs+mMAOEe
vChx2yBfFcUz5o8eb8tK51V0mkvDMwpHS3IUfUes+iDgBX1Ht4sicYm9DqxzXcgm
hTLpv733zhZfcmKjt9Q5udVvL/hZQ+l3qPf6WxTqNtalesYE8uuLqR7FW7EUCA5w
ZiLMPTBrFSgBcOn5OligFJqrJwoxjqLlrFice2LGxK1OLzAkIKRTbobhv80RVHyV
OA+0wT93lmNLjBqOxifKlBxGnnhjU9dicWjMYqb9NFK6GLT7eR4F9f3Vmzci3Tur
+2Z32cq/o/BqOK9XmiOjpXt71awqY7VRokbHWb5DNCUCSpgVW9jV5c3ZRpPsm1wG
aBGSvFjN/VfkyqKXgKnC6rSvzjODX3j/lIZiRQpLSjh2sv9KX1MfY388UL+xWjn0
NYm3TZmI6g6QJCeCXN/w64zCQOm3BFP+MsCdRip9TFnYp51yAT+mYdAk7cm7Aam3
BfDSAewN69jSUe2zIwhFQGocojiO6zzywFVh6lpvRn5oOTntWcc4W8Iz5MrYm8+f
ta+aOoHyQlriCyWxV5Ye1olXyes5qE+S7aKvFVtU0+B4yUuGZbQQg+83crvJDK2Z
agV7kFtRzNCsTYYL/OpDliq4bLpxXNfjmnZt8vgqDlAwig2VZh3n5wzFFWbet4XO
HNiKXTj8t/7aRFdHq3nrSLPGWlRrfFN0BYLe/cpEtKyQ25appkUBAvch9i/wMrEd
O+OoI8KhJGeeKsxRuGTPzTaWU5rDJu42Ua5cx5SJEUgN/NwXExpXLfj/CkOKNvfx
a28o3JdFLAGSDcsH252g6kcI358LhHHDLz9Qmj8iY4dfHjElnHQornQ0TWH/EUj8
U4vgCoQwlKTagustQGEnaQGSsjjUsFSuvWJN4COn3dSFo1MOYZHOJrfE7o2XZ7Un
8S6hsTGBgUVJRiR4vQYI4NrvIqKpr5WEGkN4wott4eR+liJW8q6n+9HWSrCLTZE1
u+FVVEXSSv395LZjgv41ea8nnfJlJ9NSBElMdKKV8U6Z5BMAcc2SHTu7WPfZ2VoQ
fl7ovdc9RqQGgefwKmPYJI9rdYPAjoMMebPinBKtXCtxhMYtcsZ4vGoBY+dW+ZTM
SKDVTCggQHRdws52kamGFGnagbF0bzHvsdjWWmPMTzAtJA59fZzDBSxxFzk4zuaY
JvYLCxla0PJmqfaFn4TPxr6aU3QQz7tWD9QfhsVyC4QxYhdDCYbPToYxq7bAtFSh
9Sw0libHZR5p2m82JV6XEocU8rsW8nF4jOPaLxK40iM6bjHkDIm7g7t4hzSselIq
jti9ACmmkBcrSSNAAo+HiGLofOCWnV/tfs66DiY1GpKAKRQXEqamJVjCivF/PJTi
El9BprgVmJ/eTqxup7hPzkbfMMXOp6yqsXCJ5daAiPT85hAVM8NzDc6Qh4ZC/crZ
eBnzJOjElze/jZUFC5DZThcNcZZpYwxOJxl5UxDbJB38PIA8DUTZR9BGBzhQOust
8t4vE+h4m7r768FgloyviMZpk0Uu6oWLoUfi3eL18/Vf9+hoAkJ2LQMDOo7kMtdh
jLFwxkTkG64KwJ0P3T2D7X8I03aRwbPiQcXtDpEFAs8Mfir1Nvkwk6ApAG2ig8c1
Pxhmtw+Tsx4BReP7YbFc0HLbRJP40kafHqOWpqhB6x5HnhfIkdy+hBYvnHqubM2B
mArbPHTZkJbUYH241bUyrS0R1QgPHyIsBPHbejy/KJKDa9CYODRYGK9dKTdmrXd1
OSPnnfSFPNfidzrB66K2tWnYIMuRDoas1wlcW8UUBfEXqosjjR2kucXTRZUD6Jg5
pXJQHVQid6ySoWqof+WAjBYhfaRAw7ddeNydl/TYbTgBIf4upLsuJwpQzzKdXkDc
YEXUPhqZPIopyOdXarRZl9No7ZhOUxNmMjTnEyF+ZukzkG61m5lf9f9rKFUw0zQy
YNowPw1Y/6a0j4javDI+PqncxgwooVRgX2ifiDGPZzWRneijwcq75ERbegt5ABCz
s3zuawNAjXMxTlZn+EypMJt/kRV0OEHuydfxUbXQrvpXwLCbziLY1i91qPvbEWQK
Pwao6STh4dJyOBVlRzMgt6vNIInKeG/NwoPeNKyCK3cIy0UzIvX1nx2a3PjwlldM
++hWfMeIsFyeq94pmUGAHL0PUphmLthEUGZOb6cR8gtfcbDRAY3zdHWv34uRdT05
5XjPTNdw8mTfh30QZyFjKMIV23SbJ4Lsp4bPfSh/Egl3iCRkOQMwBQamd3q/wp4T
jPCNAUG1y+TApL/TXSEdrXnNx2VtKOZ8/F6x9JWEN9UrAs8y5k588EgnkOVfNWpu
wOosKYEmUMf8JybnhupnOGgElI36w8okLHY3Xk1ZIMzbOuj2e6rRQ8Mx2+5JGd5L
TH/Whnk1YcEMv6aY612SIfemjCHE86kEaIB0NQI15nj+La+Id0DOcp0JAt3qzsrI
3enh8hZ4gsBL83aZwrMlDUwq8AKe3zVvMyULp4f0IBoF3ZvdcRiGzXGjRKMf/DYS
qt6T/AKV5OgW2ubRCgeifuTabP/K6Ag/KIZix/JQj21ntYXOe0ZkCfs5715mBZLq
eujuiDOyolaGxn2DRHGkfXF1/6PbSHUbRADH/VSJU+rZKzR6EGsX8kvN0TgRYH10
p36Avint+0zzePZmVqHylW6Gi6qy5PNzNfvvbFLiRawkaE4t0BvfxS2WY+J+apAP
b2FkAbedARW0djW9saT0Q5YYRWaiBezid0jJ1RZj0+JRCJtgv+HH0VcYJsIzzkD7
3cKkCd7pf+kMUI0ZbpkXVCRoK8i25emuUd4SFrD8Ttjesm0kndMRbkeWxHbqod9G
HYhM3bcMWn1TqiOLGJ6W9yzeIXN9Lrgfe1RwYD0PNwDIoE8qrwyv2vfJ9WSu/Xh6
7Zv+gxswQGqWgo4j0iKdKWxc9/8Gi3TCLPaAZuTB6UhA+HBFjLE9Icgv4Z7qLZ8n
Ci8icMlbJnwADSpsyeus+iiOK7teyKKKu/reFqoVqmBBwOVGeDD+R4I8jlL7L+eQ
TtOalQsKk5FE+jgslzjynvo4ATZ/cDm4WE7ktqdgPHM3PJfEtycp08X8qEdTl+uv
r83wzHG4qt98kInT0A74x/Ao02xctJ9U5fP+j/sMVk9OOqh8UltikOEwizSBW4eq
pWTOSxp0BWlkl9kCNKdiPZqdN2RauhPkAagZz7U+YQU5ZK6AZq6fp6axjVkk35wa
fL40t3ol6N5oc9hJinhtntev/+v8zQmf1nuSfEO/yUWa6mVojYOZhWhSzmhJc+MB
HOuAZAOORAxzAwRkfIHuMC50ggka52vvWw9DnRgzp9enXsFX4PyV/dqYxJoMsl9/
AAkMUUi1URrTq0h2eT1TQSHcDUObX4FlCnr5ncQ+SwXdSUcEj1MwBgONiTlJQ2C7
9Xyg7ye8QChN6i3izuqcwqvNsXyYlrpqfaKB4TCU3KLZJ2FfSk/dU0HShP3FvC5V
0B+NQYzDheD5Tkt3xNJj9tm18WYkVgAIN4JTAB2LfHA7CdCB5l9tNR0+FDUzGRKN
wdYYUVK+MOb+OP7+6roW8nNrwHGzlM5UdY9kbvANkz4gH2ays9C21aOBX6cn6v2S
J71ELAa1RfQJ1Xv+l0nwdRQCLrvNRmeCkJZMG1IWo3c1cRD+tkBEkel2j+1V+SEO
ukfX7+UMQKe6dI8sr18/FHMhYY91rqtNyLuhxMlN4RZJ4kyDePk4X1CHfVnBjY1F
kGA+T4VrROo/k5TY8njmxG38QlbZN5uIRHSxPKiZhkN7qmtTGcGH4orhTEk86RAj
IMPYHsoPabGpNyDM/OiaYhLg+VoJKpcdVajqr3efdoOqorTYSJoWA2XCSe8If+zy
VrPiVUsEkcwtuVk0LYS5CVqwV5wZUuC3vZfnDTDE49RWGBKaPqmNFdISo1hyrpPw
ObsqdEz0nFAXpxVCc7YAthlgBtgBpGryID5b6kllw1YCUv0JrYmdgFcb2JfRBB4O
ADvPkcrvOD1X3RhwZvGqROZ3ReKVpJ9S7y0P7k4AEgl5QV/2XjWutvoeAw6WnJ80
rrcfXUl/KT47T2WJXmncxdTskifzg/WV1LHVv9kG9xmwBPFyCSZ4VPpY3Gqjkq2E
4AQni/f0FXBz8AekcOGmm19qf54fabcIpBYzj2fS7U3172t4oLP3INjLklQEXnXx
+5HH/OKHZP35pYoVCeTuQ3REGKjl5FbMnYIXmcaA/hEBfzE12B93Bsg4hs2WLfhk
dudDqqz5VB9rkYI7cdX3kD5A0cX35exAS72QzZ+gxlF4tMRgj2fib4o/Tz1GrmsO
H1TbM1Y5EK6X1/xKjIEzmWh1c4QmoxJiqx5DGIUkgOGyWcCllVLVD1VkkKJuILbg
JmIvRghzQE1gW72AIKtz1t5yFnZHFg0NeeAvG4nplK8dHDh2csyma4ZJvsXZD0/E
8OqD0+daFPHCELNDwwHcP6GVJ4YmP05dHYOlS5www3DhtgfFan2+Ib7OeTfVLtsB
XCvDdkYVUlBGO4QS/M/vtndis/FiddLIUTeA1wsrXG2IjAsPo4oftmckjAL3S1Gf
JidLgplUMQWKmwj5Daf0/19b3XWNPmFUd4/vgqYIYVgcFxGvfrZTxptglwAe0g+k
3Awa5KC58uqXhAQqL/AuB7YqKVjh3qteLaKlDSHBoelxY4FKr63IpKyigdX/58Nd
6Ct4M9uqNcpw6nMdgOzXlQCQ/y6AWG0Qoj7Dcn1iqgKTCNDxI+XaPa/+MoB3DeIy
YZxDBtGY9rcMnsJS3miIab3Y6BcEpArL6X0K+/WKED6/OUOh7dG98SXcrZ5hkw22
YIxRO0NhJ7hJgBeVSAnAJsx8Xa6K18Ez9jE5yCDTkmZv25lsHyScGjXrSbHxcSsl
BN0yKsNFflovRCdZR0RZ8BDkiIgYXuqUAeUkXi2XUtawzwGauYs5beTt/VVpi4F9
BePIVRoBWjiAw2r0DDKyXBFQVfhs5PGeUhNSuS2rZb+UOdRPYyPCHZLKKzETydff
y0Z0NSo8DuIStoJodkgodK2WltqnB56G3VBwoA7VN16pnO/tqSJGgPG7UF/WJWo9
S3k/TrcWwk9M+fnuJpygqryTF75ER6CffhDLArddiI8k9rxRAIULNAhCgeDAB2mB
nM3SdzyC5HyF/YVxaE8dGHoRGiZ+YHfEapH4AjN4nPdUn7CdyND1K5Ii+75EXHGM
T9fWPrHOPZzC8T9G2g+4cviBfJr0PL2ACv5DFKn68RjMujiF9BciMUDDnh61wnZ0
NdV02W0begVZvNdOrFG4WRwMZhfikgJ0e8fp8MLEn3XwsXIR1XXkn22IMR6jjFHP
vj8S79M8kQIraH/73Rsx/rGjMvzntHbbqE+1F4qf7jX+Cil7EcE/nY0ZwSYg9WSg
mfIuMkRMMNjPRxD09Wakn+fU2KPJ5D4/QhGcPMklWLA59atDCjnqrYgGOdAsrPMi
M7JV8E6U1R8OCTs+dWXRmWlB6Sdp32lpgubCvE2YvL/KofjRErYeidPKFFtCwcZo
na4mV38xNdFEaQsvVRvq4oeVCXqpL8SJolpNIsqhE5Ve6bffuAfUKFrii/PLGoow
wTrqzlMDdZNN7o89shBN0F92m3m2fvgEW6Z/U4ZmzjMynylw57YIOCO/avFsvrEI
pit2V/SLz2qfoNppB1GvwzxWEUVdTPBAStsQeq8hD0msGJkmNFRkeip6xlKzVLqT
Ee5E2ibIfgCiPhFSlBMjnLcpGYmAgWj+RmrtJcU6mzIPx0Icz80lH7tBEc9pnQCD
f9aUaAfxwDRRqAnSeWA+T9h+1u+pcqb71zGPURs9EKRVb1au4OWJlZ45L6Svxx4E
V/om/e09gYUKHxj0JhP3HTrs3i1zMtXctuFBLI1AGLPEleMa2qfTO6lL8jUULyoz
tc4wT5uxiOMiO3yUCDDKcgtLunfv8qBv1cRhZeIXhEcEJtV3zXSviMhzX1Z3eGYR
jli5ABJsuuV+Qi/2YFULJPWhC0meKZSANxYmWAAvfd4dpuMTydEypX5cAL6XVKpT
VNybqi5X9EwQI6b4x0Q1ZWH+hEpR0Sft1QoeUyo1OWIftbPsEANanPdEphfGbp5R
oK9lo/tlKdmIHo03RrG5VZYwJ0C1EL0rByxy3SFjpDPcEqySWpHZjYFDBdgIz/+N
DeEi7CaWaLCFCwScqTJUNS6GriXnsrI4+ebhgDOQIBfElGvmIlSkkjOBoN7ZNqmq
UurqTgfoGN0PMGjeD5YUzyQcdmzBexcA1eUjKSy9S8ECmvrDLKpkYGi+PUaHG/W5
6ot+zNBYh2JXT4Ue6VJ9OPTLUzIs8Lm65uZ/mKB/BGEqLLWUWKo/bxkusb61kvmU
ygxFBtkRAA7JZQoIrFAGU8Egr3yZ9NwJlwL0BbX1GTzR8qmXKvS+Vt/LBKs6kKwB
fOpmQEtPjjmZvDYm6iaEU6DuH7T3tou55iDlD82WkKbvECKhGcxMAwlzHN9/VqVr
9e+qucjKjoeSdTCgv3aMhsShF9pAOaVrXBaJur4yuswWXPepFwRuGzBvVPa59Xkc
U5PiZgV3TKad4FXfJN5g4Z+fF6G0wDCY/CLHxXeqtppu3vbuW0QVvuRogfYGEgY0
so/FefYtPb7c4BYRWSWCRnP7/kKotQ5glEYIqLshkUfr/rhlbVQjIJZeVoSPrqAD
HbnnCzh20UhqyLJ+rJBzRof8A7V2svLp+ZGaiBgaTQSBQSIqEVvGV58SmvHehayB
BHHYeHar9JZqdNGh6s/x7IpNwv7O6/0SR3KCZj4Lwr+AnQcPk1/GcNrSWzf6b3ux
OquD2/J6Dewn/2MtFlI434fNoWPqlzIn+GoAfRU8AQcQcPXlx7gZdghNLJaGX3JG
aVW/HL8GfSJWeHEraOwgrIKEOKeVIfv3gyqyzcrcY0aO93eNwrBc3CmRwx0WsOwv
McdcRtzvrLG7RVtZybZ3jZ6qGk3RnxBdl2OuK9Fqqlqq0rmO34rsK2uPFF7yZ2sH
Y7JKUQMZuMUub8CND+oX50W11tCA7qUA+tSNA+ssZNURQff7j5VGPuViGlt1j76R
RoDJw5tYniC4/oaB66UD7VCo/cazdvfm/6YG29BlG8O0pvwxrWGRmkpi3NwoEC+5
z1t0IAaYwr9MSs4sl9uM456s5p+LkNywt3Wvdjt3fDsHiL6JedCYJhyzgq9hdL49
8Hr/0IyzoNhQg3+618/NUQYHn+4zv/OVbrvt249FbiDU7CqKfgLCVVwpgdkNZmBx
avH9Rdot9U+HH3yPIDT+MVw2ctymb3VM8RmNQYqpAGNLQcK0nGGI+EpH96Stgad+
d6poXG6taElPpcYiAeyFFRzA+CCz6m9qIVh4um8cVjhF6jF6pP8NVTZGgQ5h75Wl
bF5aUU9yHcOaQP2e7fuaFQyNvmEjN3EQnNp+/4+T1/zilnzjSBMNw7m82ZReyRYe
MpdvdEucCCl9dRguXiD0Z+twHTgqlMHweE9qC6uvjCgOCvpWcTxsJ3i4JBfRrAlF
LnnkDPpsM++sLqugEz+7Y5V5n629u7bA+p6kSfFA2GtGbHlA200dq1HzuC+yloAO
UM9Pf66oFIS0r5T1dmVWDm7BdaftqkTB04QNXgvoFa9+/IC2vakuNTfP62Whi7kg
RmAT51xPFGyTG19ygtWNDss96KuCgUf3NeUifhDrs9DMe4PFlD8T9x5yiFaPZx8t
Vo+8c+jqaNjgpxhI+CZSGmPAGIjNE0MGz9SEn0Qt+UHkmLgYHZTknGmWWI1nCwLz
KI88Oz0kgm5u4bUqkuiEWz5dktaZ2g/i9yD5dEBvBpIvXWZUPjfWz52A430CFM/q
oVT2b9fNpWavmC7bqpvHJI6jnbBujWCuTjoO/dt8wD9HPlh+iTWSYb1NQkgGy+Gi
E/dqJ4g2R2vnAJ9eOVACqCj6AGiPlvRyWzihkV1vPsKhylgPhGXz4UlGlUsJ+mco
OimWEFVnU11wJmFj6gpYDrXwjRtNL/5AFbPVlPtlgQGazOvhjZUkisYHXVVHR4Yr
aC6WtKDby0sHUlVXhdmj2qoCrxETZluZMYHXJIbUvRWnT6YEE+rlVuxpVaTCbZlR
1NWckBo6qqArDgRdQ+muiDSe3Ppa/96y7GZsXDQghEDY/2ujEZi7ul6xL2dP/Iun
f1uUUVI65x0xkw8NvUYWhD7fhlTXx5OzppgdrITHK/PX8xYv8IverI+2NYst0S4H
LO+pXX9rpT+z/bHCZUVoZwYpMqNTi0fOvNILvkeNV9N7EVJdzy1TI3H5clhfrOUn
KBPzoua39os2BVLVSNmQfqQtnN0ooCwlQ6xVeZjGkFBfHhfWx41oXqz8zrNdMhfA
+WqZ4CqixVwvPsCo7aBOdujzG10lRICjzI3/bF6MDXXhAQAb2cSCeIapdHudhtXb
39WLR41Ks9WkNgO+2SLE7UjhH1BwBvg5mRrD/BVnd8qRrRATaLgX/puqNwIxY2CC
xibDZjuzqEqGjz4+lGAp4brTQVJWrMMvOmJ+mUKyCmE+PShigSfGev5tCbldllyR
ckmIQzdkODbZxkkgjHqaDMH0UHEogiUAGXjbyyValenU4ftDmhOiaiplnp2+xsgS
+wht6s4fuEWNdPrj0bNaY8fsb2VNSeuR+Rz3rhdt44nncOezwrQz2fkINx/V9NyS
gQ2W+jvn+yuZmwp5sPClDzzBZRdGNwU48Kur3mDMH0MF+VV/pmX0QIe3yQM0XHfB
RSyYa9dwN/TIQ+yMGuDRsHk2avCRTWj+atdTo4/GY/pjR9qci8jUSzNBGB7lBdE9
UJ8hPt4Ie6kdujLrAGrQhfQkFE0CuMefUx3VyawHntw8AtgV1o2EAPLW1+5qK0R6
rWGzSHLk+2ZRjCVpCOmCyfZ6Zr9m9g37K3ONVLbv+/j285pKjHQ92DoXGvUW0eyE
KjGqPViy6VgF6K453SFbB/J+UQhBjefMkFkfDgtmCt+O/zg7WGr5I2n8EcNrILt6
Qecj7Cw2NyguzVNYmTP77megD+WLj0HHQVZBymrbqZxPxJVjEp1XBYpmvGO/pFPo
6tyKruFVEfWyfBzUTWolM9Jl9EBoL6bgybNYlx4/G7lDSnRufuo1OsA7J4d1PmAq
YylT4bFFKw+XV2onLo3RwVByQmGSVVNz9MJMCpf4jdBJPy4fLXLwDGLtKOWGIpyQ
cJq8eASpFobDvVHil4xwLsd6u2XkNYSme+pRczWf7V9tk6qx7mH58hborMjWm9O2
re22/QsgEXSei5pR42fC+i+iJHtCpAi9FeHEySixutGLU9o1y61cRP2utPOp15QZ
OSdd57N/UQBPcAWkcM6PT+EXgZu3/7BqinbobdJzbFqcL/z+Di/aH/qolt3OOkzk
Puov71VQeER+gqGEyhWfyitpYZtmpqzRD11aYr/GJcAy+qqstdcpcUmkXGwSL0DL
VWhMm0VLrNU/UaxvAJxeg6mXANDNMs0N9DJmXblLB+74y7fqvk8qNFNoV0NRBlOR
bedSRMJrzT2RHygOv/zrpZQwm4Ieg2ho9i0gTFvh6x/o/oZh+mlhOd9jDuePnmhg
8C3XCiUfCbkwN/SN1SE4Dyg+jLlnJErYuGV55uNcMl1NfLs1rJ41nsJaZO8Cdogr
/3gWaGSfo5U3hESmFU85JG0BWsVKTz/0XFTuYP90wXY2MF4WPQwnSZpLRjPl/DwR
/uyYFZ8UAeW60bJPfutLwj/eO9vcm0X5cLvbWkNMh2sI29iOIJ3/6WYk/N7cTiO2
3el6A0bndtn7CrhIYTu7Hrt+2SQkexclhOilAIiLAcrP98+2KsxQD1nDyrzjLeEt
4BToMwCe6FN1X3GLOrC9On9RUST0lBQC0FdgivNKVhFmIbZSaWDMYmCy385jvevr
NEnLEsyk5PW+p8fqr+4KWOS5rGVfbxeELzDb8N80wM/asYrwnQLAdVpCLcR9/Sq6
bXLdmiHcEdpsB0nZoYmA7eF+VOuhw6F70I3DCnCXYEhTBN16WOWcHdVRu0cze6an
zrYeBBcDq3eqHQJ5OiexBr+Xx1eEL9KOBVrVcB01wHphKT8XDmem9yLrwaphWsnF
T3dDip5Y6lvt+8j7QbcXqXnc/85sYZ36Gad5b/K5BrS0tLMKHHqJ6SV4HxMYc0In
wevpPrvDMuD81i4/iTsV7D3CwsysDP/hJrYwL7oTJzY3927RdaqlIHZKav5d0BhV
FdsBpYg6F4jFFyi4yI3CRfOW3toJDsSGiuPta3rPlI9HAaLazKqltc9ebDhlAqYJ
/QzLDum70PyvApz5heZIRWAoBj3kwutefIKabnVL14voh9qTSr5HGclUMa7JmXBC
zp5xjXl1ekRCG/SR7tC1I1U0XaYs0orHfTaizvQ7ETWl7AB3FOlO3mTqKRSWDoKk
PJljENnJZB1ot6C83bMMh3v2w+sUVa/jgAELpaCBx6TZSNolx/peDFxzxV2YLxRL
imhZzDz0bic656FpORZdC+7ADr3L9BiGtzjMSTr263j6mSqr2l0Lgty5sKD+22Zy
ZnsH+4T8jcmyrGgpE2QLdNw1vgreEAtpFXvfizGdTFuGdDMvMBAEg8bWcQ9MNVCy
NjmMTz6aieOTE9kmlIDQbAh6ogDsn5gpBnAqKlZsYsca6voznJBpiqpNYWe78U2+
1bVoW0BMU66dtcBkPfpFtEEkfEgrGxUgFaTqoujFvt6yjArHwJnYc4MTd7I7i9tO
E01iKhuUP06z1qbZTHKPyx5PFcAAXnezgMnf7ZyWHcPrlReV7GLmFgBCiJ4T/j7l
qLAME1yUb2HDaXthccYIDXi8bpa/bHMxlcrsxok9Qavm7UBNiZNQNkay5yKhvezE
VrCDYRwK6ZVVvuhh7czglb2ZDyWyqnyHV3J6y0/EAHtz7HAWp5XgVS5yLbnyokwV
nC96NyrjYV6mhhJse5hv9gdoj2qMhiUE7iJIWkiPYGZQpgrPSbPm+vHZ8txE0E3o
bu653C36bzEg16L09uFNak/tK9IHFCPLtMirchTtctfTc0UD2nafCeypjPz0wEPo
ev15+ur5iCN1MPpR/C2zTow0+3fpbqhPtN4aHxGsilSKN1imYW3yzOTnXlRS/XuG
47tIfvjoMmjlFH+gc1f4ofd7zslQGkPZX09RGZ8KANUBjRsUKbOkbCXDnvYaXak3
uOYfcia9EkQ1yyvTGlCvqjq/Xvkpoz6bY/fDOHGEpE3pEtUOoHAmuvx6EL9ldY+B
LVtZ/jZtwmjG6+UPdbKToN57TW1Sx0ceKwRku59XE7COO4fdveBQ/zfPAShJA+G7
ljbhrPQTBBWNBffmwyMpYNQp7OjwpoNO6QrRM11ZPv8TI0vtxLIiysjkXq/AaI9w
2y3aV9ovxWzWaCWiE9j3Sv0I/1RtnjdUCKKll7Ai2zmqhIvgHd4dNSaWGIw/fXlK
dbBQwC7ciNuPPBrFbNX7C1xkqByIVRZJI8L4f+tIivSWnXJwdBfiLfzCkfytHvRD
m1sgcAVlWVKmShclBSJd292897DzkkHLcfZ8uu1GdjuY82pgjIOFaJymtEXxFMUy
v3n4tA7uUoNd5HmTMaeKVBSeAohM4Kc0TTwBmV+uBBEWwSgwDTHIDZQedrp9Z3/6
MqmCqU3QphrE2fCFGTDSjCD+p+ncg988gUz0RE9CRCSbrMpE8LMN8ffWNXBLnkEQ
NcMRkgCiGU95l+tjLGXqzvw1pEvtkzrWSkyloGoJHxmRQN1yZ7KosDAgxkYMdMPW
/CvKD0O5IwSDKYmcICzhZ9jM3ztAAbWV4KdAkKy3heY1St5OqcvYg0vT3Bt43sFL
x9INfyyk3Aud2syaBOk1IY+Kgq0D9jCcqx/WWkJ5xVM10mEOewxgX+ihIAu3prS7
QDqAYqdhq1MDVC9GsvZl6iOrsD/COePYGG+QjrdRxPMHdef26IGrEkzLotiv8vXF
r+SxUfMVxXpZZp7Xq0awCEado1xNBEPfUaOybh39F5FV9dS4+2Cq9ecK7PDWQ3F3
0qk5n9aIAIGnop29IAvPUFaiFY3mcHTiPv0iJ3gwiHnoCesgxRSko/MfWdCvd3K+
yDIPAmSp66ee+cuwj+Uoj1FdoIRij8/ZKew/tVpLLK02ljMEJSvoqQWcQfn8cG3S
8o0mZpl2Qzbjw/IJGxiv/EGNAUNlk9BHwfvH9wFWqgn9s2sXKM7yyYPCkn94ysdp
PUoQa+rtGBSlH6UfFc9unrfG82rQ7wWYpuagF0V3pcxDpryqmScaAtAnNax7zqnZ
UdBxVH4K9rWyNOL4ggCMdqo3idZ6AVRr+3udmjKEO5NNvA08mWZKO14VCdI3QfmD
utaFtJZ3GTdjbnjnsAkijvjCcG/CXfnwqZVYhMxkd/9Whb2RPW0qlRIOnOESh5xR
p81kD7YZpweWMluoQooMLy0ZvJKM51t5PCg9ZkA7zAwdEmL7hdrUvycBZ6qhnbvk
jiELItghRcL4wO1SCtDeuOxk/cA8OXmoSJrX/cV3QoW2funzvjt1lG+bKMeroizs
gJgWpXhYFwZCYgH9K10pgG5rYRR2saq8uKn5q4Nd/FVOg3T4ERgbcGGED7Zj8ttT
t2bcq9rh8oCURQOeMQFKc6c5MqZbaKHT/xkj8wQHBkFFl69gXdWEfHWvI+YWmJtA
GI8layOO1jb3U1Tn9oTJpd2p0qDXI2Bs/i6XU6kQ/LMJWYIdcoE+7iOKEUwe2Qf0
o+ioP5HfD36xO1ZfJfC1HBw843GeTh9GY+ty0LNSFxVW8dOJvGK/antvjOEn1tn1
iGwUWEjHZTE6ENihqcQfErNS53a2zQ8Bk6LwnPShxuYnsvl/ScS74dw8cXZamHtd
B5V3of9LfXTcxX+xNMTHnn+nrUQqQKiBASKhG3s31zQV/a8Y05vUkZcJ8iPp0fe/
QY8/nRl/LkWh8a/AJNdBdFPOdY8fGzfWTocbLI3Uy6KbQKIW2yYC0rh0lxyhBDX2
phhbnFgY/K02diQQwX/RaVIV8mzgS4umoPInAkG3BzSKysAk3Gmpkk/rMIvZkWMV
Zm9tJWND/jYnda+ADLVrZsmdX29vV8V7xVRDZGVe8XxavuLaQUXA2aRsEooPPgu1
9BivWsQRhenNEkV9jiRTRlCWQrH5byBogOX5/zqGMtWnFo2JznnQrq6I71wP5uMB
4Iigjw9Vk4o7BoEvIpn//33/ikxaFUAgf69XvmMqnYwFTsUOQTqu31xmZn5vG2CE
hSssn1y657+ODkt5Jy8g03Gm31HqnCEN+00Z3N2w6KU+3xJJTEDWb8RP/opSCqLM
GymNvRx02HXWeyJPstyzbKRoMkcuhabsT3jpQ0qVbL5aCtHpqUiUMrvHwY+JYEIP
gCKCSIpGPd5TeZ9M9RJzjWXaBUnzfB1X+UZBp2dYPhqFffGqbX1Z7u2cSWjlysS0
5Klba1LjfE6s0Zscp/2GfNx1acJOHbDsyIKWV73/da1aZMMJ7TI5ytLRpLn1HW0A
8pwsXFPXoRu9no1OCXrciVviBvR8zyln9ZLVE6F2OjkW3HLaD7C14hXVmaE1OU7z
0DkA9j8rDAL8g+cCdr2pi2CLK07V5Wsvx6ejzer+hjMDXGSKCO2OX8kaZeXsc2Hb
oMDJ0rluFnkTJyH+CrcWUPJQzplm7etpPxFqREgvtaMRx8gqObI43qkUPt4bA4B7
qa0hD163cKAs+KI0Mq7cS3aPyjt25RQ5Izxm/HtQxy3oILx4Tj+luqm7WHzekJWG
mQmTzz8ndT88qW+xHdWz6/DMcdti/ukLvqUuOPeCiICQukARHW7LxFATWhvvcQE8
lFGHgspKXtXSoWYiQAQ4xb+uJ/u9w6vPQxEZ9nnquM/+fVRNaAWiDqOXvMWo6RYl
7vLiYSN0lR94aTWEBF29iqeeoGlDfFEHket6UxNwWqrChDek7T5eggZ/qxLyshg+
nRqdj7ffN/OdeBkLvvCdbFuqTRBKUvY7zC2Z2EFhFPb6mE1C/02Rk6rr2udzl2K2
5HRKJXhfqGbvAvn53M4iKZv47RbMQETN5JjtwgrSN1P5Lb+/YFtP/9gx5C4yqHbI
v+u0GQQLRUW5ptXXvZL0CE4vbUveYKvAClVFP7TjMMa94eLKxPtFIty+cu0FmDSs
xkmSVuAofvG5IAwIKVkyHU1uJl78g7X1boV77X5fnRNhjk3Fev7y5yb9FOpZiIJG
AnvuX2+RMH5UfB+/JMFYc5jqlTl+utY8E3zK8Tf5xz7JLkyT32oOQqhLDsGlMgtK
OQK9JcpDB8ETYhLcZfx7LLRQ+kGtAYEohFihK2fDAU5omo7AEy3d5/NFiSAfFB4j
tZlo9GWzFBaKiEY62VjGMv5nJBscTgqCz9U4PEBOQrlJiWhIj435NiMYTJCN3RIQ
GB/CetlELl9/DmMQ/N4ZaeyiYQWmwoBJp7WinjV0Omgcrvyw2UI8loBbdjb2qFyA
ygyKTo2XiYNcDJApuGx0XQZezFFvjSvA/vxWyQPxirlCsZdjGxO/OfX5eLg00D1Y
2DcC6vTAYil5QvpyjsSqQVZxFWZHE/ozlOF+wsT+X0SFayP1aPhSjN3SndxJyDwt
2AoYryYA90TEM7wY6eEFOLLak5F3MEugxALN0nNzlkgQN1MCyjZ6AMELznyXJTAN
WxJvdNaqXhRvo7w+3/qBibBnFNRgPlF06m6tDutFxs6+nh9sm+je2Jr/6U8v5Zy9
mtDh7reJUdQmyp08p9tBWl509QPA9FZJr2Ouo2FVuK1iCwTX9goZ/rtAAL7noPCX
n3YU67nFxglpqcfiUvIdS8Bsh4knI9uhGYvpZjjlXsXCpc0ty6p0U1BECSAZQJTc
qGa67Z7AIxRoTTfIq/mPhfqxgFZhQSam+o/Mdy5PBTnmewyMrRbzirur4V/rcZUo
t/cfPrcuWTPzKbEbQheG90fh90ApVXch6JeguONl8B8tAGLIU0QOa20xb9RNXIEY
LjKn4PNzIV17fErQxFaZOT9W8OoCOHmW8de4mYx5s4LS3M+T7RXVTgF0hDQp1CxR
t21cw9NEhQjN+BnKHZnujU1HH4HWpJT3vtzsCHL1x/O/tMHDadlZfg/dVtv0UbYf
5N6yBLm1U1KEKMn8VWBwO9TKssUJ+qnWSCYNLed4wdBdjpTidILZSNucuQg+56Z4
LdGZaAGJSHrK1uGRTjvhqjRCeSZmAd4Ujjg7gQ21J8N+OO6LbUxYyLmBwGRGj1BP
tel48fx5KqXckH2KU9bgv6kLsCDoU1YhpVgfaQwmFj8OduIhO57hwdgc5TylkJ+x
3vFR+9pYcKIpkmS2+QUrLFOUoRVCLEGX3HI32+O/gT+XfNbLYCXJg/DDM3ixK5A6
B2uoBDAh2+nT/6qcGV54kdZhDaIN6X+EUCtY4AGmA/gsM5F9l77MCvAyRGH1MWBM
LMXNjiO0O6t6WyCKc2BthVNY8cDFLdoqd382q169yLFu7sWRn3p7pR8ptLJlwkVP
wy1ZjiprsEdgIrotykFOoTb7IIpZ7Bexev5pYliVVmnTUzC6CpaaWYp18eM4yHA4
s2+jyhdk9k/lce13neOgFEFnDmxsjlZiRqPCKSGXrFCteUp5y1wq3EU8QLH9sQSe
yxCgc7PWn5b/5Lh5loYudjJ+TmP/mCG0FipkAMuQoHYwFieah3h/XEyq82lhWLgV
8XkxVPuKPLnKAymW7SV/3VDGyy2SLPZXhUhFd5eEyryst1ST4ifcT18x07T6AkGu
b8p2wgva+bSlYJdRojFb/UNlQA7seMrmnot9NMTdacM92Vb+7s8ET6uj/IxZ9Vke
4aH8c++cKqzNWI3Pxtw/T9hLfBQY9Dk/wVVRGXJLolRRUsGzGipa6hzdi031LAGA
hGicjJsdspD6TEoa98SvKOou8fZ6eNOP+AKwy1dVP6uZGEGvvhGzeflAxKA9h2zk
oAE84FzOWjsqWeslwWHadG+aTtg1RYVXPrRpS/H0b4i4joryjOUTguaDMuRAB2gb
tVdyFagdZvPEGIBU8fWrrWEAeGAzXrd12YV3oQI54rJlQ05cVmfnwfe0jeoRPj+s
DdgyMq6W8ZXWsCZ1ufWhgCf0XVlYcivKb0SU4lVxVgt6KPNgTQ8Wq/4sCy8mdGkW
vhEvwaFqdJl7OedJ3h2imvugK/0sy5J2PHIYy2ZQKurnnxsSDzjvm535fKMkKy21
f7hcVW6WjgG2vEXhD1jY3Tp5Y3Tu8Bwx91H6bOEsrXr0Juw3c17Tq1Xv7EFIq4rh
nZBJZ3wZJLgwEZged8K4sZ4BYb7xcmMUZPIAZIXZev1CuY2iTOnNSn5UlFKUbyAq
LBka1UNkjksNe+G8/z+xFBrFmscmH7O2BVGqKyWtIxYg50EW3ihhf4CRpyhjfek7
9H7VINx+VZhWOC1uct1SZBXQkBXpuct7tleTvS5ieRXDKB0RE2x4440h7NmrcsVp
4vJNG/ZAwNJEvrjPuCGtld1qcMnOhtrZToFj6KUXG0YAB0B6gaeUMiWcEYnk68jk
U/DVC2jAq3FzhlECElH7yePEeALbsetzPO35H81TB5UPK/CwW7wcx4pJzW5uB1Rz
DNqD231UaCBEcxoKlBNow24K67bmPZJi0t4bk7urh4w401B6Qv+QYq9IciePPRNE
hHa079uL05K89a8cdABOLjdOyESEQNJURmtuYeeeZBfIgebVcOmp9DAdY8kwkSJ8
vuz18TPyXDtQAAtBaSWW3PPqmW7cKTdzUfuH+FlmpimLs8hlIUjxSg6aNKyBoZmg
JJY30uBbZjpQ5Li57J0Pg5Mge4i7bqFgL8WgRHLbKK2UuraHUZUbDo5/q6p/0ARu
2XpN+vsoUeL1L6hXjobL4cXjiLMzGkaWyhUJ3y7KGOa69nO40O5RkBfUqR3TqN3f
vsHvXy3Z4eB7Zp673feACqGEmpOOwnEqn+YpXf4qXsBUAQm2yuVCSdH+XQ7qsBZe
D4JCAqe5sZ5rMbTcuW+Tc8/yGWvSINGhsrUTFZ/lV8sCRP8ug8WzWFHiU8JdMSgW
VIkl5Tj9jh9XwJAXelKMOUL7Q2XhGRZD0SpPJOwMp5C21V0tMyvlsjq6bo9tQ+Jy
IXGZ3tnLN0XaJSuaRwn4Z9vyH7fjislAM+6rSBg5MfXsJW7G7yyiYgi9aGpDEEQr
wVF7eyjDHmHjUzXEgjIHdu0y9iLI7zPqFh6lRIKcp0anC4efqG+9M7UrTHObDIUl
/yXHgZWL524eqlDtL2so3HWm+VbwuZF9tP2Lc+/7V9SFrH3hGq3uTV8NXVmyqYSm
ulGeir035jOdhkBSeyTK6MTS32oZpB1eWe1p8/wR8f/uVbGpKkoOTZqOVkvWUrsv
HG4lpwOsHE2k6QfBGEBI628Ed/uSXl4w9ka8q/N6J48XOgoVelqhZMxOLyTn5iII
C94tx7S7M5jRWTQqCV6NpFb3zcfFyYwfM1ggdbka3E0GRKe/Ud705gJMLQUUpiFp
8qWt9WFTUwXaMm0+bZSbp++eOschGWxAfOuP7jwghhT5fSVu26AlYy8OhP5JURLm
qAfbxVIAv5BCRJ18N1X7aoDf4jaKdG/4pF7fMG+Ra3A8ufrax0RxlS3kLoStB3t7
5Ln2JitJXR1EzMUlmpXBzi8gPD5N6tnhgO0ig6FA7Uaq5QLWy2W2xjlQew5CKbLt
BCivN3jkIsKumdrNpedR1td8TeCWDoHEB9Hvcm63kWvUPxe4qDcGndBSvkQlQukf
k47lEjny79qIN0e87kMG/WOziO1gggNKpTKgGieqUcypyJHaRvFNTNuLtxtBQkoZ
0W1g/19FcFJAr+3z4weZJ5mJx2G40I1k8FkEPnrakXhPGp5ad33RPwASav+k/aC4
t+Mh2iSN34+DX+tA6+2dpLV7IL0V7QRii/c2MlZKC+UHPIlMHyVJ9+CSsVAx4JUj
SBUy0DvmNqAFop3VC3u397Vdw48rcSJlMdnVxDiFThS22vflU+JpCht2I1rlAqto
P3FW8HlePx+eBd0MMctFM6xLT3rUW/l24acEnfXfkxWh9/Qd7rd75I9qyL5Jt4sk
GJTAWvVTdXNPHvvrrrrCUddP7pH6FyyFsIwOwIrYbjsqgQDxXSMpRkU52fc6dAQ8
8r6bIUJZOn+mZnOjzDumnSnkVs1Ees8FpRKHb03UmGSPz4pbj+KLCKPU061QK5ML
XyPiGHtu4s+gB18ZEe2c9CFxnxcxPhVJJbRUlDwd+9ZvxiJ9KmeTwCp/36X17TOO
NCi1tZn4RBneubOch2G9Gp8IO2MPCkDQZdF0Ebtqc1MQKwwQvbf9n75WgjXf0mzI
6nxa0wU8p5E44Te9aD0vZgZhrNtvg6bcXL1psbkRkNDjKyN457LuJqMbkK6VU2JR
4ZAwcNh1VvvTxbWkfILAgwi5FaakgcY/Juwob5g3FL0jYgI1/a9KjslS9WXlPnEa
VSkMuheXeNrV8oCyxfZ1ckEaBlm+tBG+owVDVHPJ91nPkZ/NUeb/CRKJ2AFjR6LZ
HsgHphuwc0d10VdptLMbVZlJ8Zn1w1rMmOohX5/W2nIgwmrx1OrD3MJhe3PJDctd
1x17KYGfaQdziyQAhZZACN/axzKF8v9isALzeqUDe2vGvpVC58AXw7cqGfjrUCvD
KcwUyqt32iVS/Z9ivepFxIa+hTWqaT4/2BYWHqwNQCEUSEClAscEGrCVhMrqUH5Z
pD1agT3r+mCcVxo0j/BiinDRSWxBoEkQQLGaTudyoX85zI2nOj8u/4bg2B9hkZPe
+WszRBJZ9JKJfHSBgFFVf8PUoXXXFz//TIbQIzMM7FwOQ+/H+HFbz+gcQikSj1vG
Ad/8jnrgXYlzQeYn6eNLaoX0zKo172eJjm3484emsATzrWbgAiJMTaF2rgGo9dbP
a/T2ECWAnVyD1rBtI35I1oa6+jA5ZtGQShDq7rG7HncYbVoLKohqY1drwFWhUchF
I1VcXGs63ywB/rimDtwU4bQ3Uaxu1ZQVFCpAricR8t3UIi742K+A30vZshmGHzw6
Z1RWJppwOwK/xjbdzpsYz7t54xobLJFAwSkvU27glwp2sEpSZcDbCkLoQFHX32zA
eeo2AoNV5zPYax86UPi1oFID4NhwVtiKWf15wJwy9jZnVwZ7HSMe8bAMoJFWwr+6
HDJudmDZ+wmErBnYw06Zw7tQxOWP/Q5CT4ogag2NYYIH6x6rWmMMu67+C7DfT7d5
Vo55jyk1xBJ5HnaJbSCs+yfGRmIDVEI2h4Hle7J+X9fqhVFQNO+ANIhXTZaJo19J
iP2rSO95iO3Giu4Nm7G9sjYASQhTJ1GGcfLpBlaPyEnXLHMQ0Ezvnu2Kot9semBu
Ob4LtJNYgcbC13vf3TLH6A+Ce1jYJMF2GFwDiQiO4BATjiYG6sFd9wfFZ9GRoyTB
acDSJiCelYyvnv2uVU+3u2i8HyTG3rzOwqnx148QDENnt845rudcI7TKa0XW23xz
WDJwWjXQrLpVo419Derkp6B7Lqhr663whXmGg65mxaxFWvAgAM8sacADwQW8rNO8
M8hwYIeRNScQfSzMZ45WK87XrqDrcWP0pIZoDG9+ClYPhXP1i0pNjyBeQSq6IfJI
W28w6nQMIRNvFY8D0XlL6CO9uBXlg2yrUGOM6ySQh1sm6B6+KRgIuMzGGXxG/uWE
aN5fORhtdxuTs2cxRTTwosKG5ffC8PwrZeLtWS7ejDBRggsPqxRundN3bnJMeViS
c4hO2D31V7E8ioNOFqOk29z+bmhuIsWQJqjwcn3lQ9iUsZMMB1oJtun3r8ie3/A6
xXNggZwDqy9AVIUKJnR6SClM9b54FKt5SofHDgp193cMcxCRNqR7hK2yqK3VrzJS
+A9cIMQWBBKXjEIhPsaP8bCoHvtuAsAlutun6zzrPgc1XOnPrpRhfD1Pkqz2EMPB
QQwKLZOQiZYH9WZ0rIGg3K4lnqr/vMea7ottWJ4yL0kpIZkZdOAlZeevIhXLJt8w
G0WqzBPuRAvQbCmYn4qm+6Z3aQAzRW5crc4hlEFM4T90XGXh7dldhGPoU+DxAkuP
9dZvJ6n8AdoHC9l0LjK2Vzes6pKT97pzxVWm4L9PIxQ2HeyTtVhDT9oNXFwKMkbr
gnUe9XdmgA4n8LmqzCUeII2lJLRvgI+/m1eJfSjj4tOxahwHZzNHHfWCMVUQKXAz
4K+JAaXcOj09pVBp6HmsIr1doTaVo5UrOToxy1TanM8gg2BgP8EqlwCxNIELKN1P
zIqPApDpF+6v/6USkQwV53ZgxGm+yqYMxc25Tvp3tzsnz4YhXzZJ0vGhuxVCUF4n
spiGCFYKYaNPHoEqe5qPM3IIz5M0ctl0WlqKs9rYESnUF2C0mJiGF+l6Yp5wicJ0
ghmkhqt0oZLUXu+OBxAJSFVcuuQoizMHbgaqvQoJ9Qqmo0umP0bNDgGk1c3KsoVU
W7t/IijUUqv9fJ8Q2Zh8RNK2reSLJwr0Y1/iQCeoN0fW8Jne/f07/qqMGaMsUuq3
I0CgHopufyhifOWGCVvyYxhyfxlbe3GtmH2JqOHofR8avApTXDOe2pqjLG4Fnk8z
1bRERo9zUUv9YUEv+tF2Pvmf/05cRU+B0U1cEz09BozTsnOIQHiVFlsx6bu0m/b2
COBmE0BlnOf7v7496M5WIqk3JbtN+QIoom4b8clU0nLCH8ypkVr/pqfgLaNlA6LR
oe6+U50bhqYTEoEKzsmyE3nNs6DkMLKojEa8NrzwFg3kTYDcwaCdLbBULnrcGCBy
5OUIdnEqkLfS1LNOMyWpytwnOgmgTUFhhOfwiML+QovozeIIWDUstdKbGLYHfHt8
bGlAXEbFHl31CpIXBqFKWO+RnUSQ/KMLqWq1KfPMEhS5GQGzWj7UAP746HSvWgDn
01mxOyBPfG4nRlC3IsItba8CDY8d+Qn924+VPkKacJOXT+jKylFTfhqTX6aAMlo4
fWpSS1K9t4DbTPJ7O1uU8RmkH2OSzAGioD6YbbLeV84GWszB5WYtmK7WsdYMGoq+
RP+h/FZVOXwaAZ92Hd3Qu1OocIrzepwR7Yaa3O9Y9OmVrvITPrUU8hS3jTYjgGjw
D9EA9lIlexm67EaiG4TXRVv6zgLKGcePNaMkxS0KN86RImiwtSxuZEJ+cPLwauzZ
6QEVnjUDyRqxQaLd7/7r+pfNgfOnofXmu8dUc7HGFFIAnVOH/mKSNDljRf+xFarY
D5f9qs3vSt/NAr5Pdw1QBpUbsldDHaXREl4M7sRyWqugoqy8OGpex4b0L79aKAzJ
VbEw0908j+VMtW3s5OUQFzZnb+gGA+53obgEFOJul64Ap8qQpK7zmalW4u9uyZe5
ddgVjlgoBKf0hdYEnCvfxFJGnnGCobQO+WVh/94DgsOmjdEhMnR0q1Q74XS/an1+
QxVZ4zppFy6d63bSt6p0h/pimoVwzPI8I25GdniLbA4ttyj7HVYAuV6MseB5NZnj
ly2Q9v0oc1HTHLvlnLCnzBkPXjPe5YI6VxctLGL7ief8F0i/pxlruWpZFUiMFmEv
Wy6I8Gqhq0RU+s+l/hLWTeyP3oBd9SuVc/RcOW5qek7omc/RBMQySQoQxJbsyS1g
IYMBAyfEkTANUt2jqJXdu8+2q+Z9EJ6MDI4j4Mg/LdjrGI9ST05ZA/3O38y8g6s/
jHfJr2E6lvdldjhDatWDk45UwQeXaQYCJP/8+1Ai0skJBqfqx9y17uudapokXP6x
eQY6MZE7Gm/w8ML2ySJfCHngboaiRAp85VibKHUVUk5H/5j5YFviqUBjEUSDbQoe
BxL1SoAgfFl1BAHGEKzsCADBvp6Ws0O+vtQOFogVCWMnVGaUSVcc0Pg9dWh6P925
qRc+Me4DIfUIc14GBolunB+Jm70gCN1vEcCDZOBkiODUaZLqz+ntainb1WaljrvV
x9GlELYWupanlQEaUcINlb9eW4DFAlGTfu1lZkTnCaE+r22Mx/svJ38uEueI8fcx
9D748rq2m0M4BVuDiRV1uRwVFGViNesxda+/PAkXMWPphqkMp/f/miT1Rmd7PSb9
WC9AnR9by+4vseQiUyA5O+t/vYRkme7MBD1zjvqNMPQjpTF2ZlbzXv00ONcgsxRf
jtq4WAQWQo6h/8j836ez5m/SzUGxPDkbmF4yR3Qz45ZMhndhjdU8xgT3rV10QFt1
SDdFLAMsg+LX9Ehkjg5DSq0yy2Vxi2Hp0EbjkNd4tzS2NgZNuGeI9v2dUvGd0MEq
u4gOS7bMNl8Fq2U9lyEaFYJnTvBxrpxAlI8kJKt9A4Q8cQBqNahECmmuVX8BQCsT
/c28nDpaeVqUoGVkuYJ+SLxLItclmhAKONS4YgBmCySSnn0BiqrX+czq7L33xyvL
qcTW192YzTN87r5ctsjZ7Msb4tYD6SeeKbb7eMtAr+zIypmklMucid1ff9cG5jx1
Glnw/TGTa2tGsKWHQFunhfBUFwbXQaQn5zZj4hPse6GlP/cwPT5HmBkSwyknFuse
QNYdejZJFM/2ghFRqDEs8zUeD+Bhw0+K98x4sG3dGA8jUWiI2H1uHrQgUSBe00JE
F5fQX6/Z5o/y5zpH6HSSo8C/E7Z8L8TNMFYTS+htbhVK47sOSgffE/UvoQRjTYa0
3coIWFVW1lH8cYBAaRegvrSFLftGJPZuhZgj0YdHlknZxIr2rpuPG67S43aXbnOs
qL91+AealV08e56VTQ2zOATnu7i58xmcl/IiF8PuWv7sLcVtsTknaK/U9Yn78RDk
tX3qRL34yrOE+ERe4mFjYx/lQVMnbEjvTpxItBKTBDpyeoqmtjdL4Gkc8Z3cXbIh
9jyxtFLdbJsRIMczUs1REQ25H9R7KhZz59d8rrw1NIl2Oz+APOs/kJn0C3S3jbbQ
9QvX4lyrK/XuSnZzVNdhngQ/twIP0/DM3kf/ewYzhoZ53dWK4yXfteQh+66/WzfR
o/i7WNg1YjasaPjvSMmi8Go1+adt598L5u2/0Kw/TSoy5UY6uGMMzhEtt3mFGgbb
NmDFjEvMC/nNcK2UgNK/VB3nqYe9ZTJ9dycw/qgntjA2iBlTNGM3hwYbNacAg6uG
lted3uy+vDKkOBFSTAfSZTM/kXkAQ/a3F+GeWLSjhJRga5zCcNEl9vLfd15/Wxyf
qU1mlpqg4J6TwcTqENDvBEw1Sg1qKcX0YGxBcl0GtQXvXzHgnupN9Zp5VOt7UfhA
4Z7ACVHbOXtvOtzs883UtMHA8y8PyBij/srjS+KqpZ2bgj1dzfMNwvsoCAGBzl/y
45CO3owhwn3WxBeNemKasXYf+FH+3m1FE6v9cckEa88QkR6BYCRojjIekqPdl3dL
ojHODsKNCZ7DsuodmjwMFJzF7nrBPuIsFJ0ES0GB/swSfUBodDVCnoQfdCowCwCg
1r4/L3rPfpyJqEMQ8Ve5PGbqLDm0R8sW2/0AKBESwMcxyr7kSo7KdT6urwh2AKel
7SWnHI37eNVfQftxXE+/64oOgaG/cpdCal/s0WTMtm/KJIozZsKhrhiKTagKybev
FPglvmLhcrcXZOFtP1uqg8HBAwd6Tg8eXHHnExlpkyKslehxvWOHUfpYflzKMEZB
zJEoA9cqMQZHO4W91nTYbvalL6/0UW/H1JXJz6TfDFNQk9Vs5SGRrwm6D4L6EKBW
szHNPzEknqtZru5GLGViFn4tEQc2Y9PZ94ufgGQAJ994aN/t4qplrQ9rpWVRpemQ
RRxWjCjBkmDTjIOg9WrSg1H0cu7RsvW9IA5+Dj36enqLDtYUAxiVcgNAKX5jnrpq
qFFL8ERLqYc1XK993lpP2r9hxAQJMYB5o0/4mezXxJmiQJZs8QAWJTpahkZ50ICf
nhHLbaOcF4/q6Fm7TbLT0GTkGMqpmZavKpDBdh8rp5hWcQ4FDTVjT8cL9N9JxEMq
njSPcNRmL+5gCgSxKSO78TqUQhXWyXmUpGU8dvzx/ReRYL7zhZJKr1PrKoi2oHbv
L4C8sziwIYxh4hIjRBNnY6h5zyoGeDx7OgNGzBfbXeQR0tUqJx6FGiU3w+0kTXJI
8UD5wyRxpRnvfIlN8b5FWyhb1+rxCC1Ct2Qv67ICBTPNsl7zxQWL6lmOrV7kfCDk
g+0K68vTvkfpA3gMk8iaVx0koGQb0t4qG7aUZKr+topTi7Tji95cZi4asAfsEAib
eUQPaBvudJaaxirAYIVDl3F4Pr1ywoH20YHr5v3UoSU1igybtkiWFZRF/eIeiQ+y
gKCIyDAWwZtMCvn55XQgcqkqZuk1MDsnXwOshmEhk97WFB8btCpdJf0op9D3z+sc
OqqGo1RWTz5TI2AABiMjGMouvLdWp9kqI/wCiF6JVCX2/jXG7/jPY9BBylDxi7lt
N6QXAmE5KjQ3YHQ0w2Yy1pgdMHAmeh485QDBmalQXH4pyv/Nutp0Co1J86cP7uQ+
IlMlO6hGEBXK5ojujPYvUBRZrS6/cYqKzc3LCJjwgG+VQfAB+NCrXUVc0HyxFQPj
FMF/9pJgHCK+sSQBfPmPHjcCR+Hf/AIYnmsacukFLCuow9nLsIiHWbYZZpjheM+S
Uu1jR0EjNzgOmDG5uMc4yjxRl7txvfjPqEGkHMmrk+0eDnez4CytdRmC29ckOc1K
i1J2t37wPd3+L/7dF/IMCMIQItpNxme3exZJSzcc6sNL55Wx+17n0C+Y0OeyVSd/
ALGA3ANmFzufc6TQKiv374IqBDr2qv39z3yJCLcBzt8hPTpAXO5+AUX1024YqEJY
TbgzLA2qsmTMWscoViWs339SYecBfq/zbXu0gVYutr8w9XijeNPTV+BM+7BdRO/O
YbDdtXBgZR0nQMUiEKKtfdHj5SdrSifn6oHLtA62yAB6Aqp4HJaL6pIffs1gzOMw
GekWIUudahWaKVqK+oaIvWwjiKfpMB6aMyizcU2SKMhzrL6iP5lSEQXhGArNR+0o
neHGZydV9MkO5PeTClxfJUQrIdDI/Myxhif1h02njQydX7/oCHdMwsYnUwTSv4hb
5SAxtIOiDKWeIuj2M5gfIhdBSBnP/oRYAINAnpmYwYqT+yhobjYbFcdbuI9w29c2
8OPlJFJl+5q0pX0JGe6PcuLvhgCyQeWUJDr9veMnTXs/ZCmd6rqprUu+nm7yrVC7
Ccur82NyGsRrufAWM4g+xfKddQSQc7pcbXY5AtnActgZrUtEnboZiEFUVSic4wqs
5lhfa4wKyE9pd0PdpCCdctJLWyrkED1fpandTEyyBuV8FYeX04rfGWZdSvx+5ZIR
06HvFP9oTH3X/CeMg8kZxHDpI8mNAzip6Qmh7qeZLGhSbbFidFutpu3Oy7FcJotT
q/OvPru54Pb9odiZALI+xfdG6kJLBsbhcxAUYflOqNuuC+R9v6beXz5hiVJixaVM
3USUZ231Wk8/h+P0SZkrr8vVPAOB9Jk1R4fFSVv/lZM5xYKSIc7+s934TmnxrF8W
nh4iAYvf/oOmP7Jd3efrPXTupzPmrGHwhe3FX3veFJpStunRftHm5hEpSmBT6QsX
S66yHKhu/56nOPIdA9QIsXYoMjqPKFzBr3mH1UHms55zY1jI0CMxkFgZ4VQcSEiK
ZZE3QIYPVCGraG8hSWvqJ/3/SYuzTbN/S+EJh4sQJK7GuBghEQm0xfQSs/GmLQhU
lv/B+VTGrs4yAp+QwX2joxBZUyWLgffoc4Ec+DDAOGkTP9s7XOJWBaHUGTtnhQin
+O1xqnb+HpKTdd+ZmwqHy6uVSZLQoOqUiofpqitQM2SZAfQ4yr4nuMD4MiSMy4iP
r4bWnaw/irsZg7wGU54FO9/D111xN54rtlni0Apjz2JUGjiDZgNOrb1tskstYhJu
e+otToRlMLOMpLar6HU5y5iPbwqkdnbNHbVvkE46iYsxfOZkMbfVm5AHN+SZ31sE
AFfdHBWN49S4hkKnchb0v3gCr8o9suClQcv6JyzbSw5IPQR/K3dYHH/6mk/eTqqt
KcaZX6hY7lyOgU65QI21xd7hnG9fj05fN5+C/6F0IBwhSEdEnkGEBo/vxtD9xh85
L4VrNiTOiJR53b29iFj7J8OVmVFLUKjJDeYC6XP260dSNMju5Y0InL690Un8bwXV
pgD5U8/FQahtmWq+JNrCmD4E3oGldrC4hWIT+PWjBI1wIfaKa8k/cEGXdqXxWnOi
ocfgGBeFu4W9j8tG+fRnqY7N/zZgtftC/wPjFswyfYll9+uBICqu3a8dABwLOsbY
zy8bbvny8Hr91WBGqDyZt2b3ur1lLkBnve5HWZOE6rGrbjJW/Du+biKb8+Lyc303
7fNqUjvVr+4d4U1etRhIMXUr0KC74Bkxz+jx9YC9AgrQU4S7R0d/j6cC5/agVLyL
rCTBvrKvRya5yt0RbNdYpyUdHx/LF0AzA5LcQJ2h7Ab/wB54HumFoHwHpcxUo+7p
nAdVNF24PaClobAgBUGBFzAbBXRArZrQA5SVYmCm7wTyroMIJmyS5Tld3aPPs8Hh
9pD3twB/K76Gu9jtj+8ZqoRjrbxzC0XmVR4LBtOmgzy3gp23LndpfFPD4YiOI+gG
ZOuuNg08v654U7Z2Y3mjxgLoyL2TZRrcw5lbPqX2Px94Jp3pYAf1my+98y5rfTRP
N6D/DIje/T0Uk9a60lt4fM40yOquV3dbDKHLoCtTbnI906go9vMhwa04jRHmh+6q
19ktXvprWanhMfRGq/hXSzFt9VJmF+gUFdSfgaoAi7yAk8c47PSNobqzzMlzu2Dl
5eD6y2pFOLoAvC4SBzsRmHBk/MYPU1bHSTs1Slms3rgg3WgaaBC6OAmwNsIuhjPt
/E0eybHuOJBOUOujE13TLqqd4Jjk0KJMPNwEj12NIzLuHTWOTQM+Cyr1TOB0XsRE
pkyBYRhp99N3jVZPBqd0QOH+Z51KPEAjZ9It4kbVO5YNH0zf/fia88ITYCzdv5E1
yTKDAUKRQQiUh7JWTD2R9OfIwBvFJ9HsucyurzVKI5YcK2KHOYEjGAoJdxMI944y
GHvXBaWe+CckJ8mO5RR2RgDwaGVTUs79CiYflE4SjkTgbAr9H9cs9c+GnusN/yP2
bXx+kKmgzWAjbZlLbjaQko1nSJAdqiQkASa69UgAPuKXLjMe2kxkSciRLdcj3gRY
/ihWnKqpDeqDd/IA0eKiKuqOtcVesRmb0g2wc6AsOmMu7vtgBsUuKU26qxZtQHGr
jTYFjtsBVZAlXW8SNZ2jYnh2Sx44go//1jgZud4iifgBdSA6nhX1yKINcII4fP/C
jftWhgp6Gy5kSkv+/qyYeYc+EJ8W1+/lJDKC0WSWHXLMf/WcEqV2UApLseAM3oi4
Z3dGF/rBsnAlpxKuXV62jqtQVRC80+gaHsmBl6CzsWCmLg+5r9seQE8Z3gbxL5ry
hVjjIDoDRBaxZUawo5f0kbd6dZBtbWiTNz3SGzykTfoDArIXpneJRkR/jBE7/mVD
vy4uWctDYLOkXpxk/Z01RWl6opUk5W4mJozz8k7XPLJk+4kWvcBvZ5lir15MG44G
IDLlJpf8olV1HABvRmzD+/voaV/JBsk1jctkPmFck2aSCHOggMz7nE/J3ZoiBPnL
Ul+4oOdGdNQI86/nTdogLizjlqGxbpOlGS7S4Jk0/b/hX1r72Sy/dq5cMOIU7tFg
MnciO4zixf6dS+KUv5J2ZuCVrWJRrdPBXRC1KSIkCQm2d0931I42UjRD8DDjR0WS
+41TQ0MjpFCyXZJtdkfeyKCkDiQW47zaqox0+IhZtDL/AAxDA01mACNlc20r8AAq
VBho3daan+TYPlVjsLGf/HQcy4SK4osblDwB3PZ1pZAz5cqrHBvzNZ0f9bXn88h6
8AzvPFDEnKzZtxWa8e6EojTXt2Yawr0w6B/lOLcWi9ejPPxnb027KCQ8TOqMZCuS
m/AsA/XBOY1Wp9aKSYJnlptQI89Hwl8pWN9nmpfv9L6VEmBtM9p10HebS8PqUZlF
ZvudUIKJT2+i818Q4XulItd39BkOIwxPh05XxtsQ5fJ6Spt2l+Hipe72yGisDTdL
/2CYk+gUORkF289OFGh8cYb8Hse5jmkuDR3wt3+bI6ZEZPJjIm1BjOwjFY/xElNg
ivYLCJt0lJYiwx9pItPu1NAZvOl8OowxlI6d1ONeqwptM8ChgukiOFu/jA3Nfjr1
r7Ug2L7SDBpticOlU+U6EAwd5qfPlJPZ+81yUakaS/v/qH8llRmmVIToxm3dgrPT
gcCjAbNXyTW/EoiEm9BgTEh3l2qzt9Bo1rfUfJF0AfkYPp+ZhBLHJcPRe4NAq8Z5
oPE1iQYJaUaJFajxfdpXo4kEJteXL+FZOd/F0j7YgOz8VXXnT2xkipNjVIdRVjtY
V2fSH/bMl780D1oQj+6fXZbLAm4tunTQEdAs4/9a//cIkjXTiEAgiQsppyzDHPRK
JFvudhDimo6AXF0/HO6yM4yOLpamJYMfF5oFdkReCGPnMhB8z0NSupygs3ZA/ug3
urKKcFM5x9txAvzPLe5Sx+WoqV/QLSKDYu4mMTVaFGlude9JeWKeGD1ckutYs5kS
nGga/wW/PFAyiugw/6tinYsw9i1zw+Q+YgiO2DHlbasB/kSsYXCdTZdzhXYAlFJD
yVZHh9bHhqwl+ZWEChZFKQskBpGQiTMgYBn+GpxgjBX85PKwhzI1CDRhvtGSXZrG
YCqQRYdGOvJgJpmUj5NUz7T7umdU+T6eTvj8sKVXrnNpyFS1vRxyNUMJksWdEGzh
1ZAAYYoQmU9vW5gcKViaVnu06W6HL86qMDK39rCNzi1Bqr8KFoQBUCs2ziC4cd56
2b8hQ1hLzog3roURnf07GjB06/MsYxed9KvlWOiEAydEdS99wsy8mBGUHUjXlMMv
ezY+cPHhlV8V3F4Pm1JP56bYEKHq5Bw9ENyFeV49iDCkamVkJcKHdJAyZZY81/GY
3WUcqkEojMy/HxV6KKz+/tVBdjfMLN3CbEVnB7JMtnALihiiMlQqTlZQSZKt/hR2
i30kWTWPV9TU6cKBq7D13ztDbMOPnbWmPQ+IEOOIkivdZPxM958TvEyDX3Ns9Kcs
U3fjsB/yK+8PUaD/7gUY26eWCsjXTQ9rBgtOQdqR4JMv70gmH3iU1CBQmgblWIbV
I9DNbO+9ys6baoDhSDiAo45eBFsyL8V+kNjZtQ0EqLLwudj5houX2g1VIUNKOnwK
d3rkoddU++pRdd+9kmW7e1hoPBdm0Q+1wl5QdvockLPZyDjcY/Tn8hBNGGo8lJXI
dajGQgSS5BTHofmp1F1j4fTzSZPu/O4CukRsVZsmdeFVlqvtEaUS578KIYTe3Rat
7areZDeSh9Ety3EFHKICdf6Gjh0jX92XdRtxeHktikLtQxophaYcVSNg9k2i6jtd
uGs9qmPYIJJYubDB8/jE5igK768eSn5CGmj5SMw+999f28rVRuOYLBKaqf2dwV1H
0QO1cYHVX86nuCVvUE8vOdI4XKUt/49raEAR/hZICurpdxS5Z5ca7eHw/PDKSi7W
cNCgvZeml77Eh26R7KIEfXex0ihDXVzVXSGDTpqW2uCpcgK9wNpq1H1ufGmeDj0/
0fxAMTS64JBfWKs7HyX/DorXhsRiQEV78N+wOYkOrO475B1hLagsIvYIyOcmSizf
5lggdoWhzFizsYCxgrz31xVCZfr8hMM/tv3x1FxtyCc7tjkTS9yovzOJbVkdREp0
s7jsM1CjUCXkwX0mkkqZ0jWPshZ7a3a8z6AWlkx4ukfH5TP8sE3sLBPVP33QJjKr
Y2awfVlTWPkr4wsLSXRl5vj1W2gtrBqBKPVBpY6QXtXnSoZC4CnymuVZZI7+xNIl
OJweJbNqnBymtScnCDylpP8g9a0Oh9xwX5a0BAD5xxq80ZdliaKVX8UushAODgba
Rk0x5iqHVL2SkMUOEP0pVAK00C5/lONQqdzAawzPmEoH3CBW8wIuWuQfy6BYBo2V
t3BrvZqT2RrJy5uSHhQ8/E/FqTLXrtE6hDSxAVCNOHKwIorwDUX/gTCqwVCguEHH
qd7P6T0HnkGysteOczciex6iL01s61OPJ8LbBmuhd6fc1hVPUBBiU2/7sSn2wjJN
3w3oa5lCcBL7dFdh1BdCQT4JcrqlHeha+lr1MMWsv2/W5SBnX16K+HrB0tYb6a2E
EtZrwnN9x+c4i8TUGfEMy8FkAgcNDGs6Q0Xzfd+c/WM4YmY4mDKaWhE8oXliLtGY
0P2JKQvSK26fqRIt7Q1hhHsxgV4pMOykuTXjReVoFdST3Pieph23L3tLDBqBg8nn
TssJ97VLasMv33yjzN7QoWdpaWTgpRV4OnDkKJkzEwx12S5us6rh9QL3u+cJcH8y
U/otJBS0KkBIMuuGOlI7uYUBHa0GLuUBZHT7rA5erY8pk2X0nowTeq1nQtfv+CD0
TsT0HyK7q3pctXWXogP02VF0feXTBNtl+51EWHIXZJo64iptF8TD8N7HTwu8YxaK
hEIWxkcWAw1Ina9nx0+gPhT2/0ZD+lCd3hqVrL0jzW7BpcFP3en+i9dPK+PknZ/O
FxWnkfgeejQ+vkTfY2WESynfouRtSFjyBLHPfZQnfQBfKw+ud6PfFAQLhGkMjPoc
DadbOHEMJo98boIl5+h4dnur5ruW8Von6mlMRvfCD8efrX0NlBe/ePTn2RCLj36l
TGf5W6MP27qFJenzQt7/zGgffYefMxN69Nf9AR9HlW2hOkEyuPwKiioh1y/38fUr
KS47RjeOpJTCVrg+NRvRFcO/i+7tMU619Kcv3Ogb55u0puGy+Lx0w2wdbSPZ6xiF
HJs0m9J+QVLeAjotL8QbjdBLXvHiuOlWpSRY6AL2VNyAjJ45PMSxFW0ipbMa/sIL
Qqw16ZHJa1wP5JTZchm9Q+7DoDPmTJBbX79+Z4+S3lfNhdidDgA9EvHmCbykNdZq
PL8HlxvU6Xi8CHlMG1suNMrV0JIKDPz6ZaCS4b84woNHEuWkBlbj6cFJRzigF87f
JxazknJwtJzF0jYjb360r/dfSUaM5Uxt+EmjbPwEpmAJaPwGtddTWcWefwJUc5+L
bLhQH0lud/LiBuJbzZ6pHjUtz19dioAP2yfQKCgxVKkLoZnFinuz278a1RpcHccI
wsZKeUZKKQ5PzLLqCwI8Zdir23EQFQVCeU/qM3963B2Bw86KHp2+MDfltgm1h0b5
QNIgHpv2PwIQC11gyhXGuz1PELGTiB1oPgXvBWvA9SBzhRPSb+pjM4RHy0qLUZk0
VSUW7y3pYZNPJjhXaC8K0Y59cT4NZF0YL09en1f5t6s0BAubMlwAMzdXuoQ7Gy2P
F8zzbpE3qQex266WRk+IhCNO9Wccf5P1Uw9MR8uoL1C7aapTZa9S2bgtZwT3EF5a
fmm/tZTuPZQJnbUqC1xLaTrkt+Fu29OKGhCiIMSauTWuOgFHJR54SziEJT4W0geV
JEM1cH5WuEUiqq9vqoNIvT/hpYuh6k8+Qxi4tWN272iVPNtKAD/Cs7fpsI3oFtYo
tc0KW47jbNlVN90908X2FO+9JcUUmOYswyHrJ2BmjoXXpM6GyZpN7x1ij13FtCTU
sYhHVFNdPbPDl+iwcesiZey4/hsq/DJhSu0B3m+Vj7hLAFTQf+U4hbU09vLKmP24
SrE+rh6c0KnSuQ63x6+kVe8VzPYkByatlvMu+bRDzykW8S4LhINJ2EJTLi+TLvDj
ja7IVcsfbhp2H5OSbYeXaSd/0xmfad1oKvy2+9ylhw4ABz1Hz/mzN5GLuLs1Kl17
RLYJTx7tzSdQu6Zf/3I8wQNkCA1mWi/8wzojZ9pk4XkvuxOLwLwPuH12ULqmSbVp
jPQegQsQPxjqtyhRGsBx5t+mlZ+TCkqSz2N+jnTHX2EwHrXmUldNJOURg41JW5iu
ceQWCogyzYb7OwNET1C4f+wV1k51sM2gb7p4RBSL64F1LxkYTLDL04DnexwgVP+p
mAJMLGeunhLQPuIR2GLyOa4wGIRBH1K6LF3ZP1BobTsvPBuLvC6YrOLxxuI2q40C
Xkk8NjA7S6xendCztD5V78pJOcH9DXEs7RtLZ3VKabNdexbCEPqFtraLNl+yTMm+
n2cW7U/48DvTVdgnWSk/bsVrAsm5wPuOsMQbN4qRCGoLBhqaHSkW2HcgNN4HehG9
eGgfr/OuaGdv9saMZ5E1wDoWuzCqp1Q9MrJ0ewNgb3dBAZrM0AU+atqYg1Y4bc3o
9UI2MJtUeKsJFY/YMca3K6QD9fkHZAXKGoo8CyU1WhClT8gVwQLwP5VtdBov2SsD
9kvdveVQvsOMbNdeGaBIGuQ4YfeVuVuGmS3hxO68G3gUW2CJ7jsxA2x6V59+LFyf
tGo3lOGAxoczObPODRLKP8So/0+BexEQ4vlhHlmrdMGiMVa5+QZ4H4PMxQLCZm15
wGair8tWU4Gc3pSMxMr1Sp1UEppeMsfaNB4AuF7b4/28y8Qe6gD6wN8zZvsMwL1K
+0awkVYTY/p+4EROKTQaKtNN6UzXVxOQUqLTUnvCELojYdWSBPkfx3oI2VGlxLJK
ALdL4i1Y5DsKjYHL+uY4Qhmwe2anlSl3ad9BN13qNHhgjWAAGYsZ/4RCKVLznp+Q
gX6Q+ypRkjg9U+FEDMAH1aLr9eX1Z5tnuhi6GaK8SZV33F3O3VCPFtP+JhyR6+22
DW5+q23BbrLdnOhYqFKAf8fJoLTje3Q1OULxdN2A5kl5IhqjUUxtU0gkZ+guDN/f
COOLyubX4tjn4PyPSYVkw159CHY0vHM4t1h7e/4ufrddgt5tegGLMRC7aw9znFFl
xfdM4La9NXwZfWDvAusm62c5uP6o8Px6muY2QfCWFZ+x58bIsbl888zcF+KJz0QR
55dLCXJkz2G1LjaOXP2eLgjYmX0Xify1XkMrdYuj+AjZcUxRx28RFTAl9xaX9+Tp
rFf24R5dEjDJSjmC4nKo1L+5dh1zq5hdt0z08gu851bkMZRqFaL5GjfROWPVhpcl
8Hd4KbxPUBgHRLuPX1Ir8kwJ/vBeWLYzo+RSAbGJEOEHUAOthNxt1mReMbZPl6H0
DY+aB3QAyuIuCpwxrZi1K+MN3JwPDPJQHgQlTyynjhDkRmNEgP65A3f05zHPU1Gs
OZ4g7yoo5lZlojzfKGSGkYd3xaFliTdJEGRNVXNtH3pImRSin8b44Af1jgamHoyW
ahJnYTniLttCdLpJMasVtkubo+cZ8lpEHfTWAeGPRBOenvISQ/e616OWRCWZZMbc
LP0llItw1llCU6ufbELbIczMfSNqgc/vx3deEQwi8qprDGpyc+9SpDeshDdif8+8
jy/6l4ayUaJb2Xlq5B1Ho5zsjKLTqyPx/kG7n1sK+bJCGYfC//NreDlc/b4+BniF
O/PI33C0EcR6KsNLD2ydQDuh1KXC4eU09tHRBjl/gnIMJZoIoappLw95GNchDmVC
iQzFTWLoMpyIt14AK3mVGpv07wTIN+gbXCr9lM+2aaHuJipiEYAfvAsZ2j9nTPmZ
gl/3NZQIO+IWhejDohD+fYK2KwTnOyTp0MFpADv7bApJjCcrtKPBJ9+M9IHWIG2L
2x8+jcMXsGXV5LWf5XI1UgFSPD/EO4Pxwc/q612Kgj58EVA8iTQAFU/bs08KUD/Q
GRPnq9sCgDryrF2iURjIrx885PtIfgZmHTc+SqOl+hpkl1sfP6iY4RZN8xJHd6wq
JXScBbOrdeRP0nVhQWgTnAsXqgyJJUmFfYoNDiAbJEXxq07jW8NJYQe6AjRMakij
D0tclDIwja25YxvTLPR9Gsk/HeZv8lZ5guKkCd0CS4BmJ8qFHVSLg+496imsFZni
EIOUGDhYOn9ZNOiIhXgaOQjgV4FiUnSI3lAhix15QvJkfkpmF6tqpDliaFvw4EXY
0oIWrqsyJyQeF8lSFXdU6+NXukPT3CLl7El8K8Co5Oiz+mlTVfXb9Dqm0URYITqg
u2tWr24Qi4BPJYnun+4jIfEoWps6GkyNjZVhfND756uSp4P6gQe83g1bLpeFZvCD
Z1OwQedVOj4X4W0EVelnWa8HPTKVxqTOeVoPhWo6AMRjhfX+XX+5LvUfq/zgFcpV
gMTwuL1GYc3iwkq8gxHUePOaYUrbUdc4DWW0F8x6oJJUtNgLCm0hjlEj71oBnYz5
H8qc8GTuWmKjVmCYNtSGDFjugjUpioF9B1frlnR1YCSVEa9mDl4OdjFQ12xnn19y
hwksI0BmxJb36obFn29M14zko/yUOT5YsW4YcXRHMxSuz17nyXNMVETQCWIuLPI+
aIyYMtgxsoveCgqiCaTxTEoEMiZVRVl8qIH1hIBZSufPb3oZXSC/r4a04LzFEO4q
juXth4OVPJyIIETU8Jt17uPzYvSA6xIdUvrKqz+G+q0sDr17fvET8atutWAvmZfP
l3ntBGP9dYI3RnZKF0kaZfNj+hbqORyL0TbtZ1bFiENZAp8a9bXdndTJAJksqn/a
IKzrFf99YMj2OXl2zkwv+9Ajn/N8CMHJKwitoRddhn50mTt9e9Nh52vn6Ywjo+HU
yLYNgBhGVSViiHW6eUQ6CguXAmOMrxzhQWtg2/C6o4xUn8zp7kUWzpo4jIaHacAM
ofNo/2Lyg9jRkDL4AUs4p9d6END9pNqqAJYUvauqtXoZQwWJJCR6atsUsTlzTuxs
Hy+FoUl5as55rc0DzSOv3nI22n+LJTj6O2I4cKQB7Js2hH294xPC/T9r2pegwfdC
obj1xsIizQzuksbPQ30IUQih/zKhrMD415IBzhL8R8MtXrWN51YnyHxPaJQsiZAD
UrkQrckVezGNLqqSIH7ENFZYH18hk/nCOK3WfRsA/3cmqBWlnkgAsydEf9+v3o21
DhriOU1K6kMlrKui6uK2qcCUnINN8ref+o0f1Vu1YekPtSPEvoWXANyS63wYEiTF
ixSrUYSlOHMHCnMQmN0/tWl4Hia+ZPko+lUYBNtCI0X5JI0JlKHF1ZkkJYBmQK6A
Msra1Ty0WMUMr2qYVHWeJwOiA298CVgpT6d/1+TmCnRwCfcV37AfQMMDSiPTJkhR
MhKYUuaCej6IWpKkTL3vDpOKTfLnqGYcFbuenasVN/3Sw48hjsBPoGA83cUQ9SJZ
1r/86BSu0WjbDbOIO0RIDmZNA2gJdG4tcuc1O8/2/GWZVc5g6yMh0JNqBnkVcOmN
uityHMt8Qp6pMNXnHUdxEI+cy5HwyRdfVYYOSvHFQeUl9/3IPcmlr312m0k+fgS+
aVkNV3SJasa/Fmyp0AeBKlJD4yQChH0CS19l8GINO6yXisfvu0y19IpTjHssDKFA
J3CytM4AmOEmWRvL6xihgpU7zLqd4aRXqGfiL6pt+mt0U28dYP4ZMojrOYsKtZzP
0nt0hWmHgqSUUMextha3uoBPSFUGyLKUMtYF3Ea5sGSIVJNry8vgCu7igulq1Rac
qmksdSpZO3tYwn4MtN3owLiLLLMMoJp8U9bE2Gxdm1wje4IHGhE+s2l1TeiCM+5o
Ubo+X2yKIjf/YzyrKPIzahRoH/BWz2BIBGFHH5D9Owq+czGb4Sba0ip+FreLVGma
JLQ8cNjLSCwaeTOD4xUDGVXy1KokdiZWqCKyM61QNwuhu2jPrd7rd2hgKAWYgbsI
dOvVropeWmDbVMdxZuYXHnnf5X/gUAjrT5v9MSVGPzEgJhHok28xmii5gKpcVPCf
AroQmFov5hxsiJAiMYt5S8ATncIfk6wX8O4/m39Q+/2Q7PvqYjxdim77draFikY0
EE83xjTMi85HNQNlwrMdQzfhUXuRwVZO2ymYp18kOgpAjDocPdYyHBfRZbU34bTn
qqxDv3ODOx42lmj21Ufzf4dezf8xAwRUn0mnuRAggTppUxxa9WmhjH4OqqsEhqiY
DvoY12FfalWfEydU9oO2Wk3emGyFpFYjVVJ9mjosAHg97Cc/neeinoWhZmEyzoc5
GoKVa6nClXFbJgM8SliTEIJJXVEKuYCtgcWncu9PWjT/SnXZ1em6iuY/UVgwqkp6
KAr9ADOCP5Wfh7ecZ+eu/SBlqcY9nkne9zXvVnypNvAslc+CAbUzi4I8XTOrrUHM
ESgEBSs5YIezqSR60TTPR9J6wVRWbd6l43GEOwssKct0fVss73pGNRyoWYyEPFwx
+KrskazT1VC6/YO0vqtVfvF22pnuYV3h6yLrcqv0GZYUidWqHD67pLYQwHC9HK65
eh0WV1uRs6NrmeW3y2UyiqjEaa/8ZNti5sP3YdU5ZOitedPcOJlCOSt+b68boyba
4ZbpJzilIIBpmBoxk8nT5EyVlqQ7ISnSwLtHrL2Si+juKNpOAV1wjnuy4wulQJ6C
+vRIjxYM4o59tPLWzlNHHbzvMfng3L3heW+6oSWwyJ6SiOP8VXYl+harjSzWUK0/
VBAiQvyvvCXhsP8wSxt6EFvpFrcssxzUM0BZFefV0CRfF2WDE8vZkGLVgkdzzExw
0z4R+mMCOLqz5i5RHdeLkJ3M1bAW/HcruEoy04XE6bmT3TbOriyNyCyj1Ss/i8gb
BAEiYvQXLW4VI+8APn86BTRwGlE3pMVyQuDCO+pU/tcHpgZPasC+Uy/ukAQzARQg
yq78oY5OOIzVcKZOOXZZVThMRZA0l6O8l1wpcwUJETQYl8vRO31/4x9BQgjq84sf
ph3ohvIhSKJfss36S7yYbQhNOWxJv59KJ82Oaae8YIBZQ+Nfv0eeMJXlezovTsbu
z1L0MgUIFdjdtZmfN9RmjrEl66JzI1M9MGM4KyuStBXyT9NNVk7p5q5Os6TRTYbF
7WTJMZEDbH0CPiUcOGoKphhoDG6UIMMv4/u2iB5fzImw6gBuDz/mO4CBkGrvDVyw
bWlyFw8qFjeyBFi33/JDWtSxHz4sNS+kj7oFIqaG3aGtnP/kxzsZSpZaY/aC1XFu
E6aHvYPlajyAnABSrMbay5BdiGam2cdboYrALrM7wTg5uwalVtxKH6QJRf8oet6j
s+Adn2yttnFR+1ZnNz3SpYk3z1H0ffKZV9bqeml0NPtjPP2V+sO+RmKv38rWK9Fv
a2JcVYKZCcr4X/phJSgP56GixQtPnujt7QNNn3ALR15z04Fv61E4dhgBZP9m8LuS
BbuTXlLjNfXCBR9qrGxF8PRqE7P5PC5xagA+7air6+OuPsZRCM42/IeS6A5WEC6M
B/gQQ4etfKeJC0Ls98JRpc0o+e5gK2YsRVGrD08Dn92bNkmgZddyth4wUL3O3MVV
2MlqXfZEsiQnpTTJwJHkqILFr8tC3ilU15i6dyxdzCAwPal6GMoGx3YOXJS5ouwM
0ax0LBnkD4Sj3J7dWeEa2Q3R9yUejDBCXrIOo7QM8K+MqG0EBSlGf/M540mlJEjD
S2CmXLeIHHeZ8sLBmqXT/QNCMuOeSwJ+mVNwfepDYh4Id2QUoDaKAgm/q9PnrKZA
PalvHkiRB+MKBaht5YsNyPk2c7NKf401JQLrjV1CyEN5DE4pVzGQL7YEH7hWBkyw
RCwmbmntmzV73mN7ujm14cPU4uHAHyK0dr9eA8/FzCdykgvmbDnpZKR3xXtMxcrS
0wo6HlvLyA6Blc9NWiyn6zKMGl2biwFl8/+LhGQ7YG43iaJWc12wKiHfdz3z8C/e
PbXXC94v3pHSmRMGDPlfxhncRGRh972pTWRSQ8BfOUiI3b9RfpeCcFYXXnnUgthz
RrK9sHAvx6xzI5yHgPDURLNLCZ7TVm++DCpejO3w3q0qZuLspThwoagI6T9sx/32
pap+azfeDLiBP6gHRY4no77ez3aN+mqlnDucGKEPQIDpjnbpmuTMnptbvH8Wwhzg
W7/Sl9rFG1ruBaTqAuJvpGxK1E3b6sDAHQ9VXaGVHhNoPnCsSJUKwHm1txQJxVhC
Zp8Q4udLz7K8lOel1P2F3LeUIfj2ql/DPURjHxtiK1wROo7eQPGlEycB5Z0pqnpF
9J3+NRPowm5ri1/iX7P56C1WgwdSpbi18OY4N8twA58MfHGOs5cKET1KlqNCoJ7w
qh2OpoL60vUKimKU1GhH4wFh0/ZOIYCRudFAjsPPqUJWEeFjm2sH1z4aj7665znY
/nL+muxBtd7qoj4qWBkHTYJVLvHKY3HEK99Gl3agPKOwk+FsfCVn5brmtw/ePD1B
lir5BG4IECsxkR6gyHq4/nPKnMImPaXYDJ2ofSxFPG/8wMGQdmLouQ955M4Wy9Ps
1UrlEkF/K7aBiVo8QLgIMkfHKtnN2NStM9peZHrRN6SoJ2p2Nokb/+EwsbdlGduM
zMIz92PXcys9D+om+evN/Pboc3ZYak8VaEMO7uSYVwf9vI26TGOyD3hDZiEfvTAM
6XG0OPGgYc8RHYSoqdq6tuogezBfSRbufhBqYf0Pr2P/F1GpcNrcHlOKJapOkM0G
ONXBkye0DuMx00utrmIM1fkToABAMwO8CJ/tcRRGvvVzKHd5YjGkuZzAz23XsSm4
LF5F34sw5ybFv33C2Svzqs8OFAVRQqhmkfcteoATqsUuuQlR2v/2abx177uin3+i
W7aWRm71PSM8T24dXQnpGleZJmH8KsptMOsMubulBWDTqKfXOj7rN3vFEv+mPUb3
CAmpa/fc3M6i9GDmAFsB7p+JJFn4mEY0v65KA5rNu1tr+3H1LaJqbBQCJWRHluoJ
Z1iB1DSJnzmWc7mbSjTiMkcDdFUtrpKBuVOWu4+K+Z6Dh5eu1St7gJrWBn+Mv9ut
kEAIMYh/iLUXq3JlADFuaDXnVU/HWLG1CwZtSJ9yOJc47OJcVc+7445idSfDmI1Y
e5MxEYZlypQK0PHBjjI9Z2z5FlhkpiuGFpVdqTaw9cQIeyuUFZ5ZnqdfMpxNeQfM
iynwzxDUXmsm4dUkkryRW0Tuu5AixOlya7ik+CUnZ7iO7qeRtmJMRXbTv3M22k9q
U8axLzsdDTjLAghODN231Afy7cLWHEoYF0Ou1ioavP2A/zAV5VQpPBQm3A0Ut3Ey
XuHx0ykbrKtSztmLEzbpNbRBXre1I28DMjV1VFJ6GD7N99JLq9SyZS10JCbX3jQH
qGJHhHWECXBl7FyHThj4zZ9H9WUDCFNMGNVWXcF1AxSbHHxzcHQ4PUgicxvJkLCO
h4VMVWhKDOT/w/Ba/nFfI+e8bh45xta3tqE5MvVBN/ixNcdomQuQppZHz5z+G/7B
q7fSLff2Xv5A7dco5awjusu0zu9eswfIEv0JB5BYWNr+Ff8+eDUfRz7omULoh/GZ
fetgRCZeUl+CtOFxakNyslGn/D7DuXtYSkaUsiWExa7yUeq2FJyc4AUsR8/mXvc5
HKSaxrYSn5gD5eQ5AhcBHqFer5GzyY0J/edLmikr4/JS/tMyTDryMj3AF/4n7Ca2
0Qx+e4AnygjZDQIXTCxs2ZtotgvUpm/397r+g9NN0STvjaP0B/mEqDkzpIwGtjtr
6FeKo8lEuw8i3Yi11oOuEbrCnxfbFwYg+yFFT78+rvw2oxIZmokWy0z3fhqFb0YF
0wHDiXhxIj7Iw1b2CqKtuooPn0rvDMhn7GAmQW7UPw5z+ck9KMFpNsknzdXGUnPR
f9UcdgQpjcif/1TcWDkmMex5hRxjEVCNDTQ92+9WIl2LtbS/00L+jNSgs67C+hAI
+SIAHgjLc6Nsx2tNwxts7NaaSp4rvj4l42xh+9ZgVg3+yXhV75XqMsxJmTA1qAwW
ndahVpNvIbF7jI780sBnElNhGGcb/mW/RxjK4aLq+02M5ixLOrTQcfXhrw4dncKy
yghi31DiUtGdQv4NGP5yR3g/ff5RahI8fZaJZ+mJHIsNi5Wrgdor5untzeuA06zR
fm1UVmjnwAVcCH2tIokPA4p1oLG0ZPhsNtHtORhPgNj8Q2ams4RdGCu0JmaQprLv
F6tm4HRWLdHTTV2zxhzPHB6fG+SiEclRkBpk7xRZSNQW2U83K+M1+CiiCWbkfLk/
zgG7AoNnWkfUy2sgnUyPUBkaTRCX+Kr1Fzkim9rZWeR/ifEdXdh6F5Y2YJASGFXI
Egi6vkJVitcLnXCTZVrq6lId2qVXKyq5S7bmHOm20vNwR30E3ZicooVvWQCqWdzb
w4A+AWn30wPt6vu2frepppAxDWt8mTN36+QHPWAAPH/X89GxpMkNCVrNvHOwtolK
vfQHVyIGEUNrSNWynHSWaTtWXfLQxVyVt5Hf5wnYmBplRokAfQrRacJqET9VCnjU
HFFwUovW1dGFDbc1KfYHYYY3jqzUWYdCIli52sBVlQIbYgaEKxslnv5ltxYqiY/c
99TnNrE3o+JMP9zrd0Dpyh2fUFkZgmy/CfrLabF8L+zVUVYjZKpwTGcuFZ+pcHle
iEzhondHJ7oHQuIltRaMWDgIQbE5/4nn3aG4DMk/wOtgwJM7hvcc68yDLLZSe4Ph
gHuAudpASIdy1n07lsX/dCOuqyw7YEttw9a+Jv20rh+xwLAHCqHGfB9PqjE6hDkt
DgRGRjZxiEflgzP38ERuucw0B7R7PIzhP1eU450CQtnIP5rgk/xkdD5vdvEw30yn
C9ZxDsfxzMg4iLY1HGJ3AvwafMFh7h4gDXkiWtX78d0iOPf2TICezVx3h08+Od+4
RgXjNut70aMEpctwwWf5xJsEjLaRU5hX9dTQKsG0xJHJ8kDNJ/SD9ml0fvphnVaT
uX16sYjoxNK7OuV3GBeJ7f/2QLVVlh8RcTogj9QKVZCxH5M+qjA4B2AxxKAcNb8n
P0Ij4PZawA1An458rx+cM0BQAJeKrxf4cidEcdEUzcPC3VZJVae7NM5uAKW+IOST
6Sto8XRb4XZDJQr3hBO6BCKYUDrwFvdr9zbyJRoKOz6hJY1NaCbyWdnIqEmsaXXP
yooiqh8wg8k9QnwlF43ajvg0QFdqaMoCsnjlD3DqYSrKxXKLtRlXNU3xB2v+2Wsx
zMh33bxca6KwFoZVBItkKe3B/E3yzaQAgVR5u+/QEr+j/Cd1eYlDdtD/8c321UtU
os/AG9s+7ECMhR28VcDOaKczvk5jBTGfWG8L49HUBa7KW1YtpsCLVNg92i7o8hCj
Ib9tfrAUC+2pVaFc4USf0vmI6IjGYdB2v+CcSJgXkfnspmr2yz8ddwh6Ve4aHktz
8QHArFKvG2RR/zzZpPlvtHs4DlDPyUgH1RqmrFMWC8ypu59MF4Rj4kU2azU+mffk
t2O1Z9S09QnaVkRFEkhsyekyNp0HG7tOkQL7nrS7Zpm5AOYaxQNP1OOcEeM+Qntw
qUy0uJl7OjEbpczEhno4PaCb/GnGdFfwYLt5VEVTAlx8tx1rIeKrsk8Je6lSE2bQ
KErelCAACjEfMQgnebe6DpsPg6bLlgznUa/PXGNTt8B3VwKDSCPvVIbdQXqC9pa9
91bpSmSvnG4K0HXzm3RPeNDcEbg6iAytuhCqqZ7FQr69LjyWWE2RJ3YQbZYATYDd
voeY8do6ltofq22bh9VtiIgk4BwUtQAOLoOqSPohOJkS3UgBQL2HzUWrjsPvEkgI
oBbwlqdqi+Pp9YmR/M8kxjLWwqq/yjcHfF1QsZr3pH0J8F7mVKwOmTEynSuHTUeu
hzvMwJ5K7TK54zgYFLY2inye72S0awYB7tS3KRPuyNYFzycBMsJS57m85EyRp+KS
6FlShVCquYcYrPjpfDyUyFx/OVgpbMnSs5mLijDYRWsw3+snaw23QU3FhPoMel5H
Ex92dTEwBvWj2YPPn7E8w51lY3nc7bV76NQ5L+Evwo5p86PHCFNV7Rqnl0rSKmaO
c6L1t+X4c29ZVNopMJlxG6phH358RWK8aDYv07upuIwqyRQvOAuri3NJIY/e2C+L
dyHwnZgpwbPah0EXFlJOPHPcM2gKMYJv+xsDMtGeB3fm/eLynr4uz3o1Xei3YDl6
wvGiFlu24Pzk+9GwMoXX45CAs9Pl09iG8EpHCZZqye4ADIifwCihS0jO8eG/aoSF
nDgE4fQvPJqOr5sSVw8fBVFPAgUzxAETg/o9IWtsKhi4/dvrws4ydArqgZAHyAil
aLMQH/RQR2DZ/rZkHh/PxmRli3Okzn1+7b3WAJkQ/Ru0C0KRWy5hTudgIYAEy5OU
lnfWOsZ3uzRzrgYonkkRefjwtt3lApk8FNTaIov9HSqk6III0Sqgk7WHT3qXoSis
6FHy/uMPRQEZxkE83fxUwkf/MsT9t09c7yLpPsKmIl4cUXvlS2Esvf4EIUlTQAYV
wr2Jxsy6fAexvKnA5oGuXinCNiqYDw83yflCpADE9AEw5SGxyLbwU2QDtTnK1WBn
OEJofuEzD9CgdSa226uQw0imJ/PG9/T6eLChAqed9iNhDW2pv0Gw5NIpHXZMMlSw
G0+EhGz0o59/IjXrfxC5gZBYeuxaysZvuls3jgIa4w8wLMp1sr6nzszqRw8NTY7h
yZcliN62VEOyIqrlMMMB0oIHZ1O+Rb98HZ0v0M1dANBbZvCj4r7FSIlm9SBSpkeL
tu3gNGSjrXowliw3kOdZe7aD2NijaWZ2s2AuIkG4IqN4mcI/vjnRkUXv0TLFEOF/
RVp84MZvXNEGk5h1r+lnyxXikZSzta40QCioUwg6A0D7eRs1qWh0yW3aIG22bPMG
km1hWNTb0hk4ju8QWa0tMrcPONPMfVIq+gh/gw/qepnulcxxYeaWq5jG5OYTe3Wc
DDgiBrIq+ue0kOeZDKJpkn305rckr+QD6FZh8DHcH/WaX4Nw53oJMIqr2z5V73KZ
VcrhsfwUK/V+tUPjcKVDn7V/FAluC1zfC42SyLaKoh7CE6ecHp4Nnfj+t2uLrj9N
e+P4Qxw1YdMO/8M7iIRfKJqyD51tegGBa+bD2nxA3O9ycnjjfvwJZePP4P4ShLaX
oFF2dEbC2sPpeHrmvLI/UXiVtzC5sISCnYTNSgGh8sS25461nPkJEStJOEak8Mwy
CDNh1FVySERYtlpKC7vXEHHmHc8OfpWUBRjipYVmoRUn/6ZUX/ohKZL6UiFGsVoO
14eu4ZOuOJINBF5S+8FJcX+D8AS7CE061S8bFdB6PNf9qQBVKuHIjWkejvxl77Vc
vbEpfrOK6yIfKEwYhz03lVrYiMoO4w0umQHEtV7SRrOhazqLucsh3l8G8rIPnvcA
7sANS2XtLqTlX7mvzv1x7Vq9e8CZj+Hsn0VukDDnRas9PfrYtyUwYWPxxY1iUKl1
1ScBlSRUeZPRpdBJHesGou+qv43V36tOX2jq6KT4aCUrRNHaOn4/63dP/ITSpSkv
lwFnsBH+YlDStN/rd3omhKyTFrIEgMo2lE2Vb5+He5inryxGCPpirh9nliLHVUaK
xRj+eXtAu1KJuiyIOo3Kxwd47uzKcSTLxMuT0m00I2SM9X+uXsKVY+DbYR5bGNeO
Zw5ONylX0EPMCDAi4I2NTmcJdSEuM//pCPHExiZTkdQlxVCNuZVe8hXUe/FYJKh9
SSVKr2ph2mYC5UkkDBAuRtPbm/MBKk4CpUmg664At9q7xNw/qwa2FtGn5xmR0TG4
/HP/suYhlF/u9cb75ko9+QQ/fWIQvUgInmtHEwIPMk8PWhu17VEKTYEnxfe1yMhH
lFYKGT4BjGJ7SNnmWt2/AY66Hmg/TErycjaKJlhaFyM7tNzg6reAt0sBE4bRQ4fE
KEk6F/3aK6FIp4K8B2RiX5hiknGPIJVfeo62Hu8bI7JpzdFrv4bSRwTYFIxH/zEg
pQuY8BBxVFTk1qGBfuzAQ5S4PbzfWInHqs1T7yacsfcRP9rrijxSUCzh+I+dacEL
IUj4Pq2lB6I4e4Tne3jN3lFL1sjlLiCDzRCyad+WjnzSnHOJItJbHKNMgx8kmW5K
HuFdXQWSHf4MvjFM5ZeG1v2BMk76BR9MLh83voqegv5f1O9Tjt1FV06aFb9D6sgf
ddkBkjG7F09PuNSUkj1BRPdnoQAbXk9BS53EU3vlOab+pX6bSFJ4BjyaFq7iI1V4
cWLh5KIYL2f3m10kGFB2NsGcqpxAEcNlmIfliPCAzJ0fovhmbbzVxK7yWXZXgbCP
puOSQXmKMshITB6quA5MBbt7PYVX4Wur9+WmTNsxer1mUrj5DqbxFt1NwZnvWaeV
F9O3IUMX/rw9RCHN2Np0c24un5dx7glgGF0GovI9lf3jmIgdL7XnmP9lxRS2H/Uk
ToDMBd8zXygCbpyn/0xrSj2ondE9Y0Pxt9FRUIIHfR654sEIntUlCeocwFW+Mv7J
e0QFsHfKQdqeiSKNzRvsEUjEjf9y+7Dr2RxvSDUBIZCSPl3zC5IppZB313lyyP/5
bOz+6AKZ20FJ9+IdCU40mpcHqH6rAhec4ztdrwUZe5jcyDvdxW265hJ8c3YM1mJ0
1rYpW7wKGJoJelwCVDXNszc4gBizcAJ9WYVNVW95cZt+KhhP8ZNtlNjTb2MHE0bF
rdNnygLgSlULrnY6XT39HiBl76OrX58QDl6TL4DlKvckk/yteAm8S+0GhNw9UH9x
sHYvYsfSrZdB7yvlO1kwl5F5xelES9ZQzDM7AiZH0M3BuTFmT71qNhUSCBfge0zF
3yX/ILTaUsTfDwxGImZdKYzzhgCqSVfPi9AG606tSV+Sq/0zPGvwcP98clTf5E0g
61ASWG874YGENw8KUMStlWUzk6HLBMx9kQ9YGmC8X9k48FEf2zVYZ9hKUZuFvqLY
DIMT7RgD3RpLHY5NR4Fb7i8VZLyA95Z4KVGgYpQkxmSWApubgxHDSS0eEk4uE1+j
K/vOy/vwxA5GyhfNq6Y8XIewyR3s7O4XKz4+P9chPtK17lXPd0d1atHHhN5BzbLF
+PvAdEy1UJCXuQtCmEmqRN3PXZDF0VRXOFGPPrGEQXDbpsZrbECwUDnor46nbWCN
BrKdl1KfODo+rGB0e16A3wV4k8EYYX21thqPLqy52/iQEvnYpw1tyhtsF/s69YY4
y33uAAEEKfjD5P/7s9f0aSx1gg2kJkUf9UUjc1jYq8xbZytf+2AHaELg7jZdTjnI
puGSORoprbmeNZBPnOVUlRccyEHhcyjKc68A7uYFcXOwT6jkfXu8kw3KNjH2em2D
DPKLvfN1FBchOZ8zQQribDc6Rux1RAf3XwCpOEqtgXQ9TwIjC7PcsrIc3z/vnaMa
cT6PnShNpbvor2mOot7xJ4JcM0JqDyrI7qUsoytj6+deCEKlD4XbZOaH/tzU+hDQ
9+9DG5l+krg+p1KDOKfdY2qUBYpxpz6qw1HLyUAyNKb0g+by8PaPSXM5GWW1xOtT
lkLVA8ajA5hsOtNNe46YUmvi3emBcTvy3NazgIQxzOSwxuS5lc0JTGB2Gn4VHEgj
pUBSddnyRmPjFv9GRfvYfB/Fcf8ECetiW76JOD6BAGdgcE2p49SksGDoFSqW/vbt
cXfPkOc8ekQiq0p0Im0+1gQg6nnl1edHX0FuY0s/apWiDYu3EVw0JtJCqm1+bc7+
75K+me802b+HBqGRhj5rWdVrz31n7XUd4eyCmC5Ol0sT19H3V6FVL2VtShS1rymc
B00d5uqpRBoPU0Ae4yio7Glln4UqMh+KtxqjVnmznQjZX/h7FgtufOAK23P+inLk
yb2MPiknKwSX/J4u9A+LzyIF/+JBAs71jUejSINDsFFE0wO9rgwPO/hXlszSSEen
BxXSe6VuWtMt8yA9fbQkuUAQtcb3j+29ZWBUJzM1Teq+zH6sd+9buQMZ2hB92njC
zaayt2w1YyA7k5ZE7nuYCVT04bP+M/B9rxcMlfJmbljRUjL68935Qjd79PPcbIsH
8DzJ9GZDWORwd/pB04WNP9bnyqgJJ9z8NF75FB0xNdkCH7nHakcShmYKG1ZRSkIQ
m9Ne4OyczNg+ax5e0DYe+sSP8stxluN7C6UgB36sZzKEFd1nPEjwYWlzWt4Qtyua
0R6V0R8OKkE+oHeWyRUmv2XCc4otAtgv2ru+cURX/p3NCeCunDI/y+rVdfUzVT35
UX2eVGLrQjwpAfVIInXYmlm20nvno02oa4Do31jr8g9lPrR/61hOMtSxuQMHSSfG
wmr5x//L4CQv8JYiIM+LcR7nf7lecF5vh5hogTlZRuT2294RhzQE8bpM3VZsM3rh
Z0DfffhFiZ0gfR3A8YuZY5CMrPUdBAMq4eFK+zSKA2NW3/gSI2adCQac/vuk6954
0mXpW5PerGObU80w9Nu/61VTN+HExMwvUqUnYiT9OilQMLqEPkS1m/mI4GTF09AO
jyycS4Zz6swyPZlWWB1PaqP6e2pDAXIKa2ez0kGGZUnxKZnviijU8lsq+CcVcgB/
RqGWsSOChZAXwlwCxvdODljOp9xW0txf3ToI8ZzI5JoqT7jWcu3R+w56lXQTI3Ln
x2ruHALeIsKzS7ePU0RgieRYBNRfFSGaiDVYdCO1ZcaT6KqdLf4PSj4VVB/yYzRb
exnvEI6srIUXIGoqzb/uCbYQpYQ0HdBPJgVgmnv4uZJJu8zNPWdc0HsAmVCWOuFl
Zh0cYjHfTa2b/AVIO4fxOFyI/mxbxD+MxzSfA2mwXTtsMWFx6iHlltq8Err+FZQY
hDFRQC5QSjol9DucxHEuzk2cUnZHUUCzEsGrgIj5oIuLyBGEB8E+7D7sMj7aIkx7
iTmGw3lq6v6nimdD1vtqxCi7OL+e9t+fmsa8sjEMxKg6GxRb292S5o5kZPXLU9QW
/cl4LALEp826+J9jqsV1UFh4JUJJqRJbTGZOdjqTCgMI3loOyzFFHKkPcU31/Xnn
zZFSjpqQu0blBLt2WLbKqdpDej08blazfS2CW0mcrw5QNW3Ro3AFp+BOTTVnvoAb
HahRif6KpmJqP/gGjOZfD3xlI9lYMgFH6HFmXQhVIHEicJcKO3wzWoGuBgw6zGYo
4N4XvFKyVKxNTExOAy6f9/la87sMopKyYlIGxXM2r4UHtd62BwipAJDBpcC+R/DN
lT+HdC4CNQ2+z5LZoFSCbJxqBX8iyq/3Yb9VXeoDk5o9sMQkKqE1IJPKrhzHdZJK
U14tsPdXVuYi9ZzQ63VriyWuDxsYA5LKI74aQq6ePpnVwEiEBLycsZLgnYByz40h
DXrgwLoxs51CznKGXz1TSMTVEFgCjS5Rp8CGM5YBvLzFo1sthr/Jjl547m92imKW
rfNawELatj95CTU7FdCZM8jBiAdUyFV17NWKrjlIJaiKhWrr2IGzCKgdJ1nOFiOo
jeASz+1Lw9LlvB2po6XmDn2+sUswghBg2EVMxo5ycikqSx7eQuv+CuHssyeWcACn
bPbKzb0CtMmJnROH+OS7ugkT1fHXW9//rweuUU8DFPRCzLgncAQuj3YOvynSJDOS
APlqxKH6Kx98KLNZIHZgA9mwVdy2KtMC4/iZouOsfMyaHOGZ//gqUE4qVZdw2JAC
DfKN7dww8RIXoqnZfxlH7lo+2ySSu+8OpLWKS2nlRQdacAiolgG0zZ+rhXKdacQ0
QKv1vT+mc2n01m+Wn664AtQ7E97bWbn9gNBmAXg/cVM+0CkImL3duj85nN4afHZd
5NjaKFxBUycKXK3CzVFAe23B7/VA1gy37pNAfSt9tV+k60FDRihTEpE7qEgf8AhG
y/5HgTTQuZzyDhrStdHVV8LtRU0sppcuewccJv5fPB7M7kOSoxx3yUbzAmN4uKCO
vFsmZngAOgA8tW1rB2lxCI8rpbH4GnCwTdm8FtnfRaGdoDUdHJNzErIJxlZYfxln
YpDYlao1yFc2jVbS2nazMkqwFan61dkqQole7vhYOFlsTBHhfX8hbo1ui1pspC1m
OajD1nqlazkI2DdxQeHEEcqWPdsjaspQ1FdFQPcCzNTeBbP8nhpvb9887ME5Xk9Z
vC5cn+KnT0tSDAucCFLwId4qY6UiHZrlM9SvyIDr1tQArz8hEYoOyNM62KIbnmib
D3c1HJiXAwzX2HKX9pmP+fYFb8Du0nIS/LxnhVglRbTKc+VoftshZEpN8RkoxevP
DxrnxO/WFVThJdR2t2/nRymTB9Vu7SCYwKiy/mjij/a8d9eoffjAIeuQrq0a0Ul/
JsONss2c3dof68JJdaiU0S8Mrk7oFoX75VN4BFAQcCgqRmR7reJSyjqf7gkhQDEN
RfM8S3hyaf7OXb/9OreWleMWxMzRWbxhtmyJ6bMvQTvgPn3nKS4pLnenGo4AjaBV
ia4JpP5DtnWATzBL+lEAgLDB5SnzrTejLT5bhcJFjPe3Kn+st1r2Ga1NmIJ2QZ/j
FIjk5u2cZU76lJWDJXTXRbu3yDK8cf3R3F7JbG9hwrATSf9aquWto9rFY0dMZYXh
L26b9rw4bD6vDdSBMPmGu3umeYu9zlpDGueCMYFGfjRxrlujypBzuPP2FJK27X9i
x5oWppI2EUd2/IbjH+OOMMSXFoxGABlMOXA6/v3dZfD2XXpN69/tREK2Vf+ZZ40d
jSpUohEeKyURrzIQdYWE0BFMvofbPO1bocNPQq+kiqfHtIsaWFdKGG0QRHYHdaaI
kwdheCBrm0MU69JDCa1xcMLa7aNhiekSonleHHFK10fSRQm/T/u19hZLD7ijU/0e
C2kshAESD7L1A7HPYC792sOL8Q7/rw33Y03Ed9PYfxJYOhLj0kBldavUNnsOoVG+
8RXuR86NDG7QyJXkDs/zPMdL9l8HrZmZ0oAL5rJAcSpSODzAeU3hhEcPYmXe2nfu
fFVP+aQxlYZhALBn2MPW+aLOfspmy5C3THbndsdA4Ka2YZNgAxkSYEyOFoZC5qb9
L/QAl3bqSoe5kthm9rdGJ4crA/vO0e6uI6mSVTEs6Tvm904sbSPbH0Te9V6mrA3t
jJaAfvobTsnGzLlsA+NukeniHBpFHZhSe7XmNRlR3mgYUtByl6ULJ4bny+iIxt85
lp9juLLEReQgUW5PqqySjRnfo0h5rlqfbpIqSti+dXGCV0GyKN4vkfCuNJ4xRUG7
/L/oKEKCoq3UBfPher2yXNp72EfH46LiU9X/x+JSYhag85mTJ1/YjqejbiMaBws2
8MjrQAOaRHQYwyM/LOtaXCFTJR5kaL09AiaA5Werq+OWYadHatXkxY14IrGiheNd
Cj+TJPhB7oM/2H7GjSdFxMyYmVKsobLLO+6l6C1OVwDjQBgohW3Q3Sm8Dzk7yGlj
r5hEvrEQP0/OanaxZUdkfGc+f/cAOPNM4V4DAJOGwzOL/U/t4K6Nnq967TGVyr5e
X+X0jszLBkvA6Q8BAEreTXmJPz0d9UcE7LNyU99fXjmgfKea46HltplwcNsX6ijE
nLXWgKJpQK0lQ2rdPwVct9i+pMxob29jO1SlqZPc92wKCIbbFsCaFIA9ISv4HGKR
7pIgGIJerAEyJlWIOaLjfQ8j+rsOK1kY7hlUwV8Fhoa2wfVAyG7VKxgXHdMOYGAy
LLKhL1PHEa/yQcytMjTIi2d+VzEy4meG3Cge9EF2Jl+i1mPfejzjtWvznlEsD4vi
vT47LTyLBP2AD8MNbtarLOWE+/06kbTb0Qbhgq1lDXWE1ykPamG/WzF6Sl5DAX9v
H4/6iBecdugiDQkNUX/7TjxzTaHpqOQBz6ezly665aj5niHGj0k2PhJvUbN7YBhC
r1mSrt/oEDFLZOPBP+ViZNJ6n9V5qqxvrHqClx4A5TUH1VPlElnzzdCuI/fSTy+R
swqvDVQe6XRLTvUCJ5AjUL2rR//rRqGCGjFNqri6EKo3/CSdlD1jaZNqGJamWPXP
f3fyMxh2sexaNBdySnqOzzlv7ijWZ4Mc4faRBrYRklSljBN6HETqtTibvYxKa8RM
eHeWuEdjAYxk347UFNenDehQnM31Lbp4AWi77tzKGawGlslWmbgCJte8WYkN4x+E
cVt1Xj4o4PZLGhH+MBfC9Tah/T44kePMltkpIzNYMmyvKczY5Blf7CPpge1tyK+i
/hcTYXcwBNhJQLiGW6kMI4GeEq3EUdcysPv04poeRqClVTfFe6hKZGrc+T/WkGxI
EEg7bRi1aZlfehgz+CzbIwRpwlAeW5j3nPmVc5ZsVNgPJ0xXRHThnwqr41nFb52I
3e6/m/cWDus4Ht+Lulcga+cWwl4n8QympLbpKFMzyEizsudGvyfaffCDpVoxPU4l
XPPNiDgN71urvybU5cYuAbsvZQ5YP4oihWpN5YpVvAUcxE0gtUo/qsysmtWK8JWs
GUccquu7bWw+zTSlrMP0afXQ2ApQWLQj2rl6UcG7aP3MvJF1458fnu7ktDyspuJK
LOq825VLP0DU/cl6CESLaRy7tyyN8+QO0PsSEESGyd755sD4FJSLl/FlkELcvVD4
hDBnQi8Rtq5asLp3+QyqWHaqSkjNsVi43PG8473c4jR+A/lKNKVNktHQx+q+QJyE
aeFtRmylJExwyG/706jYxh4+aXzUCYABPQZNNQwF+uAl/RaaQab8d0Clj028lFSp
M/5/Meuun1ooDXJfpPUS61XqVjElB/RwC07MIqRjorwkL8lycfy9MAwjiF+X9Kqm
JW7cKG4eZCsmQam7clEmp8ndXHs/Zmg5/qfdfj9w5qbWbWLPKKrYH86ijTV/crP7
l5AA+/kFAY8JWHCbmKxOzmTno/yN0xRGo1ElKuiuGtbsbrbUvXyTw5Z6gHqugCv8
r46PWCgAttBdRex0kBbJIBCKmpHE7Bj5nGM7pYrcxzIV5BrLtYkQin3bx3m64Qj/
jRKpEcYVYGguNuUzKwpzJBwDZ9iwNBM//ksUGK1Ez/Fgax/FTBI7OQCTSFI+/rSh
Z3yMnxE0A4IeeokfG1Jns3m/Bbovm88WH9af/xFpaJuo7hTgKtTD9xaTYR1FPmXS
2z7dY4q2cvGgvI77vjzq6cDVUsxYf3E1+vJ0NK6hX4p4NYTHa0c0463kTtO1wI0e
pEGfmM4OhFgFPS0+KCUS7yckPj/+gmd6aQ+1Dn+Wei8gsISjlOmebsefGmKQKjYQ
lx9cfewIu1Pk1nd7nbCKTYAor2iiH1+CctQx65wg2KhDblyOQbSGuL/VxLfdopID
VuoPI/hN5Cbb78pc07l31l6UCPUQ07br3DUnCCx3OnAmsEUctbE9yzyrx81lURZL
JzJpBTVL/ZoSLD+GK8oYmEg+yhQhAdRfbkQhODFYfATBQ0kzaMTwOPEdiqjNBbr7
DekTSPkeK2SaDYN81tFT1DBF5C8u38nAa+IqHmr1CRJGb37FvDyqjj3yvz8Prn9a
gb301DryDnj3J9sdelzNU3rcwu5LY2JJLGr8vF91P5WenHiQ4rgNrw9IvFDFtLJE
Rk5XAV52kkHuQTUoY6ua6y6hyZwRVjR5QxodG6kJCMHvhThrqbz1LWnSBqTCblVN
BEwBK+LWiLDFoEvDEMKrW2iQeHIhH8zZmLPShoQcQroDRteZlxV9BBx7cZMmne3x
LNZfVfOg5RGSqYzZvex6Y15AeHbjhrr6/I+4aUVyL96PdRHhdAVJ3+vjdWOlR7HK
4OKNbNMiBBj9C8cxRoetrA77brbZc2dw6B6MNrGScssityFsYJ0fjYRAbLF9iB0l
E5heH4lK1nWux9BiT8rrH9oBlOK2Irr8tuw8pW/kdx3wFcZGDxFJklkDbiDk0BgN
KWiMs+ry1ToyTSWw9DaE8+OG+6eUVPczjrVXrPQmRJAhrqshugcAlihaD2V33MAF
kyaUNDNJx53J9KH2l1IIRekgjCG1veQ7xb+npVjSTzvxfJ0rxjE2OQ6aBKkrbiR7
rXLO/XvACUA2VG3rwDtGTpCsvl0y/VjEjH8U9cz4xD2ncnVFN7DNQ8qUB/8f/NHd
uc8f+SWSYUFuRRUUCFlMOJ3wzoZMz2AnBr58Dc6NiDn/YLaYCl4xSIFix9Y/lkbt
03v310MgV+x3mOthaWGqwCi3IUeo7CJRxexmRpJhnqJwk/989dmFArhMf7wLP7oW
TGlJIeyTgkmF4OvYkF/tEBxMnfL6VLCpPTMRwaMHOfhCNprJ20u7smSjb0n4D7gm
sAlrhZQJYHbci+xKXrRiCPvGpRpxpR0+/DK0Fif58rXPHOZWf+Sses6sC9RcB2GT
anB0y/a9vI3/wOSq5WrAAaNU9hf8dJ8zb7sgC4O5J3OVbFMlQLuXaaoiTEAgPNnD
JrqePJGQW5DwZs6V459YVRCUPRw4DsXu+OGHVNU47Go0GiNBI74KtcR1oAvAXj0t
cTSADr5D97WbpHFdI4kfHvQIOKCxGciCmLZEqkmdVQkKaQYV0+tOlh7Y2YY918J5
l+/Uyl1PP2/SVEf8Rtnz0kPnjRvrddEWFzN9DmrCL40+ujddRyBqbEe6N9xgCpx7
K3FjnJNvUP3u2W5aFqf7+beOAhHpq5Z1hChGErJR7ReDDn4bIaIxrEN3alYyj1mB
WFL8+/lAN5arDKulMF2ehTSWDpwN8zrJXcMK2ScXfIhLBx0W+qUMRGgX0qc47b3F
sdAIHUduULkIy7RyjivvwA/hAQVCXttqYYJrFEfbFmRTmNexRTT8kjTE1z9n7wog
EaxPwNvq9gQpfUe0HRSjWdjs1Jn6IKT692gDiMOibEmVolXjyQ2Oed5oq9A5I67a
IgjLjKS6Odov8mAaUeo6SUABJlsg36A74kMU9ZnjoOsyuXty17ZaHwxXvHMRCI5d
ZD0Y/zNSNpy9opC5DVXGT/dz42q+kPk4PHJW2Oiwr1o8Jg3TrAEkLAgZYcMhapKS
jyGxFQlJbSDujDaXqY4v5Wfy9U/sdVSa1g3c6cjv/yrTIVTUt8n5s3E0X6E/PD7h
ywLCGUS4HxWCVAtp0wmi0g8fyik0xRgotNO2VriCbSSFd1ZqaBSmDp36jrBoiBfV
2xZMe9MkwRrTx4ZyWm8KPwn6IpP1R/ReToMA7i++T3UQsoNnETvR0jpIlH/OvBrn
UFs0j3CpYW66Hl8qwD5Elikimm/ToDqyo+VzZCIfBU1E4g5n4WYp4Wqxhd3vWtvE
trTHAuP/+Itsy24IVlca4qpgnhm/TiW2ApA5N+V3W5iVyKN0SqKTKqkauqBh7byZ
6zyAT0+U+yP1EqpCYb8nSAk5xhnfD8dOuNbCtnnYV6gPsOrkz2Mpe56ntJhL8bPF
kgETxkWM2rRP0UBQatEDAvRWxU78WOCFbWkbnU45Q7Y4QJUFLbgOQmEOPp+Vuioh
BcQLVMwiwRK1bByh+ZG1w5R/gRYzhuhZhfELhds5KgKjraPPbHjtIKEAndWOBweh
rjNMb9hiBXxfjTzNXXLaStn0+dHRdwUF866aqBzVe+moIizKvgHBxV0AsKi1CQ41
TMDsAYlFilH38DxaUL3fhxrdpkrMLzwQvZN/OSvodjjIYpP9WvPkM+eGrdxlxEK/
lQSUqo5uWKK9O57FlEarVAgvP5GG3QBIPBPK0CSjwz+K4eHSNjY3x07F4FQRbeSq
+xJqI71jUaU08G0u82an7TpWnsHJM+Mv03WqcUlFtxFvTVP4WFIZEP0fwmZ1SnVn
R6wpukKX9iGj352CDfoZKh/pGSHzRZ75cM+iwfLHpaqiwH2Ftm+Sge1I2i/GYLbQ
Ot8ZLt5GEL+v0i8+h9WuoN45nc5S5Ko5tOupcayRoql4lgKXkwo2yf/HR4qmlsm6
WV2fIh71Ms85BWs3a3hgml1UtrGFtI4jNz9Iem+oEx02rzhlauvAF39EoZZ/1Be+
c1KTxSw8x/nSh131lA0NdqRbtYPIrBPEG710LBCYodgJMKIlHprRJNd7yjiU7DpP
nQriEI7HirlrZRCW8TCpsUTob06AQZZZ6t0xKx8XoIznI+pi9Gpresz4U6dACXX1
Q/ZOXS2ctWzML3Q4ZRccu+M9+fbyrIBOkTWXEDKnPnub7qvcXIEqvfiEqOC/FFQk
NgChZJ77269+Zkkuytx+xDpP2vxYjusZcNA/x5m/vAWyIBBZH0L5BHl4/UDACg9Y
C8JYGWOqxeMtZPDAfNunBi+RjSprFYE5ktWevJP8FJTB613alXRILyHEOUxRPOdh
XKRU05v0EuL1D0ykjjm2WjGDoxo57uLwRNZuY45b9QbaG6ztnQnfbxNkVyWE7BQh
z6XzTE1rTbSfMidcsWYgoajj5WbE9jsuhJfn6atQfTrpQPUXgILisFJRZk0n3wnE
6T6jAKc5qxsS85eC4n12txi8LnAVpdokm+HU/Vuak4t40aLAK+5YCAMcv1PYZNTW
e47UgMqszSV1fcXkRJEurU9dV6ZWp+wO/BBa8gDSDhTwGGxsIoCKK38Lv2wFnxI0
je/sGE7eV8VWIdVKGTYCmzKb16JSwdvcqTAUXyIk+04+c0AwfL9VZ+DxU3ddGtwk
fjAZdjPlAHtoKf9hC569uzUsxl2940CU8jx8M+CY+OtjG7Cuk/sU1hkPgSivUSCK
n4S7msKd05LYNDWiKvGA1Koc4RBrMXc6ZGvGx4jX4Ts9HYY0nJ5ASvAy9frIDsJz
mYP7PXrQ92nWuxuq1RaDb2P3HsQNSV+0uRx+3r79Spleu6cW6WIk0DshTyxrhsMg
DWiNjQ/yNLivsrwNtUt+8FI8BtSdHNq6lDNNiUutSHbLXEB1HhzjVBpIEcNzirPg
x6o0JTsQzmrg7XrgElX9+SQMVncYZQSHCeq5wdeETnDfIypLAV+SAV+Czp8FFw8C
a+DWn3HwvjF416xH8MSm6beS3YSVyXJA6TAVq4ZHfAiyZxv43o1eSFj1LMCGimjN
NruV8E4OhWWb/R8Zc3jbBkxS3AT6nM3RjEnGxNL0sM58zGF9wIWGuSMEEU+zn0+2
XFn1JNWlUwuS+BtKXze1sgZEBduWKSrr3bxg3R4rptgg2rLczK1pKUmiM2c4ZEsY
H478+JhUoPvS4k7I3ewj6A9WEw7vsEw3GErykwAeoLWpL1j0oB6CqhDtSlqokXbF
4bU7AzgcKJXMJwsTqzSKgjvPUvqiPATqTgpY3voPb4/acmPXX35CG8ggMhSzDUOV
ALRP0lnWf4Ic+/RclTebESm48drv11nP0Oa6TerijZF5KBLTgVo+Tgsx22tg6fst
UZ5Sap7r0ZpWAaIcMhQOmJHxolHfrrbRVBcAjnefBQ2l5llUxT73ILCnLeDQ1r26
LToeLM2LDYZ5eCLUw8p/UvA7lq6Qwaq+GWz+vld9e7iQhvpqkvDQM8f1yuQ6RwA0
ypwMr3tv6rpGASm/mhEFRBwTL7+MZDK7tZlCeoGcqOhqspVltSTbUbpUH0/dyzKZ
GnBSecZtOnFozkFXuKeBHgu70dH3UetXJ6BboRwOJhM5Twq6wRbvVy3HIsiDGWz7
ZycNN55DmOuLrmZfTz0aS7jIQzCLYyKHnEbmxcVAiXhfUkIaO3r/WAQAGJORDPFL
IeohBoIOMTxDdSKEhc7XT0ztUP3AF9HRxnH4D8cCSzl4BXen8Jl+BXmHwcB+tL5J
K5UaD5JlDdPCx0XEZDoo0Stid9OwTFdjNNTXyVR+552L4K2WGwkuQx1RjiLyoNOF
AzDTj6yV1Iky15vcr6iiETBoa7hJPaCMQkL3/o/lss8wmLucKTZ/iKra0/AA4hTe
5SLwxBnOjX5ptduxixWeKyDehki2T5gQym89nE4f2y28O8kVmwMmko3ZFpjRWXhz
Y7IGyPOfHroRk+8VudA4TrLnj9QarS18J8tHav+fxpLqzGpyLF7sqt+p0UYSjUj3
hjM0E79bvMgaXjwFAduIWQY4bl0pspGVH22cQz9aYAG+pcnMrE3DpDCMV6RjLo2T
6UDWQEojelTtEZVtCnRmC7xNlcFPkx37uRMepc48KMdEkyWnap8Y2sd9lDIN52nc
GQ/43dDoMkw2sIHiMJ3IjtuCmzhajDhc8IxX3awUsotDU2n2owZRL0vLpjTEOja1
TpD1A/KT3FGiJ9aonRoCgSx9tusFJrN0d2B/aGFY24dW0lkNL+IcCNUPUaqxjcjr
9uHAfF+PE89c2QN9yBu+mzNLk8nLAcEV6suYx+66ggvK1nLkb3jvCVzOJErDnfy0
rCa7ftvRmtp/jRm8wLemhbWxBdSEpud2f8A5qCPji9wJNicstKQRTVUXlWlO/lsd
YavDiA+mYgdaYdIRHTmmrUebfNwafQFuB9BHPKHH2ux1r35xWtmLg/8DgVLOpVk2
RHEfHkQtoB8vkzXjregop2w5/oPODtuol9bQQVBN1EfbcXvYM0kYisldB+NmwPxl
iCkYh/91jmDzTjoXkMh7LV09zsaEb5PVjq2eArWS2Xuy31RODF/tCPvtC3dTuvEN
ey01dH8ui+CezPO8CT4P0RBWVqlJI4wUto2B9RpfEbmquiQ4AAL1T0GhfgNID2n1
rcx3I0OP/78C0Oz2bF/CsEmtPOlBJqkD+h1B/RnMPWTTXxhQIKamUn+ws4aosbTp
xqfHRsFTLQCGtiJQP/pb2cNXpFVQaJoRB6ysQR1MIZDJZV9VeTIyhh06QM1uUjL5
9JfRLY7ywo3A+dRhDqMcGzGyH37J3UWBbI4YpP+OrElx11j5L9jt+Ctbjh3jgaXp
XajpVpXXWXY+W6ZIIT3l61y2STvE6J9PNilzUiU4e0h+cjGDGqsxxYJ3L4YMPC6b
MZyYNyqtUrZAWlqu6nVGIIwIhlZWjNoAfUSo895a1DDcAp6c1GhSt1vOXiO8LSZH
fCGauvuHAOiv3kcztISZXHjXGB3MG6hyi5xlqPhNvNYhzlwAFQ10YYikho8ja8Qz
cNy6aCqnUS+HAu7mc0prvhhQ33XARJyxzCqPhFAA1tVlDlsTP3aJDnkh3cRyS56/
SBHbrWp/9BzPiE5dnpqfth1b+1U1gi8V7Ajb6CJ9UbQrSUF/kfg+ZQbnvMQ4lIQR
+vrH58VgCP1lLNXpKBUqEypf/4jjrLdqdoSxZ+ftHb9z6yLHWxW19pz4+KtVQbQ6
9BX0vwIso71Op5WM52K2wt3nNZpLTjIGt146OhNj1joUQoPq0O93xJ7YnGYI0h3/
VQtk5+0ILLjw9r2uf1dHgySe1WTHgonw8XVbO2wna7+e58HaR/0Oug/+9AP+CtfE
5nZeM/J5m7PuJYzbhnMZu92/afOe8L5nZjnyGYP1N0p8Fcn/BpTK9KBpJSfaej7d
QBvFOUPXGaWaxCE4peweiZ+fj9EAnnDxXHa+vzsyTzHKI6igdss3WVtDxaVrXNng
HljyvyIQT94QJe+268JYa+yQIwwApnyCbwwVjEKKhTFNKANmW2ybBlhvwXQUYHvS
Wng74Ssk51yyrYL08Kq1NmXKfz+lGPkmE0tEw0iEd1fnxGi5OUJ5WTfRywKP7/Ja
ox1YK8RWIm3rcAyz2leGZlq47+Njc6Nl5ACwJe7iy/nk6vperJ8+3RFiHWv9bSuA
WcAAQACjF+oKD/vbiAHozH/utYbUfrMJ4g0ucdjjvIlmkllSmNJBcv7Tc3eQRTJ7
/4pYLPLK93g6bjpzinBnDvN8wSj18X5cpa8rR7fSqejazVuuGGtggyTPIwb6MqDK
knjAWKos43J/rjdUzCzLMjMn0Jckpe0WfQ/6uMsIAvWuIs63PRLFJ/FtfD8+nNGC
RNg43Efp/r0qTBsf5KwNegqoBP+fFfDNJE52Cz5gfFzNT+A6gg9Qw6j+mKQdBODG
vFwqrVmOrQrg8iTCxCEM2fjnFllQlwDatUAOiL23MxIUrjzmpGWWe6b2pyynwVpu
qqf39o9eAZApgC3NAGYWmwN/sTbCeQWBOVsCCD1c/brY2L4KwA0XJypRz0PCG9pb
NOnqm0EQssRWtxADDuD3sB6yU1cj1btLbQy10Q7EaNMLx7dmw+O7w7+zrcC7KZ1D
kOV5bVi2ex70t65M1IlNyyKiPclNaUawdU9b1T/U6w3+DC34/ByKtjQGha/FDQHL
X2ECgqrQaevtSS5ni6huJ6wWT7xmmBZXEwey7Zf0vTqGVETtwMvQomZ02wK+RdDK
avweRCmUcceSJM1fit7kkKNWdd3WYBIhjAAgxhduJho5leU1knW5MourG6Ph/0HL
0PUCsEQSWPxScyPFsykzj/UcUQnqzvxBSYqYb81xyJQpHhsJUCKj6CXM/8cA8gqV
xyuG1xGWTJCsxMima8D7FrSWDIolIRCBRuy7QAlwsS6DkdabKtsXKM2RDU/7M2b4
7dLLGTdsgOnDl1Q3z+kVVzhloSHq7AOQpXJsjE1dlXGEiuEwYdUy/tZZ+MbXeT5o
eqvADT0L/6UVaHlHCGzYVUQKomGRF70d8kd8KWaQxK9tWIBYDW6eyQjSQ9cQZTDK
sQl7n7ktSyjPiDSXLIgZ38Qs5GK+ynePKHkGjifBOhr7Tx7s+LAoD8vgV79pDvt2
/+gsIJOxuKV7zLggA9w3tLYcKrBOSsrAQ21rw5AO6zVhvYqzx8HLrx0wgVD/bTe0
CoVSD14Y127uYkjpadGAlYD4SJ+rfaCrHGscqpr/SmQWI50UMCB+VwIng6/5ahXU
JUkgktnDDkGZFQa38+4zZtVoZW5XguTlqhjxf5Swc/iLyDtPNCBqArRNNgjXsouR
UZ3G6O6UPaqLEYObaZdm+fZYVcOLc8HvoEyIk3/6MXpNNpyMUCkfM1WaUErMG+vL
N63T4nhP2QOwlhje8JP1KKCiiWxrAgdfw9t7ywaUqW6QhYaRE7YU3NJbKBL7T434
+mxZ7j4d5q+67t/zx1u/DjQgApDnLbzSJc6uNEn4mbXnDscB1GBadKB1NzCse/b5
or7VebDrhtHbdL3dLqLwiUzLiZHt15nvQgH3h4XFQoUU9pn9nlKZCuspUuSSQSda
UKYvJBVdhZdwULOKw99frLA9tZR8wH9ZpKehcjP0cU1ub41qmv0LUKiWObMpJIEm
2kjm8R1i1Fop+ZORAloiIqM4U6yz7RCctknMzyY3Z5X2HHlM/0SivXWcPg9L/zd8
1VRQ2ijVNsewqTn6SvR/1aPMQG9UVIeKeVXRs4GKSkRRmiBNrA3Z1oXY3p9F5gIt
T0F91bSugAj9cGEUFEM0CUr+HrWKkrsWsyePZeH9HAKhEg1uevFU1aWWwcDGtLKf
dnHIGNOt3MNhsBt+NaFqqBl1v6fwFMC3AY7EUnyAISPrwC9+ir2C7ZsAMh5PqR0u
/CHEmaF71Zeg+xbttnRlriemZWlHlY2tH36JpucCe2Xy3QyedVoeThADqG4AvIcF
au5wmZNnW1vIvhxQe+18c5WqpMAsIQeg/vbAQEMvaERlI4JGGWJBZPF786cUct07
dgoF8zhnbtEQAfK3FOSExckC7r4WvtNkQ7IJWZcPdsCMn83alOOwjJgArqE4/boR
WH8/QQw9C+5RmM1HE/i+YcEe1DqMsf1eESoCg0nJyZpZw+pcbnCkgHHDhW6UCRhO
ict79eOIX9WtfhiqftDMb2OaSZpHuZo0ZWWHKdhpbwRTbnvTqOzM0XpR0TNebUGE
NTjLcNcMfFRucd2N0eEgldOarGgZgZg3NbKe0BRzEq9sZdq0fUFRkPNtzRT1q3kn
nyMltXFF6LR68zVliL4YQHo63VokgSkaOmTH2e58XcQIE/k4sTs7AegrqQd/K1pO
Rap1ZzgOkuEaPJiyP4rDD70NZwX0h9xv6ywzQmWYBFzx0Obz8wph8UegD8+a5f/q
XKld2nv7fUBxlTFL6i8i5jr7GIjQWA40OoC8ouTS/zJnHGWtAJUlmkH/2x0Nftly
KOiFfTviM9FBRvu2Kl1Ip7kimyF7I9BsfphfoO8Z1Vas1UVU5uY4gKFdY7mMocYz
UbSJWQwtuzhDy72nap1BAJlaVG5TKPlJPYMA8b56Py1dqyiK9u+PcoI2b/rgJesW
PIzmed7qgmBHacz5PyPkypII/xBY+h4E1Owx8rvDnnvEcDAX9uevsI7S1Fhgslo2
wpZx3P5DeZTMLsgRmO4sXFVQMOv27OeYkD+T/oAS9fZ/Q5oIFK7/T1rel4w9WLY5
RyB1rOucYwUMkwGQ6YBNlIV7aRLQNqKflNarUA/sX+0tQCOWrw2WRPG4ljpOWm6e
Z+9AXYyU54aYYr4O0z45+eKU6f2Wf8EohdaR3bJ3i3X9zWzddtC6o14E09iSA3qx
D5bV1sXe556EsYxN8DIbVQj9obAsZBvbtDGUWhvISseYh9TM1EnEVGl6No5hN+ti
lrbe2CC5lgjXpObECAK0e9yqK6fAM4Xqq+wvN4s3xGneRBSNjkfRCwQnH+vBrlAn
JDlIbSWJUuJYl46m4hgZEoOtZtHmNbwSlCF7GWCkhMl79x42LsTltskyJ/y0xX2O
aKx7wwjGwgW1d0PiJgnbODN6ghhVuVyWQ//5GKSwf8on9uRYA4kUz3dZiGMLYtV0
/mCEzDY//8GbpAFdnwIZLmSbsmeHGnzeFHJKdqxfR59pR4awv4KHJ4L7RfE16FfN
IgMbdEdSlru2nJmIuA6dFd+GG7Kgq24+ZXZwYa6dBVSkDl+QcuBwNKyWK9BRqc9Q
IOmv+kH+XEOSJb6hMY5/DkqkHJstby65XvfKHM613s5jbVCcRiEfCNGhU4v/gAKk
jblAZtbLF/fJ+aAtOht4xokY8/K/ttZHBinn1VtPUhav/6eNpHobH4ejGB2iQAI7
k57/1GSuuR/E+kVife21rVTD89l71Jp6pK7kmsdMcjytEkzD6DgctwwiaWDVwP7t
BFmPwrHEHLPFnCYS+ULeEJLRISIsGdA9uxLUAsYiIAij74g4blvDMtFIfTOVGijc
UMYs7qkFOmMn3PrPgF6CcIx0FdFcDMrNB4nYpDBRlfZn9kUTpO1wPVyKgfSKqIm5
nxTix1csxnb+MkbWuiP3IaomdOb9JneRFaNxpj9HaR9yT+RjFnxFwpClUFIZLTVh
55OZiNO/fjVXeCw3lJK37DyeSXXtWqlcriK0JDfuJl+nZdGbFTMEF9f3LfUdekzt
X1+OW7dQDH4qJ9NU2HEpc6uPeqT7o5ossi1Xpl+EZ4PXxmUmnugW0cuG6+nveBM0
I5wG/y09zBT5L70K7r2W+0f0WcI2a0n1jEWXp8OdGX3QdesMB6YvilX0bez5+gdC
o+yk0siR3olowhYyHSdo0gQnV8i6E6dYINXWwD83edVbJtwwy/e7QC01sJJvB2GR
fiuyQPaUjQrxygyDFQp6chzNFXdmPCtXqYIDwhSisWxxQ4xdAX6HTnJjbkIMAD3j
6/AhqzDPevwuHzFgcLEmZFZIbjUDWKt+VEoX84j6cTyfWlyMBUoHGfX4RlRC8Wn6
NfvaTKv7Xn8AnK/ju7+d08ku6MqL8450NCzZVeXtvi0NFZIad4R976oSKcGEVQmb
Db8mPSBNVu0Pf6Dxpvfwy9aC6AqHzVdoTqYhxlJ16cH7NXPGU2mRZ/pIVkhTf3Vs
07skz3WgXw0VBoZ+VbXcKdYlXLQJqtHCi6a6q9wIFsrU2EC5bkhrk8a+MptqM4UY
Xw+EtU9UnpN9/bHb3DHSL1peCrQi8iUYwrb6dZbfM55osCHSbv8Z/d/pC6So04rK
6bMzQiuLkiRnaEOVvN8adLSA4Yr38h058mbUbjEaDeci7G5dtEbkDclgrMNRwQ5t
SIvR3DVW3wmZnsXYKCRf+kMwj91n4otI77TJsdvCyUmm4iniJnbwb9Nh8cZKd3Fh
iwek57dna1/Pmtamtjwxluu7yqe5M5qYDMlzZEqk8gGRoWrB9So9+zTA915TGX7o
VSZZkLrm6f+0bYTf/qQU+PiMS362WZc9bP2kDWd5w/LM1Dpot0/uEmA8CsqmMYSY
cYhNsuyvAq1smi2ALgTsVX/IKktEZHCv35lQDoe9NbLQIejU1OwX4gjt7Zt5/Sqe
ognaklGIcM1ct8t20ixsMP1i5Vm0TvzGa3jmYazDj8EdVhEQMsJ0NYOPoyAerBsR
oBVGJiod4sTbjRGpXM1s1ts/y+pzxI4vFSvRAjhQLEoGFbS/xEPkJl7QqBmRSXRu
I+wVDtRoKikZOZE+YlvAJBA4cvckklhCKZs2NJVft7ORbPYPlzht16V0BN7ReWGK
wmm2Fuul6UJ1EMid4SKjA1+Bo00fL31MKqE9o4RtErhGyPX/LMsn3DLsL1yRLKy6
vL1wdQwwDzODDEGCeT9AcIvSuJhE1BEK+/h7Nfkgragop9CNDoAKbWFd5FYuWRBT
Z+UkBVCkY72BCU63V29N8mVXCBFYkJP0E9WVpDI1W9ZAgt2ef7xrRJRl4KXA7f3P
06vH754Fe6MnWJwAjCOeBU4GWo1oVpjOuTzfyYB/bBAHB+aVphc9rsn0da7uml4p
DgANFy/wvj+xxERpT4PCTe+PVpgRADdpe3Ob/Jv0HprANJVlLIdSXLR/LZEup3Mh
GOWGuHet3HZGbMe3X7Z5v7IK2i6oUesFyfsXFjF5+w0r9Oohwfk8VSiBQDbfY85N
Fv+ie1V6ytZ5Kfk1WfZkPB2k+dzMUVSPfFOL5lYhqme5RaSp3qBEggOM2B+pd7/g
aAD8J31kkQ8Ra17L4+NnfANgmwWIUpm8UTUdzJ3Xaov3QfFV0Y5SrKEUFU78ty1k
o2+36j7NBw8LCQdo9mKxtu1aDtdPR1TeBofucRKu2p9GNoVQBnnNz2fy0uQlr9Fx
mlHTeTs3cQIycSJ53hDPW/f4Bs5RlXV+ksoyLKBFO1yaHSNkI4GvMON9MsVeFfgB
JFsQnuNBPGB+Zjv6MY6RdGEptSXdzxla/CK8AlrReAFhxRu/qh4k75D30VFjoQPA
p4mv2lLbQdAjYkVrp5ZiIzHhrBJRl6rO9l+Or0ZpS9+KK7B4o5IpHF3uwAXIZoK/
iEO4XqYu/0YTnSV5gdJ9XU2Np7ouJ2Ig1k5xCOl7csNwl7smbJm+eTiOrgd18WOc
eGJX19CBzfYRqamMLVWTWXojhM4KuPCJIDuhAsSg2MnLrP8dilnY7NtXIP7lSfDW
z8SfUEfasYxRjMZUp+bQlBQibj5hSW5xD7Uam4WuJ9GJSe3l5bgjXvuufP69baGT
Nbg0sSDwfG8OXaRX0TBpETkKrz8PKJyH6WP1VbwUgH0xtMR8iAq3wlo215h/jgGB
rDLpo92tMd40neP0JC1AtJ1kdR1SwmOX8suWdBPOEK1lVRuNCEqZUEjAYmi4IBMF
ZpDQTSz62jHqhG2GCBOmDkTqyhx/iGG5KHsEuiP9425TKDmpLejwhFeCgdSMRkry
9B3BgAjClyXGJBR9IlCiOVHX9JE/N71dnIozCFtXr9fh/eHdBrFtnSJB0TyLMJlA
86ZjjxEgEPUYD2fVQz/JKLw3skIJIZjVAFFqEALQr+l35SAtQJYEMEaH6zl5+UyJ
MfcOWdXLrYAzds0R5whscHabVw2qMZWYVfv+LHJzXKDBahhSwNaVhG2jRtZlTha/
k1M1Ny+DWg/WRnTUx+YyjIpR8T+KUn0nAxQyf/zuxVk39KLNUXuwGmIPX/9mXsb6
wssyEZjvuCswVWxOpvROrsH+bvBOiuZ+Aqgk5Ztk0jLD1MoJYOky9Dmtc9kTk0/2
O6UMcS5Sf/OC82++VSpgUCjJWm25J3TCPIppo5Qz5rmqmxCdF9c8RVel+XtbNoyA
HsEXC2S3dwEVuoNYGsMkb+8kFavDVr7I7JCP8/k8EvlI37sHdQHUYeSQrj0LABLR
bpDHKW2Pa3JaqYBe4Ybi47FkVsut9/rTurF+QkivLrd0saNkKjhd4wOyXhu+JYUM
gdUemoLLirCrlaqoizAvIb5jDU6eBX2hgr6FvqaliAm/m/aHd/eoTScyE+L1cKH4
n0PMNTGPRwbDuEpcpmMHvgVMM4xy2VoSkYUx/Btsk5kgo1M41iv4CIx4IKg6ZXHr
LSewCQ0gl2MlkZuEKc6pmHWJADP8vkEFLmPpPM9YdomvUsKtCOvI4rqH05vxVe3O
we5iuj9q4+P8xacpUj6ZpMcwGdkNk60dp/Xpfw7cSNCNhD8n9O3uSl2ulH5JnoVB
gF7bdY0TAl7oWa1I0FGMhDcShgpz4iko/MB0UCH9AhojjfmWl1nYCjvD6/uSgIKT
C25KhTeoXxpR3e5w9eK81z+EwZZrnFHbz8L41jeeqyLthzRtQ1F3Gh4j4II68BW+
o78Z6H1VzzI/oISNMtJYBTzWvMLT0bhcCa6odGWJl2L1jZpV8GxojcvQPMiKavi+
GYva00TgWh4+NBHUTSPc548XLLKFEgGPalgM/WB5DN2IOXmOvetQvk+fQgMQDQXH
OcfpfVbXXgfBu89RUug6UykcndgZegVi/jPqT3kXwXipVFIoZYuZnv7A+4wR7QDL
MV2sWvOWKvAfHOfBgZf1WY3YC8QZi/Qr5ORvywFxR9BPQBxH18mzVIa18KmFGmzr
DzJnCp+7LxjNgQriRNfIhk8phU4Fymm4wdnlqworGoo4ZitEW5URybcbLNP1P4qd
RUL+SigIdoGp6WTVhGNbuBYs1GVMh+f1lyvyp799Hm8pQe8vtOGTBb09VtD6GD6u
F95vMojWU+I6sHEKEc4pKxKL1T6J79gbUj07Cp/lnlo0NhTrcpMJhVjFMnoIFCnd
w3vHi6wmUVowZVdjL9jOz5O7YaFqzGvRyzNP0EFxkERhQXUwNjX8tfAKPmrWTylS
ETUndvhruqrh4atNLDpEiZKDwtkkYaDCGHXu3UOjlLMJYFi9WNW683Pl1lyFGhBf
yl0YSJ5sgFKUAzHopLe046j/VP+jQnDgqEg6YiowcOhEU/xnmL1j9fDyTHN6uS71
MI+ta+J5d0ffiCB2V2cVGvGL5uS9Err3KVOL2cMkZe05h+qkdfIZPOsb+Jj6bTGj
CHr78mup85L6iQ9cDpfsV3VLPxIc6b6ztCLv5oV4sI8UrLuLdFZCNLgqGQUWE2Ft
EgM6mJLVbekrHCAzdHDgWxgIqqdT25Q+fXreYUg6GQsGi1REPL5FW0e9vlI3nw/H
ceFROHgo23jxLmJjqpnW+q7Cq87R1QX1grKHJU/QWM742XEOZYWE1XsF35xuYVw0
hRg1Y73WcXpVt3ndqLfYlfsqg/Xc6sVO6ObZWmyz5NBmf5h0ieVb1fn5AUjgYOPh
pNA56Bzpfu7yZpJXtNS0Eqop3YfsiAIvwjo4qkfHXFEjkoNoUBj04Zmc/gNrZl9a
Thkq3RLbwGLjMxMpt3njP1N6nPLRXB1JH53rmOXudzv1Cf+EukuZLNKDt9/1I2hn
76KO3nmV1iLV4ct+yW1JFHpMdYLOTRZubG4St9joyri8NvpYpgbSJDxy6MlKN7qQ
wKKlWAtLzUCTdn1M8FMA9B4K40HI8T+RYVbDGt8j06dOLjWhB0YMT5QPkMNLVimD
qlj8lM4H6PujFLu4AjkMvmRVG+fiyQpquV+byTQJ1UGREOZ6niAvJ1627WhxhJbC
WRoLkrTfzxkGJP8rNK0bJaWNM82CEAqcKSkHDAbpkcH8Khhme114GSrO7KaOrkkG
QMbnp2FgkXPRPRHCUNEIjnPV43r2sQSUKyaWjopPLIdPdQAlK2BtnxTIF9pH09eL
mnSA7JJ0HsLUGUNe651Uj19vuTnJuaqkyI4jvHhxUz9edWRXk4ZNMcMEqP3Rf3zb
Sd0Spb+FOMFGD34IJo+liFIWuMTzpWMkuKj6uGckR+KB1MtKrsGqSd6V+5TSivAc
TqnTFir17DV1d1949ja/xZ9lGdW50mxay4wJo7fUHzJ/5BAd22ZiluZAUTSgLFQB
CcxSYKb/A8yoNl2xH/I14GXjvEL9bp+wnpPCFAu9hGxlPRwQPI7Z2xVvsosYlAvs
pWLfRNiSE9y9qKMOxhwpDQVYvxDYzBpUmUD1tNjObtZqM+i2v04EEk+Vo3LQAyUE
9n9emyUbIe3hiu5+X4JPquVA7tF3Eia7Gt6JkFons+vhs5Q8/M7KzIw1yE21bsD+
IM5FOI7tsCSkgTP7YsTuG4m/YMHX9XBH7DiG/86lbzoxkTYeipk2AxpOk83wpwS6
+9i63ek1Akf20ifu1I81d3DgmOcenxBv7XlOWhb+ZXRIKmKDbmEbXxjW9iup5IWy
AO7gzJH1z4Vd8Qhk1t6kzZ+/Jdu42NVzs2dJF36CgtfKWIvfmvSd+JVWLlYnWe4A
YtJjX+FuM+Dds4N1y6i7mBm/w+eFpM6ca2jEq8hD4tii0Ew1EW+RbkxoBsC1xg9Y
n/iOIM53E9/6Mfd7VW5C0ZEs+dZhUcUj8yzMUXgsMPqBTOgTXJXPtc3FOizyeDHX
yXD+AKr9PBgu75ERupod616eQv2lJtnlYa2sUzZHs/+g1Y1RXHBLtrXeNLNQ7WVV
hG7jBFRsUQrQX210jeMwmTW+vfl9FkuMFnEgKST6Hn7dBrrmXHjLVheEr7S8jPm1
DWsOJE3u7DGWUJSdiPYt8oEArJzpbxV3xE8etGrrNEbSBKoRmlQj6ENzeaFQAOxl
6mE8sWNI+7iyTj3j6upyaWhh5lefjURP5iMZF5ZvSZO5NxmMe/nwI8F8sSeJLi8q
H5RamShOo+JMKbgx5joN3zpWtluBx6CZDbbor3aQ6C5VGsDfUAJdF0pTPumHuyqa
f89yH7tUecA7WB12iSlzK1HGiJASiMVpNmcBLQFfUdAMr4FVTKYCxIliEmuDY1s8
qvs45RIFz+W3nScu6n9t/GGBG1qGkmD2dPuXiXYY8pN44JuXv40xQ17Isw83wxYA
xFzfciTRKP7btEf+EyherNohqGsIgnPDGIKcf+V+qF7oOBeYPSJ2v+QyKS+HhdBM
IsdCWLFQzeubwqsNdrFa3kEzvmogIJj9AO+l+cNENxA/XWgOu8niGHQ6+Lft79r7
bi684aGrWWPiSpI5p+MgUOLXxtpa4Vo5NTcpI3EckfVJa7Xr5ZNk+cD26GBz1kNk
AQGyYXz+jPih3RvjNJeqM1bkV+iKKBc3+TMOLuJUmMo8BJmXlbrlwTUUFS1WUvSc
ryqSOvTAtcpfag4QsjP3Dt3rL/5u2oAqSb2poX8OXwCMC5bJcJKxJVyFEnv8zj/z
OeaA69PikfMuSevyzT5WLtXorpcQycNLjfyhhyoJ2CGyyUqXodIYhMZpym2t43iq
T6wmXqGn7IHk3P5oYIRfGkiu9emzjoak0xXsBwoCmrG++eQFg1rxWvODHXztRJPo
HBm2B2KyH4gYOANEncRlxERtaIlJE/xz1iZ42i0ULv6di7m1PJ/xHtIx9IPTmmDl
gKTuo/xxTB0JLZ9tfa5wOXHHKuj7WKkT50eDEW8ExBIFgdeMoSk9KgaEVvIljFDU
Sz+yjq7NJPMkPCmX/FwIKovxABi7KUe1RA/6vpxsCRCX8ypGvtjrzX/7cM00s+Zq
CwmFFDfYx/dsvsZdE4WPJANjALeZT0Ljnou6zm5N7IzuRsqd/qgc7aNwLBYEXStM
doaqMp7ZTagp2jXhWIfQuMNe4vdWcqgvlcdw8ntjVC0GlXPpdujlJe7MBCdxa/kG
d3qi3luzBJMqqC3ydWD9nBwqpBNG3eRGluMKWbdhQF24WT4QEdgQ7gs2iD6E+2oR
ZgGyXW0J5x1jjQe+ZCtfT/UxJ2C0u6/zGhqYfZP2EqA+M2KOgF8ieky5w9wriqu9
pQpeZaY3a84H6drwXDwCVgcGl1J1Xx7jpgh5iCbBwyOyyYC7u4jpWBWDXiAKktVk
l3AOelMZhFtUZorpzOo7e2xtKG+QOcTqoHnaf1MPQR/a9ePVAYFtHLPKS3GV4V/E
x1Am/W3qBW2BulQTZ1m+keoK4AxhgyxybJn89Ia+TP09gOUAV7WfsP4njEcxJNQO
9w9aAxTgvDHlQ6NetqCPtAwDz9pz6ncOOl7RbOg945NOT6Cq7sl1Bs0co8A4yXpw
ophTzXN+XNdubWKMtvWCX2wP2ADkvPBCR81E6qbmZu1pnabFLLtBYcypk7SAb83+
6Gksx4CwJWXbvusLAC93N+wDXCkdGAole7GwfJF5WAsVdq5vbq7NPBB7gnLD+U1/
SKAq2vpl+BeEEYZFH7tsCqNGjowNgw5nWOHKlvB0RkEpBg5GXwGDU9g2XgSxsT56
Y79C6KbLqDxVnvwLnm8w5ciGUeGAmHDJ7IFD6o49HCQ9bJj3OrGavOeIy/5r0mfF
GqU6B1hjLGx1FQAqKsYCTUvO2nnLlPhNCtITHNwW0Wj62vb9SCxfTnMWKdVNiEFK
rsmQRZ6CBCLsLysKLKoFBKUaSMPbbP4U5gAsaFG/pP6GtNKl876JBtiEooBvGLma
pEcU8+MjytNHMyUmvRRhxcerMWJfQUQ2iQS8vfov6qVNF3hTxU2y5QK6od8s9uR4
1b+Iho1QeDKm1w2JX9RXlfk6Tnr2SqpRgck4oSKt5t/19LvY8utPW83cOOlMAp/S
++rersstEpXCKnRPGN8oMkE6DKHLvBZikuJZZGY8QoXa+mwXfmxO9r572RIyDIRs
qQAN1EmdzLWOkbbaO9NXk7NiiZeHAjyeAJPji5J8xQFyT5Vy/UNXoncEIUkqsxcG
fFLb6DLQ11L2WAAdY8e80wD3vMouu+n0I9OdNDD0zrSwUYjO9JwwdhngDd4IS0Vs
vwiHIyw57UJI3tGOCPwBjbnx/SGLeZPTEXyJmlleyW4+DJPzblrqL5DxRvB+NoYq
W6zrP8ZN23cfsJNY60fn8aNPgJMSP0kqc07pMWK3zND/RNWCgZrwcAoxtGQETGIn
TByUk7MGQzTVPuLYuBsz4Gj8WL8ARqbW3j5U7aoXagyjYjGXyo0lZXZ0LMGm8pPq
cO8BQ0WYa6ieXF/797a/NCjUmBQR+qa+QbLyBwDBgw+A7QrPifXBxFgP3TgcFWdh
Rr712JoUpiolKEUl0hJaUBOhoExc9F4VLPSCd4hAtEx7UEkiziaMj9PJSbfgPC3w
YYx/U8Q2UAAnxTu2YgS7kgHj86kuBdNWKW8xot5VGv3jmZknXukvmOWfBfazOUEk
DEOpaijISpso8vztYysGoEaPdu17U8YrvWCUAIZHrNsmMvZy0855+aBMMf8cjIov
AiSdHVG1oaD0pIkOscU3xGi6HvSjtDUKfx9Tc6MRV3u61SiwKxezKYQAOH+M+eSq
jNmkis5LOWkdduDf9ui7E+OEZJmOPvM5h/jFeYbtEL3Cddfwg6VveU+s1teEhFZ6
WaWIas1hd0Mf6a9s6L+6G7YRJ2jaAF83fX4WncbEHp314D+A8kwd5F9faPBgs+DN
NpxxTzDySImFHyNVf/43iCPxJDiP+MOdWaMMDynRuUEOLRmyNQ88IQCWW0DBZ0q3
8ksNTey1kQt0WyiH1qoq4SjX3KOk6oPliCSTO/rJbXmBtuO7bNRyxOJLA8ZWtnIn
xLyB/qZjeARkY2qtOXMkgPIlvEoTzfm+OZWJkBpcsztqZblYQKsu4uijCz6YY1tF
WiICnF9uWIi6MX/r3yoyHfpDxwYlFFP7OrvL0nrd9AIQi0XqDs/5+nhSCldIlDYa
0nJwkPcF59y5vEUEr7HqRqP6m7m8cy39lefO4pZRtBODqUayNgehTIsn3frpnbCF
T+DHf6tMsGt/qa+Q9/ZK9xN1CBivBC3C8VOdXlzteuFrWPoYK3oWGRPJDcVMs7zr
UrBzCQFIZeh+UM85axcRNEJ+7bCWfOKLPlQQRaGqRc1COCPJ+2ktu+q9nqZ5odVw
48GhnuoY1yx7aJysCpVWtB8QJer7XFUye8zvfYtfeQ2sA2WVU+B+I4OGqxB+rBQS
B1fO4/mBvCkt4s9tHjdup3xs9aALXb9rW4DMaM9dtjh2AdBs7KIxtoxD66PVnRfd
eC5PicYjV9mEZbUTPy4BbXyZjUrUlWiWaz4oywdz0YWRXO94Nkq9inmVflH68XQm
5tV4vFzqyQ7KRWs++ll9ni0lB08yySzqTnllQl+3idZR5zU/IX22u3Uf2EF1oN/T
u/RDWyX6F3EIpiskwNKJat2jCuOhOcbhTgs8QrELnG/Zz0a57j8GmnxTsue9CKL4
113k8f+FFElvy9OhDEmOTa0kPNVEq+onWBN237F1s0xBi055C73+NtYrEz6rHh4T
T8Ko3JxjEEhq2fw1kqYdA7e6EgSGex87kevozgV0KzbfU8K9XM1+2lZjiyfJLjgH
SoMMcN7tGFyBJfbdcYKHdQA/tA/6uwQrmVS5zqizVbc8lLy0aUOfDiay05LUckbC
xMoQqSZ7piRctiLdquEg+BVvUY0gqOutJw56Rc4oMMAEOLKoXBl8pTw4aqIbhEQv
2F2QGe+AWNeBhSCHVa+iwTwOqvSAEQt8feegdkHD1TRBasea4JisMOkfqP1yV0X/
vLcSrLD2VhtVnZhlvf3vq3YwurXSGzdSiR9xX+veA5eJxbcnMHvjCwVd4XugCA0w
3gLl3WD4U0/trgCcOdL0EFbPhoGUGMR+mKj+tlWcL8tAlrV2OqIP6YEdTBp5cuVW
0Ps5hTmpqPJypD/ASB0GXIeNFGP4egVaxV/XGZso/pP/mi+d4PNecbRt1Tiph70g
B5icMmP8q7FMTQggVPgNKoLm2wNosV/AUSWNU7cg/Yy9vECx1HNUCTaSEmHnbkac
NcYWTeJKTSxV3xAis1iBAPeEiXu40Fh29z9uW3FgW2F6fcyficzCK4BijuHTjiqE
baFHxyVTiAVKcc6DjUCbfOuumYhG66FtB6wOT0cfPeeTo+g4RgBEzJ7jHtCXnrLD
jGfIHhgFiiMSBR4sEkRQMr3KFvh203Lq9gEmCUYH8zRAeO1hsbIWTaNdeNYYmMR3
Y0w3Qf+D1iMZvZhIKC+JxRuT4Rp0qBBj4h2fyVSSWOq3pOH0n9zxZt9Wbn6lnK2b
KzMgBuHIrXy/iHDt0jydk7ylz1YaX2tMlsqFVs8IPpFET48r7SVOJ8EEJOz+beLZ
gV/0kwupRiMJz6VvqsbzL6OOX3GbGPDnl7DixfdagCsNvkyl38+BDXBD1MvYbl4X
MnqSkJ3Zgi9TdgxBRDgRBVSJBiRN7ZCGDBxJfAo7Wqkb5Zx511KAb/x1P9pRFb58
GETuM12Aj9rvAl1vKRA6N/xZrzJX3nNSwIMA9EBkuyPq6v+UZAdLqZEpnUQsqLZQ
IC05jzcDQqFYscImpUjLxMIIy52G0b1RKmnB1H0sdUCo/tL7NklZtIQx0KOvU+M2
ntlLsRg0JnocwTmfco0rQ7UmkkqjkH/bIrWVkgcIvO6PwfUgbL3BZUqZJmvl0wyY
ddWmAyO1cOni70h1KhKJ3D+DsovTcRwFtcT+oOoDPtBsZsLfjiKE5FvCceP/InyX
lgy/sB71XXWAoh1ns0dXfKEIGKVhnbmguW7lULG6/nhdM4wCG9h445+UMC+nk0v6
Sk0xHJVM7h9pf/ETeGU1Njdm1rRFcPUmsEVg1sGqBRffwxkP4OmN5MxerqpmQerl
0WKdotlBVaDgbS51RTZPpdv+GaHRSj/YQBpuyJTSzIxAVI5Z59qoKlG8RpgSpKvd
I/j/b5jytUazq5+kd0p7vlR3drx9FYYA6wCHO8cd1MtBWqUVAaPCrmA4RSsF0Nd7
U1RS7N8K9I0iPhfQj7AM4/be83AquxzO7JtAkPtDvEO8xqxSbU17W7ZqrhwK9fFA
/s9xJUyPO3/BhwiRf0JR/dIGFHskXGsjwHkpiv+I3w4X0+d93hm53Z+M8yGBUrSa
HIbWwAKkpl/BnvTdRLStFxBFvHnYUUijGmKE1mw8iQuais6AiiEIK5RLuv7f1qzd
42srsii+QR/XCGydDeRgENHe5yKUZKctctgYyPpwcC+mEosNGm1KeCBGJigA2h47
poCmlGx781VgWcbr40sJwze+kMckSJWCTwMfDjscgCAk68ncBrKe6kQhjVXdH13E
cLoQesu8hfLpmOZx9+wSUNMjO+q2P0q2vh46D32s86Qd7I7r67sJis0M0DcEPoDt
yU4G7Wc5Cf0GRX75PTrb4Erie9/QDAOigmW98++iLyPkVAli2jnMjX0hmuPkXUDm
oilMM0Sl/g8N4DMHnkdHafwcQsjbtIQh8DZ/9/Rkm2QJyo1TdE2qO5jsn8sunOhs
SNFyPrz7N5CV+I1/Zf83raojvUjOvrLCNauj98nGLTcCWDp+MBY8TXvDlruwpT8p
N7Kcqra2UYjbiYP3GWBLoSka3wKlg10Esdh6ysD6sP9/UPW1hiKnI0d0KSu9PWcC
wepjlytXZYkt6l7yS9KJYoQp6xzQsMFuRnumwU2v3n5ySasY7ve17Z4jlpSiH+n8
/YOwz6YFuOWBGe6uoEGPg/tRB1ocaP6uVJmGh7sa+z/cnd16EyrMsivw8WD8pH/q
QsbH6ezEw0yQ99UqofXlVJOIKrLDZeIl99K3CHsNifg/5W9SBybRuo2ElmJq0H7s
PN7ODU/NF0nfSd1we6eQosmWZ/44i4RtdVDu6w6OHKC7SNs2zSnfZr7FPNzuAP4V
ok9W77wl1QTSdjrnInHYX71mxc7b5hZ/AE6vYk3Ra/N9Pi1iKUeUTG3IwYSJi+po
HME0plfmu8MxGdqeNhUfg/1jzoM3Hfv3bTFscnePVUkeLP2uR27Wti6LfaE6JAs6
9EvHkJ6ji1oo3BvECeLnL9TPfoVvQDfwjbfJUs+cwbSV6yWEwn/sHSJcVHjywl/1
TBKomBm3Md6N0/opZzRFuqbxGJUcRFr5GBEcwyxQyE1k0UtP105dHyCkeLA5k3uo
54Zqihn9Cue9cNKYZ0E9OIjluD5J5RBQnwTb8YYap3nd3Ff3wcZRLaXzz0kjQA2A
juK2A58ok0f/8pZgXPIeroFV6m7Dc2AGbJzhHoCIWPA74kb4bggVHlzAwgjXJnKL
P1dowMnTHG5CVgcuq/3Ifpqh8MmV9Ur0n6vVTtWdYhyLUqayy68ZPeZJZ6gi7dHS
qcZeu5DBxaHUGZrXvt7RwzJ89Hc8wYHKYHCns26KTUdq6+9EvzrdZF5lRtdQZ3ZY
q+Ph98o96wvEdOUhSWp+lqYixqXDcDSqUPkffGLS59IHO6MWEYUaMcoTin+n2vzo
qkqnMMknFXRtTxxGa/XSS+0hcgfAKu/5JZdTOHO/UHq2Fd90TYbI0+sZLSrt58Vu
QTqXwlt6ccyPndr4dtFDJKzo0nTw4d7kbo+tNQVYDD8SaEdssX+yvHu1qUDFUDBY
lGNgscktOuzgOseJT/Dj83FfPghwEdD7iDj2uEuR79P/JFa4vfc31s7oaLAH+TY+
2StcSzinBh/FW5HTlpdP3Jy4KlMA02woACSnLDlNve5TBXfoGqhOQBoKZ4G/tB2K
kowT6Otd2A6UaebJ/8dlCHajzkE/QeuXF+dTXMyd62hQT4Rc5IS38hBnqL2jx5ta
VQdFgij8No2hZlppVHXlq9OkttHYgiU2Jc0Fa6JuJ7hGzbcSgFn9KoBrZ6LQnlPE
ShsoV+yMJuoLRKcMCbDP6s9lLTgnHXXfVcBu6REEF3d/mCJhfMLGh8ADfbkOAr5s
SB7vcfRxvw0s+85wDY1mMQhUnH8rELsxVZFqYB7LnC2aW3TuIocv4a42c4/ehrbe
cu8290LhYRtm7LXXon++DymG30b8BRPRH9y20xOorIkLU0asyB4M/5k32j0mIhMg
TayE19Vp5+bO6udyz5W5+LRbXz+v07GVwXQ4FIM8YFPiWs47J5fle+0TurchmRWl
WU1C9MgW3cDW3YHH2MQ5ui6kyhnV9PH00Qf7putl3C/r9xAK/rMuiEWUSabEZuet
w0oEG1NSsPgQBYKKW/GaABza/gzl+/NYrIUvgZpE6SNy4KD1DqtXDZB0rxhnY/Yg
vGOCqRYn2peYz2OUMVNcQJ+Uv7Fd4G8Rsl1RmK79F8yWftp47iKeykn48MPSc9Ei
QWTvHI4NuC/oVSyipjGOC2dZbDlj4Eag7h5HfF8tzG20usN71hGHwCWHIfGyIN70
AUDF8g3Ok46+hwDtJr7/FYeQgrBTuE9gfBHd3q1bD6qqX7yHpXnw9XOmZYKynQ/v
QaPsaNJVwCWH6vZQ5DDJVa6yfcyi2OnfCfNXdSoQhwXq8uPMBoSZPSN00PVEng3q
7Hi58vuFNzsIGPnW5KtZ8hCBBIyO8Jw88XKAFgjrFpXiEl5YIZnXRKVkwNJFcav9
DQASh1qbCM4nD8e27F9N6R25AT8rTjrWv2msydJjsDKR3TlyTaeCicebP9n2dNSG
57VSzB3XhGYnLX6F5foJb/HEs8nVP3/loRWFJC88xRL07O5OOWdmWrgwfQVApLQx
MClLneGFMRVQqrYNoD5iXBywOOWIRs2FZSz+8fMqrn9s+fiJv8HNtPYz/zQqrZBK
5cRo7qKabssHgXXthubiFano73jRYV+1M5vSTw7chHNJsDiguBU2Qemkn0KfmnlV
0uImusHDTDOGz6ZdqbnCOGBrw0PtekXyeGDZS3cBahppznU+M6P619E+j8ZfMPUF
NHwBbxrmGfb4TlEWyePqjVAPifCbXrjmADVm5rYI4/3a2vKW7AzMmK+LQER0Gp0L
oCReK/s9/5b7Qrr7MlZLHZRuDrpmalbmHiC6gjjxWFm69bwfoAhdbsBG84nwnk6R
Y8KVsaFSnr/RjgipJ9zTo5rurcGNRpXfeTwX/VCFCC43XZ+ykQlO0KpaPqd6lbnO
Q9TTqwhGjX+/fAnJs8TPhcIsvZoVmz9+iS6eesJElzH0BqyOyxmbex0Knvoeojrr
7io5pKRmnA/9Q2NGHTGZQ9unZPH23xC5Xg/GX4K10xHkY/wbpNBTsf7DSG9hAgBv
r5nEC47bqw6AOl4F6sBTthSC89ggiXOnJxeO1xYXNdlLeO5H7bBRbQ7jFwdvGhad
vZ4b8MjfZ4CLUmMqTxfJFt4PHeRbxXrBfwdBdgnEFZudj6Pfd0ePF0Rr+TsQoPyQ
+DjBrpOSu2PNI7Rk7RYHjGHG5+TmDdbhvp7Mm2zKr2kfCOk72v9aqbRKrut+lhYz
YrSkDHIRJLvL/Gf5cOZPMVaUHhiGZ7oGNep4OGJ2YHa0jNi84ctU3nSFLaY0jy9F
EARZeRqHi7f2qEj46XY2avIpUZinadsM/ubv9asm3XR07yU4D3ZerDoespU+P478
dEz3xKjFM8chzzuaSzYvthywbXWmT6ImCXFTXZ3AVUFNDLy23+2ZGgNbDUiuUrmG
XBZpchyUGM6RhJthHctnqwFMt2tuvxxcG24Cqf1AfRaouI/O45sPNGChTz1Zx0e6
zjzhTFx5HFpVvgknOhvnoDB6Oyoo43p3dsESSOnxiEmK13ODuJsOeB6WxILIO3z9
ubZWwt+bTmYnP6W9fAmxJPyZJXliphdp/s9lrH4HtMz1sFhmjudWxVi0HXAnBvr1
863FAKCbMNg+pMHUTj7G3G75JrVCImLeAXNFmbxcL9R0iNKiYdN46LPTiN8PlPFY
S9B9/2PAtSqOgHlv+bhHETAA7RWDGX/2/uJhUdWrA2PRkmuwWM+3Z0Zka1TclLRC
W/hTvF/ttp8EOwvcT8flLfacrEV+I8NmutaYldv1T0cPLgeKZ61OB/p/Pu+1Ej5O
u+iNiw+kd8Y0xHKiiFJWRTaDAZyZR1zfGtqUA3BPSJ+MxZChc027DOB7WGb3Kq/I
3vb4ept4t0rFQHriZPxvL31xt2EDWCiX/qNcQVOd3uawMeEVL6u5Y0g1Ku4GsPz4
lxOZZc/54SaAWxykEdjKKzdIQG9tF/ax4CXGuShWgmXwzDMArrGStt4/dqmGeImU
4vXvTXTfZuVRgfmH5o15fYqLBrgWrnAXjbH7Zc5KePMoLd64nPiwq7LrOXeOLHE5
w+eLMkwGPcgPLUwPVbOTgO3fs8VU+0dqLrTmVkB/EHFeHThEmgfLf4xcZs7/Deb4
bCimgVwU+UZE9n0GXtkhqmLneey7qkVk8OmfHDRB4ohZlvxb/ByPDNMHK8dYzJ1Q
b/RK+XVe32J2YdPLrbw/h/zSqVe3jja7YnbmSjMwQX9cdjQ//BEJg+KWOSPesy/Y
1uF13NCZrzGWmOT94Q2AqNi3bWV+inC/kMQ8vcepBttM4qrYFdJ9CbKEg97w1Eh8
CBH0h5sl5gZWNtJ3RVgeNo60AuHrm+Eh33iPh2hGtDuAXuMgiO9JFwcIy4o+xv+D
GvpKIJCP2RNhGVQPZUv6lZTN7TnqGm7jr1njFQQk7rDgbNhE3Hvt65Xgyp7ksKT7
KP+i91sSspBS64+aLsfRFCbEqIXfvkFL/ZzyyRa6W/Qt/kqYhiAjIyhxxMFhYjSK
jsJNeXRTO6J3JmgHsaqfYsNXpZR3lEqtsakY+o6Kh00kDCizl8pgLuI0WyNR2sfV
C+UfqTpmKJHnnBjCyqm5tHuL+mXYmECswLfbmAUOV6wq8GtLKZynovhrGTd/wzjx
25Y10AxXdZgOulFQ4rXlmIXwxLIMyduefUnfZB27t/uNlxAWr4j8o8bwyDtQ5s7D
OR9pvfsDDq+WaN/tykMaSYv+NwEXcAi2mhTVJQVBs7M/Sma/3ULLnyGc2VIf8Nk3
r2U+Ag/HYI6SDV0tZpq4JA+tqY/pBoS6oiwDk1RS7PyHau/TTU1LBZ97tU65Py2h
0YuNrvj4vtyNa4R1o/4g3GnF8l5iN52YcfRgvf3C0WEjB/Rk/89nDYiAe56NIhWo
jQ83Qz8geXAbs3SOodYwaxCykqwUzxMf/p/9nDsRVdzwkBehKwmg+zMEhpS5h5ky
M5TJpTNWl3Nu3g+1ctO1nbJLyeJC/aJwZTjMeFBcYzJR5o1GFM3REdzAsomxQa5/
0dHTHY1AZUBhVMrVz4VoUQJkZGNfNAyafdppxgaQyoluxfBUoo9DgDjKA5NJ9cM7
vYp5eleRhemb9ciYXbayAaBQoRY6s3vZgBQuML7oD7BXvlrPJRRpTcGqp7gzptAf
QD/BRqYCu92asKEDlqLrp+cTgOnm8WnSqbVP6De9/vTELyLUR4T6gflqyhQ91SRX
XFWSPKvDP/ep51wLGH+tPW7pl8vj6SMzJROveRFmXhjsl5oxcb+3ZnAqanG5SGcm
gSSqOo7J2ntTNgFwDz5aRBniGrj9L8pyK/iMfbyOBkVktuU6Nq6NgJMbuNOe9U4+
3jLm3DB84beXIFnqwnPbzW5/S603KWrSnGvyeNB44r91uG7splk1Da3NV1w/VyYZ
dwVPhRoJOLLEQ2jIEFeg81d2ZYrWV+76BPwocgFk3tBG52t2Zxynkh3M0qMmJdTI
llXVkWN7rLmnU1pBahFylaJEsGAZ9UvKXtDpoDDSvPe1IKtMTqyjBk99YygKe6Fr
C72TXbfd/1wt6cohLUv12MV6CtA/Y0S06i7+6MSMyvbm66gAtWm5ZuoNKH7Nr7ya
585fHEwiEKPY3H5RnzbH3f2nEnesRVqo6Mzzs2ExMOsmab1dC+7avfkrnN7/XyGg
cmFhUB3RDsdDXa7zE/v6lc4yKX/o4W8mu5h8RJM9luTeuRNtxP5w5cmRHhs/grc9
CbTtqepWaK18Csu7ZzCZkju1MLgUBlWnpGE7CXKQY8F1iJyXS5uqHAMkN8WhaW80
ZFBjYxVb9PE9aHl8/mdWaAOgck/OCrggeS07cT4hDrsGKZJBte0I+SvECKjO8jqt
Y6bX0GhS19jNsCuKHDrmxIRmnBqb43MUoKmXqlEdoeesnuQOKEibryah+ZR4F97k
xbMkAeAXoWTKmwFxh9tJFpIw6JTWqe+4qh3fSjT4XQOW2GUwDyrfCZjs8jU4/NjB
SVUrtlk7tf0ECb71t4/NTJe/IVBlW/DQOtX8ybYq1lFOGIEw0hJ0ZazFySkOzo7s
ZfDufldODA8BUc5V8Esg4zqxwSagIOOaGaAwIR/FgVGNOEzQyD63dWxc9k3SNXd3
iAGzQ/RMW7HsWLUWdq1OccgrlZqDEVrqTEl3KCcQ1FXQDBbwnoycoKz0oWEYoxnl
8V1TLjJLz81RvDn6qDkKfDaCZIMoLzchJOdVkqpdPDsqUlJFgRgbRnsM7wE8R4FA
BZtr//fhkgx/Jkv0XQFJnIJQeVM+a42mzmTpRmPto3lz4/ThSFb4SX4v7fGmmIQB
ux54XNCY9wEwDj2XPyzWlj0exVoLKSVzQqY4IvtlWqj/sOWa6JvcDnKydLE8mzKA
hmxMQtLT6EL8B6+EVSGhuFXhJQ8YKzVt8Er2fQ3Swb1TrQZWr00FMzk5gtRpnlyu
Ely70RPKLRXggs9Y6V03WA5C3KQzVjaHXruhqdOchptiS3k2fI8swt/CfU4yTjEs
iSzcoB4PH3YpT8q2W8C87HLYsQZMF7Sbo2Llo886MWIeKFHFaIFhKJcbqjzjVIPa
XIs651wWfrDxV7NEWwfOduwzcOFsk4vDtD74B79FZk1VAVpjmQw9A+b0Uz/5tqCT
51eqliqMjPHFL4U0yni54/aaKzeKvu5Q2uXrmr0XRbuQ+Ef9ajM5YB9OwyEr73IH
+25EUzdalgikBMoARv0yW9PEKwwEGMQ+2ld/RhCO4VWBGx/HODiAAtYJC4rTdBiF
g4bq5ZnyTEr8dVVtmus/moHpnoDKgdVfpseL/WQUyEMzcZKYAQAZNzr5hiR+s3ut
ywAs85CcjgzAvNhd2hpmihjezV83SrxfxqB/V7OcOmapb03KvgkIFnG0E+1ykyQM
TnyZHUAX5l/DtplfNS8YNuBU+uq0Te+kZ8Lj7kxZa5umrIVw9fW9Y4pnLHAfsje/
MTbgEjq66kgHvEdaMC/CCQBrrQpbvBzwgQiKma8OFB6mmexesZgb7ZWaipdOeZHi
xBunVYQWcY0ko0Jff1kfZWR7pw2P0UD7Zv9Eo3hFajbKUyv0wC2pf8KdgEklrSam
f/3jiSzdLoxVaDNMrLvzNmTxQz5mBg7Aa/3Nm47bHQ6IWDRyenvp3E0JpJOSQZmJ
m7ISAnabud0/uhJhQD31Ar8dlUEbuHECVsqLZHNMvckET0gwJCTiDQ4vjeyHiDk1
n5gUADtEfkpoDUUU6NYeQgZSdNO9NnHaAYrLtVGqCTGILRBIT5atorS+Akd8oknK
zf27ZEdU/wakv6n81kNAO7bcINn4aZi9avioq6ovob3Z4ZF518eqGTueYI8E3Fvv
V4TvkTlgxuzvVWzlhNpeBvovFsYedYwGfi+wakjZWunAn7wuGpE3Xt8YhzbgbIBN
RADb7AmMDRB7KXvJXWGbVi+2c90DffbeXiXJvptoaYUOjxmGaDOhjplF4FL7o+eu
V205+FZrPig6zjyB9YEDSqSdRuig9uZz9GvFKNH1qBVeMhSs1IUs9e9pIGkOKN6R
MBli23qbFKMXKyDS2rr19rxKg/Xvhuc4UIzTyElVCHBz//SdsD7odw+/jRm6oLt5
xFoiyeMR0hNvbftGPQBIFSbXa++bJhXcbdpo/WldIwOWGOru5LxWCY6n81UYh9XA
OPIC83FyHveqMgDPlU9EYwEIDEOAFSjEBkeerNcM9xP3b4U4mUClCovOXSgMQ1V8
CBl8oFi2M+KEmQD2nYax6/cakaaPojCyaEa3GlOcZTSBKEgWQNkg79pFB0ReJzTL
XQPitIgWV7+F3zGBxAuF2Og/TjEcPwly/evLZOfu4Wgpl8+uzAyA/a3PuoprtdhP
R68xS3TBOuAY6zucvGmqC66AC78alK0Sx79x+epZMVZPD0djhyNBDWS1YXbeNshU
6f2PMQGgDRj8z5r2tZFWn8gTWZ8QFR4bnSE0w6CBPLDBNlkIKki2ZsmpRkJcWu02
g0Ms1PC8WCBTwVVFxm4jJHgKm0NAMmBoxkQueKp62VxuaHNe1tTWWLvbKXnDJ49B
7sWIKvsw7JjMUArxpCGQ6Rn9kES4Lo1sIBBjRbzDiq2sXfxtTbeu5J48qhJ9uBEh
mS5+BDMANyTmB1v0MXjBlsud54arjZIoRv8oRR9voQs0zrM3L+90ffzz/O8eSQbW
BnZKj341dMA4SR3tyViiV+8KSRMXwJXVvW225XIcnC1IXfPSbVemTBb1aJiFhhdW
p6ZMJ4f/dDQ4K0xge0Mh4y2UKqjhVZiZ+v5ZitqVhpNc57NuHWeRCBeeZ7E3ZTPf
em3Fslhg+4zdVkyaw+EXwO5lncXdfKUm0pvQhBOp19W1i6thaidoQr3sswWqQ7KV
j7QOYgTwKpnm1CRPMuUco0DfMr5gVpM0zikg1WXZEDjrRjerZ1svj7N/coWoY+sw
0i6M86vfKsGnRlwzXuQ7EciaMjSdyXNHXiU7Y5kHsSM52vAClwt79umjbZeSbKjh
0dvPexkCukrGKD947DlTuPHgGg6VWdABPYDpPLqwATFmrvcex/hdmYA9fJO3uCmh
Tg9BowGUmu5u6q9Au47ajPISAxYtIEXOQUtiBA4rXJCKoNY7KqgU0qLBro4xlQRy
25e2Ef1/Gm1ajbc4xFsSunTFwmLvK24sFVL0a8iNdNCMsKzHf0DxI821oil4M0BT
zUi6kfiY25WnL5N2BojgzcS4q6WI8vR/phIhcas7NfdEqTJFAt48h5pb/SV2fwVy
pGwt6KNIDIIF4QjFpIUmm3EoV73U0nt35BKznEJd+lO/DqV+SFfj9llxEgwRXvjk
T3xIEUZHX0EH9toihwHoKxzTxJMuz3ZQycQox0+ANnTeICtUe7L7JTr7beG8mDTD
1AUUMvK+k/A89NARtr8M85PnFCZkZF6yXYOPRTWR5BNC8nvzQ9eohDcQxrSqOZQP
BSmQ4pNDEfl9oUMYki8JpcHkihawf4NOMRJre04PaGxl/1iR1fRlo0C8/GB7HvAk
LVIoulNR0cB0QDnWzvDuti43uyqr6ccHBAgIzOSMtHHs+hzKZalQVG2MEudIct0r
46OMDBNnxdvS7UTZMqO6UKiIqQFzZa+ACL6dWQD2VgJ0Y3urY1cXRG1HNwoEbQ5H
c44vFrm4V/5eEcxPi3Qj6vA05q1TC+Z53Mj2jgT76OtFZ4DEZ0+kViMR2RHG7fG5
sYmXiMseyE2N6RB8wbVwJvk3UwMh5w2FP8dJe/EuG2uDzOypkA6pFES0pEsz0x0G
0Mus0H6knY8TlknDexG2c7kzzjBSlexmTOvOfcalgwb8FxYfn9Mkc/F7AK47QQm6
yNh8gX1diQRQwTYi8zEM2oICOi3vRNMXXRNI2K4W2a/2Yqi1F08M4OsCBEpTInuR
Gy4/kpYJVbNq1toRYxipfFP9qQW4IIrtxhf2IVqXhPgxP8dkPvxpALJj/GBcDUN5
Zo4ZwhfdEvlnppLQWja78EkKPa/cBs8qm0D+EzQDdLisDfg0AyUmojI1yiP1myCl
tEfQ55dNPBzXG+7g+1k1pR/lsc2jwgIIdcjTCzmOPtxgQpJMdl8bBoaSPrsNTZSq
9KZNP5rWT2z2+rxyfboriMX6wisBxeHfvO2mwt0ZkAJQTSNcC9u/QB/nf7ocAPxj
Cp0lUEh0uL2POw4GzDwXkvoefNszmNOx3b0Xd41zpx/7TyR6CzRhjZN9g8fqfmxy
72d1P+xBasK5kHTU6xHE8HT23ktxkBU5qHpneL/1BeTEXdCE7E99rbtlwkIUWDZl
EOLJ8+UDHwCxbO9ZewdetxwO+DMTc0Ba1jNQNlN7Luym+X3pgHvEHmSAdL7aj41Q
CTr7YuYaQSxOAr9/FXR3/SZw0WQGun3FGcSn79tQniDIup260k+Xvs2rSP5nYoDG
3fVs5pEOcj1DcfXg7yK/AlQTYeISzG7HjojaNTSJejPoiLLmM1CS9F2M3be0XScK
/pmjcZOVGqLG5I0ck/A/Yff3HxZvmH5rbt0RXtHOQndHDJzpDvbQmON+6xjhYgeO
UfwE0dJVSzQa7jE8zCcHpQl9hTQFFlsw+/nv02JPPQA9YSW9Rsc5inKoKOJtYYbi
I9GfITQ1tMzr3y8GsxfkZoVR4DSAisMhHxrlnHG8rhOKAlx7LWXBXbR5yfAM/TSJ
gci7JfkkH/u46jwWfrBEyP5AD6+9z2Jad6g/RqdlXvAulZHpnVcQQeOCzxfX0ScB
8f7ykXyUyyBLA/hNvuwkA3ni0xaHVIN/lr50BxTLdV9sSrPbVCLfi3D8GFV4WjCA
adFFqQdBT5cHoTn9e8tDBOl3ajcZFqIfgDotBk6eruk1jJ3ihCPc8QUdubTRUVTB
P1I8sb7x/RFNnGRsEU5Rvi4nwJ2gQ0C71k7FahWxGc/0jAsotsOM9tSsyzjEFa6L
5jCmk/Z+G3GF3Wr1shNQNr//u+kqyN4CqqCSdV+k6YZaBb9vjdUlKW686QesK8BI
NIvfb8SqtAGO+cFckEq8OTiWZuU6bKrtylj1tNvlaEzJRqRLiXVOVoKqdWkt3n4o
Zc1shcxyMOl9SGRvzHoHEcIafwRue0Pp5nL0Whtog1T1Uu+E7po/IqpUOoP3i6PM
xm/GAt4+E7eYivkNV3cmpVFQKU+pkbCwitErpG1pPnTztxZAx4KUfgjTkzXbP+mw
+8FCsFF6iuBjDC0T22RJ4m6Iz5jtd7maRQA0lIOJrDZh8Gd60jWjMKcy+K1oCJ5+
aRRS+nLLOt1uC0AHWfgdsuK2lx/OWLtxUrGqwCEqAl8GZ9ubvkF/7YPJL98hacih
rQTnbUtjVLOUbl9AQjnNdcAxIAZgNDh2OGT8/oM8C37lSGWsCHF0uF+yIq8sWdaK
0P91JCCdTB7f2ZkvK3pRdsw5qQ1jN8+QGUII5C13AQpQo559KDbKzoyfbdLWRIrV
N2SAPwIjmBvBMVSF01rXKCQSLhet1wbi8lcGLdiM9vibExwngkwGpy/R5lt+V/PJ
ofLFRhUVC8d7oFtbUlVdfIjATseIBH1iHj2I5CUJXduxlgKlyQ2fDFcwmhH/vSL8
wIZ9YeXQayNXl6qhJofMrP3EqwDi0+VzOU1akqSeCU/wSjQlqotv5ax39JFzXPMM
d08gCdgoALoLv9yEq8uzUFeoE9qVt9ghtc7TLqBartkKjthFkhhFFTcp8RilvN0a
lMLfrCjt6/6bn0uCxgeA7FTxxP4O2cLR3MT2GRFK1mEjJmPeCvAwDY7WDjyX3YNo
P9zh808OdnOMK0joaCqrpiEwz+Oovxq+eEtGkoey0orIg5BLt16eospYQX9eT8Lg
Bi7F7XuqIoSVR4vh6mWS22DMnewJjUyJthN4ywtUBsqlsBU+vqeDO8UX8hgUheoy
pkDATipxOmguO39FYx4WzM9UrJovXf6v8tk4Vvud6q9QgdjWicBvN+AdzdpUJkXY
gS1E6PHOz54Y0io0d/lCYezYIK7ZQ9zVnpsyRw+ZR5JUZSDaPiun+6Tu2c6AAYw5
5IMFCTZCdAp9o7tZFOAxA/Dr1VkJ+gO6IwbDuW706JVBJHD45IyjCkh1/L7uuRBu
8wEsyRZFjzDtDW83L4CGvd2TtTXGHDWRwHUqFwV/WBwfjLrLv7aS8AgczGqOh7pO
V8OznKBRu71tOWYEK3wVKZMDGZKKQgOAd1DIrZBkQWlCVjExGQ9mlCslDqH/soy7
vFDvM8jvu1dGsU2WZAyfkVZY3CnK17wlLu6pfOwcjLwlKUi9P9+31FhCAQHkH7xf
0gF2XwoxzBC5VAmES6+eVNXj9N+WEBKPhhPZ6sCMG5jrz5pJWYbd86h2t4HYfS+s
1k6jDuK3fzQ4yr4G3I67kzvy1GEiz40+ZfrtZzuPoXPpuI6YJIKjJjQnwP5eCtJb
+blrDFQzg1OyrhPKFcH8coXnKQKamt4K2G86CX0QcGQGna/Qelc84fhZULUlYj0D
UjK1mBmnRHNSIu24bun2A0/t5oRfihUZvXpoOPb239ilYvvQWJ364Beuwo23RXjz
P1HdRlGI73VEpZO3P6k5xbjxBaBmZpZjOfI6Axb1ktlgHcHZCu9jXrREpBRDPpQL
rnKbq8wT1/1ds3YgSVFt/gd7bRlqSjR5C7werBIs3X2olDBX2v5Yp9nbtoIFWxIC
NuiXGyCMSol3FbNYB+Zwh/98iZ2qSyo0wAq2lMozDGg/UEdyhCJ7eRSgq1WZGseY
SwbQLu12BQnAT8/46sw58nJeJLWFsoKbyLUPIn7TI/8k1ZLCu8gr7YqMdPg636bn
12+OLPzzjeaO3WslZmxw69hPmu4PPjuNAo1t0WMvzhFn65k2W0cEG66hPRk0wYjh
ucNjrVmLLrgQzDp5Roac8HCzW8C/uK4hIDQK31YdLX4LLloW+2NAwjYzgdkmMnEH
ayXRVb1M1FDJ8iSs0xOGbQoLCxKnx3kv28kscLPSn/HSZmA7PSFlUj0CDRjNwpt9
66q7T6PvqVH5RJuuXXZW3fXZO5FCsnHrEd/JUh8fVN1O1JQWbPVy7BFQPbNmUTRz
TwCgDXynwy2GEoZQ0FKYIF0pixA1oWWjr/UI+1eeiOmrcCkSS29RULUtGrW+Iacr
7GH8GdzF7uDUjy3VyFtjJem9bPRYHcUTSJkbBenSdxRZiqocTpoR4n8DTwfIJ5xf
0XzxcAAji+J82ToV31pHH2Yy31UBFPfmV5DHp2DMPDa40+vif5/GVNniyH17LaCc
6hfRN0yyh1YBMMyEv209f9X34u5Q7cHrWMZ/BM0IaRRBrT9lZwKIG8xCdzaIl87i
z7hGwf1f9WB6KAyNkD2QUdfoJISYo0ysEb3ojTgggJWUXXIGTn74CdhbhekeiHcN
9Sga4XvBQmr1QyhEZvrHIsyaUwgMEuwywwngEweqH/7St34P83Lz5sZStfw/QnpU
1JE3JDo/OvWgGyHKHT+Xr7bmwapUIH+dOnXXD8ftkxQ/LBjsHEn62jlAbHFWWbWw
+h7skjM6L/bY/uJrlTMTSmIN7sTIlyDfLQAZC7McuKPWc4Hcag/dASlsvUzaM6QQ
5yVXM6FEBsGfFfpwa8Ze/Js4EdxRImUt7CGYOM6gxc+CvwVubH5eG9TmnrDV7d82
j27cSfdS0XI49MndaOio/5uN8h+yc768QrfPT/quAkWDObxCrmerFm/yhQzicPS7
gEtjaF7f+pc38qagS6/blp/WI7UCPXH62vfL5/jiRIMp0wglZEgffWxBz6tOvYIt
PVgNIpct4Q1LApXJ5scaffnUIkCCbcNfxSXWizNhAOjP/bccS0ToKBXhJmAAXwNb
OzgxxNdBopkMZnDgOabCZJSTlA7kjn/Vzyot4WmcuXAoBmf36o6EgCLPn0zxnYM+
i683bZlvGvE2wL12WtTOFkYsWF3sxqudJMxRlM6y8Cfc7QEDxnuWXHZzjVLEsRD7
GmUbcdIYcEnoTV7Jx7tS/PH6/Lc/Ylb3oAHcDWoMiTO6hlbCRFqbbOBdPW+Ei37O
cIOfB+lC7EQ1mkHFCa0qbHy5Wjq9ZjomIX4flLaRPqqYmpELOehN9Nw0ANOCHDAM
qdxfJfoRpzG/puL9tk8rPsiWzryuNnDdjEdXwvfUpiINUxVbFCjzmtm7SEocPnyq
7MsPVPWGvbhBoolWUZmKRRSuSMveDK6N7ghvFoW7SEaAPsJ5+TbM59Ia5TbAQwbH
zvuH9LnBHfom+5KIGRUp9rMIfTgkSdvQuehmv99l3KdIdgsyEwXfoMZ7soMijAan
7XYrRP2fmr0iYRecwQroHsA8UxRgqlL6yZ9bCatrzNGWAwdF8QhFeWgt9OGJ6q9M
bdalxQgLTfKrsQtlpvPAcHNNv06qJiBCXfg1m9ZV8FXXVvoxZDByN4+CFL8qMvoW
RuDvfV8NArfYbhAWIiA8A1nmtHbcjZaBZgr/FIJuSjLRkR+1vTNR+xgqCNBXs+ah
bpgRp+znoCihpIm4F4fG3trjcZZfPXA95TEOmgc/C+U8BlUcdJgpVWMs7hNh+uiY
qMYqA1jF311iR2ttlnxah6CbQaq4vFRtwEBpTgwy/By97aHogTpX/FUiEDvbls79
WBaO0R6NmXANCkru9Eo/JTjPD8giMf6alEGBA5biyZ8FNAEvaJ/vZ9PkjteCWlj0
mo9XKkkbAN+WWjng4zVB7ZV8+fQCZ44khAoq15cm5jg8FgR/pg6Kx5KtIvf1e7Sq
AZBCLbmv0VByXv43YKH9aoXwerfJSxTSO2x7XNWL4fQovo7cboQ4pY7IF2OkU0O3
BXKYiS10dkmFxS8Fv01pn5qHN661q0gSbjvYpmOoSNq+1j4sGHSOcKSNEwhcMy9d
lshIY8hD2D/HQnpSU2t9NV5ydeaDvQuzfkTujcwqBCjU21MYWzHa0Q9sI2yZ+nJ9
9nT3kYrnica5UsMcYgOs93Cf9CR4pSw8T/1r2PHvg5tSRmlbvYt++2mq5qRSwY3F
Zycn3+N+7iDfGvMIzh5Zzp0BclTei5I7faw7twUeCtLnV9uRm0ar2gYkvJyXs63R
oFiwrr2XEucrEtVa5Zq/nxW7LiZWI3weGx9jgrQTG+TkaxLSVxronm1l6sU+rdPM
0dRwGx+FSFFy6mCWb0H6WQf9IxmyYqGqPEsYnUG0YC3fBX+h9WRxyKqEd+YQ3p7N
ICPfPn9kW48BvLe3KGBXlk5ivCD2hCgf/kXDzEN0AkcsERVvu+mNeCkkUxrQh8GF
wCKn4cxCeqYVrYO6d9UJ3/Lkxdqf+5KOMX0FZCgqTqjTi6bwD/+za7PUXfHgei8b
0O3j2J7nXftlweqScw8lqGnlsUOUdNZoyaeMTqtwRsI/4KxpT++V+AioPPLt82q4
T77JcXiYOSoCb8ZwI+2QXJ/1WRzJQAqQTt7IDA4OtFJZdADIwBAVaE9/YPTHlMig
OuTPRbYHhRBoJuTwVLRo0RiMRkUUZL0q4DZ4tRYVXpJZed2QD0QGnRyBPYYazeOQ
deabPnXCANuSvcgi8kLD3ovP7A5wCS9ZjqmQ25Y2ala93hxWVIOeDqF3IzRofLGK
ZOVurKNACfmG7yIp5ojAwmV7XQPeOsGipX8KIgiStNIeaQsvBvX2AHogfLE5Vxfi
ss3DT8aG/TwKzRHc3VhTtGF1S7anyjc7ZuDZ5Wj49ylDrGo3mU6PSsNf0cjZbCJz
pTV80OsBwqUOJKvYdPDP1DxrCa67bsfnpTCyGdEc702Ry03uQsqdg/T9bZXudmR6
yoLRNKOedoAb5GZSdhafreIhTrfydc85wRq1XlPdS6x4M6uctez6d+75QcizV/MN
NTeScL9EoE4mC31ggRIr+xFTsD3ZFulmldG3m/CuHipZWFu0c84R8FqM2bFflO8m
wHj+Wu2AEnI3PwK42ptaOUeWxYP9ZlTGfoyxfjG8/+tLBxvFX1FFwawp+C4eyr0S
ONrKTFmUbAP1+9RsFsuNonCECptDk4hqf3VVcX/t9sa8/Bz5Cs0pCVLKVwCWxp66
Uc+THWn5uL6ckYT/MgH9+jKLiHxf52ns7nIa2tQisdWMbSSM5apnZ+E2X3XwWPNP
1+SEAgeyfAh6akMPWkwJGCC6txDVO0gGlASQ7mqhM6be3RDmAJKobXPfvwbCCtHZ
tjVLOUIDDz3W8XH3yYWk8qfG55VEYZaApY1yW1LvkeUbHvYl2qymfw/VqZ7CI4pb
7ZJPEUaGbEN3ybvt0X7IwlPRARfEmOplZ5fKlWValPyDQA0Qr7Qg+NLpm6QnwJwh
a9E6+M6oOF0dVsSh3i1fizXhfXYeQgktNevy/eLxbwB+WteT16ZxewSzeruuqDl6
GWFsC7IwxHQxh2dawZn50yhbvi59i0HTysezX4sPu0CYxSIqJ2m7ulBb+7GZ5C/M
RlnNCndBMXZt6Yxo32qqZ9ZFgJaVcyUqe5SoqFW9N9Q1d+ion8TK0DYPiP53Kn9h
1zvb7n4Gf9pnv6za/M4+INk1fBG6qEqxQ2fkdjocOYaVI6HJ4fNa6qUKwIw9CCbV
ryhb0OqLIhpVDAbh7aBjCOrFQXutzEwZ7uYks+DlDRSv6UlfnpEzZQCn4Fy/Fl1L
B6IBe+JpH7txFJuTItVM6H3m02EVlvLY4w8pjKx7SW07aKo2dbqiXQHTWV8ilzjJ
OdK1wSgTqN5a48fEHCse+lp6lbARsruI9xjAZOdyfA8tW7seNdprmm+S5m9OAYGn
wg9K1Yb5xkzqCAN+tEEUNtKje3Y/8abLTZdNRc3XsBDHBikPaLTtKH5AaJlBc1Wf
4mBL1yK/62izdxY8Pga4oUK49J24dwnWh/fq0QACnRFEpq2FvshVYyg3uzNb7N68
voJ3zGA5SKmnH82WdiLZgUfHjJo10pHury5CK8wSiEpLY12jfxo3vazc62wJPGy9
NaYKqTIKgnTUo/ZtxT9mO+CtmRhBxK7o9x8t9R5dfVd7hCZKhsvF7l2+d2ZIAHW0
7YvBUfHjrA+U1qYaGPynGdiA58XecIZsDoD/5hRn8U0yrVZ14lv9hv/HJ5DdrG8N
Pqw42cFPKdImc8cPHnG7QoFrdE44bMN61s9BaDdu3O2aefw0rRJSISaIUvVAe9CW
SENXdplg2BUSpnapuRtmYFyrA+3PAlQ8xTouIDpOqbAU7GJ0+YYDon9EjxD9lFFd
bd6nPxzWvC9j01J94CPuhLx9cxwyLfbAXhyFBpB4gNflbe8LHrEK1rO/ihRxRplI
z4bIbyYrKhnOwuC0qYwCQDy2Nh2MiM4Z6DTWb4zIUN6hLZmwuom1SkSOSjg03Sx+
0wKJZDbiyJ14Woj+VllgicBY5o1HndWTERpkK53FY1LS8jvXlhy7gTHtLJpxef29
PJCpdNZR0TdJ6LeotY2sg8Gb9zA6apcdSqzpTl1DDSsz4iQsW+XXeNVB9S+a2DAG
kFuciDslm4k3be1UOqqsCX0xYJa9qlnsaw5rqat/vXatO7YhHgjRvkp9/il0ZVuC
drU+80BrwhFtFH7omcmQRdYxcHkDbhBGrubspUaOUq8ZI3pzAjsRjk420fNSxHQy
39wIfWUF2bcLTXunOzGY6eGznra6jm3jEXQbicTazyVWeyOzd6gfZQw0o3ByJGqY
ZO/vg36JPDhdJOTfDXAmBxonSsdR85IZ2GHW82FTG5nRiyyFqDOC2m9wVyLlGJz3
bu37kzS6snfnksaHqgmXtZJ4atuJ0lZwReGzee2nZsyLXLy8OXuk4RE6IEZ4TSGS
t7MjFPBA+tAm5K9uaEMlfCkzmr6QFrxhjW9cexO0IOs1DFONEhA8qRgqQGkQ24TW
Gp1P7lPbF2A1KUTy2gLf9gnWR2LxkK+7JNXv7kAsIGsFiTc5r27SzD6DL5Fgl3FP
6ev7L62uoUDqX9V/NsW+1yQZgANmWKr0j1hvILMOdB5RiH5zR25mbJVaNEZK5zqA
H6f/iLH05lttkx0hpL6wQE8h21aZw6eazIvPzXM/V9yt5yp7zi7NPJCv1of7oxh6
F8kejqXRZ00gg0PhU6/7YeXAAfXGbpQGpbmGyAU5U1tssXM91hNnr4LAPXzL9W1x
dOCswGHAMutMziTTFAw8kYTFVpQvqOLQuWFsQ28dpMX6a2G8rhheDcyZcUqNUB6y
ZGvQBkK28ZJGwNrYW/P6P2QgQgVdts7ftLi7kon+AXW8guBKSrq/nryfPjo/vIDK
hFZeHFa8507TgurEC2PouuEKulbUoImUanU/HAA/fZ8oA8CDcD5HY2l/Ll5CLXUL
pBuLbxxhE/MUjtzvgVt5ZTVcWMT5gPV95kKYScSVhq2CbqdWFsvE17tgHx9KjHeW
7jAu8PVNJS/Db6RzE+YDt51fc+aNHrdmEP5fFeTI0EVzOK3BikBEqLhjN26btAOV
RCLfz8lT1+xkdw18gWtR5zwQPv76kpHw8GxQMrjAZVNIeQmW6HhX5KsB1l/WQ7ts
Ar6RXRVe8jngbv7yQVIJoL3SlPbkriMhrPJgAWzEw3Aege6jnZnI2PFupMBAAA99
w751tHlsm6B5tL/7GWeE4UAdWUAEp20B1Hu+sNE7jQx8RCHBcM6HPmdVN4MnzDDs
0+zieMot4/ZYM0jNbisg0zdne1ckkUaTN1aNr3iJlwI8wMl7Kz8uswJ+taMxP+bC
Xt1nbLzuX8GR4mAa4dpkMX4icPXo5qFoBvWE08kKKzJXCGZlL+nz3yOhCfp55Zks
hxyXub4lzG4lYuk/IExYOv5RxHOYqd7CXbBoRbjyepwKX3hiaiYeWd0KVkZ9muCO
M/0BZuGUZAzUSk8R3/PGb0XNSDSxpMpjTZJAzJzCELKKee7MpSdHsbyOrGvykOht
Ts3Isd8LyA9ZhV+7taENsK3RZZF/jWm4d/GAS7njOrzQf3YF6rCsaG/Axojrskuu
/AvPQW5v+Ln/LTdDPOvd6obzLhodUXAjbsWlY4YJygzKF9fKXBkL1Vw6lvEbhuQu
Uu+muHclmrggZtKfPABR4LJAF9cWJuRp+zNLhGoYpcESKjEVPbsnQLE+4AaY0svh
mINbom5SiUgAFP31zA23eHym4n7oyFbWLhHk8u0bezbNIACkmlg1VKbSJly3GGrm
1XEmgZvN6TWSFo++fVf6uDJRBfDNpO4oeJuCojHQSsKFQ2h8xjiRwRT7B0kLRVPm
3+KobRX9cub1DAbQix+9GC7bvz71AiISIZKMalU2L3SAyDUPVrn6RQEGvptasXdz
45ZHTFexXbtTuKhTs9iN8I10sMfkPiw0ewvVJhejbIC8NJ/RXlOCoqvo/MUM45Fv
1hYa5K4Ni0AEk5f7BDRR8RD9pADLUVVyYosg/Bq46NadBHh/bUgPN6MzVPIcrW+R
4z2e/3arf9uHEmQPhYaAKStLC4mXGTn8cWkXVKUgiB/2fG/mDW9PzYgpWzzvBWtt
dSHNQyXx0/KvJP88omysP0k06vdVTWyU24CFlfuFqHeAPv9S2OWiUgJa5bN9XbMx
SeqQ6FSyHlkaYTAojl1ncqqezbhlqtY5tSoTcOTeerrxwzPuXEKUW482lBd7aP2t
aDrLQV8gp4Macmuoc66NB7FgN/UQI1SLzEAI+09Eosv6bBowbh/dEF1L2wfZrMzk
IklSrxVPn9RjZNKI90/KC9PBZXvNr5Cwl8QSubxnBltAdqvP6S4fgk+ZZTArkDVb
BXPnPHNdlzyOBdEzRsuOh0elQAypxA2pA8wS0zcPpDJGz3cvCpCXbpBmiddYKh4a
cfsrzT3BBJplXJJ8VY4/r6jjvBYjThkVW5bfyep87q22b33o8vVyFbvD235q0DmW
1vmWv3Ex7ESiaMiN301HsEcJS5xehxYWlByrXPUKxJKtWZ4cGk+3ABlGcum9ArUi
06UMKWaNjuvqs+Inp7FvHpZ5YyVlc32KL7YFcN5YudDOxXaEj23qs1puCCjWa252
DSMCV+yQL7tzyeZVnFHZy51wQkk9qz8zYHnQpuPGv0RSgkqFLjswZC8DWQf5E639
80Bzbz5AE5ONT7/66UQ5/TShJCEBjAg9KT9omh2+x22gzGLjSbuEr48uiCVXOfSV
Gip3BJkeyxs9NgEWh8abo0XQ+DfIE4HuEF/TGRXAreI3y4Sv5rNVZNT+PXJ7z1fD
Jzl/r9q1LSPpEWaa4G/VIfM5GkvLFKp+nrSr7MmONRWsHW8+IPynNOjLC6SeM7oG
qmqU0qQn1dx7CSJ/dLJdbhECj8Q+GYpj+8CLQa7arfefmxEHz1yzhqoqyEJUotNg
QeImOPxZrSM6+/Eavytol4TsMH1wMM04LFdVaUIHS3v4vIXfADY6RSQyCAF84Nsp
8lPWF6+jd6RLrQcHPc9pfnF/fb2JVPnluy0FnEY4Ah1VwKAyEDD5ZsTqLujYxZA8
E/9LUZ2h0uFPaU6HV0/EnpZrvsPkCoc9LNLwdy13W5aUZApavp4V9Jccb15ugaHx
89p67puEZ1M/mjPubCZUhgZPDfPKqmQs1kn7bZdeboJfqhwHnqwyMgF7PhAHNQ07
yJwkpBVcCzubz69XJrhmuxR+/8xXWSa8trmrqgPsWzt6qMnCuWSfiYBR33inhLte
WcGyK2pW5HBwTVUZDakKLQK2Y8s6Puwdv/E0x9I6sAqzgnA3Q8xLQabWDnxL5/oA
f3SyH/prTEaBDy5GzzNEDvix97t7yVJKJASFFn7ENT27cOKWZ+MibPcs7NQsE0iz
oc0tdyj0AgiYKiN0489PCefMU+4WukQIwF3oVBflu5vO2l9zgwkAr8Bt285e3YRO
p86qFWG2O/kwUJ2kihuSftDv55Gpid4pJSY7NlvCb7ToAoofWF3K3799K+7AiZ5h
8rDts+Ax/cz2W5pxwG/CxjAzqKq/CckOXoP3f38vtuGQkWgVVk3DKRo2+FVvkcqt
ZRn0Lmp5XXmG6roAq0Ls96Yob2Nj7l2hSooj+PfhdsWhdWQ4eGJsY06TKwLjvuv9
0FGQGzllglXCn7ygw6i+/fhZ6GiOgTyGPXzS5yOdz1DltZcoG/omSnQ5ZtbCBXjo
8u/Uc18u3QeU2nE5yGoSZx1f2+blAtw0W1bszOV1nbeP2HKJbjJPaKCX/gZ2XasR
wnkaEBh+Vecdua1W4tXYXgQtl4bkJjzgzDxfO40cANckP0PiORRNwA/8GNrVXBI6
vD1L/Lv9DdjvojQ0SudlnfbPaADYKghs/sWosuHTv28c1cs19Qx4kINqF9S5Bc5K
o2d92yKKoNboxLZCmdmhbSd/tPpkmqCink0dlMX50NsfgMPEGap9F3Qtz8gfWSq9
AAQC+XHQRFYCY2RxDc4/oGcQuDv5DnDF76omFzTbTp7DWYHaYGu3esjT8F8klCBP
7FhZ3RZS7qVvigvIZcueb6elVj/3mQ7lYEwDcc6Z1NEIbBio6bk6OmMmufPvkKf/
yM97ByJJxnInVGFPThEXDIadCi8RuE63raOC4BSL31+zXpNZL6Etizy2FOvkaqx/
kDWYORE86oTNSKcMyLCq4lnVpVFCYYUXnmDvvDwroFG5heIniA1HKhckzszDFzpw
iUiTcN80IYltz4ovTOFYX2CmOPteBhWYWxy3TlLR78oAv3pFvoquOwiWS2S4i5kz
16AaVKwJ6wUwTooOMlB9ms2Z4RmlADeX7UBRZ3tVG4M1+hNBji7VeSoiy4jy9x3m
4BPE2zU7nhW3IOxryI7NXEWOIYvsUsRL+WLAEYSARxhRsHokFz/4fTlbZtJSpEEn
FPERjYHjxK4xjt7j6WyfpLoj3sz54Irw++snrEmxKm2S0kFArOYHHqWnv5Qy77dP
zunR1yJAwTw1PDoV2FOznQ2YDKr3JrxQi8WTP+zvAcS0W9W8AnsZDWZK/cQ/ufHC
3rVLtvTD76DIgOVgA4ET7RJnKpFYa6zalJyDV9LOI8H46YbecjrfkeReFn7bCv+V
ToDmbDgCeBeI3JHSVK1OgkEEatz5mMi3fkU7sJ7+bWHkQxDXRkdSlf222N4X23LT
SkREGgJRyDe+dOmeOcwkjz4TnX5/B9FxQX84EVgdPrwtyW2MKw03JkK4DL9HTuv7
R0PdX0plWiZieQsGyjDfmybdkwHY/7kU+LB3ynGbidKLj/aHmquhGl6cTSEouVWA
IYfsdBhDjvpvViK98U1RxpL6l7AJrFna35SlZrF6xVLIqEzhI8ZAtMggEJsuEMDz
+nKTaZt1PVlAklDaCVRmhmCxLiZGzjDdLOCM0bD9L3dQT4sYM/LVbKfcWUG8X2GT
EIf6se3Njkd4TQc5ZxlS6r+Fj4Lr7xdaxZQaB4bVIXZsfQI11mGSna4q6YniE9Pq
w3iy1q5PQt/sKf6DZtAb6h/SNrgwvIkV28BjlNIOKc4oDfSPNKz4MDLerueGsTid
sQucXONtP3MJHB+jvy5nJafaIg6d7fI1HEsFZp77ZEWPtjGW91wEaeihjL6uWyKo
He9nErl7N/tesuCMPLLfJWx6PN8tCjp94bTqqD2tm330Cf+T0SXtcegkLEkJ5Y6i
iN6vZLTryB/wUg8xsmL08RCi0x+4Z0giSJyR6/IvC3y7w1blm9qvbnfxBXSU+b3c
1AE/QV/13AFkbd+cSkdtALQ/0SnPVXH7UdI+G6bRGfFA7BPt4OQ9/qQYxTFta48p
q3DW3DRTu3uCKCqtNoFJcWO9PvPFEwLi4K0g8ciZEv3h2RAKhctYm8Y1kzhTBh6L
vfTEOF3GUkAWXM2IQ76BdJ/LSaYfLZCJ6lL/iTB4v8ZRFKrMuf7HE64pV2P7rHO1
qqQW4rlOaNum4QpmGoIbrkL0GbIKUWogBJFK5Xv6y7BNA2eUjtMPK4EF9CDV5H3H
KSctoEzpGCa/c0fe7xPRqC77FCCmhSN1i8cRCD5fbPGloh+pxz2ftxRdGLTrjF08
HTG2a5+FSBnPJ8rb0rrDX+mSx36EnrKfrY8fMLLzsZNwtIQhmOIdM4OqPE4FgGCf
ZHCRpxHSCnakQ4LW62gIQ5F+TPxUfv6hXS4weI96JcRAtUmaLfkBvrr6S02OYDw8
WZX18+3O5uAKTRPBgNiAqmbD7TllGFELVN716EhRnQ6kpNOaS5nqShlHQLWIjmKz
rFaKguZeRS+F0UdXJ2QwMIRyDfytIXxMglDZ6yOWmqbnYEIxoDmMxPbqxIJ+AWld
5fIWMOrHKoa4iD3QBcTwr02ifOlZiWOIMWMLDr0l8/F5/VPNIyhn8g1J4xmKZKaZ
Jt2vKxvcNycSxzKCpDvtMAzGkkfrsTdIQM9grKCW7w0MkzzZ/Rxr7Vn1hp6eFnQT
MrzDiwooRMnXVLdmJfEg4T8XRwrKfk6kRUrllfI8KInZI+TrJ4BVQ8Og1NSldd7D
IKsqZPjSCTao9r1TSIkbeZ68t3ZpfQKGUy51tGYUlaStdMKTl+KicPKrkncmwYqq
6jt1p67rSOyGwP7/KcDe1WuOZrzzAhhZ8kgXbusnEyEMbvzA/h+rHC/PFq7OxRJm
Hk1lUnUudN3BHM3QfXgEJAFEnXNI+HkD2IdH6m8dqhmBNDf7xIFRChdKEtAMbupH
QG9shZEa+Y65RU6QOabdaTYwunqnAWqYWnciwGp35oQmCVPIMaon8KnRQjdxj0Z+
iLBhrdoNCm2rdr97MnMSery4nwdi59BuJAmJ0bkTU5UHw/AsLH5EJ/8WtUifblXx
F9J8mOEsk7D3BcWrLvP0lkTP7lZ0QzGvFLtBx6TGaSLphJpIBqO4adSck2l37lTB
+z55kZTWTyiVIgrdjhsLuj58a+nPqg/OoLaj3YrW8PxsqDTjgxPA+U0ywVtdjGMF
tgDUQ8RFYOnw/od1D9PUyL4/ubH/wzKw6plQmgxz6wjz5HJkfQuYFWaSZdIYeK45
mwzts9MsYjGbG74B5nKqQcHui2Kv1ekJaJSZGjRu0DNJ2WYNe/ZJQh5j++uaxU9F
5cMy+hLme2bIKZO7SBBpHoZvH3+wUK3zna5/0yFEkL8AS/jeC7O7p4GeihyFbp11
mqgco+GqAvhdmkc4XGOMQK+oxERJLRKHB75pzRRTxnzLdmCAs4OeaPo0meposEWf
w+cQ+ysYVZ6ZiYfI/gRlHOa20Pgrrv/R+hVFwmpIuk3z3u5teH34D5PKGbc76xZb
3lnssorVDcwOTDNfNDopKhcDasFPN1r4C8Jv8WrfTkHuAqWwLdgGn56JYr7ZeyDh
WGwNpmyNfsIobB5bxp/LLs+rjBhsmBMAMxxGP562xGuJ5ObvbmvxzvbiV3rVE6XV
hOikTqD/FlOpZVi5LjnFGii7ZvnfQUxBw8xUPKuBYtjAPkWtwXRUSWy3cQb364k+
0Fy2GT3GtrioCoJV5D1WMkzjwq4pYHrJkQ1xhXmDxsxLbid7aRooS656OZx9e1Hy
clh33qOUjkLNsOBG8mcXG8faD901IvC822r2JatqZNq1R7T1XNkdT0WEvCakvNJw
IlDysOJiyiaFJY+KfsG7Y72RAqOhlLg/iRFs2xSjOVyMgflOwXhjO6kcPtjgaL+P
C6qitA/UzFB3kWQvD2zhpcgRhC3xCSAg+0sIZctCPLBJionKuQ27bI6Dx+R4LQ4L
TnJ/Ud6YRQUTHqjoJhOfER76M9OJDpcC2FCT5/T6416x9xf+o+se7h+4wzIgncLl
tGULF4fOhYpxSqSotMnIXUwtRHU+2aDOd4PwfSz3fzz7MVElWfJnwIPKg2R4GNLu
UbG+cXZ2dVx9oRvJdf0IX8BRG4qMbIZ9mRpu9vYCu5cF5h6d1V3n6EFGANhbcft8
HVTknvI4lBgenxatj7mWpaRM9l695tHNf565w3V8F1Wxb+I2lMFo3QccXf1rq8Ew
lrYs+lL8Da04Uc+oGvB9AN/FILuJkyLGgcqVNNkwZ9j8RHNb4lIeVk8ARFjURR+7
FbuMR1JUVL3vWfWw7glgaNraHg4zmixjH67Oe99OTe4KFuFfsN5yKI+l9FgSLgPY
XE74rDsf13hoAKv0Pm+Lmub5Ze8wn4Z4uKfjrq+d+36Zcr7GPvqnpH3Y5Py/rLut
RKMMtvCLHcPZarQPDYDNsuTDtBeDFvc4iY5QDB6tc9x/VIR3KGJnfVP9DfAA3lKK
YQsv22G8ksE5MD32JVwNN8BIC/dX5hcFqe1eb7SXFpmPYXLqvotwvk20ZOYoAU+a
WAH94ET5zPN6qA81WNwQuIoEujnd+g6O1+eq0tqrug77msBjuImo3Tboktreu+RB
sy22EG/NvGFpc+Ecs1MZU1+NMRC9P5GF9eIOJP+HgXKK5I69dnIhxfQxM4SR8mF+
4cXbsel2Oi8oSTVwk1ccmyQ8oxryplhvjgxEqsQ0h/1uLwJIPfZnJSTuDX/48kI1
+P5upmsvrnquCotxkoFQ83v79+3O9YIfvwr3ubZOUb34hwuA2jPvCO4Pj/m0DBXW
MSYuQ3lkc9VamdddMagRctfQXr7XlNFvpsSIikyZSfgTOL9F2FCYXrbJ7PoN+74j
H8qgSmt0vDu9YEfs1e2TIQz/QH39W5IHOrfRQQhWyK7q4PMChA29Ga23FPJoxoEV
XPKM7/I0CI8cljdemIafru8u36vRY1YSgEMYrPLiTXlsh7lJ5L+JNFG4VcBRzvk7
pxykJUhckawVvcp6IS05tW0iYPO7W1X52Gb6gInQ5shKPzuErOjyu2I2fsaBmkmO
WXkjlhZM3DckY5YD1/tBdvDtKE1TXc7CE6Dk6oEZret256Yjz9b6xl3dyN92BmKC
+VhB+wJCs+b3E3uOiKsYfv6DLcOf369rVgW3ppIu5ONLkJ05Gm39YpxJ+T+Ilbzl
z8AU5GP0uE4ZNEUrFNn3HvZP4FWk2jUHqDxTH1eUA5im6guUDb+EwXk2tCvHN6zq
8nc2a10rwX5IHvdX5fv7hl+Myfbi5YxT7MgmjAkFJblJ+AyKuTekT+iwHuaKktzj
h/rjfP/GW2+I1poHx/EZctOIAnPr+cBSOm9ghk0JmqOA+Ss0kjsf4Gzy/voYspMY
ACQ5AAjfJVOK6lrvekh7+0YLfSAb9BodoUyOo2gXto7R/mOpC+1zgixcAoN1dzC6
Wo4HwZ+d5Fea6A2WE5Xmyrfa1yz4401uNWWUHYRVzM1Qe/a7419ovDpRfl1K1qWG
MUz/mbZr6Mx/8cAsykdh++73KEjMeOYERgMBevrszL1dsD50FTAnz5OW8guf8wgR
BxJPoQQm3zgsyAzK+zJh6lH/p5xoSrtYKKGF2HAdkLbYq/KrCrX4EZefjFONqqw5
H9k1TJE0RxWkVfcPMlBDqKqY5FzS8eOBvnSZiTe8v63mJF4s8nDJ3dHp6inFynVc
vLqnecmpGhsqOukAexuSvLIvSoSvyQv2IUK0iAVaaTjbAGxklshY/dnOUrLZslAV
HlnMyHXi4DmNbVmNC6Y9TPr3w8Jo5f/doH9HtBRTh5qv+haKDFI+AZV/Icgagctb
wrvMACk2QJ3Lfo392x92VYtbaruk7NHmnY8WcyPzF4ZB7x29rXjUpz1rYCEQyf24
EwKk+6PLJ65uQDSGYjTUfPotpMK9phxQeIzib3CM5aIcZ9fC9NuVvgqmXsxabnA3
0fLH3ZOGWK2piAwSYwYdtl+mSZH+OWsmrxgXY6Z+NDmDcc4DDGts8FZaBhQHJ6Lj
aWKvFFdjoqn7e+sPQYuY/n72nlBrd2QrBrToUn1/CeCJXIZ1FbrIPeWP/Sz54CS9
qUantP9RuMAG0QQAmWGiQyTn/kYWINEFMajjz6WeKZvp4Xo49gnQpLIvC1n1aFjJ
81pANncZ0jN4vhGypuEETfUkE4nLFAK7zOcFCOalDsR+Ecc0ISP8Z3u54rR+M3bw
0sK9obaMqoBNjsaEhHBfMOOsw0AmIhtO0f9Ea2Zy3Tk3+UdmDFAqmpxIACMsITKa
hsvfOklTih6KA5vxBb4PKiHZaVHhYm45YAd2gPbYynRs+0auqeqy78S+9t7e0YDc
+7OD/x91sdT5uv45eFxYbbeScURNQP+xmL5+Qzb54q86KFBPQV+fVFEK5ss5QGg/
W14Qpw2wAESWBSBAEBXeFfk0sY9aVSHyTnk+un9A+AYExRTLm8pxI5uPFMykKMo9
6yJ0R4J6G26mYemEkqgcwm8OWHZHKBIfE4vqPEcxU7DKSNw/1G1yJ9zue5WfWkb/
b1rNRs127q2vXkOmKb4XQC8zpbiAUf13wnyI2Gqlf61TdPd9qtpXpxa9uKRxMAqE
cnx/gNN7BjZ5PL39dSzG/aHQK3cZ1ciD129YXXsdCY/BK1IgIj2PtByUkwlLJGLD
pAf76FGlKWzeAr5T7j2W6HHOF2lVdeuV6gMk7nWOnR4YC3DSE4v3RpCR4iT1x6dh
ScMbyjTD0MhWgRU4/QOcqOmK1XLOmef3VLiARlICTCpVibkNhWvYhEIFP+ndlMGz
W7nJoH3gbblDZkWcdBu3TzoceabSpwejzOSCbsS3LzRVVTNUYEgXociXk54tZEnX
KHMKvT1uVuihhQX8ieq+Pgr1a2cP9RiiBRpOM9n+GPRHVUeX9yI4cGyYjnPXpp+e
S1xcJLAS3azSnuRQER0G+YHUlyCwHH4gEZn9GzS/Z8PP7FKlHZUmCBYdcnmoYSO7
5apHphd1aMx02Ot8sGVEiUwynljheqyIEosd9T15ulkeKpNG0HFocYJAhgj8xL81
Sp9wak4il1f9DhoNSaHH19ILjC4QmMrt1XQq+11w7fiufxdQ1v/zTpYBOg3w/2uC
d5P5CkXNw2Z07kffZImsamg7bvXqFG3RD5IH1Z/dKg1bEhmbzqY1RETV71xPP3Lc
PMFBRK+U7eXPziJrZsZrXk4CthFIE0k3rHqosyah2a0Ono3Ez3pnrkcCa7a8vTQF
SAJhihGYe5KfdOCv/VNQiNaNcFIIARfO02oFYD6DW6ztq10HmN4AjalVXxcs+Kfc
MqbEbe3BdrfjcKygOa7xCBRX9eEnu9SFIc9zQ/qoB2hTS7NFVBdmKnxmLCrYch77
hM0MBPlt8PwE3ooBJbmMzXwO2GxtzHCk8vEf/vpBlCOWso8pkxUmim/gANMtrHb8
5eEzqeSaNR+yymthAmwR075k8iIPK2MVrYTL4sso0EdQlc2+NuKPpyFT2bDMInqD
VwMUVaU+7R7BLeeuDnazGHOCtmP5Wp93Xpsv5LWzYoAswCI1WMCwtSrGaadyPHqO
p3J0BVnqzXv3Mdg384MecORY1SFvXQwXOQVYP2BrWnaSi5fc2YitqXPYPQxIJtoH
5gFpLHYoxwQ1bdN46XDs8Z2fM7QxoePv1v7UUIgVy4IcY8pizLW9Nk4e7F+DqRqs
mAYoYpm18w5mFw/9gsGF/swVMv2k6HrJmpmsnOuWIAYo84FxbWcFxxBGd2MZBeSM
o1kpn6hzbJwcJMRcg+YOUXAAeemXXsJkfawhFpewZVNuIedARvfat1PmvydTtGyR
AQUrNnA7egXb02vZ6zr7qvtJDZrOG07HzE7W/IMx4MgTPxhvDzImWbay/0U7Seru
Sf6e68mPpfs1fzY30tvpLLzPo6paplIqsLw7CsonEx2pEdzvgtVUm/qfnQz38jLr
k3rPGpvNw+DDjQe9fh4TlKUhnwz+zRZUIsCHLYF3OOI0db4TamRu/dAdNLfxxj9p
j3U58p93qDvKo5Fuef6DHNlgFCVQW24+zB74jqJdBHEjyHnaF20GB/MGefUatlo+
HmPsa1LoEqRJqXpXR0HC51Pjc41TS7sZBsrJN3KzDjVxZegTsb/mc1GocEAaVXQ8
a1t8nkPtuKk+Mk12mfbrwVu9IspLKcOez0ku4geAJzyGc0cJDUaMWKxyvLNueu9t
SUAw+vrOSCmxT3qr2nbx9+gCysqxlxIjTLIuYQJR41zOG3Y9QtaHEdBDhBdbiPNs
3suAXtV84zosIj9OJiJMleC2OzPtjIOgjDEclVkO51NSSKj1gJ34KSBJHU1hTGST
TKJwuZDC5+IL6S4SnnTClGYSSMmmZsQBpZ6LNonMBpqqamsOHCF2Ph+NPrFedGVi
cs9qJlB+AsmDFUjUYHpaiAdU0ilOLJHYZ3LvEH4HsHgzzod0+oqN5s6hbOpcD/Z9
xu2XKc5/WkMzOIo1Ud2omvnYOSqcFpv5OpBUogBU3PYWG82BWTxW42Tubr1yyhGq
lbtXRqym+d/aIITYooLfd5a8Hx1UVKWZqceJI2n0II9N+6knQ9q0EKS5ukyJby33
tLRa+B7TEKGR7Xqcu7/+OclSiUhTEM5MXPo7kewZ0uNUfm834RPBiCl4r3GNG7XF
WDWo+6HvKcgK/YZjL/b0iSGM0TPa/gvQPAQGoBnJmpPHoCqTiUDNSYsDgPr2/Sl4
3nSy3zj2lwXvDXDqNWXEtRcNo+sdxHUy2Tk7YRXyA8BKY/s8F71w6KCgRzkSiLwi
R4SPTENAmL3hR4A0IjOMYCza4HYiiqCEbRVc9TBnOlpCKmiv4AzZ8sidmdCUsDik
g0P/X55hVD1PBlAVXjWwHxEdr7OLYM33/eVWa8ZNFG4+hBza7VLOCqATf+Edu0+G
C/ok2+dWR+ytfrg2k/YA/Br6P5M25Z2VRC5BQacftcXh7Coyjs/IEz78N5civHak
xdGLzDUWA1OrWUj+o/OtocFEWKskcM+xsdJhwK2Qym4eJc5jvdiwvG7RXv+YRcJf
uQWl+eGGiEA4hj5yBTk+8K012/IQUITKbVATvIK5WeukwgpAGoA+hg5J2UXEVKU0
clQ1Qu5Kw1Gpr/8jGxYbYHyXi3Y6fE0P85kcXo94/z2qZBNcydmQb4UNSX5cIBY/
MReUOekDSaj1apAWvMd1fAVKuFnQdzbyVjYTvU7IVblF9IIJopFhwdsmCX5TIEIw
d7BxdVXzrDLucikTBylDiiMzFpBVgCBW9BWzS3I5Z3Z05ZgwDPA899gI5ps43qFz
AE9w0TqmyCMp7b3xHKBdmvx+oG5eNgvhvAV45EofY9Bt+jZ6NMjYOntZs40whk+e
LW4zTDJceyH7ci8j51LY/cLt9yslGYPcNvq84BFa4ajpeb8pqkJVb4MXhYsEge3+
cef0n29Va+few56GeFRBIfT1HJ+GyBt6XgrpXmRDWpLqOpdaRHXI0sNRf+7BkKtL
EsGbSSKfZOBOe5NeJ7i2tuHlyC7EQBolRbrBJmPwf+oC6i+n8JGQrOEzfL1y6Xvn
78pQMiHauWGrZtE1in8yZpRrOfI0ILeGuL/MEnCh3Uct9BT00N1vU+O6QJDC8pPZ
+Hd77Q/O5Idz+2aW+12cWz7FZxNhR/SuGbZLR/Em7qz/io5Hy/bUbbjgUGkxTEIx
lOITMLryWbrkipA3CcR9MYwE4IOsLmpqkNd7LgiJ5U0/nOqXxZ65D0Q9Bzk2CeSI
90V8aPVZXVf1J5jkxk28qz1rPad7sNaZUD0WlxjQiz4CLRwCNUa8iHITBx4vvZn/
FzoVJMh4229g45O3vKlXHzwLPM3gVJi1bFWrT8dD1clJWDw7oELxKFO5t4HQuy/2
7nD8N0wqiUncv3dG83GHBZfIIYGkG+m4vd5YwDDBdaxmDUarcGMiQ784pNeH/B5H
6Gy4RKI6b8JZesx39u2fvfsRatJ1Xd1PRg/jPKafKu6m0mH48Q7LPXSxuGi0/wac
0+5vcgiGjQLj/iPQZlt14tiRjTLswl28b0Ih/Bk4BEHdBs/kaWt0o2ize0xCwtSJ
62/8zGaQZn7cqnOY9OKbekd9Q4PELxnMgAiwK7c9PpXi5Fpkc4ygsehi2lk2hOZs
ktfl+DtEBSXkygqU8btCOFc5CzvNmXbwN7EXRTsOsuRqjAyvO9wboTQKk4j8PoPO
wGVYmsca3Z6/AMnT/yNsFxp86MhuhILwGvndxkfuiUUTkTjf5q4zJv4Dj5rsuCMa
k+SSO8P3S1M871ebluvLsMcMIsyL9+Bu1+vy8wBUR3XsSe6lSKrrko6Ow8Qsa52M
prafq/Brti8wWerJfsXEaqFkcQm3MKEJ114mRajqZrT1L0+hFhw0nAuxPbl2TTVr
YVmnLTQMnU8xkb31RT227neCHv3bYMVoiL8TsyxfIWtF8WmCckEBtg1TGf5hwEY2
LiAvbSvmJ6ULoBu/OYn8LZPUtMnymtfdYozWO3LBsMMHWHAd3zH5R9oO2mTKxDNQ
rf65RZ4EA8afiOvGpSz6BLSHK/N888iiXZiMx7SF3jeParcL5wYTnPL8BfQbio0v
RPD3UyBgpdkYf7pWa71BCGCHf95fL+/3OCAIIX0DU+8izdFIYwbWYP1Wi1wNTlKq
40ICr/naDM9W8TqNBTQu7iuPHwmuJNBTiQvP4sGKcYnnDW7YUISKOoxpcA05rcRo
U0F32RA0tkI4noaKU0mILtveLxWhKaRWsoelrhNFPc1HZWCHQDjZ4FkIiwShGANO
luUtr9WHFzDvt4Fmu6TSGKdm2OiSVH+po8/wCQiNn4/TDqxlfDKllNSntRjGnzIk
GV3YQwo5Rrp7MTcLtazIqMTBJn6wXmqyDTjIeEa3imyJIVGx4XTd+/0uOzKxFAxV
A/TOixBt5HslcTl8eZ+uMTj2XbWuUvojJ3yNSe63mYuD0HDjAxPPpvjuGihleNVf
JNkgzi9lAmJ6ZVKQxJZt9QRbNVyTKa0H68mNxbBiPkA/cnutTf4p/HIofj6EZ38L
zAOfK4G+cmeRZQdxgVAlbj/tO773MxX/htzGRVqOJAmf7tKgeYShM8CnRwNBnJIt
OZdB0V3vsARl/fx63IwAvGv05/xB5VUq9bb77j6W/zVwetPyFIwn42fPQJyNRUuV
+16hiaqo3AkHXuYuapdKN65Zthf88RG6hwpoPlJKdftaIHWsFICXywakRLlnmtIF
W8/IRNfSPlIKUDt5WXxHdkJ+C1i+CP36RS4RQPRr+z8e8SBSd5FzePWAbL6+NV27
LsQcac49LNvk4My60qpfR2mifyoS2gB/oKU9MmeMVq2ZCU5uzc4a3MQQ0U8rvl40
n+OlnpfUPXqkwKoz0PPUt6wih0p7y71CoBcV2TfEy4CMr1xsqBtL7+VBML98wog0
C8SNQTeEQEpXZgiIKVkICzYbqkzvR/fGZ5nVtN5BOd5wsrCBTqApl/m0VXyaNZMF
FvEsQ8NndcFwkXF8v6BcDkq1mrhDQRx79fuymkcEeyZPyng9D7LoN7GVlTJVkhXx
PD9h0Q0+PQehvINAxbi1+USGV4AbdNKlWd7tVFFMO3NINRvAvaVT4Su2pWu9BPru
BTz12NAcwX+qbn/c/XPSl7OlfVHcoV+zR1bGs+kC8Bfc3X+bPhfJGYk7OiM0jDW7
87JJQI/ntORWKEZgN1nFlY8p1Lm/Alj9q4dYA9z4H7wDbV1XwCrniLLRg/5T/CfV
V8q5zV2vPO69J26vcVUScLWrDzzivS48V0Thu+yYZXELqNrWpbGhAywnEZZt3foD
g0UrLfRUkhDOdlit12O6c+h/rtBAeTw5foLtJDt7l9tYavo5g0V4EkGLuHzS86ZH
UNeiunoaM1fvy8yJbGj9UWRMvvGGWyJmy+wleomT5f4y7OoT2tjfbWvjBy3xqstD
4b0GyVGUmQ6R9gVboALteBLpXzPaXCSvLGXLWHnhbHAA1sUqV7gC76gu19OL+erh
rjPtIV+L0t7TzVB/nvzPKqn6EtHgy1XA9a8pexfHbamEtT4nldVmiywGOky+5E9y
a37g2Ci9PuC5Z2Tl/jfIpXUOIMiBvvkmBTOcwamxHqvGn+6cPpya0j1tOplPcfGj
OfFx7EoAUM7c7BeJ0879ayHdVX+qKRWyjyy/pOxWSvMUw6fI8dmmo7rgiUqfvBZb
eeSI8DgNwHtFst0kcMNlNU+/DgKnIvC51FpS7q4N9nCWVqgrwobMYX+3dCEoITa0
fDeExUIRHzyLxRqZbjMuHcDRk4OGEx4Vp9fWdejXXnzJHFo3zVegCQA67OlYL1s6
zc9pb0f3hWMJhDDFAfVmJHGByFzRhrPh9PrtVTFXdmXAh9y1pmszwruq2dlCxyuB
gzqaDF/UNN3ARWSQd++lSlFV4XrU8LmTwY97aw33sgvAcGJNhXImxdr/vwU1Qp1k
ufV5a3zs6IbTAsvGIJTdFZKvDOyuWzbaibVY6Z57qwoFwXmjuVxMZAr/JHj9LNAG
baCHk/1Z7OzvHZVoesCf9go497BnONGKE9+S0UCHVoCA+XI65lT9BWNpxHZ7Vnn6
w/79v+2p5qvbSCco8ikGaDtXsI7uxOtftF8CfQ/+shpp/zZdeEmnl24VFWS5EEVM
GWThBqgxc0XC1Iw0yw/l+YBmKuR1XEJhz88IzNVSgsPAGrAJ+dvmrWyFvfq3rC4l
0r7/3JSjE+cIa1PW02m5Ossd2UhRE+VeNIBF9xMCGS8vM+DzUROve1Cqtx0smVyx
9/6Uvb8sbZD14LO2rfjwewZ9g1/ClGAWwKOs3kK4ReDZatJkYoCquBtIkJoBcwPf
QSgsOqSFUtMJ74Abza0O17XXHPVSYOtLdO8Dnav/DwCNzrsjyevlgJI11SxCA7GP
uAUxQ2qtIAcCHVluSONpGoi5PhVfx9q/1xxvlMtEvNHuCllTvt9v4VHhB2vYqVX2
nldqrToxU605Z5XRk9fW+mzc1d+Hu4CnmI0my5qGcP9uj8NJyhVodOlw+QHZsOgY
qBRfacTtnxn3ErsgyveJye/VRIjmYy+Bym3lUx2FZ2cq4hLYHsFqi2k9yMlrmrUr
6UCjWYoHHERhWaLmTlYF5Jl/ZH6ApKcBZFreGsH9UMB6H/zJ96aNFe86IuqZMYQr
LE0i3rrW6Gz2xBDaNPfUM8sNr1dlG4FofNMN6mjy+9VG7mUiXPN2xwltQhPdU/7U
eMrZ35zdcKlJHrbuY6bygUg61Mj6F7+/06phQrNC2sLUyzRB+FQHhc6QSYQ2xPDb
uymJ2oBMhHRFGBnSIQxIBxdXZ2MNN1iL3i6itYMtcTfkc8lsjzESRyHq4rGudNZ+
k12VBC6dHweRyGI+gRAUrp/la8IkUXU2sCeUJ6gPLyO1ewACJjuqFI06En0AEOG+
kwzgk42kWWm3f5h8q9k6d5V21X9gz7pLHy1OjhD9cYuaCZdsXqMLaacZgzdkbBBU
xDmImyJBVS0IHZTzq1Sj6rnbDsJZzLvH5YehRWs0qeaShy6c822d5iFCdFA7+SAN
VQE2HpBSFnU2MkkKb2uRC4UQe/mK1tv0bgR5X2wi+4Mi4xXsYS90aF9b0xbVo8UT
gBvYLZSGm6Bl5ScRz++AQR7mynMHgrS6FTSxqDGP+MkE1BkWa6Kz97wAgGX8b1ko
hvvtPbJaoqhClyf+ILAKcDFV+hPbUIIdLnajusuMsPFXSlGWZhExa2UC6le89ph5
rMv4fX50NC3No3hXTeDun0FBuavxIWk6KRu0f3tBZfOiPnkC3B4m4OUMJUYtADZF
dhsy9S7zATIRW/f2TYMIu1+hjWFLaeL15oSWRp4Da+uO4Af19WZ7G4mzovWdLZdR
UpwLIpCGi6hfJ/d9B6Gu6H07JWSxByUazYrA90/Owdzt5XNLJ0DPgLGIdRb2BK7w
jB0W8yyE+7PSyXFREoMsqCnfvDFM6+lAH9T/QZuSTVHskQqUQEahVHe4CnTzq4Gi
FGWB62pHAROzo+M/q37MRY2VGAEu34Rra3DyrOPJ37iunS/imbyk0LN6W5tNC42z
NZheGi7KGV18QQwa2guPceRQDzjldShwBlLG9KMzmeh0Cr0ifzCEiM6UG2P0EmEF
59NCMPBGUZ6GU4pFkEo54D77OIetB/h/qyhjkcqeM7EXEN8MhVrKyLnIPANNIOJB
rg8WkrdasgoKgY+S0gmmbvuVMCm90gDqIc/LqkOy23xUianqkxgQRwPrTpfpp4Oc
69VNuoXRN0sKdUOJZ0yfolN+8wRGRXfUxTKft2IwAhMk1xAH1AB18IuA5xKhvavx
zFyDoG7o6YMVF7AoT7kbuUPHRh9c0S3T0sPst1DUIC73CSTtAAvqSgc/8oLYJNvy
5wmTawdP6YSuC9LeUgXTUyg9mDJsui5a+QoqRQost1EvhA93sNH3zm9y2F3vDsJ3
2yunE0toPv3DaLezdN19/lSaHPmBQ0DwBZvvanie4u5hCHPbE5Pyd8pbyXzI9Fmy
/3IhBXd2Ui90O8vjEXsEA06PA+KWYT8+WAco8NepS4kzhu7AzzGTO0dCAemxEhYQ
ORhkCJi8s2IcLMACVxXMfyK5SNchID1bs+028W0IghJsbilXr4NlxzSMOuYXx6lf
UCOLRLxRgLEkQQqhKsyafHB486jLgI8VTocz2s78a41wFXfpTiq4QNNznhlgdHMe
JhddZWUybuBUXHzcKeJg7AxI+Gq2I8Td63CLAJBgNd9JRkaWl9g8bygVTJSOnVC4
dXSkrVkFEFjo36hy96DVnSqUFzYqnOgFI34yxS4HMO3UYfAJjOTqpnkZUVCycpf0
5Vi7chnbMnfJfgCproNCl9o014sAcNXSSO9VpFRxLPJdiOM9UQ2guVwLgXGujPq4
EOHs6iYkkCIFZgmYLDILTSMpAQnv7ivqjOeBtRwJCEHSHdKLM8NbNCawtxpfVCB4
mHe8EIZ2Srqva2mkgBowzL/j74XAekX0FkoKWgMBJtPfJ9EUnb4/65gqro8fhKxV
vZbvEP7KgPx2ya+aR/s9iol2aP9mdalpEGLypq5LUMpbA0CmBgP71LMuvIsZduCH
ks+Kvr4qBTAAoCPyYkHT4iyQg/7B9Q8+4Ik1dipruGf0AQDX7eeqaT7pnnUk1bOB
ScxhCuO7ugHeepR2W41M3rvQh9cWSYIXMZ1CW/QcpBiwrFBtKwANhFW0pgqBl25b
wA0z4DEjatq8X+WMBNI5Mbjtm/m10ebeItVB3OeRd9fMPpwQGEmjo/iy58NyAIMc
wyEKqfClKaTdi3DW/981oLJv0Pxm5qOLVtlSTZ8hIB3vCqJq12RMakGSMxDpEH49
XHdMEoKKRCJqdjLUbGiOICCgSKk4IcXHo9oBWDJFVKwyBug3CcVPQCXwRBFzK0DC
4fT5mkmv8RynHSVr0P9rQPicnJCPUB8UyjG1viFeYhCyVPXA2ofA1G60L4PXNH9v
acFyRb/tlAbRLsPyOcYHI0Xdgs0E5f8k5W6s2WYHGRZlxiolXz7fyccypgJqBjO0
UsV0NDEQOeUsgLofqvYW7CdpVEGg55IzBWn1EW6m6qPEAxx64bIsOxTTE1oPQ9Dq
sR+rVeo01Dgrk+kTG7POtDnt1+03tesJRx1stU6ElMgeZRb44pKf86eYPzbL5dmk
WRvIokVZygr1vssc/xRuGDDPhq06LsBBtFAJzuKfbLHRW8mmLYEj9txw2YayI6Kp
0lYTmRjuyEk72JkDz2X+eOzS52BwPSy7EOvZLcceDqVvoQdfqea5PcRyma+rTKqR
sx2yDRB+pw07ypd0N6G46ZWSXUUsmCum4ujhnwKB8/v6MCUtqyaKOEszel+jTllF
Dthbqc8Yd5awgs++laxFDzzbm8Sr3W6tYP+T+QfrfVE5tweR1XKpbdhbeFiodBsA
U+Yxe8+cZ6nLJ2rkJBPSsBz1jBk4f/78Pf7vjJcxI6efA4PQT1HFUH++WLFkvNXR
fZ4vNwC9nyx+sPKuulkg9bKRl46WjVn2+9f6sxlbCwzfTSG/RuHll5rte+1fRMzU
MST5Lk2G2EQy2syycbmxN8DkM94m1v+buEvUNGUfvZB3mJX9qlA6B4TEywwx0MmC
EBHdB8aZ+hlebfVs67zkrSKsK7KCv4ZiR8Ry0okp++2D/skl/O2SfuzlQyIFlp8T
xjlK0SEdaaFyNhw8oRP7SniAEMby8ZJKSJV2xOXUyZ3eBldBruGEORSeXnuJ/ZrD
mTU0y1mmMMTeIKkz7gNM6PMdTNZMF00AovBi1nqNCdiEJFi+72ecGt1XhHKsMuaA
Op4gbk9sffR22c5sqmktyHD2tnBiHhkDwSrsJ26QO5c1oiNGwpEXQEwHPQwFZQto
GQTaBzwHhDr8SycHvnJ+JPIWq3VrQW8eCw6dW7SOfL5NefIRiPVYx3y4w1NzCpT7
Zmh8EoC3+UXpQzMNM/QRKV2FQ2/fpeVzXBBGJYQhYrfSauIr3sZZs4H70kKMEA6i
kp9qY0XR0+xq/3DR4y9Z95hQq9hTRD0nVXrrsO0kLqw7Xm35lvGaYbsGWDsfZ2/P
nQNmZUqirlQhFlBi27BIdanqEp+qjKGW5EGTwbq+0Vcmd89uxErcQw2tWQ23SbBq
6rqGeRAMqs33yHvInMu+A9q1uJJAl+81wr4DgIUO/bKQwW+8fmEfYkA5ykndy9hJ
J2ytHBo66/iiKyh9QDSLLFhgUJZ3NvTOsOFJmsxf4hSOxF09wcUB7YbGWfvkG4gV
1i3LAmxJlJDeO83Rwll1eEaVMyHE1KDLq+izN2jPPtJAImV6UHvoHg3n7SQX7Zjt
igPYrDx0nnZgJrLq2aNi8lEXaYCoDX6zxkcjWG3sjrZvL848OM78WtVQJbm7lMYQ
3rkpg2E2W1BLLpefMZjI28n65s8IjRuz+9SCeWeMaNHvF9gbjaDgcffbmQ5dMaf3
iw6OkoUJNsqoUC+v3cSr9pSu2SEZXqOsxIMcX6J8zFQSe2bllwlv9WjsqqIIgTwi
Kbbwm7QH/6TnSwazEFsocn278O7VAXG4165KAVINxeKszy7EPt6mP5sJTWlngsFK
3Aky6W/gou/Zfy0kd5CC3u2DCMVUNGojVsQzJDcSCOK62dtnWIsir8hypH7m1Nqu
43thsL5helhAvT6gU3hlz+vfZh7U9M6Ssa6UXGD7NVNi+FV7ux160MFSXNJaBzlO
bCA4Hrvx2WzlHqYV0Xh2qd3imcRE3lupNpCV3YyzFwyQxCK12n9u4S300EmQCJwj
m+0lLmhiXHyH4IEJaBigH3r1oGqVk74TSxalB7rs2y8oBksyNCvWgBB08DlECkKC
p9oDfnFBm3xNIGTtdB1uD5jwgPQFw5cpYGTz4OJOPilPFbhwHCj+e01sRPraH/+2
RVodLmFbvN8MEU4tsjwFdlYQppoA4kzoBln4/NS5aoTkHW6/Ahk93rk1bZmghIK+
xujJi3DyiVIgFYpdq9fwnub3G/B9L5Wd7CMqkG8e8Y+HAv/nyGmfKnqsbDtU2FOK
NuU6TQ2bJBH5uECabe+fwUxOgmoUc8MBM5y9th+416CzGfRXXUKsCR2Pifach+qp
QcGigIzeX9t2MAsHOcStnc2mRZB2zHZ8R7en12nm0QU49X7W6NNfMQcKfe31fdV5
loZ4YD2rhvhhTFD3pGcy6RCju8cmRoMPzpcUcTFHqgjBc//lwtk1yCaUidDNVRNS
FSalhy/AABqYcFZrVtApuA1Tj1G+6CthrwbEiKMe/R9wsqJvoprqTbt1gx90uWhG
4Rf4DR7JGRh3/jjBWAEXB3CpTovhtgomGVhOGQ8130THCxtBaKglvt/tkJt9eWs+
2dmjzs74WlnPH/G0fXZ5s/VMDfHFyEBEegQKfhX49xvSMVqjBLH4kc/QdTNoLKsS
B8cKhfNTht4T/Y7haWL+7gpM6qnKuAFymJRz/Hm3P7moMIUiDRXjCDsyB+9Orza5
DxfcfcTol65FaCxuKH0jQyL0qlBrpK2b1/jCjGj2ymzd4A22MJISoB8WU2K/y906
TyirO0Dc6G7/1Jwd7jPfv+gw0uqiG04stt9y0vGVIM2tfA9xpSUym5mVKqJDI4Q6
R/XaKhAmho/BzQwcWVuKel3+HmURNSjIkNKoNZyK2VPwBtTCaxz5QUPB4Bs3wQY6
NGHVUODt//UE6u/ViSWfeuUCszde2Fk8pvR9yUbsiHTruEm6dYPxG5v7L208MP2l
zWqYHv1WqDFCUwqX3YPkSHP+5bA3YeSuLyJxkLyBfXefYmw8gAkEq1J20wdhxvNJ
dftfVsfDtiFx98nN3wWdLg0VU2sOJ5jcYOtlsgJ7NWN2ygih413xzalA5xRkdqrX
4sd+OWihuFlcPK9BwJx4opF7bg7Yrl+wKPKQq430+BBo58aYhjZDTNmc8OqzRd8K
8rg6m8z/IuW7KPe8kUdqXII7NvOdBmbbFcbQRM9ACAOuEPiCWzfkAVDW/GB0oyWk
rHgfulhz2kSykxwLJ+ol3+qtDbTilapS0LtjvEz6uwq1bGXTqWzZctnY6aLTtUT3
yrWhoDWz3ziayrJvDywOTIxjtjhBDMDJ5/CyZbEyFYe5xCeaRskbg3DNWpKm8dJA
nEQhjPC+7Q9IBDYo8yn8CflSPKbG9NwfmDE1JhraV0+4n+swy+hVaGIKY7UJD/Sv
+H6V9fYmnmwbpu1ushnzh11W4VMVTzzOa+jkEeSI0yGzGaUZ8gLmR/5q9HOXzV9n
fo+hsti4mo7D8uGoKaVNPNpAFHGpIU6ixeveKW4D6Ud2Dw9AGwidUawPRQhrMU4d
mum1psWkDSUlcQd9UB7KQfYkVIMhe9fGS/L+Niqfco6p2j/U8/jYBq/BRcq6kmw1
3zg7UbQnM8MEldY7MU7wfkwC1QXhKEhSp2BoO6kFqOg0hQxn+FPTqQMI00pnvciQ
GNcpN7Mb4ADcBhxkspALvpB+GGr9IeTWE3vq7/7kSy2Do965oScMNyOOMRItI+i2
TlbR+hsSexNjw7VEwFC+wSlSAzSvzFQlFF1lcHGlzzUOV4lyt37I9y+SkNSsTY1i
lLSc/UVHhldaMJ0qMosej58Bo9U0ySlxU3UwCe17Fqir/DVY9kqvphVNr1dZhi4i
qM49nSsO5VzQ7IdwLFy1orPs/SQ6tuUyW6Rn1YBIlR60LmVnKEp9bGSnHQfVCQEt
R0p4ypMjTjtwr6GzapEyhtY09JT920td/3/ZViLxZRxSaI7rFrdRS/zt4W5o9v5j
wNAQZxP443jUoCMIz7HtuIicFo1tvT9q+ZcpmGhSTS3ogYacZddLXrsvqJHYjvu6
AzLFcx01zgw6telmrscCdyYFeyR9gjZQKtKbxJ118a2VbtBVact27yg7soRavMRm
p6JB38xcelp1nkKyjDDCd3FG7Bx09p37QzmwgyZyy3ojhjw5BqWb42ACw2nqb9gK
PrLDFIO/fXTVb4rOLoj57K0HMrZwhQPc63fwqr3s9XxRqBm9HJH5NFarRo6BUG8R
7n+fladFxJ0fXJ9Fw2qNMppy51YGYGEZC2uzcRtOTKOBxL15PE3Zl6FSEdoPXBng
Eg7Xdvoc+z5RqhrxECkl0druhE1hlOC3GyowhB+O8Ze8oih955yqHarmKGM5W2nu
VVXGXN3EeTD5fkCekneZdMnTzqdbD4/azVHaxLbdXMj7qHuD1vox+qy0U4re1aD3
2vOqdOJXBr3aNYifGc8CM4O9u5EVl6Je9saM6DpATdIPWQaFFN7MAVfwTIssqOCD
ktdmyADF6cyE26iZnTCZav4ngWstp66jVX/8M58q98bc2IUvw/OLctbU6pvOvVif
PA8z5yIzV27W1VQ5hw9BPEB5NTgY51yS//qW0xnVKBIlUkG5WPzueeENWhHyRMCf
l8AySzTKPy8vk5tksftbso4t/68oCEgxn8QfJ63+rVC32V6DuJfobPxm1b37V1jp
2xlcyHdegYK/Y9X0F3Srp4psN1vJeqvMpASSfIjmsfKLDJM8VUAhfC/9rx/u4NpW
DXtu3Qc4f/18NYjCz5U6mZR+RdWxrkW+HsIf+hlgiSH1P479yEXMi75ry0sTmvhf
sb4hJZiF/mt74UsdDsqrYqNTuI0kWOcdvSZes1TcANSBRjAKFX3t9T52C8QXk7po
bVCSEsC1EYXqOn3HzIoS5YVJFhz9F15Kz9MWEmpAN4rfjqysjjFdOEd/N82QBAzf
eD41Mpip9il+UzegKt3Ay+SAzjPFt7NkjqHZJQuJjeKeHuWXMMkSjw5stmO3LLlV
QBQ53O0Aw+pKbOK8DAQqPMHI6K+3E6GC7kWX7JcRxFcFx/MgKRJgEdmVgjnjjF47
jQ/Wws+GTzTvcvlFyaBIjk02nO6khZlfZjNrV3GO+6VIrA5TFXF107wrl5ma6B5r
KdmGiNX+3qq45uMtJ2SsA8PJKNIHubKCjbMN49Tyyn7Fg3z8oXswMSIiYbpF4lIF
XQiyVyKb8d6cZ9hjzcWW2WP/i+6PbNxgFxQ8p60hIHq5FUnV2AI/nFFS0SDJtpIZ
dlF4hwAqYgrUMPBoevxNriGzqx0Gp0lgWcjJ+cykPnQCzvWWCyAm/3NrPsQlOU1s
k5X6j4OnCSIRskcmQIFBCTvfZXDh98i0D/06kyloKlnMtDQ4gvgslDksF70j0Oub
4u+SuWA3/5QdniBfxMIOS7ko7PdNvc2leRaNmWweaSSivV2ETcqsOb6k0mGQh/eg
t7qBm3Qs6U1Od5P0GSloSr36QKlLktNCChb2rFdLq+E+dkQJBsfS+FDKy9y3cQ8f
/QgA80qVFqBVlNHXpfAvr2/PG8IQhdly65XJf0jvc1ogl36lvvfS4kfjqqPXoJce
5sqEDnXXo9ft/nWuRKDTJ+jB9yjRdLr0i5KZmDrma8x1LKF9hM0qFj5VaCCKcQ3l
20q474DWYFltREhFutbpB2mQ8irle0lvVCA6gbMBgcEK5jzBD3MSGGXOq+zh8BdW
52IpSkOcWUicfjjhTQXmw1IBZRuHlJo/gevo/fe8TIeW2HfrJPPoI+Gkmk26ZWl6
eS7rHtL9kGQ7CqgGWgN0wCCoZXETc381KE5RwVR3Czx/6Mr6i4uOlXPW54f5AEFX
mM/+d+zxPATHPuRuN+UAV953TEfULHT+G3t55gi0fLE5KyLmzOEXyPjnNvX2GcNJ
39JvheIJ5U//1CvZPBO9n1+TIegUF5CdR7kaeXviah2qC2XKffP5ZbOZRxiYWDHp
v0+eIOG9Q1lXb6YjB60xhjN8bt85Wp94RrB8/GMOAebm3fRW1MTHSbFAwR8npkyq
ggTMoUgKDGC3wWUKRkcAnFMpgrhM9bnDbbLgI0Hpnbr07LrnU0S3tgyVJe1l0DLz
Kz/jJDlcPhLDDKnRxYYqJYW+AVhm6oUDD9Bd246t6sOXLmNaazecdqP4uA+8bfcn
09ngOpeLXijYP5BSPPOm8/SG0sZF/0zr2JBe82gy7msXvWTQXAufigrlLQUJSXxN
SwQLQYbuCDf3ibb5srtzGuP/ABzB0JRl98mEhSaKj8gtfsK+Rld2awDTQsKRKE+F
1A8zcTJ6nJHELippJwin7jSqBkv1baBYRlYWI42CIVHE1JCuVfOtuztrqrsWBTND
6ErCGfUG4WX82RwyukkSpk0p0Gmd3uAooA1P0/6MOA/4uaNV64pZ/jmmEiJE9x9h
qGUgdEgD/ROR03KcQMbdGkmLId/AxfGiELIfLuvkG+Uyu4E3To8hiTzcybJg2L0T
HcMkebymqQpUkWdYbutNuH3pKMKq7/Y84YrS7o6k6mixn/elbWXZFlv9KhZ87Cj7
gf2TM/laFJpPPZDnAqgVMjnN8JzPy7yoNWl7ZXo8VexFcqg24FTqwlEUmcsiOKVL
Zh1VFO//1XmXioCLfQBORdXYSAJIgEdTnrDWKvHh1bj7uqxMoFSVH/UeRf0wQeG7
D1yroOt7+UsDszaF5hvdZwQVhINoN4jX6ppgwv2C4mJiIBeW4JYqjJG8yn09nkUH
uMfhaXdSQILxZ9T1C5pvhVToa0R15k3zI4hEjktdGaTJI1QoQQO/2EZL0MoxcdAn
iaAXWiIj6MfcZnP/Jy+ClR7xA5qb8uxVHSYQtUGu8FTlkJEXGmStNJqlJllT50uU
Nj+2bVhkdZV4vmN/AqdgkvrsmyGVwfVv8A+c7jUdtbvDMG3jp34qyhWAm3kNGK9p
k9m15w+87rWrKSR/Ykm/HIjrWU8dDKbb/5oeBJHvj5B9zw847stSasqc3qtk4dkk
iefqE+ahmVJItVWINElxtfYm+H71RskdvaH3ta/LSpiO+Xsg4zHup6RymTXLvxW8
BF6R6/oB5119w0ytMORGMKrt7I/NRwOv5ww45g5HbWjEZqaDP9IRofJ9e97d+39A
epPqekBk1iPCl0oJuKcZM9NrOifCULP7R8vFtOP4sA94iFe7XfNu7ybbe5vlwzM0
4g1/9WVIU1iodpmfM8ooAI98e+GIqxwLut1dtnLJ8UuTMSBrUlQt3FBuEumZRXlB
H6QT3Q6zIZrJsRXKQ0KeeXrtPdO7J/ayZnzEPyP7E5C7C3CVmsy5PzqDdFCPcM7N
UTijEZWqp4ozemcIjXfWnb4Hwl6Mbawu3GLixjKnmmACockoD4GxCvJ9otgsa8b1
BAauhZoACz+5G6gIgz0Hs/1aDoqJnV0xWAyD1xVTFe9KmxO7sWl27kplllRyik8N
3zpF6Ks9sXSLN8B0cXeHXcsie5x64nGg2K1BzT5drlrr23DJDmHWTPoFudiJxE11
6Eu9XrdetKQNzgJ2YDUo6dxuyblXiUZe7m+uT68xS88On3eZHRIHqysXG2P4cWwi
gW95pGHyqF1ZiLfQGgVtiboksBP7QHqXkOVan6ipdMn3EBYTgHns6dhoRWww7lwd
7XAR8iszbgx9Mub+dU2p3W1aw2CUr1fiVON1bE+eATlaXOLohIS8HvuqsCCXo3Uv
gHRkJoUVUT9WJ2K5AX1dUZVzaQL4pA1vHcZbq6SPWtBcD3UcLaz8VhsE3T5lu137
bMR3mxfcdMjsIcY8J+Y4ADtgwTMMMrxOW1mI5OKGGWprWsyqOzAMk2uJixTsOTzX
oLX8UiptHCCgBG0DXTdarB/ANYGCCPneRkeTGQWRh1Hcrpl8/mMMcLxXxKatc8AW
9h9wrzBM6BngDF3/89rlX+Wd2bUZGyhtjrpY2jFmlpY66Kajf75guqVYYRVfFTuT
32ss58yxnr1T+G7Pa4b3HMJE5kbiYtNEzlDawP9Bff/peh+SBVyQs+KEtnc9tLit
mDUDnLinLGoPaNZTnwHCabBY/AM/oSXQyUC8GFB0lr3zmkP13junZr3BZIBA5RQ8
vQ8+YdMsIYsezPvVURN3Bg2ZskMgdtbXWNQ4BrPnM5xmmB2lbSe0YM6KQBtQLL5a
lnda78a1O5k+7sH5sUXYK42mRZOKesR5Sxs7e+iO7Y1NqR37qBTtwK9HNyTEjEID
BvBvM6vmwVg8tlCEksnlMB89B7WhKLYUm1iImoVjvVUw1tZvKpJmXvC84sEHa7ec
FLrYL7cI9Q403t+8BurkjRghaybwKk/uHb5RBSyjhWqfDMY4EWuhHih6gyvWrJPp
o3qE1EO0T8ANMfqjCgcw3IJ57q/KKE+m2QVd+suVHzQ2D66Dug99g+PA2QSyi47d
DP8KYGP/r43ytE6ET8cLYfXjl5KNVbjluD25ftad38ay3mrT30iZ+9BKjYCj2BD/
VOOy1AiWVh9e1Sjd2YWWcn4R58B7zTmUG6YVbfkK8jRSmHBV5fnyqGn2S9VTpVwn
yPslM4f8cajgdO9ZQpvZfhj0rsLkXjGM5o/nb+gIOQ9dO5iBwhxZ67eI2Fku2bay
pZskisYXIGPQevxm3DFfc2zne2aP3r43BbbpDeVmWx7SyzjAl/lah6MU9ZsT3N5Z
0zUKLdNg3EW/cugMvJN5clfzRmD4Qcivk9uHc+39vXlN4tv9QqDL/0DMPrdgFQ6c
nsFQPvfFTUSI6wKMCTMM3CHmpc4DlU/XIJo7V9M5p5xQCt7aZ7VaCpvP8GrmH0IR
sgGqeisYmF7CW/ceTqqbsAnfkI6/njAp/v9ayd28A6HxGV403Qm4p4rDyNoGnaH2
gdSML3GEqvzmu6OTsbIYrYDIDTbaEXnu7DULc2lgaoudQQmlkn6u1jCEkrnx/nwT
fpbuNwp0smHx819GbpPs7U6PiqEzzy4FFidYowj03UJJSG/VTwwEe3otYISr7YCH
nniCP9caYxWLu2ZWWq9VkMfL4XX6B6Ubx6XV4GxRSq32ArCBtHHaQ8n1AYrqjHwu
7FfL/HKPs752s5ecOJKnwmxTXsABSaroW5gvSHVDfX9ZE9B2CsQVlFVpnYBOPH91
EReO/1GupJ3Ra/BixEKpOLwAlQFdy/wHayGXg5tOgVZJ1rhTGDTUN+YXIp+MyNzI
QseRX754CZ3UZQER/Xv0vmOT0xG1B10LSw08R+XBh0hknRSzSoT4aPUSGxsYBkCC
dtZlBfQhu21gI/XdOStPA9rJ8QItmoxA4AI6Kny+KvEjSLu7hNBTwaeTvYXG6RsA
fvDj/enqGeNqGnxGcXXp4oyHH+eTxmC07LEGi0/NlC0Q50T7mnyoVsookZKFViqF
C3QKmRdkMEOIrGG2eupVplp/fuw6kLLRBIKJdPb7cs2t/Uuf3TVwmzm6R9h0sY+3
3KFjbg+76/kfVSh9A9JERLllik3EyqQTEBE3u7f/w4/9Xhz6J8n1KxHK1a7nZ6gE
6E58kr0I+OseujSeMTg4xqxbzwkR17JfDVSQ8DtN8smTzSjjyTUuNO6MaW6xgPzV
PB6P+zV2v9aniGGIrNGKol6eJOn0A6piQ755Nt4uMD+Xr5LN5du2wG2I3IcoTzQu
bkAnkvtVULU9H5k6LRS8oiZRCvjqj/VqWLp3xmNn5QTxUb/g+F035mMC26MOhX4e
Tf/xXCU87RCqJ/s+dBy6xYiuY7TXTSIDjA0VxfY0FuF9bIXHT0YaQgddA1ijbIdC
vPWKO5kzNtJpdu7k5snXyVDLCBakcdqOubIMEjYXq7nPCAUAhW7cxKzVfrUzAC2i
qVDTqu6Y8bSz/kHJhIbNT3zvQ4UcBmeh+e3hW/LR5u936lbNkd4a1HVqPdi8HOyM
b4SqU+7KPGLBQOhi0j8WVI9aS0uZJgJEmYMiw3QIGVOQ6kjKkuszN11ZF2u4dn3K
Y+lUa+JWxgiKPoomLSf/NWHuFavcEt9xnouv0GECOhAzEGemeRdIF3s65luTGS0N
KvWKZ4f1r02Piehj0sIYH5vDJxyyVSuLuSqe6b7UV4mNezHGCuCMzgdFQZ+IuXO+
XfOmKedKvKPAshHNbcCvBlj/f8cid73rAFhH6JOvAxv8p7k3CPNwRtWX3kcRmwOB
JPTNRQov9C5HsDQXOWdkSQ56UMGKy6s/bFU6rRj8hhCNczouYXfsAnqCqJpa1W8H
UrQpzf28pxYjwN9DKnhpn5J+eVS33Nz7uxxNGPme0uyJ+kZXN5DsnvSq0DOswfWs
fLCVYSCGQdVhn7mX0T9YPtUJL9AbbKoqTbIkWhfPl8dFZmdHoW3sOzntYi5d5/rF
J2dwRg3Q728WCUJHUZYUvus7zC+TLu/YlU7b52xrczODA8M8W+4IVNbTGORyuBDl
dtdi1mpv37IQpOR2Gl8gs5q3rPErVO4VzFVi4Leu1flOYOTsd4D9tIiTefH9xJCF
d0r8d23KjCHBtm4oUizlPzuxgTQi8QIfAnZomgPGHaM/KVhqXX9AJ42yXeaa2ULk
H9m1SxSA2acQa1CqIRS6VZ2KhaBnm7wKDGv8EU1Xrd8M7nDtb3tyh386OktfZjsV
FQrKe2fGzxZK+q7CZl3Jsm+q7Pr06ByqbQRpqrGydBiuqu56mcrSQ+3LSXOtXoP0
yUbAbOCGET6Ro6a3+40Cq87WhB7rfFun7lNgeeTKaxW46Cd74Nh8cymA7ev73YZV
8Rbzg7XmBxZZCoxMi7ag2beARW3M0NyWYglqA1JeLFG8LL4SlKSgXQbFBbra9n8q
iuD7CMmUanloLz6Ogw1JDjsiR0y2P427e7DW1h45ERgO/nl1b+PrJ2QOTUeL5whR
lED6wh+gvNMmtlcGN+J7yKkMBlkVhZM65CqtzeXXxxMsrPmmZHGcTHZgBC6OuG7S
kYt2JbdpBCWjFb1jNnRO2a33fWNjv11ASNYNWYLNjzJeAXikss3/63VXcTAspMbw
N6W5PmAPEyd5rMfATDpQiDATcruz1wTMh5w4LSVUx7MgFKwy9hAHU7OUPuKeQ109
Y3eawniwrcMeF5y2aVgICnIUL4XSd/x7TxZCJOuSX0S6ww7cwXuOo2mdYHIDrU2F
e+qGowteG72ClgGACScNyOzRr+sw0S+SCGzKUbMC614tbrxKyoVW+aAhKx4gfyha
3gUJz39Z+D70IuhWY/X7WogN8gUvpfOAdnyndLE8Qty13kq8ki2wuvAdychjzIio
DwhKc1szXg896Mk8VYpj3L0hT9c88jH/4+8qd6SxBx+5fE+5A54Q3Dyqf65o757v
Efdjlg6WXDLemrAE46stbpkEjrqWEpKcaV0nZvKxYw51fW7u04rH92gfL7c6P7u5
QRwZR4T8g+1+qqrWMmZF4b/ViO9AZOirX8RGS+t43pLvupY25/fM4QivYrw7QOMa
5EmrNsfkknjD8LuvNAwK5DWbbWP+gqtFf95OO9OEyto1yk2kBwMgCWgcPZbqlX+P
qjNfR9jiKSegX65CNw0dEXX5BAP4yQpg/33sLYAjFPL+7IAPQjNJ0NakW7c295Ou
yHrGLerILsg64GbfMxBgIb4rzlSIlgyznstKvIFadvEHq/Ep/LdM92OQ6T5huE8k
swOxnFvE2t8ugC6phZVBTD2szZDezBFD+QhbQk7pNZsbmr0nnHsdVz83KkDhd0qg
08zkWvI5659Fv67d8PZkOwvDyxI4AX15MtKqcdC90V4uz7BtdbQPFWOIR6rjdeWP
vQ8KALb9FWC2Dy6RZ7kuopqPe8hq+HRz5KlxLKll4qmbTX0ebiHmRc+fs1okYV5c
0TDfxHuOQ3oun/OX9bCHLeZNuckhLv4YuE3OFm3faI20g1q8wT/WiLQLnYR3FkmJ
Bm24PWnLvEWdVXzGvG8uBFdSW6At/qMmLQVgbvQLoULf9yE8idgi3DgJIWMYKLoC
a+raq8YXp2KVKigxpgI2n9yNQ6ytFgYLLstb1VKl0KuNvvV1WpiCMf8ejFT+Zceq
jkVC+Wt+/xxZgWkYk3cMP5XQXaWxkh0amXiEHVCvepn0dUpP6Xgl8NiyVYa1ye2b
tO3Mkv5m0zujNmtej8a+nP454z5z1QpNBzISyHCyScBPRvW4blOn5ETSEAbBQ3Ke
IcWqMqcYo1NsEbUvmFpHGvEUVQx41jVoIsf6VyVFLN9MSbS7koQ+UH0FmEc5b/Yk
hU8LSQZuvNFnajRDUIo1RxWqQQidBHFsSsT/VSW8UBpjzWp5cT9wqOGrlX4s7XqA
7x3zzw338GDckgOVasJafD6OnKJ5/Vlo+vOX7CIODeTInr8joPPIpo/0GaPPhhqg
tOvhUWAzDbLjbjcMSPBcTVzkz4H7QVKolz2TJvqHwamg0Gm33d3CVQ/WQ4NWyCRA
J22dLNwbEsszM7tImo91cDayrTO3I804TwvFyAw9RFVG+Qh0cc3mE6/CGwBHQ3et
dpEFSYJEKqB7WE7PlT3QdfP7ppK7CsWU1sPhwOQsfko1jbKkqoPSJD3lJuyBPX9D
KrZJcSPjBTs4Nd0Ok02W4CQ6jRNfW8u5NQnXX3giyaQ4Zr61QHaN0fod8ZSs7ihl
TVCEdZdnk8nj/v0+Zh+LVDR05CrAjZ/zya/ZAemvIgYHj3+YFNyiWprFEOSuEO/S
69R/2YslR7Lkc5YYXTxDkbd9lxgQ2TbrwlFxiZbmP53iQZGWj7i0QoHLJv/9eygB
xxTz1rzahe1StPU3djtOJ9lYM9/LK0ZkoRzzhM9w6+8PEUOhdiI262WAVj8sJzHj
/sIndOFh5bFjK0MWdrAlVl3xXf6/pUDKr/eHR4MnCw6geg96Yp+MguzxJadA+cwu
2YjPGgJ7UFZ2NMMJE6bN5RzuZ3ZHg5ccbtBBXZNk68+9fD6g/Jv1fSfOdONPBWUI
GLQ96JiCHMmFwfxGF3JpWlP/4M1dZQnAUC/6lpV5qeamOvy08RSuNCkqKio1thAy
fAXtuRMXNXW3kTGnKKQ1Z0lWXqe+aGS7aDYTE6GozNU647ajGz8ZvhDsLip2wpJw
xMIqtIxton/Z/tkFBzrum3GXhNxQusMsHPIUY0fhZnw/s5CdDpMPNsUlLXiUqCku
Spyr+Kt5OEiSAe2PNh6+DbTldKlG8agkHE7BI3Mpmefsh4TptyfSDC6BWnDXfSy7
03UhwBQxbSWNjnBwd8bpFXz9aEX2Z2ihhq4Qo+hAI5Fda7HKbiw48peydDWGlNbB
EkuvmMirKwWzBJM3cC+Pbbbs+jXvJVM6T+pCNhrM13nSRA+A5BxfswvE1T27vKNL
ltfNA9BtUI9OtV0jrijCzCxV/xEl2OAWV3tH+7GAFdPkHyrnVmWQ4jFIJgl8ZEpB
FnkiUUO/wY2z8DqDqRHv+cRMlHTF83ZLAEhFfYHtSkwg1Ce8qHdofwXQkyUMHC+u
mAkr3hLLhBj7aAdWuRpYLR/VYkfLoOO+QDN+nJ8xt32IDmnIxugf4f7xpP//N3ZG
nodGRo4hqJwpjra031JBXmcAFaW7pNBT1ha8xPY3kl5hWpeTA9ZNcdPWDa6zmQl3
EYBAcfJhy8ptLIu36FO/w/GL5fANv9q5pVPmxPtpgj2eoeVskgX5QM+Bi01b+ZZZ
YqKiXQhZF3TPSIuA5cZsD0q06eqhN8dGtI97prCa7B5DkHm/YSMZw6lqIeocyt0X
mYa/WqRj/l0EKWqzzdkEOhf4/M7N6lMKdn/tH5ymLM1tYcXc/R79EyPqmhMfahPn
dmp7bx0LdF5P0yeKfEGSVQAZ1fMWofC6vJGavVvD+XiVdYvfCU6odi2yM+PTQ6JU
9orWrT2ZwKfP78nXR1WAmwPkSMAcXI/8CqLOH+pYFNeeTWWibYUb/O2CfY13Zlfl
vfsHa7puJam7RZissB0Aw5lnMlbVkZ1u0Sfb4vd/rscvbMzjU6cA9EcGmJpSitpx
bd90ypQ7yria4BzlvsWUX3BfGdWtEcoT+KkKJyYqyStoVE6USrtoeOBwKZQXxjGU
bbMwBLNgwsgQ/UCUhRiKi5CT9NTzxW5Y7nIJhPNE28mBAttHHCoz8f0FVjIdDIYq
bPiaezvSI+c16+venn5pdG5Z+uvv/1JfJIiLuvQzoKjoXggkLX6HPsQDz0uisd0q
3r6BvCk6psp7Bq6FFbYgp0DH6hnDmHwkO/gfcg4Thr8nAhnNt9hu0WiVAQ41eeL3
mDi9JoIU/p2HmFQFxQjw4N2m12c4znyP5Knjb1cb/7K7RULbA+lhQT/aMdAnu0jh
DEIciNgrsNDFwKbC5XweUrRIzdxTIXZwyG4UHNk1ko894NYfMuXGhyX9HlodskVW
Ob8UzYb4UKJMtbmEwm2q2C1s/O9Hj8By3qu3CLlbXUnl80yYL3kzjlSsyyNsGdvI
+6FG9kAHItp1gYaCf0NDiD5zFCRLLDoXtPP/6DyXqT6oHatacAIDyBJJUZ6MpWNT
2mMR3darc+xEEdk6w6TTTfJ38QtBAcxr4iHMEog3jmgY9V/n7ydDbXiwLjpfOPsH
BlsziDG3uHDdS/3pTe4yfQwI0IHNvnDdCG+i2hHDFlkg23fxxxd8Ehx4ALnJVSUr
La/OGVlaFxLmpvoMD9hh60n5mbwG3NDLPAivbYmLgtktJwrhsxz+3Nh+V+OeAr9R
UIpA5DOl0+ZFOKUOD1Coh/dCIKT+4MyymCtzF5A19qbN7ffmkOsZNIMCe6LageDM
b6SLXGIAwZOljf2Tyz3Xb5ZP5hIt0IG4IiEwkBRpHGJwaqRu4om+JR9Y9PNGlnmi
6GX4QxLa4zNkCebwhwRZp+QMQuq2KxURRo4LcF9nkQU8ojUaJGtdTmdEC3IOP+KQ
zRGoT4hUhDkrr1GE+6zASHotftwCerMwZV0fxuyRVXb1FIHhNuL3BpeWQPS8Cz1W
LySmyICK4SM3ddjNmP5biBgfYx7BcCsRPKwiF3bDmfWyL5RvlBwlJLxYuy8zIEaM
mWDjDorzlNrd3TX1yd1uUevUbcUO4GDqUKm56aagXLZLAgurMx0+GDdoKbCBDl1l
g3xdHzhnJGsPsgxv72KBUSPslFt6zMCmRa5Y4XNI/TkZiHOczLfWdxHhUZprRNjb
9h0bveosvewtl/lhUcqThlOy9p7zMIVSgkyk9AUdgEmHXd+I6WhRBX//BW3y2wJo
yBf2xgjD1iuZmuEQXtRF+3PH8b1NE3mo3X0MvECduQr/ryreghpcqKuQXsLHOa+x
fzaE5pS09h+umt+Qws7HMuNVauMMoOeVYszlC4jjlWEp4EgBcKAvMpZRIAZEVgjO
uspkv9r63h2UGS357YzuomJg8hn+EVMRUKgoINintvD240fuRlC2eVg3pcW1cGmJ
Xfma6JiqzilEhiyqGvYBhFeMS/KCnUtOQSyLxx5RipYLT0F/xtoj3tfhOoZ7J5ti
jsnpnfomG8GJaeMR/fEKwTpYSgLR3macdFgCeuARHT0ZtORoMlgSq+M4k1J305eu
JCcqfx7qwjm1B3XGXE3rlNPERlRIjJ6tWmnA5t+rX0IdrB9oYV7Iv7Ob0jzs6IxB
q7DkXJ97VFDsIBXTkOVJan6AJdJX6twjRlhjU+54NgLR1KsIVSH1WRjkwxmWkcN1
XTaR7wu4BAG8Jrt0TSPnCYJjgMoIBRzd2eo0mvPS8Gy8I/eXcR42k4KtzDPV2vMa
iu3uwMJYVpdYcgU9kYgCbM7kRf9/XDpYVXAlY9X+VBAd7aywovnnqiUP84mFZTpV
+BRMybvGs3VvR5/9TEpeIvF6FmmaL4+H0HOCTCtK+l6imsvH+JhLWo0h6SWoEn9A
h+VQUxPl3NtzhGdipDrvnGvyT+U1oTvCErms0/BV7aPTnzy4/JJ6wm2tKU+LuHaf
9Fz0Pw31obYFOhvwza6Q+77/hx8MO/vGg4czbDtBHdSNcAzX9QY3DsYQPvdgiVQG
C/oKLx3W6EBq/UC+z5qF4ZcjXovo/8GH19aIhkb+iTLLiQtMbXygE75p10gza5kv
HCz7uP3kGL//OF6w+Fcrh2RUtPh++OWcBYBi4dXm2jMgDrDoJ9ux7djRir/fKMLz
qaY4YDK++hkVAyI/TinG2dHY5Q/PIfzn6yFf/QaSqlPIQf+fmA8K3j0FgZfI/gYa
N//0qzhjMODUT7IG9RNG+8ZyhGVU8WUl/Vp00CjKE82g/XnVGMGfYvaWWmkiZ0lQ
EPcNL6rAztjYWP474ovMiEN+oB7IuSm6kssz/4VR3BQrNpzZV4yDo1hvV9mm7y4O
GFaIGRrLeUnfL3W/7C9cevLDp6noG0xl5uS8lgLk1lniDl+ph+yePwaz9yxo8LLR
7QDbprQihy8vII0IJPzj+MMGoaQ/2wC6nE1F5GxeDurrXCOvcsxL380ZXtoTVPNu
yqsJoBlcU7kO1LJFqt1zHn43qhr3xObRgNJmEnn9ORy39k/zbpKu4W3/htTa/dix
PdA7WBpSRahs1RVCJ1UPcoLhdPq+D0IptAq3/ghLxYqSFFYvzwJ2IZF457WGrESe
NVHdsAjZ8aFIQIae0XttIBIFCcw+8aO+42H84WM2ot0wVQLExv5LPmVhxRiS6vPz
zKQCay87nPzj3f4A5rj1aQ3SJ4If6ONodfFvbrDL9pzlskYCUCs5lB3wRTsyIjNb
TEDse4MLQAFJeYOAe84QCHjJN/+Hc0FwJ0xlyb+hF+19oINpukcG4ubHo3tWKHSE
nQLY9Sj/tZw7q8L4B2u6ouJC+OP7Kleh7Ftsk+NTUWXlSmsTiZaJNSa4b3mLNWXa
fdrDjNLzdktlsN9TET7vW0EihlGlIxTFObr4ncoYCHvYWzqG4rbFq/4eATiXuVkl
asP7yFmlRMK/fMRuuvHIlvN5xq3KTb886hqaKO1NifGvwnfFvZonkfvxdkHYNTAZ
5gCnl73Jo/nRCq+C55xwHime/PUWTpQ/aykZ87GiOlxJKAt//K/pzobSf92kZCDY
8N5PFUazZoEFUGg0G6xeDuuzP6W2k53Fjizg574w/wseroAfj6Q2NjWHq3jJYjLt
sGV/rkaPrQMM/8nQji42w7svrKy82wViBV43f+UpuBhIKDnkM6S7woAbM+BbCtb3
cxQnQ8Z2+7tikEhGXuWmoNCaIeiQmWtGoJa2lqw3LwzwavqlCbvTclK78M+xxuiA
jCco+RJr7txck6OUQwqCZtNcXZQPE2/icX6gM9osYdAHI/jzgGimI8sx1wDTUbm9
Z1r4CB1JLNcmpVYmYigjaCaAqMV+Ihmw3Ri5xD9JnFANKsFzbTUHnNK5NAJbu/We
uYQCfA3wC7/uFS427CEjl3KqKnq/TTvgybSiu2seudrQgGoxMItvxJfgS8CIJqci
Fgr/Q0tdvlbJ/7kgI0w1lkjnbIUG9oBKIZ1zPSB6WzEDT2p2hEDIaTHhAJvv62BF
9i37iTDsYRdPafIvpL4rx8jVo4Zp53XETBjiuvCH9ajv82BfIespenUGYLjrofSb
umQiS7TEojSZ6xLshWpdT073jb1PtPpU3D2qowazC17NKDs+IDMmyblkBumXKAx2
A4Yl33+Nwt2nocwSRIhmh1ZCCLz2oFGiCkf+AwLpPPaNasZMHv+GWSdbbbpnnhnB
GTmPYtoK6FR9tsE4WZyLIsDDHWKTxrDZ2huP2OuHwTw+AOgNLA/lAfhSlxDtOiFH
XLO681oRCI0vkPo1eAONmozI/2UtFaW+UbAEYSqzAkSb19IMR1ux164toAs13cJK
ObVk8CfxeHBgX1AIcgCIuvcVwraJkzxI8YAcEu7r/BQOrUlZjnOmYWFX0lhGplF2
yuGg9ki7a325FbKiddND7wsz+coFEk12i33eef6wbvjsoSHv6/3uVrAJQmLCX8sj
DB5QqgPVilUL4goe1oEC7J3GIu0ZnkO8AYxm0UTMpxZ0MUIZr3yj1Lroo1XFM1zM
O8IjRTo6RWRfop58fdG0gEdEKH3611vyc2djvwe9vHyi4RR0ngdEOdjZ+gc4Dk7U
Y7yeqYivbkPhAB3qO2YVZ5DlO+Qf1cwzN5palrcCHhAjVQPZhX1Lb2LhavthF6q4
q3b3cHaR+dx0792xOSODMB7yyfi6Mzb/8ADZqcRGaGvxnYjABHCSuCWjDoRJ5PtY
BL+sPLMtZ0pNey3cbv5epy85Wy+NRZ3IzbDnf3xnFlf9AlRZJ6Bf0lg679wNrcnv
Do0kvAvnBHkVO11A/bKNSr3RW65fY2EHp7ouhfqqS4mws+hv2o9Zeo0pOxefYruO
n0/JteuKwQwyFViGXU7G/XYK3KhYqoQKyow06Sg1DbKrIgHEOsTh5IU6HRfI78oG
iO76D+WU3bN8KF1casNsBX/er3jcYGFFnrnb3nrE33y9DK9bE0aYQVrv79zFR7C9
F0bwWWSjbXRrnX/yyk3rVT38ReZlVh68qHgW2jca47ebo29z5hj1hGP3jxhLIkSN
fGxRraRHxrJpKhL4lMTX7sd6NXUOwW3RplfgUfUxXWv/VMHyu46jnXOp1yYP6amR
Z+QI2tweLVfFSvBD6eQJjBlNLp+ZPy4JHCd0DbO/ajkansymn2qmDljFP1AWLG0S
bf1FruNNVwe5D7JmDB+CSXnZkuqpzYFMNtrcklkUzNl6dT+AJed6wTJ+PneFhhSF
dAundLbdI5juPnYUPFE6uwYjTCnmRBllVIFuTi1CvWnr7rTx+OV0FGa2NRvRzeXg
//HxFg1Cm5RDaMvLgTe2PBl4G+awJFWsYAVNhWiGXp6mUv1CFCZC7FMEizBsYjHD
hunU25CtXE0WeB9Fv/3E6tkV/nA4kjgdVUCHpHFlAzh6cn2UM/eNHT4bq/xDSgKW
XND/3HtinB2rOD/T3ihwy4YEShNMWNichDTV5WrVWBVSxh/sr2Ju1uBXkNNXZFvI
Js+OyZx+LnnI6sSeGEW6SyKfwk9h+wv4QvyrfmewrXjVpl50Ofz5gRWdUF/7498w
W1a0wuekIRuOgZzxOSwPjsWEX6GU2GzD5CaQauq7wEDHelId3OaB6KUWYrSyh7k3
NSw0733ZGkM0xEfQ0uldyilcBP87Ze88dn90LKWu8q5X797A7rjNdMWz1lACGwwD
XwjNDGhze6C81I2D7ka9rcyHIO0uLek3yEyh7fEnHpruJdo3RqvlORgK5yKiv0S0
sE+tRFD5i/xGhbV6Btr/vjGNtgTfWn/yu1Uot2iENGieMvku1BYF1CiGJ1VuUEq+
or36XCbUa96lwK+gWEd5mhkWJ1G3lUEkimruHupRLa9+JSSUzfV8UlQ2I2S/Qb/i
A3A9gIqSjSwHstmNPZ9KDDyfLI30m7l/f6OtOf/VuKM06g1aXIANykakQlF4f8au
BMCWGageTR+b2u17zK5Bq2+mEa3iCNXVerZrxF7bUacAzaFZLqaJSLJQURcwnDM2
RK5GcGEBhiSACCw15lon7nUE+MPmWCuQJkrvOZ+//YNN1mnPRSn81cBWoSGnEmo9
by/sPUz+L8zDV3jv6UdjMbt+Zo4aTei9KSBFAFnJroZg3xBpCY3+HYX78SvVK4OQ
VzLXYjRDpQi9ieVruRst7HnDJ4N/EDopt/WGIl9SNLnM/gfL/Ida9+P9qfLP7tsi
79PAz/y4sgeGZNP+pa7Xdjibycgn5UlmgrEh/xrbJ3jfYCblD/HNnInmhOFJ3HbN
sk/6lDa2MUDF3KmHr8ofG0gJvF/2BMsSN6z4nktwtrcwxyf3HF13zrtVOutmG7Yl
JdMYPKOswq40dCTack1GebmkKAM265eGv4c8yuew4U5j0kp12s2MZDuXNswHn6jf
qdcKCxRS/vSIRLSERLYiGcP4t5cAoaoQyMMphq47Ano8HdAX/dZMhxkeC/2pYx+j
QAD7fv4TEEqZ3es/kIZbI+jKHIeCi9+/YQdfVPtZKQqdemha4byfvA+vreQAplkt
sMndKHHQYb+f+1qk7NZnaVnir78xwKBhfumJ/wPJ3JAlqMGSMpQknPt7qG8pZegW
dYIgeLXnyj2eeQQaOP5HtG8JqbnnIi3uGrgxeNkzCY0Q1VS3AD05HRJrAyG83dVW
yZdye/4q9IUyHlQGjuu/w1o5++rbb24KlFJWouMWmERygBNdPd7sOx0aeHSk7Q7B
7xiB1xwD2kGyp/6KhdY3Yd3gNuA0l+GHhZKl0ed0HQhxSfibX/xwlNGTozJGOCPp
aBVTt9nACzmJblU4HTF0kBblkiT3R0kvWhJuCWmH6U3gcOWFBDqRwJxTlS08sxFo
xXADJj5rIA76kNjI74gsqw4PfMxNFe9N9jgfmhBCBxGqMEZc/cA9pgTagT9lamwF
WvPlhHGTtkksG93nBcQ8QrEfgc0CSzTFNOijqAZAktjLZ1NbnMhDVeHv/JBG2Ylq
OJZOLNz/uokYUTjfiFqjZj52dgZRtqhvBrBdFOSyb6hLdKqAS14hGLJhxaymV4he
PaubytJHB4w/5ZHk/QxkipzNPdmPg5PizgHzEDlqRqRgHcCWHYSndXQWsaPm/CoV
sSOml8Zs/RlWjQb10Hqb8M4Jo3LDsLSr0rRLYEZ0rBejHVtYFIPUNvii4+krtECZ
SPSRhmTiwiBm8I4y+GG8kEDwKmGUMRhueY4GhtSYHJoVu77BEh7HVdQguOnLAYzG
MMnqmEtRPyQBmnCtzNAe/2redZHvI8ouqUAUKl0h0e0jW395c4JR3vzYEZ95ZjFI
xJrxrinQyZVfr0gTedAffar21uDGuIdP+UOmoXWxJZW9CivwlwCUFt/8D1VbVTIl
48ik4lnzUKqb1NGR5buxlw8AA46rvmsrnC2TZm8j0xDDPn5cPspV89O6/+gj/7on
PE/pFi7S8eaJmB48/Bjj0+7kCP8pg7Zfc9AiyXz1juCQhve34pYNv4z9DA4H3Saj
ZajgGJmwDxrFz5QakrmeJdkwEvFM7as4RrXUsxBjY19ErrBUGF0PqY+50N3+3WLB
t3pqOUhEDp3mib9QnHGqFVieQ7kTajwFk62EONp2MTXAgEOXKwuRB1CvHVCu1AIy
B/DJTWCIqwFUQn2v4V6Tdvwi0nggiv+I+N/vrNkFkfrg8FXvZGHSxibTQMO2xFbd
643JcfWECIYYeHD86elGk66XtmfS3fT378QSZeifaKokagykwP2lwwVW/unYXN/a
RyN+BJxc/drCNnFepUc3yl8oZuTCo1kaQJuDO/B0HYRLqOJ4Ngr4TFWmCs+2VIQ3
UVem/sG8JINoelXJ2uEPps+Vj9ShxLHzmxmdIbzLwpZ2+hRBNtCpUJtGjvHlzXMT
jnYIdVSqlG6X1RzxYqWpQOMNAEwtOoRfqK4mjm8yps+TImkNKMdfiS5QPAgRUdf8
IdfT9Fqyw1M49dlgQgsL8ynirTl6aI+cKHI+dCIhjy8KomNzUfJKO/gaSXjjXRAx
3rqpvY1lDU01ZioM618Erx+RRapqdu7vk6fwlK8+3GaP3YRqbeWc2Q5Eh+oNvvdB
5PtFhPo9yf/FE+gnAzJMwamvo6/MqOkbj63kqIoDV5u+UX/6JW+fDxxQ2P45A0si
2wAvDVsDfz1kik9/qYozFZysDmQuJTotnp/AUOn9fWpmhH09k8JGys2t1U9M2Bms
ynnxpd7uG2eEKifWnY9sR24NmtHg0Nd0ayrp1iZ0GF30T0Uilf235spYkc0ap6jB
245Y8AUJh0MeeXFv1YrKYSUbs8PPLiO1CJr8vkcHCfA5DPQP4PpJ1BiXgAXTHZ6a
kpJ2YLBkjBDVCpN/NYj18FT4nvzBexex6dPzsDbjC8vA7/8Z82yRMiXYfE6kFSLV
sP85wB2Ep0/zwFNrMrEq/bj9FI/khCADAW1SxUraGzbL6y3AU3Rmfk5s4lOqa0vH
gSRSGWSlKUC0YVZybEl5mfhlcfR3XyptQ3dfxofhK/elUmLVwbqCWfQjBtY9PfAk
exDaAPIN5OTLwx+/IQrX5L42pw3dMgHpcsZb/yLj7uIC84nElTfrSgIr6XHcdKDx
n6F6L5H0jAdp2+sgCLgjN821PCm+KjZiM09+hoU8pRmA+0eCEThjFtosAY0cJ4xF
13QQAt04EaFO/wFMOSNzZboF2Xzw3bH31lkNJ+auQPiCtTVGKv3wnz/TPzNyLJa4
MFCQImpTDWNTbyl4O/GBnpLUnN/eUOlVIImPgOs8WqaSaeLWfFmhuGDUs/JU7o7W
qeTJHMXP4TpjVqQNvqRdY0ZjNXSn76DXEg6xO7lGx5vBfCgCjOaKt2nlfWfoc5y5
BgyKx1aDHqQZ9HEc7edkHz5ut/ihoZb0SD3C5nhdP4Owg9jWEOzliZAx3PJLVA/c
6lgLZ/IMPQ7A6T2VildVOpQXbJYW+JGb4ZW/gFE54hdg3kZemvHqTq6U44Myrpn5
nDVv5gc7oqpOZ17MUGkYrPzDrpvaciMSvg0WUAF3YOS5VcAXKNSEKe8+qZyxn4Yq
1wwvOgGT6HaHieRp30RdBTbK53L+9Cn6AZtEAtWUDnlR71RSuOjCItoKuXolOrqf
s4D+I7gL19tq3Xt/5G9BOhbvttTuCzX1Cbxu8iRW6nO27S8iiUdL9XA+eTId1XXl
Ruk+/QLskN/cUvgIl4lnpsTvHh/OcIdktvKozEWpoHuEasmBFIiJwkpOcexsBy/p
pgGtGEdOuZEHOpKcriAkpOj/lbMVQxJzl4BNvzHrHY7DDHomNaqYFHLqqru2N3Ip
D72pK8R8PZfqvtkd+HdF5IobZDT7vNwWGd+Q17tKTshzF7vP+ofMiKVlJ7a3nXEZ
FAMi/7SfJ9wUj/wLzvAp+e5JE6tXg4aS3MOHLFdJgeIAsqD6ZBf0b2zR1S30O0wl
zn27Dt8W0bjTYi6rIBAXQTs5yshmYPU/Unxl4RYBZqbAKrZdDe2pLNTSMxAe8jfn
Z4y1wKjnMZXKW/Yz3cLG+dJ6yvHem/y4ARl2x0ESsHXLvnf8PeBipD4ijuRiL0s4
iSwsnWoLXAWRYWM6Kd35VPZT2qDhH5MQ/0yjRLM1e8KAH/KQZc1aoLC+F77xubtd
xkt4LrTAJ3eabNzbV6MGwFUqj5So953BrOW/0Qfy8CbpX2FKHL6xU3mSA1YxZp1i
ptPuuUmnO1SumSTUnY24F6SwMgJ6/vUy1h3bfOEvBWznvtFId7APd8MJoCQNvPzP
wT4fTrs7LEBMtblq9/vSQ9qIsflWbTHcFeEHuMhjThZCT33fTmbdTIjldvibySHI
Ru/WIrWE8NUkSL33ZJAu6eD59K9r2Pbw92ZcJH41kEKIgR2RxpTdg2AWzY6zdZf5
FS3+c5q7BHmWfBLjgevRoE1U53Asf/r2ZYHvThPXkH8SN1nsArlv4lyY5OQnLBMD
EHYahZOG8Wt+oxZn4CcPVQH8RHmBHZm/pQ4IkIUz2Vx4lbY4bTAQPrMma3F9kdxe
DYkaCKFyskEQiGA9CfQzbRtTSTpbd4u0glvTsq0TSoIBc/jOUcHbCc6yNLEKvW+8
/GOXXB6yANu3eGPldOKdSCsWyatnh7SkYaagDoqOjvNm3jjWg3KuMReIUpqr4tvG
PS8OkWf9XA+HYh/JKuDI2x4XWMvqEmP+KCdxUDu3HHsw+jadhDEhv6G6j2MIhlQd
dLYDTSm992rH9p0D+YTCo6U4eGzxpE2Yv6kJ3pKgUyNP71w1YqoqV0tSSpyFkPkE
XakZtkeqBnmw3aTmB8R6I4FzBYg+KJjNsIBZaBPLX+jKAfwRqKzKQRhCh0qmbgrl
piX/aoZuWenWCrIDcsula7t2rLAWbmtop0TMiY9zH1sxyugs+iDGnubhDyY75+xD
a2Zgy16m3/LfHNDS/bTgepSDdBLxA/9REe/JaZEZNFn9Dty83Y8CLnZZd2L39L6N
N0eYkYUdNS1M9N0y9NytBNqOqsc4+xblB7r9iV74NDmL2D9qWDeD2UrmdexBZcSv
Teaj0HuXDhVbLWTcsabF0dTHSVjfEt07hMVSMs9MoS44kpt1EpOXJdwl6rWxImtR
VlUNx0Wxbm+4RX3hX8X7JtZjxbOTa6V8WbmZJIRfkyzS2He/maaIp7yw1flvHMFf
gEy1XTCYHCHtoyd78UEkY6mgAov5xqdizeqDiQgdAHLclTrZmcjtz3Q0ojDyX9+M
bTLuwHUSWihVlU/7bA+0Y1bkY/aJ0U4PUCdOtaMkCTDm47hBD7Jcgp6MwuXAcLie
sOXL6qZWWsXhoEVmueltI/4Vgdrf9JUtToXBqHoXtzfuXAKpKjZLvSVR/JWU7FYd
Ukz9FYneFkJWvKH1PJWHqlLWsP1TQGEsylU8BWBp5p4OFsWfeMpdwLTTii4i/r5a
F9eQmPXssraMxfdlx9kZHwDxj/+E0P2FzBYfQI38+Bl/TxUkbwvQGJlbw6FCcG1B
fazmo8o1r5Xt8btkRaIpEIGTDzPztBflUsYr67bRcCwJ0blpwhFiMIpRH37KQvN8
z+IRlXGQ/7EhRinBg1fxz9T5XddJvNjlATG4qgiFQrttF6CEGtzU+1aKMF7DujwP
OFjtDmDDOul9r899S4Hpo8gqkEpEYAXbxV4IgFaSs9LVWLhLEAAN/MEMrtzb9/vO
lZqwAPxP6i7Hp8kwXHPLvdp4TUOwm5Jug8uoR0+4XF3ZNPfW5BITK6Vf1R2euvmf
++kyvNv7cGwXyzth0EYH/El3UuF+6f6DeI0wGHIFvFLSys5hooKuzPlGa6Ev+nvl
93PSWzcDHsd4Mji8vHUW8itVJX2c3k4yUhcBB+BBEyJf5w0my+2d+AJG3sk4mmnj
I7itrOpNAST4plmj8lp4wVP7eCieu6r9bh6Dpxwa3DuZSt7pjplZsCMY9o3fdkqt
IJH9YXixwgDsbDAqMjbpXJbfnCPuquMSEf3oiiQee0LAI/DK1adgw0ODZrS9pCpd
pRcbF1526SwICJdYyG/2tt4hBd0Z16Yo6Ez3KA55+PJYUDmQnXezcrNj+8PcrZes
fYyoYK1d24fFXf+kcy5xb/5lOlzAfaBjY3fQfgXJB4L8D2yNjgV/vNfI3pnVGu5L
+W9GFIjOUNV2UAHIKmcLObQYGjEzdE11W9Heu5/zXp35ej/3xq9p+Jk7cJdnjy6Z
OOlWfkwKyWayDlJun9UnGasVCFs7aSYN4GlozvWHZqkayL9mpF8qOUgGbykaapCj
nRNQvZgMP9cfu6mG7UKTZIBRTqk4yi42RZcM6qkpeLhHSFBSaCIC7CBB+yJt1IVP
UZO4oBeJ7HapcvSdsfVaq6+sly/Ke7+Y1J8+60gPECyoLkCo2pp1bsrf7XmyleDN
dNmJQGdJK7cmiWV3lFd4c1AJdiiF7CvnFVBPTEu6+0IE/xmWvN4zQL6bmZJlgww3
QmKAvwQqtuo1GmdR8ISCk1ep40rn5LF8w+Zj2uuoMBD24T1OAcMeJmQEgIWBUFV9
1FnEa9XiPyRmGqkArdNr2jemghfhFLhF8wUyltEBaZZDrcaWkeL9rn799jcNjK78
B9ivsJoq2l3u5C0/vIFIFndaiUcKcATi3BKRqOqsS5uksYQQMFqzXzg9KF7kRven
eunr5496aN5rLZSnl+t8qpRBcmBXRKiTqHsnr+9R/T91X5sl8sKanGa01i/UFH4N
3t6J0cWqJnu6fiZ3Yd31YMBRf3w+oH9OeZ9kBMVxXid9az/YY/KhYYCpMGvyXYMC
8MSQIEhdsFzT8XgWw6AwnRYn1VM8JSnPhm6Qwk3CGyix6aCzFaH101iMb7C8iBJJ
xaBRiQEzSl/1YhEV6TZ2SG0e5WVM8DX4kNTfaJjK9FCgeacyKktuiq6AzQDdPKP+
CyKUQO/btIZyRA5D5iNo7k/5ADKEBT103kKpL682uWKb73KHUQHSV09y6ei8rVeW
QXpNk+ST05KhaUVzpU5O19x3S0z2tUpVYRGRnhep0Cvry+KTQwBHBVWlT0X04leA
lJhAfnhRRs/LXrWXA29CyBaL3jidUteIJPokSIAnj8yAfEmaoed7h36kBYnH8UDe
0CsprONjlYrTA2n8ypTOIM13xbEMgcu858JZUh0y6po/xeHNvU3l0in00I4e3VWi
tKcGz0U6F0o+d6ZuLE75QNcCZMgMBOIjz56zt2fyzc0kITktWMyEwr2u0BxY9EZ/
sICOXJ5Ea+A9I1p+NzBbCw6n3jT9OLnsPFXUroljHOalqU1g8dvtuUEXC5ur7WFV
jX0N4GmP2sGR3Xk9ENdTlcFqSy0Ce3GHVveJ2WJvk3aCC98f3JIqXnQ47MVruxJ1
cIZqZT05B+czUWoR4Lw6bDfymxg5C1j9IGZtOIGwpo3x7NdyzkYrNGmkEcZ0ovEU
lqn9i+M7klgIKWjd/a1dYd5I9R3lI8VR8VfYh7UMX6nNclFDQXhT4ERivc27Yah4
rsUiS4PM9JGlZ2ImH5sPvsm9hSsdlIwr78HZKqXDt1PzXke7uf2jzu+fxZQQ1gmA
wW+BFSH/KQe96q12+UNZhe0CRF1JgQUkEFmOV3giSmxQ07pnBGaIEAFR3QIN0glk
3LPxucKLBrT8X0aMLC6qOB7F3uLbLl/hAp9V0ncnNTtrjXpMPXYzdSYChiEOJa/b
uxj/BzvOZc32z9GJiUYu/GMTG2fLeSeM/vDGrka4ywtem1ct/iOK5QihtRMoeAOZ
loMwl25cUMPaBY2ofMVcdIfmhi5Pahy3Hfvhct7HOmy4DwvPCxsJcIIkOITK1sg4
JNMi0HUCbcCEucPVn8EZCluTrRijHRMFjG45lyxZsMucRnt1atmbK5pr2a+JQ3mu
rKROgGkFtm0WbnsMjGL2ueF37QLchibGLC2zMgH/OYr9Lwo0/tIn6Dx/oLBj2/Jx
pfORLDQKC67Ii3PHxlquT9c4S/unYbOtG+DUdXz+xya4KcXHQgBqhvO5ApbHInKy
xsircEuhr35GQ1AAMVMbupGG6tPubMJ/lbndla5ORer6lIx1VkjCQvftVSH8e4P0
y6vfWHHa+4z1YVL1UjMN3wJ6w5PbTBUVFXhLDnhQ53grpOalmymYtVa3ssCoUZu1
4ogsCvuOz3+Q3UnUfg8bPzLRJKNkFNHBrvXXdAtBUAxsF3pakP509YYEDyAubD/0
eZQpC6kVAhU9FnKh6IvkUCrje/9x2fPcLajNm8NSCdEP6Q/9YNbLqA4FHuSYpRvQ
Xeeym2dhEND8ZSKQIQJKccXUAwO1wHMPMQ/eXl6M8ZxVfe0qiFmzP+GVLAFdSelQ
7rP7457g3ypYQpJInQlXtmD25jamQWoLztIlccacBRw6NeBdFkm2OiBiLkI5v5CS
QnHU78nWJhsDfkHWc8xnXuWD0Jsp3eHdx2CiEDxOhB//358lFWXFclcIFU73nw0/
wFMaqZWjzUJSgoCynZ6jtJqmxPndismd3vkCGPslpVK0WnXrdee1spsQR+SP1oij
E6HCB4lax5gD7j3YotHURXR+RbrK2bNPd3Ig8/TCfgtPfa16dFfJwoNbgkz0s90t
cPSss/7JOR3fsK/She6iKGMLBAabo4jstMlMfEisbtbrGDCONSsGHzvHOFTRHzlE
loVrP2ApzmRhj9CgYdRGUG9Q/UNCwPH0coQk40DhaEjE1WOiOHWkikVxmGsi2JpN
JcWu5o8pVDdGM4GifQLwHy7P/sAqLpcjX0N/GvXpCXb8kdUyWfRvQEK5m5c79rUo
BTmXUrM1Dn8SEJtZfoWYXrq2Ze3FZT+LQwsMTHAvZ2B6plyo1cxQtVRI4NDfEC3n
CYAWTtphW3arIodbP9IIBWI0jXKz5lCUrvJRiS6NDzoHtT0msN1gAbwX7CTx3JBs
mM37wRkj0fjTh1mFsNAVS2kzuT+/43aGgWxtRZXVZOGZ7MDFeYW2hhDsTvVhCGOY
bLy/gcqFI+xO+e1Z6E+UVeIciXwhOtp8eVic03EQLXnJNo4XXG7+dnGdYXel6Fag
zRniOL4bm3aUAM2icxlAiZwrvsz15Gq7UZRtI/Ym6oKQcEWX6CSgwRMVMdJXrCgr
oHW/DIP8xqZEJzq83I1d9LbK4FpQXGTsWsDCv0UPUG+Ay43bM9KOwwRj+vW/4ul/
DUMqLXkV+JIHSs+iUrs3n6VA6pbeQG8qx61AdV8XSChBNrXoPJe6gpVNRsdsqitn
FeoxN1qvvxp+rNir7PiOVudyCMJTD30Sl+fxyxAvfGpFcFssHrEY0mlvYW7g+IT6
xzpRCoCjtjJ967pWOs3J8r/Y72wDlSo7lbivl/3qS3eAFsDN/bC79vXVAaj5pNkL
+RVICnVF4z2RftjvTlLRBJxa5y/ms50NpXJLtSPsjEdz40fLR3m6tgS+JdHbM/iu
aee+3MxS/WyHJike5/ACdxQCsjmhs7z4m4L5+u0hoPdv+5/jakwNnSU1pbk1IV9q
iuobHnq/YXoaafWx26GNbWbwS521DYFEU89rF1Ata71q6WjPQrgiXB4MTMFnpdFw
ME+c8F2l0yfe5fYBGOS8ENXFrInNQ9LYMGxigWEGyKi0Gex7rVi3XtsREOc7M4Ds
T6nbuBF6ouoDZR0Mtg7rVpYr4dWJx2HKZPaJ45gVcyb7241ShRecDV2Ld6uo5RKH
C8IceQ53RzGzR53+UMkdvcqYu0m8c23IglzS2vSD1kOAYtgjpJWKU+XrwECqQLKk
6gHVr06DDVYR2q6dRdBrsvTzMmcNZI2FJ1eMoe3YtXZAXYrNZGvoP8UkCfSC12EM
TNGPJsAY5zLlI6FwZNAS+Gu9/NT10Jz3ZjWniEP6HS4plHn3T1Ij+i/OAEhItDW3
H1wLZYu/8jY4yW3GdS9zvMHPQ57oD2FMPBOrIC/5+r5dBuyzv2Oh5pzBR82bp2Of
wUaO1f6bYVtNVxTQY2u3V+Okj9Vz+D8Uemao1oyzzKj7CZbIhZgEA6x5kPGYq6eL
oFDK/JA0HEnj/fYWjfjrkZUYcvkZvDhGUVnTaHa2fIfLdV+VkTjXyScFX2QDYpPI
khgFzpF+1qZbmtO3bd2Pmjy30smJFCGc9p5qpQetI9w28UX0w4TUrj9GHHn3fjiF
ph3wpXCmBWNL0XTcj9tJYl1ZYosadc4pjoYEpBjhOC9MY6+b/Zh0DkfQm0PVVXSb
1MTyXe6+pXQ/3skRZDbZo9c6EPkrlLYV9wAS/gcG/A3BBRDIK1ZslWcyVVsw0J4E
Pc77pdEalhGOm8k41c0k3yeFVAfQ2mG/wtVtbeTWBS1sRFlyRywqq8FBoaYVtywd
xbpq9DgOQUKmrghopiRHR/Kr+h754NilIjfuwsciWF2coKce8LaXs4cfBP7GhuND
QxFQPh9UzCXEIFcGpfUKqaZCjeUiRmgZZsNs29E9dr2zDsAf/LTFXjRqRoYcsjiu
vTUSWqnJV68J56avU9+Z5p+4SMFHcPXXcNIcGLX0Yn5UlEqUu44KmPtUUywGx8nQ
SY/Vyp5CVzlOB01JOgA4MWZJeChAvpXycgSwmAf3lH8mOClVcV6RDdZbENSW1Nnr
cnFjQ8++9FmxX8BZ5APeTYYAIq/7IVUd/gVgXh4A9dix+diip4mNVYpXcM3fIgSU
QypZfI281xvfN5XLjaVfN5clIdtlNYvsG04VxxO7P3Q06nStdsUQCFsy2F3KElxS
Q13UDADaLZKUgrk9stbohNEQrZO3PMu65CCMgP/1rHVS91Ve05thpWqs9A2ik+JE
dkhWhSqtg+Wb71KZdqmmoEZ/CcEw9xoQSk1LpPy2LLn1JaHuG718DEubEiq69qvG
gm3Ytm1W6PrGsPcVv0RaPl2kXZnVFQbGsxVLIrHRDC4xqQl6QrdvRnPBusQb9r1D
7mdAGt5lHzquP7WHotq6nEfa37moWE7LNxGcGgLtOv8tRQJx4GlXjMyXAHyI5RnH
fs2aVEXgT8iUUmbPWrvqNNKp6Hkn0ipm4Wc7Sb16Y9S6YPfo7al/ALQK31Zxxbnk
5VOvh7+N1Ec6KBCqsIzF3xGsQeGGPq4BTr0bcQl0rfdGtwdVoCpiUpOWGH8N1MZO
7afrdePBe5c/Qf58pf2oce+zkvnNX2Js1nSYqTOaNe5dJRq5B9kOxZaRVLV8HwmK
pXSChYEj0qowSs4gTBLukPpFMIxK+kRplUBUwduC0cNGdbSvw814ATsEbVBJSdDa
cvQVENwyLVEukn2l8Lr/vC+dTYe/fmthVYbXKElFJrszf5b0OGWoBd5YRQZpyTvn
HV3NJW8SAc2N5A67O90ofT6RYoOIP6i5ZoW9P1/Tz7TjVBtqTE5jkHEsSFwb8Ot+
KceLvo2GLJH+vET+QFytef2fcnapD4PUB5v1344Eia4umS4cYry2fNo1UlW+8N8B
mDslGAH1JOJ9DNQlR1aYogbXOA+r8Uh67e9VqovunW2nM/U3blSMDL7RACNZnne8
cbMx28WlU0Qha/sZZ03+doZqS30nNRKp435wFAxuJbQNLMMtbF1ofrFw3vPqNuX7
cV4isDNqR/7Yi35tzrN4LG7aij8FLeeCR0InwhMJaOSm4quPAepu/03lukuGmH3C
yZosqnvaBmAz6q8Cz+s0gCEb9hZeO94wF5Ez1L9NPyKMsCm5ZRyYwOKJbOlPRBL7
Htc5Pe9UDlxVTIZRQZCzhm0F3nS9J9TEd03bt93Jauyc0hYTk6DnDPdDXX7eRIyK
GMxOvl1cI3sMTj2NrG/DvP/WXlpn3Aoj7KvKBbDaMY47BZOQ/iRJ8d1YQBVn5r9J
V9A2w5rORbMIULtluPNriQATsO24gObvMrWQLrVcJUiK8L7X6h5CThyVXPDJaKmD
8yTDKZCWag8yQ3NxLfp9aRrEPRm/wpuVK9TgeHVNqXcDK1KKZ6g3GYzuNFrke0+l
i5seqMDNv/NcAH9l+q/BT7NihIoyYZTlfLpj+xnhROOjCjC4N3JnOvL8HR0jN3Ao
flbRlyCB/8TSlB4p5MqmoWyq4WZfMeWx4cyElJfQwGoFEHkssRZJhYy2rf0BfcgI
XTYdyn4jESXG2ougYN70iNWY81che2tS3q/Bhp9/lcBByr9RW8B+LJ1076jYDAPn
/JQbdHwtXhrF8gZYJgLHVl6wWfR0uOySOljdW+8w6eYOWmqGJ+DAAQJ5pV33/1dM
9f5RpW0cy6I4Ky6AtcTH+CHlnjUlvbRuYGz47eznrVtqdg9VD6CdtMFyABOqC40W
NhsuO73WhB55iytTVCppvZlVzHdl0UKj4/7pEcmw05j0JpSsbV3lwRGNRcuzSU/4
s2W52BnUMTlP5CTpvC+IAOF7kbrXUS8U5q1xAgRQ+2vtcqVrBS4dCmJhPiKf+fmf
aE+LYYDUj6rH56FeS+OuFCCy6iRtl/5Vd3853atZlBcrW6I4Qw/vhL6gaaGg7u2Z
g7mtQdsGMkbtBK5Ui3aOO66nmQVd8Ska+UiKZSsnNreQdnYEsqGFoI3duK8UHni0
qg81VfLyCHxjV9I5boIgfD1juBPT5+9oWUscfjTmTTv9qG4marFNwhzeSv5LgN7p
ahEZiXL5g+ghYClsIxqvNGsJzc2HUAKYNkGk6Y3PFS3CPQlwIgdmfcB7UG6lIzFk
ElZvuCJq6R0aYIfEUy/IXb+2E+Mnmq/KjZIUy5ONriEcmaIb5r+0T+c3xAVI16nO
10eE+WZPycUE1b+0MruG23iAq+a4WQne26mk/LWPKrgKjr3HUjv+cpbyDZZ9GoU7
5cnpneo2bSBHE83jYgOXwFDExHa+AQkvq4SieiyhfuO09q19bxsYgtZpMiBnKmIH
c1gZVr1qJDCtAUbqwnEhIkNGpQiq3NLVV/DPk3TlyuorgTzW8QD8QUzF2apYkpcu
WD7RZ02dcOCt4UIy+s00n1MhQDNSrAP3ZgC30x6IDKEN50PNsS8YlmUe3UeglsCO
IaD7k/Yl/tWaiJCTyiUTsxeUl4+N8L1I2Zi819vpndVLC20sKHoE1AsIhKHOE+xv
DvNyJGwqVtbrIcjywZSqiFhd3bo4Owk8MfQkWAy5yS3NpY8VaZKDtN6cfcGBVm+L
3K5Ac4pRoZ54cMY+66RHksOwM1B+fr+EmL9bn1uoWGgvL077JEBIQDJ5SSkR3627
lxb9qaAJvF4don/SGN/fi8ROZrVJy7vgE65jaVNfAuypiTJLM57VcaoylfJ12BIa
cDdsvyvIuUu1pMP2okF3pAPNHXMC0C1irPo4KSuaagdeKXsEfBnLz1kreTkfvHAJ
y6TMb1CtGgPw7Uh6F51mliIavsdXE8gY+fwqDyplMHOBn6AtQamOnHWuuu6yrqRL
eABAK+XWxDzzw7TkP2kEykWnEOnAt9f5fm0iyDv7/AUFQt8Q0bHmQLq5O0YI/bWi
y1IdI3izx2LQ05hJUca8yWvidEUeyT5CLcvYsxGFmWPik8vCcr+lzVCXbolb0pMg
5HoeTBxKqc2+qmH1nROto2Iakh68Aq5BfO6m5ZOsx21A66WX9DR16wbSGdiKS8x4
Xp3n1jUnmiteFKdbHJ5fp8lxcZ4x9vc5GmmlJkvEkkEOIrIMvdC83YQvvUajwn4f
C8TwreZOibxl8s/n/ap6KZ7JXZUHuIPwM40BnktqgdaAGF0XfL8eprAgd9HhymsE
mXCRAfE/GRnLelykWvjQod7DtWQFCB47RkUMZenvJNIz4TqnvEgn7kYGGmJss0v2
ZaBjar6AUnrlSlvgno8hjZ7dNoOONzUo2KZ7J42H+Z0klQikTvdXMkbP6h7aI44K
hUbFDxo70kszvlM/QCyu4ralrJrUGJ1YKQ8FMuoEo50FBOvxV5ffzBLrJmcABhXf
1zp7NmZ3UM3xduTInC8/zVjmP/Eh51zuz6tkoxhgiKd11FHT8D/gUhGoKuIzSDFG
2Xa2/O56BY9RazGnK/9HROiS2Ya8fyxUHHeRaH0yKcMcFgKWGEcG1hnISBJ/bvd5
MRhpdimwmfsi4Pp0I6Z8u8RNUCqrdf+L71kVpFoLjHmmgAl+Azw7y5EdM8pA7q0n
QY0u1cA2ksZ6GsZq+gA7g2oKsUf3Pafk+bBGP7i5IuYbm5vjGnTEVRKiSK3FNPq5
KrK8iqvgizw3/DEq0BHEV08Rv8fpEMDXIIc6Aw2wU/0eeXOqFiL06phiqeLP6g6W
1ST1wPGFT414oT3ljx0MfnR3GhEQpx9q5LM29Jj/5+oT+DqUOWBC2DQHzpY3eN4l
WkQ4k9KRkp/9SusLQn/HC63xuUsH3WiEbVBuSIxZxKJP6fKH7jpJMt0HJvS0j312
t1jXQ6QDEVIl68WogeSyL5thMefGDETTUkj1y85bncfZuxJ5C0oealJ+HP76etQM
E07VODq1sQR7vFEtySalTBDz4RNza1R0uyt7fNkKZZK1BqyJBfhM6mK0Xk/z6M46
TDjDZLl9uYmVNB80TJ8MA/jyzgrio8kYHRBGgEyMSmyGhQ5m9ZJS/sVRostxqe03
G5zj2wcB4A00+7hMIhxCeOMTtq0xPdOhlnUWymzfdf2XIBw+y1rZLCEyQ+iyhzmp
fRUkEpkjjhrfQS8MPme1CvtaOsef0ghVqJL2hk0y9WNWN6RW6cs51gIZm9BbzOPX
6dNhJ3v2Znj45GfzJBAIYXnObcRtyu3jRXO2Stjta8Cd6DbL9RcLYdeqYdBzRRBi
k5bSNE9CHwfGGMre2bOGhHVBSO3NxPKT4js7zBC6IRn01TWnl5YZWGkHr+1IqfvF
ErvCkwrVtsIg2UfS2aV1SvVrjWMIj9sapY7/Jnb5q+qPS5TX3pi3MwNFdkWTPbXK
TibkMIMVqj30Wg2tgemyz6xDDYr1zt5kCJDxEqV2Ue9F6rDg0cpA66MbudJyU7eO
Cqtzv4JM/OQw9rWkUax9371F4XGcJpV++HqVgtPN1ipoKcgwP6oW0ys9AYDgQZFu
3RDutacfPpPcvO1sdHrv3mWUAs0fhn2lowaaySIcvnS7yJvUPfMAP8O6k4AKGeVV
2ID2PZ1rnGOuWyWR+57MmP/NvD3oDnrz9xQuhr41etCR2OmmWDhGYGsZovngdjpf
z0c+ksMuxo5qJQTLYvDoxjGVuzSq0KaR1XR74+Qil3MnDiWg5h5vCXsXGqlHZS6Y
3TxZMxWApkj02HBUnwTSBaDY+7spwBo42wXPH7o7/vA0aLysaW1pLr2zc1MGS8b7
oojjtS+pg37QXa8bV9O0qcY2R2jadkIP8eVBAn4lD2yR4b5pheQGksfTVDJwHq4g
ugPMICcrxTkji2cqQVOqdyFGr4xZPjW+w4wt9C4/eLVfITpkA4Ze/pEnq1JHG1tX
dwNlpZ2UfhL6rUwBTgrtD+uoy5DiHHZx1gsGYnPOP8icIWIgbVc6q893J1NE2cLV
wT1MPQ1VbFkoQBpfzg4agsv68FqYlfUWG8gq1YHAJ4rzcwETzDneO7HVr36DMj0m
pIqH8N1+J/NDPhlcPxy2gxYPiITq/tvhWnIZ/UEoEmI1wv+2cuiNrvmGZ7VYdIYV
oEKxoTuibRtbQd3OCSGpcCTedFFenG+dqvTOMYZL8YgnRtd3E6EuBStBq+DKpoEM
RuBscePlAOhDY0SuJ3o8vl6MYN5hUYr2gMbtj9burZQlJRNP+CO/TRo3aqcew12Y
9BBrboMtUoH9bED3+XrXVjcQSmjE2JpYDPo0m3iCI4NrYXECb+DhTh5Lg7uT+nna
cIP0tc9BVV6meTLTrxauCWwKcB8z5PjvLzPnP9UaeLpiUXXWyeVKU9ZPd6sDvFvD
wvY/615slL5tAnaJf11qSciWQ3/snLRu9xvFKVFzdP+TymNF0mHCG7PnUZz6a2xj
VxkUQ4YdEMW0xmZiqIgvHrEIaJ8p/ccgLa6bnZK/GdJdkIiBZa4AjueinjAA1IPa
6z+KbxGh9deHk82WoyaA4/mapQUxj+zcrV7mBoIGtBhI/JVAahiTzTAFkosQNvdT
8Uu+Y5rilUCrOnsg/8WOtn8Y0nFpjorY+EBd8cFy/wfF/Z+R9Uit6pV5YUkRnEfo
ykybHYe2dvYMn1tp5aosvYGpYqS4jcjpsU5qjaL0hMvYGAVeaNpyl/ZQj/XeQiVE
yglz5Z8jZtNi6ILED39eq7iVtknEbHjzqOBE+y5PBKnw++4lQAks9/U5LkWseAsT
iOdkuayFgbfA4W6BM90CVjuutLTv7F/sh1rz/zoWeT+Mj2qekq85hStP/pMecXEo
xXSoznWWQTk04AVdYCX9XlqikywnBtzKHhfqBRpChiz2+p6NY8u3DIV6PGayo3hu
Ft4lhcoQebphSdA+7I7G1GQaCmhrNvOpxgGLGvxRSlvNV/yV/a7A1nc3MCqNPMaf
h/yu/46i3owt7ymvOxk/4j5dOfYBcmF/Br2rdr5Y/J+Fbmn+x+cSkEEU/lDhI+er
MKjpplgc30KGgFDwczhQwAEsUq+vJYzIOZdT6F+b3eLN2LmeKzW9JhiYMblCRS10
TqX5uARysZTfol1QJJdyw6fQ5mfwjBKN1uOCUGgzWIWBZuAZUWwYMc6ob8QisW8K
C14c6VjGQ4bu5SfYoVms0yISiyHn25RgaM116ymKT7kbX3QdzpkP3K9alybbL46p
jyv7a+QTz/W8PAufKp4JqcjczTS0Se9YFGtZExCgsSS+9oh5fBMabdcDeR2iL7aE
p0YhkH42oO84YJ0YJ/5Tqiskpm4lj/MudjD/yOrODO3NhJ4nBMX1TAFGUPnsImW6
pHBEiljel8Yjs0gH1msDNk1ldMYiLkNsp/tDRZr42KeJOQGPL1/UYd5/7LZKP9SX
udqjxQWY/bAcaOwHSKaw9F9K1Rh/Z5sMad554ltpptVp2wheXUIfWtH5UCnQ8QxN
ZW+fUKQ/Evhhh3shIlOkGBnSZ26jRzQtshsJImRydPZ3hJEXknOVyVzlYtEOOpnt
pPE76DjxcBvoTsDNrnzSOygxl+YzmYUiyIolpw9OS8o7J4rJJHJ3zo5Kz3B4vGg6
zNP/g9CrZx8fOJ0K7dN3hI2quJCta+hMm7i5BRdLqSZTvm/nW64RASiP8UZY2sY/
87OC8XVInrmvI4RacrmqzW8KvVqitdOh1miFVYv83mi8TqJY6JP7x9cyecgYJXXw
dlYXLTJRG/LOu2JXBR2G5yGK6Xh4LJF9h+gixdb9O5yli5Rs83djIxdJFdm2/dSS
MZAr7QzzhM1yFr3A2iJYcLqq2oqSvWPts7bQGbjBQmlPLGGmV5mzZQiJEhZamZZM
yDTjR81zILwy9kVDWtISCZ3/yQchZIKbmJp+TFErDWN4mDlEdSGvI+t+nqpzqxk9
LhM62KJavCKb8w5mpK5YTK+6+9uAEXXFzdRJnOgQQIKVOTzlqj1GrDXkFTiehsrV
Z0n1O0Fw5eDCCfgaMLVNiOLaDz3ji2i0zFwRLqXpwoz1cFVS5r/J0Sf/RvWNn3CL
h6PzDIbuZRBl0ZO6H2v+2Bjw+kNml9ftYUr7e9qiMAD76UbbF78oRZmIxe7N88DH
bIRN95WdukcvJGyW2DQzZ++6fB/0r1KLAdn+t3YUBy4rT6mvrspKw0xlIoRqED63
SeVX0eu9daDdR40cSPmN4xSeadzN20gx3FoqMCIJ/P4u4tMvmkrubxoywn04bWbW
4ztjCRiJ375hJSMGRUHrmp03W/KaBsQKxB2sGN2UHzmBYb6GHDK4ij/lHqGvWyxR
8cKgzvOjS6oxvk+sAhgmmU+g/us9DKnT2CmL39HlliRD38Lj/yhnnDFJRQ3T2NGl
inQrgc88ZVuiU/AlChJw2RFp+19j7VHhQWJ3c2DK48GqlFC+GAHOVLWCrCV5WoUN
6TPprCOLydBr9HcISJ98oi5pDu92rFb2lAop6bHluGBOexlH2bY6Lw9kUd/t+zgr
bm6tQgxFEbF0YsmwulfaDFMu5rcWgV3FsPN6zksbh0wz2u5rfH7nv7N3YEAfHS/9
28v+0pL5DXYWXsE13y4V2RMBfgnq/8sXf+Qaql+V5fKNm3lsUuzcDFYduXKVo4Xf
tBz/iyY9MkEyXmysJd8WVrTiu2EQB2KRNF+lL852u9NklaOBZ+cwf2SK3loHq09r
T6sic9P3f+Voie0n/OC4iE00DYPvEmERs1j0Tzb3AKrtYBhQ0btIVt9usKRcbAnN
HpZHzVxG9OqTpbNn1u/tAcf8PCAg9rhjVoo+d0T2OtNrJ0ASYVpGjZNlK2ooXqOT
I8ysbGH2Bg5jzUs4JspwXD3OASyWoHGE4QiHncIvMm2UuHXDK6LeszoENHh8KZ6V
A5e3JGpq4U/YgUO4dvYecUUQtlTANvZUMvA+MMcdfsCSYEfjDVao/RsZMdgbPmCn
eYVJEEJsZKSGVIH18GL+KyYgDvnwMeUewv95WOv2R0gQwGFA/0ipdaSz9eL6Xemm
c3XVWFauK4QjKv1PESWFU2cbDLA6nyAQsXj6xbFmRSXzaI3hqf4KH1D8m6BFYvqB
RS6R7We2khgrosJnPhZ8lrjFvuqRxvD/YHL/edaXOuTjy7umqVlTJPC886o54IiV
76sOlNEg7F2MS8r1I7pRx58y2Ga09QAwu15AZVkS5oRGSZgT1AsnW4Bhkie9XgyQ
JFaqwWyaiN88k4vDJQAbVSDUpIdjXaspKrlgPJCTiCqsBvty5YTOCHEqYa/HJt0i
nFdRf9kRjKsGPBL5JeMBc311rM7oxlLcvtbx/anQhT7eV7/l4sWe8J7YNDXQtIU1
9qBmgNB96roREwDfO+6D8JaeD0YTzjh1wBhwo9v10UdKd07x6y1CUEKiOA06BhLp
wGUQqYIblfjR8Y5Og7HvuEk4LYbRi8lMtip9O2XWG3w5+M8o9VcR5B6z3HSAIrnF
2xPZe+nOh+mc2FWD3y0eRjO8u+46D0HA0kVmnH0r0yyl2PzXskwQkU471837XoiN
ggUdeUg4874uUxC4nC2vOZ9AP/QCjRdx8Rk/q5/bb5BI59CA/DWICkXJx9/1risT
RMq57XkyDRqGLvLhF7zySTAGEnv2K9+0HYp1QLeoBU8XOKmIcXJaKbA6qbtU7pXr
mPJ5CJ33yMmSolCEaaMUQ5FbLiT9uHq45Ch7msm5Sf+Zr7PicVCczb0kZId+zlwC
3Ba3IhZjocWmje6EWF8INGPJrpHmB1RvdZaSTfWDrnB6fgxyVZeFMEVaCq5nbV1f
CnxaCmqEE5lKkzoUQNB16GohF8hkUekdy7AXqt0tI17p7NJGDjl7a2AFF+vhFkoY
pkYOmPwy5VT6+a7Aopf/mkTVGcNpil4RRX+gYs3z7rvhBJylK2nGxcUKT7Bj2jLO
pKXhltIToLlhj975YHBht3gMTIKnrcvQPCCfdkCqCbG96Csb6mbgeIhy4ca+gANo
thmT6Z+srsKt5oVO4BKzm+gcGd62PnbGXFzYJmkkmVZJl0kA8x0hxu4XrEAPbDdS
RjeDG5MvkOaPpeuRva47OPdlcYQdldLFzfZ3ShRhvV99HrHzglwZ/SGUHVKc3sT3
8fi3O+7MqvZadszPxrzVh7zDl6kthK1RN5rjw7eY2P0Eo4URvf6O+8Q4Mx9vCDkR
reE1k0+40WQY8ywl+k0R8od5Zl1F7uL4OkZYK7HOrw5w2FKVnUWYWBYxFGUcpM+U
U0ciJXXXthc0B1Mv2txF0ocFFfU8ao19BbuuQEkFoNdBbxvkgql5jqrtvYuzeSiI
sTXZsJ9A7PgM65DWBRLNsjyPQ4gbu4ZhrABFaGDs6y9wPMF6u3RcllDJw5tl2O9i
CTOJiWl0GYxQ/G0GNGUp4RWI1XzN1yKSkxHW3jFxpdVj/XcCMc0dvpRVpIKX9AbG
3unXgw2/1DFEBtaWT9wg2NKf3kAkPJbESq0GWI3abTEAeJf55LP512RXnRj2EYw7
UOm5DcqMm6liLQRQQTY1ca3S79TY6ioB/AO0UbyEFR/Oo8UEhW78CyA3RetkbuNS
5blaLJLGgXhDS04y1g1o+J6l2eQGsjl4QJmB+BQSYWix+PLuo26Y4yHuIoLFXWDO
7qaj+iqG6ttGLvZRPVtRMmU3WrdD2yoWXNb3zoeTQfWtTOkyr8auE7Egt5hvI0pK
B495azeRBYV/Bx/dlB1JucMFG7ER7fjHM5qwqEW1SPUa1rauZBb5UKOZgYgCLBD3
onTvFRQhWvZMFVSuXUUKdEW3Ammmt50P4o1YdZrRnvIB/Z5v7RCMGg3/AtiD6rjW
HMX13gNMpkQYbLq7f0YPO3lDC+UhF9BX/98giRhAC9wuLGB6NZdoEGddQIWdpAIU
C61Fw6zgkNBNt1sNTlTVwcx1LapJw1JJkIhmZbacQVnqDyBuML+sGwKOwBPxTbsT
qglqkIsSgopjbOLhH+0jea0dvGUSAWHAqLRi0GVGsIXftgjHLA6G67je0DZ89pIG
YKh9tEqpX46z6XKMNG6uABJdH8F7hfL7+PpncIoB0DC5V/MJAhLSEGpy16lE4mSu
SQaZOBHHsZgMcDPGdgsZTWplKUILDcb/9e1r1Qj2u5Yg3yRySxc4WYJ3E6dQIHUk
ZaBfhmA9scaz0uf6IwC2eoGPA6eaKKsN2ZE3DMSgh9AE4MG3tGoIGCphI0xP5/Mm
1YLwWdN7qrNa9nist29ISYVtrj4JD3/wBAqKcX3oQ7lUniG9Cha926Y1ASdFSnst
SFpF16LnGvsCa3QoQwCL56MGpWnFs0ZBs4P/n/qZgEfqaVksFKVynjuS57jdrd0V
BSXP8dZ/vrPBolZObEhbyIEbI+qHnb6RHE8OnXSuILMXKkrKUWayqXDi3St3NoW6
46uIpcufYsu24TSs1KIceehbaJwADzrCZowT9yuao7uAV7c7JrtG9LZlYwrrpWKG
hXhZQfR54WwlneENWlblptCWl+KarDBIFxaNQVAqdXM4pCNXMMZUu1yj1moruZVr
p9Jl71F0qMrQH3Hu87AeM+18akKWS6Za2k0iu5iNR2UmD6Za9VM6OdpL7tv7vMhX
kk2CyrDfXOkk2uTXDXcJStN3+m+M4iSP32Q66meQxEndzhAQ/KZVlk4z+/rUwlKb
gVo8IAbTALOmJQ635UWEi4Uxwj6D4oQvEFlFJvC/yUXk+4sNHKLyrjVKnENS2qK8
DUWmMs6gOO9u+h/f74LYD5lg+42lYSHMDjwqEzkJmN/mE90tyTbpb//w8bc+9IfP
Blc6PlYIL9nDCrQRy3g3JBbOzfmSSV7Sqm3X+sdbpGfHcbQ/jGtfKUbDYe5rnTkT
TyxtSUsSNHozr+WiaAXsy7WuXa1cxQb+UKKnmSwoBIFqvMEw3uAk6LVyLnGExmx+
G8Df9Nw5r5Dy0SFtIhR3U///0thY8RfCQH98xRQB5Ofck3ObKQB2m6ZVYi+TylTj
CUG/uArehA/RVjV2rxRqN7NWDaskKyQu2ULcHsAelHa+vFEt450B9sFVTBmVyl0K
H3lklQIYVLfDWoMs5R22Zi6xGCvv35eMBSNlbtzHVKfsKFl0XdLcDmCA7B3hZ8Os
Qi6ge5dn/YVQ6+WVdQkk4pSdPDQhDFigY/0uBTcuqceC1YRlev9jMiNT5FLIC1Gy
0l+hSdrzoFyIXAj8lAQTLQ4P5m/faqzzIORIY4fHqlKQSnfWcmss43jUmIxqrjrt
fJN74fQpRGw7DBapfwF24ysEiAZsMlU9oXzzJNkZxAJOBAuvXFy+Ui6aEMnqVRaX
y4sJVklCt86cyRdvQwouXfkiGb/xzMHiU7kSDH7bs7FpmxC0T9hq0M3LmawOWnpp
/dcts9L14+QONsp5S/FVfF6Bmi4hIVwJhX0nZWQ2lq+UIT5x6zW6N26Ob192dbvc
r+QpSASXZbuy3/rTYrIbJKPtUJuEhc0LA+Cg2blFeepNniT9R1Jj4NLVg3tj5K8u
b3l0Iq6KhoT2ULMFIzWIap7ceWkU/DG/l0w97CzSkTBo0sVAYKR0v9I/oEpxe7ep
VC4c/+ytmkBHY0RfYufM4gWv3kGTA0syEkH+3+fgV89JXm69Zu2+8zdLfPyRpeGm
0CXvDu9yIXAFSMVFWoG6tS/ANMlXIpBRGaTmwX8xkJKV5rVDnL9EmFmodQOEsobw
RGHDajOYef1MO9OdAZvQoAfnDwsx9IOlwrYTJzGozPXV8vHdyKo67QufJeLYWZUB
C9HkdszLKSCAMhRTSLTA9L6rzvTCRPhW4I9ynzj7DBVGlcrmdj2ESs/t/6IDNuuu
Q2eT0abjEYkV8eYzcz8MkrDT8zvntk6AOS3caBSUfaqVzjI1Qx6/qrMVE1tr8dDk
DZK8/mL//1pI/KhKER+Bcq0nby6GwX/xon7ozdHSpG5ZMnHfsISsSPXWxwg9H3Dj
Kp8gUSmQpdT1Yu2fNve17ISq5ft/f9V01JPj/yttjDDKVqedvyxfjTHD+XymXsrW
zPYPqqt3FeLfbJA/3OnVFwtAPCMlGA24UrGryePzMHAXVMlUAzx5vFnXyWyORK5D
67D0refPTcRlsMQRNYpCv6FT9XZxxd7BCPxbI+WvvKur2QZ/6Ltd0uaiOMl35c5Y
Uemn6LqobCxUvMbb/f/ZOTPGzqAC8DqbtQCxei/CxPVYbAnVkQUKVp3wnNrHh/DL
pOamq8Uk4hF+mKAEqVuqm37RZ9vm1FBUBOWCvocP3+8TfqrKCMPNZAL4We7LZx6S
ket8c6QozGlxK9OWKUWJE6+fdhoN9z/HAs7x7oIoV+EyFn2HdqVAoZp5bsS1s/tF
liBAbd5128mJaZWDyhuMg7A1xTkBppLXQnxaW5ydPVL3OqaqwY1edat5eChAMxJc
G3DMLHfTKAS8pXkonAVJhwmhLlyrBvVpC2wku3eBXfn91uc7ncXcFynlqkWRjKje
+OfGcPZsh57sC4+HdjrL/U7ik7H0+aHutQkiHbLTarTEdyr6MIpUhf5V0b2ZoolZ
PIhUJ45U754/OVXEIL3jH4wFJxuoQYDHr2LtPVILA8KkmFP3OOJqr5LY2PjK7GrB
QpquuPMkSPeT6aY7SwhFdE06s3qdCxI0/ZtA3ZoTeQhOETSXeNck0yWFXJZETiTr
sHXTMRSRumqcbCQ21ozf0PabmTI5gz08jWel7jlCXwZhDmm1SEUFyqFQvtrf5EaZ
RojsuwvRzXyqfmnchrj4TtP4QeW5jJ9nYnnj5j4rn6ESmLfLBvzZXyjECPp3gi06
abhd4PLCttgduYtX8P5wsWyAw1szfFVZb4gU/FVdg687CaFtQqL5PqtEPtGp0iLz
CTti8Fz9P/AdSv9ZNVnjkXgWpCZU0W03vjJouTsf9m04OTdrxnUuAIXNdTghNvZv
6DCHDx5PGE7YRh70rqjdonllpxlTs7+C4F7eIBhpsSmGavedqeTRuKyXQ9h3mi23
haLqFsdz2XJu/LNhfErqnAEMEOozk4PEPzz1ZP8rhTN+IIaVY/bfLwhK94pGu6Kb
UJeYwFEeN5Moux+/ETv+hIgC2J0UMy4w8E5AUydy8fsJ+odame60bUuwMT0Z1JO2
1G4xKpkdmqOX4euNz9CorpKCvfGKy7tTKs1sHIIaTfDJOhBNz0Wq1iLiy6S9t9OC
1kdRHVIUskV50DO/7rJspSPAQrjHYHVgCQK1vcR8nDENAG+q1Mlbus+pirXOmpBI
5prLehqaVmWP7SpUBVgOXe5bhKxC0ffmIOoSYf4jpuBsF/xxUhiMKWcQY1HpBKBj
26yK4rAiq1kwgwgct9OJ+vQgtL5XJnHTbHbhMi6UOIQr0oPDnvkoxlsY/2w4e8ZP
8vO33el4Df7DvlfJcjvIEl7bUtBHZLR7usj1581M2ek5WCAaVHLm0zoEGH7x4SVl
DfV/RNzBq+4iOd/eDB1UIMlV0ARGSVkyU2DPMlkDTaOhq1Y9PNlHtQnStIHN+la4
eMDaj0v0LC0S+u6f136OmMw1JRMe5SQuQxFQB/88ts6RLET/moy9lY7Uzl3oKn/9
7JYgEfGxSkh0/fD1PJwXV3bcxuzVCq+dFYYamAp9IcGISi43DHBAl+5WukhjHCKx
sxEDo5PWpF0R6lgZPjGUBIm25xmQ8chkeYBnAN8Sxdntldoey+srf3Hl6t6PRNf8
VVBW/NvwzkLybgKN+dNcRd85CAiwo+U7WZWhE7rCkdkcYUpd2I6WJImqBEKAwd5R
fEScApdKnKVG88K7+IHOSHh38JLTAdnL04xEiMb2cg6iH89z8BkwEQDSIzHV7qdI
X7j1xHcYtmuxWxzf5JcZ6QGZ/7RvZPAeZTdLZxvzMyD7TxQQMB7pQFEEOLjPSwf8
tkuLjm4McEsz5WUpM52cxkWP2RcmEi+izykQLVdFeQ6pjOGZ/SEH9AmQH6Q8ISsg
IDxLAVAyjoZsS5w648S1kbuV6Ynw15zCCXcTIVpaYjF8aVIkhHl13mQKgV4MQL1J
yuaN+i/w98LSuWCrOsXHBtIYaVJuzDTl1hHbiyqSVZ4upCgd3QjvSJ14CWo9qtQz
QtqcfRydi5Ib1YGeTu6NTE4iJRCqM7YtzuzHjT4YnlErh9utLdVC3qGPbBXzmHJ+
Esd7VcISjInN9/HIlZrk5eSkH+ai3u7kovpAl2p4poGYYhf+HMAwdBbU61EYiNCa
Azo7Fv3gCxeJyXnBL2JtBrozer3TbvIVWDA5YsqZkUNv75UId91YNgGWX+0HHe8B
Cf8DiCraGwoOuM8fOMBs2G7rWy683uDZ/LF8DyjrFwDvNVfph3+ojAbj/xb1tzhv
vc2pcOZRbCytVAtMZP++mtLk4LPx2dBKLWKP7SaoKZ9b5QvBRCyquaugfExCHBNm
VxY+r/hHEZNnf3rM4HtqJTU4iAe+TME1Y6eh3IZM+aKUOF8LhhXhRgvA4HP1k+e/
O0Do/B1KI9ws3n8vFYV9hJH8SM/Ae5C8VTtGSd2IOFBKxE3uAFsivIgrNr+t65kx
0ozpSXGS0L0T3w+D1eFw1hlMesVrYT6B/DppY5o6pvIRFikgpUxzeisdH4sBP9lt
HPQkKvGxYz9iX1sbizRU4eSF1MrQpN0d5AWPoalA3jER7fctncG9r3S+4+NwU8mD
cRoOib+95BlJ1+UDk+GUMQ8p+JqTKfxeD9Oq6jzh/yQrV53i1uN0mXXwpTTZrMFJ
7BEmdWyvgTIm3p6mJjTF3Hdf+FN5d9iWnkof9uYxMBpGZKjJLtyjScDywJqt5OfE
Hk5FVzhc4HI4JTembIgUXkryHI/Bl2YNtfEAK07tdruQRKcWav8xa5spUzMPY8ck
dm5UeGVGnHX52MSc+VgLRamDJN3XofrpMcftc8hdyGHlIL6JpGlr4s+hPpJELwV7
PfjsrdnRqXxDGTfeoa4bWeHdcEi59txDLBDCur3JCtTjXLtu6wc9ZvXNXC/L5efH
JvvzL4+68VQXd8wMR4s2cv2d4jfzvKrTmwykZ0JIBm3gKYOrZMRoTxpzCb/NO6xz
ZQ8J2GxqB4/CkvKchYtR2Y5kAnFbacgf1urk/hJigjjmVb6xmj7k5vriOZaxlpZk
jICClZP1njYN971e9P8KMEh6V/qmpk6N64i7hgjNoGRDLCSN0aB6emWyjdb7g1XY
y6gYmXSsY9O/md+aOAkxkFOGii068zGQknEJWdagicke+JFKf7L4eusUbV+Vv9Y5
X6PuAPuPSaJVRvJT8gtVmtEK9EeUoDGnaTPdSFjBSzuH6QvPVf8I0PDGYgIevXsj
wnZrORbwEE2FIYS7HALpgiYYc+EonjSw06k1HgRYFLe0zRfYeHny8vEsyJkq2Tkm
eso2u8QALx0eRVNNL8WIuKhAds9FYk7mALDm44ohlF3pRFKCtQMzsq+h2jh2DrRs
OSkHTeMSnxvsMwh53Zu94y+2C6CbbDl/THNXkR0TTTwoEUu1qlJ7e3qLlI3OpWkX
ZvR8mQm3pVMEKPF5U4RY3Pj9t6F5KAkX/pxOaVUs7yei1yma/8CfaVb34Rkbolve
4OqGkJ6rmc9FWDumy349RSeVl4RjVVOcx4OxGjirLyA+XcNlrE756nfEgSvRlhRj
smle06M4CVg7kgGUw03BI7M3haMpBKFx3EfMOOTU5v+O5Xnyv8q63dsaS27JUkRu
bSEmG75XSF0N0WSurAx7yup/cVBIGYOw9Bj32SJ+eCsQFsInzmhP+5g/YmywxjQS
gWHEVq+X5Fpl1h9VszKAqfnwP0DgZ7V8bKM5iXQ3NpdQWLC5TUnteGFN4bYAJaMs
vfCPeos2jVnIofqtAm8kjDK0vrpPXFJEN8f0a/bCs7Vy+4puJwXz0EaQtsgx+TkT
fouyNGF1pD+GvHInSX724upNIWZn655kqZWQlWgbYTwsLC7lOWwqucz8wN2fxh3a
PfDh0sT0Yspd7AbhOVxd8AFHHJtYDgIO1W26gbp41LED3lhe4p4WOoFeW3+ZWi23
AUTjceay94S9yl3Z6kgTGx7f1RH3jJtxiFy93PHcZc686lbw/AMDZqcnc4WLk5jG
u1hNVHL1ZZMPlAXJn9vrh0g72vHqnZqJFCrkbEubuvLtPu3ukxGJeDXemxoNxFd0
Jjk+N6qpDeEbdiSoPKllHvVizGckr8/7RNq5Fpdq2b2aq9Ge7dSt68HLn6M/WjDm
Ya2O2v0e51yumpTf8/4z1EwVCfIvuhKbX4QLPwb0TmxkJ5TTtRaTZY5zNpjEUZIS
NecbR4C2nw25INBTx+3duGcSQimuvIgNGD3663pmmeAqDU+X4wLaHSWknPljd4w6
LO9lpgADA1liVOpCdajFJOJ0dq8GePELhVUAJ+W+WMnfGCENSmWi37NcJIPOc+wC
CF6oNzqClUXd9gqtMyyLejPSDgSZuCMueiP6pQo3J92wAIzzU7FAa7ziVCsp0emb
Sg+1cg0KQS60A7dOBa4J6/bGHcBvnOKI5bYq8R1AOQrTANVAW176+qhWHk+yoFaZ
s9mlA71KgcuJJu14/P8mg5bChDrqsC94gCwOYry/3/zwsIpYiHRT/qZ2ZdlByifA
0+ERFYKANAMoLqhuc4+V/xgWkOo7gJA86bG1aikeeqJOn+uBpJsCHR7bxKDA9W3U
iIpwdEvMuqBguh3XOs2m2NXDYOG3m85BDfXvV8g2UqZ4uAhyWGml81MG0WMQdCqe
ZoQCFz5zfsB5I6xPNe3zopPHhH2ZmPI7oJpmpDZuJgu23K1Lk0/xAMtMbKxqDx6C
niGCrGfamFlsfwCcO8hx0AlVrQ/qQ0yUE3OgqytzCbeYfBB/iva3LoF5YqcmDb9U
h77FNYlcotTh2NE8j7NvRCrd9ZOxF+O3yApP00gEm9Kyu6Doq6Vfop81fWtlteuS
PUdgCcmBqO8IxcvAHOr+/8f1RTmxhEvYYfE5fZHeEgbwPHPNNw1EmJBkkwhZFHGz
EuV1fgYqeP7kNjGON8Oj+dEhlC4Puqup8u0O4nrNWVrr/bGEHob8K1Wz8U2jnMKE
sKoO+ZLUe46iDTPIDAkXLgE+f73ezr+WR/81I18hOoArrwjF4Oh+wJAMq3H8xjgK
BLvJsQQRQJIhQLDxZlaQ9e0bso7a5zKUJFJTotzVtCyRM4fQ8pZzxEuAsTvdoedB
YBTpipJYeCoomB2BFMHp2tz6S3yV1dLH4loTLiHrtwS/o4HBv+39pFpozTP3P0Gk
wnWz+gCtEvlLroVaTDMorE5AGcxZ86Ca3Gxm4YEd21fGGDVFvcNWpROlOjiaAI3C
HXh+5/BLhXdLzFoUmtnUeqOziXzfZA1/QmkU7mhDzbXWtm8fZNFL1jacF9HLld7r
qVD38fIjSmDe3MUd1aSDReLGLrhYGQN2Wbe4bupWHjwNsUBZ9JMhiX0GoN/pHHaN
qF2e6NU/GZMKBo/dOvEOgwDtxtkGB+WA2SKh2Db111PN+VJ5oLhHIBNHpsnHMen8
XPFYDXRBR53SdlGkhxSTF/3knYvfRgU6k9Z0SlBuco59Baho/ib4eyeP1s4PjYyS
PNEUQgHIuZnEYlLYRE4lUWzJlYv+x5qMscZNbPW7iBohhaxsmh24/kMy0xUn5QvO
Dex6HLfp8TLjw/VdmsuXxcGMyrO++wyrdDQo+J1A7oFda6O3z7VjyiTqbPRWzjZ5
k63tHHce2oeA//DcSRTYpKnXY0/Wti1ycdIx+ckwQoQjq8CuyENGMvOIDD0pR6I1
qis+ynKIlDfwrXO2Je60u26KezUo3fviXKCMZLsXEJbvsK9qVnHCkDYjHe5Qof0a
OFh8b5+JdPrwLJte90Cssn3NmwhbbbBzjE53PQQcWhEk2m8OnzQWLzEEahJJG3pd
gRfew925FZgcLFDYVf7XAfmtkzDGRUvYCkrGWX1e18X91zJE3pD2TNWKBuLu0oa2
qAgX80Dy5LZ/+nTOFZjE7hLU0o9+COragRubTQJv/I+AdG1a2r17BVLDI1M3lwsJ
UPKZZvrXP2VwKvgWyrfzNywkVwg0LrM6UH0/HXk1v5kKvxRt5QGmJ2o0u+ovGmjf
WrcewNWwpnUpbb+3nAAjF3awiP+BWvk9A3MN+dmFRaPrAB6FSmwfl3XfoF2R21nS
otUepMeT/vhLZj9iaTW0brtYBKfWFnYt5Yi0JVW7vXDm7UgOg0yYsAh+XyjkrbB/
0y4Y39uwDO9W3KcYQfOQutmoRCt1FDEnY9ZD9+phRg8hOZkJF5Y0A67iK3z182mK
7B90TDoYTHKtIaOrDHPrb8TfWXYbb2uDLhouVlWRJZwEOimyV+roz9j0jt8CwBf2
CUxlPgDWL5CSs7Du1sEPnZ1TbfS22K8Med5gyuXqvH2JxwyHULgezfBjRUoHFt7k
yABJF1cvBg+AChbRl9ZgtANKS7shHsS8oD8MLbFZmsrQvpYhlmNhLlCKcdbt2ATM
D1kbdBjEclSn7fswRbosHbauySAROXvhQ9duhMpx6OnmP1lWDEKeNkzD/G8ZeDZI
ySBQ+IOmRCoc4PnT2DqbBeFA5iA/BkPeS1HW88OGNdvgtLX6KtLJ4TAOkPtl+GQv
2wL//IsRWyQID5cW2qltJotqdsZJIYqwfo1w5FislP+sTYBGbgR4tl4FQO42Dn8D
iePC4YkaXwpv5VLa7uBV8k0nxM6sLte20HeWFX5eUFGPsYbstzKDY/KKt4YH7aGz
b821v+PSTjbcn0k+MkFw6YYR8A/Zbr+6vsa7Q1errPXm/Y1QgmtW7qHu/3FHFV4X
goLZjht1LHz9vlnng9JkpT/wwSVSWUAUl8FWHYhC7hu2n2QiFRYW9ChdFTamAOiV
ekyZPjdLzCAjTMd49C7pljvLDzuEr/wTY2TmHBQs8kvXCBo8tZ2oR5OJS0FYIqTl
umb1+zhGSf67h8lyLtxsbC1chXe7BQMUIyukWdLfxSgC6AZeHeaKvMUcyd2uSR2a
lxs5USrXX5DOHwRUAamQdVLkFlWfiqazYCSmbuLKwXXsfOAd6ZwYBbmhXLuSVSUJ
v2Siyo8yHeClVXrhhUvgwc5btnAKjc27wkvDp2gnpvw0ALAk2Pxf6SL7duHjc+f6
Dl5cY7JHu6YjmeXt+g0DodPQ1rzi7CmCl+D/2PKD51Urh11pdkSmjxNHgtYxNRx7
TDWdS7UclsOIXGmFEB6P6452GnrRFc9xSpiQBSo8PJW6qZlWAJ8nV8H7WG92wUKe
EZ5E1oUy7rI+bw6+x5rfLfiTgFuTuqXXqZmh6FtqzV0eG+tozyXmXFMrZnIVg0GW
0amosXGczsxVWqnlwAUTZK3T+TQAQxe79OMVOd0V796d1d0JBOMb4FppbG+aI9DU
Uv21cl15DKXGwNzCm6iZdwygWaeH1t/EYdVtBT+KVBODhQbI3oXkI57jw9OggrvU
aTMs2RLdeH6FprJcYNLP7LEZ7cxLy3SJ3MlMJDkdqk+2zIO8ks3TZFUn0qqsjyGG
DNJp8jweb8j8IghIx+Y7Jdty/t0f1dXQRJMTKEHLlbe9EggBAPNzv5Gr871PUeRP
3lPFzSfwfh46keNXa4hBo0JQUwLeCuM+UVObrAcLu/zR2HMDR+5u4DXmE0wSrFZt
VyJ9Yed8W88qMqGJ9V2Ga8/1eApzDBJuOcGsAh4eu1WhK3iaqxVcht87uK7dVxcz
LjSmKjfg3TR+fc7K8qkWtoyp6bvvByKii/YBsZeKZO/2u2mTPX+ShZgsiY+4tQZh
BIUGo2C95JHalDFTpbbkZqjvUPCK8OBk9OOQ0v3goPChRpAmvOoAsaVqaC3akM3n
1aA0AdhCWvWuDBKBfvfQisArwld68njR2kXaQBwxd32RPvqHbsyaCUeef4A4RaTP
o19GaYNgB42LxBC05HS2CRBc+vdwRQ8XXbLncHlZGdgyfyyygc/QE0cfKsfg64xQ
pK1Pw5W69q1OwiVfQGH/2gGgX0nqVR3qhIPbXgGCmZ/hlmAgEOCNrcw8V4QbDLKv
dQNpvbF+/qKD5OBGfFAFne7X104ipJm+SsGuhyzqUL82JA2Ks6pqKSwIAYffbli4
qV41+2Gam3RS5pVN+C9OyPhgyatR/1HLx75LHJHl3iA2MQVnaGtEr/k9DRsOEmc4
86YH00I1+y4EF71P/3mrj0IC3Mmxkiy2mz4zmg7uuFiJUw76fMT7qsDu//aClKpJ
OSUd51AbcdP2kqx8J5p2E5kRHgE99SpW0yD/YuByXOvC+2t4cyD+hEJlrr60f/Zf
MMepnV03/Lfl+2KDE+PmzMkl5vthzf/S0lWBkHWRLkVCvH5pvsZSh7vjP9iIYffN
6X269hgFS2avzN3+Bs8RVESdZjGNIlj8LPlUWWg4iD1tJKuTmyZVP8s6rd1gWfOw
5JtFFCLsxYo606Sri6NK8rf8JU+xUg5QR392FIFvWSqb9+0ANdb2oDXABfijUART
AI/YAiZEmi4/W3kTBzukCGLHly8E7TyRwmRCq8kup3IVuogqzPEBejAMZSfr4ZNI
kHUJbD0bK9O/UDiXDLqhBYwhTDjGdtEj2GPPDr6jBe6WtFtefbBPsbfkbVCuUhqH
Z0NEanwgq4jLQFSPB9o2hnfAg7ioNWxP83s423aCO7OpqEf6W4hbIaApBtJaYNMQ
GbtaOUDggSsujOILk9/OZ61nEGLjc9/qSFqSDFuI6Af2mqtGc0jYuV9KZKhuqHTP
HSYNZF/77J9jxSDHIz/RP4tvLFO6VrHyjLyQE+9Dy777+ePXGK0kwjskBv0Yjazn
vMXm1wVrhBYui62gwwnShzJm/Kd8ig54+extlLRIyjrG9MfCwthwTBRJCEUhEifl
GhGo9YYSXjyLspK1tdCcTlFERLHsUnEfmvZT99zpEk64M/549Z8B1P62/Xl9yVAm
LL62gCriyeff/I9XGRS+SLQTR9uXX8QqF8Ry/KKVA0dy+iaK3PjPjrbvhuV2amaO
4DuqQPAMCNlaWzbAgtftJW+ilsqHujpch1++FINSnikDTsAGjOlUN1sh9KHTs3Eb
RlU1bNWLcJqgSmNwfj60kbldbxSJe2tdJDk2WfJ0/1I8o9oVEnweZXZ1pDQjsDuf
xASQEpT02cY9bvgDvvAgVbOsu/HuzM44KEMvjIYEIvnJuZb0nSB4eBVKRM6fuW8A
+n+HAkCYpxY2L042YKKsKnWbVO/AP65KXSyoiPrGS4vdu4XlqCYCxBhxzC1HwS8Z
u0YqZ0SjWhjPJWaRMxhR94jhGn31JXTG3UfsFzSPJwOKMzl/ORSWDIZs/pLg6YIn
E39xYj8Fc0dNSMOmTwRPs4A0KNF3tU8VZpF5Ggj3rHkU10DKhsO9Sw+WwmR2HvKi
lQfAPJg69Xlr+BQALKV4LdOiZOsMzVF9F0gjA9fqHWyufIEUHlLDErZDnXYvgM5r
wUP4Ch9Ig+WMBl6ypWODHsFP8AeNchbpJdnB9z9supwdVUgZc0k3exRThD8pQbtt
Z9ttxaYtJ6MAUQ/n9EhIUr5Kbnbrh25KZgWHtXt93XNGshWp8Jifu+WbbmRm7qqY
SIHn2CKBsVzbFok5mAzFAuZPLM6hXr/T828WUbjuBJSsdmPhSoWIByUuw/mDtHxB
rfagWpPTuJxCa2BjvYPD5GBaH9lR5s91p6bfsK5ViGbwas/EJwhxM54Q6ig9zlHW
9oluMy49VBBh4wn0oFERMXgxAke1c4nBsHQNgfsKH1HFCDXK6Tya6fBdCXRYpekZ
pVKubsY2ifWSZLaugsxKGA1ajX70cMBa8oWgB7Ztt1ZOICTjveO/3FhDpXx0hyP5
qsStkBpdmPlNLkkTBLV1lolafwnqQAaKJGimrt/xFFkleqRCk6/o667avjDuq9q6
/OK9OQsnI9H9mez3TjPSyFo+Hx8HclbyizHPugNC6mm7pBYbiGTkuHfv3ME3HuY7
/kH7JWCvzoePRF3Q30r3298JeABMpthhOb2aKyvWk3ifAyagAz/EQ3oiaUsIt29a
8kaTRPDo0jJ4r1dfdhLJ1HXwlYxB3xphVA7H10B25MeG+Vs1S4WRvDCFNxzmZN6w
bdtcq7IDg32yQopiRKR2HgWENKpsLbBHiS1I7/9kS7Ep5DcvGpdcnq8KAYVrbRT5
Y1aeh0KedBAN9XCuMcyQEmqVLNuafTYOA9+v0umwuKk0IpChGcw8Jy2rJrGYazpZ
diof9YUmpcpHbsC5QIZ2fZ626l7dmxo2WkG0Grxpp7oJ15nncPH3l878mYAHrJJJ
bPmPgMnkzj/yE05cTn/Ke31wzEPlL/PlebVrxhdojxPx/tlCXyjvfSTI5YSAQixp
65AzPdok59F0Ql00Nyt3Gyh3mzhTVE8r1x7K5vHLP4vbX4zapojky8i/UzlFaPVy
Iqm4xYdX3Mp5GCsbcbKPSMI2sU4VRg0OGltO9DGTEaY4Emx+VRQC4tgztESZs1wM
x8ouzGZ903FrjcMcW3XzLMP/8Ae4Fq7RDIp346G2ly72gWGrhgF2xef/EhRPPkRo
Ncs69ynbeDaPYvU6K7UM38kuJyPFlJ2sopyw9DL3nwXIxYDVm9tt4qFrNMkwDPFY
cPS/3Yn7U2wHT/7aoPX/xznLqlWQe7Va9a+2s6NYxTHa/2ZBNIL1qs0M/BI13JDL
mCO9kgtk8mUQw/3z9RxzGGegVx5TafPjVCJqjBTp7DoyHWEfFgVL+Jtbfxu8Wtsg
ZHZV3x+UcMRFxfVfp6XJWtpNTk+f/EPIyhgZOWcaRdV2P4PcoP6KP/Xlb26w7NWI
7nSDzganRXIkuPbpjeyl4rAAAZr5C4Dj2BNG89gwYYEprBBfz9HYp9oAvkmMUBWl
Q8WgzyFQfrjOlpdzP+00P6JlAYGvIuCojD3IP+NkrHmJfUMwVQ+Y5Jlo4cLkOk8a
CSAZHECCcrrbfv9qbmRKgKmMG0TmS9Ywe76KJ6eZTc/uJ0XkkLUnf+iTE3w+4t/5
/8fsC/sOEoa+MU5blDj2dFu/X192ZXHPxgImxY/Q+WxUQXzI318MjkSHLCKv6+rW
IHG8ZzuLsMnGL/xsSlLzgM+X7NNnJVwy9PQmuMhk0kZsITjSTz+7336seTg1x2Wb
SkQ2zx/pF04sfTdlUfBNToOuMgmAPBcQFQ/DN2bS2ODm6XwyR3rHDXsqxpnCgj0I
GYINCg1Zn1oX9nitPWmpBAGxgJBBLy6WQKQUgxhOVcSC1nG985PbWUI3KaANuK0t
f9PS2s7RYRhbx8iuosPl74RS79EDseMOtFoKDj1FzWFbTLYEMcY3lAqM+5HjjVrg
eKtMQwdfQH2OBN2pInH/m7btoYGnmqQ0ATG6RyJ9YcRbudT2w7/Rk/9+sVPWSnCz
5Xl8wgNubUbS9EzwmHIJ/rMsSTeBiU77yPMklwfyFnqj0ZuZtNIoj0k9K7M+BsK8
FWe6gWqxyMujQ/cO2rUtEKLIpEN37Bu1KvRmP2TsB1cSglZ5+VV6p0pjuU62P1fm
VsY/ez+WzMvwVxC6HOweTRBssYlfHmokUL89bdMwN8xqu7eW38m+IN7PZJ/xFXw8
upV3Xs0PF8JJM2fnCZO2V0J+oqiFyk4ajLX02vQsrMG/zfQbzuK85/CJyOwkJcIc
oJGqY+5Rny1tfJvcbLXFVefGTY/s/L0p45sjd4fVqYIRiq6tXEuXv+Aw78SCxdZ5
dhLbK4piW3hvdzYXe0RbV+VoEQ4iVcKmD3D2PRvhRbZu2AyCq++CG62uHlCJmWaj
T5DjLF2o+7/GIpweWoWT0FKzDuY7y8Ovp7bW9PtcO7J6fMa5MycspyD5jrTXews3
fHm04PlhII4DQv1Kq2cLsuxi9HGdQ0y07x8p453AIp1CVbFQZRco2ZjBw4jJOTHm
gk5FZYoKr6z1A0Tugvz6w6wDKrFfbTelCqUK/lfaetgjWmi7Q0OCKuBvHAkkTaOe
W2Bas4evlNdEamgb7sJ33VWyRxuoq5zSPXiOM/Ul1pKRJh7RqDtuHPQOO/jUfdSY
rl3Q0PWR6rmtAtFX9tnNDPnPCHg4Mdbl9XVEPKtj9pimGiLH3PRHfcikBCAK8+y1
ZTEGcXojQ5dC/VtLalMRbgTexVMudiJGo1xKVnKD0fxahayfqzm/1Ie0fwF0FOcV
cszOtle9iIBPoMp4AdSSp228oCaYdXK1+OBjyggBGNQ69IFrX3TSo5B+4cY9WZFG
+QZptBKlBc5lkRmmRg322IlfvodCnkr+bTLoCO+mSgbjoVOXLdZWRNjy7/yUPd7s
UTw0Em8Iy992Fepg690v0R+RmBVwteY0px3fWsW0mBeaLM1a6tKEIkSl/cEhZzsm
cdUPrHeTwzGmOnt9GehkAjxtnt5vUGSAVj6zt0NzcDNltqvPhixrppJATvVhpD3q
mR54jKZSIyjDArE0FsZzxa0DnKasllVd+e6lv4xnw3SZNhaJSqNmGfhEWeE0Y7oA
RKKxZuwJurnmMG7Hay6rlm5gSczxBGRV3rFmHuUhVhEb38cM4TcTgeCxNNgbE/O2
5ZjXw8QFYgxDvARl46VKuFiH1V7uw+ajaemngBu1T20SDWJlcMnH0z2+wN4gk94c
rjH5kc+sPPHo2HNYY8ATnLvF9CnjfCNV/sqkz3memkbXRVdwYaou9RJTmOLLJe71
TK0Zd31seil+MoPiOqG7kKIWWVBKpmbptqHWDT6tRKXl11kr/hD4q5XtxjvPd+nV
byQOv/gxWv6Mm7xmzhYd6zbDZqhPA/BasBbS934HyI57CUPDrZk6SjlRrUuFbdAi
0B8kbVt7VGVh9IW99eYOYgEa0otTUfUufC/yrrhr5dAtDWB+lhU97XTdNfLZhQF4
ev12xbgBI7zcQlwWDHl26jeR/DDcN/QD/qhdjU5EYpYUJX90GgXu1ON0Y1i7mfi9
vmg/wELYfCGUxZw9SOcVzFcrjclUB/dnCBFRG9K3GI16Jtt4PERbSoavSRPCvlzB
i2LNzREsOPODtFynLQOfT0/ru8cOZzZqZMF5I76LhfduoL2Hr2VUjqxarVTVUI3X
aHRs99E3r8/Xxdtc4nd/sWoZNCZV5sz4+lPf5ZM/IKynopzAqsse3EIyPgu0gvdj
Q8xrPcKUUFlmHUHnjHwvW1b82cBqTqhSwY6wl0j0nfEKFnOZfkkCledaZWFNUvFa
KsKIYZM5uvUOC8/bYxYlUUGBCIAhxbEQpDF9BWoOP74YjVip7/E3AsmPBfyk/IqJ
VJsFNoe5TRI6Rjf0P3ArQYteTvk2FOkRVtnOlj7RT48flJZg5O3MTwD6noN7zh1i
qqe4EUD0d7AmGRX8QVSlkHyXPmVOfH/afEend3a8pSE9U1fp5Rlvo9k0MSFVvyol
FaIQlBDW2DnpTodZ5tXAzdYRFJWbNDlmfNel/aLA/bv8rwSPk4itzOwP+EGMTwzC
kVQ/RapqSnZdhxK2MJ0+enmCYz8HYi5qRsI+0dRw20bCMwRuxYDczVX4G2/CegKD
QMWKnYf9oRn9lGek4/vdKZ+Z6v4bcK8nZvvB5lk0uvtMWbZ+d3rTrJxGKt9sefPp
6LNHGfNktI9OAUK5Okm9NH2j2rm3KmOa+Ten1N6HW7e7ZvSE5f9IBYAJwisDq8NT
V+5A0YW397cvMio1tlmUdP2+aRWMr4zxva+/bd1kaiBp8aXF12QpbJ5cMaBRU04e
LkTxhmEq3MAK5l2jkRWD+Y4FgUAG98DjgA20CU8j+j7efjiuPTYAA52Mz8zseI1u
u//L0QiBsc9ee4wS/kmj7hCk8Fmh9r6vknt/Bnj3/9sQ2+hBtO7B9/A+gSj08JbQ
SjPhxCYsN+EaqIWNIDbqG3/LmH8HSlB9vgSDU1k4uhkixrxboBbf+iu/VtdrAILL
JsAqnES57WIeDZnf4FUeoAKn7k47Mw27dzNKo2zmdkHIoIkQR6nWi7C9qIy8gxpt
GCdMKEyqlFLpmobaD2/EIMLz0Q30ZP1/qmV4l9mqIVmUm7VM9OrAr5txyOLauYC5
PIazg0bdNwUrydH+7qrN+wUGl97JxGnqD1SjHkqVBeoJD01aGndEKDD8/gmUduBq
k+u+mOOyvrPDpGC49S5SPzpCwzhbS9/8LNagZZACLfDP4Ms/L0KwOKFGkCc6V2ak
ZxvTVhSf5f8aCoI/E9tELLPtvFKooPhwbTt0Zzq7+0+0HfEgSmaW7DEy6f9SKfy8
BmwHSGvKay202TpMPe5zNIBQjTvWm3ssqH98cBxXPHcHoxJdqK/nvE3/IaoWG/Dj
fOvFzIcO57MBX8/w69FyDgjA2vdkoGiv40bMyrbHpWnP0nJnJKBLZa7csqABC3RW
tJRWTX6T3xlgAdhPIHfX9NO2ktKcD2BPS1n6MqPA+4lQgcpdlE/4OIZkrk2Vj0IU
DX+vg//qHLKpLXel7oeZ3fojpWK35BbEtdh4SHUPN+7rentPvG+kiH+MIfWoKChd
vw5JltSwBdKACiOi3BVmnoiWr1RTGtDtPYeIX1ScmqTt7s2szNu68klkMPfX+7nX
OJyahOq0FKOItUw5ffqiygrSaApoCfDfyebeI0v42aiV1rOKDobz5Y4x9MsXVG23
kmUE+XDJWiozwnMLkE5qCYA0icL6tzAGuE3cxPVsKPjmuOlb023ms5fL6IaocyIV
nlioa8/FWf0rixATGslnbmEF7d7d5NXldWH2gy2tTiYQeX4+h0E8+3Db7U3ZLI+S
ucCXhZ2xnQqbALgsvjPELMiooSrSwPuFUAJJ/x8+K3gThN7xj8618BJJsHejKDb6
oFMR20NXinAxOlYPN0oh4Cj/vL7F0Ln+HU9AYHC5PiAltviyZup2oNfE/1ZYiOvw
y8/zBhOwIbTYHN4xg154TMOrrH4a7E//kHl0MlodttICrqCV2XiBvH6Xuom1daqP
VcjA5KM3hQ6kTxkOmfKkYPI6f9l7pKP+naLLTNWEHNEtZgrsBMmE3LBRgiLm89ne
gFrlYoUMQMJtkG7FY7wWby15qJsvo/bjwQvv1PWHgcw/OpYTqJhD23hZ63cWEuBl
a6PkSWmVFEXw2HcRuhcM09Ji/rVc0oCh+k7XgPvVsIAg6K5PNEikX23+HokARZvV
Lxk4x5vJoydUx9Jv7PWIFSGqTpwgpXxK4O5V9839Thzx5Dkm/xxC6dAArAwJHV//
BDSzUis/Bog2dpJJRKfcK594jNapZJ6UjEvcUUGzIS/HdqFg6allLxCCtbVr/Rq8
+Xrzqlgd23HUOzC0cDhLRRILxGVm/lq5wjaQ/Gm6YhxF5qqmguZUmSabKoU+fK2D
/bziH5WMCPU//iypKgZ6rNs3tDzzJoVPlHXpu/hXH4JUeqbNwO2+gp+cEt/65Zio
VzTZI1OmA6fh8CTwtipOQ5YMHf7AAM5Aw0m0J27NLbPSCkQurAqvY72GlUoZisnQ
PnEEWVYT+QwuiVxTD/b+B3xaWTaWbNQGx8T9JQzEUwWpGi697REkNhHkZzBLrdt6
Sg8OEg9k5lPQE9u43mBgiaJ/L/BV3F/fR6PMfJsziHkYirWay56xPWNkQXztkUNh
4Rhv439m4q2s7kR5zGEYafJUvZHaubseZtRdZOPr/jynGMJFpNYU1JyFNERhNX8Q
rf3h6RH9BcgzIGu/UpchVVKMT22SpNlSwMr3Mf1uwIV3hYJHtIib6Oqn/ody+Hns
nNQtdTaClu/9zswy10LLRgN52b239RofWTJLHWjS11X7ae07k0wcigyluTg2X7oa
bxSjtdbhrXUEBiQeT7Si7/VMpPKOeJ1FP/fwm/W1YwtIWs2trkq8deE7XOuBi97C
HtZ7Ox1WYwzjmozQiYOLca4o92yqn0zPnvJOQ5tN3ee+XgnTOh9+T2zJhea61w8p
DF/8l6IIUSgjiayhW/N4bc1G8hsqalvSgf4QyoGAuodQVc6ABnZ37+zFEUIoG4c2
fpwu64vwa6GAnKFkzU+rSNc5KeeT6+fnrguiMbSruYxcwhF6A2p77bkL2Ih+0qTv
mpEI6d8lOKtlT5g9zVUI+DicMtc9Z9DSI044gyP98kiJgBeFS50ES/jK/cuBtoHj
R9ZStHLmOZjqHIw5OokfN3nsf3SVkQbUbxyk5lqqRDQ+5evK+TP5FcapzuQogwUG
Hxq6OOO4MBxiEuSrwP6dUh60NebpE4LKuIBctrN911fa8aPswfpFyd2Mz+N8sndc
MROVzK4beHfTmpLG8nRNx2c4u65ij9D3KksMHduWUpVkgPP42B4F4/2Cs5d+TAFv
Xs3ZcJUfZLpnjK1wwt4vSa7Ija2+kGX7z2L1vc9yfQbiguo5rRfAdVPRDKAF0Xoh
Wz+ivDWjszHwl6qDWuPytbmfd2uxKimCxI2EJ3udz8QrkB6YADr3CupYSNNnHGf6
RkF8xbyJQ440jdSjgXTFIkLzSxgjodG7hsppdF0BSU6HCFtF+nSpHDx5cfvlGp2v
dANVABKuKgBTqeIFfZMznMfRGKs2LCw251jH9WM+V53XNepniNpGGS/chkf53pJy
Ki2dFSTjVnbnf/rWi+yywWWV3uMcm6t01oHG5gSjKy1C2Pzkd7+Y366vSxHi3Lbr
QIvYRvy5ufj7rFvJfO7ZGFGfqOgtDfdgZw+jDmNO5P1oL1i+Y3JQk9rR0qVl/Js4
ITJMcdzL8TV1zT7q47gokEUMqXlFbzB77BtCbftVWuX4rDsTtATRQ3Z2dOA/ZJQp
6CZFCDnBqpPK0+z6oqF585DVZdVYhfIAv5/Tlj/4aXtcNRd8kfi/SQhzRlGaB7Ay
l6yePOTILPqXNBF6VqLaHBfGFZqLUCaM4rdqMl4FlY4rcd7EvS1p+PgNV5OCainN
RbOBcUZXT+ilSoQP4nP+f4dW8uhiEIZac+BKeD0QOwWpf5fgdmA2qVwL056y8L8D
Lg1bQkFQAZTCUICb1dlOsRVGs4YLPSBzFc17B+Oe/2Np1SWAgzg1WAaRYo8kRb9P
zU75+ZAOp1QmJk9MTki+vSemt0J6HyFZswY6JsobF60Q2IN36BXDXRNjq3UD9yNI
Ha/f42sS2MqbI/J8XUvwYMUH6O/Ftcye41Gm6R3rVcrCvvgOCbn8FFDLIzySAapJ
2sJjxzDJ6hFlOvP1IeoKcpHMmUn00syEz3uOurFyVR4zPhVsi7iKJGWfqsL67u82
ioH+HKMp4/q27Atsj3qnh1C0dvxeC+FePiyqcD93yHMTnBBUJopx51zCs5PBLj0Z
Ju9KZl026z/zzLxkH54rySVv/ujgBRzhPezzCYmn/gya455R3w4Dgpi4QBeNLDdQ
rr5xj825a9vkTnM6opBfzRXhX05863P4rvJuP8aGX/KGPCXMVSHOJox/AbSMY+hr
aAcIgd2CV6qGshkor1TPvaYUfWbFw4YKY2NqSBoTCZ6TlaUBgxSYekoYhaix6siR
bYqy/GOXPFr32WVhw2Rjc3m1XJK3gGFucX9dMjCbHhCBsrzghZKk81wxGC94UNrY
aF9aBdSyTBoaQ/7FLaB0UUE+nuOSKNo51B+Qm9vyylKdF6wHS15jxVGkdQJnheoz
M+MHDyG8dXpyI264n0sHEXJ1csK0y5YY9QH5yKEVM2BUN757NLP5tCzc84vW8oyh
Hn2Mf8H2GilZIaY0f8ndAyYf/jEKVPzLGYs8WD2XarcrlXwR7a7NRWQIbDMgcab3
bbniNCQYBc8v6F0JvhTaQAVru4tytYQYHn+tvDGx26eeEhP/HLghlBW35LtalfE2
HZ74he1yA0enmyTQoM0ypI8pyvqinL8InpHU3QAQRgeGCtWuPBPcWqp5vyk9CP4n
kj4g/btQTvKVZiIR+iOuZqd73karLAsipcnVatAS25pR/L6XqwIDT4x7sBp7q92F
J7DSEcdUH6U/1SUzMgF5idwcnKkMuQaQC3IM8n629bbiRqrFPzFj+SCx96tilnhs
abgvUoGugQY0RbbaVRoM8TYiq9rucMHK4G421r0uyp3rTmGzCCPVYuGmC7kchc5G
Ts4jSQo3Q3ZgI92/C036eFiiaA2fJyeOK3qq5FGBYIMtI4BJdqpjLwGS+HVjq0FK
ClVfAu3HPrR9KmZ9Kvc3u133IbFunpxBUemdo1V5SM8nZw16AVJ+5QFx+0x+SO3H
SJN4YZbMxClD5T/pc2Qr16Tekrb4qmOOiHwd+O5XH21r6U9Pg5diFuP0sb/ahQzb
JGon9OjPx/byp6foY133Xi0ue2O5OA9LLLCc3uusJZG59OyLk2EK1GKmt1t5Etxv
XXmMr8uRAlALltGaAwmPYblaa/lucvqxhtxgtGy5haqLsuCwOmEy0GytSLj6ta4W
ItcEqdU1eFbQ/NVqse5PrCOlVkHUlJ5v7GPF40eGUKvO/zAIG76QK8l7KhUPz93t
0h0j0wx8sKBJEXK+5ir3KKkmCNcABcRPy4Bms6XZVigkSjvKrhcNBo+b1fRjfV8S
Crk9QcLyJcY8H4+ErjhAy68OAPMekKZkZi7Ip3S6g0w2TEtajCbOWgoeSKQ3HLVI
ZClW0VX2twnTJpcYROQbE79dx46KSVJNnhG/oVFcJv974AVQLgHHxbHCwWmJ2q9O
qCiwOZdeHhZf0cR7Tz9KnBU/GCcrOUEL5+ldzzeJ6AwKkwsa0a+dgPRnDVomlQqi
acGWPex9gfBB7rOSLjhKbZnS44rKzrAqS2v+ikuXHZ1hfw/SnOWDsUa8AfFwjcXR
xtc8+ZKxLSTkRh1jKqJTxWgtZXn+qXxLr+/WvGU/gzyil+flTxmh3nfbJRq3Q9QM
7ZyIBuQ5FiH+qeHtJ+jyQ7cmynlnFekQqkdaNkpasl5g9FqCTJCkfDPFOsc377kL
ZNDfM1kJy4LorQIkiPsVIt9oRSGu7s18tf0cxP6wiDP53hFyvF7tQ9XB0QsVLy/d
VaojKBoVt40kKHgOdHV4TMvBzzd2Cn6g2uNAuHzMB3lg+FthU8sjPof6hUl+kiMi
V105kT6XHH0YIHRVrh0Mcw9dW8ju86IAmQe2dOKxdXNinYlPeFAx8cvF3VFFlBUs
HtKHRcwF2xUyzQfp3TDQnpP3ZxqaTglZH/dyH3Du9nH8841UuQvF3PjuStCydT1z
VCv04gs1st+ycwptcOrWKWtZ1y7pFRrv2bdZ5R6v/4qchdlS5Jo7kfJxU8ymlOpO
33dnRRaE7yCJVxdEAB4IKdK99uSog3o4Vf7uvGftOSjbc+3qzfIV+mVc7vr/8JZY
prlcaKzu1buvkoK/b34zxhQnqjT8BjHPxvyE8X1rDRq5SWJSYmS3WNVM9TcSfHBV
656SBJkImHaGtnqqSUkgI++R2DNzY/SQIxCboUf8NJsrmI2TJSqgzSgPQrAqmjL2
8pXUvfdG6yp0unOPplpeaa6ojOtV9SZOE02ZdX0ot2DJnXRisAitCED7EOIy7HYS
WElP7bAtWqNLBr6m0FGrAFKdgR0CQCRcG5YsafNRGWdseAE6itYiPbIkayyQa1q5
PmpbXIJ6lN/HpNWEYWwrou9J4TH4pbzUO3XPEmTdGR4uG7EoxLEKuw097SQZWWxV
wWa9mJ9Ttkj3qSYXR7d4wulaARGSgrvZWKFrg8SSgvJpkP0HbyL3yA/FgK+H6GbV
DJauX7jjUQ3rcLJ4RY31+EYdSb82G3SBBgOYWOmjyYh+6NUb0nG73w0Hr6/50sCO
y2M0HVAh6Tfedx0hk/GXouxUHJTbq84IY1FzxA8oSyR/mYFayS0H2g5a7lYF1lS5
fD7YD6ZRbfJgEnklmdgL6JKieY21rpNWHG9E3s2LzAZTLuwtaVxyqQpZJAm4RYc4
DjblGL+jJ9q55ybxRFqc2aVqRquqo0p1nGU+xepX+h3mIRbyFsADtDMRbirkgHwa
ONg26vQrPCE9GsRLWfUZkuHn7naVQV5jC6/BsXDUBE+clOl8ZRP7GNkNvUXVdwKu
9+1JvBJqDnFtgI73yLJqFZbpiPrLWrk18bNL8BWNEOKN+xN8bcovqMaLbfOJnlez
8Kc4l9eDdzd8LsMw5a1DeWsb16u6yvWoETndTPMVpubi88bl89/Zlf7U8r+IVxum
7ila7ua165J2JLUTmCAxdAIvkyyZcsOUgP4inImOt8q7BTg/9i3W0atiHyeMklr4
nHh4wbyWEBEGZY3+k70BbX4O6GpYnjLVKzcf2ONvGtgpkY6eETUH0eMcNvLJyFwI
XnWc9q6tvwjy/8sOXtdx24GqiSVsyqk3Td1FMarbbPy+aMpX9WHFPjK7W8Xc6s1h
q4aiuknMWr900QFGP8K30JAlFKjePIz3cZGXrty46BLm9j6UPY0b7MabNHP/miZS
bpMCOvQbmP80IFPg1lCqgvcu5ahKIgSM8/cZs08w/VpxTzPnq6pRPZZeqq8HTUFQ
qcGSPRgHx5K88ntKPwdeTvtDZyoFLvSqudh4TnmMdVNPVU6zZmUkWwZeU7ymo+OR
gG9o9P/EPNpP1v55SHwAtehGe5Q8c6nsWDv33CO6S18i+EkqDTsufl4GCK6Jw1Tz
eDa3chErf2hyWEWRG0fuXp2ianzmYomDCBIKyYvzq3QtMu5EThx0J+mvWumu448+
ephHgG54fkksIA1wYeR8dBbwW/nvVoJP2XfjNP/cbDdVhRu8yFyr+iKhD8hZQFY5
Sac/647iUpqFN9+I0mqohS1Jr6IMshFz/oB5eBc9X422CN50QDD0bfTkrXcee3F3
qjou0P4l3Eu1MUkmU4PllskjVI7WYSHpNOTbnxlj7ReSEgjy/XZerrMlqVqlyFR1
hBr7mCWSjJVS3n25tKVODPLybW5wajfc7elyxg9rfLbmRi7qkKB6pAo4+BC++bNu
ww2zP3TMp3v6nqbztwtTe2U83Rb2ks2oTF3auCuQk2YwWqiahc1YhweCUj2ldXFS
S8HcEL+1PkMW9w7wF3VYL9Fvh6MRmbQqeh4tPOs4Zm2RnKUaXpZBt0h1J0ejRvzS
SJbl6aI3bNA9CT3ILM3UyW85db7Gcq4m17QsslnmWRGFS5CMz1fBr5LQquMu3Atm
pdf2QM4zCjufaajjmv0DlhzGp+E/u5i69n7X3blr3QOV/fCiOYmjDbXoWMW78yvb
HyqW+4m0NRhC5azE5+FENv+RAHeyJHYSBXyRy7GOITf3ABFrP8OShpmMZOKCXgls
wxY2gHwpXr/OfmREFWhcvLu9SaaQotN4MWwQKokO1m1qgVgsUjE+O0YkgKLyt0vQ
gH0pzhnakVhsIDuy7k1XtQ/qEy6Z1OWMpMtjs81nZbax9d/D2cFIXnF+EjJZu6V/
ki0RN5KFnXftU2DuBDJlLf2vEdmUUm271EzXtFg9iKStfliiCtaxZSLFom5+68Pg
ktY+58NVxj+NjXe7VyuazS1zjaBqAGLtexRxbP5Ao2jvKSGQzFVRPTMp/VRiQinl
d3QVadLif3vKHJgtF3+9Suxnjlv6GmAhkFcRB/neCPRvbszz68//In1rHcfRaPbQ
6P8up2RinU8Fh3Ja4B4sQICGuRN1Q5S2omOtRZPQp/1I78LGMS21qcb0smkqSVtB
ozbM0XsUKAIzqpr6TePijIQtFuTmvL2JqqYtcd9/3FQP+PEnXSqrkfgcQYx8iOu4
stXcs6IreuXGQ0BR8UOVw+A+4U/O1pRH1nB8ImiSxc48gfqGxhxkMitT1mz7oiDJ
26eVKbFHipnY+cFJXgzk9I1a0zheRH3v2r1ylEQosmLASrQ/PC2lxhBiWcZxKeip
dPa4uzKs8a3aIZB7lCawK2oHRWmODwk9OcOGYmVFSsjryQsQ68P6SeVVQERsKcjb
5N2SxKmWdabkrNucKyjtgiCl/rPjc1pqvd9kHM5w8crB7WTWShmhgD6o/dSJ0IBp
vni4VHczkkgt8u4jn8++eTgr84OnNnVDu4CAnx3MA4L08gebSPguIWc1Y70wVgSq
QHT9c5LkK3ciG+EWdADye0vRJHzbTUB9NmPmNhaDSfwYVmzH6jc2UFz4X5eQZbxU
ru/GbG89MrF5dI0asKifJiBez4DA6zX42mG2ia2BdKv5tDFL2MnROpH7ut5oL992
qmf+XQPQIk2Nk355DNYBOXBc7jGFAp09H7nqzYuq9rz/0alNGEDZZ8R5yb37Xp3x
LULTM4M0NTibFk0uqNkx7P2FPk+w/IqtjPsoZnD8kxgKMQXfvcttZ+i4Z934Sy5t
Km1QXct/kyxg1pRq0kgHQAEyoQwveljPKnXDaqPFxrP94ysPlwslRkmV9moD7VBL
syFgQafN89BQMSId8TeCM54ZZBV1RPBI8t9ScNt2ReUnHS59dGuJMzlGWO5PtSCv
WtN7TvgaCKbVfX4Req3QsdtGJ1uLD2VtsiUckTAXQjFYW6NqoUx1HIbxo8I+hOBb
uVJ/A8ulKFGfqL96FLEIzTNpnXNbqekR5IATLHufmGP1YK9aHAFlVnbrokH5D5qJ
/7RwCLUAJhJv8rGT2SlhDlTtgORtC+olgceZE4oGZ2PnmB5muuVBjnh4L//tp+4D
6Oz2LLAu9AeIVa5qyJ5m/W8s5DwsARvtdv8hCE0k/i3CPE7siOGYyrNriPCI7yIv
TIijFS9r5cP6VMNOU+6SC11t+JHZjxZscbADkM5kVG1UXTip7+jHGrW9HnhT4Scj
IJmE7pf9HA49OXudD/18ZXhCc7Nrz44yTrk4RH76iFQ6KSQ/WXVQ5mrYUARph1jC
tovsEgrWB3Oo1aM+IpCdoN6t7bCBrQbwCzd/LnAvLvrqF7jliYwqPmSQ4enE3655
47/988OT1W5OeHfZDq2P1Rlt4zKklZKN++WUo9S4L8aUkNDmOy5wOND+kcBl0kX0
G3RwGUlFs0ilbKcR84345SAJnEGRjnRmp8u9hsOd6nnljkyYIjbanhyU7QMZwqed
c1MuA+XM0KW2Z1LJ1+tkbmU7IOQ8UcE0Z+ceKSpcjc8YGm3JZkwL25LQLE08numi
x/F1UR+KD5UOS6HuNbrYV5dySEHMsSno1rDI96kG5rKIPfu1MQfCiyWsKzeLcKX+
7NsAnytFV/hjI14vdu1fM7hCJ5C53PEhGcoXXEg+jewlXhXNuE0BzC3hk0QvjRCH
FUgFtwpPTak7TrjwcyjSVFY/w/u7vtVbmpWv9eOtAA6DRmPETcTx6Q2C5BzREscQ
OV6rB4YjMnOd7Fkdo/hTMJRnc8KglzyKppcmKOLsHhe8VSu3eEyk1DbUqvRE8X9S
2inm26T1JLwREuJpC5GQRLLvM5T+adIPpGT5LOyMu174hqJM3KsqsfQb+U4Rz1L5
iRisR6mLDQND8CDnAcmjsZ5dTwtSHIOAFJKOpI+dcpcPpgWaBaSofjLKY9D3Pl0x
IZtg5Aq8mGmeMvUkmFn1lvb8QL0108qp01oShYMr2Oe91+PwVSxc66QjwqXyXOCF
JVoN3z/8MEZCWaSNJAN6BMd5hihWZ6g6OlaHhohmM4Oy70BZN0LESpofRmtpLNbB
hOIAC8vDDh+qZmlC0d5x31ewzBMjqGrTBqGPoPXg38qMPHs6NI3ySmxdm1ZdJsg5
H2L5al5pfiZQP7irQDpQs2vJWn8eoXHNM1RjcGAfBY5Vp+kOwUc+sxBQynTmSog3
FrCK3isZpRrtj/0ZYVaCtuXeVFB8rTSs1NZKhOBjNI4ljWy70VUFGkmvMplfKc5x
aCn53F7ycC5lGCAI5vJCJSGrOHTU/FE606y2YVBliRBGTn06eogQxhaDtEGXflHp
fF+3SaZVOKWeQtNdCXmjKGbg0C+0nyL2z8SDYd//NBRR8yogfn2hZOUeiXZqzmY9
yFWX84k+aEJNXt4/Dxegv0uve40p/pDLEgTsDu2F0k0eqmU9qwfX3Ccf6PQyPScv
rZo/C0bKH8QlxJpeV62VZN3XmZ8+JcbfimOeepNb3KdpIgMUWkCAPBqlvCRQDB0o
s4xAmoOgBJr/C0Oudh9D6hqf4tdG/q3kgd1VWOixBnoRnqXVrwxghbIUrww667PG
adQj8qRTBIn7kXcIwAXPTBMbvCwveNPlO1tkXiLhUXSeqOrb3QtsgHCNQ+6uqGSa
klIfbAtNqDcF3JooJ1WtWKE1rtKTg9L3ZBmjf3mwtNTo8fMGn5OjuYIx/FcksgDa
fXURx0k6/LA+hjzZYXc6z58bn7tNl471IW/JQvTVqbbZvsxE14iDHU60+hfJ4dcU
X7fUvtxwrNFwvh7AmmBq/pJZmRq2oVxtHDG8vr9w9qgZh8Qc6EOthYMLiLT6clr1
mRUqaIQSuJt4/EuJbi0wxGE41O/lWV1guDRXplZerchdTU7XF25qC8+ttAmOmELV
hHDHa/3cdhIv/uMGGuz2iULcigjZedBUD4dEWJewU5wRCCwDmJFqqY1exCj/9X36
aNEw1jmu3TWbrb1jhI0Qz0s2jiv+lpVZ4qnnDnTqcV+UbzOfqeeUvrZuve9/KMs1
BHhh35hoVs1KC2ioBtSxfrG77iUBSZT3Rv0pL1vdqcvKmvivRk497S+q0GIySBnG
vhxDp793SUQnhXoyHW/BHxIo7srrkOwUPrnPGlgJ8fJpOhmKQuAk3GRMiMoI7poN
sv8srkDv++G6fCIy4O/nnwlPEksH15mwhn1KrZqSaGIVt/ZrhpWrvtf4xKxUhLV7
Dkxf4hs3ly3FghiepL33cb99h9B/2uOBEk7ASYwwM68iiSNCdgceRflu1CBuyBYC
nxObIQ9FoZX2P7mgv0lRFgAn5i1mCyWi3XavYYPb45KhKusrRWIzdmCK9Y3/R8lH
4jGd77o3n1I10Ji1U39x946EWt9wWbuj/C6VnqizExFaVmPc7n8MeXpa59AcT/Ik
+GyrAAdrxsl7w1C0Yg3hxU6laQ9W8n+niR0ocH2FH19k2Z1PqqaU4Yd0d5QtjDUx
K3QBoynCQl1wt6eBgoo2YZ6DjDnBo5J+zRWM9r3FxRn91/yzrZ/tFNOA02shedha
wWuDEz/gY61WNlQO76KwoXAArXDj9zdf2effCTLv2YFhYshkVyUot82v8QWTv7KI
oDRwy1J1BxIK80GbZbeXLsWJqIUwA+abAc7qxFFHKuoqvmPPHUSwW7jnBJvZPg53
xU7SuFmWAkz5KZnWgzDkKGVMWyGAmqkLUNpS4z4QSx7NGaJ0KNLtJsizY/oW1eOX
xs6D4x7+wTEaUIycd/5gT0qCRz4offHKOHadiXv5//3EzTRwIe1usjafxRf3DpwM
BaLwhLjpPaCftXOVDIuKdGOo9cCuqa8hq56LrmLuhaJFxHDMZKqURF/6b6lMWAsS
i6ay2HafRnMEsdQljUCZ58w0VR25XqRXKkCcWfsCulv9k3qa9DoNC7JIFvzeLI11
4MQoRqDoFqF+4smZRXpyCsdukAq4fKw5iLnXnFXXhVXnA+96nfSbPTvqpmPY0P4M
St2MmkkCuhzeImNMvaJo5YnFe8pY9JKq2duykN2aLcmgJc6SP11uTSirMsdHQltw
UMN8klkWBeHbvddR+BHaxBhm/6q6JrwvJ1YC0CPxGliUdfo6wWUyhNFQkDGmQQgk
kEWkQiFc2MCqzLwVJci2J9Ze7vZp+71Wvr7SR4delusfeJ5esuwuD1ypz5OARAug
5kV0arpxXS7RYumRzaeW5KlaAkNHpZ5cAbVkpiqdO8iNUWEq4x/4OlbYxPPpa9hN
6eblqWfptUZ1GX5Ix8N15eqUQnywnogspZrTNuFUd1GGMqJnH2Ljwe8MvObZZXSx
W19yaf3fpjMeSN1dWcCBsoLHjakS9OTsEIX1zfzG9ijz4ZdFvAR/x6AzB2serg1Q
C19ClbX0EfXRj8joa4HsXYPyMkteG5jZh2CgaSojHG965IT3g7P+LCNgHXXFyROL
Vps4IwEsNhBwTN0PFvYsP+6ckM5fk31jFhsYc3eM79rhQ8Z/B70DSU5lJhZ51Cuh
x+syxPMH5qlIqYh4A2ivdiqdBcc8nyYSCyEC+tSwW5OZqWQDQSR76vfqGiyb39+d
k/8kJD56qDw82ujDtuXMxqeUl82ricQ0ntLie6pAdA3sFxie9rllJqOJEIZx6uCp
pUU0/3IPjb/fc8YKiSto6R/05ySanF7djfkYr+sYVGkTkdur4fh8fh6w6M2XeWYx
hYBS0NGnhJjG2grW/yQxxEStD+Db7YG6P0CEDbiDGUxyqYHfP8lFX3ZkbKrbJJ5D
QKUYZX5plaVeV3xZRaRI0wwMtW8jgDcFav8fM0ielCrZpFjeiSF1o8W3i19wO9AB
GRSdCLRxmXVuWfLmvPTuwJsXxN3KYdWLXX+F5YGB0tVADVBKbhZI+g47mBma96aU
J1/Xe6Qhc5zirZBmYtBvlNrSjMN1j7EidGqNVSNXtU3UmaA8DZ8K0QszVqG47ai0
9fWrah38V96+Lkk3QaG8FfPrhVVKPaXlabca9vzF0PZBj5LSSiqqNNTSwHeXFC5t
1X1XhMgxswostAhxr79XkPsDk0+wdpcpkJDA7/4y4nM/nyWy6iNVFmOUkOMGHQLD
ZrL9XYBAe9kvtfByN4+Lw/778O9lwKSePJXIKiFmDAcHbzk4pGRgTJ03FTN9zwNl
gsPaNuKSsI62agrmeJ07DCFhPcMgxJ2kGzyMFb+pHkscXUaawJLJZWYVcOf7uvWz
26S/VYFng1+ysxSFGYoB/rtqs22WprvXveeStEzmudW+mskdXyBagq3BZjBx2eT2
fp8stHGkL+A/bazjPUlUUvCgo4fNjeUO20oaMuJ2sUmLfUwNixDgyxuFbRpcDAQt
qPg7/Of1t+/4WPbUYpZCnGauYXX9Jtek/5M7LyBnZaNtlibyZwtbOTX05vuZTIL1
drm+bE1tq4tYHlwH3hEfQXz8F8FFOShyD7DbQCClHxZfpGbJiJFerMIz66oXLpzw
vrOydRgcG0yhoT08Ej4B5CFCFuhA2gStjC8WJWGY2GyUjhWHkwGWyQ8KgbH18mMx
6F6yapA7xmkaDmUSGM37U3/WMpbZa42MGoDh4LPmSoYu41Sx1RHwi1g8GTJlYaS3
PvfVXTms57yHdsdYrhS6W93xWosobGkfVLyQk/0M7Vgv4zWlayDeZypROLMdQqNq
8y4VUHTxzZt0Ay72Z0WJMKr+9THJ6IRjOsasgQSAbVdgN71DLCa4+nmoy/klMsfU
OeQ7IaNwKuIl9fEDGzS03W1obHBDwKu6vE/Mp9QH8V/ElsTQoofuK0TS3UAYsaDq
wDfqBxup5lHuJrAzqEsWEGcta8jhQYiBLnfWl46hDRoP6IAH6q71IGgYbs/Yidt4
0nLOmfv3PPy1b4mflBx4chV3j1qrCyy3z3G4eI7EGrBIu8pEt+DFXp38hSB1D2Hb
uijOnpQiYLyblx971iDEdbkVDMzTnxWHkzNBr0q0pxKVcur7A3wj2s/eA41dOf9V
wtSabv8RGNGgdr1MzREJmRQE4GCNtiy5oDkrQigxSDYcU2JoJz5J1sdO54LEEu/g
Iq3NzcaEDc0/u7+fzQHScRkaIzGHOMWNjLxeFvuXscSbDkWtcmd3WanTqWx8acsG
1eim1cFl6VexfCzwOw4Ge1iy9g+YaHnGUwHXPcj6rPIhWOIS5+Fx9kBWWzoTrZt6
GlBXLGZstrKvl81Iba9D0JsELpvdMYavZoLkMojAkGv0VI40/tFKbZMiI5Fw+uYB
ivujc8mzdnHDyVEH7pzbrh1B9aC75sqtYb7ECJqEinnKC108otfJ1K2vcOya3la9
YEojwu8nn1YDRpbpcOKW4BuQ2o4o86cO1j/+ta2b/B2t4uARQKBtXBPGcQrDBRqe
kS4nCxPASwIoYiateR9b8gf1xbjO9dQx6EcggLK5GSSDFXZB4NWc5lQ2ErlfE/Ro
S7sZr5fHD7wt8p7TZmigEoxr57ttSbcHtWyftAH4FJYLu4NXt3e8qOeNw/A/ZGa8
CZl5hk7BHOPuNXrZi3Vk/kx4o0ziLkJdT18lA4zf6qU3PqcY1les754Hn1/iZ3UH
8LWbiOmWIEWutE48LrBmv3lyUmXLL2YDAqykNCenIH5QB8oKdf3h/TrHr/t2dGU/
t3A11FbaqfyJXV122e12VuRCUPZmjSc5cU76HecJoUa1gyCAzis06moCcoq62cdu
CAz+6zt2IoOpppgLGjbM9BqrYtRYHCXJqUfEFmIceWuPjuUOlxzqFbc921w39O5U
TluVBmjWiLanptUcxvXzQKt7qxH5NdUBpm8ICX8sbkLOTor9tbo/hCfnhb0Cf4GI
Tk5ksqwnS86mCB/+pELZfda+omXjb6aGYqcy66q2Vm2JEizFswa3Mq9cXWvYpW90
EFSqTSUYh/wLfIC0ygifJ6j2Qd7G37yQyHn4DT4V3e4GFyfBaF5Yqs4T3oJpiWls
JAsk4hAAJLKsp3/GpQ9s7MDIAZ0Oj6YZe0YxjgkiJvkdfFZ7fmI6XlViP/hxoyVj
R2631jrL1bSwi4xGdW1L4rpMZCO61tgSwaFuXj6/HHszWGR0pSO1iSQLP8Xk5K4+
Pf1K5vDJpMtp3Zta+YrqSMQktgpujgd3xC1627jNwSkk3DOkX/GGtxzR2mzEKeY2
vQLjaW/9vi52HX/nkjd9Sr7SwjUNwtXJS+t/CpcZ538MPZQ6iWo7pwhp0h8zXuH0
9FPE3ZTaL7EEUNGLSne/sGNVF9E8AJ2ffRaBZqldXOd3eN9tEzEylY5H3Iu+yaJf
xEHsuEJovHfsQE/1jJNkBXxepvLSy3TqtJmietyQMCckuktTvtSjm98jgUXHfios
jpr1Cg1ZNR1yddQ3jEku5cJ4m6/X1DFaul3c9sv84OB5eHhjSDxXhchEDKJK31PO
+47CJX0vHR7E7yJmhSkzrO4pk+AKc5FPgcuRG91KJS+juYeo/rQj12C81P6LWyBU
IbycpUV0NPA1SuYV6EGZtpFWm6lX2wo8ksQPDjRJOd8eF+26UESXRB1w+hUJeOyZ
glxgvSVpSm4mVvfZ0Z4wa+U8PJpv07geItH/bmKbJTKXVJbYby+I551nz748lk5P
T1dd7uwq/TFtArjAynpqpsvC7pyOuk6+u0QylczI3KlfTD0HOwpud5Hj3jjxGIVc
T3oEQ2AuheX+epM0hlJ/0fiB02/lAqh2DKif7Dl0KQnlRbSUer9dXNq6xaX3TYT/
0z6yvX7HM1KFYCvrfvyzzl9aUzkLJ2zwb1GMpreBT0NrrsGDyXmoR0/dJwLo6FoZ
FAFj65tUCjp+p9hz3NMm4gznZ/icASoFa/6mvpBzfQr67g1te5Z7T4zt4bQIbzwF
UB/6kjipi+DXsMQZcRgNkOjcNVFipA2sHbozZGDswFE+uAgqJkGHbYC++03dBkKY
3zCaQu3YQLQHElmVLR6TZyRWaYbruSaL/CZdK5llYsafCbo9lmKxWnE5lpW4tTPP
4yvSsblzNwppiD8rBj45X4wi8HX7pVnEZCd3WbqAjw2oTQxdyeid0MMt22VnDxRW
0A5NVkE0PoYPD8lSDs5gbr6nigEK5ntFABdwF0R1kZZ2yPH132ATyWZDv92I8jCn
430Gyn3Br+IEuJqvIJbmxfaE6HOYMDtBLWRAb6O22F2znaBu54Nw/Pqd+hitL8sm
TpfyHHgYQGC8+tkaY7eD7rKSTKGGsXeRNFTsEHKuUE5QI2te/ixW5mui4MGiHoVT
BjKWnRc6ler9qhf7BkcZ0ycHUOahXRbIV48TUXjC9i2i74lc94Qrb2fyHJafOTCP
5mJSQHGY/40AjnqshNmVCWpgLGjUZB6KyvMjJ39lP1DDjcwa/UUuaf/5gw5eU159
FxlC4Lb0tP6zfzDPe1nNMZsyb/r3y9FrShKGK3QEewyBc0pB87q6pMEKMky3RhhR
FSqS+6W9oJ766ytuYgzqq0YuzpxlY02ZUJmBDQ7N+TAw+iipOqwltrr3qB8hnqj6
efSvpDdamGgPmjydNGzHIkTqFXRc8AT8kItosUDIUbzy3TpKvWwWxrROuK/K3cdL
nZqXQuAi1QgZZuFIdSY1dd710NSxr/kIRkyGFIluIGI3+RyAwMW19W4vYi/jZyNB
T9BoEd4nXr+JwBI7Q6ipZjkZ/fB5SoCLsmwedOh3htno12vsHM7VAqbUjSNFkGXJ
M72aHctgYMLfKrKxXtUL7kkiLMSO0Ao5Bh3WEF6DhOhDrz/DNliPh+Ya7w4pjVv4
DkcMCiDhafn6zO98Acf6WLpI28/F6b2Ir8+Voj5/U1AKWb0qb1uWBgut2Z4IepHo
szSoi2PktGweamXibFZp7j7MtOU44/hy+DEmRYw/yiILk6k9oaXFV73VCrQz0c+Z
jy9nYUCRl+mDfbq9YxWtVosnnDxHoLA+pqcMHPfLqi+mSjQz5c/efdibp9Yz8vXX
xY8vFrAhCx7nubtJaNxBofnDny7xSSlYArNoU11cIN1ghxWZVb+AVyJqmaXg0giB
JVdbZJS9412Lede2P1J5Dm6x5kli7L2aU4d3JHoRRH24sYA5JObSVujtfptHno/R
8aCuP/4fRxb1peE0x+de17YzH4GhisTQq8EiGtsRvtl6+HrCg+H87UO/JF+YDFGt
hWRAgljSVbUHcsXeEiuKeAn488zRNueGftDiihU9nXa2XRulrWEMEp/Z9o1GDHTq
qn94L4Dk6XPualT/SL1CcUn0V1cksSNFaP4Wgb/rxQ+T19ptTd0bKVQ9RknVXmoM
ZoBBjQ8uoRkKBjNCy3ZuXW4VK/WLKHhC5FNpZWgAeD48JtNIvpETLAN6RYdcDQKB
aUQsWciigIkTIShvfeYXW65d86LdIc2TtYKB2ViJi/NOjjJKNrIMcUKB4WwPtI3w
VlqJyo7iw2CgrZnflJMTV/eanaaylbXGifLYeD58drAqG7B5280Vpeyj82dqKSRi
3+EG89figgia+6EhbWah1JbCMOfEQmep6KGbrpslp5hSKgnfFKS6cVDyaGlkPgf5
5zsgvICVYNGE/PbhYGNLFT706r8ypbE2Ejoe6n8E1AX0k9ECK7cbqnD6oLnXE9Eq
Jv4yTDnDRhF072tT+BtVDHhNCY4o0GFleDC9KaprCVyghdZQh1HPd1hHWKEzJ9HU
8KEjsAl4mzKzi3RWTeNHS2YDwD0/nuQvAusasK1D4TKRFrouaiW2TWwqjjCWxJGE
fbvs3khfEeQrw8HS4j2bob10uQh433gdvxfzd2pLWBPpKvwfUA/jCEhzOmU9yhb+
LKAfbtMGuIXl3PWMY1Uf33xd+ChmCXHY4P//ONkMjzf02Wv0BX4o43xRMY61sOIL
HgfyXnQFfs8pqFAXyY7QP7F4dgE8zURJYePvTeTI+mnFXvM4UbHMKdYn3zDBLDcG
o0+wsQffCL+Nh5gKagJUfM7lyT0z8jVlu8F/aKNf3YXefL9j/b6HhJGrLtgLHtJO
hLCvbnhOYbNWO0di6RIapqqMZV53HyOMYqoIL4bs99tzpp4FJGcsUR85ovxmyNaf
hnCV/ST79gn9++z2jGkyh0SUccxJkLlWguYRC7kDOXyy3BTOJFJ1shPMB4XBndo9
jLIOCWEoI5WGogskoRiKcbME4u+EaypFlV17LE5pxPMo6TN1yD/06XKkE3PjIWjT
/gsvdyhvt7ABxUjWu6jw7RoDTFPvpKHC57Mh03jIWAQXAM3Mux1k+yjr8L21k1gQ
/2EFuJz/sDd4P5OGD4r5Y6BBU8+h3jgToqHj5ktd7h/ibL4q7wDgEMMA5H04hztn
rWQqWBoFO8ME0hVsCP1VhpmK3yC3waOP1wEoA00t0IrnMF1/7uTdwP9dVAL2QjyE
9b41GnFnFe+P5AnEapYP4e6iQA+TwRfInXrjxJ9dNSjvKCPZove+k9j2/MlMURvR
QDpY6ugbtMYcW7PPyJJHW8vQI5rWwYKv8Yr9RMvc3CIInDkSHG6xQZRLHTEEFCnZ
SU3H3yjqnvzVpQKj3mSoed48V3bALmTROEYqmH9tu88rvDNMjHf7GhdGgdA4wsrE
dOunNWRcmNp5ndZTJltkdEw40nDCyGsDBZ4XBBlMLJ3jeIT8DmSLkbJZ3ykkSMsY
Chf1aQDhJxz96XbYn0wE4sahHO+/9mMMeKBqzGShwgIp3bBh1OVUqjee6V0g376H
4H744r044+vLBXOoYR1uZSwHs3dQYf7XymTZDU4J1TKkMDQ0TixLuhoXupPpNmg+
IR9MzNC9Y32+zlMcPjVOKV1KXyDA+cTIRLFj9kNpCl2zuFplK8XbTWOrvO46vVLx
c749cEQ4Rail4b3Y9NRovtlU7sjSFzOWrPxCQAZkgJteYxhw3h/FvPdx+VkKQ7R4
iBL19Meu9Rs0cWyGug+o2CTliIxzHsc7jALgzNfsJlUE7cbNPt9xv9xQ1LYgh6Ez
ieuU0wcB5mLTSsGZ+NB4JFQ/CWPynqweH7v8biQaljQZQRkaRVNjqsYVOVb3MoUk
/iEiQZ8TkVWN5lkDIm6//RrIyoLid2KgVW7NVSvpLVuy85iCkZs3J8gpx7d5qqo1
PN0Qzzx8Mp4Y4kkRbj4yaJKvwuQ74GAIlnnhPx8a87VwcmmAznZwxXIC8bZ1ME+t
6RclUkHxQa3MGKIWVv7Ct2fYIQsSJoKaFzdy/CtiwlKr3b4G1ch/6KQrS5FRvpv8
hp6paz6WXKdayyPV3ol58+uyJvUlyoRwJXG++WpV3z1iXuqamTPpk0D4f9uaekxJ
QqEpSZ2uI9tz02hAo/ecJ+pF6A5fZC/k50kInRDfutlDMQtVKuRgqvc7QkWlQhoB
xBqgvgvm7OTRAjetTBJ4Qq2w+Gt5Y/UxmOuGW59yvl7teKK2qN1v/0OnLpmD/4E8
T7p0idvtoBHReFcAWxQH2xwQgZizySTD3QolXy7Etrl5CmgMxzveh8UhVUCoSpD9
X1eJL5/TUXu3Syb51S1Ucl3nkWGu7C6dGqHeDHozHzuBtpEXNeM4akf7ftR0dkaw
t5VV1hp/kEYTiJaxVImLcF4l8ozYti9yYE5N/8GC3bd+s7sW5rhkj3f/qxtzUDNz
wuiYhXAUhJssRdnTb8/shQVSu8DNpkJgRURkSafvu4kkVxXkIu20hn2r/V/DNUPa
pqupWTB0bCS2nZx4ICnZgHZdink3nU8eDbgivky91y7zSh4ml8C7Ry+xb74Y7EiK
4pU+lzQuN1GP2jybhgp0mP19KYwD1tlvrKeZ5J7XJSCLE/TMgZFnzX28fO3+Nr7v
9+EWwyhmD4F1Qx7KXyNdsXTfalqVncAzzVskCJwo32od6ARmjTO0SyZ86pzoJGm3
kZZEZHRX7U8OLYxzTv/V13TYAlTiSYWO+fYISVWARJR+lI+ishNfTDrRm3/Nf8Fv
Wk46QIuVhRHhd23dJ3kg5esxa7Q3YbU0cFW6juI0rxFQ8m6Ujm6KwQRzf4KM/vht
0svhP8Y5tALFhK7A8pztZi9FE8wInWmicEtctsZY7zSuCFwnjgkXTpsYq8FubrLx
xY3gS7SQPCkamyv9H7zhYQEerb7rcvtx4k1Lc+2SDfBzn+4jpzCT74dnBmkxxbQ2
ebLU1M0f4hONMqUxhbJuSSLscL5T42O4gIkIWblHj+6bGE0yorJftxIzjmgPRp/N
+8BeLABqbGsNKROGV0fTaze0AjKKzitSn+2NdpcqbF0hMiTvyKdYySlTmeHGH1Cf
me7/8joPQYlO9Fz+s6BdXaZDMjFK3VC5/tJvYPnsYL2iEhlFQBbRJ6+BUK6xJ/0u
Rq5F3VGovz7p3WmAcv0B2PxksnAatWuFrXSvH2hLaFzTDYfm30FRbDXwRxDiFeZb
t3uuYuKiPW0eBP1/9lTsqYetSB4P3i7rB562Tu+OLj9BsPk6oQ36vZjMLODNUv82
Ku2oFzRNI1FCTuFtgfRP9qoJygGJdriQxBSf+w8dm5rX4Nln/GqtMdwrft3SjWve
SyFMisoUtDEv+c9Up9eWOAGCSPlXY7UaFwmZupxo3159coEIfMa+NdGJJU6eazwv
dn/Hvq1Ws1jvf9R3I1Ky9LW5fQnT36UWQcRQO6jMWhQqBBviyzKcr8HppI7Z7IUg
Y8lAvyV1Nng5mF4aZgsdHrFxUZqVgr9HHQgNrj3TBsBGfUIr/GmjiG2TdJX4vVUI
9f/dndepXTQJbEmBjDetEmhsExJGektYWpK8kZ1xaDax+ATbB1JB3wO1rihSEqEw
WFrMHBKSl3Z4KzczMWs1Kz1mWTT/w53RfO5ijbtHuvf/zZVGe8RisDfeD4ZgIYKE
nQDnqPWM2QZj8DLZMiZnL19lP+0RCBMnBpa5cGcubO7WmKot0Tq3E8i0pWiwSRwZ
50lSI9/rx/Uv/QI050kAGNPwiLbDpk/zCMhT9fUD84NGQXO+KcIENPPxkldroVpY
QEIcRNEqzA9hPpHcraxRkCwPNWssei86lTNLKiRWBTv7uDbbbi9T89yuERKeNzPf
2fYiFfWQ+53izKzISRsAy9wdZWrnqc3iJEQoPHbdmyTOA3Y4TaC7+J63G0gZ/Qm9
sQfw4RPyHMV+Q+sD4d0V39U/1+N/rNKIfEMwo+41MGwX/ndQveLDcdmMluM+U98e
guw2/i/IV2jMYEy7Ci65OhoGb42ZRqqHW1GmyDZi++SXFdp5LxxreZkW06w+o/Fz
UDM1tyMr5mhBI0X8sRTvYOnw4872K2bveB+QG/8RWiU3hao7ZyRFSWEm78qRkq51
fU/vjVAh3WykODMdB6c+13nXGG2i/xroG9CCqWEAbI9jgYEutnJXgrxc9e6yexiZ
BTyphMs2AeGRGRW040UReFBcODKM5i3r1gpf8XV0PT8wlMB3RoxPODUBEu5wLNZB
S/BQABmKZzU1Gs57bjhz/37quo8xfOA1GTeUs083vFK3nU2Ida5A1QNxQsXmJaiF
3gdcyDsLPClgcCwC2DqAnKNp+4nXcQpPVVM/gD8riCwDIgQHmiZ3uo82V6/7uJ3J
r5NfBqt5wmImXVvazyfKCY5eAOgLJRzkAUtT1ZNMFnsTi8umqOLEm+g48Xd0ceeX
Sj4ayqj+zplN4uknJrP8TlcAPPu3zJk7tqiIij97g1tX2jzn0usV9ohZWtFwxnGS
+tZT91uwMKEIGBF5ZRRBCs8lm7YhHF0/DRtK7jR+P46ufde50eyNubNuUy0g9los
8ZiU3NDydR7hbgM2K5tt+uS9FmfqtZgEHZRvFlx09uJFaMrh/rIZvFcq+k0IVWbA
4RvtbNw+nzuDZMzz0eLFRao0c8sCswgLpaNTVvz245Ph8ohFt4zI2XT0QPET4wru
OINNYXNE7lO2hyqRtm4GWSaCOUZ1XglFDpkoGU3vJ8gk4UWCmRSfdRl5YkZyHV/P
J2S8fYKhbIhRKHhinvl6IfZbZwC11SCnzK2eVjAD+L90DJrK5ZkC9UFWfbAep2Zd
6+kvk45vI/dGzpokl5vA46blcjHE14j08uXtoRHgHXCYahzWXHSfe763XHgUCZfV
8UGQiJCnD7cuzdjVW52v1gzoBbOjc0/dOO/HKb5QljZvSiJpENdYV7jg3TLh3cMd
wywlWXta2OVgN5MIuzzttYPksK5XqaKWboHodDTkqf2Ox4JtsoACafk38oGhhnZW
OxwHuocZa8SUf1bf2TrFFcJ2GZthIv6M9aEZzK4UxBaRcXaKq+TR+5hYBP93QLVD
OKiCEg6jwUp/1yggp9xTsMgrR3FgsoMFBZh0a9KmItzUiL4TF/NBpITdBKpSwB9t
Uhh4V7/XUdIEyoNfvlOnB236oJUcTGdao+fshKwlDufrGzwQ5gPJ3TUl3ZuaqLdl
FD/dWgoyl+CvwKvacZKvyGsn3bwx5jn+dk8QUJvdzmZ7hhQ/XrcGabMxzx+Vgz2P
RsWCNHAjqQqc4o9iv3Ws91DisAFE6q2FzvZ5oP/yJ4/tEOy+vKUbKW/YnwgreE5Y
I+3ksOIw8OPpP2LALV4N4qGz2XNhA6rvu7I45GFrQnQxYjtvkzNfAnARLOZWw/an
CDP0DjFLeBkwsnoapC+/WQlpzP37ymPv5Tm99GkxD1KP//ytRxHw4+cK0s3/+gOW
Acxes+8QRAeM3Rsq7d5DmwewdASG3kYZrjgjp5lVQ4VAecqTwp+y1VjkvZByxOuH
acai7JADvwsk8NUvWo8n8Z2negrDywo3R6vj8np5K3ZHF5bu9Qywly02nAR0fVUB
HcRKXal47m8jsVYS+T9DVANIB7Rhhkj+rT3+HVPUVk9D+U97BERG9GURYmkdGMau
b5MjlRzDaaeLCXa+fpPdH/R3iPODQdDiVRbCl8UNshdeROQTMAEdO0+fc8f2bmAt
yBeBXGMifCXpYAcxgVNjkavkE7Qvt0ioFA1oxiuYzoJPTusiLCDg6AKh+0hUUfWb
7chgJPIWNYDfAxH0IbgWsuD0rJIM46s9FaQ+9A+rFI91+CV8BnOukI9LrVMhA+Qj
Ap+TEj5ksoXTeJ873eNp5sALwnLfzGXp4S4P6fk08ydUygDrXD2yIy7lKS48zbBD
GzW7klZC9OU0VN0RLZlYUZ+I5Znm3610oaEkhqftYNSguGzjzinuNgjF2A6lSNvw
XvVRgS0LJslSPNWEjDETxayl4ruL96nYQDax6IGctUloJ5nfncuDDecmltA3sX9q
a2RD7gFydooAKg9pgUV7tmJMClRSZscYW2J6ATtAXuGg4A650n7FkwuUFmPcW7+I
bXf0laOZvfjkBkzhsezpJ0DVv0l1cdt+kgRgXqJ5C0bJVInzxiC9GyPFF6B821zo
p3KdNQphabSO9LVMkIlO8iq8F4wIAXEICjPzd6vIvB8SJ/WqVXsX9YQ1XCUJSb+D
8jmpo3Di+ukeZuSF4Qtwp8sAt0dOYPrYbv/bYCaD+vQrcQq8ea+AlyRMzDukkXzr
E8mqVH6z1DQrou8sNgtx1DuOGxpEXqb6v/6qcN4pnR6bfZ8WVs9fu/zBP0aEvqAk
JTU9wOTfkUiLIJBRsSt2oey40fBS8Pq/t845yKHZt8STMESuGtc+eilchxmIv4/s
QffgIJu+KWrofViBxmlZ3Kg/bLFhLiCQe4QBIoMaCV2HTe4Ihx8F+jTqsxGuzRRO
fH0gmubzB1jwYURGnXlD4h+uzb9Eln5kPxONstvbY0ErcSDRuuCrnwonvlOgSTVE
39ucuqZ1yTdIKIWzaX47Vinz56vtWCvv+8dJ6kwH8P35Egf57lgyOwiNiAAiToPB
sSsKjTpCPFIAhHSZqyxWsg//d/s+qlRFeUcGO6dTQkzjqhvU+upIkcpyzubz9eUW
Lr5cX1RYpr8vOzpzBFZ2vapVlpN3WYp1mpJk8pTiiq320rlU+t11E86WPs7zSwY/
2smK2nxYQnuboR1eLrxPOPqDq+5m+y8q9U9KXgBouhqH6Lit7Lybf+TltNqeCSfc
30Yw91YCURukdy3u9VTFNWT09QDIcRSy+yVMzWhDsqveS/pCdRBkneD6DG1cgJky
WkgCTPwzq9sbgYdF0ictyptL/fPm+AsUh9K7W5Vpsolxb9/6XK2X/F8UHjqwEYS5
jCu60bM98rXTMWmCx6BOnMnQnx9DS6sGG0jnuRYnTM2h9x9+xmpqLBYblchHQt4m
j59a+Z1iz6WwXioEpwIap4qBDOZjkCQk06QeK2oxBUN33qEJhFDdNDHsz57TAeGk
M8E6+xAD8ugPFbVSeM9F5ocn2JTtTksHamOfTYd4V5a1KbSAkflitH/Mov4zV19Q
p67BFu5/SBLbl7t2WN8oxRDgSTetWg2MFvJVIz/Cp/h+Yze0V6mKCpQRn9QvmMOM
OKyG12HT9Ep4LFav2foawKcGc7vQEKNIAM/bZPNVJHBM1XTk97sfbDhzhOt+A8cG
PfYyaCD7Wv5jdb6GZH09lfhh5eZucFVWSbGtx3ed6gjciKCq6G0CgCWYIw/l5lYl
nULR9GGPMqfqvDE4vrWyDwR0WIjmGdILZcio0JXXu+rNycq08T5mf/Dl9Qm6BaUN
+OwYGris1DbkocNsTcBlLO8TM09wKJsKKv+PWuaLSZWDOLj5Z2hLw7rpa/IXOJsl
zPUDuXY5COA1eA4UwZHh4iKC2j7/o+zr9TEybKG28w+F+Ck1IMJM1Td74ouYhaIi
ZYoYG/Biw/HzI0UDvThUmug6wK+l6UUymNqkupCF2zGX7fXWIz/hA5DZkvVaMjre
VLHu3PpzvpkM9gcCn8VQ7xiZZfVMbbTnieM3BaSOAte9/fxw4cd8wu1UTUXjjele
7lQBOux7UOVz082aPdWiwWK1+T+6UGtky1Qb7b0AXWPQjWtIfTzsZo9JBAyyNTve
vHZFFbvlmrLccraYT0Na1riExruRLx48xWPwSlBi1Oc+DAuBH2XH9Xeon1s1/4os
LpbAWVYka/NkfEfEc9J9HMC52m7b1wJaTaHn6lnML+qzG/ZVMURF6cxLXT6X2KzX
Ld94glSgbuup52Jfuh7eKowFRce4KV8yyl/Um3IBEZpZNbbumcmpvMVyhIlJnlWa
C3Uv3qFH0k+CDLHbnkhrhXqasEfAoXTe5GwSh9KhJAKE+F8/Udu+YbafgFgVT0tt
+bG5D38TuEstrciPB5boBtcSDbW8oP3qIt914cNnYe3748CKldaWSwrr3EGGXS+q
fXylTMH3xnPDTEFPfiwjYCvfHn06kHQKQQMhx3zVCZh7wbXv0Ntx2sBUGVANzkWM
Xr9CcVqICwmq5u6GZS/ExutwSVOPUj5q7r9WhqFO0iQmYKj2jVdlYJGwgU1Bcdy2
W3ljnG8LGdj8kpYrcJ+/OcSAVufpRq7nXtyoptEHcs2m7nQNibnKFDGazjLrC0+h
qVgQ82dURMxNgHAbGYFABrnPUCuyvkeZUmwnsSDJut2NcV/PwDs7MaKBn3Wn5DDR
MTy2+5yjAwphybQOoBwJM+oGCUqJyAqVnKHI6qBN638byneIIQ8ToYRnKZrQmiv0
ZxF+rTEYQQMRoDkgYhErTOERQi/wxe4DFoXtNAaniLpfplvurJq4+DmGuiwHyaLu
OyVM5rTwW7lsB+OQURuQDczwYKoYWnt4bAijdqwbtC08lkkt2mUgmHyJZ/Aak/OI
wCdGeJIZmR+sc/df2EbNZVcQvGJ2yN8GYbLqLhpAITOeVogIeozIa5qKl2UhhpRo
AtnqXAqv93HRKAacKW6NUBKRPb0B6pzgBnKSkTXC+tPoCEz/HAkEYJCxoDfwh/mD
Ezyk6Vlsd5LDo0jd08AY1q2Go0nVaG6wP9DRlN9X7Ryy5Z1AjaBqMKEdB0JerpPH
84nsZA/riGCUFMr1X2A1jwZR51RoaJP5RkypVjUhVUlW3FUOPCTuLHJKb055Bb5C
RC4p3OEi2xNHyF5g4K9dzj4mtULYJa+KIDqdmKff4OJ5UfLoYbJBHS3XxbF6nMbd
6TTUeMa7wSOtIaEHD+NJrcbDYil+xKpf452jgFTWsw0GVok4OmpK0saV6RsV27yg
bHhf1aBPpiVfrKc3nI6fwLICLPp9XmOZ1VTQmjLIJbI2KNSBbsdrZP8fGcSMtFyv
E00VFvhpjJDO5WWIJ09PPWtQT4WIQYXi4VGGQ9dmzn0HDey3dp8ZiZHfHw5ePV0Q
lKw1AxCkq0MQZZ5pygV8ss86Avz9OA5S5jtbLECxDK/Uono6kNMcq+VZT8mu9Vks
lFQ6xrx+0BAuX1wMNXnsz543yeitnpSk9Qj5RoQ++MvIoL8UOe2t1wn+QTggKJV2
lvfvGIIW1EqwwIYO9My1IeMieelF0ABXli9Pb89U25ildK0q6wOg56g3tDpJJsXy
iaOU2Gmslk8TWNuFnZMuIF8N18AJkh4Vr0Z0JIa2UylZuD8MWVV8NnZT/9Z6naGT
uK/sbixPj7S+cvC6bOGzZZLFH1RHt5ClZIP5Qp/zLzTQXYfXmUQND/uZAhwgjoeW
V8MEMZHJDV0/Uy4Enon3v2rTAP4hfwBQl8zO+beiaC3C4n/1xsj4aH2X50N2wtXj
ElTSqoGmDiQbn1CT/4Ogm23xPaGWEnBK/wXUz/ajMftJylYGq19484Nyq7Vbg+Tt
AGqUm3zZrK/wS3qnm6IyUBT/6lq5uaAy5Tg6p64d7ce7SXwzGlzRiQtoF/6s9A5l
TSNh8/RZ61LpwOZF8nvKVWNGfxSpTzvL9W2kYR0JGlZWIgasQlL5YqDi3G+CMlFh
vECxFyfMq8YSUiVsAVSK9nrXy5bRxdzTX3Yx+vnaGtSQI5U4ugO4LNj1gPLpwCTP
VlElIe9wEZ/mCall6VE25I0yq12CdtK87JsXKUG6/zMA8bL0jL30mzcudiNzRqAI
PkVnFBB0qxL/VW6wdUuubo1U/T4rGWHzjXTBq1M+RzamFDnp242CQulMgi7NZA2A
Uks1YodlycNz7Xhvxe1DSdQBFnrPVPtp9gZeTIFaR0vJqXstJytESRNjB7ypDkfT
BkjAUbSbDl5e3nysrgA0bg9k1D5sxWgLJUEH4C5rl369FsqRcH1y+TYlRAUoDDik
vZPveXqHiyO3Z7aUhx5T52yC3/dgGDeO/N3LNSlQNF5pJ+4hQ1z5MdsIeSbrsiD7
isLkpVJ6TjODQpM4aO1A2lTY21VuKJ/cx4QwCVA/hr04I9BcJoD/Yq/o1566rY5h
IUXyTNXsd8LgyK01ayffHVLCQaJi/FpUXQByNmSC+/+BO/ZGaCRu8DIDa4r9DMTa
7NrigVpwScIqFgCaAlaePcVzjPCmfCi9QSIh1wJx3RxYEBuZ8LdDnCJkeCdmn7d/
xR31SEuXQ6M5I+w99R9S/sCwTmdIXjSBI/POAy9cliBYOytn3Ps3a08KIUj7FTEx
tqGTei09REcc+1ONeKF8ygWmkGfWRsFY4QViro7tSARSw3xELmYuq6p6ghw1wqy+
DAgGgAvHVxhQrUXY7RXblEtqKvFuZKZfLI19Oa2HVmzTxjoX1seq0ums7VZGFMrx
N7LmxVNXXDX8QgAEkfzeOvs4rLm+kj7j1AXJClflx0lOy3Egh8M9cUZcIQ3b3ASA
aS+5+6Z655HrjDCAMKQJj1C65ptT9Ft6haUxShLYSWU50wFxXpAVqmhAnNJQCJoy
bXgBpS5DM0St7yNkyO8Rd9ZIc0iBALMZCIShHs7+H/PuboFzfCOZrwOkZrPBvAq0
aIb7V2MpH5bAZSuj2BhWkQazU6smZS788esD2Anl0cPMFfVKa3HO+vEEYQ0WuTXE
fs083H92dVaLSFhgIjrFfNbubKxXNIcXI3OmSrqQMufZ0/zALdqolgNO8SsuASpp
Qu42MDtzknAbm6HgQa45/f6B9MzFZeEbPpYISw1o9qLH7Jyz1AxLAhk4NIPYbAPc
kat9an/2m00EkwU2VoZB8P+fZvTwh/Z/XLZhjqaZFXBOquRv9e1VN+PDgpghfv1b
KNQp9N88Q1X5SSfm2aURWyYcryIAZWhP42aRtM3v7Gsa4OMM1YDP7G2p1+oC0Ktq
pxdbeNf3VWAeOhmcAImx8soqQ8z3hjegdOuPCUkmf8v6+7jXJ5yLfy9wPAi04SZD
aLuA+HA8KoiPND/2wuUpK9fYBq2T0kdwmpomNBATXphv1hrlQAe3Izqn4hPqh2or
iRlMMJT1AklpCkcFStkERVaxZBgopRtxADP5IfRkZd2xnPr8Ooxix3vWsabAPFPY
DvHd983k2/DLR1C6AJtuRHjnjXY7X/9Pag/O35pEGw2pCtpzOmR9rDX/SjRlLM+Z
ZJecpXl8OmAmRxx9wCl16UrB6xAGbCcrRZZ7wu9Qr0/i/naCzNGvflNtZaxBuKcc
U+vQ/ZkHmD5P4hKd2hrFYRhkgQ/jee3p4cnbjb7DsEDZcf+qceFFX6tI9GbYtWhF
Igl1nm+RUZLhTjoNV4rJisj6rgOuep0NYjBy/4kqNZjKjHnVfLfcYCdbyX87JzeA
yiK+Z/lGxGcGYycRj6Wqaubt91V0Vg+j/sErdWQGoNNypsR7ok4O1Ye/XhTQZ75O
RcF2QR8x+66VYbNpwPWN8vs6j+hX/Zal1Ve9JGh0zWtY3Lu+6585hPCvY7scLTD6
LZayEAktziHrQYqG/WbZplxRhKh3IdRe7k9Mxv1P6kil8I//zsYe7RhpV1iSvRZq
GL6Nzx+/cGKqE8+LbKrq7+I6aISFVms2Njfc4KcWNf7ZDSbJhr6wfHHz2z2k2h2A
u5g0Kq/60PeDqbDaY6WtNW5kdYqHkdf8r15neZNIjiFedjtCLwlB8USeDnriawdP
L5MKx1K8VJCdywgWYL1z7V58S7LhQu72cKtRxS9DgJ09ukZVsd5WZGVjWuLwlIWc
KCQJ1qDEmbRFVmERvyL8znZ1O1vzMHawyof+iqrmIYVdV93KlQjxph0dGBSa5MKr
NCJQx4maL7gxebrtyKDLEwzGdd2ge31tS0L/wJ23K+35dgxJSRd4lOyDyUitKnoL
4iFRcqSJ1qhe48zDnwM6vMgy/aQbDHAY7lsPZy33NekZbf78asDExM3DtlUL1OAn
WJqSsXxuA/+oYEPjlSBZbkBdwNJ3CRW2GraNqEzaoff9R2V8levrAPgUeFLGHRJG
6Gpmv52EXx/HeDo9AqhsJ5lWBfTL4qplhoVslKLXCouID+jtYCMSm2bkscVXGFDk
iVLbJd7Bqo1tnwLbRdcNV4S+HBODHla6ZGOmB37GaT9QCHejOHkj5qfur+RF4Zqt
s6mMCfZWeAaAA+ISE0E4eVLZA1844KwArHZiOxzbNy352sxszFKwWBHgxOatUUpI
GYry77ErhwtGVrg8ckNvxgY6flawapAr4SVMeZljiiqaxnIRFmaUdPaERBvU3R4R
OL3dBPJEkPPX+b9sM4KYzm0WBD4TH/WmttwlcmPuqIeAsh9+HUpZ19LWuAWmBSEX
95FTwLoWzaTw8SrlJYRH3JLihlM4dnJNlQ6hPpxxWOcnqliUJD09qmdAgJoR/qIs
MPXDibc007SDKzHVjnXRIvpI1Qov+n7hdq11YJdxsrVYZH2+tFZPukd+7qeAQX5R
zFlpQyTVZhd7NQZljWzO7HYyRLEXqVddcOgW832fus9M2aydM2qYmS1COreJmEEZ
TCLOy1krT7fVQWwhdlyRMKs7+4r2iDkxH71laN5iPdXQqJeiVqM8wBU+UFiRsBrG
hiMH2OacAa2fWauBMDQaX7ILNp0lqzjUqnwW1HAJjElbrcqNhOTPHQRCsQgGSMi0
bFAbHGqgW3jYbU+1kqicuZ3BsHqd1KhSBjOY6QQc/u1hVzLomFbLUVRWejdEo83l
b93JALywCVXCZHIheIzba/1udVWQ2BCr1TMeSGjWGgFAmCgRgjtqZS/gyRVKpI26
yWvs5KjwzZG3I7FLmK2BRPeeRVl3t/yj725S8U51yhlwO7ETVlLlM3XHzpw5rfOq
9Mq9NWHFossv31lluQ24mnLiVBl6mXIa/eYlEEa0wk+7Nac5vHzGBULN10Dzkahr
skkPEv2qM5B4YFaDbv/iG9ReVQryGwNrT++dmjnbKW8heW5kThCyq9CDLBc1ECyV
J74oG4LnsbjJfj9Zvx1eHYOkHlB89lP8mKA3YOCKIFU1nvVWwT0YrQk6Ok8nhPwz
R+Nj1yuAVRzPSehzfemFh0g0elupTp5e1KfljBWFYtchxVToxLkqmzx3PRPMdgrD
jyXBJBJhvCPkTZ10MjIn4ty4iLJXO1mj/oSeC6AeN7dEwiUmGQMDF+GiVx1fkQAB
D3o76irl2HC4nl94VCNZ+jiFTKBXhsVJfnh0PkYbiZ8hRcWqUDecjEx0+auRV6LI
htTpaRQOGeYrq4iqIVdjxNAoHzu4CjQI18V5eD2sQcEMv0G/0XWLgACByjwDOm2Q
H94QM1mO/D8SOH5BcZl0qWsygUfwoAZ7HqO1ysKHnBdKTYRJIzk0VYApYiBY5S0J
alNV+XCSxMeEwH01KNcYicr/GFrIYn6uKZLQs+idX2xVZQorVZLZiy+8GnCYphxR
heWBvpPcqTGA1ejRAYs0aF/SJjH++haaXYjXqCCJn3zL0OXIJONOkyeh3NTbeygH
bmRMJWsiTYTvKsIpGPA5JTDWQ/r88wFQ3q7UN/RUWYhp1WLqAWeC8tk7leBUiY4u
GZSKPgyItrZaUdzDz4p2UVFKTJdJB0E5EkXchT0c4Bsva0o1Gc4YLU5wHJPhL6EB
8s1j9mrEN+grD2FQCOjO0P8V2j9wPPJbrjOko4bx6WgFWitd6ngviIW/Iwtp6v/t
pqMXdUnSVBATxXSOZmmnncDQyTKfd9ApJ0MsX9hbHyPXSMYW4By9ubKfbBkm50iu
hKm5T9Q2KZM/HN/ex0VuG0BnBLf+FGyL2f5Wc3vqzwyVDOrCsZ0nNg1tA9o2zuny
gi42PRNKVHaUts8wurBWIzxFFsb3XF+dCbkC5d2jqG3CWb1oG+SdIP62A9kJBD9n
2JVm92csq/9fXYOGko4F0rJOMSCWTmf7wmtHKAmZERmIqSv9HiOtTsRfyRHQsfhG
y0vZPu0OAMYj06hflnoW5um8QO3f3NiW1a46ruuIkD7ECWMTWt5GU6gsXAwpPqCc
8BTvmiSfcGZqn1dIt0iWOiALxld+49Fue9m7bXbY7i6NHL5V0SuZVYkLbj0sczSG
eu3xoVnAEKzWaSfjXl106y/ThrvMvx6sxQKIQRR3h6HgJaHGoWuPNzw1nzSBFUvX
moFAx6QkuBmaQusXThN3tInU6vpsIf/sK+fQqgKo1Xug3tZdTyPYV+ukAZZepEoy
4ftMHiCSz5Q6/qIbnJTyUfIByqMlNWgJsJoaw4QivFJZ5waxMUkw8K0qil6qEj/K
C6y9SonkJYNtLyxEVfccBvGLx3H7DMKgCbC/95Umh3BGlQ1gcAVy7LAdiddccf1e
ijb1Ei4pEOG3HqFe8r4zLkdZfDKlav8OXdhN8TWMSh3vJsVBkSKZqms0skM4rs/B
zbulovYxSXCPKoqkDrzm4Wu4YLqX3wG9c8iDXvrVALmMZ2jaGL1sJQccD7mVLvX4
74D0QJFl0PwTxdwAZzHC//gdOI+ig81EkFVjrGN8Uop1gzm8gxBVcJtz5ziAkzOR
0VPaFtq1doKb61FBKPwbkMOxm56M1OzThZhpIlySK/dfWsBedvG4Zp4FtRCVcbTP
g7xBMU8v4bHwOy1unxbfLrykyjGuquJ+qC33fQ6fFjdBHy2Wvm63NDEe8Xju74IC
dPL+/O/HMgKjMbrGY9YzNNisNyjHXKUeQFagpO8XzIe9zodIGuuOKgaOo12cfz0V
J8wzC+JE3HxORx3+vEK3YZDHNmWG4JAMicpuCYk6VszqtyNPBlc2jvtq9oESQe4c
NuXv+cz1A0wm3M7hNXCTJHsUXxidfA4Hc6j9dWAVcyoeLjSYSz3bSfTFZuNZSHRk
hE/8bQKijlaMwQvl3BvFoxojsN7DO+6yAnhDKiWo1no2fxm8Y8/NNfmyU8uwNeXq
n3SX3zfSiTP1yB4nlcLEBXEvQ+Gc93EkRHZS4AeSlmLK8vFS2nnRFBGq3c7M8+Ev
6OhZXi/S6trNYZDQnONRysS3uUkXQ2fGVL9TkAp5bVgJUTLb/cQJhQxGDddt5Ocp
OVb1jMLSFXF/abBVme70XtquE/yv8y3LAivWMl/DSLArGwtiMZovgKQYX1+9unR/
cINVHfVaPoM8w6PdcgsMJCs97VZ77kVY8dkJyPc9GTCMnCh1+y+AfHEQvlR0VBdz
GY0/pQDkAn5V5phxQnRiSBdlnzLxjFyro6X94XgRrUnvrJ68F7a3By23rSkEjZyZ
QTJpy1BraF6xHXzP3mWYwJOw/+n4RR8eRhBRHGtEpQjdyx5Be1CMT0aLYU9GDkYL
uauQibKNzATPofpn2PGpJQfqMT6A6x/SxvZ9swFZLA/NmrE9zQ4zFPUS4aSpBHFB
7j7cSJTPuhssF8Bha0xFJAcBI1IM8DNWvazTIrtPQL0vZWm6bv+jH+1HeoRqIuQy
XrZd2p4lQ1Ed4oG9HglPUsM+vbjrfYVvYWYyd2x2HLeTtjE40jwER00bnvtmCCHm
c7xzxWS68jJZJXoPt72vuf305lfYUGsxBNBKTyaYUH+UIPjvzoTPFAUXREdpTudT
gSMtXK2roDSI3UQWHYsUvnDiJjoC+dcHopU4fwEVCoOXd8dtZeW/LU/76zZfIxDz
d1sy8nnjiDR929Zf8yjOnulF4jTTfZWzP+aafSIiuHsp9L2FxqxfKWcPptQV/XyE
wkYIrVpMtUjFHfzogGUwnaxuzdVrAOWpNuuZ6/dLNuwkaCn2m2Z9h7GfiDUEMlp3
okam0d82B03xBUMfglK7uEjg/URI5qCOrSGQ8VSudtCUYWYEpL5vuRcbjFIVRTLy
ygx6vUrGzknFBOcDE4BAx+qzCvxpCjskt9Gtm9h5z1NMmwQ2xrYBYl9AysPZagiz
5azO1G1wnJFSlnaJgQKHW1X5UmUN5Rl8pVe5/UFWN/plQomNkDcGzQgCqNP6CLdt
T3MCbXhfTvhEjn7GjRPn+dvT/SpFJ7xGpbJ7B+okyfdQCRadwTVgdk6Wax6mrbe1
8LtQe/n+6ASrKgi5PE78d1xyHie/+Y7laUGclg1g/HQaSnGBxGffbEV+D4DgnYMP
PWGKp1ljn1bw+RBQIdVV7IIhVo+lLxSYI6GufdYa+Y4ELdiZyUGzp6y10tSh/A3G
SC6zaRbUwgidoqLSKe1uKBjPgcyrEAf+lYec7Fryj3OQHO36CtAYdlP3khtnkvay
NIJR5JppaE/sOSZ9KNZINAb2yosCnxRafNNuRXLZmgXC/meSyGpvEnA+lXh83T29
KLKh6MIJL+AUUiuYQvWwkPCPL7TbMmtulj8bivCs2YOsvmqEH4yL1/9+ZWfrdtZE
hpNSAh47vMPEZoeN2BApOzNpJ39BUGOzLQUFmkG/2ZFrLBnuY7rM9GuQIXF4IWXw
rzXeP10V9f3z+C5DZv3l/FSgHTtYs1JJz5Sw7pgIMm94P0zhG5+mkxenKYuH7pL/
i7x/PhsJCXcwNFBsGVOyrscDgktNgN+62YOODH/j7RScSfpT7X4jY4weaTd/5LHv
ieII9DqcmDRTwb/T4yiRpVT1puR2dy81rROUWN4mFJnI4MyBcSe6p9fpnuQpmEKG
cSuwGzrFTwz2ZMjso/W/5c5SQN9guvGmO0n7+En2Rqr60wHlqs5ChxGA+hSyB1oE
UIZdSPsZfVCezx6pVVi3i9bmc0/Y553YUiXZXYXAJfydMiNaieeEAew+CQaNHzeQ
61aS8UA5YLXzUtmpX6dnzoWObsA7+ZPCfdRO8CAM1VNYok5mVs0ekwtILn+XxT2M
wXM5nn0JjZfiymNWJc/AlUQ9R2u8G8i0kv3IhpdEWuD1rpHEtxzkHyXGt6ocBvih
v/J6VvCu8vRtGLfL6CjUDAoq8xMvv1MxSWnvohOYwwTUhd9kn1wKClwwTqpuzBeH
85ky0nRIgTkRZ3on9yMxmaJi9UgZc5iWG0Y6h6BydHq/R7sFPE6/rq/XikYwy3hi
HVQi/JN+AEaVonA7CTByRjd7X3OaOYLhgTbe/nkrOQZy2OwLf3rI21Z1uGdhiHyq
KY3JjX2xOFNZNClrTpI0qus1RE/Gt24cTU04ULudA/CxhS4TsQl3oZDcvYjh+B8F
ve5bxpuZJWzPUjUlTfCaVE/5kyJUk1ytLxw6ZwtFDPq8icpPCUjsatmx8WA0DfXS
UbbMDEXC4d0eWts59ku3GoLz0r1u2D03mIU1FrkU2uBP4ua//W812NdQmiJy+MWD
wh9LV55C6asIm3oyH7yOtC1EQWoYA+Qz5sTPNzYtbH9FbCGBynKW+LHPSv4m5lLS
S7FV5ougNM3eRaVcH49gKPZ+Kjg0B1WtrQyZJhWuEoaFOrujF+Saa50xGNHKrvVj
1hbj/94Z4L2hQ7QbFKpFKPg9HPJbffSXb+XZS5Xpek+lVkSo7zT/AgkSv1JEUmvD
lmigwK5f+bsDK3dfCwmwfFokjX8WD1Y5El2KVtfhbFPfzy4ypMV3RU9g/GK4cEcV
To/dgiVzWDXwCoDwoZqocrtWGcgPGjKLjEo4Q1dkIjs7S59SQDwJA6CKp2q/pU35
/6AmQhjqYDxEBqYxIVkcdPB4XKcEFVoQr0B5mGhp2Xk1xlupqi/w/zZBEIcPR/jK
rfXwORBHBg2GnU7mfxSzMCIVHBcmHi/qjt/xmjhjIOUSpzFHeUzF2VwNfyan54cc
rv4Q2wMiSOqytfxioYqDUrjrlrEP+hp3jZdldIkOY5Vf2PD7NqOJwbbB3EqaiSK0
k4AAnWvdtL4LwhS1RBZn5ZFioU0Y5vSxHBWVG5LH5CWQsxluC2d+tEza+jODitoy
2gAB5qa1CCde7uoeSAVjbpRylZDeMOhCjOVrH3nlwxCA8GhXvqXrH0ccYz1MmG0s
bmqv9uaofL8KVIGZSICQteiTG+geIHvlxNq1ILP35y77CFfSvf95XEhLY16LRnPQ
iXonUjn0apaSRczWtl7bRBZKrVTshpJ3IpfXmtkZ5TfDFMi3XXtcQfzeE+ga+565
l873zbHyBtRbp+V3+ayVsHRfyVi0T2JFqPgkjNW3fHAZFea3Ih+WM6L/44tWbCht
JLthTBGtotJyCg25cKyf4U0P4oOPwXIDyXpYCJQ8pTXq7Vr4E/iT0na/JCPIb1Rg
Z70lfvPvSgoaq0BBzPhsm05x9TqZPHw+Y1QYmvdKIOFzg8tvLmhNpYoF0mCze58y
idifck2BMbeWZyRxRGGb8q3Mf0kuycyq2zNelbsiffeAlnSK3DUfzRYHKjtsIUL9
3Gm6eajxnGzvqjjCRPopkIY6aKV/k7biFdg7QfEHX6NDTAMIwkH7dWk8KAvpO4Ry
HUfsY4j7K+Hx07tbDuAzp5MS+Gc1VL1DVssqHzDahm3A1DPW1Lf4u0e31YlG/j+E
uKSrmYWW22flpLWmOHOlbZn6hmE6Nij7MpjEiENyxlXnZ86IjKeRnXihXJ4b6vX6
jglqo5+BgS1LGCpRmvGTL/mHksVBZFeSjBYCW+hNDzI+34CRFT3CK9VT+pzQWI2X
rr+dFAGqfbngTN/XtjG0jekEpB87GWep/n1EOEfOePIOTc96WVGisht/7lsZVFqu
DKbXPaGCxH8JhggDP20ptH/6nCC0R4tma4jjj0H8V3OMdFK2oSPPTtS7vHI+JtoK
U1F6/ogSBETP/c5NlydD5x8oaJAuZ3d7eDnBTbbkHW2x5lACyGX3vx1JrlviaQug
uvIgjRVvf4iiNBKS3WqV9WRgF5qM7ez8q7+UbJIp3WbEz6UwtmaMncYAQFrXO7G7
a2F02m9mJbgj4y1eXGK7WJRAo+VHlFPhq80W4dJ3bO8STaLK3jVySi7LGFyw60AJ
m8HjZC8l08QKFoQ1spxkQxTnwwZgErciBQh3zxvxJJIdz2d02iDUOpeHvCCiSUOX
d7K0RRhT25G3H8zxRuE5w7blJfUeswu3ofMmnOq3gIIpmJhsTdDOnCX/bjlTsI1r
fwDOqpzXw1ym6GccJBhwJh7KSGAMwEMHUet+4oFJgXPOL5gQ5Eth9T+FpdFpkJ9G
llFkBoRqQUoB0M0z7dc+RT4dbrtgGA5zM7lt8ukG2P87buD7xvvKmwuXF29xROgh
phHbqumwDKPICPCE6K5ED7R3rlBGeS53R70m0PpVZ0oV2kW7wM5xukI0+3YwLznt
QuUIzzvZuhRuTZwtxq/vhT5AHlfd7JBleQqQR3gNy87xnhkc1t/bBSRIrHx5g0QW
L9aVR8xO5nu5YC8j052+aJcVJvHm4t4/bfUbl3xDG0ZcFCS7SB7UN1U6B4Z8X67S
4piaBqckeWo/FiiJe9TEO+Lb0kPYHCIROCYcigewaE+e9R4REYcqrXnRgSFQIOAZ
HbpJnNzJ5p+OErFtFNmmkayKt3s/yMb98JbPUNQHguRL8S6vsBdNeo6JwGQpuVcE
gi5pTZmh0gjBRpG4Vp30F32gkWLI70osqlW8WWk4MDVXw2w1sYSRbK2JKS8iBPto
/jkPOoMBSvlHx0de4tySOnR6bBYqi/cLIZOvkyQ5BP5cVKQK9Zx8PH21ecEoNgLl
d8E1eTMPa8LfbvM1GpVFgEoGkDHg+blmZOHvoAhUn5bFejRlE/auC0qBzz3F2hbq
MazRlYdBnfl63xJg0j/n4AaxVh3IP/yGhhhKMuXOLOEQL5vSzYn1ylAjzNcyAIeh
2E2KKZwfON8Zfz4yDNSRcs6hZN2OJ/k6g+MmL4UnsecGyPBPiEWQ0jGBsqu+dIqq
TA2Q3CZ6nSzVPY0kZDRNBGZpw0T5uT16KbcYc4dec5M9bAp2x/WNDt6QQ6Mo0525
BBQRuJDPQbR3TQriccdrmH63SiewepHplh1IB0eXfvNBDSxPYttI5fC/oPhgeufJ
0aIvoEJaK7YffYP8NJ+h9kmrDZNlLE7QdF1qznhiHKL2P2KcpNMVhw1F5hSWE04K
a5m6Ku9By47gV8al804+ZBV8Wlt78LZzpi3BGI/He3LHggZDz7tRy7Dx7m1k2bsX
AnK+vZu0m/D5M0TRReaLTiP7I1PbSKejLA07maBQqjpkep4dVU2DjWhF0oGqO3YU
K66UWpI5Zn0jiDj1UztKtOsgT+yRAyEDU+Y2Ja1U7Z45xmQdKfy+Y6Qr10HxgaVH
EZ1br6N1AGuSklFZIw02AwQQyukBWNzrkSoSMCRiJ/pXY8A14dmKmms6o/55vec5
saIHLjjo0Ky23ors+7cC9FqSSt+GW+zU6dypCJHAnUGo5V24jEtoQBxAwA/Q9BVX
8YhwhvOMy8X2OnzDtkDRAFCkJW6BcCC93ZNpouOxoCysWgmEjb0VXeu11OBb9MdW
LEROY6exn+ZxrwktW1azhvoMWiVBIfhMC/d4d9DhqgQOxaEGMvMdrYRSjPh5uKi8
NzrpzIKrHN26dN5QEVGDEDsNDTc+KFiMZUvgYEWFmyA9z7G/798mNjlLbgAx1sMc
1ufREsSCvADyb37K7eJHRb/NTiHhetVi+ewSLp+iXd96M7fwUYYoWDSvyj3j4TDU
yGT7ns0uH4Jg5qcIjY9EsohdX2vl+MXCOMw/2Wf+PUmc75IIGLlTwKQw03JjjWsW
37sXZbLpa3YetMabAf0vCA9ccU3dsJGIqa84YxmLq5DWPnVkU48sNmZyfRe/R4RA
NiAM+G1p49ENcLpIhLHzw7Lrr/U/+Jzb5QrY442amKylgSYYzoIHCjXREQbx59I2
jy7PsjqC9dV/3mzDrFU0FnV9XslgbM5HkEoYNzcqDsCWkN4p9ogkCimjIUr8ctZ/
7OLW62RWeMq4izWd7oC4kE3syeMvCX6Sqh4z941AL6BrQ/m1e30zEL1+AndgIpPH
5ljcyFsu7ZQriksYVqi6KcuDn2QHRAn4yqljD9OWjmBrgIBtnV7UBxzWjXvOoOmV
N1eDCk1RwO/mCgA3zphug6zFWQAmYD01A5iST0EqmFnzls+XTCDoQOyx5rhnYxUv
pCPtPAgXZGL5ZeE7yG4Rhp4B7ovgOFC/gBcZPH4g31qgDdOhL+bDBIp6VAk3vyAq
yrAEjl9JtwagqbbFZa/mAJDH0fjJFdZHBS060EN4/RgUPwVwrZwD225YABk9timf
oWNvZmHa23+AdJMs5hBQw/XWmtYhx6Y4pwzkpQSW9/mtk+mBfFb+M3p1uNooYKj0
0AsjtnaUQMe1WX3IySd/rbzsvwV8D4Sr6FsRnXaH3zkUky1tUt7gZry3qJGKlmbr
wk1UJ5c9YXb8mF+2d/KhBrw90NkVzeUlGs/U4WU/4s/6Q0vKuixya8O+AVXJBCTO
tCnVixE/IZxk9XVX0oBeQMdFDr6HRsdNln+uXwGSgj/cDobkgar7O1xVqQ7/DrQj
Qodjdzql+uHxaMimUoPAw3n8gNzkU6nUr4rK2W8RPlucj/LadcyD/TdHkKmrEVXX
7fJPQr02ocofHk650GHJtmQBk6EPiz3p8UldsuPOFyyzORfq2xOj3V9cgrtlervw
9ItjXwFQmDm1vKdUYsEia9PyAabdMNTxGqgQhasrzEqSulJcOFyuihywYYi5Nyb/
zjF89MIedNidW1mGdTtJX6FuAHJ+e87fIdxdZRWJfqEIH3oA3bg6I7Ibbf5hMi6N
zLI8/pbdntIkA+Lfs+rV9QcSLxfJW0eULUihZlhg47IkT+U7FuPF3y40dD5aDWd8
embyUvf1v8AsOxfW90an0eMJZbTQW/6AVwEN+OXNaCLhlPkqH3xnkf5VXfizQYC7
+nkvRTQiNElX6J/tM0yBw1/xbvglHfKrfme6fsrmuVgk0xNPypZFZ6G4tFrasCPc
VsKZydrHP6VQaXFly/imC73AKc6xgsRf3WuJqadbSKaiaKcqV+QqWrgTq4rQlUV+
43aRuH2Ybdw+w+qa7B+hQEWBvRG9soopQ5C8cqrp+r6PFZ41xlyoEmdvu5mZIEzX
ZEj+Z4Zd0f6l7GTtrY55RT+Q9Ch6gq63I9NI06MxHT6Ohet5eTPzXS1F/fWg1gDI
m9qChw38H8btsiAJXuLSH0ccurY9JW0/dZl9+i5ZYQlnQQdQsTNEbKTRGCs4pJmJ
nmZwYaQ8qeeJ7JzShIeRtf8waLAEXjEjA4pfF/As8B4F0DYByaC3BP3riFeGPazN
0opxtyKf79NXpcOnw0lOZKPtFA1QQPe4IRxtDDOT0E8uSXQcQ4+X1lWjz5VUwuh6
/HYoCqdxqnzbvAeCWNLOS7WSQj6NbJCo9jyfDRHConLOBS1BpwHLmeJNirKWRd4c
4nQ2aoKV0yLF9O8bYG5Qsq0mTg0Eqx2WRMBvO7jtzPmDy28EFrflEi5Zj4k2vCq7
3NRpZF8PoaSX8IXF4RPAVFEkscdLSZvTGqLp1dT+QD8PhO/P3AfRqEA9DzK1XpU/
pRZCD/1Cd7AnJqKBIeap2tkNBkcAdUZl6Nkku0M7PalFDAh0pJRSUGGCKVaXxGXY
/gSA/Trya+LFWKMIXXqvTHgPhSdynuDcjBgjbmcz9m7EZvPodEkks9SXUS2AcxY4
lX/MXAhy/Z+Hlmg/6V7kHet+auUFzNZODA3i0f8AvujTDgniRjKo14AYAHIrwHAj
RlgVciR3Gbv3ayfSygETv+UAOJ9TWyYqzOj5mDm7UhnpTEO1b5ekTgqy2CxyBgQS
Q/i2VSc5xgfm/YPBWoHuDuIZDeq2Y+fuAOrj6IWUPHlahyYZvqY+BcxbqVD8BzVC
uXQ1swgf+T83nUux1prCQMh2ZvdAQx+YyLmWZod9vFMew3Ov4vaI/Pga1e36vDUE
z/UTNbff61PFcVuGFcY/5nIMRYOjppPVOon8c9uOgacHDS7n/beCzgVh5bsD6kdu
t9QbXpjZ3QIB+ctDkS+AKBsnULOwWprEjJXiVzFY0jEVM/NY5xrZ5VwhvxeX5hgF
TFPgeY4qPVxEWp/uW1UMlN36bqfuAeNg7g/r8IpZhdly3biiKg2vkW1V190i1ZZm
CwB/x5/1ZyN0KpWwpXe+GIOOg5ZR5a5Yaj/ujkHwK/Igsg29Ym3DK92vnzcVndNY
iv67W2WsYRMHWu2tsJBkSqGrbbUhO6uoDXB7WiPomd88RqeyiGb8WGkCZBiOWCYQ
Zyg07wnZ985/pEkreISC3fFG5n4xUAuxUcjbaESjDsirQdr2WB3OO+p5Oi1mnqHZ
nXrsb9OlicLbaf5I7SZlbmSTdLsHBy8lcz/m//B+GqdLU4yEanVo7No8WRrNbXlo
vvzQMC1jg/20lEwcLzcNzw9mzy5J2m5kiodpWlmK0t5NE5lgpHC5y1fIyooeyOuS
CPTtl6/UZtabQ68pubuGRBiHdLg58AOBLXNpIQUahaobsZmWskEpJwNcJXpX8NHC
N4c7/wQpzC+yO8X++G388bswg+lIBfdlzf67PRD10z4z9rlE57TjRQJ4206bwlPs
7HhGjGFm7ZrJilcSiaDN7ECPjpZBlmPKu/D5u4wIDtOXhOWECa3/nEGm7mYlYz82
+9jQfjIzNZRgClpv9yB4FiEfgcM1SDhU2gPpDLVv093ijWDxn4oFtAkma1EPz7uH
REPHTG9iR20A6OpdwZ9yDGIXFdB2BTOMmBXOyMYUEi45EnG69QaXhRYbN/rN0UM0
vl3nEzaygdJ+XFwllmXOs6yAuvjgeAQrT214zEKZdi/BA1445svpk++cMd3AvjHN
8CCxV3OV4euIKhgVHjN16x2r8W6uxoYPyo0Yda53sjgStJntzO0jQFUlD89alguP
vCJPQVzHwn+THPY9uodfZ//XWGLPxZpm6NtywfFQ7nfALeDrdyReB2IuxYtS7SkQ
vSQkd+++5osz0LIDx9TzvzbBCSOtp5ThjDo/OTbivNUDINJfR3gtnLh8y2/0fgx/
p3TMyKZ2PNziv9fdWkXVveA8rZ+IG3VnBxTVRFPdLRl5makMv/rH562KdoLayRiL
7jMC6KmQWIKfUu/jbBCtRpD0Vuu3svvqG5y0KVzOA8X2eYS1r5GgKZuOApkXJeQd
Ai2kwEydWoWDjX4fvR83+VF/Jh7FrsuXyHD6TkkGvplIizzLRrf1wBVmJXK4GwqL
W7B/pULTLNrWoiMwISFAULESUFBGwvVM1QWi4a1kpYS7NngwrMFy/Q1Wi0QYEZqQ
ePFDwT/Db/W2Qa79S/xCx1ISDxOToXOoWrSiKWZc4SQPh8cwqIHfmTMyiJm0abQQ
ctDFdh5mw5OHpVd0vcmlXKly+TGmri+kMmXdtIDrba7vg9A9UDmCA9TqYXganesk
5Ch+TrylDGlAiKzwQZetubK0Q57GtoXmCxr63CX8rRkVASVcV0BGqu5bC8KMYW3j
wmqUMxpWa6Ra4M2Ik6Xa4Qe2K+zr0P2e3XCqDMUK7LzSGVbq7vQKEmGKAOisekMk
S0GWLHTVo+8VLSG1yffKMd5RQSLuTHqgtTfvnOJDQAS2k4NzFPFk539eBJEtcX7R
3VEv6LLmNVmuiH+sRNBhSG0Tgp7AAZM61JijoZU1e0S8NwSpOmAXlT0byQ1FxOAe
4A9NM/2S44DUZN0xPN6rAXvoABJe35QcxHnbuu5vwlh42DBWteXNELq4nn5wlBmb
S1hO4GwIVpdj9N/C0OU8ivx2XTmhb69HAw95vnWgtYc9Mx+ctpVQ6WTNCHGUxYl0
sj+spj4WyTwf7IIRUuIPlaubly1hoabZNFvxmshFKD7mOhR1uEFPkxk/8UUMMsfv
wdh9sRu+JBMrBBF28OSwEyh7g332GJYEbhzsNUMDkxKDIc3oAdj4Y8b+Wxeh1PQt
6iLAubNZpaH14f4CGGL8LPBpumbivKvldStWBcJ8N9SiDyGSLzQgd7JEd3LORoRJ
glpJ5nd2ggY8iQyYPbvLWeeZjZnVdC8nN31KDIFwxCLkx+Nk/I8Oa8QN4Z9qGtyV
j5MuV8Z+c0TNDgemS9yrcHr8bYlFelk/GIAEfQQr7y4RR6phI52NTYLMvW68aK44
0Id1f2ccEY6P6rxxDjcZsqAoNcvHrvI0lezXVADissZWT7XfZdNA/Eul+oQ7zDv1
sy2MdSauc2jtIB/Sjs9tfo2/riXUL+HrTFQVwG/3aabfICLR6q/wX1GSeFG5+B0L
RlcUVeBPlaQax+Tfg80O0pkoHl8482sPuUCBxStfl3fA3n95yM3xh/L5YEdx6Csm
tHeimnqXQ/d7iLY1KDmoVyHUfJASiOi6oNjjvG3aSiPIE7SzIKI0p5ZeWVU5CvbM
mLc7l0osZJRea8zLE01cMV6LVLG5kKvd1NIBBkFkYUOkSq1F5GPyg/xAoj5WNTGn
r6/okKh+EW8t84QoYA5oKXdookzf2yGZzwGwclm2tAzggQOGkbySWU932NSuPBKi
dcZHLrYZJI1SmsCLUbfaMroRJerW3ois78coVL9gISoEbpH5Dw8BJgAl/Ughtc5S
MMyGNZ0ckofxKG7/dt5j5XF5Y7LOp/ueVdyjvol6dT93F3/W4QIKls8i2mzLn1ez
X+bkZZsZjsdRVxdC/TMteT1cHPtaiqGSl8Sis/7uTihHL+2+bDE/aairxHuBL7ZE
kjlJYCe7NcU1Zk4o0sMLN0SsITxY6uNYyIkBrVbfM9Y1qTZfkHtXeIyXwIlq+KyE
evnVu8o9w3pSAmYHcJJEVPB+7azsBzLzobFbr4yrmx/gbl15h1rn7zsbqAhlzYq1
8eM7701SIstH8y3rlmVZYB+7O+XU7wZec0H/BYX+0UlAxZr1MRQKqRCYj1bIP8YB
8FcI0gP1ibk/Nq3+qbKplSLTH+ZAJP0Jf7ukBiCf8tmTEzSY9cyOFmroQAGKo5lX
C2OYDeF8ubo0ziYzZU62wYJ9nfSESUGDBMPtJMxjRghkV31eOCxKiwq5P575DRDq
CCeEV6UouHKvUhjJPN/gDzQsizzJAnRWwdChUNlL8I4+K0qQcXlC95AT97NyW0rU
blX89ZV3x2g6QftrnTdLiKchZO6Ijyq7cWrR1oXNDkYGEPZ1jQdsJvEp8SdHtPUh
vF1ECEM1ctZKo90YcjYICzA8pk6rZXVqH9/V104i+8weyT3KdBAQ4vHGmniv5q7o
9yTn0qjInHh0oQw9LH0AVFKr8P79nr1bZseHutrV5ScHlPwhCyREJr2BoAwQqSc0
wmkxAAXsgsLLssddi6eJqtJucQfjbvM70FOpdoVD7Pf2/lnc53PEvLY32QGXvZsb
aL/EWzL+hZZsSRCEyG0FE/MgR7yVH/2FSEn5H4BzNnvU3745StIOQRIlZKkIaG93
WYZDniUPkebU9t/jEONEqYoiYhPnygduIgPXPfBvTXEyw9wfLqJCmvTirzYFUr7o
dfp2zE2qh+N34/nvXwoyl9KA3SIcMV6P/s7AGJcnBvC+w36UxqojWoId6b7DN6FI
VnGA5xRmGrQqRDc+0rv7wGJoSV/B0KIRac3H14qEL8mNbtAQwDBQiLgQ9oQIDDyE
TsK18yl/enfItra3v4oBlDJXm/XUeQH/lLNt/CXHUCt0AkoFZfdPJWyl8jb+Se+g
FQYLu4yQivZoJFZJHsbFSEVQNHgpEsyF4Wq5ot9r6YcRjj/+8PjOGD3PzdsgipBB
sLwJ4fsXJhw3swImRGdLpKKCB/y7NqY6DoknOCuHMiafs8qy6kdbEtJh0LCRhhyy
dBTjjOIWnRyZrqXibHsP7jAmm9TCxB1wHgwiwGn+4uIqPAyNKS2pXK+rrpVXLU67
J8jPW+FbcA4ucqBKaDa7gUKywOoir1zVMpFR24Qw9Ios7j4aNkBYqJYtC6cId85r
IYoGH6m+FIcvYfd+Mkrl84exe/VBa8HH2qNjMV9UbZ7XmZLj9IUco9J+AASzwiNS
8oL7XIy1c9q5hwON+0GBQ3+9BratiFgVxDS5x56u1yBRT96UiIvanC28v1HJFfOs
iZMPc6f/qRLjxoCbP7K+yIlKBsmZv43pe6ffB/rvaD/GYgEAelc86uXjFbr5MoL4
euK/OjE0kwri7zf45SSMNQPK9tlkXHQAws3nH1UBsdZ6ZP8AppRqGY7VKw6KErFj
XKqnrO5d1iVScaoZFMKh9KlZ/n73xeHc9oCMf8MLNVm0HyVKP9gO5CE35+451w8x
S0vXubIijnEw7WqEZx2m4sqFFhG9IqmjEnCLGIBpHXZWsSmfoQDamSx1ETK+dcrX
w9YVKC3BcOJ+oK0vWHFSDla1cv3jAQLyKrY0PKbdpoaDAzNpt4Z1VFl42wK0oqce
xg1mDQIi6WifR4813YtAbOsv8AOGxUrRLovcgwW+NjVgu2TKCf6psCWxnCZUjeOz
dp63EHvxFyySqO7m3jkWe2BeMXo3GMz1+xXcJA4CpnGtOWfb1jORG9SEiReP6EF9
QP2mGb+80o0YBuNWEMFJ45j13G0XwdY9ahlGf0MvwzLrW7uDLk/Ql+Z8elS5WeD7
ag46otm3YC/T8sQN4Xo5t3/gYm5TM5ikFuUkDxVJjsGF0yOWYydXw1Xo1WA3pjJ7
8Kx1zPkN2zCWKPip/4usHmMBYPcBUDakl42jKW+alCG9mRG9raNle2iEMDkb/OEV
7hdMP4Z9SsA9+4LfKoI92D811+pjBLqZg3weHUbb3QdGtYLIZzkgjkLukrut/FTB
jM5iclPxW2rMTDukL333kbqOGk2N44P4AFR0U5QboLtBqHr/x++8UDj/DAcnZ6wf
zTt9QFTB8UihTXx9Ys8wwMWLrFERab2AGuueznQOXqGTlBUFfoPBYCLJIEdNM+Yi
432irP/nIrnsev83doA3VRy8yAvlA+SSVM0gXZOa0FaY24cAzHFxrZGPjid1mR2g
XSktB4vUqmH8xAcsR3t0Tqy3L143dWZWuU6R1J1lGqI29gB5sep4nMaEdVFK3SbQ
G2VnyMmzo7UcBpwHwWSzoaCuFnylJcPS196J86W97ihT10krGIzEkKVCL6Ifqz5q
4oATrzmnbeTsWjpKI354YHYrzPh8AKCk2lJNrwXip0Yee2ACrOXRWXMrvJMjXsAu
9aloq/niq4Ka1fDv1W3Q6AcTFBHPSPJUEnPz9tpX1y/Kz1uHDl71zTnVei0XoA/v
7nn8J7Lof1GM0s8Ki1aBt3Jm6FcqhARks2CVY2J/10lirx7Mm0+V86B6wspQWUfA
d9zeWmgrEgkFwmTV5shc79DAMDl1iMtToWdN6IUJa/BLUNgYXmOkfUxsWUyPItN2
v6OL6x0M/yBOAtjqhIbLdiTVI7xTRktPqNt2niSiQMl6eSZHRSH9PcyESzqMGNKQ
ziq6O1OxhNcgVNdSHHgX//y2McOrpLW3ceVyiItLUPLoSmuAQxKSMmWsjC96OzzV
hEeGKRS6wiVni7llOs/iUKh93Gw91Q5YAfuD73ylm6g1Tr6y1JNZl0qETi/O/PhK
CGzt9fWaGtYtmpIuv50ehUPzX+K4M7WHCG0RROdI6frK3pwf/Egc+iUnkWQFwMNC
57J32qePUsdY5KleS5jm4WzpAMGbTMAJrIXWjb90DsN5Yk9fI435uAhGPTydHDmB
FjSBJguup2Gqqy1fzuGodIiE/VXc0BUdoPlNS6AYMXFtrixpa9KE9dA6MkHVqNDI
+p5k5j5PvbkkltSkIKPZWgCOjrml6n4MG8mw7oUyzxUSuZ6NRmWyrFPe2fkMRMMy
clQN7GHWOtS/sx5oeEtpKzsAIsBewyQzWoWyCXLW0eqvo57lpctJ3+xgTZ0OucF5
RJcFy5hXHQHEy4erLAZaSveFxNkGfX+wQWUXu8myS4gZZhA+9WyvEqOxJTsDOUQA
t1+Yl8fQs37FgZhwbBYVR1rn7RBG31E2FtGHyRth+EaDbnAL7uR22fhoa7rFKRpC
Sgm/ZvwvnQCPPgr5VTRE3sJNUrWUGAtriSBCKOXhiA1oAAm/E/s3+r2y6+ROihF8
uevTKSb1Pqv/GYjZcs+DhUaFNvpeES60pQ452cQToeYCt0n3Vz54ynyhRrqc1mb0
BX8w464ZstOqpPB5zoZ5iDnI37O2aAfkftbY9hlsMeSin5QCKqEl1DPh7za/FLp/
gRaPJLogd6UrpLjqZPUl3Qk3ke/qU0ql8JF8asHyJFuZzQInWUWYp27MNFTORns0
c/zrSt+9sO3fBatCYab4KNAHmqw8uvHtpuvYw3ox0n/r6Q/PVyVFKoOLYUgflJSJ
MOy5+6NoPO4qwcfHgQKX/k5HczV5xwJ5blTa3y2Xt7u9alh0om0nsMaonSbLc8PG
WSoiBHjMkmkNQytnME7pOetBc0Uoe6ldVc3NGn1tl4+r/a7OTS07PEHO9krmL8FL
QY+0qWchTtEhk5KnYvD3h73f8xKboXChBxWpx/HdWcfhyUpq98pvXfA1MPVUCtpo
T5fFD6zrXYJ8b0CCxG1hSU0jHBsgcSDlAz/MGhYaCRAQHCSP5EuETeUPm91OfgWg
RoEH7C67jLnS3z2Ob+VvzQKx1Fp74rK/3TOtX32SezzrtIJwu91mI4aBiyh5cRKT
9H8RpnuyK7kygPrIk/chYkNSzY67UHE9v31Twbqnpz2OUk1s9Ehbk31EV7aawoLr
hgym7NNcDNND2MsFK5NnrN+Jy+7OjfMQW8Jsf28E+1KGEnnu4A7M1MVZcxjc4NDB
Do4sFwxvdMwDQq2G9aw0nzkS8wV2m6xmgzHJlhUY5gkYDIfv8Zwf/X9vCaejYawf
iM+oIJyfSt/sBNocyi93jVYwT2Mr/90qLlPadlWdwqIzWNeU0rdwqPfnvexNril1
99zYWaFL92HCaPFfugAXZq6/vda7sKlYi3JjuaypLtH4MJJWhjLf3BEgbUolAghn
4yLDFQelF9K7npmwSPK1nvgoVFQbiAqpwBtNYmxSDp9Se/T2eLueZ+TZB6c+05wR
V+7Tl1e6shoJ9BLIjGLJ3FZUyHhiIwQwGhCGQtcNIMsQAKnu8iRJ7LIacUDLNZ91
H33XRX1QPDniAAFnLS6L+5V5uczm/EYDYYGHwGs/3DH9tbBjgtrhTfOWspBeKkZB
PvvmFB+GYV3iIeAHaFLyGV7+ea/2UGOywqrDk9gWjkeG4TEmjNEmWYXhFZwTW/Lu
VfSc3Mf1THOKzeRY5WkKHA+hVeGeUvCpG86x435zuaypeGTbimzjLJycV17yHlKl
6mDLK1R+I8IxSg0c6i4pz6EoN4cHI8zQ5Aa1hBKbPfOYM+EyfjxdTkvl6GNXLdvg
YGHYQGC4ws1cO9h6a4Xvt9vf3LWkxh0zo932deRy3PsK+dX0urSx4NMGxaG51mQJ
RQZGuWnX79tUnVj8+RaBNDCH6lMQhdKXlG+HUk5DuCbE/mcCpWxYxNKxnzuwEu9Z
1qpFshPR2Ma3xaNQnl3SajxsCJN6IaLYdRua0BozSrwQOdBpM1jKmukInTwWzHj+
1JoJ57hHSBOo81aKZqe0rDEasf2djiJZTr/MDs2j9gKQiQNtIZMqDcXEXUmV/thA
85Ye+0OLmiLLxfzIxJKZy9/3M5daIfwlrXuOTsHqLOYvHGGFJ/OF+teTLckSBnCI
FjfeaAkZ19oDBOdLc1y4sL4El7m8Kn7Us5PbKbyspTcJYVPXTe1k7LZcrDoXy1cV
rLbil6TlT9qNcUPjAmg8MC8gcEGu7clIEGJxIto8NQ5Lns5VCJIPdkMdn4ejBPWu
jVm1NSSYAhGRCRIItLIUGr8OgwSWargvdFND36Ve8YeA3UiLZlIrG13iXbfdJiFi
t7xvGVUz+94vSQw6qzo7WvSttoUdXb2OfXuF/PpYYJSO4l1o0KTn8tGUJsnW9xqa
BctGYDernyuSwnwaxFpmXR0euiwfHyxhPbXFavYTDrxKUchHFC62Rwh+FgAn3SZZ
0l02zErnIArP+e6OQ4XRry8C5+0H6v5RgU5jnUtpEBPUAXgfiEBdZAxAa3L09Aas
v5Ago0LeP05NEt0oBDTih58CYP6WnRFoeuYr6OPUggD5V4DhYuxxBkfrodYZkyK1
QFSJnQn8ONZAPt60z+iA3O/qIiMbSsy8tmXIJyHdOwCAmfy912v0kR35z8UBRTro
YVIGdfVE9bmgtYNz/mb4MaeZ3dC3SpRtgX2L0d/iv+KqBLJllrHg1wFY1qQXX8fT
4HP/iOIWKklAETxt/lB/gAE7abXfl0tMqBS5K/55xeA4jvMn98cl8784IHL0r0mU
AkxkfvM7q/4MXiJ7fZ+3CsDMuaUeEtbgQVbA/5bbReIdjXTOhTj4v0BG018qHOoI
HKfD9PluCzLOhMQ58XBGexZ/LlJ1pQWrQqIRfpGVp6VYl6QcytJlzh4CzUQeZpkI
QJkrP2w51lGKnJhrjF1epfVdKouvoUx+A1TvgNiQPRBdP+FeLecSeRs1oY/56YgB
jMCdc3qwTdSmT108aXnzrDbWpcVr4CW+wKDRvprKy0rEAjPeWK6L8lx451UjA6iN
ksjvgo5qu4WHfURaCQmVqY7AVyzQ4Q/6WaRWfCSV5WLbgIGbyAljDzGcciHDNXtg
5N6qRU5sK89Hvx5w8ihKGk3WxAeKYUQJbUkcbN+X0x2xrHeffCmDio87YV6gkmmq
GQ7L7fnbNBYrAvJr9B2DO1nzxFGc+CRDC3kA5nV/GPmVzzEIWH2zEjp5xo2nH/AV
k4igRvXYpZaK51rhiQG+EIFqcpgCVoPZz4bf+mKhz6FphMPvBMe2Six8Z6WR0c5O
o9F9vCCQajjkN8Npp3mI1DacChr6UWAwysoWLMrvZ37GpPwrtrZB4GHxtmy/+yy/
JAfVYLmgfYtCXBYC5/juxFbiv6chft/pA7b/Lg7rGCdGuF7/RsGwHXzKwUk50fzJ
mevIkB5MGAYP/KhN68C6Gd7BOqXzF9TMillj/xSBU5exDeZ0WOZqOEyeP/sjGgAg
p4fv4rH1vvzQpATvlPgD0JP4zUU+7PDhlQWURvjs8ry3ir0N8vaIRGyk36D2LxZD
eQ2vrZahmGgysszyUqfl1hy0cQC1WIHwCS11T7JK+9geWW0zWGJeuxbao0nKTq4Z
deyDstFsiB9KXEoRpB97yK/noT9Yzjsp5fnO2SY7LTwJnnWV/zgiDFnuFdIiwd+c
uDYjpoyyG8whOE3tBlzEz5R1YJL6xCffENHQcR+VfRDM/ruPpLMOumb1Fj/FI6Ci
37GIrnzqlIHsiyHeL4SQk/FgXfJ6MHX9sVtK/hPNpbAi8IWiEWAQIkKa/yOywoEv
I3qUrsbLWL2H17IX5n2PoOoARd3IbTH7hGsjUzWpnSt6QCKrjxBHIctyQ2P1iGLc
CO4GkVEMFVLQXtnhxGGOHgkA9KmnUasSivGLKMdbbQyJWe6M0Kt2rIHatzX+t2uS
U2HQ1gmsG6foBVJgO2O4LWzWSj8snWVaWOCS2YshchkhWjs1eS/W1WDLA9/NHYLi
SG9/P5XglW6wIB5izzxjWkss3ooC3GRqneuGItdMlwMbai+gJxQ9PA/Cy1wOcp0A
gLG2Y+K/myogI5YYSiNqQ1x3TWL6sbzg/nbeMgevVXu4KJrx16AcKb5kWy5zaLxu
KN+l2WG8R6rk39epGkqfhE6OJ0Oyf8v0SxyAu/Dp0sXuaVe+dLWH4toWvpMsNuI5
LmFwpWrA9bTdB7Nqa3NiR7zHzPJUPmlqTHAADIhH9XBJpjJtJblujuHWuwJdjE+l
ZmTQVD7OflgwUPSV0h2eY72w5GuZoAb9HF4g87SgIyAGsUHuecQ/CMWZYxwfd8SW
plZPu7BafgiXuUr+uAKctKDaSnc6WlsdDMhOWC2A7MTuttPWt8Uq2Cp3vzGMSSyF
dNHSR16coupkA9RRNzx208v5dj/6S30JOOHiPXYtwqD//mKET3LWB52brBvgLE3U
BOleJ5s/U2cuHahEv+0LjZzEzkyuOfsNKF4lSVclYExsu/16wiFZMzwUA/ipZ2AP
Dqs8lkVPtFKOYMDLf35Qmn4MI5wRGh8FJuujAyoTQzsVd72KmDp19AqtUFH8Sa3e
Ie5DD9NwdRuCtfM/SWkhnd382e0QC2CwteVv+s9bU5Y+O1XzmrhNNwgWUX2jMEk2
sBoNEvgz7mkyC7QIYSbas8iJYHdulAz9HUQKdElGDBoS1qgKv1TyCU/XQlpRjjdB
GJMt8VsrmVu1TSOZVZvdxR+Kdgqk8m7oJx4+czNB5JGDgHBnVAtYBYlNG8gJ1uf2
fouO7iLIkiFGM7wnD6PTeYJC2PD0zSeU0bG+GYVfcgHsbTK23MrIt+ESuxZwHjO+
Pp+odlrH+fWsKYD+vfSjwkfTHdl1Vzpv3siVMch//2b6iXhrUFKHgWNiTTeIxsoX
X0STtd/XC3eSn2mT0iSw6RH6dZ1XOcFyy3Yrn5IRkQtOyIikLUFnCMPxUQzRX6Yz
XGqRMQyxfzLuE3nN3fv+QRmgCdBMh7Q73MDsNsSZFx8dhoGCnSoKAiVw4/HwZFQp
p6P8SoyPHuPg+n2uzo2qu2g2ZNj1NnBse8p0NMk3Fvhe2QRwfkD5bzx2NXsk1cvO
P/7rTJPBS41lPT48QEAcX/0taA7JIDS2cQAn91zFNjwI/sCrvr/bpxPGtN+tee2j
UtIEGFfBysmKyFhOw+l6gYG/1ER+Lzh5+uya87QURZfiiIA01V9uGz/8CyH1OVWQ
WPah6NJFbrDAzh5tp6F2b15l4N8p+yOs9pEwegx9k2ANwQQi5Li2+4iFYwsK6R/Q
tLzgwGNWggOWe8r82r3kZtb3bRw/Nlzu8sbCAwOTydvZNYEQuZc1bYW93YXLL9tU
/1IIXUhCccDPgcjRCEuQuK+UFxzBvQ6HhDTsWjZobtSvVon/dd1fOy+qXjXLUAs6
daLGxFPe7B2Hlr0tJAGRMHsEB3TisU0U4Q3m6XBQpJ41THtWtO1BM0oyGmo++bQP
H7LyrLuXckN4FSiCH2y2r7jul1sgLLiOpcHTb/leP7xm8PgCUYl4MgTno6cRwwYY
vij6fYXyj4vcTKSts3VGoYbsnrb6zIbWY957dDo27ilFjxvaG2QGvnMZ4syz6njc
LFx/XWgce+YJZzcQ7n6mUf5H24Vp0kz/LKc+803HciWAuLaqh3Ec+Bu6NBtE57Fn
355xabK5EZYWKXDPXW8cJk+egCk1qQknBh4/Qo5z0VzTpLi0tlmWSJJmrPTCYnba
/Dbx7scLeOCfM6LGU+gI7y3PsTfGoAF5IjHgbbTk6LYJ9MzPcoy7ih4znHlfzhYP
v00qu0nXy43OflETOV7TkdH2zL0Y7e6RGwX0g8msA4S/RzWM6MMiXYfjgOrsllvI
Y7dMx1KeFZsJRThNadMEmrHZeJKS3KLMJVw2vOcEObMBOGcmrqS3uW3HkBdQB60F
jyFWqYgJU8yqenKeEIdROqZ/MRRHShe6eewUrLpUfvn6MAaHrAz5VXD2UFT9YrMg
0/wIMJsudRkITIEMtnpxn4D6lDtCWbCdqCZwYAofFxwI9xn9raaiJVTss/NRuRvG
ja2O2DQXIEU5klziVQWiXGDXT9GfGxXqUuojt9Fa6fwCkkhjHR3iv8fB25pv5PyC
O9lslmVcSm3PANbdnAuWBLE8EFLdORCuuVYOpjnN8Ywems4iXZeQ0R1nbk0PMIxp
jm9QOyTOfvoLtnLbMqWpOkYa6hTfxCEWgZ6ST43i3PrVEjwEcMXOp4gAvLSlOhVI
wEEBv6bgVurKiv6ONFZybd2UamEJR1YBJYs/tP7HlWbaF1lqxtO+wtgje/I9RPMj
6jPw2bdd5XPMWK9/iR4umUDqmUPqC1Ei2m9gO44GenBk+0PDq+qs8QbGXRPaQG4E
8kGIBZRICpwLo4huWl14C8uAXdtTxgcDHYyUA6urFGWvW19EhPMARggaiktU9pW3
2UjYk31EHUb2c7I0iW5EugTwvfk77trGpEfTZcCfd5lozsTDAwSCRCGHwHvR+ETu
VqxEqwrmn6iTok0HQxWirCmeBjQhk47zX6DYKTv+LU2Jn1ARxraMHMLXNqxbDCu9
aEsdda/8wWnga4ehDloDX8vQpNNWTbKfuSaqg8J+FJ91RTvx1qaUMlY3HhH011nR
y5VSkOVdweNuroEPElHnf9VOPR4jDEcbwlezXWoI6frdI0/5+tF1D/tjddqmSvwJ
YMWn4CGwEy9zJjekiuQ6QMQXcoaNHNDfyfGwmh4HebA8b6Yzn4vt86VD2xo15PAk
1F4OXDz3SaSlL8NAIcvRHYOlVnjvI93ebGjX5YlEqQc4FRff3URW1kuq1FDLb7s9
TMABcFIyHHMhu7o4cVF6EsQ4TKMiihif+vfF1qJdFikQSkvrqUmHNani88WCkXIB
WHdzJ2+IhtP7/qCLl13LgFlCe7qJ4PGycNhPY9k+i0s5ZA6xOHXPeVGdw1T5QN6v
lTABh4SE32IF+UCcHMoI/tIIYau2BFRt6TfOkh9gU3M4BN4S6rZcpNaeCqtYwlrB
Rupvk3qqYAGDTL8yQOBePn4RJMJEV0cwS96AAnpbmWDlgLJWHU6tfiT23wmI10mQ
8fWCwGzrQB8Xk8hBn2McWnt28wChlk4RdKLpN2cMgvf9gh/S3pNGVXv1S220HdK3
VGKPQWQHmr6Grk0UU4R7a1Lmn47t5PwQnCI7XmaxD2Y+Nwp4c8MMio/M5TKS6YWe
Gnvmb1tejjp2uDRLkz+9tJHJmUGG0KUSla1YIKofN49I7EznaeS7QBgymzdCdtLx
AWmCiDlNkZw+1ZHPlUvfTWIeiU45ZiXbovPkoU/UCfQ2nvrD+e8ZM4/y6R56qjM0
JMaVkT2NpXoVGPC5wN7xirbTECuILBsTKBvgiNk/wlWe66RmqgcHXIRBrlRJR423
DQSzotI9dbUGckOWB7p2kiFm4stHSzW875qSMwg0A2UIXb9THaOv+Owfb8zobp5N
xazZPkmnRG16/Dxyoab8TMwkGyyeycCC2AdZoWTBg+AJkZcHBR7t0C6+n5t3QlVG
y+Qi2GYEdr7AmBL+L/5tiTdQQ6Y+ePd8kwzq5KCuNAi+HRXO/s1UWVLyNQkSksBs
jW8jIZKMlAkJaQp4f/wRn56y0y2BrpS5QmJmQyLOYZ/tpRzrs3rJuJUFg4ZAoU3F
LLpU0e8V68+Ay1r3oPvSLtBy3lkYnC7ZlWav0hVRldJDPs8HNdcAh3jHx/0+i0TC
hlQ488XwII3wGuYmuzs1xkhxFobfzptNcOncJEIyNrhFN72d666mKYrPW3gIlbsL
winC5V8LdFVWs42Jr6jE/DE9E6FgVYLQQ91KVPFu+ypPkzyR3kruHXmKDNhdrftY
KSMWoj5UW1rhQfOnnEyAOAcYL3h8VbMzghSmZAJ891xYC09Jnw2bEBMV5ZMME3nM
6SXrGiDSyOy+rWGX3zZNCMXmposhIaH3NQ6XTCaWUNqH/nvQF22hTIcBhZCdij6g
021RIhZqqAcOXEv7D1T9//J1VAw9vEGG8wUro9cjYKq6vdiO/q3TybWXXR+NJvRZ
CYSo6ThJuOOc1xdZuAgQxsEOGZaaVQhAVNeEJZIVcqY5jCaZwYszkTApq/lHK3Jg
/3np4Cc5K9VOgSda02AokHVCSSaLlyRRprlvKOps6i8jpRW0eHKgKPtzEiPBP0Ah
ojLRfwbf6sn/JoUGfJTq848PFlLR6pi/R/q10Ch4Y3CqCNkRK8EjZAPJv9x6AvKK
K8excq/hlF3BcJhB0Vd0Wn7miQWthBjfIhXfNVh4yEqToWuIa4ZQSvAy+u0dRt//
4oZb0ugFugYLaLyQg3UZhjkXpz1t0Jmk/pDU7h4GkQNtsnJ9th8utC71TE6FGrFG
2ODaLW1lZbErk4BNuQYl7jCOysXtACe1JWeVpAGVWbSGU0y1rIIesO1QQ+uIkqcE
ugGDfhfR8Tih3731jDEzwfIfzii//le91MGk+wU5eRSbCnev4WxQKML0ZoDsNYKp
8uYx1q2uPI5tYoQfqTCIa7mBy3FqqZUqD4EM+F+ES8jykBs2ToHJN59N/yx0Zeo6
aWztfOEZTZiHtLu77t7GQ1cbTYvBiYlkt7N1Nubjhot7PJKmGxdvBL8f/mi+qNZK
A6rOonVV0MBek5XP+1nZfW1KvyEic5EjEhzSgE6XZOlOqGMeh/9mefE/rO/jx1x6
EuxTacbWLxLyHsMIRkQ0DGpeoQiNqsCakg9Zj80nG/z2iHjVc4hrqVUE28t9xK5A
SxHHQafS/KNUzHjaUMcAFdGTwgAf3Yfgelkj89ShV2bJAnLPRh3LFDVHPHs4qz7k
7GFQvKX40urAKtysoUkWd2s4sXYTP7/L0PjNgGuUZvAt4URf2uPMUADU5q9JEUPQ
JMC8kgSIoMbS4n3tmKg3/HRTJZBN0LMgOcdtRhHgp87tJBB9RewghxUXBt5RnTF8
Stnf3zHno6EbmtmV6uE0c5EprwEicbvuDLfIcAZXF1iqL+4IRX6tPruRhLLg8dx5
p1d7O7jXOOu6kSWR3D/MUNwmExys1bmBuDcaE+vFauOMRa3iG4Fuiuh/GKkl/FP9
s0lkktQLEF0w6F8eyFMIVMlFwYIbruMO/gqG4HEWN2GJyeIkxzVG7Q3vjCuzysId
c6lxdKQsbesRzNhM7jSWtqorLZnDO4PQBxfo6dq0xkX5vkd4My4eZXigfCGtuHKK
DuVi946/ke5lfDBSLRy6x6JxN1fMOFLh+0xhzpAUtRm2XdIeSNjhZva3KZSdqwZG
NEiXVVs5fgsX/NCPcWgZELuXnhp+MgEVJAbVTmb4nNMb0vEICHXen8V98S1ycw+Q
W1OYbXfeTKk5X21gLqDD9rkx9xpwxfclqh10nqavWFCIUDM5G64IxyeKhVeB/A+A
DrGWcfN0lpCqizTnrrvB5vkYjE6UNqirKibKKtDcRZD1tOSYVfrnhy/y2pKQzG9S
jQsCIB6s3GzL1OJYOPGKRtJiMwah/nIjksFfOM7Go6y9J1JsM0176NFG4yF17eFM
sJ1U3ikfkluu9CyGyYaKMsT+Ti/YaJP0nlyClMc6mE5yp+48BTSLtzVrr3HXnxqL
yTyB2+rajSAGfSWGkrOQ/FUrowDyUrGsPyIDnm5GFY5jjfOxDIUWNVDE4YEmS8l1
5Pb4s8jgqJia7LKI28dG2XkQI0TJwqm1oq0RuARw9cx4sOaMYZ9gxL2P5U5CSrks
kPSf4vgBn5OSdlFm1CtCM2Tg6czP1jmUY90q9ZJjbiC8a/1nCKx3K6RfTaBeZ/Io
iTGHOdpZ8hUxEs0k5hCEmz0NApZCL3rDCHi12y5psy7jX0+diud92KGFYdUthyxL
+0vhqycHqMctgG1swEtL5xsf8skAA2rsNezJx9uEaFCkJqJxiCH+otDJS4jZyd/z
TlSgbKLa4sk7HScjSf1ndl7K1chbeOX4ikNko9xNlDm8ftCBHF/074vBYqsuBTQL
ciLDTi9j26HBO9RJpfP2S8ZJxdpW3lyO53sG1G17GJXb28+y8+9PVxCMtfv7tF5Z
6WJl1lT9II+V9emsfxWplWBsXA8PKs1XzmMmVha5fq8S1H5YOdmd0jEi+JoRRE22
iWbjVjfnR2YL7fwaPMF1H0bZmpP+wOVsUNPoz0A5DvkZkbF1sVT/AetG8yqXw+q/
OB2OoPAsafGg69Sb3PHfldqzgW6A5rKkDPvgKhF17+klCNV23NOquqDNp4fi30/t
aXvmoTExr8QQptuhfPDVZQsIdbkQ0KOqGlyBo9jXx/92N9ybvDh07lwd15p5ffPL
UXRTeersw9wUMm0+jQXI9K0w7CJvvetr8J23xLWfNWEAggphMyfcuLihhQJPkuy5
7nfcNNRch5y5G+cWTVqzasz5iboeb+FpIECiZi0PszgC8R+sG9n5Sv7ytRj5mx8v
kyxdsRTsSmEB61L3U6wGf3bDnzotOyc5ycs3P9AgPHTiIR75vuazVFncxDgzK0tA
HQHjBTRkZOAHAtZbQGJg23oqYdOLn1ohoRD/hKMVOI1/spS9/URHp3syDiVUdzJm
2gZ6WTph5P7lijKaLIeR8n1bFgkmsDX9XbVCQIvXMRP0S5sP15wdzVn5mKDIgZoM
KHBR0Mtl+AQYmQw/3norfcvWJwjcPNCGlAbAZ5qMRWfANDdrO+gtYAabSrGgZ32a
kKrJDgBK/dtfwXhKrdTUCfgbSWnu9F4p9MEdklfeIZVPotZ8IriyxcHjh/6qi2rI
tke/6WDok7lg0Y3axXGz0wt2PpIxdbV5hRu33KS67kbQ8I74Ze6ERSTA8IIJVKBf
03pa2dBWgXVW28MSz6VsPKnOhmUhNVepfkaU3fSzEkphOclZiXyuOB5Nl3DXrRUc
lspQRn+6AOtJ1+aX8UYBQyHaMsJHoJv5bOA560ZFQWH+HxIu7XhoFR7EbRgJBhdM
Qg2moQbmIKiyONt2Dd53p0Qabx+59bgGKboDQcKadQMvpLm9pNl9ua7Pelo6ljPn
rzw7AWp8DmoOHXd9Ahy0qgyx0tvcvxCRBNUIZHq8Ow1Bv8GiFPr3k6UYBQeCZtly
fXcQVEFpG9h7CvP4pliSugzyRcu/ed4oZA8mLzFn0pyxkQwCX07jK/KFn9tVqHjY
ZRGXS19NKvBHU2aeBzFOzYpEtcq7g4BLqgVlALMSzmz+jfmxODu3l/dm4GWIVxyl
H3Z3qR7kOgwSCNi4UOeRCJPBcXQBfI5aGB9KvfA0JtHJDmVzm3IVPG16uuEeOpgg
gWUVGp1oszQBklg30SIopAsUa3+TBe1QqEJe5tRYn3CgCxse3FR+ZS3KB1n0aTnK
synLyaxeJCxv1liWIIYik/k0tnRFWxN1+T2VtHDi7EWz0Pp6ed4naOj1gSJqIlzN
oxkm4G4LyuC5jQtpgZsdZTGitgvhqGf0Pd0Zn8Hi+AsSuuVveiP0dz6rusBwo0n9
9rTL0SFv6vlUllSOvM/mJa60pEzp3BhvwbPXnpf0E5PEHn/AiE7njfJlfXMWA20d
CmVvnVeuWnep+t3wGuGKfXioAPvM5i5Nq2MVFq0T6x8UbqPMTZJz3tHeU/i596Bh
7uvDwnR/7DgXdIV+m3tGnx5YBx+sJLwxIxR6ezwf2QeIT1oekCXyPhSdA90MmZjl
AW7i49eJc3sZRaYYVo0jpKBYmziUPEbf0Dmat/QtrFO5fAmZQELu2lJEuFAo4wSI
xhPtK95DVSlABCcpodlpBCLrsXzgtE29AF3n7453MAHYfNpT2m1aXeoufwhShccX
ZHXJnlBnAz8MjAYCfvG6sHa+YGqEuoqQVaSYU5mVppYrK/K/f6vVmCqJs9YscF5G
lU3kmlhy4kYK8qmT4bm3Mb2YCIjB7Ps3tOKWNZEiThVoNjNyXmCJ6vTrmB+6N+O/
PdZ7cU3W/+89d1XPXaef+xdu+l/pt6UdniF8rKyG3mgCYu60VItYKwhqugwW/L99
TgnKcw/gV4dHlT97PhpWeM/YGfdCqvNuyHnY7mDnH/nPtqjgSapBp54EXHeXpLyF
eQ9cM6aOWgqecsde55HBZ+qNxHERXKEjnQztCFn8IMKXyR7TN0z5kqLxMqx89eON
RwH2dBLNhe5Nw95HQ5Djbrrg63sDIDotK6x9HFUDLdoBQXA4Vb9yNHvvMgtatJWp
h98BRRpXWPBQ7UyiQWxLFFLLQJ6CUr7/SEyU+U/xx0ZD6xIrMqVO07SUFhg2JSzC
yvzqRo9UBUVQn7FN2ovsFX2VhM1NNXTGdUiTIfy5NDhsUp11Co/BPrSvdTY1tVFV
y8frXk/QPTY3bPvRtfYX3HHDWdVcUVm55NhqgvM9Q19ojmOybfLL7vysLSHnfc/k
lEmp3tP5KgBC+WRcUSI5scacgQzmgTn2XxKgOk2VlwcNpeWtwpkArAtl2c6BSvL/
WOuJswIWAPLFDe6EM9FaSWSb39sx6pl444ZIwAEDoZw7umVWzZ8/R0t72nc+ehlC
IRRHGDDnviM9iXUEaTfoWjdsvilcAtYg5wunrVQZgLglryWYguyUiOy83So+JDB1
xL0ZeZ17Twn1zps5KmC/25HkKF25ZhaT9xC3Z9a+SUtDtNBnOy2Bqaf8juWZd1op
U8bNEi/OstVwZ5+zISLpGcSACc8OqsVFG3skyRV52WXuTfwTcRY68O7HKdz0zJAP
b1Ja9QT611qLUmf/gfXYQQLaqlYZ+OBt0ZeXfKu9TCAG2pUsWejtx6boFoq/Ib2l
mWIXPC52Re1QDQp6s1BBg4HbGa/xwi5fhk8qKpVfLmKQaLJqLFnnAOJXWQ7MfGJa
cSMSngZVFiqNBTNzuV+rnU05xzSw099o6jwjQoOT+mnmn4qYLoZhYCv7XbohKGMV
eYwFulxNF6OujKpIB7Z2qcO/A2b7xVcdXynzj2pqDGSJCdcaZ0TOrsOJnI9p0Aak
hOfO+/1nKnST47/a+Tv7wV0md/nMun10sllZ7KnUmm7b4V/7q3PVu/K3p87siTwu
agvjzc9HyTwdBLOu9EBaXAtuVjxHsQ9v3mBSXrKFuLcnJ1Vh/HJOcFPHn3YqVLTb
mEQIQLPLQnipY8tCllKzZKtGqzqC56OA1N+ucF7S8ZSnxu/Cua9gGJlgaU0SYbTO
QlgjaJzJtZPgJiLYWWhhEkA/jMEMMWNE2/K8/dIG/1hn7Mg8bEaYjhkd5rVXZupE
3+96vpqSsd6cw6TXXmlxqvf7Hqvcd13peXYJ5cGEKBH/NmujNgkyk8Tt1jNd5pml
U4dY7WwG1kbYnbgvcRyZPW8JKGZgKcwjd0uguQCKJt4ZsECsvyxz4pKmrYDrF2TC
3suSmVhEvBCmdYuv6QupN8/QbD9iBk0ShIgq3mS4jWAibCvTk6EHaEs6TGrPDagT
gaz/U6xqx1A5ta3R6i8QVQKfA/Gm93nLjHJUXcv95oheslpNkJ1yRFIVLIbGZfWL
YMnXPkDlX0iMjGx/jbTKgY9PjtvKTSg9aI1tsECCvub7gGVwzOzXpUuKEEtFvTdZ
mPLDWsBDLkM/8tDSW5f/eqdC6UbvbVX0BwZaMDGmCUiOKEyRyDuYH3In424QsHUj
7XWskeweHb8BY+xXpvJEeoBM5jw9gODhKZTgHVDxLJWzb9wHBA5CcNeF5hm6DOI/
LgZIpznM3EEIkreUojd6RDfeyfCJ/NYbGtW+obUz0VQvyeDEzRpDrYTbCIfFgyOs
mkkA0yNmVL7IlKNJ5OfAPi7BMB8bBgjIQm651Km8P5kpT6IZyVG6cU3nXg63S7mL
dO5Qd1D/RQIk94n2ZKB/LXaLSOKx8Dmkx8kmECnuvRKz6Z7O5kZtIHgmoi29GzUp
kpjuK38WEu+qxUEaMaaMmwfDw+2QlO/M/WF+gVnFWQeD53/OxluLqESY4ikyH43n
imK/pmhjxkfrNvICqC479tXxV12UPujR+a01ODwx1zRi4TIiBBaW3YHWz7CABnlD
RFuPhphS7WaBjP3yUpWZbRoAvTfQiRJNVonUHWlZgP5xMl+uRQ1PqDOLncwW0Fnd
dSmmFMaLsjPzCpNrf53ap2iS5jBQ0o8jZ3+YF5HOcNZmTHIB5Tx5COHlCe4KNTFe
adBSA1VUDXKj0/ZFaMNRoZvkxX0IkOqSmRxXaD6jwadBeuuzwvPlKQ5eyt9j1fWk
Dash+bpxj68AftIAQ8S3b1ImFp6s0Cic6qtbpIzX3OK4KPM8fGFCUUiSAOhyTbzM
SLzsyPd9l/Q5/qH3z1X/oO/Qz7XCIdnplYRPYJBAzIijEBLVw3JleJ9TBLHHQ0mX
1nT0a2DyT1iyaHL9A+wciS0I+tMwbaVAZWXzGgrCu7RRb1sNZI9B6xfe2q4pgK3g
RALrZQRkJ2gqgLAAh+kyUNVY0BrMLD92hgqmMm9zXaZhkl0MBM/3BwAJmu4p3S6l
Oct5lDSKjaZhRvkUJw2CDaOgqoIU87WBUAqnhIw7lOA64ZrJSeaGB9elAdwGTMAy
wekd5XIzRdKOH2TnJWQ/IbT4A5QVZflg9KTLTlx4RCEO0iaJuGKZ0vWBsGHOVqOc
mZPKsFatQEYLbYH//KdR5NAIx61MKL35f13FkkoiM0hvIEabv7nfoDkU+vcR2EZ3
+0BHPnv+o9fpx/l1WWDTcF4H2qFCfYCdIqYPM5rvuJNrk9ckaYl5ER6x+TaEVWg0
i0oNSMDrPEv3YZZorVA/MKJzyR9kzvHPI2/WAnRwzwg4iGlbWfpBQ442MRljYiX4
D+1vGMmZEimBiuL+GC1QS/P7dM9oseaaqQzci2iOM1I9vJhtYFkSHD2R0ikeZrmx
1dFy/haR5hxNMqkmgObSmxgzcS7w4lUWEhWWbS7+zttB4f9Gw648hK08tpJSrDUv
OBNexOAqJ/5brAJ6zet1RAXNG5XUaHWB3QDZH0qHSrO8/jPy8KFVSti6PCm8ARav
w+NSzMipx39ZI/AG1WSD1x+DcfzAaJUdBVHKIJYL2t0Quh9MEwzBVVQ1bajdRqZR
kljiJMIxYeB1C12JKgteyb7CINCsF84KNlY3Uthz9RL35PyYLzg5rpHtdqJypNKv
PDT2howV/9TSAeMM6RbJsamD1h3oky2ZzzoiW0Jjtoas5Flw+ovWtu0oLUl0aVCn
wsCUtEvsgEhnnEUKsmZrIrinHln/vUpocRfujhHzgi8FeJnOafR8INq9yp9lNBER
K8pmdoJz1p6JKr6qtasIm6KCin+AtCnHyb3QoqJmUiTRg3jGw1h56VL7O2Tkh/vm
F4qDKWtwol6MU29ejk8xMp7g6HUbowazWk3sRtyhj6mmLiUq+N1bC6YIKja9fhgT
6vph8ZrTGUaJQclNu9q7FhQgOpJ/KPiOvmAFbqStl9+yRRJCehBA7GzgaN0ImWV8
kRb3xKh9fYxl3mHpt1EVlWGXNyANhwJI9reBJ1ldutJRMZtYD6tNAI490H0AUXU2
YiT5wPlDo8U6w1Id9sSTvev3OrBjNiYbIrXMPDkSoOOqrUq3Ili4cHNUf7p0fLde
qs9Ix9Y9jVVtu2Vaq3w9DTRLG/d0f4SitdemOQX/9tKdQ7jl9fxgLXESCAVWv0o3
MpgQCq2kgsTasYmhkJEb5g2S9oGHMRMkvrIgoC0yRgwkvNVbulbsETqvl3dcF0Gj
c/JG5aa6nqiGJohrHaZofpOqcIk6w88QDYZwazJDZ/0ipXgMaM8cKcrMYslIaSZl
fHOyeMwYgiTW0PksgfwleSd1CLpNdLC+2vnxAUM7wleAwOdKIx+u3rZQaG/sz4dd
4Gkz2RFE2W3fqsgt3M4/7gtxlD/Z6FUOzmQh8ipomDBfWAj66TwAT/lin3KhuyAs
RpQbmWCP6tFVCQW4SOZQg1UUMjlkjq2mx3Y5F8Jv8aKNcHgXDKm5UAG373c6MdWK
SY6SXS8UieMZnK334Bq01rN1MsrugIMAYnnzn8ZXOjnSvTIURXeW0zPZDoTi0ePL
hc2yIHFgaoNmuWnogNdGpO4bAQXSPVnrppKNw+HuqGpa7OLKZRUaXeBs1nAjXbTu
o1kvFFWP3YlneK/4xwfix759nxxZjeNVJm1XmEOpQvcblZ9xqrrLIhqlWIdHpk/R
WKOll4l/xZYeV78+iHb9chVs5I/5AqZYmlocjPK2lBgyihg9OIfcs4Sjki/zVP5j
j08LR9f3hULBLiP7RY8m3MEyD7At4tp8Cza6fqB6mE24VVd/c9U57UmfXvaU/f/8
1LBAFRWK0KcMtS10u+7Y7DdeJGyoTydX2jDgCsyB9cIrbCBw5/kd6rbaoWmho/0O
ioaOpZqoZnHHbVx6rkzCWivM5UnO+lHVQnS+E9n52RTRbtwNfdis85H0pVufEy3K
u5IG4eaWRrWp7/U51q2Gtrr3ZofNutKRUnHNKA8qvy0vWEnHz1RJCM/MBgvJCjAI
Rvz6IQXWJe+tr2meHT2ek1IwFfrNaaSo1m4Yynb73xYoiPQpE57XTnm0b9vvvHkY
ZUpGSEsTa4qVCFbkZA3N4sEoSV5QrDIi/dceZD+KgIOQwEfdKuNMfQdeVKiQ31G8
LhLouyWjVWvr7u/CK/4J6cQw/IrF3b7zYk1Jas5DDJWje8oRWPhTETvXpqBXV8L2
iIhVdZzjHzF/R1GyEIlX3EJUkCnF7ISc4ourVk14zWcSou6fPbjUHdbcK7FD65gz
mBGOGDTcBqvBkCVMCZfEqvyGT6FFAPW6b8eOEyYVzkT5UAOFq73Mmz/9XpKd8Dkm
jZJ3jh9AuaQidZKxInLA2wrPOAYMSMui7C3L4wAq2mVSkZwAHbwYLiMZWeDg7rbp
v6AHdftB1bl8jHrdKcLMuHr7buLXJt+xiyMhUqHVaUw3IEINLtEcnAbFXQwsQf3B
dcxu4ldNILIBm/gvpl0zxuu78zK7JRGLFDIo+91jl4xhZaK/Ski9bAqdAODatNVb
+rEdLaCAZ93N0X1wbXdO93kPQ0hUOqja6dDBJN90NigAGE7sZKTtl7o2hxaWDPOt
jBmDbd3Xw4S/PWiJGynTesBZBc13zB31vHumxDCuFozetL4rdD4Cp+Esj7irz4IS
ZAGxMduU5JaFxXHUpd/i6gZXOZC0veZ7EjQ5PJwP+7XAwwGbgMy0h/h5iMzCIgy4
7gM1a6bvp4cPE5WXbagAHPGD3voGxmzVUkRqYRdSdEK9+ikRD5MlY7lA9fsovj9N
gKQb5qNmomyMdJi5qJkg6CH2OYr5xMR0wZJOidax0yGRaQNZxHn1rPRw7zzNAkcG
7pvdvisCRn9QKa35+ESr5G8CfVM64RiGvMaH8+4xaWzsmK1BOirPEwLnNTrdS9KP
k30LJZ+4OwNpqnP/KZnoZ8Otp3ZBl5xBZ4aV6L1fbh2EawfLC0qVcogZCNxMbUbk
FXqKmBsc+2JkmSOJQzlgfUoCJHjAzlUrMXFrz4mgAMS07obe/dh1Da06M632mV4b
xXX4A2puKeDVFbCEVIZciqYlrzDwhDYHsClWHEV9CVO3IE/Z5xSK3uU9iJxRVDgm
FbGSJSdbv8058euO0wMFTXkDBvKnc2ulm8mi6K9yvfvOFyGVvrFsqR2yONOO1mF5
kv1XhaTYG97PmjJPJalXS1a47UkWBeXh+9I0ixX0yJEGA03XtgXH9mriLaQYkb/p
QByX2NOvq3JwsRXQEAzC8QYVS8aXV5VQe/sNucP0hj94FEhca1KTxOh/OXgRivBU
QK+B21tLwxY2HkllMeAV+LlYQa9AzXtQUAWEWxoKrV74g2/K1lSzOE59UeUX7Evv
t7TXHVvR6AJ8/SGkjNeqrFlK49sZE2vTi+goa6lWgdnt+F6uN18D2MA8tDzSVK/1
rA4ea389YYBWpcWyVinNFzA76Yk4sps5B+w60B740mCNzk26a0vNIOLPPlpUlXdw
z0KHVk4Tkgtd8eQJhZoMln2ITmedi6jOPzEsVdoYFgGbW3Qh73C5ANERwuiwSMDd
nkFdUADwxuGmEBtmMkQWvXd5fGmtqtSc4DYTkJp7dXvD5m3zwvGVEPNGUms5zfGy
PXsr/97M+Emw0mbkwRfLCXfa91LReByBdnFYFIfdAzVd0SiRMVCKEHvF7mL3dIdH
hqxZC/bva080jqhrKHvIIoea0IQs/AzkXSxJJd+MaeNftdyXNhWyIYRsZkDf65Qb
Hzv4HuuUGoj9xhjFJEjCogHDOwwqUSO6dP0ZIY+QK2lfjRim8aPOuAybEXCZTZRj
KY7LFpwMm3pv9CmcHJ4J0wiqLcxZHYYQoKn4/WmwGnni/y7qfDt4I77fW5njSNGJ
c1XlFyJ5B2Ffp7LuczEa0TDIEKx27gYapdTfHdJn8JscImgqAr/f59gH9wfXtQWr
tMpopgF1jQ5jtRDoK+07FhMOigUjkdHVTsUCrSoCrRCaxJSvyzOhi8SD9fVpwxNo
N9JxnURCN09sDJah5/kmTg3/CedtXAABjGaTYhXkqoqSzJ4gEl+aT0wuiQld6eSu
B5TprzUq4HVEGrqdXPD1oFd0lb/aAu99662FztR1FcIfqWNWxzCVn6QdWC8+z7Xw
1RBB5bi/sCOFpFxSlo2GNkEmA+OqfzO4EDEuqc/IxBfQWabjQhS1mekcHJp9mbAT
KK3IVw8F5FODcPgMxwO/b4ztAQA83WKB8JOzZCOwQ185fNOp20f+RFqtVzGsDIrx
lX8UCFcUv1ncxCKpRmfwH3xxpe5rzGpt5yE07wEUud7rf7Kuf/SxQt8e6ApN+8GP
MlV0wiKai3ZVok2JxV9csZ0Bl64m8l7g+3DfAq7zPngkK7fp+UUIEpcfypvDs+no
FygqtTkSZlpT5nBudRHdKRqC5R8gKGveEcrh6NOxF8gj9ZSCfWQGifrfTOIRxAl5
XMk5Ouprohs5HeX64EgPBdf2akQTyVLz1mOEzI5tz0LLxt9MqD0EJVd+zb97OcQj
HmOzwYyEq4e+FC3VCGNqFGQiaTpBzfyJSi4ni+1oYE795rAeUi/0RxzD5IVqqN03
GdwxxK0+bcxgD7q5mKo9PKhowROBabhmRvulpN5gPYgLmrUmFI4lKGsYR2hmYAUQ
EjCQGAcetR2t4SiMYnObke4TvfErXKcKPPLYxKMWge57xwhvkG6pjuzFEj1zItXx
Mv47/yv0nMMSEo+waFe+iMnVGwpRjL8x1FJHMFMae31a5Bmp60BeIS7kVuYAC0cY
iG8Y/zR7dWHSQaospvw5s8qu+FpL352KLk5/Q7rMCU8Y7lnheWUpC6td2Gx+nIsw
V+UK1Qd6SXNvgQJduI2a7OJyNPGg0KNNWFDYlhjlLDpV+kq7t4NwZQfORjmlyPm6
HF/9f0bhNiOZ6AleDQKmzu/Hz/vmlKDIBUySfFihro9jIXEj2seG71WTidgy42Ri
lLShUZUzwRLkbNTztHcpnK2rKnTXo67U786V9imnotYKU989ahyn/CL3pK39vYRN
k4T/1tbT5W9vbNlwjhRLKUZRTb5d65oDIy4cx/tO243vwJws/Wb8RJ0j3Q1C1gBz
GOU8U9MDoHPPOj1dBsgTelRLvrxxkgdO0L20hqae7ljbYfyuLvVLV4G38b0foWLE
PttZocu8usUq1IuJkqOIVWfp4RbSufFRdDzP15EyPrQpPDaiOyZSARmBjHLl5bVp
MyKhAeR7cTJuxbMumTT1EbgoM47wHeE0BcpcaSafid9dnEHwAx99Nr0zPxezqn76
XIhB2Lw8+cv8ehk3mOtQQ79XGEC6JaFWVf9lnLSGQY8Bwtb2PK9S82pdOj48AXM+
p5tYm7QEQqE3Zo5V2Kvh5q+RW8GIkJnK4aaV4jITCWDuNp+aH35o8t5+F5LVaDfI
zzPLQP4wa6TZ4SDUYOfZsIbM6pTpmW1FChOSQleMZj7BR0Uvj3M5Qie1ETwV8ZeH
tRN7mCpFobLSKiAQnqXyBAO65WyyQP8k5drimB/cdKByQfNPFyb6KO7czKE73xvK
H8e/qjRABJV3TfD1QTe7yrxy07MLsvYAZ8LWO4aTEs5zmpW4Yxiw9iURbmsfEdLZ
wqzAM1ubEgIMcf/aNxzNCFHDUTe0+1P00lgKIoSWjdFCxZEfdf/duIlccWalETew
8mIhd8/KXlSSKSwcuYi4WLnqN3fNSaVF113Gn+gzD/McsYPBV1Z92pOJuIM9UEFC
2eby2d5vLEM3JZkwghJD4a/bl4u0GR6IHZ57ToZoxsvSz0WHyRhveFxf+KQ9wp6l
DJCCcrn7WxJhjp8zhxB7cIBHbRjYsFegyI9gNEaYsmFPxathMxjJTzv5Fn/40hyU
kirIYLd/EVK97YsDUW52vNom8mLslXxMy56F1al8O5gKkWjZfkfH5SaPmUI5KV3F
k68XS5x5/C1a+7ykW7LkcnKSytIVJV/0GJJUKFaMKdbOIeQfLQ7I7GPARdEv8gJd
pM55Z/O7O3DT/LFEMtFuBC7qkGSbY2aq8L0DG8n6eDzH6BILcjcj7iNejhkj1bB/
ErIRsw5tqI4MUuEirmzcyqYzpgMexMF1bgN0Kfi6fxyGVPvfFcVVLQ0lGlvOndqw
hcONWHjCdFqPEy7RHIlFDMLfRGImCSLm/7svOkoKbo/uLL50g1Xt6YvJxnoEsVQ8
lWGAqnVDWb4GQnUZ/xDy4LjDyCyDseDyid4ml1esiy1ci0PmZ8g8qdbkTuGO6vmL
c7X7DfZHrvlNDalNenCs8KnVB3dcgoSYhumALZ0Cjy7nx30I9ICnEnc5XjQGcR2Y
l8WrREFAPlo+JaPDqMK3SB8MyVwVgTofYUdK7+cPQe5i9ydJ1oTU8X+Vwl1w/Wmr
BJWhM8m7tsZB3CXT7FEpE56EkS6l/avdb84KpfesvejG6jfJivkgdsnur98w7nyF
cgOfZtl9eSwpWwur+x3WTlTwKIHYCTCyjqqQu5dYLYTPkKSOVCCQq3Zafx1HH+G/
56pLxzx8OpHhwk/xz8aqaRX/OWjnbOrHzfLNIdPEV6L53oIitORS35uObuBMguRu
yx2jQZ0nkNMreJJYtI6qdPMMzEtzcZhtlie5KpgW8K8twNEpVgvXowrAc7Xxy+0B
Ec+B/pP1mCC4OAABws2h+oTRZI/hvvY29rqpdrCL0byneq8ebgWX0/Z0XP9OXeeh
890XYqaD367UXIZlbaxo6nyxcKfVvsuOUbpTvsP43HIfshAO0GNOysv7bDErWsw6
rmIgKatzJ5XdOiPrAQuL6CcNb7MW9rgPZRBxYjBwopTe7X9I2x++GOeNFm9UR4F/
oAO1EKp7+QsPaOT52lFpORNZ22dDRlx7EL0IMnpxO4YoF7qt38kGv9p5UlsxNcFY
gPavsK1YKqggeQ++5IIC0MUCsqASWRP3KHrkBXCrmLR52xVGt3UqHaYaPL1eLy4g
VlK2l6lbaagjLoYbKuRX56jB8y9vdt3/eXnMU1b8RcjI8iw9ptdnR4iCkHbpdujo
A6Y5CXpKkg7nDszr4Jmp7YpP4I1Jxe9FS7AGSqdVdCHeSV/E8gsvPW0jlOZYMpaF
eLWdgA72+UYMLZ9XCMMyZbDO7QUk75TqB/aBYscdoQaTylE6FfOPPpLItA7rV+U6
edw04HM2OCPo8dmEQ1TOWbvS093rVDmcw3XVMOGPEt9i7BbVVfAZ04fldFYf5w3G
0gLQ/9SLCu3aFtf8uwlXXuG++jEs24DUE8ArQ1JtP6gcjhouRKLj+fb3zlRvqMrR
PDf8nzeR0DAk+MtDuYtO1LZb9YmMTI+rhr5uq4dQX1pg0zteNMlcLXTIEh/woH2Y
B33GIQwXi/UKATiNZaXct7dVOkWKfQctmBGnphOrkifrSmqzWKPexiKISrAUH52o
G5hGX4Mp+nRZ+aq2RqyQQm/eKOTjZvN7/htRxBpxhxnQFeLNa3cehzmfyFIc7o5f
miG0Tk2xzjKaJRtF2mU193h+1gAsvhxFYvn6Hdu0kQ8Xadspn3cXxoYbEWQupc5+
MDAOqWgTLvA5beYYIT0lUFsZq7c7j8tGX/rrM/1OlMCy4NZN2IHrCmSxJe4a/aM+
nV2uqvYg/tud3hcBAw/hpGZ0HZyUCR76ZKTYBIkh6Cl5+dvPN9PQr0249uSqVinW
hZeyHAvJyEJp31+HPFHy/yALPA38qafG5OPhvmluzOv5VIGzPB4FMH15jVmHGK8H
maXlbrD/FARxUKKuYH2/CTfF+QFSz85hcQsaFnHOObw+FLL84zda+g7zd1FymIfj
oHa8xxETrO4yaGs1Y8VdUdAYZk+9oJBvZDo5cD+1NPrDyY/FsuIaO3+SYuaEZaHs
mgDfmG3R8UGoZN/DFyFG7cLfMtEXqBy7AqziJd7U8/aT+B40DJRbOXVKS+BnalrR
mwLAqwdnlyTP/mpsCjjx3Ln6zKj3lKHGOVH9a8wHCpLOnyr09VkRq4r1zzROWvRa
tacCLadPb7BGtj4MkrelXLeXLk6RTZC0X0RtoDWfvq/t4xXiojhXl0OZijOmdO0S
67gPw83cnlRs5yxZKkd0VeXzQgXr5ZoAJTcsIyPblmTcqpi5Urvp1b7iQUlP9Sw9
Vl/lNy5ANKfwOHtS82fNs/ea5EHbsc/cUt1xjkniEyDQ2IFfRl8Id+mkb4CJQylV
Wnv8pxlw5j/LlMBUR/ZQZobNVwh0k3uQJ1IMicr/yNBeXsj7pFAu5APyHiUBzdGU
jPoyVK88qaKwdLhKnfPRt8q3SL04V7dgr4EFJSJvcxnY3r1sZy5r7pXRXJDmGz47
okbyd5bGNQBVZwxhARoihe9U9TlVQy24u/6GNqq2u/lv7O8AuVypZ//rzUGsrHbs
DxVKESjV1/u8mqRmB5f7qjRSv+mmzNrHmqHUdQrQ2RwkNVZylBJd+YvvfkhA/M52
FatSJAX0mN4LwGwk1xoMJ4VZq9xO5oaf4AbEqaoNMx94eK7PL93uOWPPgrP+fw4u
jBZjcOipUyf3wnqvYUQBmSScFsYI6E/ohCklQKMrzLpFc0H/PLCY0ahwRZMTFESx
fWLCVaRUgi6MGfVGxWNeds22OQkLZLo0ARU5xDLjfEy0Cw8/hoRzW/MIViEgIDwX
ZItHotndg3+BexDXX4pRm13lab8H4GKIEIh8yaWndpW2yZKHatl3q35cf18txaCa
rDnpsyypFXgAWlwmUZRqx9f44TgSq1V3hBFP4AekWXeIQpu/MELOMUzKZF+8D1Jj
4NcRpVxj5NVEYVUxQaXic0mj80nTmSMvcjgHfnusGAO6zFyxzt5yq593tc6cPu0F
JlS9q/i3wckzNO9/JSXxquAZqQEojXl6+Oq7JuVMvAGbfUM9aQD8g4sIAos0YhTS
tMwSCxnGDoxlqRSTu0piP5uR8YklkDHNd10z44V/uvXL5P2L3fQk+zGUm1wuOilN
53rAU6MrKQ2lqwcpGoNsv3vp3Y3gucz0pa+mN3BUivCCeyn7QzNYNclRTW7X0Rd/
8jIvs3JBXREocgSVI3CoiSkQ9lOQs7tcS7QOBrPT/QJAQuevT9FEh4G1DjaJYzZn
7qtjX80nn/TgAQUtL5It8g6gWd/tYXXFAyCWXR3rJz3rPeADD2J1b8FRiSeCprjl
HrrHmT5YQxioMNyQc+kOnhsyYzI+v2U0xMW1yMRArLgy9hv+aDfLQFCXqZK1AkcX
MzSu4vhnqcqJFoPGZKvO4+Wi1Bbh2rQCMFxzNSu1umy1YfgvjHv5BdAgnEfKFMlL
JhQwEuTM7oV9lKWOrCJx+G4hM6SnzDmkzpLiUANO1V9gqJghIE9u6R7dmouB53DR
JH1JS9cgs2ezJCM+P2bZbGPma6dKfdRhuemQzqKoOb8YGK0EA42/ajeVM5qQav5m
9/fp0BctHIE/h9SUSQ4nl3INRBk2KZdzZwSZZJ4nfe+eSVVTLDoCGDfRTdnBSk+F
3b0pF/A6+tignlf+LLnHK7adcg4qIp17iA3nIIBCa6cVycFvTIG1ZmJnehe1cNAp
DXSjCNNIhqONUdccjsnMzxtqWhvovYiAa236CLQZHPvUKqC1zfFEMzrhQh67KZGv
0A3uvC6IKnDslImLbuVRdvxPl7eMDqS0/e9J9PNqPcryZZfpgpw/8Z3XqJXJT8Dl
pt/kVJAHmb5NUGywOJDoX2Uz7yC6NAeQSFNP4NTWEp2aOns8DloARTB2NEdbcHvS
rtSbgy96YP5SViYRi3ghdO67ulk+vDPHX3BtvtmkxuCmr8geXCHBzW9PZxsKi7OB
aXg25n01Y7S6eDvYUKngo14RvUyqIzVvCxOqYPIUoawDXmqAeKkym9m004D4Zv4x
HdY58xhfiO/fvsP+E+yKL62wroTMsNxRNrNiBSQRWy5qh8Wmq5TFN8wF4XxVzsEZ
weRUUK05wuLKHQ3cj8z63dqqiSlsJmXM2kNe9cXadFLnpV5O+92pIjnkIFvqY8MG
PG9P0gxJV7SbpzoLSUsNHBIOhJHJji++wwgCNXTTeApiIyluIKVma9GfRbqzR8yF
1cLmikVswUa6jXGsJFKZzYqKaMQrtYFT2FlfVhJfsxM6l7pshZCQHMe1+7oQqMoh
+FdTiroomLQZbu4lOACN7A6bjbJXHo4fRORNHSlMYXgnaowQGNIudR08a0t294IJ
aHsFUTHZTQBGjFJ6l7o1gxJG53m0EujmIx2Y3D+Okpd60ge4GkDvmj/o5UfrepxF
QrXBzgar3b9E/FdGofJWWpjWbmUx05ma3ACYnzRViIv7+qllfb2pDIlvMnIpTC7+
LQHveF3kCdxdtxJJ3l/KWopaJXuneqqMUX6dU0pgZ4aD4Pp+9neEFNJPN0OXY5UJ
8+1tLE3BYhGCnCziOLTo44nW+ZTWDSDBE9I2jwmlf1DOdsbKMlrowNTbe4ChQax1
+M6S45NRlpywxV3B0e+Qea8s3Eh151RMFc89al+zZkAW+V2kDMXofnhJJ/MITgJP
fdImnwgXj9aL3ZqiZU+Y82THFiSi+uMiuART8oSpiCDWBn8ZNQi1XOzxPCTpqRHS
ij4Ir5tfJNoQjYzYKcu9t8H2SOpw9f8VY0rh0lzDp0tHaR83eZkAe+Mz6/gYPD2Z
txjjLKX8pkqNqSqPTBad7d0CjsVfHRNH3CwE0/gHHIMVnrA4uqVyafP4aJ4kvHlM
MLcokXvpcm6x4p5vBheZnGBDwvSOCTuVg0/EMogR9VmyYK5vgElwwBt/nC6KvURR
QX5+astKbJyAWZpHOirSUilIqoX1ZD39N5hJe5KODXyXK94GXjNCFwl5JagvuRBd
bey3ty9YIbpT89ricTLfuCxKRGLuqHxQ0gFKFtyjoP20Lh2l4vuWNQ3zd+qGG25s
eWjjYU+nwgHpMYsopIQmExAmgJqa2wrY2SF2X08zY/yaaTVwdQxwlMbUTFJvg67H
a2vgTClqbpGoJn8wIQazxm0dOyXLQ5Qn+my9FifAoDPEf6e5FpC1YqISZWbTiguf
HUl3vaWTeTBKwwiSx2JCPgwukPOg94XJdeXfumvInKtdRWtBSARwkwpDbKZEiC99
UdIsJxFy5iWbW9lUaLtGAtn9HJ2zRWzJ2nKZnu3yW2+VQv9QLIRPBVusQCz7RAq/
jW3anudUmvjfuXJKmkpyQtc2egES3bSGIVdZdar+ARDC06fSJIX7bBw4RlLKWw5X
PMCkHdtIE6El9KZT7zhJJ6NfFreS8Qh3IT7xpvBxzZkaEX4fo88N4lVQAxSANNHT
Flbk4HvtDIVTGKhQhcu7GmgZrPKe2oqxcvYYXTwQuJJwETCE3hTPmZEGFjUYDL6I
psun4/dI0wDcZMj9K92x7Hdi43Ryh0cX74gdNg3bI9BgUcapiwLf8ee0lcmXaHib
f3I7XETtPzkH6zoLLaxU2HXSyItPfF1CJb9UQ2HLNyahxyCfSkQtkTg8mhPN78Sp
5oJ0JpUqv1E7lGwwDwQ2tuPsVsUQCwjneT4Ap0wy97A9sAcmLETD+yW8y+IrkahG
bTx3OI4szHH7LBxkb+bJQ1NpfG/hx/BpAf+50k9znXAHGmQrZixpAi9uOd7bm6bb
28evDOBDo48gle0+DfW90mtOgIKwvUCOYW2A+eT3iKID3QpiEA4Y+6waiuXBEPVy
GCxvbql+qVBa7HwC06MSbHqQC2Fv94l8lWNI4k77l0vkgk4CezJyo3hQm5APrHZz
gHVVXlM+mx0fo+pdbAAVsxucupQyCEBLu1lcwe33M5Ue5uWUDeJRQL4wbB63FhYE
oBW3tEToB3On9lKydbZwqrXgLYBp0mQctM0e3PKw4FprFVeW24iOIpfHwEjsJcVU
qOAO7CteID/jNvsLzF1dnj1IVtwFQuEDi912EmG10ZCU8W0uSMPpJXOArLJGIl9y
PL/v9c6+4ZlKpC1PIIQtPQSmsdYwy3bhrCXpR2Z5hQs/PPs/AZGNjNjAcYW9d0Zz
chl+ChTerxpSV7qS0/LJmg/xFtjmbm4FrtJsiszGESlT6KXR0us4d4a7spJvafJ5
U54+Gu1jRscYVU1GMeJ8soYXjua6nsQt69W0SPvElMJcwJpkeM5AKWQ7DqD0kvJZ
a3wxM8ovnKna1Z8syNJaMaw/x19ZaG88f6qgUGeeIgo2WalX4x4fbtI/380IuYq4
QrJLiOy2vm3H0b8cZcNrfzbA3mY0G6iYkxPm0waxFI/11Dgx4jIWI3q4Z/uBzZs7
arQQcNHCu2E+PrlXtN5Qia62Zo1uSuOq4ZAKy2tfBJ57j9TnDjh47cmFAc8TgV4R
pyoBdyqw3st/2ryZVqlIy007/d48wCYc5IfSk5QqX7UpCbvmJ2V2AvD3Q8Je+ygC
dbcXthLc/lgVLRncUtc9F+FLGTpnluSX8R3KDv5Lp7W34Z2XuyfMnqdn9CP8camD
G/VmAiTYB+/OV3NHfa9XKcXAWenbLUORx9r3LzkTQSoApjFwH/sN7tUxPKEgmK5o
JJRmZZz35r5RVLRccyQSSEWbWwgnks8Snftbw0HMldNMYPU4w+0qeo/h/G5oRC+m
mH3P0WpXnN/9O35awXs2BRCLqBEXF49sId9ndsGdMkPfWy5OOvR0CgBZni3Rq9XN
1e8T+yTmahiPDTdIxbrkGvNsrMtJBphmI7s/p1GyT1zCRycP8i0pQLGUMH0KQmO3
5X3Xh93w9mTJkTLW4ayXywioldCuZ9zR/6ygQ3PaQRv+gfTRJIQHpmt8MTTVqAe3
2yYO4py8ueqwWpnO3XV0ERFCJogpK3uaEUVFma5VAIOZMhV0T7PR54ZMKeHfOdRU
V+UNDeWrb5yyoEVRpfW+T5xJqGwi+9JdGyzX73r6dyZfhlQIYfExLE4bevAS6ulN
olxMR1LPVZJmkT5vUr/TZtqwJklVhxX97y6RcruUsaVJPACqeEyZr4Z+llqnbpfj
2QQDXEwcnRe3uW1dveKQKtPwYEQ30W0lAXvZ612rUs/R7hAmmtm35buT/lYAqnjo
CHVIHFcM9Yr6h7//1efMXWqh6QNOaBFi4OZBxWjDHcQHNNaM9SLw6Quu/FtPEGgu
X0GiH2F6ngVP25Y8CJaELZBlm4RCpUh1TMEW6jtZTMrtSvhDiqKI2ow4rgU6Vk68
orgSyLoKfq6zpP96ivPGACrJGfBzaKycN9QHMz2FcEHJU7yaJRsOBg3GleHgOj+L
rt5UUlMK7KB6y9ft1y1LzIdySmJ6MFXBB0HWmvqGXJiE9Jqwgd3picdPdmDbxR2b
UURuDFlSBuBYs+h/4fHJMtxQ68piWitx6pd9Jv5v2pQfmbWbHL+Fq35Qp8YGwsHq
59MLYrRLHMNBQOk0PxEJHWlaB2XT9MYhL57NhtJLmC+mf4Q1jXmnF1FUX81DYT9H
4eyCpw/MFasicnB+MmmUEjTkNWtrV+qdAzrZ4q0aEiPUNzy/1vVvx7yrjX5FntHm
9dXYlEzobG3MGhTfCg5CgxXfBuBVH8mFJWsUwOgxbm7t7A7eA5EHGmPT2zhHOBxq
hTHuzwtZyt2My+KRXyTKYx9WRTwM/w4HqWio1FVIBeOC7zyLBYCjsCtpqY27fSz+
zHkA0pVaJdH+z6UKzm0IImuGYFBzEl6k6nztsmzz4yNBjAx7twHGDqvzVaDwGQ47
knnzq7w6Eyt0rmnDiOI1i3uq5N35llNWJYsY1D3y6dX/m5/JEy9lRyJux2A5eTYo
V9bBjY75Ooq2ReNLdzM5lagioCKOmmvdev+15uj+NHzwbLalh5DhLrlQJ2DcsyXF
ROhkuAs/xEtEMv3WCvuS+MeUhgeIjl/h7kRJrruq2pQbZabhHOoiQ3/ZhIe+a+1E
sNmib/shF/rDSJf+gnsiwwzAtGPrPRavUblVrDbWTUpa4C/vXFE97SlmJxMvFoKy
Qrm4/MLZFZd6Xz+p7VRf8E0Ov4mEjfmPsLoxwFp5KMvYxN7dgsNL75BQnSr1+t6z
gd9Pe4ZScFUQuYTUymSTh0Nqydpp8+h/IfVyalNyT64czzu+iNE2BX1/0wAgl+1t
Bfg2dpkGdCqc2xacwN63HFyKPxyCvwJ06RxAhiHV/fQy0i8ETBdRKBAwTrcEJ2/2
iHEgYVE116xaHB7L6nAoaUyTdxXbVnziRCmVZ9Eg2Mwiw14CHMvBB9i51pv64W/K
9gcboPw6KTjJYdTKOSuJUpEYHCNThdTtW9Dt/raluVz0erto/osGAONeXiXoiJBT
wknNSSHfcuulT80LpDxHiDH7TIlfni6VuXxX8bACBUQ/U4fQZY9AlD8w4NVthtd3
IRfPq44a7Tr6i7d+EoTam9xP+mNlEqRjDegAo2L7H3iwmJKnueqK9RXPrFylR7uW
a4UOrB1lFb7ov62Z9B32gJ+5PsTgdSwcVaJbSX3ZgvXvZEn/BlzYzrHUgXsvf1zh
gLvKV9HnmGrIAz49eEKGAwQnY7uI+5lkHaIOWuV7+tEMScItzR4VASkvycgMlzWv
bcS0myIhbqSZ9f12Q5cDQ7OBQIt+nRcwArMPWGk7kfTy0oI6KRoQdh0NF6F5CVXw
3R9loMFhs3E3/YCGR9hAqQa2hZJdlWllNNNV+sVs9DugwjFXUIm6Nkwt8pObSPlm
qNDc4/OxjNJ84W/e1tEC5+ht0SJrruWrl5vAe8SvdNekqPkn7p8jLsLF3ys4nvH4
wZzajTR3dcHdQEyIPIU4PnUQ/VAXRorHDAlZpXY03aEXc0bPUX2jwb1jzWTwRPXG
pxlTp+BhQRWAVT/RZEMkbnV31UwgE2W8Ajlxw6oHclOmtH5Rf8TyNo2GnY9eGA3j
MXUoxW5ODsFCRijbiixKzY6rg7hLEwXsSCDQskLyl7+fZSSoBisk3clW/DV1gQj4
abZeewzwXLd3uSiciB5LYN54b4FcD1++PAwHHvRQE41U88AOGMo6ynmjRdsX3XTd
MKQe3ul7SkZDJJHAF4XQdH4eKrElavQAG9+Sp6Uv+qbX5YggYqmLWtXxKhI0JVFM
BU78FHtkTNV/utzuBgclJJ4N+uDooxqiFmcjrHkij1V8v/Qi6ngkRgOuuVKWRPJj
xO79CBuPHQXKfxHnDWzKK5E23mNyYrmJLOwVssdM3rrfDmx/qeu+B8ycEXeKX4ey
SghqWfgRqf/+KiwGRTJmgsFTAYUO5iA+gSAsqvR/EdzK3DCUzbHh49lfUth2vAD/
3HB6irSfZl9l0nHmDIvYPiEPwqsa93avpzBRB/pXG7c8PtKMPDif/kCaZX2eQ4wX
v9uFv42SqF8NZX66bs16t4cqaHgTU68zsabQcM66P7ND15Qfwhd/1ogj6e2BrM+z
TR0sFTjQUSietxkRPEKR5rLawBx47eI3neWo+WrtK+Of+/RZ6vL9w48/FE/WbCb/
cNywfJya3Nlfj4Hhg7AjSiw9l4E+F29G5rSahBLVVu5wAGpzmnLUiepaNcP7jUN5
lIifoR7u3JcQgvGXtn6VbHghONg8TteLC178wVEsxzLjnxGzdqGwzZ43MfmJtN1f
l8VCZEWk2Bo7AZhBgQ/Kvni+xdBZW/rhhI+xl11yaXgNgxylmG4iYMtNkOTExkd0
J82irryd+fY1OBjpX6+GRnIqqjMpQAI2+kQUg4FblRP5cTc68YIDdCiBbk1fZfeL
7W9hRfM3Sg2HyGZxMVdIuMriE/SO95iTJgRVjrhPWXbF6iG9FdVVjxA1G19oRYO6
l1tUzT5O0qQsXyxcXvBRAgC7MS0NYVWfniUXXtriIrCiamw476tw3p8gusgMEQum
GSYsnoea1xVcBdl/iCf31vIN6PceWhhTm3R8giV7aV/UIlgpyda9A2HODC3Pkyhf
aljyHYOnEZE5AzWulUjE+OL6UG8T3gZue/U42ohqNM9vvMuXCmyQ6OQ7ht71grPd
+yFFw3HeKO8BjbfG2STlt6uq3QMEy/a27uG4qy3soe+91clzAnGho1ud0HiPSwK7
fKI2v0AKrSAy96i/jmvxOgJJYQk06Aeq+NVXnSi49+pkI7xHuLIc1/BmLUO+GM2r
UE+nHraezTXXAhLw7cJfOa7GvHBSGzsQ1zZCYkyR8rugMO34Bl4UMIk+rBdXB225
dGTPtsuN0myT6cLu3+n4Y/GzxfcHZniDeB/yo6mo8K80PW/v8dcDcLJQBZKDlFSl
3XPXPlqbecVIZonRIpurpVvoTMZjhkcGgCPX3XT9h/pGDv5dU6so+vz9MXbqoULP
jTZAmS6Sd9TEdpkkZWoargK/oRuu0+qa2KqyPhXPgTbZ8Di0ieKJd+hBoEvx3IUY
tBRDCuYgSmkSZQyZrGyWdmBUnIy8z5xkN7rUDdTASGeEJ5Vk+ixN8mxmsJ30HjC1
ssuGgcuM/fP+uGQy74km7Lxm3CSB/jXe8UhobF0JXjDLD1RZXoWEW0Sd/Ve8RVJg
043qzBcecffmIo/BtQeemxKeSJmvDmty3uxQ+BwaaHOjVhty4yIfmR0Dew9LPAf/
dEmqeNcHF0vUz/RsWCfqsUizkvidhdVeHpJ3ilui2q5slhRBPovFibDISMKZsrnS
FaQWfFikWn1fgM7gGzyM+IHxp8DFWMZHGyDKruUN4cQnrGjDXHO+Hn+k0JcabF+a
a5pmP4jE0qmchP3TYMb3WWEXyS9UjiWp2Sy1/jW0he5BNcPXMT4JBU0wBGD7kQnX
79ZL3nLw4IGqRUvB58KEWsiL6iz4dsx45MkD12Z1BgZwELr4vh2Hv8EqSrSTSdCk
0pgvaXFhDy1CrORgKbQdb4sl/xu+d04wHksUaSH7zN+HtizsEsBf3TFtXfSRMDEX
GlApsdlMSr9AXlMWED3QTgbtf/83+kxGjjZrbuiD95ffJndPIhnMzP9+9ylPJwcP
026HqTYll3gzELxrXdePrwLH0iWa2hqehoMK5TNeJkUsru5T7FmLO77Ir3QVy5gT
2OLskIwtDuF82VUEgXFNpTl9DwBiV+C2xwh391YJ5Uszo/QeTsbCVq4IfLQX9X/P
9zfgF/TVldxTYzbEctmBcVor7yuiNzN9whVpwHtto4qPyF+KsFps74/W2CnriOqS
Gi8UDrqDm1aAvVkLvFWdEhzIgYzbxmH/QAM6wKE27GM3rifys90NMpT5dAmi2q+L
h01HFE2z0YcS5cCkflfW+ik/AirO8rr5wHd5ErDWyp6KStDgu/plZmLOXFObbDy4
h2Sb2xPgE5cK5AlcGzCU6LSheJBmXQcKstkKIMrvglgfEPg7PFGX7ylT4zJvUc99
90WZ94+kOQ3iiiI5cO7Y/OaidMgJobFUSXBxCCnJfJ95UOu5HlDpwhGsn9qjQ/tJ
83Y0OddUeboAoSpVadK0AYb0gTS3aXVGyLANo3xdQ89cyfhMIDJlZa76ck2iqLpA
5KPTUcXJd645i7drBBuDh2XNtJRBqEcSAJ84voLRQEokgChDfo2/JrHu/qO72PHr
92e919/LvgPuRX3xcw3mzDANcwJqSDYoaHTU0hf3L1jQo36MWJe2LovTBqLuIB3X
frvsbi37CUuq6ao1p+IuDDsWehM74yULhVX7i9MshnLvpwWFuGHeqAYZCLTpHvHJ
LQxhDpp+dKUECsybHj+Nlp9cCm9F1TlqtvsDRobWoZbmWUB+Gib9JXDmSBK4hgyO
LYBTChwz+rEVVQIPh1XTk76zAw7419Z0b6xIPU/q+ktsb9NJmsgK9veRoswmSiWL
fdCcJaQ+fzqXX3++X8YyQ9iLf0JthMluTPQKgB7+nE/FYsVJo/fl3B6prf9T+Try
tBd6JWKseu3NUlh92kiK4zpSGgitt25t0Uc81CMoWdCJHLB8bLUVJwvQWXkpQDly
0niIZQG+aNJXBldKqANQgQESVmbUYS+sA/X/Q1Xf+gn8vpoU1V5fxO79wWzGgkB0
i/Kzq3h28Hr3xgkU6aiyNZa/uwfeBwwh296l5WkO2x2c07WuY5az4ti/7HnZN0yo
wl9gcArvFDkoOE/ywgOopulkC/QYKQTazVpM1dyNXkP+Wsn1X3DyKji/8VveDCLW
xBTkG5L7k7s39K00bF0L2D+O+p1AlBNN1FOeQdaG8leh9ccZnrnQwe4CA8K/Fvpi
tL3Fb7GO0/80eC6hNMYHuzJP4v9LRu5PC7HkI04IF53OsT++tCtv8q5SuAUtKumx
3nmxzo70gBikAUs6qYtKE5ZLgpnYeohLEeUEpqTmKIKl+EvtAoe5f8fa/YTxVuiI
U1zxmC1oPbut4tRyXh3mmoiqmcsyFzhV1bc/ZByCjiwGMVMNjpfloPwjGXXyNHId
S4neRI4I6CH+rfMaFYP/d30kHaFS72y+9K83g3cpLzFqvQWgnDlTfExl3YObswTX
S9LkRRlfItQtWjuF6ngcMRkuq/QaAl3LPtE6kzYjuUkNLmwvF6C9PmtxzV5Fr4rE
pm8MQpr+7VQlAgrMAAd+Yhnofj7ApMRqT4nBNdfpp4gQ8+60ooh7atCJ1bvYan6l
Wu45gt73tvRaSalt4daF2YqlXBmiE+kT9YabD3SFtVbuC4m19Tp74TC0R+eLyExA
5Rd2sq72iF3jHo7LkiLXbOblGh69WQhxYHE5xE4Rlj47rAeC8VHyXH8PggULFLCh
Ud/PkoOzEKjvkNjkbskYq9T4orn1GngtQgxpO9bUF90ZREsyEwjpdzIm+mrRJQwk
VtDSKu69GLu/EvnE4ogOa/tC6HgCkEunXisH++hjWIrcvBBHlp1Qlus/MVhtGRfv
5zd+B60eAzch+U+dTsBONg7vQ9kHSx1xX7Hj6C90h/zw/W9rAsjnutSUww3rN2iv
t/aItkgdd+zAn+sK2ERrdniZ3lIVs7+DT43yNO51/OTmpQcW2kDQbKMuipbvGAi2
DhtCRgng8Ihet7TOY4LTpv7K9D/6XAr41V7oJy6uHknbcrXs+NoDc0rrxxAKBj8E
zY3HESAz76cGN52GzWZ34DmRbPBMRBLSTojTzo7znVFCpuXPmSwmCkynAUGvHG+8
32vN2HnCPbJDt9P+KrfN51HVUGA9Wl/s/bY+yAA14zVmDbRUH5MnVpzvJC/e6QNC
pbQvucCVASEOizhKAcOZhRje5FmgLDAZLP9FTjM1/OmtUBtWNAG5sd8Mg6Hc4xjP
02oSkZrVlSAozhvlMIEyeL3KaPrmg8hLDyBGqYHWumOJZ1Q32rNmZzJJ3DwYngFw
ASzyjGXpAbpJfVP2sDNAn61ReFNG8Pq5Lw/Y/OpDR+WLpUpzYiNtjXeIRFGPOxYW
vPHpzrQMYjJ2dE+eaxVmhSEqg1zbTFZ6I1z9Js2oibGb8entjeP3j2Vd9zKwSrvR
zN8m0xSWnLF0IBy0DE1KtknDIpeViqbd7EMpE8RPAuNmTvMFc+Wj59tzny2bNYg9
Li9yEXOOqgnvkhyhdbeWxMfgIzLyyZvsDDeMa0yRu7sL3ePT90+c+nrBDJK0FKVY
zIm9og3sbv7QC6CnuxDBwVZaJdtKk8bTXQjz5dF1VQdMNcqWDe2D/gFgYzzft8oo
hv9Vyepv2CoHZhsz5WUOMjwZBebyVZ1KKPQPBPIybzMUA1GB3BMRnr8hviVfJrlh
KAKytD3Vt6lGpWnuHidqY2HW4DxzRZXadTLDeEmGquvnxxNh3iVDHGG8e5tL8RsP
+ISpelQB27NRef2kJamVo+CFjoKaICCW6yPH+eqrXR21AK9w6oxixQf+S2xjkNUw
bjIqkK8wMc049jlTvatXXzlJJm8QGYDDQildDM4LKd/WsYgbXxVROfnmClxPaQ2k
4FO+QnPgt49AiPHWr2EAbZu31EhzJkxZg7ca1KfQjrVqytSOdNu24AhTNumcwJDg
hVCCW1cY/A86aAsTD2CjvfvG9tDe9Qvxs1Hsbg0G98GVuXRHxT6S9WFIPuKp4caJ
0xdeiIFc9hGuMiP5DxM+2E9X3KZdNUp+P7zDjhc4475Jy7shRJ6RdODZJ38LvKBG
p2sdrJDyLZ1O8soWeNS+a6qQskYaVRefJYnBjh/3QCofKC6VEs6oWf46+uErFafe
iF6yT6+84a4cT49FovvY20gkzCbQpk4JCpljk9gKjCkCRwUnAFQl3I9pfjEqgdWo
xyBdNFU8w1ubkI07+2lsQb8SIiGo5KBrLqvLTlAUQdyUce75Ld/XOQYpajCbxX1l
RcMdQ4SO97JfPnEdX7Fi3Th7l4OCSX8z14fmhz5F7ar69otpi+6FDnBO+hes0V3K
PCJkTgWzbF6LCyBXuRx3eInCLO/aHvGDXZP2w3vS3m6KG66dIPMq/DyVUEoETae4
0tBXR9lAgMPId7qqKuau5epJAwnTmLc/DnkQE1TzYyEpTbSed+keS9hx2fcB77tI
KaEoWF6796LWxaW2XYsf/52x6bJ7GvdT15AgLsrHbMBFKjqtTdZvVb/wbc7dhARc
Son9r8G/CUjNY6O9ov0gsivFPPIxNBrfMkHsragjEXDV7JhR2091tnqeCRDur/Lv
SFWgILpn3u3ebj0JWSoXY1kPn7lOPCeVPd7P/gpziqyb2YVh4OzZlMtS+wgNTeN7
3m1IwUt2Qn8PNiFD1w4tVI47HPncg0BzN37u850EmuHawlfymZnYOsYd3Oa7xwka
XtIKOJG140hLNbNZmQy1HlKO1I7AljFFK7DeRr91RHnjK3ROrz/ygArHMrW0Zb/p
lH8Bng0BQF0icpq9Nm7sbmZvn1FxMnguPqt/2jLQWvU8L9433MeKDLRQFAfXRPP/
1+Gr/lM97pDFNu4YaEYpPHdeA21n4MtEw9ovexvlRecId2Nm2dowzZmo3EXnN2+T
m8fjV6k8CAp1D9cQ16ZUvhDED7thCa8NpTfSYOXxdtPjm8ZfkedgVSbRvrEZQ8AH
5vQki5ntk9CZrSmxyHYLG5tVb2El1DFkJ95ocdD+Mm8Wl/MKmQwk8UQjubH3b+1q
+heCm5KqPp/KfD3gnp/LgmD8Ud+sNb+ARS4h+cqudBVrGhB3L2zSdvvQ8pELmgU9
tsugISUmwHvYW3EcDC5DVyX6LmC3CgeFPUnx6TMJQ6hQF6O1cougK3O835k7bVt2
0FjB1hdQSZ+13hm5aH7tvz7Xu7LJun+8vM0m31fzN3I+d48QkqbOBafg39bmEs35
dgicpE5iz8Yv/SLN1TUACqJ5X+aai8AhATyTWs16VL5wKHxESvP4azDZItoDFBTh
9JvusOv7OzXYiyP53O/jfx+uJ2QkjIb16BEBV4qxzgu+uwXuCiWPGU7dwmwN5P/3
iDpmtBUtqrb3ezB2SXp0ko8Lw/vl/nQ3zK/T0texV+qhFDPDg5wjXvpqLrCjmmMU
HqoEh/BIt0Fk+aSWaSiwl3Mf3GMMrfTZc9BEEin8RI5jxcM8Qugh2oSoayErR54o
PvRf/pIRA6IzRkMCcUv0H7+4Dd7TJ5HZZ+SFAdUGuO2xLXW+lkwlpnYpQD2floPD
DcEyAtu3yyEvR8iJP7zhYNMM4fVARaHt5+BUvUbRudkQ4E1c4ejjOO5hiKHg4qMN
RLSvxi4/1knj+5hAw2MIiJv2fjvqOUteZuU/KPHRFRJaSW4p/j7N40tBI5eMHQoh
rEgOA7RTnx6hsFCo0njUxokP7grbCGCWmzyP0TbEI4cJ6bL+PTLloXSfFh/D7eZk
m1IveKof2TRDGN1aOTo6inWafMkDbxyDkK6fbYKtm+EsAHyupsNIzPr7/Yv9sVw5
vlWweYleAufxR1pGOXGGMS0qq1fPFTpJ4IS1M5mekJld5Jv48sApO9DKPdT1EISi
/tJ2oSohH5YPOH4NXgRFR8LzuRVoGVKkSw83HRTLI0bRf5joLKZi9WKCEavHD5xu
4KyzTdOrpg8Dqbt0iDFkk/j1qetds9wsOJQPdkS7sb7MP3UBU6bPT4yK2AJoWyfJ
Vgm63Qb0AyhrPnihBcMLQhXUPLo87mSBfBoINMvfpjaj8htQV4j9eQec4tM4dT7P
BOGy6NTxgUAW2ZjRTQOxcE68DqGbzYSFtmZ0/kouZYatxzBuwXQdDZhbkolPEyGN
hpxad7XpP8dMPQ6RysIrwVujeVLtBcoxm6h6wNl2GT5RF0KaIuHZyHqo4Zp9Qw4K
yIG7+PddIsR9jHA6f8H7HM8m6muxXgfkXwGaIlUrpLMJxJlqwM/btU+HVqalU4TM
jW2+9mU6J4c8BYeSABudfrj2Kt32X8TCbelH6wkQ8iIO9mPXrGrNr/vFHDPTM3h5
0Q717jBNgo27kyI5r0sPOJQVNlD176RlgT4NFUwNnHMcisOPCollB0speppqU1qB
C504gj1igGTOQzuTzAVj5nLVX7shkDeQtW5Fj7NHx4xAGf2ZazULuThewIOtCtcn
agNGaUfWTa8XYHA8+4vR6kGiMvRJCSK7nWRubrEm6Ek4Lhg8OS1hqTYgkoisxvQA
f7l87URsip6V31U0hDF1L0kSmhRkYQnDVeYjVyaOT6LNTEGUJA4gkxqwP4J1pX4/
qmT24/CZONIeTvcL7AFrNrw6CfEc8pl+IXe++FiYE5jZHR9r2pDsiYlS0W1SGOWn
ZgFqYAg+zPXawPJw0xSlpHTDyDJSbcHl0c2qZ2UvTgrEXYzrR4NeQWYKvYQSfcOi
0tS1C/nlXlYULxm5leik4HBjzoBMxBrC+WlN07OZwB/7Z+16v+YaB6VNli22C63K
eise+IrHfwl98sA0aiMUHtRBoDlwADhUi9cwmj23cTltyK2tVdfqGOpD78VloI5Z
pQGouQ6KvmKyM/e3D7Ge4eWO6pu52BL6wXGb2vJzLFplu1LUtB5EzyBeagxaq+UN
ffpB6HfCfKgO7pXu7wKOZVgeSD52syLOviLDNp4X74vGQAaJ78ws/oD1H0BoUGrp
kinM6X63TSCvoeuwSWNo/ioKs8e5yYA6ayDsUUVZzvXex/BBckxAe5jE/mNnDLHI
FCiAc8HGQu+++dkR7ET2mX1klHbUVO4cPla0LXG5MA5JopQn9l163fPjg7k26S8H
HIV+AgC237Tf5PFBl7MdazX2rUMjyKT9ZTHm0yOeYDpiRzKb3/hjKWH2wTwS+FZb
zIeUFVWZpeMNTJF9Zm1DImJhnr4FUB3LiuGZbgPa1WZ30ap/B+AoqDgLrFD+529F
05+ZYNEL73T2577ffsWvLBeEb+zRP6ODcGsEjQshN0BXDF/KP2WxXbtsBCnol/9C
luWDHjr6oZHgdTqUika+cArmGN2HecbH7xWstpVr9AeftdGexnriwuXYekns0bvV
zbstcfNlrsa5QhUvpNzdhn5ju+VhO7ORXMZo+0yxpWBvu3gvN7aL8bDh3qCnljUy
e0swN0Gc4RrbWK8s3w7n6vGvMJgz5ikrU06arcxycQ7PB48XoERWXwidwPqhrCM4
L3LCIoaurnbsf+LRYSm5unmmN4AedFhVAbHbrTt9973ouVqxn2WRB7vcKUzAbhHv
5RZoV31xGhloNNn37+Q2kLygDwmiKTATXWt4oVSYtW1RKNwui6wlyvtLAieXupdr
bkGpX1j+wlx3x7kTNCLH+EauzdOzdvkBk/ZT/SHkOIEChSYf7L0/HlY97pL7HSS5
s+2T51UmFAEr/n9nH0HIGj3i04I513HB3d+lbj6PRRVqELijkk2Je1ugXnMKFSKJ
pIqF+fes37lXdf8Msn5kkNWbJvto28Emj5+wuK0uorb/2iRn4QQFC9aCQ7rYoVM2
Wblcpu4hTudIV/VvGrZuymcxromGvNeteaWF1ODTVPXi/W/vqqT1bUkt3lhHpsrM
U4KUpYq1OlGAUKS4kBTVoHZkMS+O+Mxs/LUnF0aO/0muz4OKlgb4reEHiONjPLUg
WzA0DLy83CN0l8j/F8bQYtpeQAXlPKiq1FafFdAAw8Cr9v8MgrICgG8kXTWQ/10j
MAPhuIs+s1z66CEsFtF8AO2QF+l5+hSuZCxdWt/VbS0obwUW292+HTXWPQrWZRUj
rlsTFkHOXuP95JlGWKBBETEFm/rI/pwGQB1SVXTiT19nPd5aUJ4hVnjLobfPdZHj
t0K+cLf+4H5kMKjq74IO5DhDUMIHJlGLYmv8TSXCBVyUff60N8BqZkT09pVF7RKV
LEt2dQKSpMO6VKwsOVp8D/RHAm6jTi6s4LngdzJtWlcihb/5ovr/l5pfH41cl5w4
/lkXALLiznQfHEc4+kucKKJgNYOP3ibJGjL2pfRG0vT/eNUf2iL0bc5MFmPGwbHG
daRBn0XlAkBO7+EaUerbFPgs8lO0qsuAOKQbSAUIGKfZeXAJNbLay8bX9hbQnfxL
r7BfW6QesXMdriALBw7zuo2A026zjSsIPyv1tC71h5fARtZJyFE+mhcr89IAWX6u
3j1ly9BROdxtcfLntc4GLm+U+xHaPSLNDdlD5PC4UtpbDGXfvP4fN0SLHSHcOH8C
SPl6LoYZi6Y3sbwidYrt9qLGFQVSSjsaeNdh+vy8E0scFqNbhnUaTy99/6p9uqHm
kUw0kqrtw7XpOS5qFku30oA12qa6Jur50ht8Vau2gOn2saak15FKb01H1O1ziP0A
gWngSUx5l58JN6pRTtMcId+a/7St6uQxVozKH9i/jRkLNus1ogekKEX7qZ8tBSEh
q9rJmEUbP2v+BnBTEMbR5Q8Et88FGanXrjVXW6vdg1qo31Vug9twkulEBcNss9zd
`protect END_PROTECTED
