`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CfixtTbX9KA9XJPsOyBwMLYxQvdBiX1eRBLOTEiAYeQlCWRuPw6R7yvU6w0f3oQm
ra/RQfJT0Gj6OL/AGYhhlfDN+ireeoW+55QefAiY0odNh5+S71h4sIROfQbw1nQW
5QCgVrB680Ad56qMl4FpwN948p4ynjwcKKv2ETHDAXE+Zbc6422I6+1m6eYC3dXh
uW+1bRDUUL+vMBtjHl2+QHNw63o9dTEp7m97CmpQTmhVJS2jBcHZ9UAeLoz9Vfuu
hR4wD5EUXrBAhcAZia+H3qfBK//TcUFlA00tWA3l8klBhdrrFz48HLlSZDskyYV1
GA73rHkvoaKXPIRbvlwTfkVeQzIOh89a9xBKVHHxy/5wGcySXlNuCVFPqRVl4Qqm
5X2khCA+8lcSlbtsnR2VLD+bPDCmYCG6yMa1rSDgn0p3gKA/tw5szA6b3ggCG4jU
IY3DWamoVB5+pMGoeHDKuDUKmV7A4+PQUxquhZgKYJEA5styNOihoEOTq4a1js2O
EgTTX1mrLx24JY4zUCKILBuZsqOXdI1YaZsHvw4qmAUYmRWIxiLQqnBRug9CMR5k
3A3LLQ3bWtHnnm4LMUDo3sqVUGH4jYwcMx+MDwKHafVBHInzHUOUU0I/JEKpjl15
92U/6rJZXvlCBujyGRtwGSI/WVx9XOK19YteGUi/l1M+qgl9NnHAMbWE8oawHlJu
m5eYVTUt68gQzJJiV+/LbyBWHjD9P6heYF2QSTDJECqh7sxbiqyVyHWcNqwdy/9h
2gX2nDwUZn9il81H5RXTCV2/CVgXxxYn/KARsRJBn0pYp07tcNUPVhbNChPpDsSw
mBh6Q/QRFqe6btHcF+Ov63mACnbhPtmgIg8nDOAa/Do3Ue/RjhsCs8mBVMSea5Hp
I1Gtd1Vm9KIZYmm88ngeu93G9A8umbyobsFEJu+BJZtDwo5gj/r1zPp9pdhcP0oE
gVo+QiW7xjxHF5a9YqC6K+aAibdOub3rlB2yhvbX/p2jLvJghU/BJ68KDztg7AIj
Ib2MYqMmUpq/oVIiybqh8hLXzOYTFFSiImITt7miU6UQ9Qwh7H1ZOASKxxVflhR5
MeDuBXNbL1nnEYHLlP3kvAg2Hq0NYxavonqhptSg0O5/qk41Ltho2kXdao8rZZnc
P1cf1X+tdFYew8Eysm5Euk2hL71ZxYwb+kK4wgoTTdo/uFf16Er8sNbzX4YNcV9t
5DuuRJMm+BMj6HsdaOMH4DPY7dVW+FBxhDRv5vWJg+SR0PzTXy2s7NgnrlacOafE
PyTD+jngDVKLWZEhotpGgsDpUvijO2CrafIExacTdOu34rqrRPppj/1lUu2oUMMM
QRyPTPnfWe/NqfU9LQBKXOMw7jnkZ05/7XcNj6G2/roRUeo7uNSvQRLRDANRbUDL
iHMOc/M1gNGFvMxkvvjiaPvYL5qgmRsSxRSw9KuTo9KYyKwYTey2gro76loAEr6D
MgxU3ho+Lu0kPnLo7l5a/kMLnUYEllMfLv/cqobmSzLAL0B/D2+QR4cH4RiRE8RP
97poxD3RHVHoWrpJlm21mhkzJsiVtasauIDrf/8LPzt5jOjA9f2EEuYU9uf/uIL8
yFVl8Hi/v20fInu9E4MA+LQA7DOgN6UDK62Ge4vvff4IWIt1VmnTHnTOodgSSp6w
q/rKdPqwwvbqVKjuCtINW7SkvGztpFWq/L2nBKyPMudZP1uhvnVb5q6A4XngaqlX
Go5KqnkgsPynpggGsKvKVXcSD8zL0MjzhN8B/LQsfVHFJmmZyQIOXr1pSdKCGETf
M8etDH2Lc46Pb6+KIxqs6gCPQn0FX2Gqt2SLTrAZxyAMvC+xTBEe3HzLbqcz+9ub
n5aS7PeMvlPMNRQnOuKEbhbFGrBxueRR09Jt5fZ3JSphiUVKBx7g1fWGagjxvkGo
QyKyMH+lSvuMLLLsCyfnJmQyF5OxAKI5u6XNYJTy4+tTm41Km8bCMVEKeOTG64/r
0L1SODRUqpqk8+1aKOQ31isb4FZSl6CjoX8kXVJONzwBMxqC807Ra5oYZ7ZVscdR
lkcUOTbQ835b0SNXRo4gyfeOVqHipWKAbJV02KSbVANAjI7ZhovqIuTj/nTFLqbT
8hbyj+JawbkEOg2ZtW0GPT4aJEzTSeKm9LQOQm+lR+njpvEOctZ3RA1aagURIBB4
Y9WEsTVPZUdqXsgFazcycxUq2EG+1lOOiZQ7fgx500Jm7OqBzoUOtVBxKhotRJkl
3NOoZ+WE/BeS6Q93QjlSj3Wz9hBIkWxxnEIkZvwqw5i074uqtW5w32UoTooGvscs
Kb7kLIh4JQ2yrZAWL/9Mvs+0xxllG+sw0x4+zpPR2EUgK1s/BI+B5OGVnt0OIwHc
9m6ombyFzuNZRFF/uT6tz3RcGP3OgXqR5ihqmAw9VNKhcf8O25tv33CyvYzinhy6
mfCOEA1iv3wkRf/+RFAJOWVL40ICpNOvFfiorV7w8lKlsktkActi0tm2KAsSdn1x
wEW3Rq1FpID3bYqmC3ugjFhmS45Uk1YB8B7P3/PVbiRj4zurnMxVtcfNxlO0pBuF
7h9SifAKY1rlFe2YwXGAoNhYyXQQj1BVBvAuD6tZHzbAnB8da5h5lxJCIars+633
BTdOcrBfyTa5GZKxmK7F6gWnLKZsuCL3VzKKAgSDYUS1C3a2Z5xH+VQuwzwLZQKj
tSkLu4mGtEbXEz62NhoyiyQwWgq1+ZYQ3/f/3zj7573vQBWjPoU0hikuMlUIiVlK
MPweDMWpsQMjZFYtdaise3XnLLOVjc5MS1bl0U2gIoXqIQqZN6O0FEdcF33pjYif
MJUTdMeu+ao7kunXudZ7xFlWoYpTaCHmXAPmaGAa2ZYW7zwf8QCg2zmuI6Hg4DDo
01G5dVecq133eD6K99rr+VynJwvEOhKoFmo01Uko5R6KhInK5A5uJlm4sKG1+nHE
3ty+XGasNKbTBTR6L1jv/YE7hhEoEckc3g48qNmyHa+AMpDV95/PCGzvnEfdOIv5
VfsFdxw74wZ0brnPOvD5+uZ40O0Tm4dZXn1b6LkHojNh9+qyARsQSn4wcAk4Y7Fy
gs4Be6fj5BOk+RioSxoXUoAHEmKoowDeujb8mAUhbD0ahFkFlOzKmLFHDIDcwSRs
1uwp01wS1mKuI5+G411AG97tuTDoMs1Co+IRP0u0UQsWM5bB0Y/Iqguwo85+fEK1
wLbF6xZqd+Xj9qj4aEP4otItijfkF70UKAYQaTV5a2lWqHuZC4SOaunrmXNikDmO
G6oaAiiqeDcAmjGknNln2NbZyGTU3PnEihzHIm3uOzaatq+ZtqnCbcYqEs4ISOf0
YIRrKp07gM2EEG7KzbXHLEp0B8L8168PblqqMR5TxOv+Hzg6ammy9etO1jBiYmcN
KufYv4Q/xKVEVr7+ap9VxtyRjyJ+uJBuCU/5lZQjA2g=
`protect END_PROTECTED
