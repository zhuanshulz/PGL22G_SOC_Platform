`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YVrimSdWafY1ZlQ5uYWuZNjfcCEawtnkRTdCA/G0+Z9Cg2rW3WaYH99xRkp5D59
cTweJkg1HTCYw3HbOFpQPKec/lmro5ytqRELg6AiPmSP73q9rJyijp8btgJAi4lI
C6DKaIFyTYj8AMIJd1mI5XcynsKZzMJV/vICbqt1F5ekZW3VZatvstroPSicM3sv
1e2uiuawfA4JUfC8f55g7wSyrvt6JSsEJ1q3gabtPmfOyTsvMDGsof1o1bAgBViZ
sKUSQd34UChuXysDLuwMMYBt+U6DK4kJJqG3A+Rwkxbx5Nat4d/9qaMl4KNZDuZq
kCR7I+zhV84MnvSCJp8UoC6xwVeFeT1E+EAvqtiVeE4iivMS3rTmxEflsDN35AA1
463C8GzEkEJGKwxusr+0sgJFayiol/r+9Rhs5SntNd4JtYa+vIFyE0LGjCzjIikt
hD1ageM2pU3ug6zlMQm7tQXyKzI/WqU+pVNwv3A+mkduAbj2OZxltuXrv5JkP8kO
z349nP0KYuIfYAdyHSEP1Q==
`protect END_PROTECTED
