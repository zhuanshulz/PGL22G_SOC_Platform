`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wyVTfFc3QWXjABODG0un2yllBoKX1mG7hiWDJYQ9R3mTkkCJ1YECtsThxcpj/4Tr
zDCl1f5ETsdnrJKsa/FdAlFSUU3DB5EUL2ygxiDjNoF8I6NRGbw2t0rQhXrjBhri
kVvP1iCkKShnB9iaHC1P0xDdGBGERO22AWg8QkSSwY/26PwPOWjt0MGSo5OMgmTF
WQOo0imgDucL9NyBYrZoNPzxpMjkbzZH4miAhYPm5VGYqFYTU24NkcVA4dqch1Ek
jygiTFHZGLzis7HBkuf22LEhue/j7Bl39ap2ndG6GttInU6HUNzPSBAYs1kH4w9T
ZVR3sCP4QbFLEr1psf2M4cie7NR6tpOk0YPLRmawhC9cSRRCyAta85xw+AoNBHj4
MCcKcdC6TowAIFYj+VcOX9wvZGWDlaHNnwTqSI8bZiYwxO/258aB9t8nyoumUX34
AW/giIXhOASXeD1YsSXOzf+CcsCo1NbTq6HQ62rBGZhp6DUeWHGq6QqTwDxlNAeG
/mkDec3ASn3OM7YGuleQhW0T4b1SfTNwPv26ZMvHSJSYDl+rxMGl2HaqbTy74HHv
N2MECRTOnmFaEt+wte8HEbIloxcsFG23g29n7hywApi8i3x1hAz2G4p3bZrUH5FU
ZKtIJ2X+cpz9ve8BsiqSr3KRwgcJGhyig1g4M/F/lV3VhjpvLpyCY7kjMaueJFZQ
N+vLD80kY0kTGDYeEjpCGC0w5hue/tijSj/Na02QfG17rzJAHY3/9N7mcqVvrnZt
`protect END_PROTECTED
