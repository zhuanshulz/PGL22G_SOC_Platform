`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Id9ETU5bfZambwiEfrqqG82goJFYA4mK3NqCIy1uxte7oRHYfW2bkj0G82AJiabO
5uLLr5bYDI84M0oibNCkycx0Iz31I/TIZWGs3SjL1MsLbRMio6UVX63dOYusqX8m
D6fE7MHjowGqEjvCwszUAf9dItILYPKTYiA/5yDm9r4a2mZYGRW7TI8xvFP23Hv2
3DiH86kHsMLvZd5rE79aKA0kZ3eMrvddSWUlJuQIgq3QP9cSVvnkE3ZHRZeh8eld
RqcP9Re/5k18EGoKudJvNF2X9Th//bXG544SSxzg65/5VsUxxGxu1Njy5QNf37Ma
dPbK5cnLv1isqYoCwj2y1BtovhZtI87PoaSkQyn4nzsxay7urUzTDd2wd74akClC
z1aaCM+MfAnJU+pI8JBt/06CdgQtwp0VjDyrRc4fiNIDUlY7aD8LoGSXUCwdjRGC
7wEBrYN1x4h5v8ZYxXfmHxO9f7tEWSAeXUdkHZ3zD0DKk55ztEtTr2NFDZrvueee
8XG6sDKGjz/AMiecAR0FJDwJUoFuIHGevCo1Hx2GdLQS5aLgWox2G+oLSZmr0RBW
ZnrFNoYOE238c0SCbeUoSGqy/PJ/jPCCrImWvz7/JetodAgfUbCpbtLVZ+Fo04jW
je03QnhBqHXwl9X/8sZAbwUj4+IQqySdFyOhuydEfWa68VeiDbODtCkNhQVyg4hi
N4wvVeoX7d8exkHZBjYNR3Y1El0H6xi+LLkMxtQ1Rh2ih8lsNkdd33gffl2mIoX5
akPw/kTbDDmk0bz9E+KhOnW/dsPYYESoQCD9zOZnRyK8K9h+M4lTOLmC2W9bx03G
`protect END_PROTECTED
