`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHXylpHeqIxqiScOmy9wbs/Ib45IIs+1xMcZcCGwauchtMniT9PbvrNxb8E6AxJp
6klH68Pl1lBZp9Qq3mlsLPaItKe4SC6SZ4zVm+QcTdo54/Jk+jeOaAtidTvrh4vZ
Xl5LRsx2Zyc1Pm9oZcWbskFKcsSxSJriDthx3lK+pAKGZoOnyRecqPaEMI/E3iLu
quMYBCHZSSMqZPs3Xa0YaRyQjaXCKXwMPCn3V6Y1u3KMBLqhUJjxX0CqutAiFxlS
xT4SSRd52E56rUn1esk4WvJ8czBhCwWf8UPmuDBTd66/yh0QSuiFiy8jm4xiygnK
DD5mBxkL3WGs9/qibqCNkVTPurSatObybLe5vImEgjfzMl8G1XIZe9JryICX6RrK
7YPQq6hStgtsW1SOExnq4w==
`protect END_PROTECTED
