`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjsD86XUr+ue5iKhFGZANmNAs9ERp3ZT47PjMxjE4brB12HsMI1ezX2+2EYs7cAN
9jJ0PsjKITuuNgoKMt0h9y07gahuuvcVDAYPnafrEoMI8KUwFhrxHms1jBdzbkxD
oVcj3oVyfGo6JuNLnx301FHWRhrSGKJ89kSG4dcZNuqhQ3fIF6k8yEb8BO1tPQa6
05dmKeQMiNwipzKCTWlyxg7gpgz+6LzuE98KW9YzEtS0olaf4Rn4bRDhQz+u3mK1
lM1ay3LFVkZN1jqhGQdUn3GsCRk7K5n7YL/XxAkzwhyoB289txSeMfbr1u2aW3oA
khDO8qBSY/F/af2I6l7T0SsqvzA9IUcf/Xs0mSiGlasrVdu4F663BSBxvLhvkTvK
C++ODz2nswfGC6mDjJbUM4ERFFtJ1A33VtozVZmAPaRbAaBu/TwwKCJ8uyB05NkH
KH90ljKUnd4Tg4inrQqNnunPFDvvyf8xre8okR0D+RBcQju1LY5P863vSX8vQ70k
P4NGY7pkf0n0oLdW1d7BYIcxdMJORmuPlIo95+GFepmrasnvE/I16zOn4MiwNrFg
xX2ifQK/rTtFGi7RTt+ywK10ewpPOBe4BkW3ycNjYcKp8YJRVZrrrChUxQM2CWti
PV3ffhfAuWDQFZBgWGSHZQxNuSi5kNi/kqhy+S6QyolXL/QOYfc6jeMorLxuWeYU
/JQq4P7TRGIb8DXvnU4jfS9OWw31DbV+nMMk9LHbFLJ+uDLJNKO4Z5v1ThTnmzOB
UIf19yJ5GIJdEXw7ePb3ku/6nwJ0IGytCsz1WMxv6zr8lhvO6UJmnfmCc1lWMyS/
t8SoUNfvOQWfnQTGcfNvZkzTJ8VY2pnMEYK0WDf5du1UbV216+ZwltNBBqF/wxuy
vUivNsMtUY7Q8GNF3t9t/BdW4Xu9lxZrwG9EFZ9dklD8tVzSCRlajtEGJrtEnvOR
0AiFWmiEc9tHHaGlhqVZxDjWcLzSxj5OMkaok6B80viPyF+yNsAIe6LkGUnrkDKK
OTo4ZGOHm7V3bXDQrO2RKb8nY8eGY4QFZsHCXCdQ3CWHm96xNyEp5hj555tffpMf
/FD87VdfxGuUqlS7liGggOnLiQbFygElNuYihrdcrwyR1gs6if8FedwdrDDxxPlc
0uaAVkoD070kctslYGdRj7qZRBRrcPkj0kv52XtaxYGEdynvCLFtoogegKsPnxtD
LPwyIp1AIEvVdXhyE9v80IyP8Hma5ZT+CrNl//vyFEF7QryVut6UMnhDAV8SaXQU
sg3GoHXd7UtvHzHKVTSOoDFCJj7urL4bORpYmd13NdGj9K5CAp8JR9qfLIhY5+qZ
cp3zSGbvqyJ9LgRXd3PUqf06LgyK3KjwkeQGx2NqIGJm9DwiPDT6MEnqlBPue3wA
Wo7C+B9i1zieP+FJv2B6QiiOoUNbebd2UDCFuNov8OY5tECgaP+Avfz5DecBHTm9
1l7I8mas+540VQk9U5vySlwh4dU1gov9j5qEXXJIXLqMw9o02UBlx6nMa8AjoTLb
SMNFlKJpvhs9YSKenT0Km8xQjx8sXMzhANWghScW+fDPv9wEeVP2GeW1XTu1jpIP
bHS+Hoj+VLvBawPvAuRaXHZk0soCaCffl5s0JFLzBUvproLrGfCUPV758VouafCP
BmfFaRrJcZ3aCuSIJObg2WJhzCwH0LMzMth+sFbWYL1c9inNuzf5XOcPhBcYugu5
SGFiYymXJrRbZypLhO8ISpjbUyGnEQgWOBSr8yMp+YWNEiA2XUbw2JDMaCjVZZM+
i+s3VYswDy3CvYbfLke/qJ63XFHsdXAYgKLZb6WzKl3ATACMxLCL9/oz7WEC9E5T
rLT8O/vmyfA+imC0xFyrSvVsvyBcif/J2+Ju8mZUDBOEey8/7GPy4Od3MzvZEukv
jW/yGea9auO7vGep9fPrhRkbE11fmavdGLFDviewv2T+n+2dXgaoTUA5vSuumCp6
9gJukYyAvPAduMVFrT8Ijn2v0SmpByb65Ty0B5iydA0BKY+JC/0Z/Q3B1Qg+Cr7e
e9HqvLfoB5ot18Se2JNRv4nxKJzbKJQLj56IujRuY/eVDI4m+9J7ZxyhchgAwrcO
5Fs9qECwJdIAyGD8Q44uQ2woE8hlEgbf7bqIip95vJS2GrEX9agq8r30BfxdSuXQ
Mwtz0BOIK1sxYOlw55RFIJ3NvVqX/wXpX1CZBbF/GZK2yLb1AUDuvhSty1WFvcip
OoLnD0axHPEhjp9GVFU5sqzffTOTM6G38skYrYgW4AVrmCLcC4h+asUX0xf4VZiQ
p18M21+l3LseXnvbYMbF+1Nw4M+XDRv4s7QquDx5A+fnjEBBXG5QhwOxdzazDbBT
aEHxWaYvSp4S34eI2QIZIjw1e654Sktsxv7F5po9NBfDsDsiWxBGfRho21UmUFvk
OAaUES3Pa00EHV1XyyEWMzhCTlXEDAPJGOVjyDbwwrPRPnY6x+qe5NylwBCmOP6G
UcAezfK1/mA9C8PuNT67x3L1vLuxPdOpbE0sKxHivfqwn0fl7P3Ov56JM0WlHzi/
+9nlD7PJOB7XnhPHvN8Dzsjh7G5KlY+vf8H6L/NkUrGcQNcdxt0roTiIxn5l53AU
2rOjNCpOszFASRKp7KfiKZm5C5u07fU+WEFb4eLc4GozqUjpdPLh+nMfZkbySPVg
QFkjRUc3WGKiEgvvgPCbOia9h/dKc7q0mpvx1+l9i8w/bIBWjw1f3rociQDdoBAH
8KbTUZ/xw/6Ow2CW0Px5JJa6kSlNdWiVU2jC+WjFgogT2DlNeOIftsYX0Kvn0Djg
qE/YUCOVpW1dnHniSVdbwXdm7gpVFOdcATRNU508xQukkUH5jvFIswsFO65GL10Q
wS4S0sQMq/aFjpAamny7ypQsqt+ha7ynJ5m7HIn/f24tm0hBOHi8obXoYg+01ynL
9f+KM/63VTdWd25p20DTAQHDaF9nxVHPuEYHGIqO/qyP5fBo2c7Qp1rreY+yfTZ5
JJiG2yz3Y+4UWMpfoUtMrQ==
`protect END_PROTECTED
