`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmMdt/S6wBfIclpy27EK94osrLxcV9dPkoG914jIeMJn+KM56iAKEanBlV/H9jGd
jHGf8x5TRgNrsqiOyKMBWmJrC/+WZExkZsGtEU7oEx5WN754KcD5SIdtlWh04gCQ
zv47nf8zK/JCoKmVvQDzO8Lpz5BMCmL9phzhTP/sNBL4kD31eyHVVj+lhn0+KyJS
DeobFxoXEEYLJiBEoOzI7VMzi+Fi5v94pCoNqnBZfZqZVh7qhVS8KGhTq7mjLjfs
bwNfm+0f7Eo44r5Nkfw/RBoyuqpMFSxTmLzl2CXnAgzTLxJEvtFSyaj/WxOxMxHq
Rie2NgojGjDleuxPzoXBxwuyp1r7jClCGoJQJWOYnMnjmwZZD44eGs5gbVCCQQnT
poF7Joz6hMTxvR+9IEtArWpAL0+A0dWZ6zAqlZs0p6HzcST50bddeWUscvZzL6Xz
cMoLbQ2gPcHbegHOZ2pkA3Q0MLqaLy6J+Gj5vgUwmxsYpAo9ZNSjsgJHOkfl2r/H
eiNRW34iMRbPAyt6sOtMH3nS+qWLn9KzIn8rmZHFPXS8uSoy1PBAF59m+O/hDOdB
m78QnbUiDpeXcYXBk06VpJ0sGsQBl8WFJB3SB9tYEeNjV5lZ0Yxr1FB0mp2i44O/
rzKvkQYTmjkK5rmvhsed5Ir/Y+kVzb+wmwgLsy+lp5Du5c7dvoyt20WZ08aFNBQM
5T8oj5xWuIvZUdqf0SusLCgy9DRP7pCX7bwg0qst7oJfs3kPtDtGnRkmdyb9D1Bt
`protect END_PROTECTED
