`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QuccJIyUDZ8iMCMaDsqoh/VgXAqzZucaQhUM8znUZ1hvO/scXHKc/1eiNQnTAGY3
Uedy01UMWoP/PRnjQefyY61VZ9WP3iDdKU1TQnoaUZ3SN2q/lOxdb9u/kCtBP9rz
+tZX3HerNi6kLpghJ/Ua6l5H8Gdmvw8CGJdnNU45TRmOIYST7IVEy6zEmaVUsLQq
4omgVmLxMC+8uxK7flgKUfptDKht0jmXFRFIo7sZv79y4OxJvigtT1dCH4DyLv9B
x8u1BtBoeT1mp0ZcM4BZXbQdz7iXfTM3PUfi65c2iKj1YLbL9EVP1/WLj4yktZI/
VHiWc2ceC11m4SQBNwfLy3A7K7gALUiGgWGYL5wdcjunaMy0Kgk7AI+0ePubbFom
5MnPkMCtE8W8stXET1L39y5nyOKysznPdnQQxREEgFOoTfqffReVOdpyFd9272hS
+kl9IvJ5Kc/AVhHiVC3DCS6B2qW8FXnFX3GmpKWzy+TuddwPD8msZW52TK6MZf3D
VupfMyDVCDKyu2Saddkhbl9xJg7TeRGHt+x1OMgn0MM+Jy3mlvzB9oxtoxjDxf/w
4qsp7koqcSMNI6QHgibK+XmcFDsHulIhtqX4EMHrqgpvy/j6KB2OcXKPROD93zAz
/EZrVomHBsR6xuER2Vuth8EErXIwsoqeojea444V1Ox67ycPt/nqYJ1dWR4GNI+1
oqKMElR8YKFrI8YrQJXZYK4bfvAFhDdLWStr2tgV7IVqMbzAwkr7abbdoRbIBb5X
PZVlmoMsqWu5SXSdsmNTbcIS5iqADSTNEqMGZZyt1Jp4gl/myvcO6um8+lB6xN6Z
9AGJ73hbo//Byzfru3EKRURnfJGhjPylyfJnHIcmPQGj7dX7jLNdYfK4LLQ3q9Gz
btX2jqMq0j66mfLKbhGtgGWJmfe4NZyB7phLMXQcC6Pp/H16aAibF6IM2Qsoi3mi
DNOs6mMnptvKeiF1PxeWD9L/WqliXem0teGFmv2/jlc7MoumXjNdfN3GxD1Ay+Vd
ZZ+ddnR4uc7yYYri3oq+f3EXqBpy8hg05CYCX4jfzTmAl1ExlshNJbAX4d3FFsKg
xcXbL4xsB65m6p3SLyuGnEbw8j7HYSoPr2oDmzj36dzBmsWHmYMa+gUN0+r9v6kE
Ug0K7vWmCmzJ5cn50aSIJYXAauI1LpgDOAqGrmerO5gMnlTlzZCLFNZ9fExTK25c
0VjhsXX5108bnz7XuPQuZwFIdiBttV4cJakOcUWFuxHVjoCYd6IDc6Nd3apwAWeP
Ej+SNeM0y7iM2C2IBmV4VHxhFW2dnv+P79a5rhNJEDhmW1z8iMR8HppjJ+aZD/Ks
bf741qzaHJrNyr8AeAlxxJ79HUxJ/blc2GfSV93DQJ05s/pI1EWJVqGv48FvOEGR
I6H0JgEBTxlMACaMvr207j7gRqQ9fxScaiM+iR+nJPsMLSILcPrjCFTjgm9LsMNz
9BDxHiCtOBcehcfYWIMGXjTizAnrRjOWPuiZaaaqKzVAdUN2dNLny2TsFUKbVrmv
20GMHHT61hyEnhzzvSU97HGpakBCQYb6BPfXgs1636bBTZ25Pa9w8raUt63idDtH
AYjsCsgA1eoNses24Tz71DMVvyymIA/WnRMxZrRxekKqA/YeYvjbz0D785fRx6t1
mMeNwr2K8RhUJMhxaQEIM7MB5lKaXgDjsVyKtBQETqR2NdeMeBpfmS+1qZmt4rjq
7sQf4x+VwWgnzdEr2uxhq98ikqDU61bbRoxGDEo0VxTyHgShpzbYTg6FqpRo1Hl7
LpyPrEvx8Vn0gwCX7OswYFUgatPHdN5n60lRXq4J3IZrUGCk2atqt2jdF4J1F/0o
9SPqUHBvBPG6HNuCOorjxoaddpX1AeML7eCYe/o5AKPXxW01F25yWnO1RllTsYG8
r7fwSPJ+OF5OtvzCO9uYnYXrxP0+vw1ZEEW38D/yCkr13dhlAr2706vIzKAnIS5a
5lOhA0DQ9brS2Jzu2A0aYmQ7B84hfyARXCkGhspcyvJLmqP/g3+P3Kzea7i01UOQ
t/3kJ3Ahh4zWoRRSQ1SCyt8Grtg/00QH6gr+XwTJ+uc2WXo2vrjAdmfpLH0WIewi
yVZv5+ubhmyphbRJiTEzpS8GFs8NFyrr88Uwk9XjX4+BoJmiEeumcLVvWlu2pGqg
W9dfvQknOHhSq0XjKoXHvm+9rDDGbaWeStXLJJ4jPku3BE4kPmA2ExJxzGnrPLOy
0EKJS+VGEQpBFbJ0L5z6WnAqsl2AjabAIlA7ePfYuKPjWCwELnPPugmW2Sb1LWZr
eSDbpQTu9nr54Ae5ITE2hrq3OdCYhGzTs8QndCngDv+ZUTgKfChH2kcxkn8mXWbQ
SbTKBZNKn9gyCWyR1X12EhIqGy5NsAmykqSI98fGhAwYYMG/40RWP6xH7SDkFwQP
OAu8cLdM3wr8x+7eIDB0FgaZ4y1nJEzkEzEx5qvPbnXkzQf7HX5JWomuNHnEuh8U
raYOllWMq0a/TUl9dFHgeZIoTCbUJh+DBKyAoWy7DkRO0cO8yDDtLnlfa7JcAH1L
wZZGAdW8Jn4BoP4/huZtJP6dcwEQqOgy5xozjkUSueJ51kB9vK2arzT2b0R7Wn7a
9E+lSpx81Ap3+r/wzPsOdIkarYQPkSxgVEHruj6lv2oi8j24O3Ub9hxnlfn2A5rR
HnCQRlLAIDc3+FxG+8CqsQyXcvxi/wZhiq36JLJPZ8YjxOnjkH1N67UUMUBcLEq3
/1JzfVkXDzo18G88YLcSnL/PD+MSoTP1AgulNYVoNwxtElslradf2JV25XxbKJfB
W+W7QkcY7YdclgJLbfM2SUsf/mNg8vrph3ndbk9telJ0scYNCAkj/aeI+wcaW56/
IL7zcsImRqPhZki0HIp+OCOnuJlk8g9T0VRzVPckAWonvEnsJ9K5IVPprg/6kAKs
vJOa7skIGe+7bhmQVxXwgHKsmFOHCAEpxaAWgfdf3ZzDGoFFKLvDVvyiQNVsg0n/
TX8D5o1ScRWdesetzyH+ksbSjKhgY97cni2FLNwqmIxxUPykhPUy2r2AG8SBJmxF
IJH+QaFonatvLGkVVrDXm6HAgtaLFrg5B35ifckeomPXMiIen1CXwlNQfFhCd17t
F9hAK0RJ4UDRzxmOps/O8mlI6jx532RFhM23v5x1slZOsbKsbUwV0afRNx7xtDCr
SQi+uO8nE9LHcnSxBp0uNQTggBMyudGXdB0U4X3/Fd8RmxdaZWPeglsBpAwILj66
6wV+gOoui8xL/rBMcrgufh7ZkqBnRS61TMBrq8vQSpHyw2xFJhtgRJlCZcub3DXg
m8/oLGOgsKw/memW6GrqXwLGbUWJ8YLgLmdxGFLnOzvPcVAV12A09/o2rtJZUenU
IiJESIt5Fp+iZovCsVTKlqdS1iTDeJ4z2Y30/ZKKZLwDsn8xuwGd65U06e+F56lU
Zsx9pak9/sJ7lhZuLp/p9eJPf/3uWDsjk6jOYMzQmoelv8ic67fHIKFuEKiYAFNB
jO0ElWO9Q9GXg4ZWPpxZncQvzNwEQp2jwWRr230RbuITsnG+WCRi0UxCVgOG7IZU
9Y0nXWXeJkieKy9PtVTUS2sx4kg32BXfrfW8Spvdmq/jVuEcwwnZ6l0twTsib1Fb
5jVBjjmIugEs4mkm/kVLJ+l3z3YXUIcZJOlS0B+dgMRRwkG4Ijbnu9loC1jhxm0W
9/NTxmQPdLum/r1WUeJdXJyfsWp0WHEpD/iW4ef14uaqFVazAkMGax8lZPDI1jGx
BsVMKPMNnpINk3BqEhqe+ZB93x1yFngyLFgdS+LawxYKQ7fkUMX1prFPkYlW2DM2
EY8pVug6u2D/X7Wm2NqsST4KQEBcBStrzJnZRS2svSfp6TExrBBcd+/NhOxNAb63
tzLfAOWvtMh5sCUusO+sncTzjLaSSJedUaUFlixrTfQ3Z8aOMBOjHqHylWsZo2Vl
MEh0rIbel8lCp/wHc/C0slM2GgNDnkHJaaBJbkRd/89q5pmHXRCzvabFs5cK/8lB
wx38L1mseJuMAlACnrYIsks21Gyb4ylB+htXhW4DFjksbXw1AyALddOpBYIRuAGP
J4IbP+L7SlssqWPnqEw+gQorTt93p0sLjN+MQbSrgB+fLL1OmWSt7AyFhzMB+ek4
d80dPoWazSvKc23wgIscAJU9YwJz1FrAa4tzG+IR+Q8JcVbA2JxypEodWACiaXfx
X8t68oswQEQneQpiEWQW2Z33D14+WoiARE6QaUccgV8R1zc66Bp2PSOyj2JjZWpW
C3y3jqIhJkFFCo8JQKCibUJv5vsxAE2xriLiJrHk1ORC0RifZD+ce5UKUqc/kEJT
pPBAsOKlKbDv8TA8/5R0VIi5L3tpfeZnmwSeOgzaeWdJy9YXSpZkQt8IvHlqQaFi
PK5YqTmKXtc7Qwc5G4dyd861WBsTV7lhxWWyi33qq6Kaf1JgbfCxDq4P8HmI4Nc6
XUgda47lxZfRhmli9jaUQCfh2TEeU3DuQA6hkPuid5DHvsQVw0SDn5qcFo8bjrZr
auujdZ5rZWF8RlwWDsbKxe6Zi8/lJyL43Iiu3nMY49EZlIQYhDhV+8d9yjNNBa72
ylZCUE02vKD3g4PiUKKe/lJcFE9/spPrnzB8UaUPvJ8BHqemD8dUTv7C4rL9Io9V
9900/WTjPmoyUgwlBeLeR+iJjTsJcALU1hySgzK8SSTGUbSHiMeVhn0xEHWlygXF
tOlLaTzFOnnnHCKMM0ovz+2U5j1zCchzeM198If3yIlUIkwSJiNEX+JaiB3TqnmW
AG9mgxNHtuE77l/cpWa+ygd0WiYR7a/FiGshafVIJLptvuVbG9h+1vK3Y24/1FoN
BBF5s2/p4JnoXjo1Rl81WzEotQGiwDWxjsWzFR1MzbV5BKqwuekDB7K6wA2wCumA
XMq7JY84tEvy5Qht/V8zxYOL/ycMKtoToCxn+FY8ptn/eNzvW3bIzwnBdeQqpoSU
Eve364JygDoHETcQZ/yTEmSKzG9xyvJB8CDzbaRQdWCzSdWzMXbVBSpBghysNsFJ
tG7/kCQVyoWZgbzo6qvALI5L8X3BoKw2utw5jm+z7YCcICqWk17fGCnPoA4wxQk7
MtoVUJwy9tLW3CdNqaum2NmLH3pTEKsX6eEAQFbM/WETzUY4YCRRA9L/VSZeT3B+
EgSknv2ENe3CL+ObG+B3UaLMOHeO5PV2xcm1zPby0NU+WXlxQvsO8SAanJAzXjb1
b3J5XhN8k1M+WNo+D8O9k9Re/S3d/0GDeDETvxAQr91Wvu98S1/khHSz4806V10R
rpsfBQQeIT6w1IEZZydTQefH+OPvs7HHAObw486CRnHkE0Pkx2ZIf0mn2NlrT6L4
o5w8/bHT9pORiKJtyYT444kAM+XJCVs49iONVBQWa5BCKXQDY/2hh6VzegQFAOqz
g7P9Cs0tVRqiHJNC4XsuktbN8pLx34lweZPTeSnEsmhHux9p7Fx615tzJpBqTp9c
/r8/PwUKaJQq3A2DUOqSJUSrVxe3eotCut/kF+3sy062MPjlunTSO00TvWjhOXyQ
nKNJ5gCC/72ac7T9u0KyDELySDBkljvmHtvaDpiA1XeSgg3vuMuOVOrKkOqwJIVE
+wj317OF5OENkc63D8470YJECei8mqHKPiXPuF6SCm8ZAa8tBjHI2fjnPZL1hO0P
bdDOO13MRj2TdU8vH7HJ3E2vfJtTnFKlwaJHHCIvrujbbTeIIsNhbGNwciyZn8C8
1Tov1DZ1OlvXENGAttqJGElutDe+kTsOByq+SmPH+mdSDXy9fWFh5dZh46wSDu/K
uShCXeGZOBO9vvain8751S+8xPZbHbdfwMLwhv1X2LBvDQ67w5iISVX0vtGqIE/d
HiDmUgTwCtPHHG+vhhHMge+duDQUxjw6BgHnrF/ji62ZcTOAYn8tftJlySUkfGRU
ESrYhE96qamckS6LEBJ5HRQ0FXkjKGSrqyxUprGdiOpHbUrlWL3rMJgdYTWlaktr
EXndb5J+GNUiaYfpG7zd/XWxBsUNiwdYq1Yo1CfEb+a1VBo2qOTm1FEVN4hCulV0
Bi/i2W9pEVFtrqAqp5r7xmGXW+1l17fZxVbuigyrJmmOSMVLlXirgN7N1Kun5XoF
Ggy+Fsz8Ux8doiEQcER67Q8sW1SGoRJ6z2VRncbfqt1hDF2pN6pOsMeFggtZuI5R
+P5dgNlb1+J4FeWUOGYET+ndtGd3QJ/PNPhyBuTDaDmYOW0QRDymgJM/QWZsX0QT
vSe7iNE3IidF9dFO9N6lI4WJq5r1lJJ7QK4zJ4eKlhklA2Fp88JtTFsNCByP8A5k
O/CUZ77g6mZQPd5CFh+TjLZSIL1BRrKgm3t/IWPaA03+ICcKRyZ8im5m/O2KuRib
+fYT6lzOk0yudtx1TUMIL9PFUKubsFRuHISksf3m+bL559Y+9LLYaXpLE3Gz3nb8
0XEvG93Q1hhSr5PsWSGQJGJ3oylokerkEXTDGwkqj/LnP0OA5LCn7FiClBq4GWSC
yfASADelu96d03pkRdQDPV3xm3uVxnXAE8wOEdQ7qMIteOu/mE2+N6qF1vxZg4kH
ylsopbhXv3Yxtpao2R3jlkUpNCZ9LhQKFya2CZA+7npqkEdXTC0i9gbYDGvDpuMI
J7YJj3pQ1q0Bk0j6F6GA0IwwdwlJbXYIbvmiUSxR92NLrYarU/ay0lHGanEQ1+io
uDWF5gGJ20MiS9yfHtDA8SadGMBYjajwEPz1PxkNVVtytcz6L1GHqgK6AQqyV004
ny8qs8jgYqhwca9TnffuvQfVSqv9V1VY82zudJEmxXpRp71Q5TxwJFZZ03i7J21j
vFqXa5I5LtxfOdeuzEzsJmU/K0I7sffHIy0/n5kksiwMQ+0c8TrM2Bwiqtt047xA
XZw4G+JVtJ+YBecrF+1rlRzz7ukNiF1BuD6RX2WEKKu1pFYSw9meqey3i5LdA5rE
YkDg1Xc3PgIWCsOU+NFJ7sZTQVNXFWM/aw5wtWzIZdvdey6PVcRiS7bd5TR6D2Vq
J34iaFwlaunM9+xLnPNpGlRCweiKdLFPfLsfH3KcImOmm63KRL6gU4QiXzoAvcU6
yDFF6TBgrS/lH3OX6e+Ovi5lKvjGyyIHm+leR11WwOCDQpY2NwN7dYtFk8pL6+f2
/Au2epM1vE3MkCMVWCkHJgCBbAgwHuI+NOYD7lyijjadTnNGMWujWEOtLWN65hIO
5m5z9GX9+SjsFf5xfmLKp3dZqUA55FAAk4e6Yzs+ijpHVP4a4dxOD7pNl783GYaP
S+Da1OhLGGU/gXDmEp7Z/nu4XtGOjMiW9wHCTjD/gblcE9g+J/UErRqUoWo+MYUx
867cidgDaL11WeFWbNDo50CH7yIrgRsxnlgo/ixEysuSeF8veOO9bIGyBgmwp5tL
no8yrdjc5Cktwx+9vm29aTwjEIXtCCzBLdLWTJn3+FIqjbrnkmfscA+6l9P1CH+A
TG/oDY1kyewYVUyGLbRoTmcyNBOMhYcpw8aCYd39xCM+LcztEt6l52RJSy25D1nd
B+U4T2m7jcrLqVB22SmPyLvfsgCcE/eqwPhh33IWpBtNn6fa5n0pyYU4HG8J8TSI
fbZl1n7wLqV1kr/QAWjhrC0X2PD52pO2jXzM9DOVtOmoad7vweYpV5ICjK7suW6z
uBSxgoktSmJVpFIw2Pg8YjcPf0NUHX02Dhf0jnqrQfvvJxi58NjtgIshGfWkms+T
iJgyQa5FFUGBTw/fqUEtSn4nfMiNy3saub4KAxeSG7gr+MPnYEg/704L4nX2Ux6a
UXbh8AKn8dB6HvMjFvA2zAcUzTrrFAQBEYaRKG2quNN3SPKFH/5Hjpn4lLiynkt7
LEQh7alLYtlOqpjhQ/N8/R5iInmkFfQFnTTXS3zbBK8vRw/Alr48Sh2d2pIAg79C
FayMWHdqWfebRwQh3W5VYk4ME4UQ2Zc9EExFw42b6pMAkhH85+MYmB16V+eqCmju
GbAosODx1CS2cwBxIUe3oO6rEOt9nJ4tGOg6iTLgc5K8mzq2XEG8ddUFdIq4mWOL
tUoa3el4ogmTyROe0smYyx3y9NKah9BoGL5ON9CvR3Peo+kU1/e5ARRkb2ZuNWyu
F7aj7tcy/9jwQnXpzXhM3KUDnziOHmxeshh8vmU1nEvN4UCmR203c7hUBDQs6OKx
OJHSrUdDrPBB0NYzkp+vJIrAvk0oxYFHNPPeDqL6AToAU/vwZaS8yy200zOYdEtR
VK0a1ED8I65i73ImEtF9LBoFbH0VDvyNETInFPHfbbKJTzUO4PL7udamw93yWZD/
i4BW7evHe/aLIfPB+mVmJ6dupEzrEHw9zosslnk9aK4RXwHbV3FT9KdiVHEhDHiU
L8Knz0kuV3/OjC0xEsDTbqqleVvy4rPhSeQkphBA+OIUJ8vXzKevnn1JeGLkaKBo
px1S+inoVc+iliTaruIHogjFxgpoZ8ikRwusudEhBHCe1MEyAF4yV4Bpvo1KnF6q
egjD/bXGpWE/84jM2vD8CZaLaMATSnTouMGtx+acz0sPOn2VjRR7nrNq3xxIQLYX
S31uSKKsvuZ+HZ0TyrBYw8S79Bcx+h6aXrk+B6zb0lJLTZbuUn9JpHxFeEEtaJb3
wrCeVF68uT4vDfu3Hq8Pa/n1AusWQl2GO9+0HgcA/v91yi911I2v045YxzNlX0zW
PBLX+nhCY3qgNiJFH6kNuw16N2RvOZuJhQAalcp9H99XmCQLSUQZ1zuOEgmlr6tk
LiWNOuY9U7rblWo/DKwDj1JYSYr7hbJNt7TvhPpMoWOLTz8RVZtUhpNO4BPkv2ST
xASzbmyEfS005hRmiAtbSa7a+j9IFk2vdL2m9q2Fs2OiH4wcZXrC1qrvA5XwkDiw
q6fTVXQY3pLsNwNOCgquON44LGHO5lRB6UaS5j6H5afvySrUs1xk1HdoxJWrbXyv
s90HVNYFsrDEOfK1dGPaJsW3Yo0x8aNdfnCXh8lk70b3xpvVzraW2Tzu0QeqIxUD
QYVYmkw0MDsXwgi7ynFstCtDsmDV+Sxdn/QQO2d7ghmZxpSWKNJalxg6X5GQshQi
k5pXKMAG1MaibLyzTbG8Df3gjjgID+j1lkNOrHkc959scL3BADu8pSObPuYSVF3F
U55iR/sEx0qI8gPIDJ4AAiots72VoXpd/YpCJGSq5aArIAOKLdOSLuPzta9v853Q
BKqa1bIEL33LOWuU674uU1uq+kHA+MSoCr8+HbNlygxNRCbWNkvbXqQsYzRAqDKx
oGbWUacItNBVSq1fBXG0IDq+a10Wj8ox1msk4yNSb55qOYoxu/3V6xLmszuJmV6l
VHd6Xm46j1Sj7l+YK8VVB+OGJxNJ1dw885qEUx2YkmWFw4b/aDS3w4RgBuF5JxwX
OvXRFR583OPr5HuQ6u0JUODO1ewwvEzx4aHHKUZD1UnxIcDGnvhTf4/sCo5jBKEZ
tvJ1BmpmKwxOwtiSX9Is5313GYb2Vu8Gms3r/Bh3hzcpebD/W37s66FZdFG58w2P
YPEjfirjSKtaZf+u3TvUwIkc6txhxP8cm8D9nFsVHbo6Di9e/eNNPbyLmOnpEEF6
WaeBScLQaXOO683IHdLJ/wGc0MQYdf9pnbz0NNVJo5ynyOKfBqdM41Gc++9BUHk1
8LdussPcy8MWHU5mjH36ErdHjW8ht59KQgtUoi8tqwNWlZn421q00O9xGPgiaV+b
HGZRsYkt0FigL+zcrfMVwZOEeuM0EVu3O9XwtMOSEeWX46Vi9x+M4x7e+7PuKKap
daGsYSQsyhNQu/EoGQ/GnhiKQsp8wpdz72mlyZN/3S0/3Ye1TVF7j1Fb7l3sQyz7
qSCs3WGUx9iyRcgtqXMOgCdPSll+qS+UfVbtwNbiBA5aTd154kNbP9JIa3OqprWO
5v0Q7sHO+GdLTyFsrwKvGxImPj2E7c3bkNRA4xHn7vFUwnCAtgxMEsVWVgmF9LMZ
rlD791ekHEtM0CB8oqfJvIe0wfUboIsH9pK5VklqHZYLvPVPr7+tO9rtcUpak41D
c9N2CUPDwTvhV6YHM8od+NBt7u6lFlHwCbhtH85cFHcRhwGI6yeQ3lhaineOvbe+
3t4GHeJIezyL0vWHhkO7K44CmwxkbQ85gnCDpu5IQmzqZtVbn2ur1FbjmH/g/eCn
J5rdNnAvy3GCZVG/xOb6M9+bMHXhEacI1rzQ4g4OprDHPjJNVaiWvrE2djjeseu+
iNO277fu1VH4kG8LFJ2GLCXA7oelTYDyzmImfI7xVZguk54YTK0fIP2n0rffihRf
ed5lRkr0mJk7lWVBMzI+0PQXiKVaXMpBYrDA2IeyRAfICVVJhHMn3392NbrpwbTS
xrfF/AwVdkdXQYAv+ValPgheWOGx6XTjktmpzre0qqNv7hsF5fxfqgkGLH/U92sv
4bADQl0Ecmtcy9zY2BB/sjokafx8pxGdzScyG9GYEgCdwhG3mG11ZUVxX3XEvy7C
L2p8xAhyqzq1ty640ShoMk3ASncxAJDGCQY6o1CHTHGcWYe0KYam9AbdimL/CHsj
Z4wWoVWWTUxNgI6ruGPkmEL6I4IhJX0+05Vk15p1eooOtjbPErARXKAfXazVmMsU
ogFct9YQjKHtrQmQWbU16rsKXaAmg88Fq57XODImPl0KcvG0Oo49M3kefCBU94CQ
1S0W6YN9pAIvbs0TiEqTozGpPzwLj93MYbaQfSqQksPrsH4xf0NP9aQ2cnlwbbZt
bjsKpUVstW1njQMOBJy7cWyf7kiuiZHow+cb3nQwHdLKVdsEcmEJQj/BJMQk16+a
tp2/MgeM7mPXa3Vi20uhYXruYAbkVT5AA4MpvGtu7kZkLs0TlII6FBDpIRwPLkQl
hvqJyGYP698JqhlZZKeGRiDBP08+gUTaBLaE3X48xCJ5fcea1pTZXnQOEZUTnOew
`protect END_PROTECTED
