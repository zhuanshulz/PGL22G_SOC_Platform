`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MGFQAvxfRFymP8L1D1TlGhvMHdsWJk3vGGeNwyUdu6cZgFdtr0Klz5hxEEqcI0xW
KPnK4oLpNM3/8z2ikhbMVMCqAwFNJNjyHJbSavF/xltpvlwieKizoNhfpLH+K0g/
+T2pYCwJ+r2auGOg2VfCt8RvPdyrfDCFbY1SIQb9HJLqLBdaGhx7UoWrdcmQbOyp
hvFBvHhGCfnA4dYrZYH6shRONHR6o3TJmbdz8sgPR+fH2KmWyFsddGj8GQt1vKJx
hLbK2VCGAyNeSSlfbQs2MXNrqvdmb8fReUVyqmECJCZbITWEJHcaqz53CLGvOekq
UWlucasuGQVmYLq12Sd4N6xvv0FlnT9Wy/LNRhCjecGs/RshQS9m2PFQlSsbBhEx
U7UMkl+xpRSRy6+Ip6QvtaiHrE5S5bDOuY2+3QtfmoCDCu99uiTtd7QlZJvtyMSZ
tOPXpH2h0Uq08AQZHbvJSXsfYuZJTbWmeyl/rXcK6/j6qki2RVNlyxVRz56oJ0Dm
yvu1qViePeQ18MDB46F8JY4U3WwQWj5+l2pOyTjfIGAv2WCS6dg+mb+88STcZ54g
`protect END_PROTECTED
