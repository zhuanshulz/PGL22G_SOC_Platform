`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
36EwO+x79UpVAVGIvay72PgWKt4E3ZdvKA2Dsto1hqCl9PtA6SnrMuQmWiFlZa7R
dEMfHF4ruBZ+glqMqPfdNrOoAo3XVPc1f8lKvH6U5HGpu+pluNlkDA1v72edhc6w
LCPpL4FnBtQb6U4SVt+CszLNQKFoAJOgBdLqloJivOj07WwozhrYA0sNXIhfe5VV
iYWKmwEYWc+Hy2fHdf+xnhc/NilP1Ca0ad2E2m+xgfc+R4WEG19QwppIav29uRwy
+myvLiGTkx7Fr4GD0i/0Uo3TKfxuqG5ds7TBkyvKQpBv8BR1wZ8iN00MzgbYWoeA
IBnLsh/c0VwWrWsRzMZJmz4eRx3pvtWAbCZvO02zDolCbxF1/wCBo+uAjbd8mgPr
eP5EX1w5Sg47sJYwWqDoMyAgfER5v4e5eBol8o7YZauOMnoyzjQa81G8Lvo9Rx7D
DpcLcehxBFaT59R5lRlhIxP+cmb6myVOtG3Sa5/m0DUig6bq3hCu5H5lGHvjyI3b
iWB7vdYrteDKVxb1VcUIH2nE26h5XNvHhc5vCz22iqkVxueuepBZHf0LCsdfNxfG
VeyjFCSphvUnEYG8VJgb1mghyAYBMAJBWQ5omCuIffwt+4KQdIrQkUp7VeiUfAON
9VjcwmQPuYkhuPW9aXqVxDQ0qB19oMDOFU3klwa1FO7LLeviAfduidpnSfNoCeGB
8IpwC4x5Wzx59leobmDQyXb/4CKFMGKZVz2dSSM1wOxqSemh1XsC4aDO1sTc4zkp
Xfy1TEH0Q9FDMTuUg2LGv7su8o2+4pRxzmTxlisJnqgILu+r1ph9qJsDg+VPlFTc
laXWWRUTe+1iUP9pYC0ysk7iQdmzvj+XbbL4doahJtVmc6+Or67+m9RXQjvuO6k1
ZSfnF70SFJge0rz3LuFfgIq53lhMxFWnyOEiRFfH1OABgfVv67jR7XOKwrZbMAzI
NFZr54jNtGb9UacGDxMHOZvA4jhGQAxpGm+gGEQRRG4EvSQ9V8xhRNKrYG5ncqfP
1F3zLHlG7loV4VukSYzZ/kt+BF2OmHeaCzlSwLFN7b3L9/t7fyZ1m7s0Qojq+PF2
EKRkR339htobm9i0bBPJsi/0bak7YG2aafapvH65suLZDvRdLGj9ltqadD4rU/rH
/eqGlpKoIAxGmUJvV+L2SSf7sU7PzAPE3z9HHAd6oXJWSZkxKDDGHH8ZyGUbRLvy
scoEJC7im6NEhJJNryXK6p68f7dM2WaJiiG5YUNQjtLah8UU7lml7yWFEXkc4SBZ
zKD/b1B/dJwaMFCjnxmEyn/L6iaBb/xpA4nkLNs8+wI+VGnaypl/Lf7ZUG1oCPiK
diZuoljQCc4ycbhP4p6Bw264yNFkBdpOxFGMF7a+jbVBK7Di9RhidbbhI0lmpbVd
4EEayE4MUPq64pVDhtlP4/k/1wGciFWRKYqL2I4cNGe6jwOnyB/U80qmVmOobkv1
TnNDXsE1SleytEtwAw7SZoul6YDkjsWJpVrUSF6r1lqPOr+XNx+HJ0gFe6hPLxPR
nZNTktsR+pcfvDk+WrREI7S6mAC6QSYxd2z5p7iHb6oIYI4UG8kKghGT3AWpwDgK
sFlwZtyhZMeIUiEecskeFRqAFrtPaWBM0NvTXDAuf7M6auvo/7dgaEIBo1dO0ukP
9rwTtX6eIUC5JXC+ZrIXNl8Sh9N/i89euoay45W1SirHuTXJbPWDGQnVEgQaByq/
AyWTa01H1dm6NoGF4R7MzXqsbPwHqJJ3Kw12QpJ45IgKwFk+iM+kKmEXKUeY+Isq
ShL3rA8ZVuzjMOajN970PngpkO3izbkAMAd3CazOfmopSD3zWGXeFD8BT6hoU0lR
7Hu2eRlVAHmU110HHOYlFRy3ZbT1ag4f4FPCwY+fJ3S2UE9we+4uMUNvbalEs6f9
HadDrKAhwIG9R3/kPuvbCiy4I0SB1n5vePecweMvNcWAC/JrLNANXaF/gOVdbtrX
0RdSh5AP8ZdHDSQDBDYyDkIpddqMVVeJ7egmzsa+2dhca8nyqEMR+bIr1SdUaFUA
7EQXwzTYOBEXLdhfHtHdFGApROWO9MW3o4BX06dT+TRM7HYieVgsEQnAZt8Sgerh
EOLzQNKl/r51OEoKU2SaEPd+7EZuGnzRqa2JQwD8w5lIV7cLvGsjhrW+AJ6YVROT
hODYLTYefWamEUnIPcYb9GKCJTpiNnNcrdQ2cc/4tRfyYSsBLgAA9hm8KlDUJD9E
t3vnyah4YEU8OMOsczSFvovjgebmQvNVTryIdE0zjN9XJ9O8k2ILo1FOicrWYg4t
YiGJdjO80q1K+Xx1C2vIy53ZkWNKNKrA2gGPl3mmxMdxP0Bt5MargeNoC67pm+x5
uvwMr7yMQoRK8DUiVcDeFmF5oO6Al1Uu6DR9lyuUdm6Z42H/a35JOgCCkfrFfyc4
EKenS7jm8GunRAC3hKCFaFle1f6TFFBhKDVdntAUi1Pvhh2kmXhPv6jPRl1tjfac
8Ri74xyYgslrjYzoXgLdbhLVBg2hxhL3t1vfumkwlHbiUvBVjZ6gEFoxgDDiFWWr
js2gHWZaGcUP+h7gLyhQLIC72FkCHlww+e2edbY5zhFS/ZdTugrykaxB4wBs0io6
z7Sae8P6uZXFqXYi1wEJSpSuCWhqP9OaYJNdBsu3IXpgIty4Bi3enHJoQk0Zttqh
5AN0wddJNsUYjEDOYjJnBVkeaUg6XbZ+0nO3MM6ebrufYEgo5jvcACBLf2yU4sxa
uML0gyYHcTOz+I+W28ek8IXSJ7f/wYzF+MoGoIMFQrlcRBH2qnNFygzG2lluk6g1
NTk/yKImQIA9kcl6kMBj8RmBNb/b6dyoIKnPD3GCvs/CDVsYK4+IE3FIrxLds/xJ
JgXajXnTcWTa8KC6SUoPcXhKXod9r3fU+FWlBm5EcLBiU04dOsQYGiCIUNu+Tj2X
ReTxqJHfpOeSJ3xbLB6J88Huh96t2kCBAC7Z7sVHt6pNUwq30+sTCJYNfbv540fU
0bKV5AwdshF3nPnesvufhhMhTJTVq+tY7qui6jMkPbMfXGjtwzZMOGHQ2db4cif8
8yAujRkIF7tKOEgIwzAC6C4zbqKJA1IjaoSuvBB46Sus9bhHFjN0iBM10c1n/O/f
6lSeeqBimWuCw0M8ZW4WowFpvcZJY/W3eLsq6lGF4+lBpLMdfyuCfJLhp+ybFcy7
1sqhvMOjHj6rXmKbdGotFHTgq/I5Q4+4u2XqnbdH68QHy3MaIBULx4roQSHMDcEV
AG8L679okAOC5uQ30m3YwToO+LYsZrlRyDSJPulLlh0DTKQwdbp99BgVXmOz5SU8
OLeCtBxjKFYNBvZje+zRsN9LWBPwLDPNBoKfnebMa9rNOp8jEFFG/IRYcU2WM5Qa
2Pli5FUWAG1VJkCN0nmVCPaNym/GEG0mr0VhXwrZVuy1USIXa+qnZ9uuB2Nj3nfP
U1iDx2gG4n11iNowkH5XKinl8ftG8O8PBUzN6oV051ASGVWAsL9m6+fxyiFX0jXa
n6MmwRVOQbVpu05z/LlHGZYwbq9PaSWQ/+qEtiSpToHt7EON3zgbmK4aLhy36rCB
b9AYzUlrOvc5SSxkEhKfaje2vLTWb/rxGbqxJ92S5ni6wpkBCTdOxCvIAHrgPBML
YoPiduiu9QOZm8rvF79Zj/K/k8bpmL5oT+1Z+pdylB1ysC87VT4i8cBFflkkBm+g
EwOC3ay+Zmg3XZMR2yG9G9Yz8bKVtUPata3FU8GDNBfjUGHW7AirLkz/Qpg0McAm
dJSSOfz99C0KE7IcyHEl5QvZKLpun977a80770gFj4V5XFYj+xEJoufdTwG7LYPe
F4uwbqj/qIDViBF/63CDSkY/h5LbvmpY5tIi6pMWkQbs1+hzuDlwFt2IRY/EUITC
O9vHkB7cD0SVUdb8k291BLxtpyzpQn8e2VgJcqCTQl9W/uJe3Yi+D73GOOS1KNqE
X3ylXtEUfLo4dL5hhSf5LjsuFGoN6HLVEpEJzPKjeL0uLrG2bWpldGFZyD5ChNBZ
+SJozrMXjma62fUcz30ULvOZdxtGGA0Q5ZeSzM601BLr0pZp6W+a4E7KulWrveLq
KMr9kKNUF2dinWzdmNRtbX+Qhh+ADkLbRleI4G/l9eIWFqM/FkVkxEGFTUfi4ycd
H5VVwhNXxCz/MQsv8Kuq1Eh2ZFRNzesqU81AGLcDe5fYRy4rpGVR8H3LAhNnc1nd
UIPWIb1LeA9uPWZiYnQPpo12mcqRSf1QYr0uGtJJQ+fJ/ztqkOEAtouL6xePmrph
5i57x6Ima0HK4v+ISy5TvNizp3Eyi8GSs5rT+oz/1WbjR4Vh82YXQtjnvEFgNzCe
cglAoifju1fMrHODyPXV/l8zCGQPkdR+54vDVp/SXKqwr6d+mxRDwWBCUJwrUanF
DEPuQpFYqnNZf5sCiywRE7PZBNG+g8FcU2RQOpHTzjRbOmFrvvxJD0cnZolVHiNs
fKUE5xPak4SHQxdTDGBq6ic7ScvOJEcbl36ehKCGDjNsrRp+s+iBbYSSKpzgcvnS
iLQ7WBhwo8pZ2f+jfFOrGA8u3D0c3x7qcjQTlEZBIeHZCtTMm/A5VQt1IrmtGg/S
e6weBJpGrb7X/wphuHo1+bGCANZqzIOWbitVm8LKvBa7OECmY958QQDFl5rGb7Vh
xrYRq/g/6pyJ63GH0+wJiyx3o6J7UCHCpTrw6srl/JIdt4Eiej81AWD0O4REgxVc
gqEzXLOS4fgBaqndamJO/gdEn/MHxXiJre6fzgHCKuzO8JTb8iHJPSlruud7Zpk0
+dtlHEAZL8HIeDPw24oRoJZngABlOdE7U+qrjbRfl7f5786YybOQgpEF9MBW+MUo
8kPrfOtCcdSCNyw9bpU66nNCaQ37Cd1SQfJKIp9X2U28nnerc1M7zuVZb4uIaryG
eOTi2ig0TUu7P5OYy7Yr6ZKs/pTLT1xj+yFbVJhQJV4JpSOM7DsNI3MwCP71z0qS
QlNHFWYBuCgTSOZk+WQbX03Hvs3yW7hfxo+je3vom3mhP5JwhdC1C7ocqhR80y2V
bqCb4XraW72C+XdKJbiyylpGltzWGFq8jtOLPk/QgceodxFrmRvZHd4E+qVz1Jdw
FR5Jeo1HJd9Rd3zV9OfEGlK6qB4MNheFCJ6kz873xI7GRh2WgI4P02TADv+zuQ3W
nED1xCH6tD8MnR1QF1tS1NLeqPVwYYAnH8OdacLY3kEyMRW7aQJQf6qSPiG7rrRr
Y/GQqVgRGuxJb75YmvAXvbxBQcZopMENScW6wVSyAFUgGKXQ+i2UYaC9xP/vYxUf
ZKP81dlpzJa6eEq6v4l4uhe2U4O0KqIp6PrIOCXSv1wkbRehbVs9stNNjrrKdO9y
Vwa10EO7/9pGXm9vKwXKdxYa2pHFjtfz3LKg2OIT87EPS5DalN5nvMhE8hJcC8Jc
zGzCdDT+4enVT7/UI4HohGZNchR43/2AdlkH+4Cc7ouShe/WJ4RzwrDlE35zs74q
i/0RHqcDm55zU2l7SwbnoWCFInqKWR7xGaejWwv1MMTnd9wSknOGAw/JEdUMwdmg
1fpNQKOcMGHLSVHw6gV3RQ==
`protect END_PROTECTED
