`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNxHAC9zSwiEG/8lf4QWco0v2IK66nBDP5GL6Jc/T61CRNw5W6A64sbuuoTm1qoC
QxmouBZik9xV4KIPmK2g4TJee/uLEReOkz5FOAxtx8lHr/49KGRFvjDn/CH0IhOz
UJNVT12jL9TPXtDyHEbOxbw/ARfFWWPN0YLccci7R5jKQghaQFrv45FhqXZ/d1Oc
RdR07/8lrRax7WjbhpUYP36O/SresjPczGBkkcNEvRdwYhoPuI2n85HQzok0iPC/
IAqb9hUuh+TWJAJp5rlxsS6Km0/YPirbHG9d+StwpcnphLVnOwU1y+3AXsKkI/O4
0rYqzPCAV6YKDJcmuVIWKJHRrMOb7vq0cNgdYuMsRpiHKDR1u2Xsfl7FVXtd2mxu
zFYwlpe055n3RzMlAI5fkf1LXncK7AHK8+dygzIv0Ne4cq7yQLEEK4DdWo6DkSod
d+zikguwx+2456IZxuiIrKrtK6BYA7vYjbPcsmx02QAKTNb7Rw7CMh5ewYgiiYbB
Wwj8O0vRIK3+CinqbHrMy/Lna41QByxklPv9wjTRYNq079It+rJnflt1+5OxZjIx
TiRj37z4oBH3ZLKyxPGkFESl1Z71SXe+lu6bj1pJ5w4ljQgcrTXgC4WVH3bOQk6N
T3Rh9v/nrTqIqZS2gyO++tFjqa+Hjk4IOOBrbFrCzH79VXFoVUSvRRKxAdQeRVHp
p9qNUv4H8EBIkExsVP2Osi1dpGfzTTChXacf2f/NC10Xf98FYnkde+QQXLY7LZm8
H6SAuqYpNEtVunMJ8bENodWUCSXdXmm8rGfyXlcyAJT/6LKlO8fC9rQEpy4mDeGm
Y/mhlBJYonfD7a1NZd2QHpFOMk+lZekNbmHi6WwWMble+8rTrw333J/B9JZ8ncDq
QjqPK3Vfatl8P8WXJwu9hxJ4GQG4cy2PsgH5pA6G7gbClpdMQjpGYGKo6zidPjN1
2LufrFH8NPI8kvJ2JrR9gH9/E0UJup7HUEKfFZt9ozS3lSVTF3TNEZTfOB6iB+iZ
OzPAJraJXjaFQuJ9a8Syks79+dyTtFjF3uKLGDIX55QJCLEtM9fcCl+Qv+aLWvh4
Ll6+/owcPNNXrzfNrmaxPyS+xsPcGeuRCcQXuboA50imOkX9IBIib+VOqd0upZ1w
j8z6CxjNtuEbxIm0IYisLIL7xwp2HTOOwF9RFsax5Yt2BBaQGyQ0+dw/ivWUgf1Z
5wMmsO9YsyRHbzDvPg1JvwNtjCLkVOQqR7x+wImSX8VgL6cAqsGa9cWXEmWnq0gy
cBZX3DMo43NYlaHQC+OhY/oYt2dq/7dzVazLOleKdJUSXpKT1U/S6NE7HGJmo4pS
MjZ3qnlqRIWfgoq4BUx5MGAbF80wta0V5gzafbwFIzCjszOUyJ+7V+ltdATTmrCX
l+yYtClb3EnUBZBqbivXqeKl5Vocw2SQzWtRgMx6FMwb/KJw57D106iYD2YxEPO9
pfpJ2fAvrazzy6gQQHL0hFwc6MdHT3jKrrTZeWKS4M5ebcQ8/xIEBCgi8HOIJcUy
biA18SCDc2JufqaItdpRrIzJ08qMf++pHgyaZFc02iNR9itDQ42XceNF9coz+s+N
F2sO4JEWlaQeZFuh1Hxe3OSdOI+siLLQHj8yHLYSOBCO2+7KETScNG8REg1MB7ik
v61G78n7FuhhXjWlkPDTGwlsd3gPQ97Atme3Olvkd/WyJGoQQSNbKmyMPm2WVile
s5yC8G9NQtapiQrt25Lq7FkSgQxehqqxxZLJhOyjQ9aB3IyXhyNTYbD1QjhwNoNy
`protect END_PROTECTED
