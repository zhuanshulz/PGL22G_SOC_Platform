`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wC1rBmveHKalv++Gqt6deih+k/FCuau7dFfbDLT60NPNs3cj+lPMNkPbAMqb/43
p5nZO3kzeyTIOHHbOYeqjDGxcMoSSl3AOGIa4Sc+ElYOtWxPPC/PhePqJ0Iv5yux
S8HBiz0q3d+PbjvrUXqHNwoFO5NSZn4bzo6f/owNYCBXclqiOW3XKjaNp06jbK7B
HkSv+MhVq7xrePQUH7Q3g9yTS1YiRIJftT69vRmN07icZ1nAd+c0oi6mHzs+8HIN
y8xhS8i5T0ZX4qRrYR7c+6gXFpk61bQ8olTTD1uD1Xtvmq8EIjrRYhPPW1AZyIFM
caGp2df9sSv/eKg1llGsLjftc/47UQu+VVIST7DJ8EpsySEdsZbczAZmfgUVn9zi
ZwZHKuZZ1F76uK3R1I96o0ZOsJWoaoRZGBSZYrFXSSAIlO45xakcE7QqwpaeoBEo
bArObw2LRLpCowExDcnqEWyn4MfhU7cvh1TBBr4m0v3ad/Y0TgcdXx9TiEHjXBBN
Wm4Fu0wf+7fhPMbhXSmwoeEF9t8libc6R9joxtJfyjk=
`protect END_PROTECTED
