`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ivmxdx7j/J8HrQP+EYYoLUMvZRwWN0E41VWv3G9pIPhggOp0wZzAJrxQz+c8AShX
6BY4htfdmqF87I/W+F5r9AJdOLBPE4LegOTcjySThGbogBq/57d2IAF1kS+6zioS
Gonc0v3tajkjl73zXAWc69JtlGZb0P/7bTeJNTb2jABuemf6PDGA5FHj2d+0LI/1
0guhgV5vDJacA9LVpr6AHuop4hIaSOfwcTBy/9Pi8q35pNaM24/8v36ROj3iWQ1c
LJdYZ/DCAtxrsNYrCx6ap7uG7U/5dp1/hkbzjb55JiEB5oL5SqB6ozMJHVYmjUJ/
9pq36WejQmoCvKB6v/XMIu8j8dloq5QT/CyiKuE6+pBl86oG6VnC9ePyO1/0/X39
U9SCJ6DDNQdVCE5yK4EBhAAZe16VNOYROfnNrarWfbF18e9FBLjksHVCeE0ozIa3
vHHlruz505S5YYw9HY1eC+1irLGHXmMWCHpgkVp4UBfKuu+/FnwSIVI4g+/r5hgl
XCnSEMZrqXa5R5ldE4CxT26bklvGzTEsfVsAQ4DoGtglzx1VU5g/i2vMQYU77z9d
edtl6JyL/ftDlfzTqPq/hq/8QZcClwjK515Gl6dj5SZZeW9XXcCttzMjHTAjf6HZ
3TynspyX7C6/EoNXSoIedmm9ELEDBiY8Oaa5nTuUPg123xYoS4GTn0CNQ8QiQBsQ
gsEaySXKRLRe3eaEsbIGeWX+wuAaoOJEGk55NRSlrfGWK9ALz54b93G4iuJqNhyN
kv6B5fzayZ5oLuQTtlcx4CNiTqksexQ8INxT5NOv0qvQVqSBCvV4ki7LvdQmRbff
Rahrv6oiRW8Ff2QWtskU/owlRPuiGE01kb84LYfIL44yffSFPzQ9coggy1+q2zvU
koqjciVPCNbObZO3bA45nJI2H91phacGldv2IL0Iv7FbArVGS5nEoNKLAYRp8ds6
JIDSuaOQtmeDvANlyb9VpATs32IPqXTgQ5Z06pFuv1cQ2Q1AUwSA3+6s5/8bEdFM
7/Ab8Zf5gnsaWJ2DakGQSXdEGPIwmYs4NFGuCIcYgek0OGAixYmNEVZYA7OCMvc3
azBF1sBf6vryyn2YhX3je2P0Riiul69U2SNO4GBqwImg8A7xSwQKFN85o0Inin5m
odKr7PI96eJvRChoedrQDR66IBSMio37JzYvcsvf69WANmImZIOhT+qM9xj3GvLt
kfXMOdTw+ASD3jCCOVQAC/9BQg2lQUhfIZhmtg0ZHp8W7juJ7jmT88LPErhZpig7
iGUkwjCWhYnaDlIUyOGG8yTTN8UagDPARZLSBWRT15zUFODvq1wAawMDfj6jwW2g
RDyT0eWwD8YYxGaKTsxjv/kthqskB5wjUUtjL8N7z5FYokSpYeM38+Q8F0M1cZlW
+1q7HxqmXiXt4ryV+NHTiBHF+3MSHq2vQB+iKS9GIxAOJbuEFifpTQvjcRMfs5Zf
14E4oa8q3OI/9UxXNlqgxqpp1fZftoJBFGpsKrpOgPfwYLjY9fm5jHn6w/QL41HV
cpa/t01iay9ZRSJRUZrePDMrpAzt8H9SgH6T2waB/kAKi5stnhnjPnY4m5X+OZMx
k0rED3SNK1lQC0ZGdJ3BbvtOab2zj6ckNb+6CxeeybgjTvCZKYUHCSKVzlGlfhuk
8e03orL4B1bvdZjDZoX6eOv5VEYiHiUYbUPqw7xyP0XBM0QxiUJDy+kh+EWQLfUE
Uwok7NXbyTE5FGa0sXwELQ==
`protect END_PROTECTED
