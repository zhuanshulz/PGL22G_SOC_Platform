`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ha1LkrJk0Ey7Ohcdr5vr9c3AKaz4pf84zDB2xGu2ul0ydFL2B0cPOO+0P79Qgx0
w9J2gF3BYRQaTTqy59iP7tRmVW8hlVjmZmGxZZE4+wAVJ5CB0LH6lIHIX642iGG9
JH9SK45ppB1WS/+xc2xNOP0XQ5jPcknQmoZqyFAthJm3i42EI7C76AI/9PGrydU5
+SZL4dlM1PlCkm+0Y3ZVG/LllzZFBn3WpfwFS+O9kJ6okhS2Q4DRwVJN2IExhIBE
qUFHyca+gk6qQ6YBiIVVOctcDwgO8avqaKsy9H+Df+Ht09XfWJXQ1xikx7gKKcTC
d1w/t8IKycBovDcbllDJk80qNPoU0vL04kv7HzVXT+dnq0YxN/NP+EbCTN4WHE/2
NxNWyIJRFjMCa7w7xdAc66TcUO5EfrolkJZ0w4utIvpk7rsUNeUB7/Uw8iB4WW2X
ZQ4zFrfGpvoxGilZeL6ihVO+1CArnlIRyOxEBD6rw0UOnz8/iUYfRLritm+NuG5y
EYLzw3b8P6o+d2YuuOgKvXucZlwOqOnyHEC6KJWhXh5wpGd+b4pZySdK0hDNLo1Z
MsRR3p6ZhlsEIhDJi3z89xs1uy6kFLE8B+qFPRuWaOYNP6Io4btv+07IVQYyWlKi
A5gSHjVPbH3ZLXWOdroDPUB7Jno8SdqResM2cUeHJeD7d54r95mX4Ln70577LqDg
N+Vr9ORXZdA8x2lduBrJyKLk4xsnLat41fHJx6Hfo9Z9blXUnXCFGsbsGCJ5hFMo
bsSSoXe1UNQmgQ+rDFsx5Q==
`protect END_PROTECTED
