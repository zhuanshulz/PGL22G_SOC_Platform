`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/S+qPuuDuAv+8AWW3hKaZ/I8NmYfotgsLTB5syEIUkyH/ovZ6rDs0elYbPALIDw
Iy7cVvidGyWckTlEEKZ4FYk+iayjvcs1qpU5pMd62A173IwhdbOT+/8j3S59VKnt
CA7Q6YOU1OWx0y4lLIvgyCmd2uq1wfa33ffAXbDxPsy2OaqIfe3wbi3bvICOhjAn
+XsziSjDtuPtbjX2dVH5mwmXG0E2WFhpKdDf7HAzFavzDhYrcKrTvtWYhdUstpiX
etemM65O/SNjnSdOVlG8ZzDYX71JHqDusixG7y4sa0vtyK9XqDwR8nmKpE4UVhfa
JZ9SQSXa/fnb/7aMDojyVlLsMBgAs2zMYTDqk7g/1DdKZa/raljOfb/qY2QohsMT
CTTqLfCGlUJLqnPCzGu6wvNOkJQRy0FPFXCMkQHdjPUdgUUaOngvzNrpgN3LUVoH
fHVHYktfCVn+KSsWnlhCnY9DHgVGobsfavvj/fFQ4m9q6GJaiU2pR1YKDXoXo9YY
xKEZjjnwGlB1VbNmeMzyBdpCH0+5o2HHlTvlx8r95qrKJ68g/nDZ70vLqTwOHilm
RYJKaMtiCfjClW+W8sMh2t4D7s1HXEco6ymTiEMH+UFMxRbhmfXcF+WWFgp/40WO
uRgNutD+Ga/XpvoxLko9zQfJvwamGfYsahKr7cavc4GvtgSOw8TlYDYEBGgxWTgR
lnTuNkWQm9sqk9IVi6yaJNHE5HdwKY8DRpxDqimomkQvuyMqDcow4iz+J5Uz9WRh
+vhBSbiF8n4PxLmj2gid1IyGRxI/kOnooi6Ob1PvzmOQGKoJ/IqPfdVunqOgdMHN
gnI9gClVGdL/pczeotXb5YX9FdUYZ9oE5mb9JqymmJK4mgA75KOnopjtz06GeXme
6O7DAHjiG6FCkjanxteQVMBYIbzaka3PBwQ/kVuwcixU1R9RFr5UcF63R7P4mSoZ
T00mpK6QDvqzt2To9PF4b24nUxztnCRI/r0OeeBVDPXWB4Q0PmUo0gDJGVgOv5mb
0RWUn8qAsbF1ywzyeEr+569evv15mZn+C99c6TYWUj2E8ruVJDNdqsJUb8vxH4Ef
xMlRZuaY3Uc+XlfzpH4eL/NwOWngCCe7X50JwtVHRgNTwTLMvIepaUSWKdCf+p7x
kR+Jl5Akawmb3ksCrtgCtqKBkPhYDrZRf/ZUfS2JTz2DA9A+lIk4Tigags5whKWm
8lbNtAXzbGJ7mxdL/talzBBN7SYU+jOd36aTUVPhs+71GAIU8q7UdTu2GY8VhzkX
XHliE/8EKy80SzWPsCDzMoSyqeiL7EMqy3ozTy05y0YpQfKBZkbPj3y4qd9lbY+Q
sBSEjoTm0tHw0g1G5N8SvDPX/+hEzjIy2w8j8Y4vauiXzy/Wh0ap72amC/ztiV7t
TiL0S6xVllPKVoGCsKXazgUIP8f1SobT4yei+9JrZcUfSScJcBtyYknbJCHzYore
G/tI5h2t+j/N8NfJt4d8hV3PpLCNqeHewIci+GnYPt6mSdp6B6OK9h5wMZgaypA8
Wjq1H7FF6LEGWKdP9+O1w+oHS7R7080W7eftRnQIhtw0TpLWl43iAGcxdQIPm2hP
/CrbVaoPcI8xw7Xx8dR5FEpzDSNYzX1+47ictOIUqT+1blJGnPjQN2EuZDVinUvH
E9etLV0BsOBA6MUOKSJXdiUPYPxlki3IBTIZsDMxnqbz8AsEYhUR4slHofGFhBM9
mYVEnqTp0U1UsO9xRSE8tCeZapJMXugfMqNmkmRaS+QyNG9SR2CpOVUPC/GOvnkC
BY88Ngkn/eWZrplyOYX6ghet9hzzFdqEB3u7AO05PkLVoIVHl5xenBi5YXhgXRju
lGyd0nHQkNrX+g+2xxUJyRqWoweu615Rblp6PMHKzHbi8bd4JjGSDBfK4hzrf+jr
C2zlHXBxnIgQpUlzLbU/DrqbbTxz23tL2G8m2y7fVtDSKUBZclLGPbDMGuUeAcj1
znbe6el6AovYT+Hr4zVEhr2/3K8Xkx3BvC/uJeGKtScZOVYIVU0wppu2g5/wt/XJ
ndc7hOZWuKFw/E1rxqCdOMv4MH3qckc9wO2C29zCZ9hBewaHQKsDHGhDkIkZv5E8
aAeiXvDz8t+o82H6/Yn5VpCqtMGRiJNSsGVcJ/wIyMU1OtXaSucSgzyrG8pfDXoI
5+QBWLhpqt6D9cRjoC7vUfbjqGBhSyPmOWKAhQf7bo/P1B9Y0TCGMSkpqICMo9yI
iJRdryJF/GstIYlcP+fa22RN+sDnjcZcgUwxVrUyFW7yOIela4EO+j/9e+qGJ9kV
AdI0GetkkSyLNoy6YFnEAOPq/7QQiMTKWZTL2cC1MPRpClARZ4XPaF9wC119F+a1
M9nOXwqAqAg5uSCcCs9jRtnyH7dxjl8wp/Gh6ztQmsbHD+cA1Q6nl0UrQnBpltws
eXq+d+lFUPUsjPTkJgzspJn/uutSR7/0Xkc0JNtpCMMf2R9im0fANBB1k2GyJJRV
hBnCpit5GFujcY5lZR3s1RZSw1LFw5e0eHZze2Tb37HFCaweAa7sYkZ3UnI4GwQ0
vdDzP708nwh4WP+hrXT/1LKe69289epzsXXp/M9qmPvOC/GlukJ2EmlXKpUexh4b
73b5pOQpCMFyblaneFZRl3XdOzKMB4Hj+KrJ5LAzb6CL8pNykYoWVLAcabFXVk4B
qsn0wPr9EdFRPDYBdIRE1Ne78aLjU/hw/ZLBljN0ETsdeEUa8vc3YGYNlEC51wS+
PgQKs0yTM0n95NiD82jZOvbSNqPN0XPLnkjuzIDf/FfBuklq61UMEfZZqtBQSWV2
jinZO1FMevCKEXc32BfIxMXgX1U/LspB0bxCyJZJ5eYjV6Cz2etig7ts6mV5Ks1w
23Gyg0rG5PCK28bRGyRBkcDhufJQZeR1l3DMn2zA9aC4EzMhOwWU4RCHl2uR/BGY
oPtRnVmPU1qbUGwh9jynhcv4hHU6IporTla7pn/TFUZBVwU4ikYJDjCFvZNAf3U2
BQ63M88OgTSUn04WJbjeOhEzKHRJ+rUb9M5phubWCzlZgQG6/ok9mh/n8H818sgF
bqGCF5ncT2wnNyWiQUf/KF0KRlf5mzQP9WDW2KIarr0tBKeluFSv3PTQXAteG0HA
ikB3UBcfCrGJ5NIRRrxRY2qT8OtbzcV1MoYzFr62njqUiOc8+ty66z7Vt9+Q+6mS
kMg6poF5ZDlU24tUj6khLaa1dcWvHcuWWiMYS+Ynj8GePHmBDA3dHZ4V8mj3Sz31
vtdCogpurmEuVA/G3Snsp4hqBALpGtVj1lOXTdov5z+DzkpUs9YBe5uk2YJbBui5
MLoRzGk8x5xI+Y3PivrpdPLukrZBDGJn6TUO3ybAjnrqcxLdyAr//eMcMw8Blsvs
nGgbn6a3B+g/CcrDWuqgkJE8Xa65EXwOy+kJhKRdGgNje3nzUW/3H33/RqW1/KdJ
yeHdPiGSiA3FNTCBwNluZov3v30wMWacyZo9NTClbkBKVDhm8ytEF+WU5RG9uWuR
1N7SirpEjo/Bzx3nIk4NuOXOI3rNXDpwHYWuA3z6I3Ai/d2q4CZe5MChYCPF9EJP
2iSstP4K9+qDWsGj0w94mhGqNXcarca+erVScp0/ry6Ajq48O9X+sFbZXfiwpXfp
6p+wfD+bCQ5pdycwAUVJJ9HJxtVPLG5YJ1FISRNp02D4ycw0cnkODXqAfbM8942/
mZnXQ460NCRSIYKy0e4puPqlXJg7tjWbg0bfQYZpkYerwkSVi9UOHtXXDnQPvC0U
ZtPUBeMrs4fzbfpLSJ2mAUyI/AT3S6t+o9/ezkEZu4aATwhseS5QoVGjW5RITG+e
pEnPfHYXZ82T5VyW1DCnTIH767lgUqwOzfN6xj9rIirHIxEn6dlpjermaTURk2Iq
5crKNoSsyC0WpXKoFcRJ7KELgcXPC04MytoS8fDIsboR2oeIkRw4zgxOuxs45+Eu
EMYy0JUe3/y0HRzt0Vb90cssowoCjFaJxU4CukWdq1jNO66TZrJkCnAUtyKbBcfD
luJxC/R0laJm436tAEcAUQ2p7Z1T1ne67H+QtlpTg3au5M/aJMGELV0xfsxpwXco
Ursh4PPBsgp06utnQEoNHs4eK1sH0Ytvh8+by+h3nGvAkbGRqRSzTqRjrcB9QEIi
jTnwlNsLQY1oPlB2OrYnAmf0ILQd0kwohUiZnZ7MfSzKI1kpp6iv2AP1gp+9nXtb
dsRhGJsipqFqHxWaRTJ5PvzSd8ibAh85lvRyQ/0O22Y3Of8Ey9SKGg7PeuC8z9dM
NxgRvuy2B8P98vH7/AS/i7stthxcE8Z/Y7wbfXYrj1VWCCyG4hJTpj2OjaR1ps8a
H/RgpGPIN3yXP3WhB0b4lTsFWOkjSbDPjeCEo9PIxE+g35idbT22bHndu/8HMHuy
kmr7Q3JbZCGq40eHU8gt26T3PsVgcSOSrkZit1Pg0vjDeLlUQstizsizaZ9RP0PI
+IT62OwVO9t+HoEej5G91y3UIfodRyEwHgWqwRo2gqYSl6A7nxyXbzeUcT2ZqK7g
eS6epuqo56d81fxb13lEux9bEkPKO5nd+B3IK9SwLZA2sZ8nzi9ygdHQjaO+IWw/
jFIxX1105mfJXxAeXRAtoB38SdCnScI2Lmb9UqYS9OJV1skUVTd+G/Ni4pB1OgOB
NfK6zAIP2qn6OjQfEjYzve5NK0fpyI2LUcxLlB5LR7vuXPl3KTPJZaz9MOHnpK8T
SvN2TGBBEAWGTj9fwbrW6+MaPr4lS9iI6iasi+CAOGE4opY7MKPn80EjDkY+O/vB
UPsvLtxO7ip/r+AmFgAJfb6E25HHWhHnj+iHJOFfdS81OtbXG3mu8XT3LOa0hQLr
srhLnj5+tgvWTkPoN6VP12gzTCav0DmV1dRJvyly9dLzDOuY3sQW9k2om1XxNtIK
CY1c2Gde0gO4QAGYY3sXDW++i7ynGTet4z+/rvJpMZTQIjcIZPSqqzfWLiNdXPm9
CUYCXQjJgepyzKEok5kFh4MU4X1jpVpyDk8t0qzuEbaDgbJeBYvs8WxPp8Zn79RZ
nhu4/FooHCc119Uw5hiR/fO6jrEFBgiXEi3EFKvvl/ybGR/zF+6YHYrewwYWNUSo
mU2p6w/BIxe4SrYqY7/B+2yChlGWYrj1T0xiL5tnNtHPPfazqxGu04cnmBEPWFqa
6SszyeY9PXrhKcbfX7SDo1ugca9I0ojiSHD8xO1qrXtytsc43jQnQvMYGBym2Fm+
2fbkEiRIsKuaXC+HGHpGgCjkoY1/3a4ruzV3N7J9qKwvgwG5sq3fBE3aKVMttC3z
i8iPGGNM75tqVOaCv6X9suWmNcbVnTWL1FDEeAwpgaRO6y/kchm03kDDLXbav8t7
uYFG6kXv1tRMEa/9ckqt2v+LjFuACvjCgPU/jyb9XG/TqWRQk4YB3BC/21oz1WGy
4wZpPj4e6/JSIyMHjt6IhNoWqh6a1+eErmqFNEf+fxXVgVfAQPt32pLBbtPZVAwC
SGDxyeMlYTc3Wo3HFVdBBQWzJ5Pyh31c3YDqSA589mVHbiUiZa2+fvTQU5AH330p
2RgdJ/I5uto208KQBrUzrmaDJxVO16hgXPSncB70phaf1ng2egM801/BfIs5eCoO
7TaSJPaIG5W1smTgYwK9tKJO2/ce7t8e5TfHdb0uNROB0VY96FdBhvijrFtKap00
KxZ3Az/r6GyYHFlbjmVf4DZ3yzw1xirorV/eudNC0HEoFNnRrJ2j5ycT7WZybnxd
piT1DF3bG6WZk/izBjulXBjwWbTBMFupIYJBlBmmrON260vJ6Q+/hvg9qlcUPxrJ
BLEyUH0RMdHh+9LJsTJhD6zmC4YnjpFmDsINEifdtgr6z7cwVD0mkJ6MXaIZ0PiV
sZfCcabvY4QEKm6FBU3wqmiLjiLLjYf4f3wkedKQv5l2YCPgrAFebclTkC92ZPMv
YaHTwSG4Dhak8wconRLL/kvUp8kc1r5XNTIqXTlKcd9M66EcyWrf0OZ+5duOckRu
1qvPbCJvBbz+SRAHP0ilWT31fRtTCZ4WJJU8C5WUvSh+rAYbjERPDlN7kQjcK62d
rBr4ZrWwa4IInQq416WrK/pbJhjKXhEoEAlrcl146GKSdkJr++CVDZFV6aNexXwJ
kC7Br4QCpKaJmndihroy1/1GRLsAKFqD0HQwPrQ9K4iHcsHc0LDG6Pjt6GVzHpJ1
RbRdgdI7SZjWSqR70SFLKWyV7+hj9amU5U/FO3UScs1OBlG4ONhOJ5QBiHFhAJKX
hpbrSerwTYIGPRCSN64FOCcS5m8vMl+oO4jIsE9dRR+yEiUKE9PwcaC1FRGiRmPb
PVmqHnO2ChuzLpGEE3yk0fuqw0UA8s0duH9v5EyqM8eo0r4dCGDM0Iu+TK1FQTfK
xsVzKZX9+AiOar+0aeZDybkyja3zjdGBe9G0gsbCtr9d4eB6zHYdWXwJ8XI0dS3k
oV/uaXCecuCD3P7FFOm0Hr/7ff07tIDvB8v/I/MoDtMyPXRA+LVF/2C76Cp0rYtN
UlgDPsVzoI/SUm/Np8MccV4pmb2udUOMnNcyXGqcAwsNhvez+GiwzDsFU4WQuq6y
ecv2P5dR5ekTHsSOqXHSrUogKLJh9wV4GiraK3Pv97QzGjFUsl+GBG11pII4tvma
JcMO7Hu/w3Yd+Ffu/37FMLNA3oCtJMkUVM/5U7r1ES3N08jKL+Z/u7xA0uhKv26r
kG77YVvTH0VNwMdwZA/HYA==
`protect END_PROTECTED
