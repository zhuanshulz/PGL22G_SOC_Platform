`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIEgTVdKOTYcVCHceX3q4BNn28v8mRPhCznqLAPDK53bwTy03d6LyORarsEsk5gD
eNoXN96pl3ayhDaqSA7VKdwarzaIz5u2mxXjE6EsAtccRJlH3JcWVucpviFoA6QI
WeaV9q6E8fxPAr6xlfr616DJlkDJ2Y0pq5doTpahO8ovYFjfOqrhUmLQTSFTUd9m
VRLlXjjA3rzmIT0LNn6x8NNjN1RWughOBOudDAnoe+gYfXDIRkGt7cBxJgYZc6Fh
bdSgdw23dI205Gp2UG20lEx0NCByDgAEZ4aYFlbFVDt92Aso3ga/fYZANpKwgo0W
8nd2hFLNCmzn90VsQ6755vsz1u983MUCblpG3oBn23QfB7n0xB+pHmfQ4PUnSIwD
L4cpSRCQzUTPiDGKAo+e9DmX258jNe3pZdkBm7sqTOWYJrABl3a86QYRdRKC0xG/
iXcBp+DLOvYV4GFBubGF8S8pWMLF15zChW5qEvacf5Xoc7TZBQPIWFYK2yKfrmwx
TEdhXwzAb3bSMGv80IPxkmZIt7m9qNbjiM0rdgqHNJwxxwGoUU4SyQAedDI6ijKS
9zK1U4mXsk+ju0nWxP3FWKp4Jr5WpetNNM+4L77GoMj+1fYDrOwTTzzN+wYWcpal
3WK2c34tp0L+Sdv03behcmhSytyKBzt5YWEdAAOYe3MxmSpJ3fVFHo8DVfxhJC1p
E1sqdai1cP75ayZx6GWIuDX9fEtCQztCwX4MEYfM4DftYx0WeuZpIVHsst5Bhv3y
7sONHetvcN1oBhHdLsShP2ABI4AV+v2h7kj4JWMqEsLVWh+Mt5EOxifN7k06K6pc
p4VW79Q9e8Xn0iX7zGQc8+KvBlRbHDE4a2Ky1hjPsvDDBqp6mjSFpaglXANYYjT1
C3+wECOPAHi3ZJ7jF6MNyVqChvCbxwbqYZO/+8jJ7CRabmsmpyhQm1Yzzgb1v00C
r7jti8npoZTJfZd4rdI61ejCL+C/Ghh73ekcTFcVN2GqpgsNtU6bu0GOFqhLRlQH
AwjDiDJXdYrqFVZvHO7AneCGcsh8Kbf7MRbRgR+/JaiF7JPhofJD29jJZ9zSf0EB
1XHxiKm2aejYEW6ZeoFigfEZ7huFRAPdyVUgU43MVXdyCDH2sRpITUSAQpOrZ+6+
E4Ere6rdZCfUVYbcvNkBjqgxyacbUaR/OrUMbbhLoIDPR8hjRTfTnyNwLFGFadY9
uZm6E0jQQlKV3ZWBEvkdQDPKTim39HI/fTxx3bQYcXnl0zYzauXwJJ3+m1P0Nh9f
uucAbmDJZjzA0+CckLljKMXkBVm+aV2JqehVi5xEQn2T7s0F0iYwzQB65c6RwL9E
LUfNqyIfNG6JUKDXJyLrhb9FJqyBZ2D7PjebXChu8BTihSK/gmyr0sN6IE++BJ2k
oE4tn1l5FLg+FMOQCcNFS0wdH7ZhjsG+Ml+JfGTO/Q8AyMpLFQMQJ+n+ne5I+5H3
Vy2EI4XP7aU9dWyv4WioeI/XULRz9cWJGpCKCs/mABm3DThC5mk7l8XONN8POHLl
0ljsNM6i0Pwk6iKJKeuWjeZgLz3gHJzNbphuP0MTyPEv7z4JJuUZxYxJxsx/QtdS
YQTat0wUWbaBjzen5kGRj5g4UKNmLlySQ7w9uFcupOT8zC+qBXM6vEKf/lImdkXm
RKLzzINKN57O+Z2XvXvvJU2nlTDLGyeMpRP/tEHSG7x598w5UhF40bwx4Vv/lLev
JVIyfHAALwZl4WOxP9UzIHJygniZ62lxdORiB6UpFQQW8dPVkOsHNdy7ed8vvmQ/
AiYrmPayhiy4Helt65NtwqTBW7UvYnft8hMr0RjWqCWlB7vqo9KBvAULSPvSPau6
vuAZzDSKkO9Y6Pq6bytRv2N5bornDOJLIJq/ViR+lNUUWpfJtDyIFi0OihD1Cuvo
AguqhaexRWQrT3bHffNBXC/bQ2nun43CsCpd2bBx/4EKA4Dawg8nq8pajqHiKu+D
kxfCJQjYJx9JEuJRU0XhUeqemKNEfCAq/qOJQT4zVQlyq3AoX7g46sR3N5TNDS4g
nAl1+0W4n0e55/2UJzxlhG7YNwrHO9D92klVWCL/wrJRoFadmBIJXfU8Csv2uHB3
tB5Sc+XB2rNnnPckymxX+swlAVq6erIAc6Xv3BQhswV0sC6zQRMSWFEwGC/jElbq
c/uS1cvvUcMg1sjEKCNrWqkhgfcUADTlQYKOh7RMjyPDvxkPalevvqveBWx6wa02
O6GXk8cVEevupFwR5dbXhI0Q9W4tGWVB5lF1218IQtoSPz3RBBi8vGqJXIkvC9wC
6GIhelYadc9PxOMLQruzVAdn1D7C5pboC3dk+kEWubsnnE/6Bc/FOBk9cfjKxtJk
cDRE6ZQFtjMUt1j9MGUhtYlzw/2DYFwLdPkYXvPk9Vo9yRvkPwJ8hpl2KDJPk0tQ
0Ks64bv50waU6l0hU0Q4B+ApeND2gEE4ycH8/XRDCbzRs5NZtiNYBMx+5uWzCs1J
EIetxGXTdrKjf+EHN4/5PsbTlmtj3FaPGaXOy6P684+fbiYAr5Wx50oKNfYjgO9K
2l9kpGQ9pUynbUu17zpNF5G7FtzBAlqrklRVdURRd7E8n3pzui/1QMbQA3XWHsD2
qfavEx9qxOuL97dQBhvDP/kJpWmyVOPdfMKUdC5mf42x+XZxYqZ6ysMPb4jRkAyx
pW4nuibRd349tx6/HvFmliU15ajCUd2Nq2vslrTsoi9jB87xng1WALqWpviCTPbD
NSQHoJLyqq/Jeet5oqKVr/DJW/3AFThEwvk7J6UO9sH+Wn8PJ+xtDsLhzcuKr7di
Esik8bzDInh5nLP0ikkQxmh4YRLXGIn+R8vBEop9hbrRb7o9XHbMh5ml0Fng7tLJ
hAzFoLg9skmbAHYow3BzciltQaqoIbEHUedJxcG2CkQB1o7x7FHKJcDfAr5NHCQ0
jfBeH9LrtxjHQSBt0haVVskFsQHVIIoUgzuA1rTtzwhIHE+liEbxEJCcuG1vcIP4
TrUwWrddLSSKt9Uw09sUW6biKy/41fTOvD4GJeEQ+/YfHbRPlw/ZEYE1QCtP1Mj8
vF8iXH9RlSYTIog131G9+8nDvVbH2MU1++wyAsVSPXe6/9SDXDrPfY/QOWKuuIzz
R34TOZkFr0g2E5fy81wk14owD1dlxhCm+qs8rZhpWxEy6k+fxCRXBEeequMVyf9a
DeP38wlPL/+u1vUSKU2q7AsgkFhsX4+YB5IifOK5aiqhUTKQWZ7twfNjmbZSYpWY
yn6qG3E/M6/2V+sZJ5h3m4UUN7zLpQq9Zq/9kpP7CnNAZ5st4coclVyGbKR5ZxHM
Jvoj2Yn6XC9UYhWo0p9wfWYzRZrD9XNTiAshi/xUmqUT9hEOdtFj4JaMcHW2yG/v
qhTReA3ziZGwourChinEBzZUuIAtyMYF6dKHhN9Asi+d7Qkf/KexU1h8H5wO5amX
s2D63zMnB2bwfmGvOBEt9kefPAlwEco9897JV7aEolLKU9IP2E25be5hv4uDgSdj
BAIfwL7xDaarDNrnzap/3gSQu7Ais8aDH7Wr2XJnhmaRlHqScUmGQMf7xqnhXINR
L4LMUy5SLTh8gRW8vacXF0e0xhZXrOeJjk0tux2XkpYp1GoVyputOosv89eg9nDE
il9ovBF5F2gBAiNGvXLUlkxi2MRPwudCbh+JUkOvG2pd2rtZtwMCwfXbF4yI2CpF
tPxA9NoL9K4ktUJPhbKdbeHyorbZk0FHeBokt4t1ofh1Gq8OGONZcLLx/YH2fy18
ppd5plJRqpP5vzbH1heMeHrkPIF0h+8u0vPdpWlXLGW/uYQXtt4C2v4IIjxceP/a
YUM5uywbVAj8/+JUP1komhYwHoNpJFgi+NUwMiK6B4/1OC1Wlgq+6pt5AdtBW5MN
nLWSLE1cY0rtfFaLb5e06chC+5qgg1JnEdYrVMfbDMuuorTbwGzdhwo78UhvVsaG
HFTcGxbL6s2fATIO8UISORN4gpZRXmqQb4ee3Z6TPtiPQ9VfaWX68WPgh6aAgs9H
3NYv8Os1NbtKPxbY3Pmp5mB1ABdNdlG+30w1pcEE+esCBCGgGGIwGhaAzhlVUL9r
eK6z1WuQh/ZrgFxOKakZUn9ppWM3/nGxqW1a0Ng+VD8ZHVbdbqpz0Z1csKd0AnMa
TxGJsrGwr2xj0ZxTwa66etSUGjKBCBKan04n3G8ntbWfIB5KVSuQpxaA29u5Rkpz
giByJpyJ6yJFngel7sRZFdr3nR7Va/oG4Hy0lqb4UpTV/eUNTNgC+8BALjGqI4R+
ne6mtD9/wWa5lcpBYzQhuwTzJd3hy/s8NKwGw0E07DWvbBTIJzOH8JCuxmAtRyk4
LHKtrp+zJCDsD9JuK40767dpp8eNEw+aSc8gJ3aYZshTf9dhqqW2S7hoqYB2fIrU
MZ8m3dLJCNN7ohnWdAYBmEc1UMdv1/X4BskuQ5mYgIrASRb+EtQZpMoqCCiWmvI/
cnIEjQFPo55tsgi3FZKfAfN6+4FDQKlbA2+FhRwQCrPWTGCLz+7NmgBfdiP6XavO
0z0LyhjJgygfWbz+oEugNcIlKNj1hKnYh5kfHozsZm1fiClh0m9Wl3DoUlk8scEX
g+v2u/abx0lA4Ko44F6c1CJ+qMBlS5Bykp61h6uaK1bR2HvKmfK80RL4OCVa8KKg
VnT6Ya1UTU9lAQdzjqG7qDCAM86KtAUIxIzTZ4LhQefNx1u3WtkzmddI5TiQPhGV
pZUYL4eAomcNw26m7DwSmdP8V1uAdBeHfIFohDHFCTKUEyV+V/jkFov+1vCwZexi
LOJEu9CNTZ2iLjH/4kap6Y4VK9ek6r6YYLd6jZiutyqGx16KOGBxqh1Ljk9RPIIR
4AAtdlt3Aa5v0f365z2ooCcjwBn2r6Fl4iMl4wp330VylnEMPIwns86zob1IR21I
RdP6ZDHSnQ44nFzEwmfwyMvOJ18PylzMj+dNEuzxREIG9lXUfiTKN03HU2DZz7QZ
03pa/D7n+EZFAro4XZIe07WStvtTCfhz7Bw7zr0DwejcnvTUP834M87S4rv9aYCJ
8KBmb6aOuN6H90jsR04kfVauyOWAMllhlpmO7jtSZy60IBbvZzj+krXDcQvdz7yR
046GDnR/var4jfyVlDfJn+0KG/AawxfXGLYux0lflTEXkF1joLgPov8hMvnS8ulg
Q/kxkFWW61dxHRLVHkjh2BRRPoovfM8k3XGM82dDFakarfbgTqb7c2jGFVZRMN7m
mQQjZWWuD9CxLF0ji2IErOIHRGh497vRxEhCOuMYv/2uJqCwJAW864iEQUFgxObE
rxO0idnRaC27iDzEpd3Kg3l0lWEVuuJCQWB+xd/BxHbf0VrCXBOrLqea7y9utObC
v4Ylh5MCX1rxPzGN+RwTrKO8VskxTSU0suGTEFHhbXhz2EpmtqdJ1587VDJIa/oY
vj/+ZSVznF89NMG4fBY390R3TT/XKCXz3/ggDIVgOQ4=
`protect END_PROTECTED
