`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mB0uHgYw+H6cycrEstIQRdgdRRNmljWslrmdK2OjDythw6PxHkFqyY0QiGGautmS
KaIcsYEoRHPMxXwFDQE97XM8qqoHegZUTne29JgMJ6pT8I4peTFdyUDu3pszRjFU
PzowIdF5jdRmZrZsarZMUlsxk0/AzvwlxR6ruxAby83iRaassORx5zSpkqOmoeOB
/NhcXF9+m0dZuRQiUxHZZwd4UjHHCWNLhPX17u48y+AAyh+8hHVKyL62ydVEEalB
bSsxx9z6/+lWDVc8V2uZ/1dekD4B+ctByt6X2O6xJEBfQ6GsRL/wQK4QQXfFsRJK
bkM1/jAn8jRMVe/Zddv1fcV5qGk9AEzrolhUI7VcQuOp/AiTZAgWcHCGTvYi2qXD
AlYa95LXLLRWRC62knUMZaxeTk3AgxClatbNNIec2Zq6+IgHn2G9jCcaCXRkkQQ9
A1CVpZAYFF7BBwytQOPxvXl24XD8RNNbnUZWK73hz4cAAZABwNaCKF/KrYnWNkwO
sHBpVYejFV0yEeAmxCIEX/ePr3wwIEb4ANpblk7WFLGnrAnSpenhi4m0vlx8mEft
cAzET4gN9FmdHOMO0Jt5tTcqvvkxTVMPZtbimGUAEbdXRfD5tnw5/ErsrUt1osBS
HLjcNEt+cvZAi/1q14lWHp8nliA0ahowVARH1j4KB1345yQnq1OvlUrJqSVPXw2A
TCC5Z0f7M0sm8+9ozjP0A/9SUaqOl4bPJQ/uX/k2lq1/lYDK10O9/dYG5uQdGrkq
lESR/a1VHeFyY3MKYfFZi6R/umXnMBxfaOJtcXyDz5HbD2+rlAoECRltX0vWzh9O
XtHz6r9rckN53zatj/AG0rmfrm2XHlydcJSKFYekEs230b65ccmANygcYikb6H0B
ksDipNJjn3gbgIa1+bBOgdDXvMI+keHxAVX6q6NcWoiYHjvTnFt3hwnx0i9/LGfq
put87LDv7MXVri2I/HnnwAk7xO4IX5kBOeDTbGkl3knIJ2Ea2QGCmTd+AmaXXczK
lFrjQ47rC0R3gUxQ0zOxTOT9JDgnoTSMepQvVhHMXS+z6laUfHI3lzCwoaVJVwLk
8Z0rePOdvJw3l9WyWEb1joCx4CovPYHTF/Cz3AwfTIkUFgTOl1l8lJb8KV6d/qjw
vF8qUwV89tCELs0H8MOEvX0Alvlg4aJhNmop6NwORVM=
`protect END_PROTECTED
