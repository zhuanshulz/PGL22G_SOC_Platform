`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lsyqts1nN70ybrh8HWepqiVuTYvOq4QU+aQVaQOrxng+bVGZssxjy13bIBr0svJV
yDbZ6gqltBj4GQVNsNC8gLM8TQq8D71lwVWi/CmaSL8RPBz88Ixe398W3ViQOa8b
F5N+Cz+6+Rnl44P0hfkjCypwO1ZSRbti7fn9LbOHtL4+Dq/BzAmUYfhVShSulMiH
WZY9gpuDYMT9RTx2gQR7HgrEYKEi493n8cfghK5TAMuF+JJD2e6NYwWzGbKZttup
TbYwjCPClSGsCl97yhcMpLiPtYUkd6/ooRCzM1UvwyLGVLXPxFejGGZeuaTIBCyY
PQ5lkjmlkG2I+PsFq8kvaIYUg0VgGUrkTtSO+PiAtzwe9M/3cKTWjHy09AMfTpCA
Mawv1H1m2TQzL8JsymZdE6xTAEoFfCWG4qUK0HK43wpE0p8IwTpCZAnEvMW3ZjNY
2UmhI7mtwfa3GLCWXvnw0VRKOjgjszhlTfB+HI6r7hvDD2tk9EiBHtgeAoJzR+Ti
vtn2D9qAQTfOOqYnpkLq5Q==
`protect END_PROTECTED
