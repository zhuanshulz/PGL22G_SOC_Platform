`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LeS5yeONLhBhTz6A77Y/g/GfzEWB4+eaZcHiZVuB2kk+p+4NsHDvEF7PQgzeI7Ef
s0qXEBvUumWAxcXEE/ned/5Ggp19+RjOx/xKTTnPYZBcynFQ4rwRzr0Pp9KRhaIC
cNbsOf9OSnyw6LgGLgUV/ld9TlaL+veNGnB5po9jLzOD61PJRKeGw4VGZVowpulJ
+gxfzVODorZfPRJLsU991yLpD8qrgfDqBLLRKfJYMkLddrweSvA4WeZlLDQPYKVe
uQ2SUIye6/VxcaWK+wZf1EHURV5NMEtqx7QTt4Fmc8Om74Eammmo4eTyVGAR3hbK
8GGUeTndCgS4XDOpD7Md5sFmNz/rbNlWIOf/7IlyazbSUDg3nnNKogskimm2jy33
ObEMKF+xp9ooFm1xb3qnue3F67Dm2HkFKFmZOIfyvXXqhhCZJyfTdih4cjdL+LI4
ue1ir/BWmz53nnKsfcVfm+Z7sM8ck+B1EPW/m3896V6vqNUh9jnH42RCmWtwyP1K
SwBUT8iBHYt3ikhpXdRJZQ==
`protect END_PROTECTED
