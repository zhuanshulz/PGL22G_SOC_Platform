`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ycR18e1PLSwVAGJUk5YV+bH+0TNiHqSIdGoKFgyf4UUMQHrpPsPsJV1o3tC9GFx
DodGpbYSF1W2zIbu6oBQa5bmVKvcefunyYRHbkZpjpaKFDxfD/GdZ7PmBZr0DKjJ
xMSRi78lWeEUmRHLc3M9S1x8Wm2qhmq3MpSszK/vyguvK8VWu2MNg8uUabN+uiZ3
T0ui0YbnZWikAP/6PA4E2lga1Cswrwu/mhd0g9cijBrG+Uh3PH3JZEnA7GoYEvtG
NgWrwWr7wm0SpqNKyayl2eUT0Bi2v7+t33KY29q+Xju6D70gBRvfhlGkVBVTidRr
R4nt1iMfCaU3M8noY3d7JU+2G69pC7l1HyX3FDqSynb1oNcIOj28mnXJaI/pM5NR
l2ODbT/Yt1YczavfqGYr3/837zlW0Ob7w4QW43f98V41Le8NTQ5UzC8YDh2IVDmA
NKfAT9Ur4vBq8/2kVcD8NAgbFd5iqGZquJ598VhnxdWAAQ0Yq8TLXcHNzNAZEPJN
Zm6QG1nLlMH9rLvMSUR0QqheocLM5sznpztWi+JG5DFBBi3l0BNSOKXsPwU4HR1P
V8EzwSyO4jIrn4c6KS3i2cJAXNvylGh7AXBYf+V4mOh8y58xY4FjwCbKgq4mimFa
Q8FidH3TrL+ERwjZ6U1GLWqJDAtg4XApAE+koUgZfHYsQ3SneBCss0XV48qqTVaG
ZEMZKHGMR4Oym2IrQpyYx7Gke8NWhVIJz3NGSLZ+Ctxj6zLjFe/WwPkoUkivERB+
NokWlWyFiPH4PkAL0/Kl1lpam/Nbf0Y5I0MFN3gVdbcMaftRfNB0P6jrwo2ZxaYd
Gx6Ia6iuKfOTK+zr/rr5R6inUAKKe6Gz5FnRc8K0X3wx+ZYPO6IdqAeJix7MajNo
wJfAZg87wyb11B2l3j3afo0Id7oB0gf/JO+GwGt5YVZ0o/cruGrAZCMv2l4Uzn0E
+Su7zF+ATpQ8ia9LR3xZmNxabxxT+F+SVF5HJu0qUeA6nSAZ7UZ7MCtmE78QIwdl
shFAJPKblk7e4HYmxfx9a+VTpIzmzHmCk60WdUGGg8X2adcjgZbrnde21GDQwBhZ
TU/hFANwx/ngWNEmPOzryX7+T2gVI8v3SHLcH/A1jXOMhRejAKFkkzcau2CMrq/F
34NoozkYXhuZcRYg6tRfecaCQ4PJy8Ij8CuWM9GDFq7Mf4d/hdJfxMhh+EeDYDDD
dJFj5XPumtCIk7VrbaW/zjPpx7PTNlqLyn0HnboEeZB6iNZwPSovi/BhpHtvkaEL
ymR7AAqGY+F1zNW1r8qdFmjfR60fr6yKZxqbzSWCYOIUAeM01G2a+8oMpGWr9Oi9
ZyHKxLDf/MzaR7oTtearGKMHU3eA6aQxnqx1PMEvoxDVZhN6uyEuJ27Ro/gjklWJ
1Rf9/w1ZcCYSbpP5MB1KN27hzxU37/rauz8QanpjWZ917nSOd22+UBt9y7cypBlA
AcAqgH8iGV1VJSVK3u7041oTcW4MLYXUWtIcFlx8e80eJMMy0poulEpyKzZ9q0SK
+FNxQPE2HeOoMthSEGr+lJGCyKSluSrrvl0zTIlRKboLnq5tYsbXUU4rGbL053YM
YNbIKp5sxajoq4NW4tugucG833wRFU17cuHzTBodc2hi4XIgPwGFf5raznwrG0H0
aY1D1SBs7ZHDInmPQmPOpxSnF0AiQDmD20a0JjB5t35u+9ES0UTGDfuuz55rG8Nu
bfUldIOJGGBpDNCYtoEJaA==
`protect END_PROTECTED
