`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rfpbQq+N/dZnXcuEEI9R/pd7MJ4/h4YSEzbBLxEg+9GnQ1+P21fiVAwYiH9mlu98
DldUutMuDl2MpcX1h72Q3qKgpss24Up1N+rEwO0+k2PU47Zf2x78pMxiix8wiMM1
u27rDQx9VlC9mPVoHBOuHcCAG5f05Udj5FVo1RErNoYNo3UKkl2fqYrWCf/SR5C0
sP4KymizydqNOIDDRjpP/hGgEo5/rYe9iccvQHKpN+jnkKYaTpAcimlo+xWtKGH2
h+MYjliYXLT4vJDFWjxA+6E1L9VnJUpwAZVVHZBRFKZQcLq6OkEW/Y5Aw7WSif8U
XvqQB6AHqAFzu5O237YvbiN+BdjaTZLldqsttG2dVji3C6rZx4iPiVcBZE68EG7j
NpNFI9dMLetIMEYq3hxr02J+BT4yexxC1rtrLxK3ZKdlOGW03ogSxqJvC/HGTrQW
7qtQ57ZM+O9GCvq5uzFNeCYD4kidzuEj1TK69vIuUNBvAdL1fCRmYcKt+rQd4bJJ
zCycBRNvjmzqArj+t5OY1hv9wI1Xt/tAc4fD6w8H2Leo0h8nTVA0uQtDuoA2WSaV
`protect END_PROTECTED
