`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZL3sh4weks7c6nlwgWd8FvvLr1LXJL6b203P4F/FL5YDvN2fomddoaQ/a37weHX
4qIx8mZyvv1DGwzzVrMwF0DPcsmEVCA7M7xVVfzE7WjKz1QayWYdXxmzaItTqXIP
n536xmv/wvKJkMuT8/IcXXFpU/EOfrYb/q7lHeG7vvtJ+GyjK4Hb0YhPpkmjQVvc
vaHGSx4Aqkp5gpaa1BkD1UncqII/Sygl3rb8HYMfxAVbapGNWECe1T1vE6s9KmZo
Gm39tPt5w+1rSEe+4H8CRzKVfypCEh2R+PVjGn3eBjLYN8nO46z16RzfXKSPAApM
ee11yO00H/DnfQnx2mRtLU1Tv4QowC+v/umJYXt4bycUJyh9UzAP9HNiTPckXrdU
ZWqvaiEgzjeqmLuXUqQjoRXiMFT392hQqYdf+B2MqSnFATMRTxHxCZrx84aUbA8U
RVtqeHt5ceULTXt0GVDgmE3hGmzCmoC1FDLkW2ZHs/D1l9NvTyj4WbMqU54DfomY
Sef6neFQa2l2Qjjm0n9rvjxOuU5sA2hqhTMB6eDRjTDGOn7+Y74aMxH5FURh6o+L
awK+pGBtkvauDlDq3SdrYwxJEJHy+ejfe9rvwOF0/4oWpW/WoTrvkKOjIOLCEy0n
ZbPE/zGUwV66jB8Ci56tm5k3TiSDDBgT/isYaQ4fW+EvDDjF5GH4/C4u6cCl/TKz
POyERn+x+mAH4sKjetIiZgHKZN+BbibH+yCCaOxC4o6+Qe2Bc9Yz8esWmQuUzKxL
NoD2qYWoebk1mE6UKCk9lEjohWcVV4nNSDbavKm33LqWyGzZouuUMknyB2TR5wDG
RjB1F88isloY02NbZ+rfpojpTlVisulH8EuyPWl+Tll7zcLy6V8sMY3RHQ3yOSg6
FeC66Djyhxv0f1rgn5Nc1/fJlycLLWOZpdFjobk4FfdJgwXyctXdLAYzF/TdPsWU
S0JhjHxVzJT2NsSjVw4dX+EK8xYglGSudviawkdampXsvLMa0NYCvylDY3Jb9xTO
WABZy3PwkAF2esrCerzIqQ==
`protect END_PROTECTED
