`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h2RRCUDTcMBecWi73+8M9B5U95g/EKusLFaaEBj0iaHWo7isF80BdQ4kk1vU1AWN
h4mDex5d8U39hELk6So/Xu4NxKGEyHXlGDXyRKZQKHdLe9Dyrjn5w/uZPBwwI66z
+Eox3LHtczbXCO6uLDxuPjQj87pyuOVs9cNy3nMBmzKfsIEGCAAxzxtw5nfsvQHn
3yRhuzaBWS7DKTMNzNBosA1wbZklP+95Np3EXb843A5g8SaYRVkKcuDs9kWz/CeH
KnScqHBww9QOqW+W6TNMa4fmxdH0qZemFrurtGWLwoFeDGhjlj0iudaWIamuCX+1
+b/VM8v0SUzKiSbqMYvslE2udkAi8z15vrqZyJtHNZ+dgG2Kn+aln+awVZOY6sc+
x9PZY3eHSLIZVfPknYW6Or+KQUGtKK8+Upu76q2s2IaHHBVgvjBq5OnYCe8SHPAj
FDscYQ8iRMdAN8fjyOpKu0Mf137hM3XR7s1ZmP6qFjJfriYT675rGDeOtxce1IsT
NYG8/9esqol48zWFGCCKO2tbBOdiC54QhuNGLRd44FISAM2u6ryLVkiaQ0xTTgap
TnqYyJzkDbGVDGeUm4OZOrMl92YRf/BRyL0K/MGliXHm+cqjZjUw8MhstAoppr/U
iOCoPPeNFCx5rBCmx9f9RUSY6KhQmi50JtPANDEuGQOfIbOCijzNSSxi3dw5/faw
RRpKQUcueGVp7AqLG7GXVO4cux0GgMn7WfOv9v7D6Cr7Ma/Jd9duqCkQ46hrHJtw
N2nG8uZcq7lJW1RMP0wGn0o8Y+qONVqSRz/dyf+dDrvRH8CkWvYTLPvHBIxsjWql
MuO+CRns97WGuiNRbUu+OG9OR5buai5Sl6BZmtIiCIS0csT5M0Ptj409qnBrwHnt
v6QJ6cmTo6HGfLG4v5fujNKu8N25blSe3kjB2Av3HaGVPHD9Xn2FgvY6tkc6fExA
uHxD/koZ21ThZDPhdu5dBZ9RXcc7cYE2FZSyiIMEKO8No317JaGUV879g5Kf+nQ6
KVfIfT/V7x7kRCLaKPuLMd4qw3mIgrMdrrUpX7dO8UeIedqzJ7tKxfSpkxMXvSVZ
7f/OlrnHJrqWziVn5oh1a3cGTN2l2uH4auhMDXWjngqXQnpnzQcnt/4Bdp26yDf5
HumgZ7L+smj7lNkLbUgHUg==
`protect END_PROTECTED
