`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccHgaG88OO4F9h45yKfr7DZ08wMNvwjgCxXI+YWpAWSODE1d8SRM8lmiA0kUuDPw
pm80mFfv7FywRjlD4z8R+XTXu9/k952ucp6wB/2LByW4l2rPiIVoJ5zkBqFCWsMX
SFTTcgqSsyfenHRwDWwM6e1qpadtdj8dPyM9RyHPJbfFfOdXuzTY8BlWNHqQgp0B
NzMrAITjiWM7CzyDkNvAIbQwOdClnUUUlnQ8+X5EwXmS2g3t1HHrhdd4OAghA+w1
L9W2tMVuTzzyUodcSeMnOPV4WMsr9QPmogkZ+VnPRS9n7dLVwpqTzfZfSIGUI/wa
iFWpcxUAot2fL3fwOV5Du7lDdL+phk3jyKeowkBBHOMR2JPneezgjC8euQrb9Cbs
`protect END_PROTECTED
