`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZOqJvY+FlHbCWRu83KvYiJKdxR9NzoAKB0+Tsy9IeuOmU4PcofdY0Egk1xmad3T
SfuX7nsUmkcT7bNVZdIvfHOY2ok8OmXSqsv0Vv6EoTUyZEf6P2McChd+K4gD7hpI
W5jpXqrqRfJI+6dBAXaAcmcz/ek2oBr4sHSlnj3y8wy0qNChYbMtrrfquPf7+3pn
PRtlQWhQC/6f2djzxVbn3CRRcMDlzHviQFox0DXCtWoI9CnboStmJJHrztF4dKwW
sfrMXDENBxLUd60JMufj9LEJCBkewcChTMJTRneDTlRwr2OuCXLpKIa54DHnglsf
eJM8Mn1q/aE3M2BQMl/kWPC1O/9fDmJ43IoPl8cV92+au1AnZcK/gdQCycgyhn0P
5G5LtKiPRfW3aZ5fL6SQTLmiRBB3oxZSjyk7auQHLvcWLl3lbchJZ34JI6qIwULg
2eq6PlDE1WtG/lYz+7dZKStYZNuEVkoYYg4aFEQTOola0B5jZSO9yVsKBixSv5XG
wrWgOZzwkgGYLwc7+C2q8zhUpMw19EKdSCYPTJTqnw9CCmB2AAX1xtT3jZN+OgdK
2PvkHGjLS7W2xlNQ1C/TW1SuCGe0IANtIPkSLe5hPxEa9o87CppDYhnibVwHbJDz
DfxASd5djz2n0uGENA0DN6gRdLbgmp+37Y0n3XVtZQcNgta3IQxa7p/MZL1sgyWF
lnImq7+yWCuzvD2C+454oNCTiYyEbisozgWj0hwctazabjAr+vG1uCe8ReSHy+3G
2TCq8YqBtqQn/BhwJV20prPa3U827+BuyLKayyBWQEtn/6eX6nAw11oIXGre0HmC
snK/S3oCwRORIAzZ26LJN67M+m6q1Qg/XNGodlbKJxcJ1ykL57Q3O4792s2K0x1a
wEby/xmMcZ8UAGFbFD8LC589s9LgofFUXZK3qb//9u/I0XYt+pp9JOc0E2Rn5ycS
aqOdzFnhRuKcbW+phQ4NFNKhcYe7MAy4jXPbhXXEd85IEEDd9PhwxpsJtDVJK8Kn
udmtQ0R56KCvtjbAco2wt1PnGoDcD9STnuE1DOvjk5eWCDs9LaXM2LA7r9eRve/K
CZO2ach3tq223CCft7ynQUClYZI/Z7JnOOoKOxfslL1GWBDXeAIQ5ZwK6yGzCKtS
+6pWTMMUqvQO5Fk+x1iphQAlmVo2siozRzu3NiQL9GWjzjCzj2LwXjNDx+6cGDIC
V31DdYlKkKtIZKfrYP0ch29l+FVcSxEumUtvXTgpUnUxnoB9CBstvbhvXbbGRakF
OZCoOQ/0Uw1Kv8PWRAI7VDPjmldFoR5qsR2Py1m8ZSbJqUnJpyc0Xj9mz9GY1AoT
sHNFu/zd1KSUlQGlKR5Hk7sKrIMfNf3ATjxrtdul/xBsJXd7f3lIGatDk91h8inY
3eIIGPyiMJveGb2jx6oHsFRJ2IzlI0wfCZXJ++rlA13TSPrQw2GfsebTmugAcXSK
wu0ldT707/1vzBV0uqdMQRmYG1JxS7eS51wAD+IbeaJaZ1F/uB82USWaVNU3cS9t
QCJr+YIW301vE1wVe987HBzsD1iJw5jj//ELhiUc8qCLFPllW/4AyiaofbUwFIDd
/viTnPcymOtjGvbHLcV3XBTfEin11E7zxujkCkvapld2t1EZqkanlWkrBi+49OGk
T4rC9BP905qGQNkPOHDw9w==
`protect END_PROTECTED
