`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1gUpXDsx+KmFM/A1mYYdks1yyQzbimjrNzIBWCrZhPrE/MtIxsEPrdc7XrBTQO8
a83rjqhRkT7w0o0+ak+Y9ZZJ889L3jHXZc4U99hQl1JYxA7njb2DRdbUcbf9Uy/I
+rGsqZgwpzjiGhr3/ApBaekiFy6WHol2+LV4sa+TtU2vOt/G9Dj1NOxQ30Pq4QXZ
YuLjEF7dactG4KxoiiBn84ZvS/Gf3OLEP8TwNAzzqYrfoK4NGzDFY+S7FdYwhQTS
TvjHGrOmkJz4VtRveX7g5M1jfqiDulqYT+lohFUf+sHC1UlDkwsWvf79n5Zktoxr
88E4Xw61qYsK3nFHt/nmpOrz4CKROY0+MEMvKPeux8JoOHpFfveTPaVHWUy9qi2F
Z/7pF4gvG8cT8/PtW6U275xuzOsHEfUgE+C5Jo5R4raJHbja0dB5AC4wzGet9I5H
JP8x9GhnOTz91oWAuhgxbIVlTTb+FhjOpliJuqPUy6Fsc/xq9wW1/v+DRcaqVGFn
qIWcj/T5obZAusCitBqIEUaxg8eArZlq5nJumMNOzWamex9zolyNLcQejhs3Z6H5
n5Bnb9cwitRuz1/1r6PTZMl2Nepn0CZIfrCGF5tQCbG99DNIF0AufLOfjqi16iZQ
AgTbKhAmPkoog9O8PWipa3XHueuoBMrxL7mMAnUPaAcTtgNNyrd583yDGibFIkXa
9NcF07rf2vW6855AP2NprfsNj1Fb+ViGBs4dlUApRkgiYBEI5W/28L+C5d8G1Xp3
8bC1Ec1ph/MdNaZaJpIpspo3/a5AFt9Y0DzW58bin6CxofQNQFmqHh1HE+fwkxL3
IuXePlHzryXl+it6Yh0OTXy1bDx9zqwSQHAr4ywo2C7H35Bnfuxg9u1WcHFf5ZzN
oO2ttJFZ3hVF0ev3LiKwaxSJg/gMbgPuZMVaxJB5PLVtKO7puobuIXNit3Pm3CXg
asn2s84/r+JV0aXu73b9z2UoetvhbdTsAYjkiivqh3yGtFMnz+lloYDMKzrSMroU
HJ94/8aovgPqL0fq8IlIj+1/Gvu8FQw5vlbZJvTqyU4bvocgVdiV3FpLbBb3Kqks
S2KzjEAXDonOqcO7C7qZLCjSDj+PPRHZDrn0xsVlhzW48qjz5SwfT7jHYwb2RTrD
mRwUxViWYfErVNVzEVuxrvsHZQB/llS8TI+UC2U0xUaQLRxxSrHqg4vgz8guK9fB
GORv7S86awzkvm6D6Lk+AN62Mjxpypugd3HYpSxrCUQ7BQLTUXqT8ZBkZKnNLoxU
je2l1YsdpSGRPzPqlWpiHzG5Rd1dsEPsr5zJYpfgSfKiCH7k73bUOzcRs/IqCUCH
ZwyI0P3/foYXpcHHdMKFDUzByWrGDmYxFsS4O3FUTLSrv2jer7i6kjcmGivNjIdJ
`protect END_PROTECTED
