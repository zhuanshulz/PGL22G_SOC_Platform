`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g2TyNZNRCanUFQUFxdz/HdzYcqQYATA7MH/PSWP8DYBOgAIdeTKy8SKDcia4aKob
lLiXXOwxiEuUxVJnDXCtHHCGAwX/mdWcmPUdHTKIkUt8m/+buQlodeCa09RPkNd2
hUJuxu+6Kpf1fySMMsRDr+ywN9uf69UtCn2rGnpOjDvutMYC++Eh1eUf+/ui5Z96
3gjgFgdeObNmw+bDTtiNysNQKajhsM5vxT/IK1FfD7yUxtvta39YIF28Vi7RjNAk
jatJHAaLC2r3gJ4AA1VaUJMeH4qadMQycl0AeHjBCFx/RfarA+XfzZdnKN+00UrT
RvRO5TB2IEU+009L7yVFBqsKw0qWtnwi5e6Y+kQGRByWuGft6fc828NAZp93daW1
IVTMyjEUtnpLzX1vfmfG8nSTiAUy2SKYyO2EyOZtZPCdSvlvef5OuHrEElQp0FU/
J652SBDcpGb4oIFmEgQt4CqeOJJzg+h1ptfdxnXhjppoSjiJQJ/jj4wY4mQfIi/I
cgcKsCDxrcjWo5EbNMr3+Wvc8vcf5F3QDh6LNT9Yo0D6BtDt8EXhNvd6EF8xiWvf
0T8/kwLbjx4v1xrAXsc2KByApgNIVGrk4F9LX8fCCYUfBSLoJkH2liiQZuLRC+Zj
0ssTAOH/FCa3V0OWb6v7Q+MucmB7CO8EmieKe/Gnso5BqudULhJaaoNhiA0iKyo4
ifoAOAts63lLNvii6q09M76HSMwIpHodPIlDOCF7+IdghJuRkehiqXOWD4I80cO5
QEfHvSL32h9Z4Rq5y/67vyp9hmLdkcADCo6nuFH2h68NV40dTu2g5Re0v8bCgAs1
VoBtecGZzMzU4bphRgNY/oeEwIHy2nQUI/G4EJkUjpqOjFGOcjatoPSbACa5CiVR
A6pSn0wLOP/b/olxA8LIFrTClBodOSYrrIGQx0xDYWoHaHtw5DT2pq43mk7UOUH5
wCOLkT1g3BunA1tJ4FDBJktMaaXXkS6whIqf3Ig48xBLdv4uzbzlcA/qG1TU7pL8
w6z6MMeHQOetUmqnocDqSJja4iSYdpI+wH6jLP4c34iPodKf6yZMBoBSwXWf6/qM
DiCqh6oxD4XruTs0rAn+l5yyJe9TxKF3rnZ537utrqghlTWtTIbgP7whTnTn4XTa
CklCkURZAEuyS50vyfyGWE98fhAVQxejFpAtblwmk694yvlwQqj4nr3DLTlPTuj/
YbAukR6Ig3iz7FL6KDa3o5OQrSjloxQC+8g0i3JfszXlpNC6KS4owYNaXY5rVgCT
ZZ1lOm1IamUwFG4RO7NdMmW2ztDlgJUnkULa3it276Ij+q8sHYXn4yELG9G4SMaN
85ikcX/OYi0l4XYBQVXf5yGsQ0iY8BYlvH8G86bnKAXO5c86Qi06e4FfKp8XZTZV
92a+T7ATABl8x3pIRAvRiDXXFzw1lOCYN1EotAF54+HdwGcVfHoSTnJgDzGdcJ34
+qdVXMyPvyBON7Rr6GgZJCtlLeqH142wJE4whZLazdfdzOHQO4KF2/X2aAKh/t63
7n/JvzVL/4T1Mrk70iT+VHaoiUg2OoOwWyJU9eZSWryQwI18f0QA5QwCA3K3Myu7
M37lAcYK/dZKsBOVnL70SFxgSxgRlabaqsTmtP/iY6M=
`protect END_PROTECTED
