`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dx8zT5TUbljx6+l/nZQNiqqNFad7NaHD2lNLsKp6mm4GRlHYhnsoBY75bBlJ+i5G
6cWKsD0tX8WTATm8vXLNsTOIFev4XWyz5Z2DnRON7GKqphDejhawqJ8Ey84qCu8j
ZMFdQF/s1tqkt4+kctpVErAHEqeFfODbVRMdBybHMQ5Tl/HcVrYpFxAoUkjKbQ1S
MDaE/7g7IXCGiF7XHIPLzW5GZ5V+mYKGiDhjsxdv//0ltQJK/rUXT0XgJrzKIqar
ptc7OrR39cP4gkT4qARWvpjQZAjf6jseujIFNYksRQpNtmk+UboKSOlyEjBuxu6e
GL5aoaeMa9QLpuZL8a441U/EYLP4SKH9DngZOv5ewC985m+w2f6XnExMfyKmy1wY
kKhLLUU6utb5rK0MQTNAF38qf82PDPUG/UChylQcDLeyqXqT7WiiMoWbR0FJCuc7
3PX1rMLNkPHAWajYYWr9nkmXbRAez11xbcEAKb2fwgSFua8ezEYYzGI8yquA+fCH
oOOUtvPQfdOL4lc51LD9XQ==
`protect END_PROTECTED
