`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRTZKXCa7sXexIdcDrPhnV2ekSZPY6KCE5R8Y3ZmzEy8wvAQd3t4HZU50/czEUkX
JWqYdotPOM9EbdwIChxeZoOoAxj/TO5mRIxQTK0LMfXLV6C6WVSMCr0505ZXdMID
bj6+7wYMkr/1it3+Nu53krv2jg4obFkZaXLJrmUJ+ch+fiAdp1m8FRN6I1q0D2+T
Imw/5KDEn03BI7bbXJTqG4w8kULII+1ldRZHjm7VnIcvbz8LDvEslxo4pL1+ApAt
2xxU0qYrqp+Noom5uX9b0EXk7F2eyXUf8pnxXpflQLtUhK25KNUZr2DhC4Ct2aN6
v7bc/+oKIUFTgZoTzpbVC5ap/Utsg/3S7NESoSZn8WH9+b+8i9o1ggBcoPa0Ue8k
MSzrPusfx1k6DDH1TvQo+TkAx1Ovx1EKgf5f5puAvCwlsxUU7r3blvr3FaiVv84t
vknifRKuVAWgRCt3hsjHENQUxmt3DEoP6KGvtP40cjl1x2eNplsXQqg2000+5Tjj
wATh1HUQA4crxjXdo2vLGk0JNhuxwIo3Ze9dyOYHzGsNvAqZwngh9/BtfCTkmm7S
y5GTzuwT0WpMlJtJagnfq6YGWlmi2/B6D68ov5B2JWAWrpN+loR9WkLbTLSIzO85
nRZhhfAxB7JLIzvXNRP7Z69e5yGXIbo+DK8DxxYXP1Du47az4jQ0lreEJA2r2ldX
hlxanm1/1NqIQDp3MMQGTV2uoTYZcp9AQg4hLh6+wBtq/eeQ+JcUxI95UqRKHsNo
hgygnSK7Hswx7Dy2W8vM9g7MSL478R4B5XHyPJfAIqQhq6AJFRM2xT4NL1m9y3p2
GIqYShvmytXPWPVskT566U7NRpKPWyosn/lo06OpwQuSXiK0AjJlEhi/F0Vy3cVM
t6TldjunwdzpA2NPN6gDTlwimPsjvdz5kq7gl7fHdvA=
`protect END_PROTECTED
