`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IALMYG29MwDdebAMz9L5Ca7pmj3+825SDyMbQWrV/N8remOLBZK54nPGeuPVlzUW
IQwZh8UqtzmUNS9ixVrpmH4muBNJxIfpAAclvxEwZv5VIaWIceYUzIdXeYQAJvJM
s8BxaCkKy1A08MF4DDCn+1BMFM2ss1GwgBylAcXysvJb/ZLzw9tmxg+4xno6eYcn
0x/lRrDUa0HdXaAVLZBJlPbdXNB+g/tnOOFipg541yuXh/Th5k2iFKzhxHmO2XXm
fUBIJp+DqgDAxnXcd0rRvBEtUHeIyrYdCvTcxU85WrjYnD5EOmFNMOaLBNezGNPK
4WmpwB+f2yQa9OVqIB9xF272REa45VGglMjxonfGivHA8Zct+oZyftjWRD2z+s2i
CzZZKwo3dV2FETSrU4DbOMDRpz2Hw1W8XtPNuyXp+CBqoRSacXOL9CvCaYq4LIxt
5fcXuL39zPIjZlmxkDQInrSwCQH0rEp3PqnAjGMTf7RijABLdbFn62wbPmkC6X+L
OtDH8w6cJgr5or9Jqb3eVrG1PU2JFVBsS2KspRfm/YRAl0sT2d+ee8MPBTkX8epp
/V72GX6/H4rvFDMC5vB5v8vi/7hY11Yr3B6JMVWJwsFqGUUVGwjedY1fCKIJcDE9
C/IlGw945cgVcPUdqpC1g7P5QrXF6QfiJKowInDOfsdd26bpkpwLEV4A1ftFE+Ax
9llKmfJ43lHFYS5uj2yMK78sf0z2RPoNrNWeGT8G57xUyUs+tcwvfVltTjoj4wfx
9snV5CJCswzDsbA4fvRf45nV9Lp0ThN8JamqKG53P27GGS9TafQaRO1QYMP01j+I
/glUcZE74NA2c767OrkQ3gO5k8MT8vag3vyVVw3/UKkKXkZMFHMLvWTsaqWGz60L
8n330kZWlSGr+Exgax8NQtQg0RtBEpErWF/cUEL60Gk9ete1N50y0ts/7lD6IarJ
CZoL+2L6uEZfMvYQVbhvFgewMcg4GCqoGa0E2KiSmGwi/7/HSan1eg49tAmsHFjV
qebGCLWNYTwqmdcTwFtaEI1nNSWkbIer1W3hTR2x8NBrfJP5Vr2bBzu3Xuk1EcPU
8vOCI5PNj5ZW4VuHKpJCAzMZmw1ArKytIf6Ti+7/CU6QaYFnoNlM5AZRhOhC2SOt
9i9VS/x6E9WpJu1FUHxP+P+lijgTBn8ThTt4cSC7FtmF+MTj8w1FvCzgnejvW+JY
MabTPbBdXd36iR/A0lEE3BIJlbE8eGgABQBkbhGyq0v/FT8VYvDkKpaw1X7Ra9A1
EvrkSzU1/87h+hFLOWzSUMxzd7BOuPRvoFL7WZ9TRsXfNF4sIDbYRRDkhonwUxUL
LTIb1qwFjlLbon/MBperZtpFxt/qmdPYoB/+eu8RaRf7lOA5BIFhxPfs//nxjCv1
l5qqXP5P39y+OBKyg+kSw+IqK+b8Klt/O68/1PqqApTOqHLpEJEfyxeX+yY/Z9Dc
kUmTan8jMtr9v4B0HJV4uWB1C9nd7DdrMw3OTxkzDlbPMYVTRHigILdfi9MS1x0z
p4PnyhEweFmtjP1YwQG9j3vGWujHxGnbeep8weyD8mY1oUGYpmEiesV4Tny74gZT
E23V9OyUs352oE2APMrg1YH8Or7OrOgS4hq4Shqcf7IaXgqtfxcvR0XjH8Smdx67
ZHnIPR3WwX3TUhiQNJXqHWdRHmp664vCXiOULds2QrPvfhIYOo5LHUB+pSieFnpz
3XvTmmGnvfDwjlMoxOaTTF8339eauk5EBFxCHF+1TqS28cqEbGouBFDmTdLVc9od
yxtONoH8qE82VfnpSClxK9QVXaHW8Uc8lqpoo21hq/kH1EYB6ljHUl0cc9VsDEx8
`protect END_PROTECTED
