`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDSUbfrfczyoX5T5etwKF9iexp2qVr9dmNinczWBl4OpQMBJvZ++HcuG3prBEroo
VGB8MD6kH53f5QVPLkzgEuA37+vgYp0qUbrZ/Xlf7QmXObgJrUXeXnt/0XiUAd84
kbc7mJlbIrFYhi23tdMRTRLlIRgwmluRldlGcB0rTo99+CLtNt5GKGjxsbJLGdCa
n5K5ub1JO0NZWegiWdmcBgWZEfaBqrR+5acgrHBeph7eEU1gsERoitlTPxqQeS9Q
dODfm1Ev1G720bHDvYapNQB0UHw4OQKOaBOGKaIJFj7gcKQqFJcY7uoPde/v8rGs
B9Y0Ois2nAPJ/uCCzogabb41XY0kEOWWWHe4CsZeYF5x/UWP/LlO8nyV2IXq843c
ePdLFiBQoj1txxNNoWivU2c+EfdbJiMvMzYntUIckoj5iHGAZqp+NcNNVjGTfYrI
z2vmDhESGhSg7ko87PgEkhkx3Yh/eqZamytxdDrmtHcnYrwniKClWY9Ihj+a0NoD
YaZteu24QdPWxH0kj8YdgYdoD0onUJzfh9iWACoi4h0HsdBqtFddsnwuFSBLIAL/
ymsHjQH40oJB1iBo1btXuykmK4kFdf3kXpI84Lnp+DR5hvYQhGD5BmbUkOX69m5h
/KXfNeStKDJk2/5lMp+AcA8B8xNPrgx/SKN6cepwdLGBqL98ts0VYmDxiargURii
Ih0+MsUL+vBrbATb3hiFivi6htwUmOIi3Exy03alTPbvUqQDtbofdqO+z9DuW4NE
bfBYTRvd56ivHsShvAHr8tp1We31qOeCJqzwD+Jf5Zf1GvC/v38jsvvE0TocDu65
oNxRBs7iVKxZamECvidIlZ4AKZBnptiKWkaOw8KBZFcvxLiXa/oAkn3cbc5TOojw
Jm6iFz8tQUOKdkqGymnd4HIXd6GrgwPkR28HtwTwntVTw5Dj8gDWqc7H3Qt0kq08
ubiZBTJHsf3SRbidSOAPItdRER5B/SPAmGOS4Vsn+RZa/+p40hFHdq/IDVxLe+Xd
wcKxZBeMlE8M8bVZvmNavfGf9meFnGojf8JUME/7+r/HgWHHqRvjWvKsN89HxgBP
3isUvllyrQjOURKLtuQE7MbYP0cbAtZTfYXfn+ifZwX+FajmFKkph2yovFCjBzhb
5HUE5/vSkD2qOfh2rAzyv0smV6vEr7IUz25uBKmBo2hHldwyr7aANz2ah/joduTl
Tlt0ZFKXb6J/c7zyr9eMluwzE8sEy8ZIxSDwIFLjjMlQqjNFPz95xBpV5ljI3Ux2
8hkqUcKB8M3CdKk1Nd/4G6xeAFav0CJqyj/yHNpSnyduQs+7ErpYfWfzko5pS5ai
o91ZvDyfKHgWMUQvWlzb4C2525qPeDiFBMsAxvc7CyDLJr8D4M58aZ36/iV5GKgk
HYfBGi6XaerS56sF+GG3rsC9zHuNOTLyU0i+LZe+v9vfyuEb58ZZsMHMCDPZ72uI
UStZxXx894dRjlJMGn25BA==
`protect END_PROTECTED
