`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m5JWbSPQC2VrpzO7m8YKawJBNkWynr2/HY0aLqKWYxaqr6v8+RskGBAVdNMgbKWz
EgrahxEdfeza6Ld2URiwRwUItWzhKBhLVDniVwRySZAGJzWOevRjp7a6wM9JLj01
1ptMSiepLF9hruW8IB8Q1T/U6oKPycRjOTyNBkgqXE+cZSj3mgl4b8SN8oIEeYcn
bqjPdno9X80LpZWyzbzGNaB7ZAtArS51aux6umkErMq4DnzIc2lxpRvNw5uqQF/m
wzobTeHA55KV2fZWvE3ZcvaurBwC1NcMvqG0aTZN/Z4yJW3e3g1TjlEA8Hppn1Ak
PsCigg3lUwcadMqlwvGpEekbobzf4tnYX7r7IT33zNlkF/MEPgK2jSoFVJg5ZoAG
6BhFEUPXIpg0CmbRPWqsv907WMxDk5Buj4wxNdZ2aAt0HT3pws2NL3TNhOhbk3rY
/4owY1nXh5qluX0ECaMHvcjcbWouxNcwaMZH7UqivWjnTG2B0hqkf5I0NOssduzj
1KHOQ1YWEgayLWRX3uvtoB4y3NJgy+mZDbqrtFAbsv7lrjlVGFZyNYx5BILFEivZ
R02RPvjatSEMKb0tFOxRfM8hPCtvlMx27AjfN4fRBzWkAJhMY8X92YcaECTSmg1J
V3xx9qhuikjjlh6D6bpY39nGNcwUjXUe4hZwwG0BaUc+A14lye6jCa3YDeSO8A+N
fVZhuXmmr15cVgSwj1cOK7pbz9FmlceXQJ1W7lWUoJvsOWjxoUaazjXnJnTzxlKZ
A3uCiSRi0q9M2vpv3dfdj0G6oj6GvJyefiVnm4eMYWVLnhdNcNbd790su3OQddHI
8GFtYUxEW3HBH/Y+eXqvlNWVejJt2ta0U1f2nxxKcmBduTBj4vSyjB8I2lcozggL
fhzUEh88Wi7uZHRc/BWJ7blePCuzyW96BWA7bBHdvibBx2LXXN6el9ZPUGxPPRNh
Z5ib9qUqAnSqBncoagiPywwMjL99MeDAhjo0/rGQnMf4Sbf3Ux83URoOKDhigxIP
H3+mgvrlzKeZNuekWsTx7T5XhkPRJqTP3FABU8P4L4F458XVW2dthv9vOw5gg4M+
IbU4akOsnoGv2dM/WqLEp0UwgM0Tk325o4T5aOtQlN0avOYcGyxiJn8VvoB0kpN2
qyhcVaxjYo4LdCB+Kj45ss/3IxGuSkuOPK98pY2LdCloHMaHsqR492MyBha2961j
zonzrKUugTBgb8sGP98alQ==
`protect END_PROTECTED
