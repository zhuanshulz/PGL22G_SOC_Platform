`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XR4nnEGBaL4z0ap0mURJuk6vb22tM/tUbo2JaR8rsHgDk7AgSUaXwMs+3VvxDbas
2fkjB7mOqjEE5qgPjDXDqW1LnocaiAKtPJNDFsERTe6RxW3SAYXwUB4ASwsztdgb
sV279Tf8zRkyxff7O72fPfRhEhLNBZYSaEquIBOY7efHFqwbovgqE5ciQ/AYS7Eu
A+LecuzA2pbPfGA7M3YDJpFK08GrnMnpMQFPbfbnYZWTEJJHsaEkD88yTXMXs3FV
78rwYF1OW5LwDftfSc7SOs6kgXetXGcUjHt9Wx+uf+/YpeQ4Vax69oJ6TaaTC2JN
Mdhljse1EbcxvhVIdDPAPGQU/k4pe7otTZJtY9wEki/IilJS6302CIaKQ9CleGkJ
zRFg9blXl0ufe0nuLK0bqQExuGoF8GJiMm9MbIZgfhPqb6ZR1arreC171RuUWdSU
wwme+PDpbQ/Bk3KihL0jFoJaVSkkXgAZS4Wy1ZERXUQi149SfL7MUEVxS9nUg2GT
YLXGUdAvO8V12DwgQ6aJ9jhDINSmRaWi2cIVdVn2KuPe/bdKm4k/eFGTnD3Hfz6Q
yTX6QkpkNw0mtU6urg0SNITLbMOthYZ4RYLGLFfGxIZInXDknwu+XNT1U7OFPA77
BEeBZupmhjJUGx+Cmmfb8ZYWeGikGIDvhUw14JUB36XcJne1adHg7TWpa50+A5ax
DKOjiR6c5iVu6r7sJ2I2ABFdFcMAR2+stIIJIFmnpBUIuaWdgbwYKNXNG1OYnZV+
4sDpT3aLIzTJripuwyLTxGHxuiQXptH0mP+DMmu0qIaRAz4Al0ac8ubX8v0ED0d9
gbBDQzvNu5s4xoSXu0Rga9JcR2Iot8gFR1/dXCbRD/TXygyujNCfke4XK9kUcIm+
i39ydJGCd4x34txvvybb+jUVUTMP6pnfe9FkWf7Twfb7gOGfPoCcR29Oa00ZZOYq
k3+KXSph7XiXJgVgfbhsATt78FTTpla+Es0mn5mv4jC0VqKWNYPrT4dBccyEPq1W
CZHyt/s8Rn2G7T+aQzkEvCtrrKOKyJIrxU+/5fxUXMbkjPv3fZ2trXZjNma8RHqf
j/Ja4zTN2D6LdVrM3dhTBJEcx1quyYBchBrDc0F/5WDqmL1PAMzgxkDJSbPHh15W
lZ31uC4/N4FdorTk428uggPBTZUBJeTPMCqNdafAy1gKw/mq0yxOc9pJ2ddGtByN
A4WtvY4JP9ilxEsk4gGfFcJfonrRFIH/YuUNpvi1u7AxN4/x7jQuPslTE1f3x0c/
TZqy/rhUQ2CIyL3uYuP5cQkaEj2odZORM2Va84PIRrLIau+mA9iaMlfphgpXkGnZ
eipPcTFIN8c8I0tPwyAVIWtBjG2BxzHMMp19RBwW3fYBd7ykDlW0pxYYkcahg+BI
/imlpCOHver+1eQmzzyhnx6iBWXl4lwbzt/92OpGTWdBtgT9PQ6vwEXR+PcDHW7P
bLUxkQ+LpauF8EVUw8oN1SZ0kMWmYKtfSP1HAy8ft+O9DUWGv95aVANVvdSROAMa
b/57vxQG6Ic5YSukAVW3ZPPq4I2+moLuNWfQ5YjqjHoRIES0kiwNZFjYIUykZb4q
LbY3Da0uA1M/9WL9tzYttR1XcE65yi5ircPqDHNXOZp+YRp40fEz4MZI8VQuYoUE
KHBMzsjXNxe9ckvyLk5VJzkoNO90MbSBB4FHOwqT0ybFBb6lqeuVge3qet7zeTS2
YiVr09unakuZ9DsUTvFMSWgoItNBt1vBWfNNMPXclwtvxFsa/9VWlII27309THg1
0wlSTO83uoFXXy62819+fh29RV7j92qcz02eL9wrc13KG7v962V+KMJXNElXwXgl
bW/oBTHOwbYcIKOBr990mJFk49aiXtD2GYT6TR8RChKRG7K2wr492hW7fAfubaG4
zY2ORnKo05bixJQFsURpBDN818AIiCezhKJKhTipRnqD/7rDu9uIFqqFvwbyTCUD
5dNNyrjR3O8ngYIDvqT4NH5/Jb59INtti5eJykPZ7+Mdp+GeBdxu1ECGlzWWrvCE
YN5ArASedOevbnJ+Sftz4driVmF7TXfo1h5rmItHvpmzb/7JziB0c3r4dM7atWem
u3IqoAGB9P6rO+QoUFMDlBuQwvc/phMLHKDxuKyPRfCBGKgltQ1j3u0zHWtIN1eL
gbu7WF2ofcKJRMZsZjifhOblWMWNOB2+QAiNHlOKbLJ1eQrqjf+YWcH0w7vgAJp9
tZCMPzgHe6e4vrXiHwsQ25WE/i980SSBhBgB7YP9W7w8fnUnfGF77LQ5kVrIf7iV
fSBaiDUt7RyF5RGNQmELeUIZ9CUvK+ygyOa7BotXdG6EHW2GW3IdGBgZu82yj1RI
19Np9uvjEnQNTVUKzSU2hWhg6iMLGAPnsYdgWCAuRtD+qYDYx+qAGy3TBDORVVYf
DSO2sGfx31DQWNqXOGqd07MNWy+62A4QtbYTsMznwZhyY3q1dp/ql33G35X0O3gB
ANq8+ck+GejQ7M3hFuj/wg==
`protect END_PROTECTED
