`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tM4+P3bHVo6lM6Bx2zHGmKwiINXS+D5I7qPhxOeTcQyuVDrIwkn10vrlPamEtCQ
Gjn2WbWa3Ho0KN8oi4B7rXeoLsvwbEd9f4yM3yz6ynl0psIOFj2UNEDLWZ+zd8eR
w8FvWCkp7MabwJe9jJqqUL8AnruhLFeXjmmjrX208rk5pulnUIUXghJYRYJvLlBX
imbwGWIF/zFwFXy/6rIVEo5M0yamrGYAxfY/2lIkqybHpsGNo8Qu+DAwueE+FgL1
KFfnocLYNg1JcgmIc2/ceZmb1FH08FY5SqsbMm54GXu9As7rH5zt3ekmSVu171p1
/XjW0wL5ED0yHD85cIX6qBEKsvLw0Ium9GTpRMrZvpqJGEkQGYy+Lfyh8G6Bq8Vf
Fj8+pvEwo7e9SI1phepzPXuTTuM8MPLy80H7EBHZW4Gcbims85IrzymczVDry6Ag
tAE8ZL9Qr+8xyYMNa7YPMLZIL06X4eQw6gv5sEFBOgkMpdA+zSRCvzvGwJJ2mvcw
b1R9BlhkNZczUGdLN0YVVZsffxmlSp8masEAt2oteWLiVgzAEpCb8/vKFAubOb5D
xzyOmsMIautSQk0hP0M8GX+Blj9+mBFu0vXfdQLVF/VNE4tdYHr5Jh8SvSuhQ97t
vMSEeWDY4oFaBU5xTIbyN7o+spr2Q/0VYhdqeydkfmrOJNX+KktVt8NvRtxkYFqh
9lDlPbBqVlk2YMgajxizrC5RGa4N9HZfaWPdeWCmizcsCJgyKX/ZnQ6C9Gdbk90L
24lsP+yoa+9fS5ybSJyeFcyiegHOIvOcFb+a7AM9UOZSlLo/p8p6q9N+Lu9+wX1O
rioaYjBPK8lMzheht+js2Xj+726pmVnHqOAl09r1IsgfgePCirZoAz84vxBVTrNQ
7IU7prxZSXWhruL1vHIHMfJ98NJ6cye0J8iuV+5+45MMbuAsKaDOdZurHog+B50D
fqe5YjpxXmmXbkiJAotStK07pptu5ziW42+T+qWNlrUZxDMV9e/j0gpyNwWNpq7f
GxE1Ioky0Yym7zKHH62a3NT/hkkwL8wUZrhftq6SPM75W+ajtbjXT6bFgQn5+Z51
QVdysSTMVl7ffRzxL/tdfZL5csqttalKuhsU+cqT+5vP5CAf0RxM59VjyMLVH1RK
Zy8GxJJq3Aly1b0uEfllBNqFOLSoETSsyNwSZGbe0ubHbwGY6PxAIj/BdPwX956j
o0AvCNmmefvmSdreX4oSJq8d+dvSPw29AGjl3UOWdsuOU/Y/QX2wI/6znnPOkzwI
fyUD/lUti7zDI7QB4M0IQnPIDQQ4+zA563iBgXMkmMyIKgXkfcr2m17HW9BrtjM8
elVK+1LIKawvVKrLaGAw/m/LCPgelbyllP94fm6QahI8RjxTu9HUi3z8+hsVuZdo
2Ais48zyhLsVOkc5HF6gu5htN2gH2kII0ucTVkr80F3TYVfs5DPyfw3R5d4PxMPF
cS2XJzkhd6ZrV6g3OKfekadlW/+xESMUusAAS8OvhgeznBUsaXC7yirUPPu9AVdG
edYNsTHCgKSMY9Jm3lyxsBaA6JXiLE2o9Ln+eKeXu8eI6sIgE4cv6T/ugDdC9K7M
lysOBYPjRqewBiP6aL8JYj+G065hWSk2dgyDQFRR1gEVk231uEDMO+YLcwf0Q+q1
QF7P/5u+NhWq501bIA4GkaTnchr5b+b/18WV2TIMkk65oBdiufi1BnWbzh+9aBNc
VJEa8ULCS4oWMy+dIOmnDlqZLF4fU3eSgjnthW5rz0PPfd4R8jsltFwf1RT1j0aS
0n9i9WwpNEtOR6GiOTi7MqU6o6MxtfYRWDgdceY4tMp0Vp482rZ/I41sJKUlRsk/
6uUYQg1EAENRqJWQiwsNY5Ec6TPv+8wUEBRJ0W5W0jnWAXb2pFct72RKTNA5l6cd
qbyCMWPZuPtBNmFv+LfJs6gI8uSwhmTIolau/Ka6n05f+WfdhceO67tIaqchq81U
nrjW1b77JugPT3HmtMZ50QqZy6n2cS+m08uLnsYpOdZ+Mx06BJ8NgDmIdZLnbFCz
MgBH2UJMDXDmz8aPcjMK5ALF8Kaaur/4uJ+tnWVtMcQwCGExcCITZz1F3M+Kasfq
4KjudLc2ATfJiqfea7Gh5G9MJaFdAxI5rTI6VcGupUHaaYXgExOPL+axvq4TMTsW
nMkW6tqFPobvtBLmJCfxUxDObwC9FbjTSoJY91eY8uprmpUWkXfj344/omzkd96U
POaxQiYUNvZpnhvlrglW9++jyu5wrt29ZMhqNSn+WD477+1y+bRbFtsolwMyN4l9
14XqcJHj3o3T+cG6/4lrU2Fa+xKUa8Y+7d3bKllRP46E3L0qZUSOcCyzxoQw1glD
lZPfsJ86miwMmPOCR1jbDzBPx5FqqHoxs1or6UOLRRMFybbHI9ws/NFQWmYvqRzi
GY9DV6f0/TrWEn7vq7zt45Kmj9DhfL/tabdGVCYiUj+NOAtuuiBt/obX3UKknzq9
4xpA95sBJJQ9opeweW1U6Wva7JtiVU9iBxlRViMB2xqBq5PLSWphDPPuHeXvufxE
ctUX9KaWdX0V3x5x7w8sJJt3IQ0Hi/DlXxUHcZdnoCPdJg9Zq01wEVbebyJcITm0
AiIM9xe8oMsZqQYLYlAZzj6jPrU2bWbzxwu7Ip2Q2ECxLC6D4txdp6axSE8zb6kP
tbetF26OZf4uqvXv2krz3CHidCEsDv8asoYmoB8wAO3Bsl0hB/N0YCKGBVzTLx6+
D9QPsqxwgxieGpg/RMfe777E/JJzO+35PgQ6XzIS1QQRRqiSjzXuGHSFa0DvXtx7
ST/aCgBqITW+BfzMecKw4tii/C0PNE8OYPSAdpBlnwbVmsLc15EzlGLMnZgAUu8n
e4GVWCcdP07NTZToWGcBS88SfiQB4VpMmHPv4f1vSH1RUdcHPKJzfMsRJPjDF5aX
bGH2DMP4HmAzYW1kMSxm4E11+ogEbO2ULGHSrvZD8jwPIFx2DV9BSxwiM6C+lJlE
9LiwULpBJPv8bw/LW3WCJGLXGj9g566++24H1DIKjpTGTnxNZb6E3qB7X4PhyIhy
vhGIuN/JKMw3jp0xMPchNPr1AMwjn07AOfE+z1kfEcQRXdaDwhMiOnwvkoS3aEW2
shOAt2UcXSfmDNmGftXKPh1qcl/DTdpHz7vHdThTi/D8Af825ucUi8669jYFxdmj
2cymFanwYMLF5W7LPsa5JL5RgKZAwVIEF4rw5RNAb6++TmgIoTUKo+858XY8PauE
rjJMNGAif5vhNQSdIsQPxRujGBwZ3nyYqUtDcqHjBX0Ygy/qp2ifzvMEIKk0RihW
TCnc6r9NEYKD6/UZnJcyfowW/H5jMqHI3wGASCrNrfVD+2fSv6cPl/0ovxz+xonQ
hFnpsoBw0BJWdw63DRpU3b1+cqXqrFZvmXB1puh641r8YOInAhSkXrRPlHzKeXeK
j99MREeEOL63WGaaTJ4y+8JTblWzXXoEbVU7FQNU9zQdBdxTxiqGV52QnvRIO/GK
5XGdos2Ne8BBUTnXbFGTlrHHbA/y3ehf2w8kEY6k7pC7yXiNR7zncOg2vpRdMWQu
7poYxirqjgBqUh/CPngWgMjXSmufY14CGyiQ813suiRRvjoSdUuSHZj2EEvAvwfx
AY2TsKtJJtxaG4Uq43jf+8UpD1xy7fkypFXAAvwesACQ3alpL+iLjHaGHOySjCQs
cB6AUWrOaRCnLhkPKEVH/oFurSJGKYb8qhWV6tTgFOMBnFOm7Pra5dMDHA7YKUna
702KEqpAHppW0+IlrZA7IoiYbtUMwLv+ZNfr9qb/TKl01YGhahBjhRpjTdBjukW4
FV7VOGMJT72onziFNEPruq8f1/tHxCGRnhGbA4iw55AZZdrBTBGoOT2LBk0HBppj
F7YP8bDyCMLlsWcaAf3/q5QWQasnO0/N1tzKBpPl13McWwGVflUXhYgqrUP3YLGN
2Sq66sJJO+xakQ+tj1FQQOnBiwd0c0ktPgcHwHER3VJS8/Rgvu9WZPhvnxWNoS31
MSZaz7MdRIYUSyrgz3ib6pgiF+ciDjUbIqv2rMV33hun7J04wYpUstji+kROZru7
eJwdYXceCeEZP0cMC9wv3/wNj8jlJwTq1AZLD4Vv3Bgpd6gr4+JSlOrae9G5fa2A
7YMMcBt89pmYl0CXyRHYt9myl7rf2gGcXHTF6OEB3m5SwuAlHSy+RRIwp1XDO9E9
LMa5cgGEGyRFREjS2VGUHugjsSqd1qZra/rHXB2ZqCbnjhLXpoaDq2dTRIJbDSP5
fVQO7zFlqJxDB7Sq6KhJdSNyMWqOUaT7yfBn9+jpMDe18+C1lpmVpaBa4JUGhwGx
wZy3b12eVBZsGv8mumWneB1s7ZDaNL34xcebhl+LJayQYWYR422q+O8M+9zI+sW7
o5sxZv4Uc2rBscjCxcuLq1jsPR+q0xNiyLf+SM6uAb5C4OV9oqYUYd3sgcFmBMfE
tO0j1rykYwx1l0CPKjZO0IW+2DVMMF8bAkIx5wv8VJD9ZeT53QdpBY6vzhUw8xId
SeUdxMiIrCNPIEq78mw74Gs33DM8fMhalkSee8HUn02NdSFhHXsudohtKRUWSTNW
qtPbajo+i0x3LLNTLyxpzcZqpRc62tR1QSxm+XW/d1/e1nH5yjUIacUvVnGdYMw6
U+uIQKCaV73qWivwPztVaVndxW//SL34uzdVTJ2a+FLlNnv7/o6FmEC4xQIQA12i
1YpXbALd9ViJPlUj9IntPQpd5EslsMBi5QICiRNkRaN1zI2STwmWuLN05FJKC2ji
TcIIh5kCEcWRm5dEB1twAasipys+8LtcN879obr7PW1xfLvyNtuFGqbKgTypEuH8
8DM2H3yZNstMpZV9uBpkhbMVkhKVyjVgIMbU+kO+qKa533rpNlf07wFYf7VW/nQ/
J5e8gn46ysz/K9yW0Hv9mS/PVJF9rgU6muMstFBA82iRqAWPnZ0Id0vNquQxjFPf
IsMOHqZqqrRPYSWlccCm++dMHyDaeMFg7a/DFUZwkqdcmRrK4cXw0AgHOumBpbC0
d7rMduSrsK/lasWYrQJo7OS3c8PFnQOaz43l4p5RBRXBWZkqEbiiwlGUfzkm/Kt7
U4e6i/+4fGZYYhV4xGGytadi9+Rtkl7F1u+pspCvNYPBdSAfsNypQkNWFPF3sfA3
8mM6R8QLocWdaUIoNssMq6iEho/+EoJJuAL91evSR0DLFVW/011RV3IUDzFC7E3P
EpuK6vMbB0PaLVR2uVl89KS8KeLJQiblxGD6cMShQzVuTXmiiDQpzam0e6MPyK9K
R0ovu36sAwqSFJ5dlEd0AHiFy/I8su+UXOB/BIJvXBhYbfjfDgTjyLxS8RBB2mzk
4Wyy9W8Fu8m+KCfMymciK5SbdLRlaBoX0CPE1psBVDkx46NPohAABLfJoqNdzGCq
ZTKIAs8lALPRarxjuXZzJQbl0hiH+DJhPS0YBm0NiYlvkf1Gz+aNQqlCkHIlLw9R
b8+d4n+5fb/n7jGOQsUyliqAnq/zKrCJRR8oXyCg5KU7fj5bjWaXw2OMOT661x+E
BDaX+YMj6LPlpvCWlSlLKJYmZj2it0Un0DcWy2OdcSYYuxxSOb3gdHv+qj7LGtl+
cKvOzg0WE5d6yqfUHgy/JXLSWflBI1dP7ddI8eV14nSb+thkLegeYavSbEXzkwQA
sS4XEPxet5oc9Mnt8aI7yDVzX9Z6mq+LxXpa8wRCFoFkGxw/HfxqufaVo8T8SG0l
H+LNQkZCfXKFQazKiW7FUs3s9A8ZomMA+x6U4KHzShAIqYcZjecIm84ysxR8W5fy
BYawZI/tC0PEtXF7uP2IDcEQ+iJuYOMdZNcW8S5ghETWF9Gk8KEhsiNZ//STqBOg
RO/CuP0m2OEwJ9/mOB1HB2bnPa0ANXXYSwPGsVlS2WFZEuxvwZ530XctKWhvnEVS
V+toQ0iW3t6oWb8Q+DYLw+MTjUIFL4zTk7jDuFOC2YB+/z4hs3TwOcxGHgzDrwBd
nkJ8YnMn/uZO4SuCrsvl5KgQgZNepO0EIRhDuPa+4K0c0IsvrmzSpqwK+Pad1sFb
Qj/710/2Iv0hcS27+RYlPtuWSrF2OcshA6OayvkMcNY=
`protect END_PROTECTED
