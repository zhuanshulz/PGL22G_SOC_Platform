`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KeXOuIbTXRRvp7Gavj85ElqGoop6PFH6No9HPmcwbq/cy47Ue52iyu41+dsfkdpp
kaUnh8ITSL5kCEzSqOx+JDkT7PsblZUO1y5jtP4tnlinDfcoQ6W66eGE2Q8uRZ7u
IF7vrQGPwLgJgGVbTuKkj1FI+iat8EY7NR2a17KdZ//P30rUdeVJEm6ch0mVWOVm
NE8qaeETS7wei/Xweu26MzvQ1rO8D/BgoWK/HBJ1xcZoj8WYzPfkivKIaSYfHkB+
SMA4f1KBMGOpAbYyuA2ia8DBQ/PF4oZKOjheH5xvMZi2nQdt5csTAZV4UqvVmrQH
WhmYAgO+867P6b+mHyCU2ySQhB8liIT14r08BZWQQeCulSRDBV0EY7t4lJyywByA
oJ1r8fAuJkVbQNrBnArUhzhSdYs4zBEQ+TuIFKaSv1oe97Rp6HkFfd+UzNbQdmmU
qVtTKMsRpIo/IL/vh7F/+HWqP2n2dXH9qX5V5aZfImYQOpiNj+/NBJTnGLUVnC7r
qNDlpwFPzQKN4daUSCzu2RAIKaC8/VHW3t9gSRlmOKD4zrOJ2+cukxOUcyt436Dw
hzcN7tZDQfbdyyFJ/e0W8ngjZOTpN3MDduCqMfnCxou0DV+EdCInQ9R80E/1J9q1
qm5r2wPp/Ppqdm07XqywSNzQYHooMGEkiS5MSI0wCOWuMHeZTzKn7GhCkDkchTX7
QycLhu392gDPXSnnZ7eBeMGQboa3ezG8pcbeP7OBbOhXkAHdv0UcnnTdyrZJNkUR
fz4HxpQIpx19xTVa26pfUCgFKTlTn6WHtOishb13mjg6XEqaVRH223u9vb+1/D5q
hxcVMS3WPtAGqSSqDLwDJ+a7p6QDrad4ElwJLQ0Ly701ciaRojieO/SNCdE6qJJy
XD6+LAM1ViZdEuo2LhH9Z97FXiMp+5caLOBNXD2PEGAtSGUNxYzmLwtZSesfLO0p
bAKojmwSSQ9bCive6WRhv2gkxL1bZY1haJy654xWD4QZVui8fZhg+ipnIsxxvx5y
xULyCJ2r11Yu5zPlm0A7z7tza+ZKqgWRKJ+BoXpRmY9DboPH/wUS+rcNWrb7cPmN
s34l8QBqMOHiztkxnrV7G44vpRgr0Ql8QTwb1LFJwDp2wMXp/MFXNwU6b5j6pcw5
YpSe+cy5GgkPq2zHUEiscTavNgXL+XUxQNE87zI5sPPrwdnfUAqaDKXBPelTDy1f
fR3Uc24jVWxPKlvt7P4Oq7NrgtDR0A89iTVf5PWNbxYV4Igfgu4DyDAgtImBOrCn
tVSkoUy6nEG7dsyF+ngmqHrLDBOIrHvB36ZarmUeAM9WRVOVrS4RJzXPrvcPL4cT
Y1LpUx+4wxqZT1L8rzEVx7AaWBopsjBlxs3/jsmfp1Csp81Hrb0CXwf3sxjyaXFR
hTmnzLyOGgCi0YMEpJb4Zgg2KoCUN7WSqenZMpyDCmlniVm+ta/pgMxj2t/CZKLr
mX8adc/4/6pdPEyCkhrxAof8RBfcJk2+fuTbWTA1zgRzgQcR7eZ1F8IkQulZPwhF
1Ci+VIOsDgVkh36vvxARNBi3ZDKuYzBdkuPXAnB3vMyG1tEvx6OspnslYAvVgqdo
dIJA9yMM3wp+ht9i7ESZ+PyK4v5Ba4GZIGDRj8vEila70ZFL6Lp6gsdivO/8D2Bt
WC30mwCD3Oh+l7iXLym9PSHJEYqOZKBOGoY5Ov5cMfR4JEFKyPLhQUmzSbF84DUr
i3jzOypWpGbS+wFYjNHKug32cKV1/AbtEv2gV1vdutPSb1oICFOutmNbSkASU4Di
QhuwnxsalxppewfsZzpabKgVnYdSzUJXx6q3VHrOOEOjKu6T0IMXOWopjZaB68tC
hPsqb+sik19KB1xk2dKZ4hN6tPPIltiikYJVVKvUdty4+X8TDxxK7xs7OAJqugnn
hDiPsmHB0W2NlCFEikHBhOH8HKrMxN62F1EDi9E62bgeW4ObXZjf35b8QREPSMaa
WiL2qoU0WTpJzS6XxJ73lSo+b04SGSCjUvMAWJF5TIh9sUxLZP7WJEp66FgGQVvX
2NlT+icGuByzuVeSXndUL87hY3CosZRPSWeVHXMo9Fsy2Gs0nPtvPpubhnk22BA1
SefZi4Dh7ORYV2mNje4V2idXRfEjUy6Rq/RnB+1HnahlX54FxGs/QHW8FhkP3GTA
baTbL9/xw+TMK1CTEpBznSl/nMpWnxhaNrw/Ow/6zThj5G0x+2v78dOXN6TGy2uy
+WfrQ+7XxPejPgnC5JItzvmPRNnsCzFwAX9LRA/zRCT/UqWrtTzof/kXBBgu6/Ao
tkwodBWSQ+Cbbn3/J1/v4QwUvKicv9Pf7DqSN2JCu39a8wT23+v/1uLsAj0B+kJ5
v7wXflqNqMdxftK8MD6Ol/M4uIgAiX6Ink6+vfcaSwzBfddY4iYXZGu5FJU1CE0+
`protect END_PROTECTED
