`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FMiDYIL7AaK9U5zh72ohm6nU1BYShzjSUEdgrFYzN5hcjUWgSDQFza/E4E8F1bn8
octt29iNI10ajPeUFdKbVRyBJ1dx6bjffFRhE3L55/O3v2DzkVVUw06vPes0GjB3
ZBDx9cqjD5bBs6NlovxHGpHlAZ0j+Z0XSvON8h07j+E8zysCyKm+4tutuDlwfHNO
67mf4TOWIheQGLxriIskkFNZmWIT3ci6STKYXaMWUUAxKY2WbZlbcqTGuoTFS3ij
Puz0UKqpQ14pQlas3BtlzW1ZjATI4ApxAcjekJVMfNOc5TYgazGpLLjIOs6JC74V
bQTZ4jBoQ2kwjwzsua4Dri+3L/CZDVwI2Olsy1CSCdk+jsIfBTeuMLrx8ADfjsWk
9eDkMVFvfVlLLKYv6/Gz0/STqEuSdjnIrX+zxssR1d/CMVTtuobD+dF1CUa/30/9
vVlxccq0Nl3vVcpel84lw6xi9WDUYIkQXbM84ekHmf1NarLkyIiNOLuRJpEntZdb
jmZc8Fp7kKzPcqfykxyD6zoq2rBMDQi+Gk8TkdpXpnQW1ZPgTMQTSNGI3dL11UUM
RPKbnJSRXHjE/tuCruCNtMoA465TEaoCnf6OOaLvhfGGG4Tarj5nFA1gu+fBf3He
VNW92dlzjhZl5CLtMfovf7Ybd5NAacw4N7j1e0LnhZxXcSyQW1su7QZFmcowrczb
s9rcNxqGIKDwoVNZE82BVLUj/z6wdByL39biNok5n5c7ycnI+wBVi+ZjtOiiD4eg
TVBUrLwWiNQJE795hXZQoI/v3j/V0sCjRetfW8riYsL5x5mPJp5l/0S1IRY/SnaM
`protect END_PROTECTED
