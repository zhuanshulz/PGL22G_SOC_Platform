`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5DuDkIK4YNiZBETk2R1w/y3lboP6kGbCS+qH1ID9k+ejqZ3/Ahap3rw0fzao6fxJ
LR9I2kdXlB6077eAJjwHbmruCq5RGrBaKyqBpN+JzA3xszKPPHrq5ImDb58BXXU3
ee/VRRG9V1IhlMsSeaUA5nPzAXulEQh49RAdrjfCPj1IQ5VSsx5w6xv0ZtZdkhiy
OYCeLKLYYBldktM4+q4yt9iloTPF6h69H+qj+lueHFXPFMVldrmyJkoInyRpvTH2
/o3yrlu4+W3e5fRpUhjthxySPZe9YiLe9IYJZDqQ8gSutxyCAf1hNvM/kf0kCVr4
VIWA4qII0aVXwWqLFwIqayKdpyD4M7UJeFdMXaoJaCCbjn3WMjnqqJgKATA3D6J8
g5qyBPnjwKtQJYjxUmiaGJGuUFetqKvRfPeNjaMqM44WpPa1GykQ5lbeukhiTZkU
Zi4u0OuCrVJjESn64l76KLm80qcX3UVHXab/e8MIaL2svbsr3LFfZ5LSKjYnJkM6
51XRW08S6CDxr49AlSIQdA==
`protect END_PROTECTED
