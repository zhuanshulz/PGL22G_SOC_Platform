library verilog;
use verilog.vl_types.all;
entity V_GRS is
    port(
        GRS_N           : in     vl_logic
    );
end V_GRS;
