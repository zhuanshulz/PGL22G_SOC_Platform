`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vuG5lz7jZCTXdJT+o6qWUzLcM1gZIzpeUmZlugmq2OBPGw3WXqNYSfvtz3JstlQ
zCQCT5cSv3owQA+yvIh8KIbaCYzirktg8H77halndx8OJbBTOT+jBIs2dhVQqGW3
vXsIsBDZ0TcXqfy7XOjWDw1FnzedVirNtGe7BcZBE0CmXrs7qX61cDIQGHrONd1J
K6/Z6m0Gpxk/QICGkEK424X7qz0rjpaBoKDjUcThlU0G0NF2B7UdkyjlLkVSl+KW
hzQrJH/EuRssmoOAVM+UKS2+Oh1Kj9ttWrzRppnZ1ohwunOnOhBXxtTPzfzUkIpw
1zZGY7p70cycg35f5b2enjQTbyLDv2cLTiX4mRrVE21AhkMG9Zz8rXSitn/rdRkW
J+IDDPS025DdvaWLytB7ZovxU1ybU8xFOyZBsqwciFka0vT6x0wzSSIZD5d72qcs
cRZpLOuJZpi57flIpOsAeOksAdLtUBhtxRhA1Ii2ysn6HYGj0qwGezmUA+ZwrLsK
2s+I4LHl0l2uHD1WoBiTFMQHxEj4RedAxn2hFgTayfWYK26SwXpUtCKmPVVfl9t0
r7Snlg1xxk7qrhj165cGuWc226YgycHCZMdzqNoaDUztQ8DSvIT4EtdL5g9sOSEL
JASbTlXH0ak/DuWgvgAPLbcprMVqCqcStA+IbOCooHr/2BjDe1dZHNjKga8N+imr
/e5aY6b11aryKI65XredcDu38nVeC7u0U9u+aYNrYN2LQAbCn18SfwSzd+EhgdE1
72Mq+hdP49le+nJL/ehlQJI3gWRRl3KTpciTFVPuPm6NBIlZVDO/a0krpiigRCwE
kuIBtP1QfF471FO1gNrNT/VdKZGrWzRmBzjfr5dzcxEWGsR8IlXLBZM92n/Kiu6i
H2hGynBGloCTJjRI11aaVr5c510p/86Vn8wxXyINzJOWW8NEnOs7Nkgjv3ZYQHVS
YApcxacVzDCtcFgDWtO0FxjQu6zn6rKzzW8vpj4zFsUYQLoKlcKn+Ijo33RAQ7Lv
gjNWXmUXG7FDXeTtsGYxa3nKWpsMsvafFPOZBgNMOhC/Uod9aW2CQeKoPGcbZvRV
r8I+uOcbu8YMGRONpJMSU2++TIKvJXxcPPEnheSw+jq4IbHMstqOGscAWze+NkLY
qEQK6Ir/600sOVV4WRJI0c5qd9JF/ZyZ0mSneAtg28tK81kZmEIeeck5ySEwUZ3s
QX8z+exaQPuC18Uud17TXfZKZNMcsP8pcdC1y5BoOApOWligz7oozLq/itkLHSL8
HvzUylMILkqvNn/aNPtUMyClXbsA1HHZx/vcLL1hibQh9kPZGbmypeOyWhnL+eHU
ITpDP2PHPKHrCTs796gBpVXYUjfNwXVWNp6ncn4o8Ep6Ek7gXAti34getTmvIicc
qX/yahUyQyGmhcolM6im6qH6Hr7oKXJAsY6bBqSIvEqJh+yWPNCs/Y66XO5MsINQ
y2Cy5rk+R5yeTncrA6syI3fOS+cAvjZsMavogfLBG83P9A7i/bSapeV3MRS/k+lv
8XyMq0HIslP47phom9jY5hZ67q8uzEd2R3ZqTfNkuGkXGRBJnSoOkpbK2vA3jaXn
HuDV+B2gFGP0mxM1/QJ6ayh+M4r9op5CAynd+Lc/WOwsDqS6guIE8NQb01heDMqY
kXsF4+IikeULzwVpel/FoIDOy0qeFoQIoFAqf5pKdNaHd8rfCdBHJqj61MPxycma
yZdglpEQf86p6821gXcP9Da2V1Cqj6Uqp21REWrmMzYKYgnwYJurNRnhdJK408xZ
ldB5Kc3clVhp+Q3WMX98+oTk9ICGyVdYO2H3l6HCFGRGCQpHjAXxNU/kIz0ZaItW
Dgv2VltjWI9o9cpzUfVT0v5JOjwm6JDxzJy/wKMSoPevoWy8QFm2REbK3f/B2SHm
OQK7ABK1Qf4UcLiGOv4QpBCRLmjsuny8p7WTNCSge+enP312hKv8ZHq1LbuA6LP6
bRy9iO5tDz3pDsnZm+nWHcwt5D2iirvCzSouJxkegk1KLI38B6n+dULiwzWzFgue
OybzY+jgnBIEvaBWKPJM3b90qaPwbHHXuUi7APfecH/GLYvAGHjcB5+sCeUHh24U
9S0kgRoICvuJfb1d9ZREY6MGyLL8F2NoHCkkzRAQFNE/t2DHKnkpekQbD7N8HFue
ODbkwgYcmuE8hiTK3EnudmPs+M8YifGs0QMRecGwcW73K9ohZpPn0lyk06MLZw/+
qVesSsQZxMGVrr57RrzJB+LY9MVRErsW2bjvZS6KOLSuWYDTGVw3CK0IOyJbIWMi
4gGgfa7YAtWTtTYpxfkOb34zWQzoCYH4UkDkORAu2aG/QJP8ABCUx0n666DLmsuw
MtbPgXJUVhjResGSchClE+KQztEu2VO2tP45gZSOH+MOYeWPuipRhpcTVYCCL2m/
bIeiTwqjyMnZpqERHkSkn0Pw5fURPqlq500fmw6meM+d9DREM+c5VLBm7aAuYSjG
fbZVaA+3OzfBDW+l+y5YrRrLnyYtPQ65XE6gv/IaxLY+mTi7xW+B1J/jp/Mb5OT8
es0xoYz1s//beJohBaADf0P7yYxMS1NFl6J4hdmSXfMo7z/ENxqMGIxFOhY41Noi
KmtI/arxYnw7RoR+F/Wp3TUxf5zgzbK9cYXPPsGl89jaVDLKGi5Z/98A60m8SBhM
DvqJVdIadi8E/y9m6+VnS9m8Vd+zGoL9CTQqE0weeTmEZ6yE5OyQoIco6PDfh7Lj
PcKVNzdNShzaNy+ssRBZnLWq0w9pAC/SkCqel1/a5H5XOkpK5eK3a5Nd8HXyGUYq
YXIvQvmHvKCqobneRIZ+h/RFvJuxzDDoivs7L1FdfoPgNUE5nPGqoQxtdfeVegaf
sPPcEAynu4k7G8ERzEls+4A/ip3gK3VNOie4diBReOdvRBrZh+j6ps2zEdv7yLHf
mKpIpegmKxHWcjufG6rrEkKt9M2+NLOAihI9kKnTeKF9pf5eI2pwQoVgDOOS2Eqh
DnqCcAotVnbzd0xOy6K4mSH4KFDC1+5G5Mo7tRj7w7rab19ojwUhd+3lNmpSo7I4
Ub8ZIZ4SFiEnEXSnLFddprFpB+A7KId5BA1FxMmT9xHRtrch9eh1Ii4rvvvcDBfk
5plbxNn5WvaD1n2u4keTi+XcVRWoYZXvJG0ytVJ0T+CTCsNHJkX/GWLHYeZdSY7h
Jv7470l0tizpNRbtKm9Cj/msTzNeWjfvOnXB6+eHCEsY2/w4URH3RvXK2RReBy6P
i3hwp/AaWs//8fIzsRjVAyPyokIe1Uze/EqWwFt3bTkJx2CfqenqoSPcJhV37ce7
scW958ySZZE1k37iq6ZjLRpseCeuBM/KVp9obP2KBihM6QAkhxKaPalQhIKUNv0Z
lGRiXx4aC5KwhJGbOWLp0X6Sq/f7bP+Nth2+d6cBIGsHMjw4nyqofEc4/KG5ykRU
wB5Txbd17ZAQtuGeqCUrETywtyWWtwFNpeTU7FPtSPDHxtuMAlk3csf9HsIVv3cz
ZGoE6FN9LBJ/Xe77WqePSEVn6AsMeUpM0Ii+ZgxrMUj2kfX/texmWmS2RCBn9M6Y
zwGKydVArdf0fL7U8LpsTIQ036MWrppjyUaltRWDnsqCbuhM5TBribpSMyBReu63
ZkNzqM+1GtBm+uXupkcWCid7Px+4Kryz96Eu6xUwTeNnOhAPZHKyYXkgBUSAI5gZ
EPh9CkvBUjHIxH5FAE/5pk62TPercRM0ZYj5tcXq5ZA1lwvwtaIorw/nDvfv0m3n
AjOUXtMUo1urDdqfMQoo+MxMNwKOnYuS3JvzgWDdY+QUkY33eR0jxtLdV+GxeCc1
ozMUViPbKWcpaAOpiGy9ScIksM7b8HankX6bgaIw3gqnV2P2/g5ZFISm2u0j1Hbb
tOw5V1S7q2WMCBzu2TksPX74W9PIoiWPRWeulYCVLyz3FatuKkXp/Pa3nMot3rsm
+syVo1gU+VrCp3qU2QyoVWWOr7YCwwaDfXGgt6mrv04=
`protect END_PROTECTED
