`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNntkTemUzFLhQd53u7a5k9N/pI5CMwuGCezmS/A2pQquSYf4FOF7CK/nDYbsnw+
NFXLSvTcd/HMliNsxaFvKrA4HVUBsQpPfnvumgkpT1/2DR7DHoe01J5VqcskKVQB
ALmi4WTqRunh7rYxP2gTq4LEiNhwlbk1jyXT46iJb5MCgO8cTLNKGM5hdk6mMrlj
bagtNjZBpdYGXGKvZJJcdECgv+4Krs09GUZUGta2Ujdat6ppMuGuqiId+E/HCws/
3bhWObF53i80QC++SWWTUOrFkGYL+EzQrbvSHC/MZlRYOXxZeeWyrZTk/TYEoLWT
39jsBHnkX0PMoSxFcQ6BJnETwB3gydj5txpTbjRDJoMyVBvx0n1X9kxMHmDu250I
/CICe8RK8eY5CPQ8nmcT0EejEVwe+Kq56J9PnzA5n6Wm22zWSME4wNW6BO80bwZX
A36LGbT9udnYAE+0CaUCYgLeEdyL/QQ48EYorpL+RjpSHgxopvuxWxxIfbGtj+PO
9h9I4opiQNebrDZqw52K2D+92dez4iVvC8ZZ65dEwPgZlQN04YRUD20DODR1WWpW
tipGVmvzofeTSDo/OivSTyj8zdNBuw6bVv4lj+ylwXLqugARSND9N3gNK+pGlFrh
xI6YZeXzGShoKK5oSd/twu5G4rMYQesIjH8GcJrI5huF3UFjNXi9RUbyHYiPGt2A
ljTosfAtWSCPbWlCkaC/6hASg828fcIdA+cml3+8WXiOYO3FnmeWxA3Llg3MjDCd
FtuziQ838D+h1jU8Zq2JDKcpqyHXi1+2vMVNBSmBT/erXaeUbjRhR1BNmk+ZULCf
VhMuAZBKxASH1Uh6yNAEg5gpME+Tp65NhGrFRjjOJoLDdNKXwxqSxyEnWZ9IVivc
lYOY13rp6VSKYreAS5T88EGCyLGtOiI2JwFmQE7K+5HSb3lQibq1rvWaixEKrGND
Sg7v5DtxHDmi1+7gNJhjrBeRDOC12j7+6G2eo0gu3jdYf7e6O8Npyl9R0RtnVhu7
4IPt3+TJiMLaA25IS5eogdn1gcbJZWZVMWQEb1u9puaXwjSD9Apoopm9QC8uWEhm
AS1slTAelXLDGATdKUXp09Tq7XKDXon83SY+lJJJELT12VDgMJnEZafggjMcwo48
gAlPIiu4ndubkgQ4kUsS2jHGhgJxGBjbglXorQmrGGl4LV+yCAsOmQ1JzpNVhaIw
c+MHRnK2WHzQ6RgNr1Fkw4NvCL8AdIj8FIMlRLO1Xkyvz8AMpCyyPzozxLD8NbX2
ZK/zGqwdvKBZs44no4epVAxBphbM81NW493zEtQ1PjCDJQxEPQPuz1rLfJ36QhWU
X/yJKeCccbMTcfAXzTEzy4/lSMe1SrcczfR3XGhSPxKmZk0c13+OeLajGIGhvlXH
tnxzgGkzKsjiJlSteDQtTknSeDJO//NLex4vMRrSuZ3+UibjSSm1RssHF5G2pqFB
JDcrua9rWtIFDEV1HD9Wn7tyCWD3MLXzG9Zac6EUHLJcMJUjgPGLKgIMtKEmHY25
E1dFShcwRNQMjB9/5cnF728xz0h9kZbr/e/pCQWsbX8sZTwhtFPw13kzsYZKBJug
MhvGZNUIwUSximpRC2xWsaPiF4LnHT0SubkrqfhpnkDgg80cLU3KPRw0WoZuwV+Y
A5XfukgfTCywLeBF+8QXK+psBL3vqZzJbGe0ps0m+axOCOjLNjpKSsjWw9HEcALQ
iR/Je/QQvl419siSZiIsFQNBdvsYRpPeKuZdRErKJzj7hLYQOFL9UnKnLaPxAFax
70dIWcTCUzYK97Ia2tCluEoDdJY5LY93rEyIAk2nbnHByCMDvuL7Tt1LTQiDymBm
BZc+ckWsCTb/LUEeccl9BRb9WZnIFX8N6bUNkJuVh9Ub9RM4R97Yw0tBMh08hppo
k9B1tx5eCiM3JpqN4tVYy0w1YP5eVE/MBeNupTaKpX11VSDuGPhL5CG+jeYbIYna
h9MN/JuHgibMXYrhv6C/QJrwBVLFUv850w+3dkejx+RicS/kUFQVQx5IWe4U/IE5
NEoQdeqxn8i+uI5Qm1dBhhB409Tt9KRKk4c1RGtv+VRTRs7TS13TE/63KZoZCljI
K832R+WUwHEHd2dNQ9JMmQqK+gaf5YQlXagZYn7nHOs1pRPn/4yR0efXTuOarJq6
2VJHWZL61J8Dr4gl38tiMmz4JioueYaiZ9FbVFznHPqw9Ucv1BN/nh0b2YHxG+mt
7J/Xjl5UTt544OURR5IRR7HQaYyMIrRc4WFNnYnhSqv2mIOTQ0qI7H5iVkHbk1Iw
/ZSXyix/jdeVx5fg7PnTSmArwJM2lZhSGm9lQifRROR6YFr+oztuL7tbtSI3cSTM
V8mNwE9fhYAkeTQYs3YdQyJttQvlz5jehBBHzyw0M2MvPH04m3Yc7gPkiY2XU5MC
fwo/Y8Bniov9/oAtbuPjATAO5mgURV4pcfPdZCN+jxdVw5wuKIfbuWL9Cg0+OkYC
E09hIK2sF65nsBKYK8no02J7DUTOKC2pfb8njOE9Yqr5byMeZ8FennJyICRZiB0N
ECZEaN++pHpvG4fi/4RkORambySwIUz1cn5Pk9RHG1lcn9O3b2v/cCRj3Lq2YWxc
C7p3/zTazb4RNW4esCH204j6txs7JQw1pHpTZEM4a+ZnXtyFyLyu0P0UQA6zq/d9
9hkVY8m+X09oRwWJ0Ds9H2OL5Re13HKDZ04p7aUudExy+qrcVjl8pUjhMnnPwZjF
O+FcAYQSxdMO6uXAoo2P7rUOWW6HAQ8EzPdICFgGarpjrvFE0lfzboBzoh142H9z
ApAKH+6Tz3dCD3to+SJ5LdkZp7ayyz+E7ihMrHWYCKnHmQyiI3GkD4pGMf9ioQgG
eL/LAr8gx8QAh60QhaeNx/VSZox6JtfZeMHViCLkJ7zD58N0IUC3DpTB0sOGjDCt
zBpPvJ44PH0/r9HWCcrkjklY0wOn19GJcBOymCxuuEUvSbzjPJGQoXL5OtYYSeT/
HYKR0YaZVAuUSRS+94VfC1fNSEqbSHQbhtwTZY5rahe4DeFCjQitxF8YJfdfiff0
44kunN0W9MOg5hbSJHo3vKPZ4UUpW9IzsQVqFr2GGOAkNhY1uSkFwWtOj63tUQ+O
nNKD0qBxfBxCTVZEEBl1+6lWp8/VoOZTV6NLrtu4uz514Y1IEZHBIXAkXG0goJIq
hpSaMyU/X6ssaefjhsYpSMjbW0aiX6VJDWTnD8czRkx40CngCd8eLfIkUH6h5d6m
HaHk3hmP5+/7gWkKXyQp2ThBPur5aBftuSHnU9H+nG3/n/KHCw6BxrRzGOIbjdw5
xY7iT8DVYCz+vy15AXvp67i/u72Vexga8VYy90rTe6tGMGmUeKzeXTv+DSBHonPi
IJ3U9HfG2vD1tcx/Et7rmjLBzuzUmPvirmXHjRO1/uKIs3WAxs6Abn0dbRS/vC6w
GYBsbtWSzo+gyrnlumA6TGH5o3L1NrGBtPlCzgQsC5RLY02U4rMJv2zrM7GlevMW
xfFyfOnva7syXSPoSWM1jK8Qxy/MNs2VyWPBJu6nK3x43gshxtHAMaPS7PZJIP1P
+bEsaPMIGqk3VaXeACR/qlkDP1d1126HQMgjVKzYDiQvvMMfG+L8dJXelEPnUT2y
EmV+IX2MhWOnSIj8eT3u0mWfdchlts7DuzsEIBeTM3Y9je0qyn0eWMzoKWBKcSON
6EeMPwqBCYb/RjUfb6fOxLmN5gaAJUeSfNoIyUNNOhB27+DVinZWu+QNnMDH5zOi
ILH/8CKcGq4WPKQ2cVmiyeVieugia8fMQXrIuAACwlFcAR2+FC9rzMTuJ67fD60M
rOXGoO6SE5oCAI1chuLPXHJUirPiCSJWbPjrZCNJ76c=
`protect END_PROTECTED
