`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DG+zyeMT2wzDGPlTTWOCmKtLbKXLguTcvV8BkpN1Cf6i9v6DkAgEY0D/M+5VG0Bb
yJyYGw6Cga/YrW0IeTnQV6IE0ggapFFrukT+p+ViOeHxy4cpwkRoOkgriVbB+sql
FrIy8HCoWS87vV5S6AjOPVq7F1t4rytzN4khg2aIilAqyi+S3XLHWAGkUiP1cT1C
A+8VI/OcH9hsat/NY2LBnbeWMicdT1mr6Xv6f2TWhvDkTkxQm1szqZWT67qogR4J
9sUbRWL42J1X/jZARg2YFp04KovSbUBpHVoAMhLkEVd156Gm2fZ6F9P498F6k/Pb
19vDsYZSWLEoQt1eByukfpb1+gn+1TuatQAJ8w4SREtkO8V/satsuSfri2P1mcXz
uPz70YgYsf3TRCJR2LOIWR+PoCXjJSlh1+DPpS+cEs9tHpLPZxLAqqZiF/aI9bq5
VUzOwUz/5FQfaBfrBOODgIX9av3aiEiAMMTvTGmOdQfH//oi8oVwOTqEoVsuRMjo
9CJs/5EGRfhQZdiPOiDhB5xQtWp2j/5dA7Gfk0ZqG2SdWvg+Y9IGKOCE00Gqmsq2
AqiawOEQ5MQ58Fuy6q3irN0faekxsGr/Om7slezOHJDOt4yoAWH+XcpW6BHG1ZvW
cvIqKUlvC9Xn7OIvdxK0pVY5b/DVUa9+qttEhS9LiE9g3MSxN3JW9Yj9QoZbfx5d
7WgjbHIFYnBOppkJVRUNhnevVo7znJteu4ZoCQz77B4lZfOmzDQonJEyw+aMfqBm
qq1cgPP/i+zHGhEIN6r119dS/WSgEPUi9/opt/hEnUbEbR4JmyhhmIphI3GrIiRe
M1m+bf6NYwweJGsK+nTa4+fVhwhRv2LBhRLlDKU/REz3Lw5811o47mmed8kYQY4j
/W+F/Htt7CPK77U8PQoE1A1R8FihcyBi+keJR1CjXzM+vdjJ+MW3uZGaXBb4YILi
ZroVlP+hAzMa4INAImE9Gw==
`protect END_PROTECTED
