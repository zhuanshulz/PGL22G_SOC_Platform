`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JgPGqpAlE1Qy/EBTsIQbr+vnCC2KAv98TCloykGmkeIBwSjeEzQnKzIdMKgxVM6R
Yz8+iYV5ynjg+4zg8V7K5kkqPcJLRRlhv581Lon5t+Jabi6iALrnuCL9hWraFmMB
tU2qi9K1dh/y0Yz74Htmx/ETYluske7lNzWbzaqmb70qIzpr/95M99cgP0S+iAef
DFvFI7OFpw39mT3IzCC2oit3jkd7gQc7qo7Mz++t25mAc9IX4K4sVElYclUo27AX
YF5VlXOcTie0d9hJnMm502n1DTfptPxjz8ILgTVIRBKoAtDH1b/jXou7GW+VHTF4
cLMwFxr/Sm252ApJut8Za5yowScz1cQi30frS6ospwSRPidikhbd+QAU+xoTlyZX
eFjlIbaTIIyNUWI17b1oqYo+6wrSUwnypwIyllpHQ5VB3B6VlYPpVDrO5C04dtR0
4r/Fa5RaRCNsKWiR3151HlyaHYwX8uaaWP/IrMtwrYMsL7f0Pe8tjgQLIlRyOL4r
I+VSOVirwTtyuN9PZI7V95Txp8igDljGW1dTjOUkC0DgJrDtAr+fuRlF5a/sxZeO
4NZm8pGpWj3iTzCnm7ZbgCZlMtBvpk31AzQ9rZ1KM+RzvK2+loYvPVVZyHALfXvc
c6+yWsIxDWI2xza4rrMG0C/BaxKWJDUWkuqwIRH1KShNtziEB8095b3djB5Wivoc
Z20yCESE8jYvkP8yZF/2lrFb86/xitwXpi4vjwL8kVc0EC/cyLoRS3OL23EFtFI3
9PMMBR1YltvuBhzduMRtR6xwzPSlcEHQVDWDBK7rZ3O3p6JiO4Tg9bUEXXGm7XXu
nHb4CGsG4gs6ZeCUEbyVL/FC9qoyR455/HoMlyKeTM1i/Dt7cBbca9hLtupy+UFe
NnqfQo/Qhm297dvDtUOVI9zvoQchVuggkFolcLBbsxuLrnNw5cbUnhCQD3+qXwft
dQbbiow5uFXcQHl+99FmN7u3vueiEqX2nkyTOn/SFpeqmsSBTdYIYHtme3O3DZ1x
kBT+hrzAp4iM4AD1YD1uo7qdui2lphf644JU69fafyHt/UfLHxZITayzHqZ7wNJ7
PCp3s9rrgueZieY+HsqBwDD7H13XJV1hXY4dtXAfIU8VlYmAbW4VmZ0vAP9ZHoBq
KaVbn6JF+EkWUrhsllqM8V4Grvtpxnmnj1kU7KdUU/6pvkk19sI5gM+wFd9a9JLz
zqL9R5Y/U2xQV965x0/ag9qdyPRanR1+ArHmvqN5+xXR0Q7XM+6Q9KVWdJYb8s4K
PejJW5gm6eLDRfIxiuzfGtv0wHpfxtk5daA6KMAIZFLT3j9Sy7JHVeF7eASaoDFM
fFcoSJ+VxXLQJwT8hra/8bGRwBKDXrCtfc7/HZ2hmUaPqdQFRVJ3LTtDwXFN4XeS
4wPoHaF5bX7YK7YPQ+HnsKJ9g+njfgdiN81M+OGGvggp6nwj8edebRZWulkbTL+3
FINdYsXUZK+Yc4WYmXMx4Skd2HRhc6ElzSmShJtufHOVo4v589xxGkel6DA1VT8T
nDFHjxss5nJ/eqCjhcMYuqwiw47J2Hcv4Rm0aTIbssO/3CUuA9H7FpQtb0+ccC+d
qgwRdp2LPIJinY7a2Ru2Nufb/I+gRRUfW1c5STpaPMP0Zfi9m8ptMN7gd7dSjuLg
4czDOKQYTfguZvVeS5hx40lqFliVxrggM6wKw+HsMzChRb+V3jxdxvxu7uuwFZKy
/ut1LYNTva7yQSRcrA/Z/Evr2bX3fUmEUqwvOUy65hn44rgjlORZypcLD8OdJoMe
Dd1vLDsJwvubbci7smdphMz9WsCxjeduYNmKOO18aySX6pTKXk/FBrLIB+QEzNEn
YRbw0qYhAq1O8QFgkNFeLG2sfn2Fm4Yy010IlXelWb6i9v22/r2YoOr+VuwEcMSP
NYMgQlvYfcIm8N05lU2k8AWMwzkRmaWQAKGwWSaAdc3a6ZWuE8U4WuSoD9X21F3g
rcknO7wxg9TZ/LplRbjSfMN9ieFvAa6lM2FiliwLkgB9+EomfA6KmJIodcBltk03
deClphZ7NaNa3jjxTa3I2jc/sf9CHy2/u52jiju9bUlxhLKwacXAK73ujkyvSJ06
d22Wq2nn/dEtdNXtl3ST/AsZSQeyeh1y9NPdkGGiR86hL3tQcfmBWogIPty2MYho
AKerfwFxoZOHW4kh2RpsVHAahPGVAfMgP+GJJYXuowcTg60W9wTHkg3TVzCYyHUI
nkG/gU3QLyjOLKBFiGpSi2lCUKDNPLN5NusKxjhip46nDrJmy+7Y8aTZFy4YKTt6
AC3j70PgViN7OaLpCPINM/O+Xw9p5Ru4cm32zokcGvY1nbFOCfsMMI22EHiy7f+j
kewiz495wRllls9Oj0oIEu5Q1NO+khlInSjespAPbcK1OOHMo3HM/vT/6hEOl5WR
fUDqDcMTu0CX+slh7C7NNEYhJnH1eAUVfCxcxntn8hdioNYIboVEB34vIUdGe0FU
8NeZf+rmEUME0XGEepJfWk6OIq8u7DVAONxTzoI3DTHLexJNFN0yiRpiAvdpwkEv
tnhPIbTmgEX+kxZDfFqjhHcVyyxxXdC4iD/53/27eYQURiNKM/Uq5wp7BVLlUO7U
ovs1WdeMdLasj+W+MUtiRiMdNOHy5G1iUFCCyRn4coNiCOaulmWn/J/+t5TjGA5t
HTPUdq31MKPRKVyvU49nSF3y0RIvHy7TypdHYZKz+gLS556s2+vDo314C4yu0EpO
KOT9XO6Xtc7yo3s4Mq5Fobllr9NNnKY1cJrLtQeBNcdc4K6BX5RQBYOTQNs8SgDf
vCkxCCN15w5WhjZHSLneR0S51Ip0af1Xp0LoP8wQ0Wjbj4gnvh7qSNJYVE65tgBF
WbhQG/x1CAuSYcubF6qmDK+CRfQWNpUVzS9zu1lsTVMACu+3dnh4LFUhTNT8ejqg
gJ+5eF0k4QPTFRjOKNx/GXvNyyX6DSbcjWBR0lqzCW0F4JdqVtzMgxwYQL79ltQK
H3NylThDPmz34c3o1XTWfAYv32y+6lSmglYJN2gTXoSeg1No+DiFaorShNHJqAmq
1D/PsSutFSsaQ86HKXBHfKF7s7ooIf0/OJVecsqud2+pLysIYsYMyDQiImFxc4Fs
/o68lak0542Z2FPJ0jSZXgu+IktR0OblWSfKuE8pU1jQwwfMw/onf0nH0If0fiE6
mqpHwDB4mZ5mD62VQRmuX0uk9lbW4VO+c4r69OkL6E5lv4fxZmQIlFQOfGm2GJxF
VO5g3PZxJRuxF5ZBkRAnX4qOC2q8prcI9EyYd+OT76MEb/jmKYEnL5yCTH+swYFu
gldvQLGl0nrfLarl96mlXF3xtuO2rgzHQam1wMJ9CYXRS7onruMhkKESjTO7bz4D
fNgfHK2tD6YSEcimsW1l56xMzT7NoMGHf/zvs6PUeXUKLvYcq6OLgahH/GoGEXOk
nWRmrh2wnBmEA0/hbRJzbL0NpFStCbvae0ybez1F2Rtf2cSkDBapV5KKt2NMuaQL
1jkkCN18EZDMJ2eRRwMMXcsvQjYsi+OHI0YnjPIvAj4aRp9dG/RNYqd9Po8rCWLh
f/iH2cOCzQ3r9DBkKZSfqEvqYdTME3Ee2LDcM9Hm/VEM8XfmTFsiuAdAFPVVkkvf
NOxeDXTDXfr7PHh18VYkPX2SLuUYHVsPHvsxg/GPkpzzsge2Cefzya9Nx5Lpa1+j
fOZa0ljWuxp0ob+zcFMUIm/VwCkoFOJUUBxSv4MNsfd5WKGuFBtpAG7NzmGH2pdF
+GhkLEXHSMrVwLgtuyuGYbSdILC+zix6oW6Rtd9c2DIFr6+jo3Mh6ikrFhryh5/1
a881J5tS/8YBjk7q73s6K1QAOFYSV8CoGhDmSqK0wtWyFR4LAFXA0RjUu9XOMxFy
LAtsVUSA4TOj14tq97J/AGscgMfevWpvCk4RfLgrsk7B235KV4MftVr4RBZmqQ9D
gR61r0jtJP5OYHRdyNisCYg+uFf3GqBGQlUJ8Pb4s1VCDtjNcHvWVzMzpLcWsPTZ
0+hrikeA2bQRjl4pTGqT2WvOCfaOGqaoEsUZqWgOCZLWSqkmU0FRe27EUfLCe0ML
EG6yTXfxMm7ehVrelb/u21jd74cG91TM8EqykKc+cksUHTI5cNHKNh5rBG/dC8Es
YWWPViH8AhLcjWD0yEWcBMc5iivcm0R8EWPZN3Zgb4mbKNvoZbNpQiKmZTElKozF
nNNFaSSVWETxMP8GqsA5Ot5aSJYkOHx/qYyMadY0MzfUxcPLYDVU5Y+++U7ovis3
cNf3xqlTh384rg+Rmd1pee9iarCp8l8bynzB80aZh7zCRxGvGReK0Bm6O9I1EPMY
VxbTSPrxw5ddXGsgRwj9kwFjvcbVA9hSx88L/Vc4DbklUUYx/qEIY+LjW2kICeVo
uT48N8h9ZXN95GJQbNsUN8/SE9ek+f+TB1KEPVQOv0eus7fQjEQF6YPgQOPL+BUD
1eP5o4jRgQJAJX9NWxmBKHY9HXESVJ6gZxdeQNnZ5gWjTPzUQEhmTqdSF6JypWGS
6A6iS83hyyq1sjtGmeO5ob8fEhyVBhZEhA7/n3zcOd6tuUGM9ovCVUzBfR5bHG/r
kvBP/LYD13GP+FKf4G5ipzf9A3kSs8xF1tnNga7cpVw93tSz40b2yP76iysC2dII
mSxwH/lZLnQskchmlng27PdKgoqMd3A1RRDfpo2DQJEImsHfMHCsXC035p/6KzrX
7uPdzniLsOVuNhs3L2HOt/Qb2y+zNogiUZ7bT+lkYHixjWHA93E2H9cE+E3hKd0a
GhqsGcRIqWMbIOvNUTXmFkkz/oqo26pKZXbXdb7nvYr0tY982TLsV26pWFg8jikw
pchIDMonuD0hrjwCNNHxwf1bTd3pIkVExx/AjXp15pmbS6BBAu8rEh/qNIhBdt0W
ma8sayCg+nt8jJzk2r1Ht/ez8WCTwxi4anjIemlok5RgD1nUTfq9PqGWsj1MJ9yM
FGYbZpSSl6hlpVULpNCrhz2voGgQS/PaOupBoRYryMoGiFNS8m+DBS66NeqOAK/H
tX34milvKSzhGvdTcLQZS6pB+nUAjQKrEes+CCTvN1u7mTVXRBP08p1RSeDnC/Zc
SvzkdZR8+ZVyiuofwCbn2j9Y3thCXQSx2Szpn+0cqbAxmWB8wr77532A5VRuwVWy
ZMut4/pOozrl5A2VcH+ViyN+VYLq5zHm1wwB0pXkR7dfK0/KJ6Z72iFd3/UvL8l8
PPA7Aab0c4/TEi2BC6mMekqU0y6iE95NI74eMLlHvr8cM5HCSPhUQPsP4WajVHg2
gh0OHZXHCpjlkZ0Y3VRUnmUgweUs1LIcO7uJFpjfKNecg368XZC0Au5rgizrDT1q
U0ZFsyOYzLLeLbrwgdhu/sOiImA+w/2j1BrqkQpVQxEOGNXI+/T9caSCRZuoaY6U
uVWxxBbOER1o/eq1AKRG4X6rGN108SEA1AN7GaZ6wLBMZWoaCEV0niGe8ZWAXd+G
QJdVqbo9rHbWWwIV5l7WXlxLYlSDdqJLAxtRR90he2vAvDt2uW8+nx6otNer9UCX
7fAoRqWsMs864AVZaugca4MmifM8Ok3Ue4h0oxNVD9imF8XcQ7I/VP969pvycgaq
/sXTbg/ES6ENUZJSw7QHPQa5AlR6l4kypP6u3jn+CV0OAvx2POeqzEvD2KJbTKDO
I6uhoz058odIxtqHPGV+GTUJRgf3ro5MZvkh6RRMrX58CiyZFkQtrCE4+4TJFvLp
lZ2wKCM0ceUg2JXJldPARA==
`protect END_PROTECTED
