`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KC6nnkMoYvDIXBkG7nRi/aoS7nbl9O5yxzDPhTgVHLktucvUyas+gNu7jIA4o9Qt
6LLnokmMfLr12cASiX29Isajpzdq5sHp8un08fhOugliJ6oa8PQcWifdKVeCom+e
HtUxyVsvRiHPFc1HYxMhFr1IwoSxlwNQxCOFHqMsQXl0o/slvpiTOKkQcbZUkXt+
RX2ab2Mhb6tYDFMsdhvVkawM1giwgqObqDJGdtjaMFnNSeOrsWuXIefFiD7jx1Zr
Svq0X+cE1osCTDdbw5THwiIIj39d8vdCo4Eapq+mdcZ4Ir15l3WW2fx34+uIe+jQ
5ed/B+pmxuu712Bz2ivcmmuJDYTd5qNPIGx2mnjnXydnuJfe/OJUW0IUSOMfFjd0
bNB6irinwxLeIGA/reQzSZ+7gFCSX2KCo1tAuiajN0ojTvCZP8PCkSxLDYn7uj8A
3KBryrFDCvL3meA4YamfC1acoqBB07A4FTA68FBbXO8aJs9aK/eKVqImcfAlZZe4
7tlLA0DBzkmNTNwKtELHw4Xn4Le0FYMfqRR+SzYVQb3etG/ZhjIwM6KaDQGxBIC1
wpdln8Xns7unsprIxQkIywydi6FNG7HiLzQNA5355K0=
`protect END_PROTECTED
