`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZC39bucvff1HHAeTJ2gxtFIrjybypyZcD9Liz6LVfoKU0HDz+/IF6EHb/teRztY7
4ilt3eU0Kq7K5mw5kTb8NXTbz++xlp2OqA/2kJeGikA7yC3Upc0LiZPUYXCupXMZ
keAlMUXcovDABGz3sa/8pBEe2jyKfCrVGtNhKAOM5nPMFr4BUyayaohxa6vqeF7A
aIqQzCGAg8AxHN7FTUQU6ITdAo6UoET5hSnz8XSVW+6KjTix/vyaVpCrJnzFKGMY
A06nACxdTmZ43pO4Dlw+++KND6pu5f/KRQi9BxrGuIBRMwlnz88gQFbzsXixyLiq
9ku+PmGbX7umiBFBS+NznUj28chTVw35BVKku9BG7e1Z+TkGAdLcN7NIv85zW/kO
U3I8GHzYHvTeTV+gO2G8CmXfhE2Ll9jldqmq/rfq0icjVO4L9efY3GKRxoPQw3mI
jvuK05ClSLyo+xUlAsGC5Qs2MxjTXHkkACLRkHZkWK6Y93gT6rd1yPmtB4uETKly
0BTsUtxXH0J4EBmQmajFR7SPZJlAimo+xAIzhfmq4OTQQf+6JETpKviRxF6m7rh8
2swx9ALPgi4QsfJUO4mw1zyzhTvmqudc0rKmNPfyhUVBrv84ZhvbfS92aD6H+JWI
VJhRQAO3EP7CIM0o0XaIwzj9zlMikQ3CQzMUzJhTNMeF4a0ZBmU43dOjPRYPY/3R
r1g69yTACOv3RSPBvdBM99G2a9LcROXfgGf3YAYMvH7qiGx+838pUguj8XXc4XP9
d1shd9eiVTfIUSpjrFgySdEbm4215uECBQj3ORNRKuM=
`protect END_PROTECTED
