`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i4F1mRgd8p7NK/XQ4Cw+fQIAhGAJaOrpp9+3omA33s2i3UwuQi2Nw9pTrPy/Mr7s
giQ2VGtjd3C5PjJsX6ZXJ3gIwble2G9Q2ULJoKFaCoHcJXdnLi1v9VfFmpMquvBM
+QK0C7cZFBVuaVRoteCcseDI701xUd8hHLvu39sTQ6w66b1ZttMwG/N5G8Yh9MZ3
grxA6PdhoXZmVIdDyoOrB4Q6h3oWCdYpt0Uf/Qb1Xi4mWo547dmGnL4K3Mteuxb4
BxZDfbnXCVDZ9tESkE3B8qoUdCPnU6wc2N1l5rttysyKioBS2tPe6f50M3+VEqo1
moU943RB93w3/SdKXY7Lh5Tf/xPNyb4SVKmcXORA2OkQVNIVPV7m8u94GxM7Dw4q
AR1IW+2Q0tIpr5TWKSl8F+nWE1HriuiJPHm4Pnl7vArbX4OEojXPXMcpygk1G5Sb
ty6U1s/Qkq9hl5tRPyWHpULSJjkJDrcRHf76nepPC+eBt6tX3B/eIzBs6x5qOMVe
1Jo3EaLempZxPgoyzB/4sDYHjt3MtK1Zno/zezhWp52KUEba0XN80YsRE1zXIGdv
0H6lUpIIfapWRy6CneLpDAGVPePGJ6oKcYk6ylpyLi3XSRlWHWmqINTeEsL8INiG
dHB7H0t4whrGYFx/GFFYt5khIK/H4HkXlpw97af+a5ronFVvT5WTUjxEfc/5Fum1
eed3kTSDUy3YvT+Y3UA3f8f1Wj0yEBax2KchKP07iftKmFSV7nNGt6yV1GvWecHk
6wT72ZWrEX9VYMxBMGNFpOyNh64S7/JXwS2nDX9VIhhNIMB4hOpnSJw/iUd1dLT6
uDIqwuQo0Sq2PWxsPMrQFHrcPXevnVjWVrqBkXcTLtdgYwzczp0XDV8eTXqyfjI/
zZwRjYsSElWrhW7vWyBJHI8Qxoe6xpFg46dKEaPDPBCBac/UYRqBro3uIqiFpgS+
j+4xSYfCsWC3OBJ0SSJaNe6a7NiRi8L9c3bo7wW7WQ+Po1e+DcFsZZScdOwKGzSr
Kaf87ESUrnq8GYlfB6Ob/fhR3Z1EnXeFjgSU1cbk2OM11V1T/c/tHh0pppGyK3zc
UAAlzaja8KFORV75TcQi9KmXAmze5AHk9xyrV8vEY91Q1fuWHmTpFneaKdPRR5nU
1cQE8lXJ2EenNiM6YMA5/rCqxdxq3S+2qxBGD+4/9Bkegc1+c35zoE2+fXq15E+C
zvfbkjw/FLNA5Cs8kJU38WVTj/BJd305kaVpdBvFM6RA+YcjNhdFVZcbKhbUz5lM
5MrKjoTbUdukjNFTXLQhjR2sSVUPNK1qBLT9nnUSid1FlzKHyJq943Q1JxKRlVTn
5LMpb7vzpVmwhlhS9f7Et3SNNXlGsH0RI1qsCcyA96AZPTKgU5BkrPyzSV2gaR31
zrasEs+B71tXAygv/ds/Bqkdp3X+RSKiDvpQOzucUJ4mlrxIEfGCmcKz2VKoquNr
KSzsvskxfA36YN6BQ8SqVdamJAo6xbZYZfubcE3sBtvog3cJvS1Wf3uX4n3MFfy5
EKEo024wRwN8sTSdLM+YW+JfBITjSUDhu9G7w2IsmzBHUVyq5m2yfEyrCHCec+ws
+DMKfpObYuq2xOxgi/FIoXJ3An3NJVNsNPyuk0tu955grnVLwnxp5Cb0cuMjTQEy
vx5+86VTgFrV+yaO+1SsbKx/9IuQp6vDrpk89pRsK11coRMFZ3lMB/DeSKlujeOq
BvH1xf4mjLT+fV1KrSmafWvfbKi6LNnTnSDYltyGuuCpD/hQkxrT714NR3GxKdIy
kN/okZPZe3f1yh0oGYJPgSsotiNagMa1EDRSWoLzFgFgOwhkfJyCUArJKlt9z14I
qOOWWXZdo3XwcF6y2bj+2HinsoghPyx6FMuRlird926LlKDLqo/o6r0vhdCBhJg4
GF8hUdznquihKQe1Pn7aB4wqxZkbAZ9i6b85zaBCXdi2CB/5KZtYmUUVLohorrur
qs2/ex+3EOe53RZ7LbJoZ0uBZ9pOE7PThN/6B1nFDf6xSs2ozDWZw7dIY8TzkNtg
UHS83/yBz9LQpT0ga5gd7fj5jDjvZzErpjgAoRldECaqIw7NeQk6t6U7eGOFCR6W
9EABYltxAQig8dSPry5jmIU8oVonjBqrAcxAPYaaAvZJvnoDUbGWmH3xuETeK11J
0838AVT21ERB1THiR+jSjYdhFiCrQxnVfu51zObNaTqv1GucztuOhilm1LqiNu/M
86JrX0YXXtGxTOyc9Lpm4PQChcdZZYvbWKilmfDQyZupoit/UlDI7XKFxh9wN+RK
fCCaCX9+4fmWYTcVzObSBwUT8ZU32vtBRD2b8zvEN1ozUOjpZkMxSC2qgde1mOLG
W/8oqt8j3DDrk4Q0USK12tiKAzHrwfMBwekLdrLQVGaB4NdopzHF2RlkdoCsnOPP
GtakoVE8uqXtThyzJlR7VXI/LXicgqxw0EZAVMxKMbe5QdIkuX9GWBYtoaOIfwrM
ZIcGgkXbniHb2dHH6n24wzz3Ow3yRgsRIOvh/x/o8Is511De6XQtYLQ9RP98czUm
XZ7xirty0dfYDrOOEdhE4O52T9g3DZWLsgXI2yHNjwOKdUEcn1zv8GVcBIuhINKt
2u63Ajm0GjO5NPvNIr6sQf5XT7WNip8qCt+0Ehg3ROShR3ZjlDcPWJhkzH6EaQLO
ZN9tEyQLP0vSS+NqY4o4dCRPlkrukuwS6SRyAQ5+jQQWOAT+YLX0iIT3PKGjPj5s
K6UGk5Mi4gkEFTGi8jljmtk2I+68s8jRNUgsrl2ydo8IinTng6yTk2rkmPC/W/U6
dgtFSDWxDEFcQtdor9cfqGDSnCh10NRsk/UYPJdPGOrJe3JYKw+GV99daWeLihGg
rHaTaSDISnbYmFqogxQmBtQ+ZNvaRy8r5LuzAsheAcu+U0bAlRgz0rBU8gbrt3Cd
081/0rC8cwwC8a7LROdmo4Kl1zEbGcWwxGX/DxteUzJuxs15QR1IvBuMiZzblxVW
dxZswEp1FIFpc8pDtueqygO1V9DlXEqoE7XbOymr+cPLBs4ejkJwEKLkD5mNPgSl
D0Kb+jjEV+eGAEvDu+IJP0bCtUBiLtFfsTKNNQsnDxWxqLdMCIaFDFFSYMDt3z34
BfPepbiigPhygsYRucuSjdyOizYCUTUNrrSM95+3QnyjVV+nJ6vs2re8SOguSvMW
75ABgG/mS/M1+uUovhRGUukW8dt012IjQ1QjoRf9N3nChGuY4JDIK88NEJ2ICybr
U0/N01UckJufrSAV7i0WhZhWr2dxrb7lHDkmFWyc+1Q9wbh3xOfOl0uKrub0C4Sp
bZSBTtBaxQX9EkZHGf4Xy+DZHpPzRj+nqZOKYIPxCo/ta8yaK3SdootNWA++17l1
QeNtkeQP4T6wZcOq8vpzAVvfvZIvai9l5bq6D1nkgv8pt6V4lH035ScfeAmnGrT/
h9TUSDMqGanTDm/dOmfsHF8k/4K7agdz2Fz0TonmME+xJslUUhdKY1bOPP+C89bZ
/UcmrsZVmIiinJTl/ykDCZcsGQsEIQBliYEl0kyUsa+zTc5fzRSgONGI6+Yrq87O
yhW2jgJZdf3a7BMCunQYW7bnHc5fXs4PPvqrekisOWJXBmnKwoRFbu5N0HJybGqW
qulxL0jwyukhr2Q8Nb8YPsu/lTSVSHVeSSGi+8bK2evqArAzASFUQwNqZDSUsYhi
OB5Nb/Ry3ImkSZGdgnq+e/QTyzih1Z+zTbHABKxV4xjDAoGfe8XgiCMpK6G/kWrJ
xn3Sv/x1MJNQiOLNRZVbVM97BAbmY141o/u4BP8O+qed+EsUA+TKMHM6Riml47Xq
9SomeWHPSVUitFOY1Qki7V29StgCj0FysZYoROmJXhP7SYZkYFGGUe9o7nvHTJiJ
EDSKHZa6iR6fQRPVULC0AXFNONtiVAQ9akW5AhVwG7LiJ8qAPZzeZg/G5pl+9uuP
jXF/MRSVvi5m1v0XZ+A+isZT4k/KFmu/BvXMxEYhttyK/mUhEXytJpgqjik6XUyu
huIQS2ttfCOdNlKnnXSjon8AChkjROdiUCPNE+p/MxbDtDHAOV52FKQAvpLAvwmD
MT7/6tslxyOWPzgixas9/V4/uNU+EkZ0KSj4LYGAsszGnQQndoO2Ky6YQ3gQrqhi
Lo9sbuiriF4bdRgaQdl5pzCmEGC8HoBIpROK3HSLcFQiSofGE7OrtNUtTHtZPUoY
keSgid8Q6ffdRK14MWy4WqdqmkjQUmrVLOJk34i20hzRLhkBy/mFwfBw0fAdr9Dx
trxRajUs6NLki0VuV6Tc+VZLkGy1rSbZuyCJReARyZSejPppGT5tr/ED+/BDembm
pTf+hHnXJZEo85wQDd0aPmlc5/mtsv32m6JtGiVieZvtu/DwXLaVZPBCDuHKMClf
5jD1evP9yoJm7HPNjNlAd2TaLJnlIo+bD8uBEYcpcht9N8NWETTWrDaw/o3pwIqB
HDcqdX8qXL18KdSsxtOXUj5Lycy3wSoGOs+5fY/t47oa+2xIbWSld9po1OlppIus
8XuiJc8929xXzFX+NK6Wj+PI2YOg4xXapGI8BCYrk+5lx/OPFn0oG3pX7kVBP1QP
mW3FTUHktN4Gb+TtedzrG81Q66lSed5ta7eSlIu8KlIncSbb04iczLEM5YdRpQRQ
Da67vQEQeklCtOwgmIGyLiamOW0lkL5UyPdEqv/ebTLbKk0zw4UJy1VEp4w00ONz
xlpscrLHsp6sVVodTSftVMS5RX540BLrcYaaSOZgIKrntVVi84YzRvqgQ//YElQa
nj7C28RPTOnsA1mpXSzsI3S9hpWXnjOFaHKEtEekWNv2zLNVsNseCa0zGyjNYr9d
c3k9n/3GWOeESrmC/EXPktUt8x14mOuvWgGPR2IDUcaexOimfOHCkM07O7IbyK09
X7muROQ1QJK/5c/beVxVxXCQebC0FiFacyrMcxZkV1OQq/sn94E3q0CtPPYDUWB9
jf8fiLeSSbRH6xxlEqlWfvGPBRg6wplttUHO9/uPke0qO0zUVG04QJrKakVNVYik
nrup2h9aulzsvRWb/N8vFUFD9h6+kYl9/VX8rjcRyhbGTJbMVo/oNz17E7ItlAaz
rq0wzFCgqv1aw+rT6VssqR/s4p/+W774g4xhvkb1DVJ6QlMsfa9//bNifQjHZtv1
LCL6M2aEZ1rG7fmNlSpbsfklB2jFvdAsrFtYoQGLTDlcVO5xxuyX4/BWg49hlQ8Z
h6083yl00qNAF307C3XVIZ0/GiP+xf04UPey5BLfiXJUfTeQHUv/quauZ4LVoiII
oclwiiYNGOjtmTKpeAqlVb3BvLGNn3zeSOk8JDxP5qmFRD+fvLQSJ9ZepLyRFgeo
XgECE4iCAoTeg00CbZe0XQzsz4h/UeHuuEFbjlljN2FpZZh61aBgTUovIFJp3rTG
9RNoohmoIvJe7PX8L9NYBhIl5d4eekO5tDkFvbcl4XooBfqddXdfZjtRfO8C43LA
pgIXRTOPYHy72/CI4c1Q3GI9r6tj0yYgzUz/pXgdg4irRxLczsrdWsKq3nBEETI9
h63U+WjBYpDNUr55ETTv5/p75d+9wU57QZ3muFDmdMm/k8ztOh2KN/WAwu0WNUB7
mCF/FPSS7PhOfPMlF4Nu5YFl6B29C8tveA32YE4MAc9QAe5eHSBR+mKrKwnIMLoU
Fjql56BqW3xaKYCJxyt/0Q7zoE8CdfN+7NTcLpUh3M+MRVLOrui4s+EbomcSes/U
yiGnb5yl8lUjzsECVgYBqDZ3p9w5mj+ALBMjphLIRn3a1vX7rPLgwG8Kc18WMyhY
0d+8pPolsAOB0bXUJpslp9xA4mKVI4Gwvd2DKoMhMkLNTd/UMliR6YbZLOTOQ8E8
OkHKEOfCtPdcWRFfY5uTD+EDh7bX6JA5digG+r3HOvs8xagwWa7wKI/gnY3z5hve
ntnYspuHy3n09f0xRDeM/SRrsLFcAhVwvZTKi5fYNJhXDy96tLtV1ceGFn6LYKVV
Q3NJ7SOAnkENpgCfbAoSQL7uAQyjqyHpIIQeMTZAN8lsxKeuf1nqH32QXVUiH6MC
BXFY5CHP6OYd1c+e+FxOsBQIcJ0PlkeNmW8Z0bLxkBjKss7MIEXFyZzTImWpsw0G
I0kpnJoscdDdXkocj1r9iEPg8bI0EDqth553+jgpo6VGrZ2eKA2gAGLPmIeifHsu
rUP7r4HxNh+AG+Lw7f+lijUFbu7Oxw7FlvcKrUPS58woWb6w9NR268J5+U9EecS/
0nbmd3aSYxTShanch0N5JS39WUuqjORS/Go0S8ncBtbZDOZaHhIuSEXiU66aq6hB
in0pnu6eNP9oXol207r/7feZ7+6XOa+LDwbeaUDZ6GJfRfR6Ui7wicx/nwpRmd35
w3XWOUMfsW+NspsIWY/wE+EV4Bd5K+fisp/m3Xu/YYsiFIiMaGqfpz3cxsSvswc6
LrnCEUlrHkxpRY/3lmZgSmf+D6ZluOkeTHhd82JfbkJ4SU8KOzXPUaJXymAlCDqq
XRpfqXx7sjo6/B/hwCq5CHqzjW2SUhqgDB0jVgnf1x5/y98JpTgV8BYDIcF2I4Yn
S6ywh8SqPwAGSBlh4uy/lWGP3cBRAdQWZ79F1xDlaIdAbmrAdsBMGV49LR5YYYoz
urGsHyYizz7wj0S54XVBSBkx4vZGqpx/h3g9APPWP97ytZe3pytGVR8khPMSMjMz
8Ky90uihvzmJTmsN+kn8l+Hwa5qok73l9EsjDCynS+1T9N7yDDJXpZsMcYLM+i+q
EQ/hUw2vUbJgTvyk/byEHjJoYZs64W3GLzIXo/z9ywU=
`protect END_PROTECTED
