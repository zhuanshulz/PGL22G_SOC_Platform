`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0mobUtUTWH18eFNtlQFPVwQxFlJQ7kxgNaB8qzZxTB2LluOuXNboW+g8MjJcFje
X+0vTin/9ESpZ4Qkn0rCYqxwUnKbb6id+zfuqyA03GQ8kkMMvA3Mm8HbqtRA9nQ1
FSN03qfu5/kRie4P2x5eqhscM31KmyuO+JjkqtqYU/b4Tkqo2Y+uemTH3PxYfrXc
fLjZgdTjMwfyP2nwEKeiAAFh+qp3HTlXCGwUrDa/kLixgUH5Y/knLom80c6p1OkE
9077GqCVS7DTjyUHyOgWCNu7SQ7X1+dKPyOeo9ODGTrCaoqCKe3nbNhAkz1sNv7U
XgAtQj5E3rdPlwS8WzeCJ+7k0DlFvjhg4XzXBBSwWupnflVdZgxVyOEsWx/v3+Gd
ixOdxAaL4Mqai8z8KUO2QXnYdCmig8W4zRBi/IXuv8ZhdBMC2yloS/xzvKigfsok
JhBVORk2WtXnMQ+5ql16u9GS844/7xaGXAyLDdeBRN/YtcIl0pe8DEqJHCKjPbov
`protect END_PROTECTED
