`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EOnLl/6O5PyS32eVGamwFiXDfkMQaf+1uF+xmuCwvpE1Llo3zdPAfRG4bsM+t3y3
Zo6KXN5+l3ct/ujvfidjzrXjgi8cqLzU0QtpA7EGRkgYC+nzhr+iXeGxXtPTObCK
p4iYWYb9fxniibys7fxrA5HYugbw4gapsGlxxAOBdCsScTt89qie2j74BttnxKg7
dVJst2AX7ZeiZh825hkLramn60YupI9jRd/TPna7FbqE6Iv4ceLbK2VFo1VWuFET
IF0fBhpMALNnXq2s4/Teu3X9U+zmWAwEPdlQRfOG24kRbdh1w3p4KDsw+PnCxXKg
MyWTM0Ed9RghO0EiTIkl3BUxwgchf/uGUTNUPHZjQGX/Be8MUEiPLjgdkMgizjsy
3UEe47WKWLppDFYK8Ns3GT0mWbC2Eyam97/2EYDh5n0iF7SvnqyLAh9E53rwrTrC
piCADw7Pctt6adh/Uoi7hdRy2JTGbLJEWhp/5XVIBTUdXevJFAeTnA9Nde5yIM52
C61ts22STGT4YGebwlnr7QiaNt1H2PLIvi+9NlNKFXQkb8r5srdzcOZHJzL2DWOv
/CLBAZ5iWxSqqtan5YjX2ZJIA5JRNy1RtNdVYsaKei7LEoF3v8Iv+378BwY/RVH6
U+yYeuZeCUrYb6/Y+cOWNQ==
`protect END_PROTECTED
