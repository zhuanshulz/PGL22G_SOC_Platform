`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pCjZ6hIq2PdjxMbe4+QEzaVCu0nX+glgh4ft64iCo2d58HhGGw5jBFIgP8k45+Xp
MGz0mk4Jk3dgpWG98CRTb4gwpGBuVxQ0HZXK/A/QmRwDTVz5UrEReo3lM1ShzHS0
iQELBNZaJNBHnpCj3Cus8cZ7hTd7ZJ8LtBHqQQ9tijvvDT4GDvW0AtImiGeiqjHS
eS78WLOoibr7N6NQTH1BF+Iz7yXqfngfkMxoLS6CQ2Xc33RQ443dDPyYtlr1MYal
`protect END_PROTECTED
