`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A0osKW5OV3wqRQVCwZAXk8Gdgsoq8WSRRmDCq9zKcpIDosm3X0zlArI7ABxPeSYF
KD2t8j7SzfyAFC9qO06EL/NtWfeM2exsWg9GgpHZS7NorSTkOw73VVW8TBzFiEDr
Haz+pcmpVHRwEc729p0gTHQIF18iEKYFfAwigocw41kRRPTfWaQABpdgLFOmgcuC
k6WnQwZ5JH186AoBpNCdUFOU4nUxonGTW2O2uZE0o8E5c0MEAocbQYjhGOcHENM5
OyZynx+oCISjVn0x7Plg41W2hewTpn0WGPZSrGJvV449gvSSHWlhG8JPxkKPK+9B
QYzbukbdgzA3ereo2g6LvdjYCUqX9GASeG34X05BlvlVLtF4ZUI2Yf5JFeXe8CYM
segAAoufWwv18PDp5XKKrlS+LbdFEzqoErd4/8+W4VZzxSFP/rPrt9stjo13LJIa
Ln7QlXw7MIZsUIqqwrv2/P3jM7k6siw7P2czsW/Zo6fxl+nmQpBZYNgoLrIQKz/A
YBToJI8mYnvocQ0bpHb7AxBTP3sQpFCKbZCbgM2cv94ZpkVLwD93qBj4xGOozfVw
ikykphK+uZAmof+fNqFlkHmFOO8+V58d7WHs33uumaBMoVibvhWjpHtfrLauniBC
hwEKzAEq5iJAQWKVFL4fbCkL+vwQZO1WuikVYcRNgJq1ZHW+YFLmQxpptBnKEfl3
GB8qJReVo4ktWD6CGAyI30NnyopqGKq26SSFwqniqD5Iv8mKXwlTPSDupQff8IAN
TwlvDhNeiILuA8xmN8YqkXKejQ8CGkqMo50afj859C+3keHtauap2tG52pOvX3DL
E6UejbO9fZpPPveZSy6N2HC+S4nf5TsU6okF4bR8UE8P6ooF+51/nxc7qJKX66a9
p62vXT657AwPSDHTYAihtu48RhkjUvRIDydc5yTjKVvB4cs7VpAWjo0r+4uAu2+m
QlKBLEFoT7mwhmDN6WYpCWyvtUuTEdeCWfd7B0sRyp1xqG+aOzGF8pl+QwEFtrgJ
Iob6sDb845gwqZLORi1PlBa2YMhsJJUSnDoP+MVI1VvS9XdvU/4M02MmEV9EmNoW
OGCvbRoFeJC85qVUEqnpMQIlP5jUeShG8H1n4fuxB/p3bCO4YTRvXxr6xQeB9p7m
fj0Ck8jjxfN9hy0hfmAPRfUSIuxYnWwHdf1dBZAk7PmVERH4SeIl6KM5n2cghxNl
IfD1WzdjotGPAph9DBZDvneR/vQKodTPMtW1b8Sq6Zb4iXbGC5OP5MkLUbDNw7yi
/x+G6yz0PlKf/sUJBWeyQgXrdfqDp4e++isKZ7VYLJ5jgImIxgkB/kxpbuycdXzR
1JhkJ2FdQbYeG5dIwVuB1kxk4z0mSxw3Crv5iV00WaJHGWpWW4Y5YLdt6mEXhcCp
ZaCUju3UHgZ9qRCxjNQu9+4PnhedEdfcNm38+fv0QmY27hG8j8d5H5dxj3r/7wW0
/qs5PldDhI+2zXPJH7/Q5U7b8z78vA6G5C8XmAzgG0re4Ie43aJpuF+uIeh+YDGd
QMGSmqAH7uHWYgGe2288hVt+YiPTfVOjBdsPZt8AwgDC1Fhjsxk7B02TflfyW7K2
pdSKz4a64rffJyY6pi6Lx+gz3z0tb7sLcgQOmItg79JmLZVzFRZ5zTi5oPt0FyXa
QapJ08I8sN8QJbj8k6MV+s9dWMmZzmKNZBugZx004BFG/UEY7nz5m6n+bxAhTFrk
NopiZC/jhVUriuxGwoZXMIaiJQTUNLOSgg96YZOe8rXqYRqeUD9N4Pl7/dSF6Gtd
8+9zm3eOqIzqpvmX4OOYFt372vWD2ih54KEE0sGgO6AxCwF2DsF7Oz1N+/y4o3k/
9mX60EhU5Y1gYFmYaixQ8RjoB5WND6jzIR/fdjTyvrUGa4Oep7Ew7J7GbMtvJD7e
0JrH4SRNihyXcH8ycTTo8UvNFbXfprzqByi3WizpJl2M2ZzGisOLSnV6C5CwQbmf
flNB80P+/0plCqWy7Ersae8LpkM/SEqKF9IGfwJRKC/XHL8HX/IJnQnO0pMD8Bpw
a8F0EAWUW4g7+PTVSv8cFQ==
`protect END_PROTECTED
