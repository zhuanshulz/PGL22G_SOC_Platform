`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Crw8CDPyeTBbQs+udAMbAaJVoS6pnccb3ZuSZYBitTwm328IStdYHYgjR3aNIJM
ezW+piQtgpme9M6odAr3S7TRJQD9kx4vKV5D95FTphqJ8fsWxrvqC2InWN8FY7Ns
+IvhNIk19HQ4vW/7STiYOdt6SolRDZndthvYQahSlL+H2hDTen3naYi26skjCl/8
Ryw4tJp8B967deD365dQPJYLPqznVd6mGq4u0BrzB9yb0AFPwvYl+6kHvL9ztwj5
fNUHr5tYkK8pLE34lIACtMynPQQUIceohcTkuf0BQcffp+vsjfqVdPLCu8effoW5
BNAOfnS8IJcL1GKsRe+hDLHlYYkE5YmXY+fkugZKsQWwGgUrUG75+acHJZ2zehsY
xzLju1MHR1CC9iB1h9sY2thlx9aafDw2S8mXGRt0YJESAXd30CLewVjblv1dEX6H
DNjbAj5VWt5RMFHf3ouGEKpgoK+0ffd893TScRH3Fez5bFRlG9vAyVgnJ1iDzaY8
FOkvPs+BmxyMBAhMl6WUu9tPiHiPU0CAVHZEKfcZx9faISZmDIScOh/v+sCelnHe
Tm7AC40ZRnxw5iTxShhJupqSAkY/Y61iOcK89u323OUihd91RdfpPlH1QmqwfrmQ
t1C9yCbzGkeOx8FPmhQ7dYMBqaB1uw5SDYdUTNd5PRgB5kccqTKO1Z/Jdi5n25JA
Avr/7dNWj7WW9xkG1c+heUHiKiGJsMxRaxyH+D0PZND0aq1wxjozWPwkDLwcWmD6
Xhm7EzRn630Tu5UC1gMe8xrDPgUwny1M7G7ATUSBKpz7tb/A6lwj7XjU5pHKmXey
IET5WFMwMceuYYdSLsMOj3TDoDzOGew/zxrU38ysVdoCyB99OWioTaLPuyaRCVrh
FYpifJDYecD7i8pwvBkDy/yeYiTbCnLZPe9fZxUSmUbJK65akIj2paUt9jH1HsR7
`protect END_PROTECTED
