`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bwr+FB/0+CGa1JgzMcRGqs6r/XjW7EeNncACOoAVSNDsS47q6vkBs9sBq8WyrPu5
Ocdq/XQq6I2QJ/cL4y4HKBQI29nf5Cn6scF9SwxLfES7PcpZtLefN8eFNiTYh15V
TOcZ11iovowBF596rX2XfdKVZKI8UVVHqAQ31QtC1JCs5YbD2ZWi0aemDihQcOKI
YkI5XMYBct2HQVrQqO4Vr6DnWwmPLeKnKHrfa2siuaGNu5Luw1LEaKxf99V4gHU8
Rk2c8BYT8XxwUPQQxbPMgz1pmXeM4d7BiKlzt8pf2JkiMbgZ5mR+6flJ1grT5/oz
RnzlWijTQMm9XkNcc/RpfGAUIesxxa0FpembbJOG5iw9aAZZcYnKixRxyceNCKnj
hl0F7CXUWOFbrDUe0MR6kEUoh4Bsg/jMy4maZrY9oiW/2CFXiUwMn/DjKKCBkvUp
qm9ws6Dpapm+6/POBO6dy14b3irEitnC6JE4QuDUKrRtd/BuX//BZ5xDXY/emEvq
J7pH/1ZNuCYqyci2chLdmtmdwq73U/fvAsdFvTiX7BdQoLKMFHyIpFY9XWNqo/ah
7VHmd1ewxzhLKLuvNTU4Q7ou/fgQhtcuSNqk9kZ9qKn+Nt2bdkoOR6/FV/Ts+aD/
EXWPk1Ei/0Xy8JqDnij17JxN4qWSdjCUUh46gY2OxheDMdITsjuinOgk40NMpXjD
c/eaWquMkLu97ivu8vCpGaqlwZiNmz8cqrxsVbxFKYVf4A+bOqGf1pjbj0safHUo
chh4GFToshoUiEQrTTvXV2/rPz0kayYX4rvxC1xjosPnKegEUDaKbDXa/PRAbqz6
/kj/fdkf7fb2j2P/HOW2Ym5BgA2s5F+yplNdqzL9GrtwhqC8p590uXYvc5WQVHyZ
xAcznQz9RU26KHK34WrrQr4RSk24xn6MAfXMOLlGt+R0cmKLvNN589Waq2hZEfjx
xZ/tcpghXfBLf02e2ZTaGC/HeXeDgqF41nqoPa9M3ny0OC4Pv20kMG0VtydMWsPT
gjVyVshT4p2YR4dWjOM+0WwjUXBkJfuiEPowMZr/WZ7t0SG9HxFaLnbdbsszuAve
z+SPaCazGHgm76C8IlJdUXtvSw/NZeDO09evOuRRLmIxmCbpl3wF7wfpSzlaY3ai
P/hARjmGYW4Zb1y+hO/UqiRuELce/Zjkj2Hy05he2PBwBVLlBt2qhZWi3dwGnGQk
Fk7cK9RifJ4uMR/IdHST3yiVz9Fz/hZ8oYtWE4aZr5Lu74EKMRqBNCcbFFmGwgnl
8XpbcQm945OyR9ZpUw3jiGrViiD5AUQcNqQqiVbATfDAeGUGh9pk8PFnC7SPSlVm
zVReYA6g/fnmHW8mPByF3vwTbvX7cLkeXLW026AfNFtnjUhvY/xElcwevHi27cNR
yxvl4BsRtbjuKX1ylMYEP+WahZ2iaaE5hWY8gUnCN3K1VsrjT7R0Uwb0h0AczV2H
2oBXXeWNHHUtG5aAONn9uQ93O5lMHl+02f1npV2bBzyFSTx0COiANrdxoeXL8zNa
UxqYZpcFGQCB27Znn3Paovz4nHQBAGl3YVVrVBy0oLSfT9lkIGUV4DaQr6jvHHBI
t6BUR5S9Rirsgn1S4P0V1m9oWXkU+r1piddzMDkJes6kIGQ0I4V4pV1MW0P/Ts9R
+wI0jQVuqhrGkiG6Oyx82laVLEemTQuF6zXhxenN5vU/T8a9aa84zRmXdnqGqtM1
nRjAei3KgUt1JCjceA6gq/o426X8qSsOCEOVrHKROCSj5BNgLw88CjREVsAt39Np
F1PhaGPeTrnv4NjRyKnpXAYy4JzFVkno9//AoIwfRwVYl5Pr7hoyKManEr7Lcj8Z
EqVy5n3E20KKYll7kkkEgc54IaUnnRHmTRfG4XS47tEg9QnvUDoEVYNngYVCCHRc
j3t06A7mzHRhJjcdxFQPBmSbxf/kmsN0Y8wnWFSIHMTISKELJMZXrgjdV73WbCPf
srPXjUVY5tiHf1ZLcqXFOxQY3ya5J2ZnRe+ES9RNYysUED3MfaLNX8LyOZGcGA8u
OTHxXAxKyyvRPt3+y99oHVzbXjETe5ojk7bI0e+kgwSkZ8oXrYFTFslEd3XZIs+U
wAs6ooVkU+XFzfPEQETrqAOR4IH0XvH3D0ds6kV8QzhlWXXNVB5zBpHcm+r9ZgjH
3Ksq423amNCTN7FFS5PIE2kMphohPHhTcPjaEqa268fYXamR48oBL+gSoFvT5TJ0
+zVAbnJ/xGM8hMyhYQc73AfluO3EI9q04mRDYrXulpJhoS3Q2KoOdMVleAjUO0Gf
YEQCgTbPzTARUF21xe35ZUzpFntvh18gPbwin/+9cyRRkbRXZ1yBYXzU1KLIX5Nk
OUEtFiLN8TySvhnXqSyz5JpWwxjyHvlaoKTrhGfNxXtLn6Rlwli4sYZxEp/Bwk3A
1j0j+eoQbqFRKuoyDOTkRedNAURtWEgMjvYDV4RMGAM2vY/wtp8IgdG4K09pTQXT
wFX7AL/DlhPgJGwdYtaKvtKR5sY3pTynFp2BrTY2nuv9axLoDjA1G6P1r5CNoCJv
eszltnHYsm4jstv5s4s0zlb3BfGd7Y36v8+0WQFBMrc2WFu8ho347fK6+XR2Rowo
cd/ZoxhTwaYOH6fQXljz+1TnV2PAYcoNH4Ah/T66RgQaEe67QO1e22Q/m4lMeetU
JM0YmK4pDoqGz/+b8U2yArfzRKNhns75SH7XI8fSKmEHJNu3LwD6dgoMJHOlrcnG
Yg8yvYZ+BgnDU4LKwtKri17GHeLsNoeM4ww4g6dI8iQwxxkbubvxImsE3XqrGYeS
rwJC5leq1/JdsHa3Lkdftq4k5gy6mDJ95AIekMs8n8qZN2DuKU2lTBunbmOoxBJ+
Bs82PABS5uP4weAm4xF8feZXX7ccuuO7CS7ZNl0mDfZsoBZ0MmzYRG9GWeEkKTU4
Yu7Ss0iPmJq24PHmQ1bDYxmkVij7u7J4onfHjqle8+D6xaaNH/WVpvlf4X7PsaN8
ZAuB82CQ20N7OqFDJatY20og6+3S0AGz8yTnNbaTqkjhEW++s7cZN4gmdI+K8u4n
7tyBrmuOx9rDyesDT9W05u9+/DDqy2Q0Oo91+7AjP0r2VVIPnIEeMfru04/JmZo1
LZtBZZrmu6uvTRdhSHEtk7vPNz2V2JMRq6MxMPXxonjTjSU3P0x5cUZv38LRLuxS
MM1e2UaQnL6e+9TFM68wIeyaI5oTlcnB6rfWuoXbPKyzAyn4s+rY7gYzjVVeKZ3n
KOLJ14ssP7wnvQYOm4mxoiXqYr153zLGdfvu/MlBVnPf5Nf641gW87U+M3W7bvnv
fyQPd7MpRh8jmpL8EaZgubK54d0vImEOPckA2mylxQsc+go4q1WMh2rwYEVm8oKM
5wLGiEHPG4pWTGD4PzmiCOGca3AAZ0FU1tEbgLRnP+uaAmWoC+nhUduSf1e+bjXQ
ZFP/gmhgDI4KA1ttK5sMLrP/bvctMCvDp5RRSH87u9qNKdoKyX91o6bagov4mpWr
+Ag/Tj/4CR/wevJdbHAhM5vIyk/ulj/uzMSpHlbqroXittkIfgpR4vF2Fw15ud6j
Dvpk1yf6x0R572s+bQfDs6ftgMdClEGrIm4k33jYLHQIHnGLgsx7B7LMcWshVRFS
qVK8l9dniDE1jXel80BkBsWwFaITmoHEr3eRKjyBZUNpiaiSoMfsedUEmAWJyOm/
LTzO69yzUUpCRzMKmccwleAsWV6XPny8mTBqP0Jg3cuRQE9/njgRaFEMQD/Ik9uT
c9E2YgE0hVSS52K9H2GdSleTvm/iLH5SpDR5czbyDHQQ5YjgzqfOnMJfdJrgAn5G
+aANdu6iH3dam/TaxTHnlgWhengmIZ/c6GCJAR+HFUYhfF0udjo3hGnDltsPJspA
jfsLovpy4l5gJEUGCYmhS6Pi1jlLH0UzM3iPA7/mfzRu7EW/8I1df3vY/zt1BUwa
pnfH+hS7oWFu9P/viG9PGJ9xv/IF/r8cGW7j5Sw/17NgEcQv1/yEwZ2ilYL+Bb08
l32kRSk+zhUfDyaUFFRBWEb8zFsXl+hJIT/DgKrTRXt/iHnYpPW2xHf0BVmFtrKi
4GlVC5oWvLsQxAq7rkuvKXV/E/KTzcGQlQsDaAekTEzERsYlbZAl0oT2oRA7YQhG
fHuTVmlARFtxPH9thtav7YVkgn7/UhARZi4DzLWbzVEOkWpt66u/IezOvv6NcnM3
/gpeFyrqKo86DvIyProT5HC+2XnWJh99A2VmFXB5TpARI7TvSzMv6X1UMBeqENFD
V7uvDOQWUy2ZGOrYi42Cq4BXnjauUA//TRz8TlHzizHMHJ1JlUq3tZif7ItGtOeR
ul+2vLA5Jn1E7AEWL10VtsUIL0xivHkSD4WLY5XZtz9nlgFKKBuG+fbYkGpauGXx
GtKsu+Y2gK2Dab7c0GUrXKxtz0mwTC/J8FhCvFK9AbubyuTPJzMMaS4AXv92gtKL
YQzs+Z7QJFQoDfTx1faOrhD3q/pzikR/8vGYGyR7fQp8W1NHgFIp9s6uneratLXx
MUhY9aX6r0njrsxmkUlMZmdGzx0LFhf/gPJbJMZVzDE5MbeYk6R2vugyBTc5L/TF
ZcXC1VIL4DFYigFltIp39wzG4gIiE57Ow5XQHQniLbcrJoT2AqVeU1o0wppy+8Cq
0wxKTh6LH+rGPTOpTQ2j+YlIiMKGTTjehmIIgagK+/F1ZGOgRtWNoA46dK3eclG6
bRPFFVPJ2o5XrQP0nr/oxuU1PWhcm+9gAXiYXSw8cqvptArhS+RgWCpJQax+jsg9
4a5yZml5OI2J3CsPnDpPXigusanfxSCBEBtb0LKZu7Yxpc8Opk/Yk8bXkjG+hGI0
u96xKfyc9jOjL/O4tW4CdGJVXQIR2omj/JfTFAht0vyURBLk4V6EyuxNMlVD9F7s
5G0l1M0dSSNN1svzVmphJNPXmxv7jnUY19Xyy9aH3t49mOCuVDo3++qzxzY6oh8V
aGHbJgIvt/SkZAusmdCj3f77+L7WM+0viC1Te1/Aio8p8HYsuOVWO/CuNMr9laum
pUNpEUO+835CZytQ/jWU+5A50vdwb10Y4Xhqyo2j7LyIZDzLxi8DJ5YJ5YjVbXs6
vyB2xCKGj4ODryFR353AoLwFgLw1EYE/c1urK0fDbgUKHbg8azB0WAz5kFiJpuPM
oa/GvV/NiWYfihVRc8KftiGh4nHUzvcatQ4Xz7jVnWgxRo94MJZrYeFzC2f7AU7/
NmbleS1bvjkPuvyaeiWOe6lYnEt4SqlFSLWR/aSOD1R+928bNa2ZMV+DQZtl74WV
tYxYM7Wet0hAb2gVq9O2B94ltcIW7Su2bzUyzeU8AaTZYGkRd7To6xIaV0+5FVdD
j4Bs++2MX7hT41WEXPA4ppQC3H0tM5WmkNFgkKdc/ww/ULwgm6iDN/OMKwQ9uBM8
BgKENJFLyQigaq+pl3RcPhu8hHioJCjPGPia5NxzyfTdCya+a1llaVfMnE+Ho6Nj
rzw4pDnC5H5Ui1+OVY3hNykac9yX8XsxfHYt5I/8oKXv3h0Va/nNo5XU6txbn/O3
+4gyuKCJv4d0zEg6l7r1sl2EqTq35Qrg91fHnWSUHc3V272OZg3jzgoTXNZBIc3d
5hr3QN5HWC1W19aAvS95F3vzSB1aT5O9uILMRYRRhckVzjoYNEZfGkK2bTgHa/HQ
WNq4xxnMzY4Z4diWlsMzX8Y5CTHxcW+XyCjPGhI2+5xU+2cULL16zQXkd4S0455F
N2km6M/H9X+JuhybhdpMD5k6jILRozI8ajGRT67CHWZHUsP829M28evjlrr4z8YJ
DHs24KDGfswnHUsEO+jtOqGt+ix8F39kJTfVxjX9ToL413bHe+gj+ngNH/Vt95JO
UK9NwmzarMmu4h3nTGDDaaS7rGLtXqvUSqMXqtBPA3iUNm6neCoxQxKj716JrXgF
nZLhgYnzXvztp6jjTHgQPVP8YX2DCI/7UKpBi5+86aj0fnqvfVeo2uDzdUzGmdxb
uH6ARMpDEDRH2KMP1EGDXdUUF/iviGAOUz/zZXF+3DQqn57DxnfHeReh668HikDu
q884UcwgSu4erI9G1164pgPW6bOd6vs6szQdpY7A7xbWXEXJS/vJfbkFgMHJFY5V
zDqrrmqdHfOyfb/IAZyJ+aB6TjeLwdKqEXTK5kGrT/q2dxEL4n60wkWOJxMPQL1t
sDXGgjr0Jx3Nx7yBXGwy67mlmkeN4RCLX0FjdyYFvVQx5hgDcfc2zi8QjrLNGdVV
FU6pKqZs1g96pru71I2Tkg8RIKRI0fpiNGHE2679FQ8zk8X7Ak/Mf1RW9le3vn+N
MfElBnEvyh0vjltgSof3V5K8btslGcMswMQ5cZGdn2eexghk+6qkL8KMk7u6bmrw
CM6h9s3N1COLthb0lF122NGabVoQmZ73zJeED198evVuQ+dMFifk2atOphw88fkr
XCvouR63r22Ms7Hiwnjk3ysm5HmJYPMFKCzP+JUzVHRfqctMjsqbUKdZqkmwOZZj
d7CwgXdaFfgphfw3hG7c4nsH1ITt6Xc2yFsxG3taiEDhrPF9aaGOB8oXY3jCUH0p
EosVtC+Ccln5MMLOxEkueHzveBOISt7aJvK/uyA4kzbZqP+ykVt5dNM+n3eCQ8Yl
8wURrqtqAoqEpQjoqw7Udr3MVuwV6ANb4z16M+7ktAHuPs7c70aXEckepa0/8/rs
TIPjL9DUYtnigdvLbhpCSaBYPDb+L/1nanitBzd4NnGcneFLdK7IegLE1F+HwbId
dvqE/jpjAsxhJb9lNPFdmBLGK0aZfPppPXeRbf+pSrqDxpA17TtiNlNLHBfGYng0
nDxbtgi5esnjNDaiJuZm557moG5ejdW+r22+AsPJJsFyofR8wGspj3ubu02YRTmD
vCE7Mny/M3Ysv5Q1giAKKSt0hkFT7UW9LtCKzD81j7ZwpvVrw9wkdyuSRTPco/pf
qhLvlen81DSVHI6gGupPhfbP5D+0gR3KuB2YPyAne3k=
`protect END_PROTECTED
