`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQ0IFQYAEi9TuNTbGG9JvSRd8Vk5ZTVOgMnOp0f2fl8qsjN3SjmVcuh7odIfdS6Z
br4wLww38JDZAlR+XZmoJlCv4VxSYam+CKCZtJM7lj24iNoAZLbz6vWXVxGHoZ9d
7r4QqlcsoVcO5h5toZOigT949KyjdA3Bn2ioq39Zx7BaFQ+gBYjT85GEKrQh91aH
uuKqR8rt0Bu/2lB00qnI+QmGTAucmLbPQGGSVxaIwvfbH4FvE1mu2WIgkG2keNXX
mSFyjB1gk9XEEZn3m8ii3zLaop76AYtttTyw0SjkwDO6YsPvqMiL/AwMQl3IBRtU
oKRyw5px7bSyVxQN293dbZLzCRzxoQHzaiPZHSFcvdFQkw0vFjx0j1oh2Y+UIMYz
`protect END_PROTECTED
