`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKtgqtnkxBvYDzXleTir5KqS3DaMaED7U4ZShiyggSMwEbDpfS6jezWOUHZx24uW
WCYwrdRqUjB0+bnaH+ghqoSxMQCKpKfOQ5QAyTJXjQuLLJRC32ptIt0ThpQKkQJT
ETVImLIVmE4drFQODK4fLsvj1RJFHrd4JTKWIp9e9gsjq5GAoNPN+LxOhGVFUNQa
fVAi2VLVN3QNMYAxBEBKjGam21irHq0g6GGGwFjEumQMnmp0epZ7si96CUA733kL
sRL+R4we1OBUsFo07ZZYAq2+SSKWxRgjmBNvRCzoK1om6zqJWZHEuNDD5m0kuure
XIZkMgv3WMLO6a/uDp/4v1Jbl9n/LwMK6Cq7MYkPiYPchiF+DsX1U8KLvbZmJeVf
uv4YomNanU8VAYlMrHhNXmUF4AOZgWluU/z/3XRkwMhqk7oyyJvZCmY9xIHUO2ZC
vQjSr6kuP/Zy2NTz7f3rXtU16uEV0oEhaZpkdVp/IXlOcUTB/zcGzQauSERLzdQH
8a6Ca7eIZVl795vmlZPHWmgrrccnU8v2Ksbmdf+dlGwCsdSrgiPIH1AawoAPwOQP
bVPupBZJHPAx66jXnojVmBmZcuN/SRDuxJ67smArEHzYj6eh295ybFHAgMbnGEnL
oEerug1LeFuIEfQVNcAkG1e1e+IdrIeLHKAWleUocZc2jClqktS4Q/alMtlfxOF2
Eq8sYw3ZEetbK5EDaxru/Zpl7Q41ZWKPaVq2+by4mjx41cy9msLbfEo6nSilLcg4
KTSZP+9Th4SX0rxMgSpPoQ5+zHTJ86Z35U3BREwMNkGlnQZkPklaogLIVFaxR8UY
gP9bjVB7VAwuvuCjpS1D8WQbwQWTFlP6FcS13u8NiIMKr/QKvXhVX/sxFS0P8Pkx
Z7uzQCfpXwaqBOeaz24o0vsYpMYP3lPx1qcPczHrvoYyaAf0/I9JLVubf3tvupE8
aG//tartrXExGymo4/qKHKQo5RdPQRPmIup3bKpeywNzGAt/m66GTbrLHMEB2KyU
HWtS/xs5BCgxLd2Ldxo50xDdkSKU9M2y42yxRWM2coQU6OB4Apskp2rhMv+uPCGS
t/nWDuWj8r41nF3rm9J68BgjOMQ14Q9ROneSffXeXO7pqYfH/Bk0TV6LxcaGPaef
dGFVI/UYCgtr/DV4uZOt4vA33E1aGqBLUudaVjY33IJuxQJU4SwDspPspiG1PdQ1
yoz7lR9iFhRIrDU8TuHj1D9Y8K48z+a8q805ZZJ0vpiQHEwqYtybg5qTaecNqwc7
6avVZRyyoHYBVMosuE7dHCy/m/dnWMTGRD460Q5El3PviPNlizwdfp3PNyRBE1ny
nxpUyxIYoyzEr3M4XNHb5pX72Lw5D61PaWQSXJicTAeULk4eIIsu8gfeTOiyqHxL
XAGxAKh1gUMGpDSrnx0SBovY1f916Nv7j87hnJykLuvNRzLssbsqInG5bGDM9iQy
DBg5W3anRh7sqDi/8WSJVz7z7ZPA34UcFtbEcsov4uGaguIYopVhl+JnEaQPd4ug
o/HTW3IY6qBWiOVkiKZb59a/xn99xyQGs5ac237qd1IYgkKxMTMKcbEcJouDTQ/I
szNTN/GiMWBCOdYp+jCIGE6CfjPfaB8AYZIsZaBEb6XBbMfrK3I8DQCjUDDvYU3D
APsS8RZDPqn390/Cw/TTefNgsWx8kRegXFnwrNsbOMzKQ+buSO9XMNtkjSgn0l43
2BCdPXm9TBqQoXjWerIEsEWm14r2LbJJxLD5mBOJ5AjtnOAozbJ+Jd0fgFgAbRCA
E9jlGhjF0BFmgYCJlX58nhKFiK/Znzta+mTAbQKvqWrzkxKSz8CDqeVGDaPfVICH
1iNj4oF+uKO+G7DltMn7Q+N7yWXPFhdc6zkRW/nuOd1uvXy0LbkinAKsftSZXsPL
nDNGdHOlbw5klvmqKYnKMA==
`protect END_PROTECTED
