`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+poTN7efBkKpmmIX05i3LwZfh15sv3XQIh4/mqUJV6ysKnc/cYmJuJ73zbAI1SMI
2YrrCwQWj4gUnsvMCBNcfCESG57n48QhAja0aQq+MvifNdp1dB/mB9Cn/TcaWdNs
sWnvKgiNft/A6RPkm1jq5GKB6WNS7I6bTw4kwBiCnXfR9NuhXoOWPEfWyJsaV0x8
D6z24KvMEUL6mMwrbW8qpXX66iUd3JlxSpE6d5QhEb+XOpdQ7+++j5j9T/t/ni3r
LTJJlo0nhWOu2Igg4V9lHzsDT6moWkNlSyPK7zXbQkaJGV2K844J4wzsjqaAebMK
YS9fNjF2KUEp0KvjEp4voxXb2lCki6bieqXuxy30YTuqZhVMeKgNxcMuFnVDbrZg
`protect END_PROTECTED
