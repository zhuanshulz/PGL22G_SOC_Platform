`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OnwLXWpvkQdmWrFTPVFDKTLEziOD67z8A3/a2X1Z6oxT9oJoLuY25YVB7ROvW6T1
I68XoN0TtTA7mN6vmaEnvjIBIT5/9etUkDi2R4stlkDLQrld8KXGX873Yi+9QwHc
Lk01tERuzrVCkdSEsG/66ljaqEtYkoTa53BXVDffN+pOF9+yT/wyQi1XftAAtPAR
OzFJ49so7v8z47ztUVELYJteZalWTzBR7UIjgnOhRaf8bkkX7hPYuDlhIb1iXiax
75I23xsHorMKUAkSkV76sl5mwuAt1kPK3bB498HoEV4=
`protect END_PROTECTED
