`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2DxPUuh8cXXZH8XcCEgkg8Ci8p1Nod4IxW7jSuvnNjV0w2bT0HJkD2qZ7SLugoah
HGCEXeOyjhubc1M/RvxxuBX26mbkua1JRXBej2N5J/dtCHu/ndyVrJIq9zcBH6CK
YcNWl+52NB0XTF7gbJq4qCxmroLEDHUXF+Fztu9NuEawL+NmbTnZWEPWPNXFMs0h
Md2m6rYQ9J8wocpwN/p9ioG/e2gst4cB/GPbYyHJN6HBWMFlQ5N/ff9DohxuCv8C
EXpFyZmrRFO8y0Ob5l+EfU2xPCG6ftHwdoFo8pquwdZSXSXmLze5xEbbAT04kHCW
`protect END_PROTECTED
