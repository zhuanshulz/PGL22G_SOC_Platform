`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eT1m3nJVFy/qJ9fhLjSgM6CFub9yR6SR3YQ5riVShEVd14B/L1dOmFxFMs7Nc32/
ppDHY9jP2gPVSBey4TThaR1ktx/USFUGtvgzIYy3IHIXtTHcfuBTBRZzeAe9Cou2
FxH0Wvu7zDYyGMmoO/CfLc3pjt1IvJdhqIFITgC6FG+pp1mIOvnntBmpgaelWlES
VJ8R86lQM49K6+2cKr4eiv0Id4ylnE+GkmYStaY3HglTKani2l5UT81RWFoDSpHN
9GvqD1I0X4HX85KEFw0+BxD81CdT6RAsmKvJmKHhSg1xiWz7GBbdrncEeF9JilQj
BpbYmzCuyw/kg9s+TrR9Zs5zzpVRL5wK+e/Ss/OMSpaqEmjUcn4reIukDXIDgEj0
Q/Oc3cUSfIzxwdAnV/aoyD1DmBBacjzJAtZRyvZAlNOCNj/xSG2+hGP1tnzf/U8p
od9WTHdQeaipcZAOJgJHbs1MXWatP/EcHs5Y0MeAD7jjkPh1uq8lEmfBhXgzMrpi
krL38TMmxcuaPORUZ7P4ZupKjHmCgQubb2vZsBHD/MZDJauiLz9GjznGKsURqvtX
8AoYQvHOLiHSXoRxLNV4NVWJK8MOHuEDt7DyTq/kuzQB9TrybrtAFDUlJ+qykR3r
UojrV2h4LpmooxjEviYAvGEIIFknLSe+W9SmtY/RUd37O/r2lMFpDJhJWXj5D+UK
Ufp5OucC/Z9vdo+NVfCzx6kqbc8aOg03Aot8OFMFNXBpFfzdBNGlfp17ljJXdR4n
OrQATLRPgM0wyQnsReRG5iekZKLxo/J+ZjdjGt5dFP7Ynod5WtFLq6EA+bak/EAb
rrP9wcA3YFIY3tgI4R5Nv7uW1gGhFhQsC+XPHRL91KaNZoU0yQnanziP6HeMTl1N
ABakouDK8RJrHUWleXnm82t9oTjSG9a5htdJg6u1DlzXjVbjtW3wFRx3nrWpworD
ZfDdzD9xODSYQ4+ZQp9eZQmMJfEjCzfBNz6q5w12/vkABuI+TGjr1xylTcVDKbFn
`protect END_PROTECTED
