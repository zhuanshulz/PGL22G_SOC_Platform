`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6/dvGRWH9pA//xMc4ZeQKX6bl9IY0FYjQXF1jn6LMiZ0cBr1sA0AnEXwSSOxbnJ
/u+g5F5rZWPp9/+lv/lFoGz0RjZbOdWI/sfVjNPsWrdu9UOTq4Bbci281sClHXrX
SQyMtsMEzfHVafUpGxGDhy8YBmLQmerY1pNOX4KeuxZh2JzVG3BThWtwkkoaEvS7
ZvMR2Apfn3z91LS0nPrC3ROjNEglNYgiKv1dk1E5Jtwdbj9EHfiMu1n25XRVZjoD
PHG8i6s2NGX3dM4k4iFXRiTvmst4wN2wRmgsV6bAjBtWwEpAVcgf7HQQTPB6TkDA
ren+B4sW83wvgG8aDyUipz9eKydIWfd9I0xjMWKuY45aUWEW0nVBPsazl6bJGw/i
5rCMurUxQhvybNuthwjmGOhnNXBzSXkiH1Tdt6LUE1DgtShkUSSxuR3MHsGuEPUK
c3Ftbso6L8mZmjDyttn2DHAS7ikp0QXmA8Y7ouWWB0mKEnfD13OcadWL1Od2El/Y
yhCedvvu0wtv2CJb/PjPajOpR4u6HW8S7NlvZERASyLX/Rv0RlE6aGGjOvcWwj09
tNmGhKSrx05dALbR6yzo+gtUOsAQ/Eq/86bmDrn6TdvpdJWJgO/ysF6DHrRZHZqw
fMDmCjlbWgqkV7NfAGcz6P6TsLgLBeFzmBiMK6iF2EWxBAPtRhCFjMy/ba45Fox7
YMSGR59Qw2bJzT7RPpTvkf7+KwUIUYII20zK+bOw5iTPqxOe22HxAFMdRiUnTKVT
11yyFe29AZfbfUtyqSt3XiFjbri4yh8beuPQXAIprUZ5utnLr21d7jy5GxWCknzv
Sf7qI8iMWy3uSeiFYrt1rt1NB1AA8ABE/2+00MutXSNPbkJPoe6/Z/zXRaXiBUNA
60qMeljC0xkFQp/wA5OaiMfM6lH36yZ2StT3ySlgnabjAbwNJpqW69ncX9N5dvEg
Zelk/356lBhdDssxXyHQLOlcDy6BC7HIuLsrA4rkLnNWSwjtFuZABdMlSZvSt6VM
08hnIUerOf0qRoS9EXrV9pTe8EcCEO8V8vpfEHeqt9fdXLl4kOPUGNdXG+6lqhp3
RSlfvdeMzNbRwycDJmStUV0SfUYCOtm86AAPvCTW2nq4lP+29lXbDEMqHRiEM5x0
H235knNWosc34MoAscExI3QS0CHbAThwgwfuxhgFu2oLRa5G59OqGwQF4xYfzm8Y
Ae6RknQVmHXpwaguqZ1qLxhgXsuTyE2ZUNjcv+WAxeia3eqNWdUNSRXWvqcoYjW6
EkO5PeB4bnDwCkE/BjJiF3o5qzj411NckigPPRbPuORq9CW8EyoJzr2GM8Ee50LM
/6sAgnu7+jKDdxd+GPL6PiT7HmfTUAtkCgCBoe+dBURTWuWJU0SsueEXQlM3AoYV
YzqVU9xq+E5Kg9AcykJcDjTsmFb+BvzD9y2dJ6ke00phGEeMaeS8DEoaI6lgDCI8
5Tcic1JqE2HD4JydN/VN41oSTk50OL96WxIhKYKK4FhA+7DNVTq/+vSH4pETObC3
oo2vWpSHnL+cQBqL+qZvWDaE8o/UtpIHP6+ZVhtsQ7AwDNPsWdhc6byqR+zfgl5F
9rfTvaMM6MIdGfM3TIpSZ2n94oPLq2xfCTWcglH2/L6gpAvwtvvTWyBxkrtwBfmO
Petyssocn1w0Ev3bsWfGipAnWLpYKZlzjCatpdzOJTV2EPwot2tLAfAyN/8B4cnu
MSOa6vqzQPSpMyo320HpCwKBxtdmMNyaVtXWJgWIKqX7i4Ne0CaMJvBshKGd22Sw
ZGKS/BukID6E831093YSUs8Fs4NpU3aYNXhNiumctVUGIjqDLfPrKk8b7pZ4vrM4
TcTUSe6ULfSjC4hzY390uTeedpNKnJYl5vyosexTc/PefeeMY5l9tFJ1hPY/KIav
9GCLbRQRYBHXQkE9suAD1OlBMhuPrf9EdNsi6vvxNFkVkPYtBHG4F3etzKB+7a/4
L+7x2+7uayMQWg93ks1E2C48Aj6TiG4dh/A/QhprUecnGJ9/qm23PoO/bisbFI50
dhPU104YBxtpJ1J0wnRUJ1dwgkWKIlBPrFMakbk+EczxWCVDpTVVlVyd6YgdA9hL
iRF8RLqqoHZsl/K0mltDUQwr6HMoYP+2qawv9h49T6aHDKzfFlVHW/b6Ej2kiqBH
rF52sdExBx6wIhBVUdMoh9+cYFN4rQ+fjmzz7p3Vk/QtzZD/9dmw99970UD1qD4k
bP/qYuM5pBDAPMPWe1Ivrf78lQSr6Yrhqk75LYTjPFbfyhiJ1gCiw4rc9aW6lkn0
JHTNWIzzLFM9j+WZPoNCynfmB3pGdzjgXtj9VWovwN5ouLK1EjzC50t6IcmQwzVB
Au/+2lmcekf8n3YjsWgnhSHMUCmWSp/mq7IgtWh6AFh8RFVo6oQi2e0Dv+n58sJ2
gYgHPNJxvKKbNE1W0WsjxAitUAHtZ/FoI8wIwrBTbmwiQTOpKET0/eQbE/mr7GFx
WPyJktl2cL/vsEUNoKVU2AHg31wCvq9XwnF0E+p1qaJeToqV0Usb2I85JbdxczTq
mUb/E80uZPU6QetdFaIuypnhAJv3rBNeAg2su55v9drcWixtUHynB282hjq+o8rd
xMIiGwW4b6V0IzkU6JKANhjcsyKWd2CTLzUXg2N55MFjQzHkXPXrwyPN8/xwSsNu
TkVFUrqfAFuRfS+rgybaWV7Cs6yuBj/usLWUK/gk1FqUQxu+Ti0q9fU0LRtVH0hH
j3pMFie4+gkzpYRjMS0KdAY1bOkskUKqwNRGTWpEdbOtH785jZaq5W2E7Ee8GohT
L340Bd4LEQHITpT66jJdZT0pJxu2t4pQWMTDFQLj8Q2X+ga0woMVYKUS/EaRNWgi
nCg3bYvrcM+zG58PEmEiup/rUzuuvoKC7XUpqI/QA1Lri9bqNcNf+TxHssRlNYN7
szuvCdvHrpEIhssxruoMdGnendhJYoHHJtwM213otmaqn980E+YurjLAILzUel9f
ufoMB1R1R5tBdMF5cBUWkI2yoHi6JzKlKJ+9IbnAydzxuS9JAjiQ5ozcqJ1H71qC
7uVZhwBey/BkgLpRqt7GF+E4hOUjNwSZp9d/zMpvKQYN7lfHMGQNEO5/Qgu7X9ax
XcPgi+9Z8P2HhvfaztOGyqBQdi5v30NH/C96Q9fUR/EEZP3d067tPnSmlu3PZIAa
2/6E7FrpzDeLdz6LC0V2kpBXLKk+ILssyqD9rjgZPknRd0i8lb2HBKUhg0u+PW0V
csiIe8BTldPqUIsYrvitQYhiVGxCN6OA6wZLHx0cZaPamP3FgncbkPfoUJKnb03c
fGF6MDulSKRCUu2R5gpgzD7EB2rONqIQnNVNVFA9w6muKWz5zpFVokNFcc17WS0Z
snBS9JbFMwsSSCjr5HSC/lnz72s8YVh75i3QicY/Heph39/k6CilhOsk8vQtiouy
ACc8UcQ3LmLjrQYcwqn7eZ8vC82oA3lm+5qGX6Kj5u91V+zsKr0fNdo12vIaZupV
szNzXR/ScSYFHiLG2KXE8wfTDztkVPDNmdRzmvv11tlECG+u0BJf8o0VXixNl8C2
9aYCGvsiKra4XCMIUEOduuO4XEtRzzpoc3y4YCT7cIg/JZeduPWgKb59f9/IzA4w
A1DyhIzzbIK03a6E3uFEoNBUk5anrI3+kw3AY+eYXDnWxv175YaELGdpSbp/VJhZ
Ab8mLzJtlWJsM7PvBfW5083SDda2/lCUrRintvssBOmz2Bwg/Eg9gD4iT5xpgCwt
r+MEBUGxoxwda+EBOR9zSqF03GAo7rCrl+D4hPeLmQ7Cj8ZCxVIuLd4+u2F51mRT
ForDFv3VpTBz3Zk4PIeJ8wRYSK/oN2BUu+PvdVmy0xUh29TcJrj8IJjuNiPrR6lC
2iI+wsaWFgYp0mnb/bVtx7AYt2hVKaAHXcpWuQX0CdSlwjDrXWwDQf/vqwweHf0V
aPwtcLrajsgPYNiiHGvzS68VMCY3LpQHJKxP1sm5M1zzjjeVNry9/FfS6TezhBtk
VC5rnqbKl+XEvZbJTdy0Ek7sMXF2wgB8uRqVNmeMJxmZZNadh70qG2UUoitDbLCU
7Fnd8dh/0vfpGH2od5qwTv9sRAZIpQEc9azP6fFUVI8kPPyMz5cgmoBBXXTllCAX
Q9o6KYGQvYh6QHe4sNfH2WBz+50PMAi/vMNBuVGzANlfFVGz6kVeyQ9T6ehO1OOC
RlMBgjUuWlhI32idihOXan7p5GYUuzYICdnY1e0hcmVZ0TxPP5Vmdsc2RRMqgb89
asYI8k6Mi3P2dLbn7O8Z2PA4hO6KiIZ9M6U2c+D2koo7LBAnw+h09H+UKava/jI0
bxUw+SgbzaoA1MOGYzz9XiiuLFmzmYpSs7oZv/a88wmZwviCmglUeWP/ooiJXVK7
FnGYng4kDYj8D7KEtFB019l1QyCvqaJMQMVdG9f52vCmYuaS805lpyG+cDFEcwmq
LJPahEiEM53bWrDBRk9Tjf309hkL4jbfdhKdYkDgRRAA36hUV4wZFbA/7o34PW/2
F1IsmZ2X7S6kdwWGMYyN3vMOAlP0dy1BZQJrP7lp0mY+RIEMp/s5NzuUwwm5x72y
DzEF135HfNK1gt1/fG0i/Eb4tIP9s4rss3Anu58i4rbKc5M/bkHevU85lZc/EFr2
KnXtYtlrSsBYf8Ur6/rHvjCS5WYF3aI6syRHDdUM7dlSBr75F8Fts7e3rvFRhVfy
LBi8Pzd0YYX7Go/5qAcHr/vL9tg9VIxwvaSHO252GLUNrqPrjmzyML2BWcsCwrIt
kyaOxpYwDlyIepfrvcF55MDJROTUpkAQtK4wKDBb9OYalssvxbmolfYptkyOQQIL
2VrFauWfxDHsw6m5Z8E1aIOJBkVsuZVSFMshJv7oW6Hia6/GVnw8qdXRsiEojzdb
HWTGP+czYidN4VZgBlS00O+1xBx2h6F6b8RzK0AN0euiuiKc8Yve3B6OhyrcmzuE
MK+GLHcSx2CxxsqQnSUmhtM+mVn8eMmAwU3nQ7/p2tWR4qSPFZVrMZGfVunrJATz
SHmlDcfVFihJdZWwwGkWVTfvnOKBhfFPUpGa5KF2tAm+tnS4QpKjl8FkOZC9Rg6N
ZAhIVShJCL0dOtd+DNuh1QLEXrfl5ZC2it3j2v1vV75ve5m7po3hzjyLZ3T0OkYr
BBKQeIAyO1leGt/LZpDW8TsshIZFHNNVIEBnS90Wp6LAuH4J3shC43MKsfNG66ER
D9vynsQ9ANSJa4EzOyUAExWomhv6KdZKrj7/u5M+UzS05xAaZDwQQ2TXzmQLtldp
9lNANWdM1s1/8dPUYbmzqm+9lmNhilmxSPFTJnKEXy+Dp3O6YWNbH3yWsx4+5shi
t9C/e0m+BKYCNjA7d9hY9OWsNMOYJRIOmz3Ycf2834tr5TbVWBbR24nVoyMwg3uY
YKe6HZHjsWVArd1ydSu8l8s8aq5RkQ6P5DbN3HlQGj05cJRBGc/4TzO0aHSkd+/v
KhcilkBGCKrk/vA3fIlaRB0AHOtHzvWuOcBok7UUzHjJVBpHiBdGjeiTDs0jypTY
6TtDx5pgfCa42xD/xnb0JjDm/DBFYe1kiQn8tjr4Z5gmC8J9yLdE31fWyh2XtDeF
YZH0X38N/fKJZuqH6vUOOgOzUoddqSHmACFgQsYJFixhXqNdscp8tWWcfPf+Q8eC
y1WoPibcq2B1e/RmO5wTO8NApl5Gx9W+KRy1fADCdg+0ERm3volFbyhgK/fdhZtW
0mvxFnj9Asf4M3j8vvMzrrB+ih1xqRvSZnwJLsIZVfNbl0CmxCw2/vJvkyBL9f8L
/X/VFSDiLBHjYuD2GMaMEcHq/IDqQD3IqLvRWPPEWe8lsTMPuECzOlwQ4PKdKKqB
Ql6bXhDKmteW0IYv22F5FpIZ3pwmWiPW2yoLGwO8HpZzdUz4W8Nmo35Dz/YyaMaa
GQGrzMF/aW0HZr0+uAM7XqcL5AhyYwaFUsJxBO/kEwpN0A37wjudKUOCOrkjNojV
8fq4UzQKsmMxqEDHwvNseRSmOAuRzZCNJJdtsdN4wU5RmpvFfuvTEpyz9kd6W+k3
isTKpS9jSN9oM49XDKqWEzRLmOLfYNb8FZKaJdkWF6NpJ6Smw/0dJWErVR6b+Xy2
5S81HMEKYZw3iILjc8mkeh8qBeZHK6/n0IipezKRgSidKD6ocTzJ0d6epYhsHsZU
ra6J39tNwHSn78sey2uR2KAw0YJ+MIfsxAlqWzSeQ67HmilOUqUHxKxPdLMej8RW
Hf+UOzhBOW+oYRYs2N1NkggZDixGUIogCmP03PvE+4xHTu3lMR+AClRzyzh1Oi/2
Q1V+sNKTQu2ACMsc6u6KCtCzYSI/JwjVUbW7UxoshUzlurkzIzE7vzDloqjqBAJD
+eNeRiTcjlNpfbJBnBcDcxdZ6pwYR2bn9NPwzwu8nXyHX5STTFNG1taSTjKUayWB
BItG7bdN+dvPAQfDqltW5itn/+QUzJ8lWt1p6yy006zVcsQ7AUM5Ouv1BoXS5xis
OSi/m0yKO87HnA+b/bhWt0pxokPi47ao2iqx4rK9CJN2Qm6X7yfPFy46LviuO/40
QK15Aes5m7yN7qUmcxxy2yPX4wR6UNH/S7L71NvOMr/8s3ZbdjWa7XGCJCI8pD8h
o3P3+LEG2dS5YHVYeZB+rSjCRDmiA6HMmHA8OrToMxKK67atP46DRs2JvdGUOxVb
JnOfL6jzsxca2sD1TiJq/2Q+ZqnsVQnM/pswG1p9DkIJr7ob/QmnTA2YRqXzweiS
DgyzMMxBEwERn0WRXxgaPSfXyydoLXdxlmX7qOdATvpUimqNkxoQaH6ukQqFLPxW
Ue7cLoaHZKON0Z1kF0tGU+7tTqAF1oU9rKzvJTfBplwVeRC6AAhjsWxu8gVOOP56
l1SW75+Z2Zh3Vj4iRo1+74nJ993ZIDm+6NMKPjUKJYrb6aBMzWiA1O3IxyG44qN7
lnw3jyNpfz9IfDPi7q0dfa8VDiRsDAUFTejdZanWj4pKNFj1765qXB67NbxL3/4j
LWgI8DJ2A4bLVmupvKmX2FNqFEAjARJ5oace2tDqJVZp4QYimcqoEZrfO5MW2/aR
dbqwfLn8D0oNKAzkY5C6/8kZuhhuJFezjgbB/AqbRIAV3kWOrhM1UH50bbN5HgW3
SBFj0vK9yOdgukLAhTjp/saTQWx6Nmw34Aj2qWC+jD9MVffTJU0xQloXrsgJSxJl
R9U6bLrlBeTT6J0abPwzfyU9K6cUyEENV4KUrxoNRo09WG2Qck3LcqQkYE0evtFV
GbaUTFTQkagDOYd8mSr37FUA0F3Z1vECcwLvWp8QpG2JqCfuC3LmAYn5qSVGR1UX
2/xprb+v2lbqlspzyEfQYN/DVdxX8N6myNgbtr2vC9Ni2FyOQKxlmID5Q95tGBiA
0cj0HzgZcQn58GPb4BqgWDjqcpWJneck/89xFs/O5XqvVj+bErVVeCsX/Xv7nJqP
C3vbKa2hepUz9D2WSx7hVFuBBjWE90zuC/lVJ6QY5mwxm7JVDPDNttsTSweoKfIe
tV7uu/qUZEpadNxou6AlKjiA3Qcs+FUwIf6JgQkG/dMBcSPaghDDrctZLeH6o69g
CT4dRg12sBgW65wZJSrzq2RtO/SY+eZ2DxuxGxo5rxa8qB3ID32rdKFMmzGz3M3O
goGMZ7DjG5/1gTOyWKJ0TAMJ85NRjR+NprmgUKjNxiv2ppXd0mCi2oB8h4q34s6P
ytVjdQZxbP+18aDrnqHX3iCaR9X3aYjddNp1m0TVTWtSWGU4IRXMeSIIvNnJBtLQ
yLU/3y9VnextOQhFt2gyoXgige0hkzpgEKx5pcQOqQBZ9D21H9GcOLwclkpG73vn
VrkglQIHOGgczK5ra+awLm4aRqOEwsxCk+NaM0GZNeM+Fho4DUeGzhSqiIS2qb9y
pf6L4dh29Jcz/oCQxnEkFMu7cfaiBb/OayiEKMC4tyTmz1woswJOhQlHUAPVvYFj
B5v98sDgSRGsk6It26q7/jjG4UQAY07I7GRQG9HNUJFbGahzaMMmxC3qY976XC62
HiDs5adU8afqvWOBWFHUFFh6pI46m6e8Mmq2z2PxCyNenAyl5eW6J1HUgsHfAqhM
QW5ms5zLFqRapEYBW9DGX5CTTQb7cz43ZshNBJ7nBbkw9H+vzt/ClPpIMv6K+Wum
oJdnYTa1JUHNkr0qt9GVatqDk35HFgC/aBcg/lvugyJT723uJNFx5yH2jqxMSL7r
IAxig1GEqBGmovYs2lcwCLiwgm67QGZSNKwV0uYjR3Q6wiC3Ok+PWYfgFVh4t6vu
0HBSsfkTv6yODcStBHrHF+m8dVOA+vLa7BkmVwpDRvKY3jktl7uVTriNMXiY0usW
2L6CzZoPdU4S2xuTQUZd6tqBrFcQsg/ogEkVFH4itzufCRq2rs8v/tNey0d+d9TJ
IrufOvMEMfaXQLqHNS8IINdW0If3gY9bPzl+5oSYvD7Q9V58iT0XUmj5BzCZY9Qe
KkZiGMDAGQFTLo7Bk1ASSV0T/hzynnsJNqxnUlUOEqHjZxRHIG0pQ/Lo9V36vmBH
kfCzHmwjoSiOYkEl2tC3owLgjiEjgF5Ez9g1cHp2dYkB1cv98Mi+F3bOOYE2S61W
473cP4DtkqKnPS/WYWmO11SaLN1GqGCHZju8jWqAN/OTg3VLcxTm9mLRlkeEWbmD
Wh4Adhxt1tqnWOLspTu1ZA8R/8Q5ljBsxQ52haKEMB55nLwZnQUoljc3ZyUnS1Xc
LdXeFl8BBaiq/H/wXVvzJgTYG24qu3L67vLGCa4Yp3WYF9EZJpV49mEE4wvoFY5g
6wrqMIIDGnrPxpwANvlvgW6SMf08boPp1KOMETiXCCimjV7Xrla66XEBcmua3fSC
wS/HeOXZC+VqQxn8F1kO8yBqzsD0feCOqIcuxp4fSW/v5muMfKj+v5VCkWbyZab8
+ZizfU4knzlEXm/4lSPZLhak5HSUW1kVaLnIakQkUH6U6co7yI0Bbnzb2J5aynV/
qLnNG21Syy3jW+/7dPbS9FqtqW4uwr0CMXfk4iwBkmtkBrS+T69fRbAQAOee0lyP
0fqw2I/OEDfU3RAmYEUQrOPxKn5A2mJzA+IUpNMN16dENBTh3Qa0b4EqkY8tucVQ
P8pW+RJb9MqFmrjVlH9vkD+jQSMbmrd/RinNqJK0+krhuL2cq42OeST7kUBJV31V
JX0C7Hm7wTtRgqPtdv79P3TuA8Lo1ZC14H0rgOzsjR/BRNpo+hGMRfDeThLImWeu
Q7/MD91YlYhjTSeocoELBfhRkLB7YpUNhWPN3caT9Nn41dLz2KFBeClVNAoFr3kX
756BteXDITt3kLIBHCh5lQemEmZglED2S1k8ojVSLajB8fD/Y7t+BhDyFCc1nVFz
325dz4zz0LwVkKrOqCtNe+XBX62B3dBDkGY115kvtAtLESujyRFCntpQBbpoksEP
8U6hL+RXigvosMfawcffi+GNAO5vasm4/fp7ddhtIVdbYKRMTEWDBK6KevwsPYmu
PLgWx2Ennjh02L6rni+zo510RTj2aDKs8ftmWigxum7QCIpOexM4xvJktJyUZzAN
ABLsGgeRMcGtVYIGXtiu9UsjR/5IyZFWHDpyDHsCkdAwOpmqJdQPtw3kTneKVXzI
4JS/9BBPFOKBs0U120A9361rpHJ+Z7rFZPF5btTEd0JOx5d72iP7VMe2OXEmZ8xu
R+fZEUxzshxa5aMrTjC0zKBVp2t7a+Q57BR1BJDwoeC6mozR0GMxr65OvPBw9X2P
DdKxKFdpkWUXnvi7CYoj5nQCkiw0SPqHYrinQFUx9+jTYKPXr6KuE7u8UkuoFnuC
pngU4Y1i3yZ8RA5AWSnJNvYdTjH5f6MRj+jcmgZX5WT09OUsYoF4I2m8uh4/c2+y
IbH/hGMjmmkN4ImkoStws/q5xGhGb9CqrQTytKKPFoOW4S5tzHu9ZLZf9NfWBYFY
D1IaOwaDrFXTryeAaHo4difHd45b7c3hnTAjVCcx59tqhrn3KTm1M2SU9leTdFNW
Utgf4f5vJ8F6sagtwoMr5MQg5jYHCx+wPwpdEJuj16pz2SuWlZIexfbr+S0G3B76
HDkTLIMxCFd502r6Kxj44tMOEX5X4L0ppDfNFqOp4tyvH6IbCFXfaqjav7si3lWW
S7lzq1U9osyz2BI41NcxhWyoP0pAuN3E6yUg4KhQCmTK9ihr+0Ag3d4tBl6XS/8k
IsC77dxZOAp+xQDeqdfJkoR0sH7qhxyu0Go6GqtkHbCN5cWcgvmDd6pvJdy9Tgax
wTFO/4xG6Y7BHHN/OMsWrG40SAClKCU/jO3FaeNQ79JRV5nnKvxXLwxG9eteZZ05
9OmDorykd4GcQCA7gzo30udKQY7CL0OCVw990nZv5O+tCk5xNf6fZf8jz7pixeq/
nfjUDs4cn4Fwti0TE4EDmaEI/donWTAph75bLl3FI1Ft1Ln3xJ+OMq5s+/iyNdZr
VGZuC2jokPCB7BSKXrhzYz8mFUVlOftXgK4b+AB3Eusa1NK26TevvtVYpD/nR0rn
mDh6zopj8kY2rmF+Gg5L5JdeMPPRUogVRU2fSKGSzJ4Gb4S6tgXCJ588LWsidRI7
tRvLZzs5NWx8bgbSwnV9WNRei0nAhNJhHzqOPfz+fjcULyo1kc0JsD0BsAKdpJ8M
7SQYdjzZ9mKDf7IFKK+NbII2WsENM96LBiVtH/FCOoOlp2WmkcvXlzfmn6IHzE+b
u/x8TiTxu7rB9Yk/c/tceoH7F51gk8D9lEsa5XagTDk/rXMOxDv5Fc98G4k02nHU
4HbbnMcqFulnRYuPQuv5D0R1vd5I+LZ62fuBo72VbH+Ke/qjTwopF0gYL62oqC8d
gtgO0ws+WYgi5UcbnXxP795lXbZjbId4Wn+FUBBjZR+HsnMEF4D7vCawZH2mlZe8
WrIfDUCDUjlwr0MR8MHjg3gHlJOPJnOzwAvLtJyNZKmPTYAcapOjZ2vDiVf+RCCv
OL4BND6zJO1wfSN89Txs5mdPJsoyybzBZ4K7wtXJLhSiKV36lEGyWsMUb4UdN4zl
gu3+2+hlvr+f/sQzbUwOlqRE3uvgbHpkUa/DGyowOUD9CeZgvKIwjhd75AKUoRrr
vciY5vETLXki64xjswBR+drk3zIzso1m8cbDMJKZan51MN0rnZShhXHlPb3MNDqh
oOtg7AUurFzDGHb9T+SefvQbTz5Lk9zeivHxnSVhqzP6Yj8J+tenp3NcsTnEWIlA
YwxtVKZ7cpm0iU2gTgfYiLPCWVsEI/lYiJRkjxj+m69ozARD/kCnGDfOuGR7gFQa
NEMRc2OaPXbxMbsiDdl+csxHjTMriMLYgjpscVyFfZdRK4mIAnIa3lJIzE0U+Z8H
P2CXJYJQnpxjiCkzZdxXSJndSCrOmw0QQTf1bUfXBrUphnPGsVMdt0VOhNd2tGNS
I1CqkskyWZyxj6x4LvXOtaLX9PwODygmuNjDF7RubiuY1ZgFqOWxaCOGxsnQHxNK
dyWbWsjMoB0kLYFbLOchnVxxP92xiAi9oBFGFbLr0gTseit4lCeKbTsfhLKB2uG+
iiLh6pKlbqiL9g6uJ7XmhvJ4KbJGbnIC5H7zwGB6aYW8XszvEsd8AZFaMlzPfD+y
Cb4n3UVVJavVyexKu+eflNwXOHIz4LYU+vfYnZvsHvcq4jKi8dLZR2Bv5joiZjJg
TdTKl2DD205B4TzcWwXql+rqtzcMVeiXym81jtz7dalI84t3pT5TjruuL1Xvr/TC
APdwVVKsjMrntoCX5jiJYq4EdmZxFFYnG3Tm+iVB7bHLJUlTNVuzmki+NfkeoA06
ZXO+2JURTgGTlEy0o9MCE7kMSLQJgIGvOv5XsqnHCrMlpg8Rk1qP7gWXXEEzHqOs
VRZ4uUPxoufrdl+C9H9iIXwOqa+2Z/7wV2Tf/5xTavwhaDjzazNyi74hl6DOBMom
D7evcfBftFDDXV7vMqH2tHhhm8jCo+mcEDeE1VI1Is4pOrnC4D2vF4gKPqUoC2oJ
OJfJqRtngy5u/Fq6LMIKOoF1rraYeBfIQn0teuKR5Z409FQ+/t8YymvCyRbcwekF
JNfuLLF9mWTzyLFtzs6SuBNCAsvGhLmPQBPZUXYQtkK/IGYApjubwl2olgYo3n8J
kLscmZI/EQIHcMdoigs3/sly7BTFCj6Q+G/v8UYovGvqAWYDuXChafd7usNbzueL
v/xTFFC4sX6PFL+g3f4WHlzrHTMwikFmT1Ry3ioelSClJ54X8Whojl7RFk4EoFwT
+/M9PEL/EMuGiqG8W/zE2VRU8HR+hL/+uHWrb+9+qhFBzhqmNUzH6cQrYkGIhCB3
VJ3RHeypx6vXL1NUuUxueq0fD+TNh6GMPN2MgPHuU+Okoo3b0PFUrTbCobBwrLq/
U2KDtrs0GZXKUWUGJZlOD9tyIUp1kWvq99A/dNjRq8Dw634zUhsxOk1tOtz4dDi6
zlRUsA9A1qk7nRKeVOXCYjLHRLoP3IYCh9UqIOzWoEHxGpLUScPtAU0omRymFwXu
2fauTh/Qo1wsWm7N9+ZjpLA0T+X+RLkX8khX4EP5BRhjnoYKIQsSBGRHxhlwG1eG
uDQTv7TbzNvo0XSgvkNXJQ4UnO/5mspHyCf+OAa+2v+nDOXdoVNRn0K7ffWgvo87
+XAoqAl57K8fqEh3D9izha6udMO03Ub1KlmSqfR+J1ItClxVLSoHDyjANTyBTGN5
5HFZxfrK760MvCKPHhCsGIsqxfRQkde9Wsf4YrCoDGNUyBEwhJam0/WGI8ibm3PF
TsOSXW1IwEHktbGmZMxcFsXdJqdkj4zv7gbKrYiEMAkC+3mZnyjEp178duWbPlSR
ZlY7akNqitJV5k2RFwGatsiTNj7m/UtITW9Zzw9vnzF7CbcKK/OPu35ghGM6X+fG
9F7XQmJOQOWfkigF7wiDdaWzfK1BvI05j04dAMMaZx50eQEhtSmuT3wHInlcpTwn
fqf7RZFHITlOUe4f04ec/IBihXJdyykfITNXNHHKtx1nHIQa9X87QFuw9jcP/jgp
v5u7JsCki/MH1a8Gu+ksyYGaGEvKqUWGZ+0elyCcKNAQh1mQGyiPoIHW/R82Qsx8
UTz+36e7kJbvdq9D4GKR3JckUnceS3cAQgzBgjAfclhP/gr+5a2GXUDdkCWft7rS
qCsxHSbIyPTrCmcXsN197BBse8oT2xWcRBL9XLk1WzIOpoJ+tV+gt2sV7ymyeDEM
Y90/bI/pHxhxF6s4uUSv0jick14CRlQu8SCt3Qh/sWaBSZ2vJnFa9UuSTT6E/Ngt
YonXR6QMpHBZrLUpnmHqO4zkyPTKHH5A0Johcu+Od4AwfCEM+AdRjBlRkUNrvZVc
Wibzuxpp3KF2UQ6+Sx2QU7SLjvMyxMqIb4C8dPxDq97qqPMlwEDoDFiVXgBR9h4v
UOUMi93GVOC4fKkneVS2nwkLu82B+9ZE5ZkATF9iAK2jvAcxT7znYSAPmDGvnGkt
CdIuwVLitJbZYo7srbGcksLGPFugeARxjUXanY9oGjb1NzqHla9lYKrC+uBL10kG
gjHlyL5bs620waKjPWwx9+OCzh1x91BWyI6rOtj5XldjeL5CnnYjwDcbOpQw1WM6
wpgendwecSp4PDikKPjaoTwq/a4gOE4LDFaU9iByB8s/gY3HJoY/qIlJu3Y5Z74Y
QELiFpdwSmNXk8m+sL8lXwALtQDyppI1RMX0BzZxzOXE6gUv4gY374rivYbiZlBv
/CLBRCCTR7EuD2oAR3IowetNLZIjghhwjrHnLA9IdDHrQSPmc3u4zCUX0pXCwolx
18qVUuMbh0K+2mosJhXxmIeyGMaN60UQS5Do/sx3rBm8+T+QbwXVtikrYI9jyHMo
vJY/p5GDUJ3TcMW5zG4AKBscBJmaJlLOHD0c01G9mFcyYFBYxeRezQxymBB26o9b
3bWm4kLAeFaQaRyxanK31H3njrXfJ19kSe0keodtAykMFKnKlQLTcZkHnJkHXcy5
08tPJgvyPbZQfPpEVwKhyvu/sal16tSCGpCOuc3EvbPXg+rrTsETOYCRQ2iLjdIf
+qZWwMEpDDvge1AB+TMIxiOhI80Jbc1LcfAlnFgOsFLRWxMQt37uxbgOdYk3V9et
pBlSqP7g9Ko6o2H9WkTb8SBn2QyholGATSqIDfDuLvvAPPFFOR+ClD/SdVBKtz+N
WGA2JGMN0rMW78WXaRB6BwuwKi+ArTthQme5COhvR1BC+shFSPGVvUfs2d3a3ZLY
+vssC2sxfie/eNOJigdXuCGHFbEwGx0crEPSs8RRzsAGBdcCeFMskPBei+22sGVM
s+k1ACZ3SVNyEwIxcahHy3l0y8XkT2k1VZTHHZQv6WbfmysrZMtzNnDSd8N4e1CJ
eob+XiLdPDSifycPpxTO+2HvQjwPUJFGrRUQZFaOdd/AVhtqArPkQkkfWgvF8ZVE
0MmQfCX37e0++xXSwTBOsx41zWtrhYfsKHB8A50MZSslJdCTG666w2p/fnfSuOBR
V2m9veHzmIlzS9TAY1Vloh7b84Yfps7ohpfsFmL1pjszTP62XFVXGFms06LpbCBH
gQT9If6WndtwQ5WZaRdqZY8Z8zKrtg/xKgBZjCunG64gZFcvnXMfT9rTkhIqCgoC
rKu1LwOva4+8R0DTIZACwYi/OD2Q403MyFB9pvEOZOtVKQDxGEiolNsAd9x0esBA
oMGjz3lVbWkQBRH0GdzFsQacexpPekcghwctt+7g+lMl2HXshGqmyNMq23ZfoCQu
4HwJ9KFWbxSt+UQQDiKuswzNlBFID/++WGYrtl6DNWhDqqkqR5sybIxcB1flAxhf
7J0nJl+2Ui+if7dxJ9sQu4N+LV0YU/f12K57FjVwiwzM+jrUN6zUOOHAj0n56bFz
keG1xf5cx6E4E9p05w6Jq8sD9lE/TR1fSUYCygIEg/HsJ6VERiT5R81XwYrpQ69s
+t9AeLNV+meXnI4X19aZ+EmZPMp4VD20B9CiGLszy3jlpnSCTZhTC5HpCBszL1s/
3TUXFsBKxOZGhOFQghzujWrxJ1ARQZcce36WZppOHibmffEttZC31vGuHNCW5L2V
cgqTMa8bYgo8OSiSsj7APIiBVZJuCICoDnrLuanFuXwRMDRRjkMWq0MqHRSJFr1N
gDEkLLBqleCAqeATF/qimZye8gD/7VQrSiUmnPTrMpT+18qpfzhnb2IhYlYdrT1e
XwLnA/YquaULtiueGjZ5epfJXTB3uio9IsT4xqt+DyvGvl2Qeu5EV9T7qywFKZ/z
48RuZK9gAU5ezPV5LlmnpfNeHSQJ2goCzcFBVTrrHtTV0Pm6twDujd8h9Cn8EVsM
uOQOVCiMNSrPOlCluFIR3RlAe8e33C6ackuMLc2USp70Sg6awRf5fCOcor3aJAjH
y2lUkNBH7jRC52cPJ/1EHvXnO4RmYDItZ63o/oXQu2sblCqDKWfLh78ldbXChjwt
R9OREFksw2ZEIcs6wYXgxCwZt9VON0guQaFmVQfoAvrNWCB7IgemsQU+OebXYhMQ
7EEy1kYr9y44mLTUJJGrteV+N2b+ItfqsuvObyW+bpdU57+D2tqU0osQjfe6+7rm
FE2upgys0SKfia+xin+fK7Mqa6Eq5pnNQdy79a2VHBWBLchCyb+oe+wxhIvDYJfK
wqZ4hEseIkEhWtd32noEJx4UN+db94ZqGD/SOLJvO/8GvVqfsQA7GmyjeYoUPvN0
3H8fNCG5FPeU/jRdH1jLkIf3Cyzbhga7Accwhw5NVKA/8VAOY3LfnWSh/9x1VaiL
CppOxcwlFoYsKpg5Xr/8S9gVVtdrHyuac10y86YqS0QRDz1VzfdFcQTisEH4Y597
5wUF5EFkUTv4k68BaPDo/fK2QaHIKchVe8dALAd6sBeVxINfsPfsdZOg9BeIJDjE
9ylwarLCFIATXaIKOsEcrlHikv0sSwzv2IP1BBnt4Scb19xmH8SCa9VqGVTMq69y
3krRcHXb2tgJEw4V60d8rzfDk5Fb/za4/RvHa8ku59EJ0er0nBmxBiCa+kRuC89z
Smo1rKLpUSEWu8ui+aTmbfaH1tmSU7kQhhAQ4qYRYsftRjiavEwOiLTOPXxObka/
A5Y+qEzkHyA6pVtnaa5nkmvJipLVPOKKYhxoK8Gn/Q8VliLctz6xO/bldU9obWFd
BYAuc+snW6wGW3iZp+8GQv4zXvLrmJlBNy6SteG0vaysE14fhg3WtR3TqA6LMEAE
jpYZvCjkVmHik2NOjFJIJ+mg5U/evsM+ti0oPLbsqYdkOZN8zmaT3SDu4ze2HzQw
apR7XyZHyLpgYaNBfrAZHlWg0w+TZc9yxgb5yElJhJXS5hGiJcEaaDkJ5DENCB9c
JgeDn863B7tQvwBsQu7RDETMYy966kFoBCeXP5+2PMhiu6DD91sglnPpWycTG6LG
DTHToeywTs4oxob+HEiN2ijEmL7DfjflyzRE5UQJ8dx/xBYYnBMJh5PXZZJEcDk0
iZVruUr28YrquhXpeVmInczzlhcTpSsmHD8HminFramOq4zC7iKXZa4/DIlypJOS
hNZdxx1RYlvl0ZDplsLSqdc+vNtLswDNPjSXGCav03TLes+PhxnAz4H3MsqmTzhn
ZTTSU5WAQUfT+xPsJta/b+WJ+NNb51keirCIFFr+bkEqFDNy+Kx4WIUtnfGJw3FN
t1lnhPWap0csoySpJM3IfH0uPhr4s44wmBz35MFRHpwCruXePwMgVlO5Ogk76yzF
6ovO9s3pN9u41vbtkSXffwtbScR3ETgCNWIVXdw2lplb1R0toYf/f6/hzuZDjWfU
IeX4796kO8lWa/AKG/yrrVZ/BPajXAv7AUp0v3m88xwqB/7x8mvjnrokqNGAdG6X
27f2q9dax4qCF8naYnkVwGsb28LnCaHOrVC0l35uX9ieTGaZCKZDlTj1vuAScpfs
30gQpvb8RtkUu34Mr0TKtZQ+0yMeRMv1V9TzqTO/oAYqxoY2gPmBU8WqDFyGQi07
HsZEC2OSQO4ntXH6utiaPqxL30CqicbxMr1m4/yhs0PBuuEnm6RU8EqAwv7dU0B1
GBY0Z2p2aYePOYWrBgjk+LYn8Z0cp/V5fn7QqJVCtXfjAR1P3F6SCMjIhGsQFUs7
7TseugZrDmtUWggjlbfuKdId+HPkR5d/vb43nIo03r0EQETMvLjRe6LvOxooUok2
KPNT1rwm66Bz+QspymPzzHvT4gbjRjVKh4gmAwWVpmmk+mbcrMmUGsBRFbQPU5Xc
1372lbhZuHTI6gZJmpexxgTyhU2Nz/UznMIFu7kk7nMtHAoKLlllWcYUG/rTepu4
2tgcjJxIIKZMlU2QZDCLpeG1lM7ExX3xco11IAqoB/rBirUHSiH03XPACTX5cssq
Xi6Jhp8ynEwuKBBSUHglJTzZuFUC/CPipXojUUYWCysKvAeenm1/T8PkIJ0N2yC0
9IdmfsL7D+D3fsS2nWXx6NBgj3///Oka+926/1RYmV10wW1WPqKjyQoyJLZaKz9i
MEwUJa2F78ipM3nSgTy08fS8hPclMaoQmq+2lgAQJF76swl97+rj/mN5Qew4tLrL
ytKkoqy+zHWKUaOrJzey07kBU4n9eNRJ5cPECCxCb89PkkD8Ql6kVLJJCeFPIlE9
+Fq4vTzKvXsb97nuw1Vz1S2G4GfoeA79V6xCy4CYqLR7j5Bduf9jNql+GDN1Jb7s
vAXR4SKtv2y9V0JjUC8L4dTjzEcp3hr0uvZqHOGsAFx34bKEJRl+I65ob417dKIK
7jzI53WeNA6P6GihmKzI70EeJ6FLRgGgpBMsofnwRLwrRBfjHufhIjttvhGuqZTE
T8ZOFIOIcI51zibprEASmPuKLVGblQNwsfvVhOWvp2XRDkF0q7eewOalo/kGgufn
Jj3vl5zYykB+yPxjWxgwtL/4MpsFb/uAp95zJx0bFvO2musP6LIqqdCbVJrV2QQD
FdIWiHmEbYxozL5uXtGGt2IVxcWqtFjS74rpQV9PfnStV+tDK6k1nWugspbRTeuQ
AMJxuXivJIDfnL/H3VoLfQPBWCchAtrZKx9xl+aPPUrJJOxFfgoe1kPsATyFxrYo
PefV1l6eH267LFbwf5SOzyoU9cXZx0APKoBfPmedPbEML9wtoNwO6t3Apc/WQBgd
94S7R1v14jbzN/3kUBYGfyxWyn2mAV2EMdVFbDnrQqQKedZhgsqN1IfD9zFkzCtg
DevTTdoCJhcwYF2PojC2A9UzvSGoPZHdFVcjSB30YgabnVdQp98KzBEySgOoiVE+
A028LgjxZPx/i8424hXfnnDupEbJykt6ydSR1Wwxs4xVCNK9oro+1GpWEbb3O1Ba
DmGsJpRwaPaeUE0PcEnqW3Nh27UdMj/NUjRlkrk9nWrqoy84Xz51nkZzmVKKxhav
kpjhE+EEUkrnag6DkFpHP8E2b7N09QW0UvubGtNto7XBw04ojq9nEQdgHYu7uwbc
EVZY8qtZZvQvH+Cqe+fXCVSNhqu4mobb/gvrkC7EjZOYu/bQy+ySOmw7kAVH790L
gjsTCpQgBLynmRFHwviN/z+gWgrOP7b5Uc/2XlgJENkGK4TKT/MP44W17u37N2dH
T6nhOV+Rlrzb3BasfrRXdsEOZ0S5XrG0tMlb6wLUeAFK0mkmJ+zBYAbNb5MSdZ0b
4238WsIoUxJHCP4Qu3BTIACLLXjXjtF+tDqq1uOYbWlB4QtC4aUSZZSbIcHdvUkQ
FBbTgRfoKP+oTNXhRCtauk9Z/bvzFYj7UiSsZmCv2sRBeRrJICPYGcYqbm6WK9dC
PODOvoBsAnYRyXbDCyebJw5X7dx+SbRmROypE5mKKAevWD71py6kinIAjToq4X5n
l15Smy9XdCzohAM8EVKraC9dVPFmGBUv+JSw6XTbII9zd/IQLa2rbUfrgHZWiCyV
gFN/qZDsIQn9BsfuA5ex34/yPN2tOqcgCQJh8UgXa9cKEmOh07aNxHSsq3HIOdRH
GuvwDacOR/ilWGRY1nbCOIgtEYsZkvW2cHHY/Al7qGz6q8CixeaNATI9TBIQPkLU
L8jHiJC5+n2HPcAhuOntfnrCiwAj9oIPpHBA68l0DRdRxORxBwe6mZZSxFB8eadi
5NolgjUxCAAxSjqdGzhn5VJTiXZ0mZqKEA0pSU7YlIs2Rvq8cSaEF3o5x9XqKHG3
BKPMNiVI6MCl8ckhJVRh+9F+M6KUydpIKQHQ67tl5nChUump5XeKBVjBsF6bcCJw
nTPDD5NWb9apTtAvT/NkSsMkk0+C2lTcG+Va2ZnpOerFXoV9gOP4R6b3+NGSmcp2
QWnfTB6p5f34aQncqypAmF4W5P2d0l6cVEj7zVfasyTZ8a5EKNzjus6Xrjcz6tWW
SKTHODta+MnhSBZ+RSd71vRbCvX8Dti6dXApYnj5WA/jPliPgs+UjdkN2cirlQL1
Sk2D69F6imqsAjXdM7t6S/dsxN7aQEIB5gEVt0VzVQLwGbFmsb9dmphVZbzVNurT
dvAmr2O7gfr0g27pH1UVD/dAISG0t8ATnIbqQQd7Pt5lXi6+Spik32YipQPE6VQk
VT+yX4unyRySjz24SXv/5hsgGlnij9WOKQ6DPt3/u0i5Yc6NHvpI8gLrPOdQQJI2
CnXkNmDm0l+ydUCbS27CWJMJCJVkqWoycwETHmihc5ehl6jQsBaNw4CB0XjYNegg
bzj1upN2k9TtGFrfCgOUE2HONsER19SRj6NMc+snEo7Y1aG7FED7XtV0B46viLt+
geuKV9CVRD74Zts0qxR3I6v0jJd1swMjkVQjTV4o/f1cnYvRaKCKhs1FGwK/uKED
uV/wauJdxhPl8laSMZ1XAzeoZsrAhig/55xes5wRU7504uOojrTMiZhC2XhpKAuD
k7cGXooIc3rED8hz342P7Gb6bqpI7G10tkPy1pGD8NddcVLsUWgKUO80xeMHTwu8
+CGQkiF6No1Hn8NeADT7StNNnQaEpjR4ZFQNOamdwnlaCh7/JvRTZ+u4yV39c0wb
jDKVHggtqNTdWg9OfesrUbn4lDMjjnAyme1/BFgNQmDl4S6+MLm4A7H5tylAet6K
/tHLx3RCb56+ohAVn3158CnQzY3rV9CcSVwGIMc4cWXbKjIbPcMJvoMe4UpOAsbY
iJWS0JvcFb8qdOi0w1r1oKaC0HUxrTu4KPB4IW78FdGf1BsNTi4+LT2w1b9e3wP/
RxS464Kyph9ANYi3E/3VqM52jgh1HLMXwemAn0eThdqVexxVDMygFK7CT14iylth
fJKE5QXmoc9rDKHuYwvIi83iw4PB/pU4OZQLJC5zj8qDdGND7kP5huY3w1UMgDjc
Qsp6clgfbuwGJizyP4ttVcLoA/UPkrwWc+zKV+2VGO3zpBYwqWj1Kj1p3azik5LM
uzddTmL/MfcbF3FzPyZHSLwxm7Kg66xFILQbn57/n8Yzj3JumPnIOpt8rC4E+8CN
QCE2i3U2dODs/S9pmPc9XJOGwaf5uqgVAITDbkODWYLTjrksXhT7IROzKO3gyQ9I
yd8aYZ3phnGrOkaS3zvGJ8vLlTGzsBUcNbLwVYEYZLRXCCKo8NM8HuxCEanuq6P4
qui6gEAS4Wd9uYW4tqX3c4VZgrRQmLul2tV8vaOL5tXE1MohGPB14JJwfXCpE3nu
XWsIhAVugVnjreDyuaP9Aj/msB4Bpz6Xod964CIpCl/KB3nOO2/Tt9p4E94FKhX7
VTReJdv5Kcek/QFg5I+UOoTqU431sJa6ruNkjlYYYqoPp5rDiOZ+HeXzKfgvU5KP
dJdeRZM5TfvujhoqothzG4/DtRnUcz8st0dRUXtzDhck6UkqySe1ZdDOcZAyzT5n
Rvc7HIuoqcaaJnTsGuwCBlOgG5i2oCA+L/rUIz486CGNKtQyAAq5Ir2KO/OTdQsG
7sBapDktmYZe+GBxmnjU2aIFs/hlA0IjvDwxWWkXGKrDtoOEC7p9lHacZrELc509
mCXmDNxo+i8Ub21twoYSHbga94TJi2Nqv6Dw/Zy+3GjVWCny0nfpsVx04ZAjQPWp
Ve0kWHiqL3XALBJUyJidlyyrYIslm9MjrwtTRcM4rKn0jiRnFUpC3W4cIpM4ZYqq
4REfAhVY35fKWK661dtXNse25/31GYYGQkJ8Nwasa7AOUerlutdoL561z1bvLUP0
hg2VJXDbibM2mxJz9KvnNZ8RqdhRQiKXybjR6Ak4b2m7X+jZj7Bb/A71wlrsXtWa
6pDlHcZiMqPJkIGrr7MKh+meODN+X2eCneaAaWBNIP6J/3uo9tjKeUDzwFnqSqps
ql3WiRMcQMzYvLIYEtxSa1Mvo1oL//B5RQYaLopRseIl//vilSPC63m6FkXRPaw1
bUeSdyUUbkPn32ENL0dhseeSVB2iHP9ZWGOF8BU//0uXtCnU/gRQrGXggTpcueeV
3eqyBqdVWz1XjcDevroXoX1UvZSaeis2bbxoVemcaelfy0soAcjz4hCJbEAD2UUN
d3sqEZf8g322DaQqvVORgFCUAQsfr+mihk9g6+zbd5bpdymUsy83qHPOtGMu173k
DcFJqZEquWXwX9Votlf6/9xq8Nlpq2AsQN8PszX32BCt3kSi4TMUzrnzW3yna1Tl
K2K8NkRQMmEK7ITJg/Ir3hfo9dvQM6kpDezMg0OQYRILCwdVsmDk4h9sUceG3LHY
YTlCa2gSus7I4EWcqH0dnWmBVWEJro2SA/3Lk9rBLdSb/y7hB6XKgKAkgJZUMwef
oV1QK20Y0R6/yrWTZSOIX/ZAknoG4FjI6lHL+lcEFPQM4fD6qij0b7vje3b0C8wG
Yr4ztwV2S8SO3BVTahXb9TjHy2lPFXZcdmGfZbn8bKjFJ1ndclvnBLw1hJeiSa9X
X1wC76ZBkOea8a+et0vddugqE2b8Ted/9kzZTSobOObHNYH29BZow2tgocfo8tUO
aJLfQAvj7ZsH2FbwdScg09rvQ+wx8iX4iu/FB8vKAQdaxIKRPnXUSxtLdoRhwSyu
pUhJT4Xf81brNDapObMvbYJupp61U5h57pZyHCeN4Vhs420wuDSOAlNFRRwgRGQK
cd+IxH6Vw08+Nbc8AJo3bDidR1d7mQi0Mp218kQHcMv7ayjnKpzcyhqgnEMx0Fn3
wDHtinOlo0IZTEOSUfT8Wu4xmad4O9KEWPJiy03Ba3H5WEOKUJhl/epEGNPOBfvN
aRXT0u7cuu/GWx6fPDNXWaGx/VwTMO8sMfUAwYzI9zO7ZCaAy7bxqSC9a2KsWwFe
AAP8qBHpgKTdRnKfnzMugHrqnc5hLdmTJzyzs31y4PgXQ4ib4M3/wHs5865UvFMJ
pDd1WmNf+MNby1/ow3LfePhz0k+7TOfV49pPNvVVfOBVWA5ylOAVya4kD0DMofiT
nvO5/2T+Wuh+DRZy5vl/OKmmImlDCBi4Zc0OP2sNENSuA3IniOcaQUtvVFA6mgPs
tpUtZuzNuxQoe+u2J4QviXYA0Tn4aBqMKCN5XlJDMJz50Lhdg4PqlM57qzraA3JB
u+Qzh+QbiprMdVqZL72upOmXHexZyFZpw1pRde+6svVJzisRLSuRUwPSog1IkJuN
JIoNEB8p3jG+u47NjbHq+bA5GHXKxotdPGWCrpUQsP57TN8NQe015p+y6UH5bIqd
pBDy6EFyiIDpIyV5HE7q5v3p42XUIe7F0UDJ7aRnlZ1bE6usyclq+tRKxdF1qfRo
iTEBCejYxg+5U0YvB44omNIkT2IXINKw8jh+wX7ms8nJIMzjVaDwTMvRvdu/H0y8
C0sOJM62UvKlfhCy92VRRH4Nh9Js4T1xPagbvAJ0n+RGvoB2EL9f/m6NLQgTvn5H
lM0edjGeaglO9ofEto7XYsKcdfH47AcHFpiLRn9tTpx+6OaqNN7PBuN1IPPhFcQD
aCAqbIWGtNINvtf61iTV29YYVcnEbqvV3B42VwTjSDas27XZgKhaFNT4YHTMlGH/
9I737I/4ypEbLZDvr+xPyVRR5nLXG6vgYsK5I6w7vk4hFyf5X+rzwiG08N24M65s
hjjdu4pnXS8R8zchDxH4Vdnmpvc51dwF6kbuuBeuF2OvrJUmIBeiaBJf2nOZ04AY
1gUikLr1AfJ80KfzAhCfHBjK9oUiGXjKKEigSv65xZIHPA7YseTrQIak5f4JHDW4
Zk0P6v47GE6zc1EhUZeRwJuC77qm+apI9DyyuVtWibY8l/hoJy3Fuc9qq8HTFxff
7uk+BrZvJf/xyH/mWaxxMVoZSwH54GgMx5cW6InFRhozQL/dH2Nb5NoafPs3SqLA
1HbVRwxlAFg1/SUkFWBPG0IeuEDNvMW78uwCxaL15vc2IJStiTwYBaQiWPrfyhkl
z+stp0q6rjQf/j83uLOTVJNY26iPkMdwod/pATj+Hq7H6gMIugJucQGj7vi9mLvN
jkt7VhrjqVC3J/YBw2z2u03BILQE8g0BlOZXAAAjPQHCh3csqp+FcXsh2hBI6tWE
bN4VzbQhZye6X4CubJ+Ar0oTbj4hU/Ug7F2Yz2QjNN87NH18rAJZ79GgzdUa968L
ge8Byx5nu/dTIk9haQ+tSp+7+SAEKfXemaWJCW88T6E7lo/yeirPyP5Co8daGIeC
eQOvZi6evcwTXMkDSNxEGJvWUZ9ZXjqkpc7chxezxlxdvm/KtYX3caCvF7zo24G2
hpqtXtSE22mGCp7+Vjeda6OjgtW+UHS7sEOLyXNwYQ/oKtVKOH5rrEoRUMmuWNTd
UoLnvTlR/8vnBQ+KAXAkMBq9i2/Fwec+XSHewXMvFCi9WxSkOSUbiCUvlN+9kKtS
eaiTbWzzte4eCMm5aRv0w8EGPys4gvM14YEguP0+wfWJ0G5NYSJYZAbNKsz7Zinq
OxkqN4uptvAYu/emp9gDvYP3cIM7uIdtfFGmTh2MWDC3+YejLoO6hPUEPj016R7G
kdQT6dZJgD4SRtqSlYCfkn1nA3uYRHLmDP0YihdW10snolSf69KKJSGEgWugy+nP
X8lvXHc6yS0BYIm89v9CQxRFvGxztHRSTPKTDQb/R3mlYwp0NRr4VgHNqcHZe7/T
02/M6ZCAabdb1ETfzuucjUM3ru+ksqazHLfoLax0wB0QVEq+WC1GbP9wZbm1bVuX
sQvbA6ZN1I1vok7k1VxCN/kfP5T9UzGDaGMea/Woex8BH6T9JLq0mwBNY3hDGHc0
a/4S9Wo0Tb+AUCjnQrePmfgYyXw/46Uzq85DE4zWpwDumHQbpvTj0l14L8UCeK26
lSVhh48gRxERTF6q1XPN8FxjfIYiGju9zIs9sNTu2TuwS2HACy2YT8bNZqeZHz0g
y0kap0qCYpOCK+yAvuSbf3v11xMWMbUVQQv/SENpZOjqVVjleeNtJShA7wOZ8a6j
nPHG1lXqAM82eJ4B/r8dykNdnNjhBN+blnoKGoYMOgKotVXzyYe7utXtD0xCPzZo
Lc4ObncZpn+ZfI6XeXwc+QhWULJUcPARhDhotPaxdgcPumPusHkBZoV8f9DgUz/w
kvtZhIJ+IjIP5wNwVmEhxLptixv5JHdYq29H3x7SEb+2a+IWqY4cUOf+0hqEH61j
dwDi/Ul24L/BjhpANa4bFlgK4y57jhS3cLtQs5fPylSzjj/pvufm7MxAr8qLiSmH
Lf7F95HUuzJxGTg5muS7jvI0jOBTK3EtXMXINw+GuOpOXRHoX8NuqSE31WpCynB9
YosrlL+oImJSXmlCKZGLwkPRaa12UUcgIxJPw+dT7f1mW8lC1jjK2bsL92XNyX+X
GWjj7QLRsVoLrSKCJEb/NApD7XKUNLunrZJ+PQBGeGggrxyi1rJUa7MepHJKP02M
r5/XJw1P6/ob/s+cXGxqlM3uNKj7oWl4KXVh+XL4qL45XO3G3CODFoyTjN/0wPT0
u9QQVq23qRUzP0GA280DYjUOaI8ed9HE/EOA+DRVDYMCCWN6mAlSnzLumm3SIrdL
cinN7sBVC7GEQIQstGDy/GgyBA1nZAOW95Jae6gFeHoG8alO1grwZu+3SOS7fyuJ
SNaXy4ODYaDUBBZfUst11mxCCMIQTENXKhzhVUE95WgIhpGDgSrKzzAfp3gS2RpM
SlR6306x4jcokfCTwVzJ97RNp0iBrAbCv2pWaVkPCSNASeedwhNckZq6vKs4futr
DuGdE/JsplD2Gw3LFZCogfGR//+KE2+HHOBQNNEsOlVdT87guJq5xEMWr8lTfK9H
GPYzZP9AFHTc6IoZNpx5AI1gcrCvrraUwxpIt7jJhxVPsfPg6Oy+3F0hwPagzXOa
hV4eVVqum/745SEVjXh/VHJAO0a5CpzoeRSostiDm+Fsk5eVmlNmKEKVIwTMgMXT
6nr4TceJmlm8h0oIMyrYyLXqqUcpNByvAfc2tKZlJI2gTT6JfMHHurKszsnG2h+l
z7PtPetX3FWAdewB3D3RbVx6A1dQZM5fZAyqLO8dP6LFVe9j71p3kG3ZGjTVlsT7
zu0eVNVKABmbb/8yBIw+BIfwly+i9ynufx3njiUTIwe1mOC6rfJWZsV2WtGP/4aC
r+8ksK5BVveQyBvM621JtbA/qReLnaLfTkzqwSKKKzykrJudsGzKv95c1VrENM1S
U0qb1fdPJkiHTtdE7hcgQEdDYL+Q/FSULQFS8W1BFMGumpAgcXkPOROk33G6Rt9F
cjT4g2i926AmthmXaMpVlthGU+XRcKGmJtr2sSVmvTTQk2N0TWhdmwaQI+H976d9
8S4SCJGADG54hxfj589nCQgZVEJi86yaRXRRBePO5/RLhG3LKkba3yLdfRZJBZSR
qfGhpnHFPn+y0f51G0qIahzbxF9nHgj21x/tf6NzBVdf82OI8q/s4aZlGXzUvQBe
BZqEpx3OA+z6Hw1poY/ad0eL0C5+BCqhFqKr/nYKRKyc13r19sV8I2eA76FnFE59
6E7NoAinEB+aKsjfiaNX/QeueT4Q6oXWysN4+/Wx2Cbx3frGbMKqOrhArwE84GWO
DJCj11AM8XtSRs4Um3XpmgkrLzWuzc396Axk3vftZuaUCNjnGdoHrJWCF/ldFDPg
AP+fFTmCa3C2VPyXyGGujhS51Tbt1D4st+FrNLPT91StdEkouHv8M/TGdZwNv2Q2
yJbA/xJJIscfltgXu7jLcz90L+jRNNNTYwYcAIhou/jvRfod8aclmYw6BieCVkux
GQ+pkaEt9KXRj2aQKP+GvL/5Z127eSQ3KaBo5fZDUh8IckBxhz+akZbZIcRVmuCg
KIAwnf2AN8e6ZivtytGFROys8ROzPDCNoQsxd+eyJnYKT4oAvWOWvOeyQCKfrxJ3
7do/+H28qf5D8BfWSH9ZnAdvZeMsyKzx9k9X+EiFTdE2EYhcqqrP8fbLJQ4AQVzY
6Nl5x+Tm3ZhQTZ1K0G0CvUma+jdM+WDKr3JnvZN/cFvVwi/Y/eqwhvkJiUDr8Xcx
1l9/pmwkUuPw/nDvAs7dz0r0jPMLRqefHzKiwFm1dknCfgjhrJpzXAMeIPKZUuAD
Q5d6jcAy6PujXZgHZbx+a4dZWcTwTJcwVTiz0JO1mfMwYBMCOk4wGszMbiuIxJAB
FAW1OU+YvenT8GbUg8aClFe5DcgLMjb3oKrw7bjgGcyeajkW6vC4J67MX90VQGgU
n2rWQAzQhwKq9bl9+D4Fw1gHMvT3wUWffiBnVNegYQF5XBkcNx19nq08O9YL50Vf
yw9x9EQbd3S2YqMeWFy4cti/BSDrZ03v6CWns0SBNxrv7wnPMoyDcTWiZz2sUM5N
7cBzJaDLPFMaV4eDKHQq+bVZYiC8n/9zp+fpnM7rCXA0CZi8xGKIpUYPHqUZaObx
chWusKQJCvl6USZSZ45DYr5ae+k7lPDgRYj4+0HJqsGtW9BvaY2RkfMoqvT9GXvL
lC/DjxHdjP4MpSukZmG7u4yi/ODcr2qUJT1x+SQTOklNi2WOG+4j2AjG5RbcK8ed
jLzE63tTqCWoWMA5IPPBvwDD6TZTI8YtTYwLJkdJkbtWli/SpAJ4i2N/A/n5y9As
kccZWFdQCEk4aQU9rxJ7BMXED+bl3RA2QdoKW6y9V/UbcONmGM8aN9hXomPBtVp1
2xxmXH0eqQMzAByxvHcIlnbaKyLxjZ1PMlVSYNjziYJ5+GM3QamgJoMB4Pjdq6kF
QumnsdC9PqCdWJu7h/kuInRrJkYwJh42rbx6aE64KePedLprN+m8mCqk76PWOqG1
6G8AySg6su3IXCxck6j84duG/mt7CcjI07P+4MW1IAWDIkU9m8SBnWcuVvTMsd3B
nKhrDFcr5NmG362QGeg1UBzVr9wilZ/fIF3zRUTBb8Avf15KP+0Jp19kI1C41LWx
qXQsay6J0Us5Tj60qKXVA/7Xr4EJbrFpJ6z5oRS4csv66km9d/0zmaXjQk46wsRL
WEOR6VYrPnkD3Lp5irByjQiWdr39IBMytX8plzsq2wZs+7unS96R50tNSc/yYLgi
DaQJtL1El3eg037up+8+o0Lo/As3kAibteDqKyyhAZkJy4v23JmQX3xYoqnseDM+
KAWzCv3TxsO+ZWBg474hwANHRQXIyy27ScXFgw5fVUwzXuTXqi3+MVzWDq8YWR8E
Fyq0cLHi8dggm9AVdMjDQJJKnrqJecNUkaCfrWL09eLl8TBPpGVb/XxhROeaVNm+
O1TuewQIW5S/CoIuGSYOR5J5eqDqmU4KKc1r1wytSABd3oTlzwlY0aKHTxwjyXAN
eQ1rmf5FKtmlG0Qli+9bil9jU0lFk8iUDFBtC0DJEagiDhUmpayN8wUa9xaHw8t/
iaU5bJir0I94NG4x8d2KjnuC6mc/jLDeOBx8boSR8KssNqI6T+1EioVDAlyu8yK+
igR4pXJPnUQnI4IG5wOONxkhzIdxzT8kYT/b6QQALUduxlxWXDoacz4BFg+X1sHh
smmmg0AZXScDMSXoRV++LiyuBhG8mrr+7k6R75X9VLDDtO/ElghlLWDPtV6F3PXH
fSN1aFAKCt7KHIBZcuKyMa+CLu7JqSw8w6Mjj38QWhFxdoWY3RqJmhJmaLBKmIY9
cAYm/zoS9R2L4ABrTcvFI7tYIsaQcfuv4PBG6bGeCV9ZJ3nGFqvtq138Ea9KRVOj
/BlFIADWOY6XG9vvyC4Y2PE7egaJ5VJdJOOglIU+lv77gkcCAiv415uOdTJZd0vD
4iySK8QF1LX1l8CzOrPj28BcP3CtMDqheiPyqm/mIS1dqYeNHK+DhnIT5eAJvAFw
wL610mYzpMRnfSKezrzxkjqZelthVHa1oAPvaJh2kAGhI61551YJprygLV90XWQm
8lN3w1a9baNjPER+f0Gldo9Wu6UFtIZ6icdiB4yLOoc974wZWH8qVy5ZRZdeVDUw
BGLfqP+4ozXWtWPckwb+0rQ4ABoQuDIGiY7i1va6suo4+9C51W+fS5RilQLow4of
5J8BOz7KFUKPR25Ou5u0fksjdg/FPsFvThuzliC4g6f0PpeCUwZNZSf1m6VVuMuF
X11AAtioQ9L6xzoATbcWteEbV8+lEm8HYBvPyEiw2Z0A7kAshYFYsNRTwSL5WxCK
Kc8MlQyBRa3tBCNeTeqkL6GxMGZIVUeKaH1rZN8Zb+pH393ak+re1g5JC+qdUrTk
wqz5ym7WrkGafDxueTPVbxCdisuvt8Nx5P0UjDW7BqDrbGDfQSq5hcAecJkMf5lz
+P6UuTmNVuLUdYckAqRKnnBu26nR7UofnzkFPzBSz87WZhkW/5HdPxFVU7IFcx80
ntJib+KuO2IVV1icUiU4YCKm4UL4g5OBjhzSgXbke8UhSp2+P3rnSQlQqhDpAV6j
KvKQV2oBAE2lMZYgMQCLTXRrPOLYlphP5KKzgQ+c4TK0YVEv0f9rfvRMGCAuA8bR
iIdixazxNXKjUEpqtgzyCR9S8g8J78gzvToVv1mLNPsF6TO68t/yWx9FkbK9U4rh
+ArcuQ3V5D+cp+GjwbqWvWBs4gRQNu0T6GUerah7LGdHEIhu8jEatcJs0Nz0+Drh
7tTNZ9oJaMtRXsdHjkB9PvnSMxYanNLUpL0PEo2j2AOUPVDfluxuWUaH1HJMpwek
GRmrqLx4fKh7lXoFMpWYtZL0eqQk9AQN/0jFgrjSefFX9vufj80JVKR2qENJvK6o
82IT4l2AqoEQDT426sXIw/0ZSwPy20vRvwxA36WRKefa4DHr7Hs3r5HSKjKmwJp2
3143Ah9OowZO9C/UT3tUcy8dZEyE5Sp3/RlFz3z5Ynwo4LPsyrP5yXPbSUM7a56A
67m82X7JAh7SpQ6zqJGuqpvkLZeuxLCRzDxEnVBKIs2SRYn4tEAQoMydGuwo5sho
dcpjUoafYoJ+QePQjMKl7ua4Ds1EfZ3MSeXHr2Ne15ptXYKQPF55vdS/PKQYD7Gl
KH/NSltcviGltnrIdN+2elWyUE2tGDizUgQU3k36BW977ru7ghDr3VzFAU8uGzzN
pn0x/2YynZABXGAYbuyuvbWNSi6yALul8dNBrM4b726sOdR+9thK1kRn6lHgxYQV
WDatGXCf/oL7+poJ/VTypJkWEunSPYz7vV3wJEzW4Pxx6Pc5y5W3kgDsqO5f7wns
WFzOLcN6LYtbg86SsupfZE+sUgJjXN0a8y/oER1/liGbqyRdJQNZYpRE5U/vchbj
qjXLStfi1vfNQoMu3aupl4Tmggsicx9Ad+Qa2QS0EMVyj4n7wP6duoi8jHMe6NOf
BnFaawv+7RvWkWjI9wb8eXxFZ3JI/FEnvwtTdEGMW/NERHdgvqYxhlBZEg7EBMRY
ho8G2gSOLlyr+73kNIyDY+Lg2bm7HN9ITCJj/B9VON98k6yEmirJJlNUZdAy3DQC
aQjVuANNq9q1jafMybz9eY5k7uaHqQuv2A4e0H+8ZmuvsJJanhlF73o8eM/W2Aj7
y/U2YDwWDLXbyq4NrUgH48ZpxtvmRfodA+dUVQ8H45Ifz+KK8Qh558tf9oI1nJkS
RAWfHDRNEBdQST4hc+aVQWpYf4yA39iC9LNSZQLO+oKTzWBcxTWqcpIJJrtypPPk
vFJL1DFX46+iqeQuikjOwV/VGFY0FEJGDn4G8Mdwn04t40Wg2BJhz+zuGjUMkGO9
i2Fd/OxW95c+mDJPHvBxI1aJZKv0OMTz0pqeff3EuXO2UtkCmLt69Gb1LmoR3foO
XTlNjy6GMLduKzk0mkcTg9YOUG6aL02v2JUHr3KEmP+pFCtGxPsFYXDCiR3mSuLH
1pMBBHfA4pjnZE6dHimXvdmZ00Dw8/+rCeG2JrQnMaVAHWwaVdQXI1Hd8lZ6DwKV
uuSMXU783JfwbulgI2+tQNyxinMIOByJWxUOGiT/16GqcEbmPGd10wtnjJaXP4GE
sKTkpCk0jR1WRPCZcgqNUcZOCfDNOeKJG4Uuiz+4IzdpiXtVZR3tg3gkORSzh1OD
F/RVygU0kpk4SSOeLSXKBLTkMIyBO02EQmQz3X0mZ1d4O3eNrNNKqKMq4a162w7d
mT7wL3eRsvre9LAsqnYxeYHb5kCYPYPvnsylqU6zFIAlguSz5igbO/Dq2NAenl6C
elOg9e0d4pgmjF61uz6QEVmVkUc5Ofi80xEcOY7JCpDxjxGsZRie+2jIBRsMFXqc
5vjL8Fu632V9Pw7if258zXqI4TpMsT+Xqzyrnvutor2szT9N2VafyNqiC059WRI9
ShOb4s1hVrABBQWekECk3C5E5175tkT2VYTpfR25hA0It0XZmiJpm8VMllMTh+y8
MpkDHIS6DuafaOCjlAftW0B0jxDXTn3ue8dSiKn4UxQAFF1JOv53d6JMwMK38beR
HPlipD/G02Kg30DGHjUQWztL7SRjIrcuA8fFa0k0Sbp5tFt7n5ZqQM8Kd3eUgzsV
eTA+wnLJK0PQCW1Byt2jwpMutTFwxJMVaTkJzVgEiwu54I9onh8+BVdfD+/imPtn
6/uZbhTiiPDUfQvLqN9MCXr/1Q6HD3t+SoglnJ8ll0RnWhogtNTJC/28BQ5j35Uy
UxoEa+SMpabjQkEcIklJdexrQgfMQZ+J9OkTKu37BJoV3ptqT2JWMJ91B1ZEpQwQ
xJhJ3dGBNSynLv2YJUZn38eG9GuvajdhJ3PwlCCFuX/gzMrbYaFyNfT+IdtuCDFb
fxyiiuhLgvxN3XQNSBKmesIPSBl2X3Dk36cyAS8QXhnnP2tf/RBqzOmN2xbr1see
TDrxtQassch49Lv4cYW760pzygEYSe/6CiTScuq1S4SCYl0IMe0CS1GRaZpcHF/9
AyfT0mUA1kkrvlVc0ltnSi0E6SQ8DLOM/nyxqmhL0VuliiOpbWk8R/l8enn8/6ab
A8o5XpvWcGP+zJUJJ9vxuAXRDsVTWC29DTLtO7iovtwrRnry2bcb47atDJgnnOqP
KM5HqqUKYQklIYDjIwskxRIV8eSxQ0HgdhXnsNR8F0hPeU2LvzivfnT9o74AQlri
VTAQr4j0Y5QaNZKV7RGf81N3OXba0XTY0oebV35ZZoAO2izx7GCVXNU7/jt0azVm
Q0eZb+GJAw5rP0kUXENr/1jbbkduaQMSxI694BhvLRF1xtQhRVZ45y1Cf94BPWKC
cyTuuWzwtAcknPxvVjakify+gFX+Bgr9IP5Z69A+UqNQAvmZqh9zzTjSFBjl6MJo
fHAWx5883UYxyeCG1E7IGECNA6Yrjco2bkwYf4fzzmwniHfpmpIWywShvJcdgkhQ
aSuxWi04kvd/OoOwzydJ0ViWjvXCv6qmys6JKU5BjprdqsYvZ7gXb/az0z2sM4nB
bYpMoFYRbS9AEiZfJpwvM40zwkV41H11MeBiP6ZqYBbZtJlQGZoWi4dmhpsT7IF5
MNvakyvuk06O3rRyZgopz7wDYQxan27M+cyznb6LNmH2UPNhNMQx+tnUa7FCRxEa
8OvWKxRbOoJvBpzIG4MjXoYLI/4TZKvYqmKS3F4/Rk2MNdfptkHnJW8UArdJVW6g
mmMfg2yVGmAdX4edF+XcKLkx8w0wWNvFe9Y2EDU7xf92FrB+LtZYV2BW6KPvILV9
Lllj2NT6G2OPRGjqIOD6y/gkEmwx7LDcyQaBR8OlDtLxZ5bYCi5MdXV3uHrVFOre
Ijsk1/Sh1/il09cDzBonX0/0/UlIEw+fxvycNvpSSpldiPl3M2xudy9xXg5dIIyc
D5zcDpVFvYvxUrHBM3PZTgdKgGRgWaGRAIKI9xOY+TqClkvAWhNr2UzaeHk0ZXVz
FSZyXiQIhLVyFIIxiQz02v1cG1dsNB8QJ0sMmkImNA2gwVgrU0E8StQpzQRKYYRS
/lDSDPvZsJPT+NE0Z3Omf7BagPW2edp4zJjTI4HCWPw2wfGgsxhW5xoC98Htsp8P
3nRa+Kr0aGxw2ML6tsr8gA1dHhFn0aY6sUUGIzGy5jeyoIFY706DCe4pqd8AAO0s
slHbN84ZZLPgPG0LGtoZwDR6pXD/xvENbyvag+r8GA2ahEjnr16F9Dz13PlDuUo9
D82gIZbLRXUod0NIZDaZiGSE26KwcPqoO9uZZbV+SmFJ6U8nYzhIWsyqhQnRk4ib
SVFBbB/tYIwD39isys9FuMVi8vChPv82kzSz9m67roEjgQrjSIxed+/I6KYCKiZ4
pPqvDZf1L6IC4utlst8axQiLU3pRKJ5kKVZNccs5hj2fItwq5/aeK+fUWEkpIZf9
priuA8KKum3EVfnDjHA1OZT0sE0+vHaj3G9FgaeArCH4CgDmsh2WUnW67y6cLenK
BRk52S6artJWMeQGASZaBWX+eZTVb4h1v9TQv3S2yGBEP9Ui0lmTb6Z2BDLIKPge
T12djFxi23Ty6Yp9cfcfDE6vtgIP3ji+FqLe/iLBg3YnjJWrhcHFTtcYE5w+gb40
4E7OWnBLP3ED1z3cdrbwRDJ2YPw+65hrU2zo1shSVAme+KIeKWHgOUt2LdYYAjNi
N7SqbimDYQRGXobr956k89XMv7RCvfEHZY/0BSgqSY5bNvbnW7SCfjqUHZOpkL3c
7F2Bw7EQSejErJLJKdfZ1WD4W5KXX5mnoMtMUHsoqQI/jwnX3Jj/MLFJlPlaqPLM
JObFWjm60NpZJC34j4H5t6ds1lMMW3IOAje18F25Gj+Cuv9LlRadrWKbZe6HuCtI
PFdqAnXURG1vMbMco2D3qw8aGqQMeUAg5yh+9OoN5AfdYJum8Wh9bFmwwAEJRgrI
DKP48vNAIR41nd7yJbYiq51TyLpelmi5+kScUTIqaGt2FdGHe5Ke2OuXrHvtwfor
bgz9D6AcjW9o5qtGATbF2wZHMyg54v+DUXLnbfAkSEwvND1hddw3TaWrWUs52uuB
el/UzMYNlrzV8iVS6gSnljYDE5+uELtwjFW3L89AeyhCAce9zyLD2y+q/1QgQ5j7
POSkyADNoRPBNJ82KtWNCuPTdHC0E39fspSd3JiGDdQ84+ZPUJlxYf8ZKecb9b+n
jJUOPbBuDpLByGKNmd5h3y5ZNwUu+PQxQXSVNJj752fszbJiTFzH6OUBRYcSC3Xz
VD4pLT/MRSsBKOp2568BuRTJuJW+3Cmgl7MtIuRgdh/qG3s4FRwFMeAoeoM19HQ/
g9UuE2KQ+DuRDXw0QeqrX6M92VMSq5e2sQWa3WbJ9WJZnnlLEUKI/zsD5YbuyGSN
S3lRanVWzh/OKPigXcbejDNNltkWYFr5torWc11+etlXIuqKxm7SlFy7wEt8iqR7
i7dnNDP9zouwysv8oHMopNoiW9C4v1RXabCmkr2HIGcKg7KEEqQBDVOgp2U+7/Hl
4XpR7ZuMbiIec6cJYyGIfJNceR7CRR1P8TkZ4QJPRWVt1OPGyQ9TvE4vi8WoD3SB
p7W4Q5jCb6/ieTGi3PsM4NALGfadUbDfjTcMdvI17MsqfZL/4vE6iv7XmVIPTluo
uyoy5f+4gWc6fAEkFnzzLuz4hYC12IXjXxYhvuIlxVzrfv14ThhBKhTc5RnNOhJD
BrK8GzkSRT4Q1TPk6MFNkyOys84htFNavxllAm01vfxH515KrlU97RUcZqjeVhP5
oL6ZHU2hgoFhEGRxYTZh6jX+smw3VztuoPVNlgN2LpHq1iagUk54HjL4UH0S2Avd
RcbwCCMf2j9sbBAq4WZPLS4QSbdJn3vNnrucidZH3fqvj/2bITZDYJcLQKPFKNnr
jBXljo+94POCZaAB875MKmlHap6PNwlITwD6mUl4OWNMi2UMRvymvbptcbFbjX7l
H77emzQ0W4MfgNBMM45eMjDbXcIIZ+mcH1Hf2BTeF+YUe1j6pspNnniksd4B+/SR
a7ZikHY5+Z/HFmBQJ0NvKi8LIitwe2q2sCC+3BBF67Kw0azz7QD3D8pcDd7ZgdLd
KNDBZSOkGYYqwESkG++UE64lzeX5ql5ymLmy5YVAfzlTrpXgLpDbYLO2ZdM6q/l+
yw6GhyTWlg35PEUAgHd+vAKkCGU7HQ9vrsjtpDM8RP1dsXEH3B2td5E2f8h2O8ZK
uqp6yw4WQGY4B2p2E8nGt6qw1XfKghWQvNa7YFR8jF7FLQbBahD8CCTLXm040Prq
phG/RnxG7LLOLx5iBujjAd1zhuLNnJfxGomuzcvgGLRUhbsOqLNxRF4CUIA+p312
Qoql21ouuC6qTe0+5yr893G3HPPxs+8PETrXSB0cpoANgKhU9GZ1N2BmksmSFyJn
PrJKdNwUiYRQB8Wz3qDh+xnx2DBxCpHhBdxyF9Pvds6em/yqEOHB9Gpi9OZsqOKD
0f0fu5v0rlCdrXT3+5wwA8VrGecuZxE+XU21h8W3X7+m+5Ci1pNRmOc2O4l/w7Eq
9jGWc3fH4JdEXMe9kPrTbYQYuvZbnfQy9AP/CfwM1WflfHaGrY73zCymcWJUHBW5
5igkfeyK+VC7aLi45LwcYoJwKq/RFET/9TuEYyMlT9DxWD4sxnnA3rU2E+hw96hj
oIIfdngUU8wp9OHeLEMKnmyNJMLNREqEF83HnIik9d2qdBhuO3Md71P5PI1AwuGA
PRgyegBtUjdBA3JSWPaOAh/LkQdtlnZhWVNBwTPdoWH7mlP0miGNfS56sb/p/XW9
R/cD9pvtC8irbv2HSalQJ6oVvTxTGOnDkv9JzVTOTtyxVFGdFi5+f1/SD9LKAZBD
0EohuxtU+S7/TABRCyihXkvCEnY/WYbmuc2G7fpKhDky7dGU7dx0GX1YW4b7wN+T
W4DjkYwL9T3GhsL/ik0yYAeA5Ill+p4W4liXOgHMujTBJGj6b/uQS0jLQ+dupduO
2lIFs0OUD6uDDkW4DNFmo6lv6EfJi9nU6aO+LBF1gsk7MAvFlHXoe3OCbJ4oxaFk
1ejshpCSkcamH90Uj6UHMEQnGcxHMV2omNFlSPFmNfGXPrf9nbNMXh6Rt4zhRgaJ
3zdOn69w4GjsSXjbdVypq+dc/BU01sn+e6cMZbumNI9FQh0gSyyjfCAP4E8bIjHr
+DcaibL8Ym8yD5wUfTxyJePCxm4s8uuuILnWM7WKHK7soToCVvxmJbBUp/NQf6hl
6S6YynnOKRIQTd8H6WQSv+mX4YQoI9AeIZSMFdo9uxC0oNXlqkFR61Cl3ZJhb7vx
1GmwXyBXaojNVCQ+8DKTRNDg1ebiB3DNvwgTL8OKhFmX8dEqPujOBSWFe+ujTshK
uUcGT7KDkzV2R77gkZBu6/oRYF7wf3mcZNEkjgHO+RTcNcMLEWp3tvXqu6JOeS7n
7MVPBd8q8D4DYfiH782GD2rFJIfrM1Z3yWecVszwzb6RZHcCrB3mi4I/mMDVNSjU
QAoAP67oNnq4XdS6T+psbMnLxhCcerIgsqr4uRqFiwQ9fjPR9WFPwMiLJiNgvpVj
5UrE5XGY/79wSwMtS3VNZ15SyBtBBjWx2O2XYk2E2q0xuU7ERTlceaKinqY8q3UW
Kl4WQ6jlLWxdlpseU9FDPI9C061JJQKGDQ2mK7B+SwgFVC3KrsYEV+Tkrj3Uva/u
jR1SKI1U/D0HX7LY+G+0sVUxWFtkWqArFS9biRBPhAV1R9aWPmmtq0a02lQYs+wP
DjIxEW3bqEjb+0KV9+lK5HHza0OyYDuA3zKi8Z5gOBsVvrLbI+O39DtSBsnclh8c
Vzk5lilQEkZ8rjBGGezYbouImjczaZ/xwNHjNGhPM2fDKTfceSi2PrZ1RCACVHtK
7XczOHBdLQSXuDAGFdsch1WcoKuQL2reaoi4rh0Yn1gJXKZKjd8xXxxdpzsD1wY6
w1F3/WjHhuycUXqFAkfhVISEp+0C3z9Y8/wDK++nmPeD7tSstvHIPPzqItXzfHck
cyiL4Say/gvLAsRQZT6i9VIqMcbqRTCQ3FNs91tR8EVUDvFgkZSeEXbCk2lkmjmA
lAUiraDXB4WPf4/V11cM+I4vMwq7Yds+MXUITah+tDJYc+xTBnbuOkXzL3Qm6isv
yQ+NNgUrT3OqageAQM7AZ0u+5vvauIDuc63+/rWkKue58+dcKQP8AXx6+ROfE4Dq
5vw1Z5eUQI3GIspHihFkwBCUteVVYUJD+9IjmkognxrH41VBTlciBDXwbuOH47YJ
4R38OkEo5swIRHW0+TwyiU0mYo5wjcIOh7R9tC/jT4EX71A071SibQ6M0LQFRjYT
ByXS58wQ9bqwPPX614bPN11j3uc0JfvxkbCc2O5aeK6dWFb/nK9KuTBxuBUWWOXH
xLsilXcdPbArEoNF0uccHOTQUhKbLR0hleAEz2/3rwgDIm3wgcw2ykrhKbYQ1+T4
Jq/s2Yc9/ryzox16IDtlr6NP1x3nI3igMo0i82I5JW8AN6fXmGTfE67nS+btd64j
W8PNOildnqFKgraDDTwA4A0H7vPWL9/DeUr73I31S+bo9ZyJBOGEVrwrIIz0riNa
Clt9bI7VKF38cDQfS2NDNDpYEccgdhrhzO3XiqvgM1BYk09o3011UycfZWqTZH5h
hhin3Vf6AKh/06HMl+NW4K27WfvB6l4HIIUH+XI6l7OQ3L6lWeLhVyqF+r+yk6SP
/Cv/xxByRmcgd5e40MNGOGBBjrBQjyHQmMZwwqhToBopIkxK5wuC85Flj+YP+q2r
3mJf8qnmdI1fRQT4u+58jPF8bih7AyW30Itnd7Y+CqBOlAO+RdJmwPxW36Hw7UUH
Uy01P7c3DapmAxcQcFxkdpxl15RJ0cK6TqmtwOHzkeMbhZ1Y4QsSLj96USTYmmEI
sRi8v9ZPnW1dOvGvIz+6IBTBqtVoTnJ89o5bNXa5Z931h+lSpnJo/5FfsRa538YD
tmKbMWvG2vtPkwEpAGAmn3kjrESWeJe5SpiCEu9Mfv0TdH/3AWLV/LkHn58W6G/I
Bk4ZBYLBsvFitFrmJB1ir6ZhkYAwab2CuVWTszewz5YGcxvHHJqmWLQFyE2gbImu
rKJAgtpsYB9tQlRuPS3vyL+08i/9gAx/7BhqHx8yCTSW3O5Mqw+X1nCsC8QzIEFC
cDMPmequH9/KzUu6NHvtnJ5/Su6eSykW9YtUiowdaSAZRFJK49+NMvw28jHEhHdv
9pHARzOLkwB4JR2VeJshY/ghBhywRotVVZ5ESqIonE0vCtYafPkovRefRI6mY9ul
JBgQfMav2R5Ah9pvGLAaASGMrgupP5Ul53nwMjxQBMaU3BQKVK+yEVk1T304ZSX7
GoiGqeEmrA8jS6rSdG1SPj7z1uonasrdVKm4llynC5UweGoTeVlc9aTvg2d6nkx5
+kee7dXyCUEGbveD0Yxn6k9OPIi2DLyTybz4M63r3qEI8Ph+nD8AYNo1nXEjHwUn
sos++Ozcno45EwW6ozIIzCiVBywimVEVpD47Yf3/LK14HotpbOTUBO1+RIK/8w85
s6cjx0TWcfhN/jBFSYa3yf66fWxk1BBElmke2D8nkmoEDpD6nvwcAlnDb4jm/dBE
5w9S7/VigN7/Z0zCkBaS0aukoHj6M/es+R54zfrejFvGWJ6j8YoI1nD/u9TTpvzK
7erpN9W7xYSLrtt86hxt00fIaNVFxX5UL3ifXbrwrkvf4v+ozaoinhA7pEuI/VbU
0UKNolHDS/QJYzNEh9D2X4BXV0iwlSA//TN4ZLnvSKQxRYRaguuO+7i3oy8PL+6v
yxcAiFP1fOCDYcj5xUPJgMuS2J1qMzi/WggNJ96D+SkDhCO6vDOfN/o4gazmjBmJ
bkTYGgXCnYBMBoerjzgv3PZLAg2Jjx5HNaxFYpa/KKMwIPDicPVbnuqUJxISj4u1
1rys4IyXVG9Lj0rA9icTMRJLYyZ1u0hRikOPlc7Ba3J+3ocDdjtkQfjWTaPu4jOA
xCLfUzbXpNqxc/Cm9acopovRoUc8z9jgu4aBtLWeXNCQlBaadrT5hJz754kfnnlE
DRlKaAltTKD6Ef/Rkx5BLYyK9dW+oM1pilty5qdfOeWybvcX6ss+RD1c8B8fjy6o
xUN/v3KTwHfo+TpnEOMGQ/PDR6AzDS5H0ucsIHti8TKehI+ZtRXu6eM26CMoyKB4
WAdmMAb9GMvyoiN3zgCHRhEYBxS9NpnSB3EBP2opJhpmm94TsjOfI0bHp2UNhGgu
DfOd3CTC2TEN0zqcDAUEGU4bHtl4uUtwZnhwja1bhYuXTT2LOOa/BPmZno30jlUA
+YOFNLWpyVDS2+yYiMxsMcQJ5IlwWeSTG/sDGCRA80Wc58v1rupMoeIjmMMQeQNR
/UQBet4njcSrlHx1ux9Zx2pbnOASz+Pwvbk6mLK+gnKDiODyj0JyMyRtCWQXpZe3
HlfRRa4u5oqwstB4dH3mRKNZY2iidg4RsoJjxhUX5/mqPSf2xr5vdcV32WslcueL
56dzMI2IARZT9W2izsgQ/dacofR3MTaafIGe3sZ5piCeVkqdyRXUjlgJDUrnrs9H
keJlbR01n4hogdIZdmV9BCp3PEUBKtYWp/DkBFD+zw358aJuVN269Djd6h1tusmf
i978k2cxAGYYOnBtiHfy9Wl6sR0xBaPTKMmQl5itVoj1BccfZhZeTXnHWlxTeb0h
NKoOvM0jpA9rOScr5b9qwbi4zAKwuavPcPHRX02aw0GRhaXWTQSvBYTfQArptmQ/
wubpI5wVMUqU8cX8rix9Lbcm/sSCxO1RKV9MALTK4cBfOUKO92CSmY5haPEOIpvz
o5+G3iBwraUbH2BS8b/68gK94cVTXc3ruDyDG0Sab2RDi4HAT5ITXodUiKBlwF5W
5jpNxwb2p06SuEQv8/Uuf6C/liADpD2s1xlluCxCTVK3P8Sbeb0IqUp3DibsKIGs
MAfqXUSp6K03/a9keOO2oJ1SMIdPLR+xn4aeiVnQcvGYouzCVCgFDaPmjj3wtGI8
SUelxVpy3DJd/YpOk78XcGPUq/6MYhiorf0ntKhVLKwW/WnPSJySlm3QA8AcoqPA
cjmA4ivYy0/yDbVluNEl18skRZHf81tHTQqTiKecpqoQQyA9jTRKKkBSIE4wxa/r
dSHJrmoDtucB/8lbRy7kCLHbFmPiX4uYnJEpeUULspQKj+I4/PckSUofeosvyjJA
3EduupQqAkGwdNarrSs08EP7Qy8X68XzUTSfB2GGFWsTNEDxOaQBVsYY/1v7k4xP
KnI4pXoQf/akiv4C+ckOS0vgWRFAdD9ytz2lhpisnFzCngCIsOhsPPukMR7YySVY
Xk4cRyrhSD5ou82R4IRZZiv/CIoWFloIslUlVAS83gn/+9G8kXk1TBB06nm7cJeq
O9VHOLILQXY8DbSxW6S6CHDgnio6J8JROJU/gSqxNGcc6PubftDRZGp0dDPHM1tH
dMK5NJSWdC3hmrNtORm7Z1QD9+HLFKfzS35d/GoNGu1WxeEAxLsuTYqmh1bBXwU7
cy0YJArAg1ptOAKgMfAu8VBYtNCXbLN+Hq+fjC55n+WBbKBnUZmUWlKiEEb1fh5T
p1Svwfbc/2tMFn+55hv2J1vGHPDCoIrU+A5UY1xQcja/UogjJQMRA7pBSbKgrdsL
vs7h6QSMFeMfnovUgS27FRdGVBntvWUpFlMM9vyYpjzlz/BrBXtLz1SmWySL+pzf
X/HkvVXy4TQSnJPWVTNB1QXmLrAefLSjAMKSa3PQ52tXSXOzCAqvwn0s8JcHpdsa
XDQQ2NIst9Hl1A77oti5tDt3Tw+yTjUIUTx+CsxCid+blvdekzxH4ylOj07q9Ymw
qGZ4lvYim0Oqe/Rx9txxVCYYZYYZA54f+7alB5wSI44Vb1o1Me+/sXnLvDffQlzw
L2BRCJPiA2kus2dzsKjGfrRMbyAtKD1e42FZqq5ljcoAKohB1wkZMhQZ3rLpNQo6
ouLLG03dt0/Hdq0sEZR8ehmzuiK7Hdnn0iqSpPiSLK9df63vCw4XToUMR29BEamR
Ovq0xdr+QJntdY4t1Cu3bJEVRabGMtxTNmATtVmUE7a8OjfMRbQrGQZYlOzGAozB
crUVszz1nLQnrEj6aoa4fOMrsDksyNN3JbeSIR4/mJ4W9kJBmwchYKzGRPNCk9IH
AGyVIdTTql3IUqP+UJFpYX0NECC00EgrHB9ebHOkosO2u3Zcs+6+64noj/iYsKRD
pUvqrDHRrobSZv/7K+Y2cn7sj4g2U4YdPueGzD/tcNRpGQX7BltbKwgbK+D6WJCu
szmbERwzFLwOezaEDifRkRYBYOz3MIy4oW8yCbv1fmfjkwMoc1znW/nJRO0nR661
uC25QtbCp/t+U7qPbygyvgifF7dNY8Pa2MVA3FD9Pn/127JVfqwaX6zJevKflDwv
lHjiNK1OgdIA3gHeUYWtxb9J0hc7s9QyVHWGT3Q2U5NTLWlKzJdLxKlkm81rgK97
0J3O1R9+V1zSnPyt2lQ/9WiYE9p2YoC1uac8GRvNXhePNprS450f+kLlLwZ2L1Fb
LUnDmKdvUxF3DsKl34Se+XwEWQ8+Pi9Ym+2d3xp60yACOFWECwCfaQCE+Nq8H9+a
Tpk16OjLxEzq+JZJGnNeQ3/rfm07wr2srYffrXI5ctWL1cdQE1gmgalK1asePLhP
oH8qd6b9uF1VuYahJkYuPfH/+30CmEDbICnRGtj6gkVFk/EU+6o49vQSsj3Z9ocn
A7LT8/3Kxrv6oJeLD4qcneAdmjpAdQte+c8PnYLTUq08JPVp0UYWKVYlajs7uDH6
vyYjZAyQHCqvXnS23Lek2cOXlnPOlitgfliftyTDEynLGBsX0qnXUVdE9hyHowsk
OacE/d7xJwiQ7tuF8PgYs8k0WqDYfJyLf580oxYxZ4TqmnoqtYMmtuebIYaLozyi
u+v2L+5aNjB/QDEkCbvIEU4KgnYk7r+T1cubYqiWky5kD2fV06D1FpTyxrbSXUmG
IL8/M/zwuOlQU7+ZF3oKO9QZzMbdBytEraBKoioVxscP1svbLlAe/T0+7OswsLJJ
VChxlF/iiDo7bTjs4Sssw/kdjz71wFoAvWRaORGjD5600QMxd2gr79i5ZdJghN2c
ZS/oJ5J6HtikskN+aH16FRD8e1pp1l4MOt3y2VDi8E5URYq8QCQYKgaQariECCBM
HMy7HWIqaKriFAMg/92RuknIX+OLy2FYLQJxDEyF4T1Nb49dvSj6zuThM/Qs/8x0
pXkO6O9SnbRC3Q7+FPjGuOiQ90uzp19ob23kqiA3x3hIcKjWI+6vEocqIk4AwgQC
9NQYstEEhzv2ijBj0AqmJZMhq7COB0WJUThPLWxMJVUVxlXsljJzF5m2szasz/ZV
JJY6oJdU/MCG43nBhXMAxiWo493RIX4bNENEfd7UAQmy7zGrbudDMheMzVTmd/Rr
JX8G7c3vqA769sqb7WVqp5wfJnHb+OJek2a2VCq8sOgtVlBQXcwnRdCwvVoJ+csG
ESls/27PA0FH2Gs55aGZPIE4WauH5LY+sm1b8B8We6BBsfA5yO244G2/EIDKv01p
dYMBiMvcrzGxQp10Fh0sDEsFSooQ/pTmDbzZdxnrgNYx71G+WS3yGhNJVGyRK9H8
IuWZ8ACtge7dVnOPQrhqv+d4gFWUlzhdc5YMgUYI0megAqPn+kn9gu27Z5fMQR/b
iHVjjFaL0cb3wE+4d4Kx9q+db3mVgsboGrOVlExsaGNR9NLHyMngpFkh15dJA6hx
fngQ8fII2ymQ7bxd/ogXT21gYcU1LIa0/tSjhS5Fliv78seduWTcEQBJIxFJY+Kr
FIDhaX5Xz5nfbxc2hQlt6Ab7Gg1B+k9S/VmEzMiqxtPSPQDK3EOFOrja9uZSUQeP
KmewrnKsQl1G2/Nh0uUNUybpe/2xTzCZ81wYxN2HbtfdcG55e3/x4wIWiA2/Zr5M
97DHq5WcRZqmNBRDELxFWlwVdx7CqOvVx7vQuemBNyZrtUn4GReeSA0EJrll9HQY
+lrUd9bza/vvEM8x5uehuHcrkM/orrms+08ACGDPhAhHFTjiH0cNUOMRgA3Dyd1g
nDuLOkPWjG0WcWqNzNurr+xwkPN09mZUkf2cf1PVhrz4dTi89idlRxfovW+PFch+
x5OiyT9NDxmjsF5j4LHt1nbwMCFnFOayE5kFPFvXzbAFQOnmk0lRuxu+GKe+FRYB
cl3z6fWDItzHxcmJ0WEuVsgkN9vhn5y6bgTCkHYeKoYld6vSowPIPIxHk1r3FQrl
DW3OJ6V7fERc8Em8oyrdZhSOmDW4wYbidSu3EU2UP0hh2GguloKiYhsOs91H2q0w
0IeGP1Fz8E7+nlJlh6h/y4bWBR9+t28rq3jw9czps4lyAbEbLr07atc+V1AGZ6CW
UvgNdSxELq4wEvW6AGd6zcZuOHabDwehMz/Qle8vLT3bz4XUlAqB2ZJCH/Vl6gmC
QI4fiABnWDwmHNp2CQiQ2GOEz3wHQdyrgQIf/dOOq4+OHqhxycWpmJnXmwGuPXi8
ccgu+JN8plM8KUuAb9sKAeCZeBVXDBJOX8G0GYkgrhCCTN+/aVoEQqTZPZTeHvSi
fopHIPCPrMpGvuJmC/k13WgptW4o5mT5SvOfwpwvm69QP5LxuvvcAdURRkT7u5O1
tM5i83Bo4gnhV1oCVUolSUH9bLu1Zt6OuiufyCbemmq81zD39NO8PTuZ8f4E+Rdo
VKci9f3j5juBRl92/HWE8etCQ2qT+NIcUsBycYumCbLQ+cuuAtG0f9pwnQvH4sjd
+JTxwW0XTG4nEGrJKTjKl44s9l2dqtqptwb9qpNvMHw3IpSMX4V25aNiCVWR3Cob
2IvuNanl1uIGLDOzD1EcUYpzXtXCe8lDmSTS+GDrSm5PzVwdQkKlbxWGO8vLG1+H
5vvefJFWdNMMVd2udClyYPM9fgQdlFVXTcjCc3InOWm8gGDfJLjorvYm64Tqodof
D4c1FRHy2XXsQOjeXAPXnTVdzfjNz0xE7sANwOWpdnXRgX0erfEEE0xh5YWnhGMI
PuDD6snhogC9yKc9lpvBBGy2rC3uYw+hvnYAuNeEqa/zyDiKJRAYfb+P0oR+OynY
HFiGQ/gwjGCJkupdlDZNVKFLrPXXQFQb8NC61Wii82UC5MlST/0aWs+44Ob2qkzO
w9r/5YiLrVGf/PFTLPI1V2Foai5+OgYI6yJB8rF/DXZPS/ABvuIoWdrudOfMKOE+
GexrxHKvz2tRZPGKZGZOOjq2jqeVumLimujaq+iQ59mShnTl8rm77sCax+DrVx8m
QCnK5F8oMEG6p9YiMeuHkZXk6iieLwpMlESu29Jk6ugkozeket/f0CKb2fqmR22h
Ygi4RHDEx2pfNVK/IUQYXvOaAfu8qT1bwubdsTBgtEK9+wEwyCr3d8e55urOjTzP
9XkGLqb9/CojYsklxXZUbwIFW0gsfyL+I4nhbdUCTBHWIZ1Q1+SNcIHxk47Qo+Sj
apY2u08NcZyjLFBiUleCQjIsJBOurSN9t9I1iSmTjyjO/67Ll/miHVrnWvQrIFK0
iS+rTSSw3L+oxBZE8UPzlz/ybCmy4TNdeEraB3BGJmD7pEph8MXWN6BaNRkUKhVe
YFeucEvC7Q5WKYyMCydpj/VseL//my6DWQQjXAtXzLomhrAapVgWZcV6slmn6ggi
p53J+P3ro6Q7qSwa+nxieQJ0LLheXMGtEzMYl3B0byUWg1JkUlXQzKP82uD/hkLB
oR3lUCLL4xlkX6c+DbK+klzgx8Y706NxvD5+5ZbiwUrvJUoJTBD1UeHsCOpIcQxu
zVhqUMIs/bjVv2rPqKoNNad02bFnnOUgp8pw2Et/jOCIRlbnPZIqsDmO5qeS4Kkc
cziciiKKsYAcc3VTLDZkcosdJrS6WTZXyBpwqMn4HQONqT3sGPM7fH1SNr0j3FSB
bouCCjd0azEr9oKe0J7/3bgOD+z85NrFLMjafEP8kW5hH99E4zDFbd+0WYPvvk0S
Zo1FYiDbqKjcXtdP92bP879Jc/hHHgyxLGsa4wGhZMY9/oCT0kebMFh25d2pepC7
cyWJxL6Gb2UIFran4W8tfrd6OvLE/5jtBezJKJKbDlCLSheFgu4w8Rl7SwNCJdzy
KEJjbwfFzcCVkfQx6mgtQvWhqyezc2ng+OSHAlbO5N6YDyQskSJYkzdhV8+c8hD3
PPsR6ZfxLSLqdHqg1TVEr3mVkmptixYTvR+7baMNXjbD2fSIM/l9yoqOBKDE9tY4
57NBF8CqoSwzq89MTpG1TCTSh2I4sLK3HQcTiJKEeDxh46R8Ckr/mjvrkZ5aq5aZ
eqAbnrETVqAANzv8A4pOQMHGMkRn5CYEp5Slc7HdC0HVnZ8kv0fC1vuUuQS2LsgT
msMFGMCvhHM4kXklrRxh0SC5kkg4bznrjyzdIIwRb4YaIePUyCGeMJEW6Eftpi90
2yAmmCR2955gOq14YnumFs3X5lWOs6kPwNG7RrmH+pdN2RxWanjg9JcEv2iVwBHS
1698DKoY/oH84dNr9yMKnSYxlFAooKfyc9X/3LnEk210df5Bc7TUCSEkDNmRdBB0
KI0dxHiUQlEiSlmS9SqLY+06uImIeGGnLfWoIXvzccjWXv1CUuyJLaKD/Q4V25kR
hm0++VOMfQ+r6MN5O7/lWTKiRLc1DqbBwPU/nJGTwf6OJoiaTX+WMl3WUqJ2gKRr
YKhM9QgFpl/I7bzU1IuSdTV8QwySjrwI/AOgjcjwhWb4lNtJ/mciUNRGWiLueKUk
NERwQlqLciYR8b3obv0AkTIcJdq+ZgFgIzXWqTGiQ/IRj8wPdE5N6LJjUc8DPuoz
DUGsZm0Eaxxl70IUSyyEsLfXxcqKR9aqVFBag96dJphwzedfplWMaDcR/oo9l7+e
zkoj6ZevQCb8L/oSuTrrjK4lgPwsc9SpgjL3yil1SN+gJQqftMmNohXaINASLUCk
ZnbRVfrZ8AqGIrvGGxa9DMES/Hs/sugscMV7O+nAMsg9hD686gKy2NIa+C3x3jcI
Tc0LzY/48NqpJduEe8lMgAjP8hlubKCAakEs7DfE4lfl177uR+2CP74+YiL6hLF2
KODG3Nm5b7Z7sb9fMZIP74Kns/+YlKJ0RCS4TIUDMnxhxiWpJORnYplLvEQ6mpSJ
FYr2u1KUwSrH9nELgcP7CTirOpRVgYKsOjPtS3YhM8Jpq1E9aCr1wDKRJt/lZSw0
zLiY9uuX8ccGtE5mQQjp9jBhzl6W/h8k92wCxGUlvJLTMnd1HQMPUrOYoXRoXQri
R+ljP+8YIX/HPYH1RxyvNdswSye7Wz/qg1gb4KDbIKzgw3ktzzMzVnbpjAOI2RIP
y813VCQk7oNet8JGBRbUDP/f3FV0xOeXaBRdyTsSY/pQPxuKTZLM6TVrcA5L3e+I
Hy9u8XkyhABF2twqhNFU0nXR9m+y39fIlByXBC6Eq7VjWkw0oP6yd3eDvGtMQ64i
uvfIsypb7KuGgcp34SRu+FVGTMp0mSn0OySMFKRGNKJVmzSiMUGGI7VgFugdrnXb
cu59RqT57IAWKnFyzGlUo+qCvJFcPCtd6zM+3svcyxFLR+B2pQArHNjU90fuuLIs
xLSM5Itudzh8F87ipyjdnb2QLH316JBRcRUxcEZrvWtMcuSbb3xU70IGMlQ5d+pA
px6wF8+eVF8CIyNiQkspY94WnCuMLW+wyeziky6eMw8QEi9Jsd4AzfHNkILnhqYC
1rhKgoZkkKazuHxi3Gw4QeiySR36P1ia8kJOXBdQgxh5fUGFG5SL30GV004cIhuC
xDPkMIzBxUZ+P4I2ZEWt/9xqpb9fgZsIV87uf81tlArae4pMrxXxFpwHrErMF0+X
B1m3dxQNcaKPBqTNDy5nBVsbIMAyPRRRB1G2818KQc3I7oOSP28PvIx9Wg9ofF29
3H51+YBDP1Tj3JITgN1nZ4YLxt4NZBlXdvzSOkMKg7hu0/9LF2zxkTqkdnXb7920
IUDl1hI5/8D1hrGnYJHv6eh5mCBgWz1v88BK2NzM4rRlTsOpFCYGz71ah6yO2sLi
YdSGYiUmxGjQuz9xvFqZhdmFmiKiNX4FZwmQShrEDCM3C6SbG8HRy7LF8x3z9k5a
0osdQzpbncsk0rlAM5Vr0p9YcwwQR/Dd5LDbeMODXTehU0Hu3KpJvvmUvJl/vFD5
hX/oX3/YBnnZii+J1UuCiy4aRktTfEZovkMI1jJBoJTBOYeWzu9dzFY1r8jNXZXd
1sbuw6Dbv5Gl147tEYRh+SwnDxUTE2zhrrPMsIALSoQ6BlEM6qxQjukIeGZZzAYF
mvDROOi9a0mawfWJKAQlLptG2v8vH/v5nkTwiSH6XLS8BNkcJE0IMkYkMbPwCAQM
cLnUQdTtbAN+ODKqkSjPH0jbbJmn7PMUeH7otAS8heFG9AmfD3GZg3KynQyAR1dx
jWtVnDXisxAm2/k+XSClzW8oV87JCP7H3u+MK7g5R/8Ln42WzRMVAS6rIVRFEcpM
XRB0+AObQspBT1nDS5MIS28qvresRFJ7xkndoAuvL43KT+yqFKr2ocvi6/my9Zsg
Xboi0qmAYPXUf5znGqU8fvLNSUnqM+ZoXuAbi9xNFCZx5KWnbbErlA0AuqOzg1D/
2UuaKDP6hP7b6g+l8hEYhNGdTqvaRAJONi9ceQI+kBkMcuirRiIhUYl+WaOtKk42
H5irxUUA962CIwZuc31Agb5eqqT2m1+5N/80iyyuS1ILGvxGl0TFtgxFfqrsrZoB
8AHyiGz+rXqPel3qxohUe7VwA7PYVMtKmzqn7w19T8SkUuvLU4aSkWqpdZ3vTx17
uTZtSEL0rID31fYnKsIMjJbECuZO2bMaQ4zzyV7d1sU9lcIIOoBmaoB6F8mrqylc
iic6CgjF90cxCAqifF4gGwDJsfBEU9AvrLfx0H7gKNlRis51Z8drtx3hCy965oPB
jPkghq83inOkJjgNJWPzROwLLRNBT8sRYi/E4VqIGQAyGIPEmM5YZ0YOculSzJnE
3IGspzYlVzw7oIs18+wkpCv/tcZxGiG3NJFRSQ6+bcUPrB/KxEvDxSoMdNEfSOzS
WBbrksUK6jGLtxRlpwH4XhOYw5q5xdLh/QnSAqHFl9yBsSUv3TXWLLzq7qX7FWMp
kxX5ylSWsyKQ+xB4fMlyeIHNC5I4ZcCIfucTRUEyH92+XMwggCS2/KllZi8q8YmH
tGfkvqwdcDBCwD4Pf7ZjH584+NW3qQ2Z2GOIAGJgjaCDJS3O2Eb7/qp1LJ+RbtUb
2I++yxMLPtnMVWvdNeQva82v1W/pWeEdSFgaSVTfo5Q9VY2vwm+l/R3KYKsQB6bQ
n6KBgIq/59wHzTvhPkiyf8ogPnBJpJjiL7LTfKX2r0cEWhUMucFJSEFU9k0iCYY2
RW13LEM0kYrriZkdQQK0EZ8MvXx4QJXsX0XzDIvK3PNrbzJfn9tpxAm83X0M20Kw
Z+EfnSGwiWy+b5+cxfubjDj9CdaCNQAMKuOsvccb9FN805yHshLcVcv9Qi5skb9U
k+u44vLoA2fLc7bSuLRp+c8Q11pZCvg5pkZJPqgLa4pWmx271RskhdQAsxQ0OEzq
EAkqASCakcV0FI7KAUsilJPIbV8e0OpgQAojwOEBf2saLrAyhSMVS8+aWud/pD4M
WLGfL4QUCGCp5N5zrX/oUBYQS82sY4RKOeezx2BPvlKG+UssOYBHuMDQ7r5lq4Bi
PmhH1+IvfeUT0oFI7+ynvd8tOjnlKJjf/GzmoTm+AKs2s3kNP3TyJBkeulCn/Sz6
/2BC2Qx0WEJapI2PaG6XfQgDKaHDkrJOCnTZlE3/oHlcGmBtxrZJZjHkOu2nCFzY
EaQRsKLGt2fL/MkV6dOUpV8wGM4ArRdwGRjzrZ9NG8HVuEvO41/aBFZ5l6WVcAHS
6C3B8yDoUQidECe2WmNrmX9V2lBcPkdFMBp/l27+Efafedsar6R4as2kRNYTyt5O
mqVfBo0d8B/JsAIy3GQRYO85LCof2/j8Y/cF/XdoXkDch2iN+TTkC+mauhogwIJK
K8pJUXtJ6eTbDZgVjjILwdFZ13Nnf5+2W6S09LLzyi7+w9EB4sLeUI/NvVhTC+Kf
8ugsu1afIY1GVd6gg1rUZRS89aiHaFYnyLTpQM+zbiPA40HCeNQ+D/Ww5eQBj2uN
pP8NMVHmw1Xnlij/tmk2CmrQMgB/mNrfmgdB/ZCiVD/2ntVPdzXH9V8N+V1ka7US
ue0iCM7RdrQsnitAkSoMQbXadT14m4F76KF+omWSzH26kkB1XDO2zURKVuFzy3co
49YIPOr1U8V29NPUrNc/BWYKY7BCFex0/xU7fENxroLeWzVdanzcpLwCAGSDz2c1
2H2t/4lNEBFbNtDgdsPOGqk63zdWGML+5UvDiTVu2fFgxGT8tDzYRgrUmDVOAzLj
+8IdNrA0JVm0xZ+ZkmLRa69+FiR8CH9Yqo0EHKW6lkrLMGjT9FBQPGN28j95UgjH
drL/0EUwyTmtIYVMzkw84S6HUoep4atHpTkWdnCf98grtA60CVh1r6RhaRot3iy6
lx2Lp/kCSnMwpNp9C/S+gTB4KSDPNmkKxarwedwwCa+rYAkz+/6ABVPIw/oDaBUc
bTNpWIfIMYqKG6YFkIVvYYwQTpSPzYXSiW8CJO3dB9RTYdskNAqk9lJEwuUUA7GP
g7HPT6S8g3Ehu0WJvn1+yFkrEeuh2WT7yb/15WV/SDm0S2Jz/gPJgumySaghN85v
3QbzG14WvYktdoO5+dVqAl+4t4gF7r881GL+hhfP2NgOqbLkcgZU+SMPaKsxiQGO
BaLha90z0kWIsGkLM3223DIxjboxA12kqyrz1uJpADiThHUrMcrrJYzfnolb0Htl
Crpwk2zPUbneqsog7SnW3mvXt2s67HINP2w/p5MObVb9pdrnHHZxG+zeiqDt1Z0+
dQ0zMRm9O+HrQOv2GyFW00ht+MIPq1N8l4Yqozyi1ER8Wp1LbvY60y/fcYbNKTKa
ou7a6OCKyb2Eazljzr+iRDrZqxb/4rh7u/Pvhb95guGfRNM49CgI1CaBLlUkDHfY
r/QP415kWk5e29ppdQLVgB4L69XRIwGtt77QjhJrJvE4Nk2LH7AA/Q1Zczhe655T
fhASoy9XKgdfK22gDIbUcpTQBf8q+2ZEQmSH3VPl6qE6LS68sYCSB8FMtoV1jWZV
3/xsWVuM73EVYegqiCaltvH+xosZ/YS/zzDURjiRT4SDZKs3C8h+QSU94u7M6DAO
7P16phGTK1BKCM3YpKO14Alwzh/Dq5Cn26GFzL/lOHvLqFqA4n/2hCUW8P+B8LdV
RmrCkc88XUHy1lJsJ3mtC9KjtAaAU0WkymacyP7QY/EwAOBn88asKSQbHsEq+Bl2
6cjiGyFOIWlrYIkDvJrEG7Hf8PHzJEwBFqDeWX/FKEAmwkgFWHcAMeEOMlU2U8Pz
VsK/N8N7U25zvSq0866BL6b6LTLLJmkLu0RM7aiRp/z0AobO2BCp6FkI4eN2a9A+
7PO0doH8asSpvrydpCbmp2LlNzRQns7b0xv7RIGjrVmasFKhRvNRlNO7g5G3ZNPn
EJVUSXs3FPB3Oi3PryC/qdssFhSs5dS9LEbUCuuUGTtTlmassWsseA1msEIG7UVI
lnLKLtAOPgqCrNb8FqgZuXr9Sd0n2EIqcqVcJAb7UzdISS3jQ3GZ7kyj9cL+yCA1
sUA9IpMMC4LF82Z56JMiBd6uI2AnMK34lt4gYPgDkuOZb87PWqtlG6Hgk+IASyhu
Z4Mg7gO/4FJUyrJD+ddITfOJvbRLabnRGn/9UTZP1bT/Rfv6UxsJlY8jN/gonqZD
XGR4XCdTM2v0+Tx60uQsHHMachUknYoA/yug9vBVyfLXUYJGfthExhhCUsLIZwJC
Jo1j0TZAP2W0bZhBwNTYHEkSCmyvFzXnPVS4Brd4es/pQUWhkaZpHqHHDKpXDSsE
tCbOmeMh8jbsZTZJPTcuj86hfMsE05mI5bVvVtkW636+aERxHcj+wiBfxI7SZgKw
o4yjMXpXGX+AEMaqxdjQM6kFfBXdTQWrXW39biZqtgEqr+oNQjXkGZVunnmaDMSk
4wvmUsE6Yzvsb6sLHmtxRVNhqBvNI2B71fSt4i3lTD4ep2W7Su9ezPq92YrxOAio
oqBvrHTpYKJ+ZXtl3sMfvSAzeq9PFWicBv8WDd/tOb5YDxu7Rxr4V2lwvXYUIrkc
goYreos2vEUVN9KsUz3rHSCEPawFZAedzthZcFISSMy64vaVzKKzVtppI+lqgT04
pdfIkeEJrdHHIcorN60twXKZkq4PbDQVD7l12GBGyGCBG4y1toL/g76UNEi37us5
8cBXo4gSEP8PuwHxQ7r9CFFJ+eJVuIw+kMHlsZex3JCaMqer1kbG+kfIbElWk9zd
v0K93NC3o4Ui0wLlUeJ2vJHAPKDP/WdCpgSTDCamTKD5fiJl1yiSbOBqtSgP6o4+
z4Is+V6o8K7K6Giz709/6WFD6TBTfAD7CFZ8rfGR5uq9uB6ixQL0he4+GGuXiAvp
JzbORbPuZSeai/Uo5NqIVd5CHBComgaiKrC/NvZ7FpjEI47TNgS3+Cix1dHLdQOe
MHnzefsF8M3xMQTUbseDYIECxD38EfzJW9uP343Wdy3jm+DJffyqhTOAP/JDxfCX
pKEswjqjUEWCBZmI2Wlj3+9MAn89kBuAatHED2lir8APEvFlJ/8zleIAbHRRjI9V
BPss/YHJtsPjNqD2CR/vuYYEKr6/rwPs6jZ+J7GceoFAnhzMgGvoFkD+uniu330d
eKOJ1bzYJxUt+U/yUpyEorkghDiCNnYbe29A8HWzSZgc91HBc3mHi5BYV5a/JkDv
ZGdwdk3ARIozDfERIhs86YdqCJqkei69pbO7YLYAxJTI6d534j3zJqZzNJwUweyX
XRM6Pdldg2SEfM2nZlMH6QLB4i27YwcuPijDnEFrSOSdhlbuRrI0nTWTB1Efm8tF
JPPEfZaGOq9a9UTulFqhltPwfnI7VsfutdsH7SN34+4lUHAWyQcGNhH3rTWtD/e0
m3il0Yz8/w6oF+X8zvk7OiEwcJBPF3GWUheYpfh3dMFXAoJPay1hlUVjVjjoZpsg
RVt3eS/bCCMTBpkpqyStHgCIKeMOsI85k9JNYR+TPEp7/Zmq5VuFmz6aSTT3caBo
u8O6EnDo7HF1dxLuauRNH89MrH3yveT0Lq6pZikbCJ9cC1+3KvZsI6eX5kUpWLr0
0/5wwXzPAPnHREnfNYdoJSK3reyq+B8pKTc4ToQAQVShSAvHh1JaU3wOlCiK5Rbg
jTBhvCW7DtxdxfAGBY1AtSeybV+J2R5voX46BWnfXVwZ+gg4qvT7TkRXskn3gtvd
ZSR+Y1aOmh7vSKu3fZwCBBP4h2LsyuwuJceEoDUSVYhCk7SKxohCRKSk+5d8c/ZW
e1ZnUQ/gYxLn3EJG60ivPR01a+6W9FmhIepTjS9UMfbVF3GZ+B1QFE6UO6zFBSrc
tkSR17IsDu4WlrPwXfLjkaye7oGOt+IR5PlzNe0LVafo4XGpZpmNgJ/rd5bwvMZs
Z9GiRswJBWUcuzo1TkfVElB3pAcR0l0m25BfwUldMvBX7P0mVYKDokFVSwM1//Rh
IVe63KDoCKKDdjAk4KKbSLMao46tKQglXivBj33EJUiHVUJLrPpJgn+sgeRgf/0h
n8RbNWpTi6ViUYcpzqIdy8jWuf9WSNAa+OgehNkPySNUBkbLRTkCG6Dx3akf2IZ7
3GVj3MIYG34rB9YSP0r+BhLv2afbyc5IlXXEB43mSa3ckBINrpnl1sjYG7Xq/JaZ
TR0OhQQO8keP0kP98Cyj7zW/zv2b9UbcdEQi7HTFkkHshnQuCgRuVAWFVSJyG37J
PNB1zRgGC6X3kq6pT+C1YSfd4bD027Lb5fC0OCYjHMAf00ARd7wY/XDwz39r5wXK
lSBF6y2Ofu9cOPQWppJUN2UfzMQJhR6detv+/qboGzfDhjLVh4i8oIGd40Ld3+aY
AKPJwNPo84OCzBAex7mihSlBegl2TKTY3/Um4CfHTqPdYr2g9zrrL5R/2tCqjcqo
h6DXRiun48zsMsRNq+QsUE0mfFQIob4ULY9IMYqRIhib2bRmeZJ4qDio6HRhrnhG
f9lPV6QG2VRMcZz8ALweMVO4hU4l9+SozhpXlHdy+60j7ldrlO2W3H6/uS4WhFu9
P9k5eOrDLezLNQdj+iVyIxM8svFFnJodsIc1dKQwFBVnRyz9jNpGCpZE7O+JINvr
BJWE96u3vM5nq7q5oZhuwnDdvy8YWaNR8gj9AIyXY6YagOf2zL4DI8xTZmYhbf29
Y7Etl2vWHXuw4twUssYnFbwVfmiOqsSL47fx0GyUQOOhsV1aHH0YlbL+iZUTLu1i
q+E2udCg9nYoWDnBrRygWyQh6IGLc8sjXGZa3SHrvn6NNSZW5ZSoz/OoXBOi+d9T
VUs4zVPfgtoiVm9diLyY85AqfbKU+1Vy8Nq6wDSsI0OrDhakO2wViI1FFcV7ObJT
NRLdCy4TJ+cxNICaCf9bH0N4c/pnzpZKR6AEX9PyTvJ0MQJm16+CT98wpqUjlAe5
7mWjw7HEkC0AUY066TdEcaEwAmh4WIHpnKPQhfw5yFiwCJPtQGhz0iXbZvJ6BHTr
R46VOraghrjsq3uH0VpoQ+8G/X5s3KKypEePJh5vrijWLkCPX2Humsj69MCYVJLS
LQrKKP2Ie+ZbxQKqaf1WAzrcfcTOdJw2O06U9PY5DGkNXPfQjSDvx0rNO37nseCJ
MLQepnG6XRYbxdVEaPwjq4Bx2bTOL+JSG8IeMp0HVaz6cmBP32BKJgF2+27Jat6Z
5+YbYmbjKUmTwjgF7sBKmxpWVjpQm8Ia0FpyZw7x0qq9AbQjHU+AxBrtsF9YJIo7
h9mLq9bQ4Y0F0yh8gbWYl/njZYL13biOEyRzgo2xXFxk6/OBfezUQK7YGdVBoZ84
7Pk4b+5BrpxecjGq4PTNg/vYvhlxcJLkq04iuQOR4Go+cueOrxBvTgnIN4yTQK35
GLv+yjDWf6XLNvdiWIIlpM0NNXUN76ZsM+I3ww7krRv4bdx4zsR8AE9WQoC8fJ4E
VlxpQp7OEQVotncm0x0RmYiCme7yxbX3KoyDzfJsV4QINr/foOSmxuhzndVzncSy
6TgHzdPmdBlkI89ppVK2Wai9fvhLZGZauGV/Qtyx4ZA5pSVAU8UFl9lLvk6P+DcX
+hipA8/w3X0/j46eQGiGcwu8rqa45nph0m8+VbimFtZhj8sp6729OwCVwGvgbr5s
SU1f6jhMjd0u5XSpVfSEgST24rDPwVH+P6a9yIQS8nquUMl0E54kFtO5nik0zJUA
pJ7NmcKkZ144P5YNP9Yz5CoZ0vQdR9M6ARqgoAhgXcRRbgWgDqjKOWjZPMaaG6gF
WKHAOW5aZ/gFgyVlBd0qxbyeIxpWcFzZnvmWZF2mTP4CIooSJz6H6BZqs/043p0f
JEb5356xc0a2q2yln2VqUnrckk8lBQQILvkazzxQYhYPz7WwXCfoRDd9czmMjRh8
zhUmNQ3AwE/vu8hIlrQ1tuYeAsSOUHg56I2DjiivKR7kahptIbdqsLSAevSTjKER
ZJxgICJIV7SmfX8fkZGLCAkpw5WukWWcG1Eet25PyLeosDXQ4Fi/402Vk3TVwgPb
QSpB/O1DXdP9x3Hagut0R329STl5Yorto/PFyZDSpKpaVBXw4/bo+H4WWXoabYsf
pXfohWYSdwzLQVplwypVi4d0hOKqlKYjHfS0vd7qUV++GKfpg0KszBbvwPTILVNa
VLC8MSt91HL5b1yzBghcJqPy0AYBgrJCvnOkrbGnkOC2ROcQf8gs/NaOv8Y4NkUv
/Xjboen6I9aSjPGd/NrdRMJL9iVEuySEh3cSYuiJbaIBpl3gVUcBMic32izNICQu
EYV/rWU1h5tRt785U9q0Vg43WA1vohoFDsRVYdDwp1wtV8FOdhxM+ipRMu4NELVg
lkQEhIfgfn4E+PwoX4WJB310pfSohzi2BsfPLEA/tEYfnRWNc9zArThjLgdvIbZT
DCIE+1ZOMl/ilZWWibBbjWWmKRMecu6dvbdsPq+FEyd7CabjH9TH/Ih+XLqhfyZD
FQ/OFBX19mhG6XxLs9J30YNHSrBzpzyu/XtQNaFDYcT/D3uAUbSQZ6hICTTEnWFh
vG1ltMXSonOc2mD39lWLDMRo3pxZhUHWFIUDDYnn166SD2HiO15dp0MS5mozpZmF
ayhaKQo+C4S1RDkFANXPbIuB9kaAx/HSTev3IOfJm7Ef1SbOIoXgMq2qpfI9sJpS
Q2vOz2qRvfZvmWqkPX4+CZMfOnAPJTQ8PztZphCUyqGM0xFMoX5SBt/53WBqslHV
+lPlye7ffK7DVeuakyblWM4uvFl9Vc2Aj51wdIbrsgA8W94Fr1Hhrjj9Xg+AYskP
u6et8AZe/SXLCwdRlUkztUSe5PqxIN7O+IXFfJLopChfsPARvB7KFkoAT8JHySgw
e8VovOpjl3UU4aWVJzErYl0dOTBfsI8u6KOWXxuNd+XE0DYSPISTm0oZcNVPpxbs
jLxBilwL6dqdFyQoBDpPVOLZbD2l0k8M/EZdapMhJney8q5zjh61l1p+OxhwNGEW
1bJzlRxZFrNWMjwY29AFGww1pLgyz2Ijk1GYu0cVuvNJLOg5vPb7hHPfFFwveSJ9
jjtBmzYW1uu3sDzwFoTqEaUjtrKCf159xik0NL0Naw9DYral/rBAEyzIqTwnyeSB
f/dwpJorkz9+2r7T9rYpvelILkFkA9mBm67up2aGXvmqTn1MfsKft+fbVuX69YjS
7cZe3OWEkfps16D5i9Zex8XBPd9iJTfIM2SZhzhsFylCMB07XskF7dJHJZJ+l8cz
C/PICYVDqkE6VejQ77x1MOxjcY4G9Aqe5HATn10wIi6u+ybDa6Z2lJI51vWkIbRC
SM2UOmXiD3MQC1L+PESwMHbbUutw0W1Tb7adCkbLY7WBEeMJbqXeLEN2EksZM2v1
d6pfDuOA/M71nS7oSDL/BNv+G16R1l9ns150KIzs7/xoESaaUU27okm6sk4HYOSz
qcdVuk2XF+TPJ0pxvoUzEDzZI+vdQQ80OqByjiiQ2qd5S0WfjBm3O7qbyx7MkQkH
dk+/8yGveiOpGMNh3N3TucAsF738VSWfyeb48moz5CTwsXRvMIogijqxpIFGDuA2
n1RN0ymdHUFXS7w+/5IsgTKEVslsafog+TyKPuPjDQ+ANQ4xarPs/tFXWN9cb2ch
p0SWH2KzYdEkJpqPUDXtCDooM8Sw37OtnQmm3bsywmYdZ6UktNj8H2utYvluRc3j
nqvlcgi3r5NUeIzD4AtcATmZN4+/pGX1kRBZpyPJwFWXsInGAb2r4jO/3/r0EHgo
E07ye7sfgoDsoN3CcsoCAEDcuPlpXq2ioOw/U68prv2ESPs4LOXRwCbyi9inRoqQ
35sjlpfj3F5WrjB5svK/6a1wmuk6K4qJXgDW6vSXGqf5VsbFs835te1Kox9OKZVE
9tic8c41kcE1bHjvbJduv0/X19U6rTKjbV7t33p7JwSMwYbKszXyovlbaB/dwRAk
itJ2LDxToa5A4VSLSgktOB4HfxnKRI6OD89UYecqzZDGCWCUhdD5IAihrQbvOznB
sDfE9/REQOsppQfb81mOInGphq55OPmNKlyYScbHi0dUk1VyN6a6JM3PiclgOt00
iV+TK783hHBVIG5KUa9QxosRizD6sRq5CtUoXI6O0wstwfU+wKeARV3dVEGYmMHy
oyEm2qa1rIrFDo3Qa7/3RQc0yfVlW0MClcYA9EdK1HGJ3iKDHeOO/g5OIYuUbU9g
BL8Zq/f2J1lKuN/Hsl8A1uhkbWjlzE/eXCV+bU8/CP8J7G2TSxi9BDpdGuX5+oWb
WcoIe7hy6oaLyVSh9/19XZFaZzRjw2Rkfy5rkvXLNMmsF7xs6zzdw1CPDtTVNPQw
zo+GXUReZWsouVX7xApojKrWmcMs7IG0GZWtAv28QJzRTJvJOguNdE8pKTeSnp84
1jDr9ntTAmsDp0qL14sSCpDauJ1HZsNeHIhyC11uWXNYll47N5fXzpq/Oocp3KVA
ZLmQkednS1n2mDcOnDx6fXTFEqNLgUUtqjtWhLh2BhazM5pK8JcLU8mVKKVGBagX
bgwomiJeR+tnVHIC1M37gbKV0Im15GdE+Y4puRUntvzKuRczFLTPU2+RPTEQh3JI
1RbaPqFOohQsqHZ7x72OQRfqZIhKz4SI2hx9GSlQq58a4x+aUhb0TJBXO7sWzcSv
yf2SYwbKIAZeD8TxEO/nXJ/MEbOjxbJgZV9tisWz9HzI6vrrC604Ls3KMFjB6v9X
tQwTtg9cdhP79SU5UAAsHeTQ6asJPg9Odq+AE+VaiNoqHExrmpUeNlHh5pI5k5KJ
tQBoEl7NT+AlVz7l+hsrZa6Xg5mWfyXFQMACDpC0wLRV6qf7zDBF118K920gxzO6
Mv5N96GamdjUyto2LzWKgljDqCpHYiTwbCRC2RUwar6pJ3z5KWfD0bskolMZx3pG
B7OM7eZO4VLGZcZ/jYunzMm+2JiEIoarjZPJN5FIv3quk4o2NXG8RTB155oACKXu
cL5YDSmRp9L3yTCujR1HNW+w3GcXQrB+O5td2l07fdAR9DjGw0JgXQFN5QPVdpzD
P88PlxcDbFeDsCcZ8WE5hhi4uc2A7TVuw1xoBlMnV8Yfp8AfVyPQY3eAto2Yrahd
jBTMuNZECw0pJvttxKBkP62E/CYeM71AuVK7EGFWDYPvbMO7hb3DkCcF4eZD/jRu
v/AJuLwTzwIsgx9QbNHKgoeWJmoGwWknt4eyMqBk9JYCgXZNoAL8zqLrClj7z84C
MNp9BgYi/Z1YqW9FFM7R7wHlcDySc0JhOgWCGxHjYCihHo28Uff63fdUyN4PImK6
z0Mk5Y6cM/6OpWCvTDw94zkNJKcu2eCmfrWVYMbkqSr14N1q4XhSOSjmiZzLw+GT
ZCA/KAHE1z2jub6mISYArg+k7ZUocX1y74J8qi4eXG4roKEtVn1drbPVFzeR42fO
UJqLQ4OBEa53NSVuDo1y1sRrF8/6cea+7JyGpzAESKs+6r9WCAy62x/j+JC4TcQT
eo+dePJ1ohai6QQDSQgnc9QYLVrOIjsb6iQqAa8wcMz0As6Ga+0H168I7V9UzXmM
K5EbFkn7mXDAKvam79xl8hsN44tYOeIWKuNq8DkW/aQ4cThqoQAbyeGLAwzTcAxJ
/llv4tcbfmKiOYYrjd1HKMP03OH9e9Qr5xR1uWiB/Dt4QgTjO/drO1MvroZniNcL
39whtv9y/rM9HayvWIsy6GAqGtwAMh/ygQQopF1kH8VefnzH7NLzaUWAUJCd4eeR
jjz4vWefdmACwPe4sjlbxxqjaViaZGp8P7lQz+FyWh4fxYpy5hbD8bsgEcU1FipG
Qkrx+NFK6zf87zWsz7ajG/1DG5/pCkf8jYcVXYFdLC1XAIgkt8UEUWb5/LOcggHW
LNU/Ol3rNAUw31g7OPNR/bXqf2iQkJebLgdjkNxTItYbxsU2L91U+ecIbvNAoFqN
o/T8UNOoIl3/1tQe9McVXrG1TfZv3KBMGivBv4qdVyjawTNPC2lAMDRKKij3i/F+
A+kDkTF4HVd3akzd5drM/PAKEkmjcpeINR3q2gW5uSr0PTbkrj7TuacTbczIxt5x
ze8hb3QAbKUn6Lki3iCfJI83cSpP6ztI/Twxpsb9q8zO5AV5NYjfp/eukF8mH//e
IAu9SXXjxnuC1htTCVne8jDX68J0mrS1xgu8CxuTYnIki0BuD0rkUagT7C2ZJnKN
OcU2EV431fr/0j3enE6HfR+KTmepz+n0Est6jdKq2gCcl8cm0VBcdze9Bwyox+ma
Df3Zi9le+Xt96ZTloxNCsCvlEa8X+nBSZ6QeSiWk6CibFiDfMkTeXEOay8FhlvF0
SCp0ypPEJPtqfpK4tSWRxfXpOXOP6wuzF/3Sdluq4BVAFlQkvdpgwOlZEwabvLoz
7//3KO+OS6btyTwLz7wwQ0T+kwoqlO2zV0lMvO9srVdGFM/LF1DQDsLH9QT4YTxi
gkkGBVVbeWGE/z8ixvr5+EWZP3KKXXXxNuOuiIDgBYv+xRe2ySwaGS41LOmGantB
8QlQXSDGA7VELImpKQAiYsc0aHJ1i+Zp6X9r46JOwfqaLxyima3dS+Mbf6bwCdol
csL4cr4BxBouSQw5w7OzRwhX3wSLdnpTQPLxB9Bg880AbESCFPK4IPOgmBND5fhK
ddCIk8r4MLzDR0rfiVs7TMMf+VCU4cI4bOSZnR071gI8AnXLv3VyuPgGKNKErV0U
KRh5RZdI8v2fuhhNLWz0zTX/O2RVtwEw/sihAeRkZC9JaEp0qyCPZ7pJTx8n0Bzd
8TkWPR4eLeUTtgzIGJ8nZw9RBRK5+a0gkmC4SVfUAbpm4WeFFkPJgiI6wfsIJEaC
/X+laygqQ1s/WD6r/p2d/7FgPkiBFJMy2ZggZs3uEvib+T8Rm8GxUY/alyrXzBxp
UcSrsChqKcB6UsN2aiilxG1+EYesqlxTt1OQv41uR8xqAFL+qDbwC3XhGiQc6Avx
ueUDF0aTWHzW/IZgBhCFxGH5OoiKMkhtHnsEQ3jNHbpTuNnBwwH28U4vIDML9GOz
rMYVQ0cmg6LaSIc/+UHAt5P2El+UcvA0unpwpD8Zfuu863B72uuKJo3lySGzKygS
v9nGdNdS2MH9Yl8Uni1LvznHhTko+HblZLx6n/OalrfdFsaISs9bkO/7dsfAXzDp
qsHmHFSAHSENy5dhZGnKGmbYuw5ejnFABsJoW/2Nqn1NOyM9dkpe0y58y6ecEvOJ
mEDeqz2IZ+60CZtwO0hIxXx61vvuDqQFMsx/srRwLtLePk1WBbQ4oFmHQgI8EwnO
0isvPLJURqzxJMM1jAoPRl0IeD4h4AOgVsqNjvKs2m90k6NwhKVKjupXHFoPJtM5
1wPrzGpUbG4jDQTTqUkpJzl0uq4sUuxBfJCPEYtLypGxQqRA7BPtTcWs0WZmoHS5
PjpaSe8tnsur9WWEycYpzc+UtJr61NE9IS50k9WfTDdrldkYYBDpi09o7Sw6jsSA
ct0jP9zEyt4HymQUFK8KF6Mi+KSsPoZ8PQ/Ia/eGDaHRmE1gXh1KsIXF1xxPpQLA
d+cJEM9AC7943xwgG3JsyZr0idTYJmULwzsdrlTgU1S0aZgLyydGdtAnKuLDrNaP
EYkUWTw50L6WWgshU5dcjY2P1YN9vP3nuQqwt5qC8qB3QvX5XW0JxAYci5H5pnec
npWLyXyJqsslBFMc3//E/CvsvFo2cNkdHK35z0VVb8RIbXXSMVXRg9z3QVpgiMfi
Ohm5Fjm18DKj5GuDnSGtcpJZa99tUqYjcYU49OGXsd10TBIKhQBnttWd4xEH7U0K
AXYC2yk2gCnMTWQnX2HfIbivqblY5CAEcw5L3we0gNgubS7AiYGoJ0YFFkBycVca
v28k0k9MZKJcYNc/G907BwgUgJQ6kbyx0XmT3NXIs6r8vT8Wt3n4qu7TmYqODnwr
NgwXy70IhCRXWlGqXpC574nsKYlQldXHALz10dhgzA4reI6w3znJ1c4oYZtPy+xh
L6t58M1y/EO6XTSk6ZPdo+65wH/XyHSSSqpPXeIa/4qX8BS0MmCxIdiqXSpYr8Lc
YqWZfZ/REhilPaMyw4xh0AVtHnFzBR7pL29VfTRZbKQPIwrOAuISRX9oXqlCcVd3
ts0luKmWWspJhhzBztAuKA3zm3FT871QnWoxIhtEEpUUfLLmAo+TFY9mezyXhtMD
StEWnFQD8kD03NrntBESXca8MzrkiB1rD5JFcWTARfoP6Ae/Ve7yu/mh30eIPXgr
nPdoAoXFykhSI1VzWYxm7utQ6o5IzJplJ4HI6R7nGpxKQf54P/7EBmnNkAv9FVeo
6/yBeU6WCikbVKRN+zFdRvdGVUYM1YNkCPwvSOD+fHSPwW9gvXbUAfxcSzYTYsAG
X1Fah1c9elKXt3HRRok3mhD/o28SDg22ZrJCHbpijFH8xrcGU0IzFCX1Qu0tRQ+4
QIXzI4fj5ajH5Gweb0i8l9J+dr+j0c0+thYGpLXYnLbmvorp4aKfjwPM8as1fpul
XQCrJfiTKwnxksGrnqQpuKqgrSTliv8bzX/dkTqrz49kCHJjoYhJKWi/yiDIx+eD
OWhBCZkp/NIigYlqn5tmK9R7C+588ceXQXKyZu0HLZJuCgmB/fnwN9DMORS+mlTv
ogBSA83QS7Z4A45BO9rlKtOy59pgKHfKOOX0VTPhx4ft+9kQPL6HoFg6z9DgLD9c
LooctlhBNAo6aWmM3KRhdZjZbM1zizwkUTDJvMu4yBlSax9vHqklIhJmLJ9yIEFE
eKgo1A3EMlUO97Yruyo66zKSnYj+3bbWkwV80lFK5tsldsKuOyypnXUrwklU72Fu
dP2pz40di7e5RZPUT1OcnvTWGv2yMu5FE9CEtBh1etlwML2pcuWyja9RVfyNQytX
q3ywShuwn3G2F/V9FGK0JE2+ozEw3CRNBgca2mYcIUJb86xuquHsvh9Iu/bbNEYT
h1w3SvluedSGcDlcMEce5FJ1nU96P8L7fitsnHankacIC3Vzzau5QvvjVszrTUjY
8424lhc4slY08WYRcNmyO0+qI7HuVA8b3vFgUl0OdI7SmLI2iggleCYHm03L8cIf
04ny9XNf3VTMGpvJoMslxicJa7fQnqy1cANQdq3WJKPfg8CRaTvbNJXOOxKctBL7
RNT3KswhsC2M+lhNa/tQ3uJ84aEcGfjgVO7j/YVV+bBCibMABmvArgdTHuWyb41k
l9PQe4fN+ef7B9z+JC+IAdUAp2QRWsWHBuvMwe5iUx+S3zVn8aDk89nwGTzw+cNB
g98YK5f+wc1kyOU0rq45WVrlXaHpkx6aqVAeROtiy7OTWxR0LWXhRYdqBJz7f90J
CrOsY9Te2T/L3ku7IUk0PTxw/SQSGYmeWtj9ef4MBdRSpfhMRYkbIUIlFba6An/G
UAhFIZSWrMxcVmol3JXCgY0OHhuAYV6rSnW44cR/mKtp+eVmF3R+4/VfXyCbFa73
0Ayw8+lxc9fuMde2tRWH/lcE440MM4eW/PzibpzjYCDqJR/VS1nE62M/j4LSbVCx
JMH9T2SavfxOCCGDWxFVbsBkafMv3RGawIw8JFYIg3vPNW4RiPVE2JZdZMkBGtxg
oZjY8SKnwtxN90YEqSN7bZ2vevBQxbAaEP6aSbwA6K9d+jdcuHg6oCJo1NSG/d27
m9cr2TEDwdjYaGmQvYLYyiO53JZjQC+wM0S/PKeeGBU3aRXsg4DKjv0Via+jXJQ8
LkNIcwIQNPqquyQScLqW+KIdu4wMmX1n7X0RPjbwBu88OT5nvC6JRHVdJiylzNbh
AqKtX6JVDU4qXzZtqK4p/BNC1o6WYbmuseMs7OCt4gbTU/YlJ+Oc+UsW3wlhKL4J
lrkB50sRaar0QKmKOPOMK9sIrfzs8D9HDcjKZwTOKSm8PRC0tRLcM9AV0aScAlQv
w3VhRPaZyxBdRNT9So7cP24+Ch5c1Gl0bTgSnXLlwZ9ECvbe3z3dwh9gjv5EVFCO
6VxCi5JYoNuKLLB8vKTQPQiPxRO071y7ruBsvMJhoJrfutjHnrwd2wrH1Ot02S9s
M8tXZ2r2+yH3yaCIpYT5XFHUij4cipkdRPBT+C76Xqrjx120vIQbbxSFay8yMODY
OsHyILPnAePjmhC9dMcvgpKL8LZdFwHmyQURk3bfL2Ro5143NrVt0smY0ZTCVxQL
EPllvP7aUn/G8Z1SgyCA89K9ixqaU/ylcJs8VKJq7/uYeeUfDWDvRBDD15bBgMGo
FOufn4tJGzMUroUxZUA+jyzRLa3GER6xXh2UX5BZNO63/rNYNPAwZxama+xlMOX5
bbtV5pUuptN5TRAhrL7F7IF05wKS0Zjo3Amivu/V+14+gohSmz9ey1pLn3I3TCuN
cdOCGidAkZ0tgNliS7yVk7ZKWGMuDzRrWOVQfknMLhQtreH8u5ojz/MrClcWg1Dx
vqTHXbEmmb907ckD65Hw1hV6A1RXSWRRHKMExZ49875oKVKrMCBB57xdQyRiTGAs
4OUgLeZRvZk0vK7Z65psR5SwS8F6kCQsXodes3rBiaHxriQG+2vtXgpsNITjdacx
WTwqAaRUf7S0MrvgrrjpF7YuhEFDt3RVqIi9aszImyh3KRtCRAFHoj+wDfwIZGne
0GceL92REP0Ycue9QvWq/m1Wq/N/3sv0Zzoi69qzTk4xzJvbcsnHdbR9imbPOVG5
lWvfI2ar38p2IBtSivduy5hmImR9jLaLiX8oN28LJwgud0z4eeQAYtUsLfbdCc9q
1ee+yGWafMIFuKimueShDlMNWIA6ps40cGEWVamJv4eRsMxKM31Rjo5T/W9ZBg0k
OIHlv9hqhCihl16wGtVJ7fL3UJ5sgdRKwuW3hczPJ1TGRAxCsqW51LVha1mtSkQv
7tL66H/pDRzjpleI115JDTDBYR2tooIQRmBKeAFw44UFbS+/p8POJJ2SHr0Pv2kQ
CYwPsPCRQQTU5X1ORMRx6/ZvoHPsH/R/QTfLnSp8bHcaE1cAK2PtPe3om3IO32vm
PiRY255D3iMUWSP6lF9gn6V+WnS0daeJmbSw54lSuxMCn67yznyWjSBNSyYEyf35
QnnCuIH9CnJ5Ta8vns/rbpcfMgHAWicTM4Frf/+xw+EVNeBRrZ65OcmLQy0KNW11
8gqihVcYOLU+HSg45Zu4XJ99mupDReAK4vYr0mf7qjzlvOwlO76WKIqCRTI/zfRs
R8/JYq17ZG5pp/FOL0s6IJ4X24lD6tV0F5l68gkwhjnH+qjfuRfycSo9TAyFz41D
jNcjuXWcal9oSe45Q0KMEKpaTPXrcdO4RY8I+jvLONkwExGkZ8lu3c7tNqJt/5D7
4mN5JyKDkibcaipAM7HUcR5d6RwNGmuk+1B5crSXLH6LAQ2fbPkQD19aitZqIENk
/h719RmpgQ87UqDeH879txWRIgAnDn6pxtH7KTD/0BtGPiknjOeW9KWgyDrcJ9Q4
qButvnztXCmahVPIlh5Nfl06lDpOTjzixWgBRIizMK0t3/l0LneAvvakYBHJTbvd
vv311a7L6syOah6owcpDI+LgGRUZMzL4GLeuTgtt177XJVpmLDrdbyLzhPP0L8p1
O2hJvO5Uu78E9kQYUXqODDuvHTrO07BsSVU5lJ8yPzbs4PWXaGzhQwqy5TW537/J
WV3fELuv66iIfZyweZFNsLr3+0GTSefkJGi3gaHPRvXmVyHCeyGntGvO4CEkoFgd
oy64oOq9+i3VeSu/0tqQ8p0Lf6iVE8jQLw6SOLdtUdQ5hFGJUMzaR1g3xB9X2G8E
pcIWW/Cm3NOtySfyNsQqYge8T83JpYx95YtxAVLlbpkllgFUlTofZs16YhG6xe6w
2nrz4t02Qc8YqTV6PPRifQmlaP8ItvrxbyRDIX/4iOrs5zGOW94wUp8tS0p4aKCN
l0Rgl6+5H4P1jUAWsF/PfCGncwz211SIyffalsHvCFuECxQ8HtT+mLeD/QhjOuJk
5XuI/mYuZ4fZ9VQnGOjEmYMigPIoVH4aBYdWmfETLAiDchD3kcBTFEfXV1faq8at
TYM9EG/LrDnHHi5q9l1yFIMfxGjczDc4rxv920sTUZCLXhDvEbit0f5qQzai0NpW
DlJ/s5OyFRGvsDORXyfnoPckF+ONZfslnTLMK0b46faWIvj836SC8bGGOZXe8q1/
S5nIAfU3ACxyykk8QY4FmdFcXQRF20q9IdM3hO60E0T9p6F3Y3njRYzRdpY2tW18
MC3T4fQ+2vHtQ3Zh+yyiZo78ZkH0iDtnro3RTGGuEUQ1kVmpcZ+Rf4aA47FLWLDz
MWOhFLjE9nEVInGJCOQ0vnOYcZk+cCqc4LL/a1/ITjreCrZGcttlnKH6bBHPXitw
+0dB7aAj0aSemIJWHTxoBY/Fgufc3hhPuetO3LvhAZF4TrKygkURgyQbPhrpo2du
aZsv/v+JOTsAHlbPRovX64++JvgmyyotLwYjjMqAACD8yWYnqhb4LBKS3vh214b2
Nx8Rr4JxdWsPQV84UlNNlCIwT92wYbmny7JCcPNylzkpdRh7bwyf/AKxHjTgZFUl
a8KMHpeFS4bLfR7BDJGrY+VqWgEQOnb97QPjzXzXb6xYq3a3dcKCqeFUnsN9b9/P
jjVprZwCUsuxe5L0p4vzsRdVIV/tMBm5O8QCH0WtR4DY/DKx8nZuSfRr1r1p5ddj
9Dql8c9fhxRWd++0SQgF0eJhe+BGuLBGdZU+qSYsCVce5yzz62NWyzWp0Y9ogdSX
krM/38fDab8S/rc5YLLy/dCCOEuvsFAOFFyJGPIlomQ1WJ9RrjtCYmjJPU5T+86b
7G45Gu+zC1xbfaVNPnNf8H9DiSNGDXQM8yyV0jySv+vT4A/etuAcuTLBfgRwi+61
oqeE1URqVY1fNiOYp0EWpRbG2tz6AurgnQC6hMOg48CFYn+ARBE0rEzG39sKpNhT
qOAAdqD2AQotDzZIYGSEnEI4zbvWjJUXaDqFAlBNWUgDhhAlYII7R6WAlIAaxiQ0
fHdwHstOIlTfehpAi/4AJrQXFjnEwVVZQgslwFiPC+MtVdj11TzCVv7fxkGTvy4N
QvgDBp/Nq9acdX1pNsim0RqQzNoLt69EdDjzmqdyzPgG0p8uZOykGp328gYhCx/t
eu8psLPsy+W08NQArfms+7CIoMqTRs2BnIjqYu/vQXYOq3WI63qBt2+Y/0NkTYsK
rj/PJ0qqg38Ji3r7iGELQaBz/c+/JyBMubMRgXymIfxKbuazjA8+9OWUZSvcUD1O
ynJJVR6glaGmgzYFxCy5GrTytwaFFqDSvJQ2/xc+DvO84Q8vq92QS9d50r3Ja22l
zAgueUm4dmr+PT4nsNbKdqlaBLXTnTECTlAtjie2XzszZvgZH+UxUjSdrEITyRW+
sUCVdEXUUOYcJURx5cF1HkjVHDY9dMH7oYQjCC9TfIEHa9BHJfUYEjZd24Jn8dbW
FBjWw1OnwQZ1FUvP6nTJu/n1ylr9VHOXlyuywHw7lBxpb+jNxThSmqWMUErUQET3
plkYti9TX/eqJqNT4cbhOY/wV2d6mgLX8hlJsrpmbVLAgfsHHu3nM1z6yfi6hnK8
0GqQw3Db/4V12NBrUUrwzMCnNNZUdItqsjc5k7p9im7yhVulbcr1axGX5EdI2NM6
QBPAltumqSTaZnr5fMMwTCe83L1+6zJ/KxsP3r51SZDa1EIJmvfbQExXjs5i8jZG
OmwsfIRxJjX30soMgDeVFzH0v1wG5vsMmoDGGUuLFH4YlRS+XIDmfRskMetaA9qK
IF/2UMF1mybqoth6wS5lDY0/Mb20vOdH/OmeODwi3d7Bc6Kl8DeVFpfSMUF14rYG
5Y/6u+ZxDLQWGg93f9NAhoK08KlPDpriDfGtaFrTwjut0yhrOCyD4bkukaF1xv92
L2iGmDq7qcmQf/emIlKRgaY1z/bmFPhT8kIFiyqz8x5ySeeuyKQ3T9aRxJrlIASZ
D3Sdk2gG0OYkYdZ+Iq/cZk+1tB3wbm9K9cqJw/hBhPvjYuknUUEX+0a/wNz95uEI
dv2I5jIu6C5vrD0LLgRTioQZJXE6ayEC5T5ooxFx5y6TPGLg4PWhiApEh1EuiF8F
s6409MsqhZ/VXCTd81O9qjnnm2V9rKknafd2gtXMWL5eUrY+qPnx2Zk5txwgqWBN
AvieZrybnt7te/KoWz+iHZsWjk1fKBtLmsVIMTIF2dF8FICRumvWSmCX43DvVwgA
hhhjIlyEj7qnM6cLz/PWkumVEEDMSObUGpT+KPxXtQfJkmZeo9EUxdpMjK+fx6Hz
FED07sTAT5+ivUcZfWJ1RNvfaBynKNiHBmaxPK5ujjjjhoj+sL4uenrQz+ehHMpy
3RWCRT/H5WTBMmk2vqyBH0V2Yd4QamjU5LoYRTU2yYkj6HCIn4Mzw+/XpgS/WtX8
lYaciyWo7Brc7OD2HKB+kWx6nXn2K3oVRYIEwpMMFhhTQSkwwqAZ1F0n3GGGGRx7
DBWZ7r5JMmDjxRJBOyIy5hf5LxWcNmgyg4a7BNK3Rzw/ILiS3PApdmvNuXUczAPo
ZXUeFflivvoWMHfYlq23oBi+Ai7xDPlEWcpcZtKPcAsGfMKLdoo87YawXG4nNVbU
IFuSBN6JJeOUnPX1sQ7+K61P0c7TL/nyEMVEs+6DKV9qggWqgzCbsgPMpy9NuLpG
BZTPar/iQeczyla//eTNpEtc+qPHEwSshTk0WQZ8jHmEEVe7i4K5r457zwbk3OMV
VPdF3j9etZg9x9qj8his18Weo8Uzb7mmee8OJu93cIY4F9CKLEU4boZcZ5TTU9oZ
Kj2/N0VytJhvy2hkxkEjBtaUcVkSJf7Du55NZeiGn7MxOYPwoWmGxA7br//EQd5D
7Z6XRw35fxHOcH5iuraqtX/wQlZxau8w/4q/NYAdhkwaUh8DSDJ7FWjZ1b4CfZEJ
wGQfjK2FeRsG3/onNCMTM2sv0pX0+DUXWVviOheVG6D/HXdqIZIK4u+bDhUC6wpd
eCKUvwiczBg2tj3neWEmlLRYuWQQGl99TtruX5/gShD6NnAFR6oTMWxnQKDlr6Yk
5TJ4T/HOdH6ryRItV1DLMzhi4BKVC2LrXHyfVV/yLnbQ+WbzxjtmA0P68bUNsAqE
S/VSk6BPgDbzxMAcB+Q3kylhJ+YUX9u/b6Ml3W3T8QwKbNxXlaLlKu3eJ7PLgCzd
iw8L+XXIyYKYS+qp52U9RXCrbugUycyvsbeiptmOMTAoVc9rJoqim3L9RTMzAReL
kjsfUW4ZUerZTPCCwisgwce5VUoqNReE5e+VI26zxyddBu0VbfukAAHKC2XzFsIx
vM7ZoxTxYcqohNKe8F5IcYyZvK4MHLQivcvziE5Fc8gTz+bN7+8Uu8PpQ4ismvtS
SzttFUssUKA9PA2kj2HmnXv15HMv8AHteDCr3mOp9C35MCwIqxTJUCaWAbs9Oirr
UeVK+s6Ohmp71AJEAs3oMzKKIOo+S4ZYwFrVipkhCbrJwESBEXG33z5PhZ5zPQda
ihQHnIgKZeWBL+NBNTuLl+aNRYURsuujYHw/OnqdyoOAcDE98kIOFcyBaoI5Uoo0
w98Io5BXfYlEpYJsLpEhN0NBoPdJLsuLp3E+pMxR+e7p8GyAM6frgBr928nxxvyk
9DLw5uE5YTU3s5dCTF0Iud11GHDpK2Ox+MJHals3sv+cWS8h+XCJWz9OVrATfw3V
J9O/V/XCCAGIWTAfPN6JDgKc7kG0QpQJkNVpayT0B7bcy7gJbRmlQxQVi02yGeJI
Pgia8cr8NroS34b7u6viJ7dbS43/BnvVbBjZ8WFF5Nf6KQBrodNUEXbKfn23n9VV
JqzO1CW09XnCxrdcrLiO+IvvNris629N5ImV+pTo1/0f9Hb2kYRbMjaGZ9hbdqfR
RVaidbC5B3CgMGEKDWk8ofndcGAx1aKMZ14PHpI0YK8/Q71XnGhq/HGoJh6vP+Yp
ckWxa7+8hwmL7qkyNBQZEPHOzaZaOjXnVNCiBuxfg/KmDnoq7L4KIrvahCj5IWAN
shewv6qwKzhTKtmQDEyAKQBww1lAtfh7YuM8WhU16phgQe83t5KqLZgBRVaYeEOG
W8XO6/CYiCjdCuQF10wZFre60CRdorFNy7FHlX56XojYg/jgp9CJJOGu54z5uGDn
I6FpzGhQ266V5oKT1XHeP1pVZ04/UiFElZff+o9hl7Omwz2M7E4Gcf/XCcavwKsd
1ljClcq3MtYBxQ2H4W80v6YEgoRfjik8cvT4igWGg0wVGjnip1o2AU8APEzIiFE1
Tr6s37/BmthslC7UkYB2iqfP0qkGrLg0FMocu+HO70VUD49gu4hbFLKZf3ByBQF0
IW0EWE5V/0Bro860G6goQ5fMy7X6Qzwm8tw4/Y3ZOkqAeUwQ4KLSUEamwP+B2zOJ
+QPH0PU2GxpVNt2Q6lu2ekKk3D6eWHoytvG8hkY6YKBSN8w6OGv3gpKUiutZOMR9
WdVY1aLJqXuzuWWbTtY/eNqscb6OsSLfHMUu64SGjVKi5inirLZI3zY2DKpyTS8W
lccNC8wtgRqDzz/mcxgc9uz1mrRTyf4v7MRVd5vWNOLHThsAusPyb4sAQfoj4EU+
5HkI1cqvcV+v0nqJiTG+c79NaEIBGRSqdkEEN8DFYFHHzJBBRQnthJiawi6TUx5S
DY9R+YKHtGG1F/+8l1aYZ40n3NrMAqz9hl1eZMA2gw97H9nyhmq0liaP0Jw2xdyF
kCd2hM99U/xr1VP80B958y3g9efJlyFt9Zw0ZfOauoNE3Ri2Gz6pGsDsnLL84wGG
UJy/yhUlRAon0xpvm2/0hcbUAG0vse3rawTbTD3P2HB1PdNrWX//Qn8F8W0Ng9+D
hl0mryEEImQ6PZDt2HRjygdNHSjPw2cwB3RPUsjw3hOi8pv+1rgUjNxCbIXT5vk0
/o7o1hzP0F675YztIq68e45Jh4IEpod2KBCcrDyv/C2x3jDZG9AOHtA93nQNDN0L
K+e1K2yBxer81PcIAfkzEF+a8JlPN3+PriR9nJt55cKUGVFBF/E2Af5nsekVFr7q
vRQr7SQlf/WDnZKnEMxGI3gAWCpuUxsNrIDQ1M0zGMl2pnYNH5+LskNfUYAM4t21
Uoq+VOePf80x+ZSdb2itqrTIqGeSuc7w/BNDvSPEtX4r8op15aIejOWxrpuLHXt3
E8Xk/w56XTl1RtnUK6f0z0D6YAOhAJFAVpTV0qx1kNAqcuw2PuamksMfa6yGguQQ
qA7EFtPZSX1kuuXXcPI06a6Rxr5E/rkBDjBPTIP7zukjwQ9KWMLA/IfHk6vq/UEY
u+3iqUfMm0rk++ZVdiRgSrXZwzc9iAnAzFoQd3gcYFEMjPhqN80NiKQyeLGW4XCs
0uwjmbGBMdQECS5XeI0+nub151Ie8KCOIZOfxStdKCMgfp8hLG5jsVqi7aRm30i6
H3HB7LzPafGXeK5P1uCmDx7D/mN8fAhXC/9eBBYlNySDZPSAcjcUcETsnB0aYD4F
PoYEY5RRcGmL+hqpphz4qX9hYdc9A0K3VZa+YXzZot4qXJ/JJiSWoPV/rNu1hYx8
A4/5JOoT7EZg6kiiPOhgS36QjOa7FDaB0Ehr3pfONnVXfqeJrRIx3qEhiniCtr5Y
lmxjKCx0jiAo69n0SewuI+7DrFM+72BhG/fZ6WlCiIMmGBjDsfILRKRARKRDtOom
vR2HAeMtFjekgszZW8NhGDwe+oQj1HksuQzB+xgwt1mg5thwJ+gqXZcgmD/Cxsq0
p+1R6JfLT1EQyNqjQFHbBF0x8iRAuLUENS9v4NQmsRoGmXwKmqlXIvHY2oMPuMf8
V1I+5Ix2lLg5KTP+pXe/W5OuA3muk3RTG8wNkWhGb8NKSwJit4Ev8pLS+/weQokU
6qAml6+PpdDQQwS0MOwiDhJunjhq5M6bzt+2aAQMOfKTO6ksjhPQbFYjoyp4LIGU
ZiaRzaXa+KdorfQ9ZQ64XmSPXl0BMZDleGL6Ci1MptzLzAV5DAEBUBWNRk0Lp/vC
u4nWuiL51XcPYodYQygmWDQBnLHE18bAIGncucclY4Wds2qn9/hSXUuOZh86auar
56H1w6DG6PgvXCnlhmXU53Px2SdaGoz2NAnUvNO3rvqXZc0l8gf1ypNHLLQvKQdD
MPP4QS9aiFbutE0WyQQ7W2SL+MzO0irK0du0NCzx81TBsP2osLaCA/VlSnCVxDD0
iP8CHLL8vJPjC3GgMc6/OtPkw+ZmuVD+vKYD1KHltzn+s8VMRcwNwIQ9HTliMy2V
txVB/g9GeatkIyfBiyn//TXsbPu2AGAN6jw6cAjIao0NgEfUKE1SQsI+RxRVdmeu
TntaCIJKFLN1i9f+jVus57GZRgKxwaKmkxUKeX/3qtOQUIq2OcKAYDEcgy/cVcMJ
9EWQml8nSdseAE+sgH0yW1RsdwY8CkDHs3GqxuOh0tiu5hp3Q2FUAsQ6t9X1b/LK
vHnl0DEzSkT5DzLIeS1vepPH4wcx9PrJ2f2k0f3qKzHV0Fq49tkYjSBLL7/Oqiso
X77JVGNvQf3g9RS7LGvw1hTL/qVrP/SuESoU94LvVH/IBKpI9auQL0qb63KgRE/Y
/GgAZci7KZWpjSqH6KmFC0U2RGQB6FHQrVE1GMXaLwFqW5RJCz3w4DF/wIQHeBgc
Ce7n5u3ch5io2IHAlVup8zubiKAYwfBua1Hf/Z1UBr5qULl+C4/FwX1xOR79Oih2
cZzQi2tJWoh1BYFtW2o+RSYyhWNC79IBpy5nHCyL4GYU/CwPIxDznz4I4SsAauUq
NJVmMSvWW8rSDLJPOEKfRUxfW9rk2JK6lTqPO3fJEFn50w09VIbtl/2C2XyzDKPd
buC1SuetTGKF8AItPW8HfQtipipLTrHpvQqez2TDqxtuVaoSEW+3zYBsJaN07h8/
TnQDHtC1VhyPqrmEzRjh2SCpc7qvdCq1DEnbGgCgK/rGmX9/52ZB6psVQm6jE/b3
B+b2ylmrWJ6dty77+N3nsHpKfS1tuufgPk718rPfzZbKKOwb3cvcYqSmVNIoJ9Rp
X8bCFtc7ebRlbqwOs3q2jFkx1GXAQP4YtNT7d2CehZ6mjazatlQhr7m5hSNsyp+y
g+CJpMT/qiaQgbzRDNJTuu6aA7AFyMpEzHXDlkKah5Nv1D1++4vP0quFjeby8fLX
rgqPbmrbNglJSU6rtEFtvfpzpJL12BpWp0Uh724XvtaGiz5CkpPptRCw0DClTUJq
FS+bix4eckC40jDuZyPsnyStUf0p6Ws5JcPZlZ+b+yahBnCs1ZWc4DZL5YOqC1AO
Sc095RLWsfYBdjbO77XsSl257rlsgQ2CkQqibkk+yOYslp8ruX/UA0U9D/HWzYSo
F6SJEvSlIu8g6te47dmeutiv04rLvrg8ZnZ7c6jnZJf6JfWH2hUXYOGGQW7243sm
9C1gYforjyBYZegBcLpzC+nPx7hqBd4vgdVU5keOY1XNjHCQi0m24gkcqRszfRn/
ywCtDvAub0YlWNMtKhjj8NyXG9QPnncyaztyDDVXVi2ZGKg2/rO+7xG+L1IiSvqj
tvlU4G6jE3fzCHVNkYUPonFEpVVgw70N6mNm2x2n5yt6nNa2gr+h9CCnfY2Nyh/R
LYJ9PJUFlHIbGHxIwPXkFc4Tl5OT87JmqV+iVkScB9gB4/WlOMYuSaqYvAX8UxUA
i1N9AwXkURCRjD/4kjKN+wr4UZKfVfsTs/2bEhWLFmM698Wo/gAW09rXUs50orXB
u8FaeUzH5xetjC+hM7u4w8g0HPJG3SSF5j8lf+ehKH6luAcay3NWEId2nep8xuUR
7PSq2qoNTFPMZrZN6dcJPGn16VerDZ9VajrgdBaSVwOQLVJAxZFLQa3CVyFg8KwJ
+fTuXkS3UmhNFxBeAAwAUpj8OAJiQZFBTgA0g7ZYF2S2CicbCSM6O1Qgr1qdHHdl
iShqwKi/ZlUuAUT48F+vAVu+XmS9M+8wZllrOK2zjHmJ6qyVv4B6ZGYQcsN3ofMe
lPV9KxzgP42L1cBJ+LYmbhwTOAQyrPfKDb1ui2YtWrpoSUKXnIsIctXQ5GNAdVA/
YVclzMSCHN6jUz9NSRSTS0gGvIy2i61ljYQQNFWQrn4Zq8ZI0E+vWd5A6UobwYZ3
8gvS7QmjUVBg40lPswoXk8tRQMCf2o/UcobKftrot4+BqAT9rqa0oaVAxty9ctLA
wEbsYhej12dfRJwNNrJyJmy3LMfyfn7EZp7s9BO3tXgnaRt2iHuWMu/Vlx6EM8Aw
fZ/0xHSt39jGy0oFZJCm9OFqgtR93dKqGv6F0zLEcatnFa3K/mVl2TFeT05+SP8g
+AzZK8H3jJrYBmwD69buKoHsLYLpis84mTuXNvMUs6cLN24DCm1jnAqjQWs97mb6
SGhwDnWacnE+pH9D5OELjalpWYaxSokQq412SGKVec3XjWvMgVDYDyynF15JCYwJ
nPtnu6nddAJiMS4Hgose1DH6ArBjkpC/Bwu4S5/aCvZ0UYz+MwcO0uTqGzwzNu26
3TRHfBo4iwAHmAFgVcRvl3oZKf2fYOM49HBkDdw9MazFQmI++PPajg13sitkusRZ
K9yWx90MN5pTHm7wRToqEBu6OvZfdtY9clpURnUPMsvRGUL/FViyBcOIbhN49nQ0
HObJvz8yNR0PcvfVRsLyFiv1BSjPrUzO9Kqp+WHLyRSB5wZdaoLQsc/XYlDMMCb/
1jNFG0MHMwmmLsgWVb3n2k8dCmllIcTsB77K/s+a067p77xD9FWNBFcOCrZpbn4+
Iny7Ijl0D1x0J4SvA1R2NgLFRWFEEwGvd++8O+KoVB6I4rDKozOGiPhTQ0d2MENJ
2nYuDIgMvtCeLGwcU8BZgFJFlsBwPeFc9shUd53KCwP7stcg0BSKg7l6pyMg2rEu
8hjex95wgN5PjykF0MA7sPrlIUOQ0xBBO5nnAk+SEA8/PlJ9F6ibCgFRaYctASHm
Q+drWxA39uSbv4pvvv/J0vXtC4SIgk2ClcNiLjiyublvJ+VTR9Ai8f9vSMgjWG4p
Y8zbpt4Vfe3heDQyPO21rLEbiT9evRrrkqFInBXYePJJGZgL3C0LcX67BH4uhZqn
JdV/gBeVXOg+ibVWm4ru8Uh+vFbfv0mN6J+HzeH4YxIaMwlalxy7ZjhEq4XqhEIu
Ka1To2m15eRnJaWvKXEqgsmtJYj0yPj+BH36UeEatE0beq3YZLZq0HP7Nh2rlogp
KpwY7fP5j0jD5Fy5F0mxqmG8B5KPkSB2rpzYTSCBceTca1ku48wM12XZkleFXr7I
P/wfo6gEE6u33fCLE+Pb7ObDEjva76J5KYidbDxp9fUcgWCe2q6kRvJUmvQ9oSd3
ZqPmuuGcIGckG1q4ViHDDxuqW/dDVC7UHMa0wpcMUTHAr5i9TXHfOKemDqjkXVhx
6db6qPDKBLrspYUKTdshW6JIBiD2T/RbkZ24iJRmEZYd1FNN7e6pE52zbqb0rEyr
Xgia38pDhG1B5PO5chwFbzvfN03ZQBijIg7wTmhSo//BaAwXX5gZ8N8R7KKioI9o
UA119J18kM9ZpBQ5L6G2AHxDL5Lk8NYk6/VUXy4r5EWhNbE4BO0CDRgx7i6QlobV
S10JLfkqGOLlWjpZxfXyw7izphS3rCbzsKZ7e+tXyzMrg451u5e/NVeJDfbPBDa6
jt68ARdlT2odrSSvZzDAluuvq91UnZZeW4rzDDvUD/+hrqlTDpu69F/LlxEyADCY
PC0jH/b/e7qSImNsPp9+2n0oPJnN9dw9vY2hpZz6Ag8XxrA+CHj/JD12oxGR6fQt
bjRNhZJX6OohQgcqWFmGTy0HIrEnryBYsbuWtBfT5rIopYb1PT7XuwSCHqn0X8i+
z+GNl3sHsSGwqgMJI9h5DuWv4VQ8CDPB6VCr8JXieJYezb3t4C/Vabukl3QKSEa/
UeSJJmPbL5dN4vwgJ33jeTEW3ZEN7dHjuAijbyJgfbLPEntQfPHnbFfE8SrSn+Ho
4JgP5JQmpgGOKSwufWUB5ETU7amuA8p/TByVEyJsJ5FDSO5IhmRkNy+jeWB6stRB
hIantTQ7DuWcDrQsZ2WlpI33+Lh294xTfVbi+E/dMQluYrR+kZVeSNCI80qC+dRw
mcL0D4ioTONUGI3iGa5pQDkhiFziDSliPM5pnmMwxb8vhJcPyBeVVZglJzr1F8op
e/EyFzJWN+NvB3LQSruKRO36/ryvhQSZWeenXlZDztjilTKXH41HHecz1FjDWhB3
bbsVlLMMaJF92cjHp8Ak3rK3KGID+8zXpzJ8FCVGgWAJRO+3+AjqD8YMJC5Bk4XK
DBZncoMuCzj5uZhs8LUcOC1k4LivTPRWh1/cn/X1NOfJfi8uFDwdPnItO8L+Ie1R
HYHX2RaiCvMz2EkXyYmprsDa8oSKiZ4om97U7XmPVBB0T9SYqVekz5sY3yyGI3hh
/h9IVSxIpHlznmF/S7oZ26Wa3HYvM3+ivhgoqxWy8BamRkBLm5ORKQW4nVlSSKMF
ottKxvMoqJB7StQWkfTP2t9TNc1ubAoIfEwg3VFyQVpp1KfZkbTi/jlSW2uVcAx9
W7blRXx1MWLVeJBSf+zKrBv0O/ZL30TIUrFAiUNXe0kmazWUe15KsTeJMEs50/EF
SlJnZTBXrd/0hA4j16Eo0rMuQSD5GbtxXlMQIf6fk4EH1G2M49hXxaf+VySohxX0
9ikPpGwRvE3pBeReVsNfnSim64zXh5TeM7Y0/mSlnATtLspr/OJmuCGdnwhlzTT/
EMfnwkHpg5mnZ1IDUDHiSB85lQvdY80OtUzRWD9SymEW5F/C2SqdU+jsYjA7qIbM
aeYQhu22Ffo5O0kBJZpjVpIlrnBggOfBjiKy4htevL1WTsZdz9XNcGhlQ0zU4cex
60kOu96/zRejhgT8Er1gbX30Mc4+IQ/pvL/wT43PyVMMWl+pnsVbmjJIx7l9klf6
HyV4TQuUqGVXAYhHKfFXRJTiA4DyrCrwImo7BI+lIqABz55fWMpYQAQZOFkpHqHQ
ZC0tE1Ea4wJ/g+refQ3FAUCWSdhVu4pKeRBIqzHWF0/gFLMH7KtNYjRFsZFhc1aH
vV8qeIeXSo7z38MZutbqdIcuM98Cm7OO+daLXlcroftAE9GJUsmeTqdLFOytJNel
cXTXut+iRIs33WjgRBDpaae0WcZHZDnJUqTrWeU3Pc2Y8TaDro8qgD4aE8GO0Rot
RiRQ5G4QMm/qG+6zRyTkLQe1zaJMBPpdZm40kmvoYs7xRoNPiqLDlmjSJ0lIaoC7
tJLk1YEej4vcFYrJCoH7zGQU+erZak6Tr9XitZf4cJ2tSBDrUnQ6duvkivkEtegY
f/IorcSz1TPfT6qBDOEePmkRw/1QzXeqBcNscYtkYr3DgMHvHmOdGHeipEQ4W1Ti
J5sQ1d7sHakeDCPmtGuyqoAqMLDWC53iVkXAPUhHdJ14ZBe6iPpMmMjwaALb0lWn
eXzPd5j2RohkTf2ShjJkNTJqLgrLUsnnyqQG/y/5E7Oy5DwD88ITlHYik6T3rEfq
2nRwmBLDCPXm3Ia8+7jCMmpGLcr0uG4TEZv8DKC3ftuUNHSk5MY3cEMu1yc37uG9
YEGIabfxo65UY4PIaMkF4pCnHWHpD52UodB+/y0isn5mZrHgwEChCjKxqUusaC2l
GJb+hVY1jLiQ0NzTgN6SYHSPAbkLQGkzEuxNr3eIQNhQ9+CmwgG2ker+q40l6p9H
Ue378TSH1X9EkQCftm8Rq4jEN4euJdBkTjuQ0jWJoOm4aEzc6ghMJrggHzOaWfkA
ZyExBvEb1OIcS58kgKpLbGlDzDroHVvH7OAiREaLs9NVVljcLS4/mhUbj2+ZPPnr
RKK0TAUNaCypoGDCFM8Q5VoZgylar+NOxeCjWsBzrKoDMgX72BolHASbDMxHj4vQ
L70TAjVt6tWJyOMazM7Rk8yhIY1wB/a6bQW53K7533E632nXWMYpkhScc/JGVbR1
br6SJoZgEPwOsO7uxGLzCUaFbNshEZh+AQZ9PD5IGq0kgOfi7zysagbbrjcD6D1a
glzpCDQwqNf3q2kt7PYgsQ5vRUkJ75J6cte0zDVdOPo76aZ6TaXDQkTlrJf4uP3L
YYzSYnCzCvy8iyVS6FC4W3b/rImgjpZ9m3SlrrK7Fp3Jdjp1j49ZMT2LWBUkOwVS
gQXlxz3KMP0akZgELX+c4QnRAbEXpNRTOSOlyiMZApuKzcEKd3ndm3Nempax9GMI
cTGjUgtGCBkzKGKmIz7aMztkvySxlr8d1/go4nwHRG6nWrI+l0zdShgL8hpQ/cqd
8539AsjBWkxl6uf2n+TtYjNAIzhZ43+DBNzarNnLRmqQwqfBGSVW/zeXBKUb1Tv1
jlO+nJCjutFvuphHg/DTyEknseKZ0AV3d2dZSiOJltXy5OYHcXye7OyfrnX48g2P
RLVhzcvG8+MmSQxNftUNW2NfGmb25BmEWvD0TTfcd0evSfonqmBm3fRn4TixZvze
1sWL8+gth84ElhlMopxrtMFvEKMlmy9NSzLWA2QMxnQ9IFly43FatWzsjvuoXqTY
PNDF8S2upjVzVOKrlvfYTU3KAwek5M/EdfUqIii6fAUxkzZ5V50SiYPLyP38YPlU
N4YOvFuth7D1NQ/AnBFSFP7tfSJoOrJTCgihmHLpSZpMw+YbJ/rL79WBd9hJA9b2
x7hk1D4s4lx85HY1X0LJcNZn6SeVymRL9B7t1jjnWls4aAbvyQKhmgArUtvULgEi
4lMKRqcdAyiGZtUZH9W2hDKR8ZUBE5ahaNAQORqLyaz1wvHgDchq0mKkNs1m0sAP
ZK8L4ZZinLefiAzn737Vfw0lbnNwLBgr/mvjg+gresJhJPgi3KhuEPqcWZGzrJVk
+FEpKvJWxsaFsaDOzx0vr80xN/eI9OzepO4VGCieg04begh4CzLn7/3m4ywksR3v
u6zr3iHu0Z21wF3J6axlUDWTtUYOMXC8vUKG+pt+885XMcyuTsuP+0tgtCV0n/s8
PY5Rl8ns+5iRFuJbAgW2pccNa24k0vxZlmPoLqghMxXO+u8N9O774t7siflyL5m2
NCq8lCXthPt6yp+8Pha25S6z86TKOIRufX5S+MPFO/O6rgWaQBdw7YeF+kFvWL78
TE8Tp1AGGht8LoVzQrElwIBsqA+E1FdwebbnnfNdu6lgJWXsuIIm42KabWGvBrvj
SRLvplsfZ3eLUQb2tZ3pnso2VEcSwe727RMqu6+Y8Z4Xw4Ai8mrggSiHON3fy/1X
A20S9iDxzQ6R8rytOwAh7cdHnoONmMcR8Xbuq4ZqqwtcH5UeZqE5t01zZhHzGfqW
xDSPxmyXTM+C6Leqeiwt5s/qEAcqdLCaXeWAeb7UqUugrZYAQUwc2Es2r/1ChdG7
LEPxxHAlezAeWZRvRSACQO22A5S9MOZSYryac7X82RvLkOi9zkNf8eD5cpkCbF1c
3Y/6FTsCP3c2ABfrYMJkzPOnW1UAytlhMNN2+MVSE2mmCVxb1j/+AMHhDpJFR/Wt
3PCCmK/ouaTIl8FCfqZLrAaxlBu2cWCqT6ZHu+kNYfSnwx/NGJ5YwuaLdR44zc30
OvnxwFAoOzGvp1fU/9Epp7k6RcKEvideIMV1G81wxepC5vBsRjeAMReDw4gKgdp+
vc1PyQs/UdrlEbrth14rytuoHq7TwjMp51bJ7SbTtj5Roe66Xltcf06bCw1MkRmN
GvdWwx02rNF2dgzpLBAfRc6yAMDhtsm+RYaNFBVa5PRpWWYYbOrdSQLVBqJlRoDf
ZxnOD2upUMzS5hhSso8GCEmpXBStGi8gvbataOlEgg/RxPWfcoC8jKvUqAZjMgZx
uAmv4/O5PNBXeLSLowE41kjl7g/k4OxJ1zkkOg346H+lNwwRhw/YpQGLLIupwoGu
wW8LHuu7x/nrY6ssfUA3RmYm6QE4cEme7oSP6pLsCfqUBhaVvQ6cofErXPmAY/Cx
aAoyoMhRFSjQEJW0RGTlfb9bdI3BL+YEgeNo7lvG8PmkNsdQ5iDnsmtE3ZB+WJs9
VsWb2uMciBPTb+0V5GiWWOvPzdJCX/flFj/ViKOIA5kkfybp0ff+z+v3acVtn0bM
U7Ru2ir7U3n6bebLude7mpsuyzIornlLf24ETuJMSkFLRJ9AdAjl3sCXq6Pdamai
qJ6cknYUylmdd2cro8bVi7NPkXTmQ2BX1+jr54nAKX2vt5zSgFILsUrD7NYlIN7T
rOX0Y1Ks+m8o/G/fTeHVrJWe18W/j+Okdazdb1xwkmNR/y9DqGk1AV3ha1nEUQ68
EwvbuJt78ClOxrZC+U4dgLBWblzeijU724Z/9DPkwabqs2YP+zZIczxN0ocFM9ap
pSLavBfcMTIGOWw/7OgC/UV0YiitA4dwBqceWYFLxCr0oMNjv25QfP8VeFe3qnvE
v1ChTekIUBjt+wQTiyup+X3I/VOHNbw9m/Y/+ib1GYQImILhJUaYAQsHWg7uqMVj
rjJAcV2+han8QMiJz8TxlBPJIyQBKWjDsukjRJrUWY/ggS4duaC17Y9XdDP7UydE
rriZH+Hc/u/+f2Y5CCzM1cpN3BGaTIjU9TvU9pqkU60Bf3qM7fBq/wQMZSop+Vdh
T1cng+9E819oUb6hOBDRMyQgLrih68OAYYBYDg/eZmn9dKa7o2MvPKifvv/IflSq
GjvUfgXBAPgllTTtKl4tcpARBhNcyRkZggt8eG8wp6EJZJg8CO3ElWdTau6/kzfb
Zb2NfBMt5TC9Be+uDUO2JXUtsEqkVrFgh/yVwDoNidJuqIZLXRMSwiC74nU+SYJx
5vP8NSJ/Zrpqon8PQ4XUgDRPW8wSuR38+GsJypYK4l/qDLJjSx7KDELbRO+vbA7H
GsydHMzdl8xl+URsedv6/hVXfWgQHtP6uRfBdMhawAuuUygXbNGgCsq0Y5tineHT
uc9+kvA5+vM2vd0mJsGoNdtF8KlYQThBeZ+gNDdniVNUbnGWq3yI4KyAuy3yULbl
SqEJ+NRR9GhBtQCDJnde3KFWx2NteDkkb6J9AZsxGIv09YmTTQnGAGm7UiJ+XAX9
6nHW+2z9K6BcoCvUt5qgd4qE4T3ZFIWZnO4WTQS7Terrh7l9Ftw/Sn/BmBfJwSnA
sNzpNui52lXPFsMdVJDKqm90wqOOd2FAjJnS1kDWHhZq0CjrpFbvbddkrNpIv15W
EZkZiazsc7fdIVHZkxo39+8y9zGjO7i6N8E4epuYQn1uAVxdHooq91qZCEy9XaOx
Qxdf3CXvNjWBj7Q0kwP850itsHShnzm04MNqiUgHZUTB1NwPFF/GWg8siZt6+79P
TSjTYQ9lEh2kzXuZjjJKFNMEECVMx2sPmaJNdGOzIeraTJywDOT0LDN3irQxRQTo
f7kI/3jBws++PTZevqOSnJPGVSiMJQGYy9o1dhkvj8/zDg+cBjDWfSjM6QAzbT3B
nj9/gBG2Po3hzsRB2S1vFupMYSCAv3KH+RuJsWWJc2Q1L6kdsaRhLlQxJiuovkZ5
c2Cp+9AQ+EF5mg4mkm5FhiKD++zBh+wbuQ9/t/cSekjofm69wxQxErCAd/uRCUqm
gWIjX1BUpTObka2iMgalxIoRaxsf7DxFX2GECnjAIJDp9ccnhbxiOo1mh51QUsjt
riHgo9iZpBoUibs1lFreEiUdpI4Vd4A2Bz5sln/4LB3YVvwaQhPkbupkTWR3gm2R
MO2Kvo/1jaYwqeg+YdyI8pBXacCkC+AHdCsvX2rnMyncs277+UC4wKxZLoneeDiC
ZL7Tc+BPQTT4o4Tk5yVvKzXguLMIC9E0yunckxNAlXA5BcDT1uZqWrmxk0xPDoXR
t4PQen/QgtFmiTi7SuANuriJLDzuvYbp0zqVuJgeamlOuvTworexU8htZWQmos+z
4wFWIdOPiIviY1Jj8w/VXlPFdHRIFKj9BTmpuGDXUQPO8uhdPKonhYmqBWjWbguU
bxFpubZV1RI3/NHymhBFvXvRVYhdZkLRgofTpYRaxnHMQJFd82/MTDls1k9LEBX5
v96ZlGcW/sXPe3O1YOPB98tey35oVbbGFNpiaNXloMgXB15+kK1E4CPYv2TtvntJ
B9U6r36AbuOVY5oDjldgOyzoJpWB50dUv1EC1tXh/CFkkoQODur8Pn1IHbzdWXyR
yE5CERpra8A1HwQY7juAlrQDAaPtpCBFMsxludbQgdwaIUDK6Os0/MCQn1fsVtUL
8lIykNhRdL625bZv2GM6x87p8FNJLtVIEq+x/CKjzkdPbiwU090X5LEMP6tk7n13
hsU6NS8RpH0oq22DJ5hY9VSX6BI+i7CtVsOi5qJe0ihdwK/75XcKmdA8oBPPS6wm
40KaVUv5rqeauBbZIkM55s/OdOQxU/I0QTf+DBWtndvIKZiQRHhDp7zV/dE0aQcX
dzA2PjoePLuF3acY9oGGuCxb8J2qSBPcNy1kjRNoUFyWbLwo2K9ETqm314TXHCAT
/G42IkhO0Y2xdQ/dyhzrpQlUrHuSEYU5ZwKKjAilkt2iVfw57b+YTfmTXGwgiiot
P6dyBBhtln9k1YlxZ/nV6MG6L6m/ODWri3bVbtMcnyH0lfC/oHydRmqGRez0YeDx
G4wAz/wJ5WJNfjuEkS9C8KUg8M5qkeRwmYIoUa59nJVB6zZv9q5oEHi7Xuf2QlY5
qwffkI9XqsGvq8DB0ehGTfsTJ20nR96AS3tkQHDyi8uY8so5Fqxdx1hyWW/19+3F
HI/y29JqYD8Fe16bFf4kQNOSLt+TrYJ61mKLF8aNeONkb9U573ujcrO8LJgCx82A
o4lPDZYQB6X53we70wQjTW4bLJJ6MWLkJNPCfAtxZAR6adulYXnbRGIWgWO4wWuL
uSqn5hX1VWt+KlINMB6UfQfexR2zq8CZiJqnUy/MKUvRoW8oaYwEePYPRXZAW1hC
sMocqFHnC6scduKfWtwl32OftjoDm81+XbCi0lStJgCojahSF1Jx5EHXJ75dfL2G
p3iJkE+rYw4ZY2Y5m4GGgFir/qGqxxGSCPpQAxzX8TM17RNymIEOVpo+zrlkgwww
aOGyaIB0L3tocvMVMdVoxiK+Q5QCoP3J0R0562bdmJcDRT4huydWh1HJC0bxUDtR
6oa75foQV1tAqmY+AWBedMq9GDCiMBhZwH/9gj1yAkfkRfJ75rmDNtBNefDuNvUg
AfzuCUhj4EmrlWnFifqMkCGnEhJW9TIJrKcNvVwPl02ofLDtujuQftBebaJ7ZSDd
Ul6dNEOzIhYwBk5lEA/cazocx3ENItxm61Ctt9ufpCnapo4O4EiASUnrN7EAvY4H
L6tkLolNFi57ThWP/zZG+W1eRC1Wt55Yp7CZKJW8kmwAZG5VtSRnLNMDETGf/Bql
bz4f7KHxhReABKUxrF4yKawQwIzJrK+eETSfDgSSygczW/EayI0yKl+tyNhcgoFX
hT6Gf2vJNXKannjhGO3oisCISbZgKIWpFkxj2yj+d7ZfpRyW1D7YaYMJfa+IAZTS
FtH7lDxov5NopkL+XL/Q0HqBUERewOt3aw6ByK7/mYFfXyFtJ69UA6igX+WF0Pha
DNZ+nbWSgVu7A3GZ+xQG9riFf4mkqXvRq79mkKgXSzV98IUXmvcFK9kBGoezKhKZ
g1j5VBE9T9gonstzAI+hBr9z0uLg3DQNnL7j61DDy0j2e/XIcJm2BBOzv8fCRtdG
yLaXGNlbk1nmGiJvZMesatPbMX/ATlu1n29/xh9qXrgikzpy7Ndfz5Db5PFfQgXw
p3Ob4HaV7zYwbk7bZikiJSAZfLgGoR5X+Q+KfDyrJ1OjWgwoRhSn4yrTJgwKC2Lf
Pfi7mRkWHvOVo9Jnid2wmjiHMCuXFadN0A2Z/Qxhx87xO84UwxIRiOIVaD1JF9c9
dCsjmG2vR77BkSS/Lqe96rGa15fcgjXLgfRJ6o4VfQiFZBgC+2OOTOpZnv3ipFI6
vq1KLpClBAj9ESoEnu9w9cfhTW49P+35ZtOz8YXJ4Aq1CQH+SttbvEzECbpXPdOI
3EGldP4HxncPYrWu9KInd/j/WhT5Xv9dxUtzlMWuZkKui7ZlAKmWz/8jS8gsSpSi
6jPQqIE7y2lwdV0q7y9ghb5o78pRuAWVOc9eG1FjKOGtc7jCAvuKAhfbPpGt47Oq
2DHKOoL698tGbZaFOrs1jXv34VHYaPRDkVHcpKwXGhAYRK1dIE7ne5/bwWE2lmsm
niKDxmo3r+Sf+YDwbhoTTTz+vEnNl+rPEuCSh6Dup8YRSXaXQmhMh80qpWY/YB19
Vu70ky9qwHD8iJ2iXI7XYrHlOmscD5c+nAcDRl5SszU6169Pd3LrP446AlQl7fNB
yvUsG4+TiT42lbv6QYmA8N5/HyR6bUjkTdMXZFuDu0Z+IYBQ6qUbr6pPUtO7Oc0p
pLYhg4A0rPXJiBlQaoJ+PICCMwXUYsBjQ2P/OExwOr9HVoRXQT4RPZXtZ7hhqyYc
j3gfRefzgWe26ntulIlvcnAfOFNycUYxi0jxRDbdeuAHzMY60PJZZoVEKWe74nWj
BkliMABuiqvDqDZ/p+dyQQ/o6r//sztqlOqSduvFGLDS+7H/XDKPqOMwbvxoG3PN
0ng7OR0c+4uzLcMaG0ere7QnzjRs8Si1lcItqok20OtoBL7EpE2l2BIicHiV5Npa
MO8LcTSApyvjdjqGOQ69dgjfIS346w9O/SAxjh8WmnZ0Rn+ASba/mSXAZRbGHOD/
lvJIKaNTDR+w41GZuKOsNShNvLace3yFGQC4WU2iVkrG7YdsOfHQrdpbzWBY9A5Q
J7vl6wW5DOc8MuqDfKkmNZ/n07rMEg/vCz79NozLPUSRodSKd8i8nWL+uWt45NdH
VmfFcOv2b8lg3VbRLtg0qPnKUd+4BWivInpe169vE0GihDKd2+6eb+bVDqh7mtuK
G6JMUJL39EjK1ExI4LgxZMQ5t7G4Ie2nV5PqiKQ4BomAoAlJ12LnYjvfumBJzflF
s3iINsDe0U2I3vWWrf2zBT0Nn6LDTyXQTatkavi2ADr78pKc58S/V0SzsVZvd/gx
NTDR1WJoatwEGCuMa4PwA423ZNWUdFhUbHyEO+YPBxvBcGKXBso0ntfXw6RWXl3A
30DO97yIZ+0JyH9Av3lrsIHakYNsBxscQGI+BFoS2EuRUlYiPA9w5PV02KP2qnhp
mHX6aklOyJXNkdED7dxnzPNsmPIIO8F9h7Jj2mT+iTmmBQwmaq44NoKOPcWpzSqz
EbpjnyUmFwmxHl1rVHjWhJ1OWcV6u/Gbv1rOl31LGUqcMtqjX+14ryMKpbTriyMe
fXXjZvZ+zO5Ti0MZWPsU9Mmg/F05jSgDctJr7iIMvPBgebN0cf6Xru8v9Y8mP0zl
VPs3pXsLtJ86p9zFOIdz9hk0WFqQhQ68wSH/OGrELUCKH/XPqwivAgYFXrYapGty
cyPUF4qqUPSiOpLeGBhkbcAldKTnSLWbCeuIdiaur4puMeDFQPBbG25op5XLvI+u
vbwrCkT/UrMUp7w1B0wfJGUkotEgjjAEjT9QTZElJom8CUbMfVMNyDBGTyR/pTMF
9KRHcM8fF2C98EyJK63tcyZXfjEM3HeFgvPp79oixENAp7zaRx9fsDQSzLzYTwCx
1aBGAyXX+cmf8i/Tlic1TiI2ZbZTzOyWdptcCyJ4fgaIaChnC+uAokCTIAmCJgNE
IMdviai17wnkWxEKqwyNrQC4ih/jpiOfjhEmDqKFdOl7dRHmPBgGFK+L9juQX2K/
lEnOM3IUmFlhk8fhxuk7fXhPssK2mcM98oN1k4xbqbTzlHMJCXkO9B8dIbg6PVey
OsMrjKrExSA14pd6/6vy/SwALfN02J0xuGpeapIe3tOtP7pof16N8uAEB3VnBkye
W2nCJsS4Iw7eB9G5hAnKLbuJ6YKvGbveg8dX/L0ywKD4HmGDrQ3ixxzMYSlizTN/
iMrL9w+HOrxS0QPEr8IDAZpS5q10g+yZRjRePazk2vJ6Y9yYRcPNSwpb0I2LleWI
qYphV2Kb9IgLJClt7zC5pniuQ2OTSHVYwDztSRQmfweTLnG91uavWBa71SauSZpv
Y37B6teVjwZ7M7bVJEXPN3XErYB907S0bPPAO4amen6cVZS8L8dpol7+Hy5D3TJA
lzmpMS3DhfJ0JORDZEVJJPr6v1lputMNwk6ajHUIVxL4JMplO7fXq0RExLxH9Kgp
RzWcBBV63X813lVPNNkPWtkqeWAZ7F03RyJHyKs2Fe7aoJeBnXzB358FeuPo6w2e
B+V3pZP1taxTh2VewwYMxN8QFZqm2K4ZBv7YBQD+BsuDqSdRC2sDZpojm5/iQ2tq
cfvu5YNu9lBBYPKnq/23luXpqneIQl5iJ6fU1FuxA1qGmzb30/2RmO2LW4QWfBu3
vapQ254wBcXucsPjjkw10zoiqWPZRxe3qbkQhB2x9QJJxcaINaR4KvVUaM92rIhw
QktdutiD3EC6m0+vWgvrP1E/3/UqaJ4hx1P9269Z/6tUZoIFtRzfPFRXkgSam64H
rCwNhuhgQN4xchwS3/ZboDrbD4cX0sSoKqvZJyLN2X0vqT5o7ugL0KkO6uLGxJwX
gznhIypp2dNTbJXqLm8bT30NFklj5KjE6JS1kSBXrJtVcEOFNZLUr52MGPMDVRKn
mgc2Z1wMxmbOKXjVmTGq5vYgs4TkeR26N6c4TCelS/P7zFR2naaolA+IUB82V08c
d/Y9xlyFv5j2t1Fr5hMrE8AtZuq9h/3XEvyUWC7B3XQCSZlFH5VSvfdxEAKky2mX
5cVOuhscuEVFhNQ8Pd0q/niOGpuI7xBZhycO9NpeBDAkpFkw2ioLYe/492D6JOOl
mAlEljjQHdZ46CUSv7pu8fpUN6PtWRPHbjssji+AwHCKuS7g1itM1PfpRj3vkKca
pmVW9eICPjxFJAG2HkBDDzEnpYlupixhQNqP9yqconYJ1g/6EaOQrc+CS7jGLa03
2SxBdlZYXUnzSFHd9WQ0Hlj+1lnlcYgX+NlyHunlokmTVlqx4ubq6+GvYPe9O2b6
lpcip07PEJ4/rnFKMV7xBz0MrCO2f+j700aegJwea9PVE46oNpSPvHTt00iewi2J
qPG2nRGoR6Bcd/A3u6q6+hIlfd5rA58QUGkie3Xc4DFv+09IxwFuDfXVJGCuB9C7
xQUM5TiC7Pt4X7jqu0lZ2mRyJS6WEgFDPtWwSuA2WGVxe6l80XZrLEC/sUq9OIXQ
OeMOJ5scktavMrh91qy2f7v+RpFAhEY2echAvNaEH0T0kP/0vmsY8Yx4BCKp+kxZ
xLp88inhvyaLy9oAroeqxvAYhXLqWFoWO6RUGWLhx5999Hst3z+etibOub0fEPg9
cI8QP0cf/DAIO0OoheDQ2+xY06nWMHnh/pqvt4QhXAnFV/ySKJ+7r6BBy9D9npu/
3F7R0JsSfJFaUKVyb2UnEzxZ+L+u8ZRylymtrgUkTFWr5oftoT06HCf9nlAyaXHZ
SnvlCMmAl6idptjesxCj/vklipAd0mAo3RO3o8LMjPrYjqvQVIaXCxl6kEGr43SZ
4CuP0AOB/HmAaE9kkx63obPZS3ArV0ROaaTqUe0fV4x5l8TkJCWAt9WlijsE1rKG
pFz1QEfvw7yJxjvexCISCOT/wRhdKt6r+Jp2CivO6DH6uKkncos0uLL1Rf7RD/nZ
uCphJoBzRnkj6wt7Latyfz3XymGb+L72xOvKdSN9TPtkew9yTCOfxrzJgaTE69OE
wwKUW3YpCHX3/KsYjHhf4rYeLphgr3eOs7yHJwtSPG8oVRCsy/rBtm8u2K777wlp
dEMxJDPTmIHK3g5BwPGsnbMZvtksCKTNFXATfRNMFI/T/htFVnQBX7hFeSm3JcRi
dZQkD+emnStlMfGu5V4hZ3dJGCrsVQySXM4HbiXTjRYqe1IdovlRk7Np6/0Riz3A
QzXkqehjpxutq7R6hAiNPrO9o0AZzpCHj524hhL0NAQRiyFP1w0DRnnIubgWJngB
A5+YosOQhqVLKgzEdmh6dGn84cniO00i6YrtQC0ZD4hmR/xfmg8ZnZ+qmic/gsqf
Gnq2sFyodDmnxLWEmBXwZXbrwxikzd4L2a1f8+dXFabCImeOQZQ8vnOcguCN0RII
bWjKMS5NY+2Vez+VCTiD7PLNLvjWx7TKuef/ZadqVd17PtBJL8hcPbKMmPJsqmJN
TCptsC25JGkKgi+Wf2yDx8gjywTCefXMxg8ATABR10xhnTihhvAMKqHAez2Y37Oe
s3fnItUu6PT8pJwuXBg1vwvYTi8d2ThAI1bnFnfwpqTSwYu05fyJdOnMnlRDRzYU
CWA2zEKUZWWpxVt0Itbv1+CYkaLUGUfxTavIHxl6lJ2Ia2uCHEKBjVJGHI8UssIN
PJLzxKO388RTJltz8vekEa7469y7dfleVzY4W/hIjcRvEM+QZzXGgqImBfB9BsDW
wla7a7sh6nqBONEybBbu4/tVLLBundOZA0M6lAlNx0g3hDqnA1AVWHaB1yQOC8+4
2BfBbsO8bihrCiVzRYFEKMLs8oFrSybjbuh8aJfrucZylo9Epl9tURFDxclqLY0n
ni+1glMUgbArlPPZ7aijokPUDGPpYLKZnbxPe81WZeH1h8FVrZgZ8lFgNnnRr0jv
Z4yditYC2P9/V1LuatOnjUOuS806C3Jr0gL2znQRMsK9veZFj34Gpit7fFzeuYf5
J2zuyscZM1qbHoeXegzVk0HAGzIEI36SJLBXsnJQUuLDltGcxd8BhCg29D+s1Hhm
TJbuhCWMUWhmMFm+0EL9a4wrov3KgWvl46QHY4VXCqj+l35ocyuDBHeSsQVw2odO
F3EIJBhRyhcag6dfO+rvapgGDNmx/ank6aO2TgER+97KM5hKi+HXQKCUoh5zH0ch
y7xN9h/O5mcSdFLCJtS1Oriw/VCxCbR7O4e/ht4suYC83ekzbhzsTG4t+kZR+tHx
Sxlc5K3CD1IJyKNL8JBaGR9VQZIada3YE55ntDGYZ/43Atl+nxxOfPR7cszY6LMj
xs5T5+dp7COknot+MtY/W/FCiStaa2lQjFhf+1GEvP+l6pLnO6hV7qjXwPeHMhmJ
8BBsuv2Cn2x0s2zHnG++/JD8VkCLCmSd3fM0nZqyQWCEWEMyuFyxlOA5cKLUHUca
QwlNYeI99p+6wVlbkWOIRFy/nKOsBwyHpRgdWne7uwxuXXirT8rhSm6th2IjTZg8
z21HFdVGuJKkoCSis3S6gJqEVnFvqLFR0iiEGDMNiAQoQLFhTH7Nvpvc1bJfbkkJ
pNOixm8AlI87yD9/tQ1TOpe3NO+vPXCLKGVpauLFuQLt5Nx+WVOjp+KY3w7DeUwc
7Xz/vyVGPxCwOvm+++m+w7bwV16iv2W1gD9nuCSK/xQGoL/hll4GwrBSDwBOSlPx
K5fRKObtP9guDQaCAv+MHgDAzZzc1AygNHzSLIkvOrB/BgOv43FYaAp2B/+aKfkX
1sX1CLR6Ah1S2HK4/VU1yvHoRJHLp9y7VC7I09CZ/ScxCpQsH5f+Owc4SY+vYLhs
w+WVWkNPYY9JKP3eQDWE8jVXndH8w+5wCugw0hCssQbbtnBQ3PX3KmsmGuXrE3AW
LSb7wLKZQ4sNru9UoFydnBt3iLeGuIAQ/gFe2CHnk2I21thUSZ7N5Qm5Y/iUWTEA
dsH7V2ou+2ufxmuDRB9O3GpgjXixYAB9xJ3l5o1glKk=
`protect END_PROTECTED
