`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zx5ndFQb/+b5LNPMC/8QCvh7ehOy+5woOhHsM8MkesM+mH/hPiCZWmEWOvVyW3kO
bSlVuYmPWIIHkCaYb8u55AEQQ9A1isRYuB3QUayoQ+K/ovDidqmxh464xy53lG86
hZ+xb2+6ONkuyj7Fj9L33RWNQ+5Bb9+A4ltNyTxLsg7c74WB70eZkSL/8MNIviZ6
OfTI7CSIm6zT33+ukPPXA4BPJlRA4KW9NgyW2L6oB6i5RhjxoFFBHBb89hvejY/7
fbGSQCnVbCNvlILTf2/0x5ozBfxeCxx6Ew2pPQrdWlNpoQStCbuPFFFQ9MXWXxm1
YPK228E9rVFU6uwjPc1dPYJtOuchmLG4kPysLjwWTTFB5f58XIkft93a2+pDDN0Q
Q/cngEDZuzQHcBVuf0HqXQPIZEscdo8x+2zLIJAMM1k2Np5PJfe55Qe/TnY8Fl03
5/DSBzApcNN+hg6UV9EFgmQndBF+wKiGjCK9QaJGu8kMLlwLl1Lw938Nz1sr07OS
cWh+QV6MqAIYH4uBlDsM7A==
`protect END_PROTECTED
