`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61dghu7VxnXsIAnFeWQyWp4RIDdP1QgYj8Ijca/m+/uB9xh4ZcUn3PjHu+/a+Te8
EkG+gD/grvziUGbN8cG3wKdG+Y2Yq41k1gz7EW37uNY1udI2A3MnYVcGo4kVRBJJ
LjSNU77ApAtg7qHVksJaaCk1f1+Lsf4+h2QOLYBQa15zVbtLFCpbh53lttitqeDx
s3dnS9E3wLHXT4vSsjIXtrCT63zehq9v/Zg6EJolh9EBOznoKXV9auFrDjcsVk7t
AmwKJONJNdOphtb8bfLzygrXojubory1rZKT9m1u+oQw4wjlxrHUZZsqh/ydwRSs
/BdnUvl9FAYWImDK+rWfx3H8ujYx/2JJk34ovyp9Fy2gUwoesxTD4Bw10XfLwAUM
lJqnOKHpLWsPvHlk5faWtzKSuxIZIZwJuxouQhAdPksI74iR7M8RJP23GXFUqwya
958wcz/JtvZMufxui/df7EOqxjvvzJU8O6YTrwXSXrRQ6aES3LH5VUwa1LYFBomX
hVIMRWnCFnnSy6vPW9uFsFBW1jQXiKXCuNylAdU34Db6JVWjoYCd6QD8DtDj/43+
Eb0veRRX/hBGqqDIqLalkpETFhln08ZprA8JMZUm5vNwzG1OrV8521dPUlOdMbEL
2WfOabpjPq2pAkXxWDFMiwaa1KMwS4QtWwAjwXTNnnlafqSAd1sbUKOAaDuqdf/C
qKabSTqn2On3YRxMjrE2p4iZFr+QdEla0YDiR8cT9EKoFnRP7uFqb+ZN+k7Z1R3h
`protect END_PROTECTED
