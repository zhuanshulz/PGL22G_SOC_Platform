`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ewu3qZ4VHZzXmZQkPPQQjlY/TEpZba30pmMfMrc5Bud4skd8da6DvuRzKUwjkxL
GShBoUM44sRfe0lYAfJgyBIvX2/qrfJJP10B540JirY3U5gtL34GmH+AEPOceJRV
aex3x5Ze82krCdmAmoyGb66ZStPt3hU2EdYZSOuwXLun9+zaL4RIWphRG2tia0Tw
7vb/gGmEmv0p8xeKQmDR7Llz0p1JocZPjcaPjcgahkao7y4cJwdXdlPMxs1BM7Du
tXsITsiT6say3sxGpSKCdZmoqGt2Cuh4z7q8Ly0sRWtJYtGbSIEB+zrxnbrlRZH/
hnvMe7ggZ1BpCtv7Ixyzna9pawVYh2J/2zaxK200Ty7nUux6TEk4d4NRDNyR+5/i
zRV4R2FSWIaB4XioceU+8oi51OPyEOsPwj6eR6NU7rHN7+VgEoI5ovz6wnGHMwo0
FawqlGHXNgRfamqj1n+Ruw7wUcD5fq+FTr0JWsoJO45cBI4hffj1CAjEkZhCuPF/
W+CIUm3/zhsnfDXOq2GEVjiy7HkeScoArk9hSCbPcL4z/mr9fN8cscFhjPEZ56gT
svszolXb4SaAOtFO35ryYx489p6hiq6J40XPkrQZGpDG9tk5e8JU2cvNa01XQemf
tw5iR5CdiVhM8/nzo0uLlkgoLgDtf5Tj7OTj9k111nyHeZ1nZXP6/0Gwd1ZwKVQN
td2ZIi0EloACRTp2pvqe+gTeQHVh5SA68I7ecr3lDaLE6x0rBVHu7yUOfhLcTJa3
DWep5QEsqbJ4oqdFYJXR2zR1osI6Bz2GMdMf1KWvsmXWAJZTKIOmOFowDZsMioAr
UlVliO9uhjhUSPcNivJnlZ7SSRJop2Dl9iK0hfB9xZRpHblNazLq6XKGibMgOTXw
Ey+QeudKlAAVecd7zZi0AUh7Beq710wrQl7P+k7cN0AbEg0HE4+imC5jCfGJgWRW
rSYWo2mCApGpLVnJ0o64zD5Fs+2LZnsl2Y9HAcGM6U7CaWuffRsa+7Wh3iwLaHH0
HcjEF1LQex+9XSd+31TXtvJOZHOJEgYy9ibHWb6OohQNU+VK6+itZVbkKA5ovjkX
stCCNei/i+g4Ibqv4wLgVDOSfkOzDT/i4I0QMJVC/0nuY+lOl2qgT3XH1ytJUrpF
qeE2K8StqepwhgOE1yklavIKaDPZaSsdbuJbF7PkpfXQ/FEe1b0YRmxowLmjLghf
iM2CrvHQhpj4UTktssxS2G756nf9bpqSlE4BnjeJ/+w5DqFDdcJZqdJXibNuLx2t
WR3aFtNFz8w1oSm7wM2DM9V+Bq4mhONk7L9aHsQRSq8AM3OtpSaXoT0493DgfB2n
d+08iMTQfHondid9F0tiWq10T/jx9wu4MEITA9sv/E+rKG6KXrX9ui29KECio/Px
te0lMAGcmPXFheqjVmu3zgOGs/7xWMrgGe8FtCTEjbgVUcLif2jmKxrSe7omL/I2
OCOnujGzcingTzCEDDU9zHrhHfFTEDNrKzp9iR5GB0U6eIn34OUwWXIewR1TnBht
zKhsJ6iK/N4znx35+Ntzt3k6Dw3Ke4W01BOiK8B2xhpaTQoCAhojTWlRfahSQsZN
wkQWR5LPnFXgwH8BSiPPWqiYOkCdS87atN2XccBthIpRylOynjIm3ueKKYaqN73B
o99VhPgh0vIsDcPUCNhyKkUkEYM17hq+SjXC2HI4dolHtStBaROqe9M2E/a0WdBu
3M+8cmI2JEaO0ZHjOZcrk8avgJS6HEjP47ru1db02fNL1K46agTRTzp4nWdiIooU
xVlpfdnsbqaWekyVBpKpv0Cr/hkr7AmFraHfGfzXEbbmFH5EjGNdYrpuRcq9+Wgn
EHKo7Y/PckS2zQ63vEF3YWECm4X1c5tkNq6G3q+auY+I/ngH6O13B9OVHQAEbwql
pVx/8CgY69SMMbE4YnaBP6HxfwxXBhkdnHkmla7KAe3QP5gDpEpjs+OXY5WF8tyY
aFgsaKFCy4Ihn7bZjASE6Jhq1kQ1xO8ZGqO9dWWWUhgElQpujwgfxi9iZBjG6ej/
If7p9TVB5wmrU1n1IiNVvwia2+Ne6iv1kjjYrjPjglrlmjji/NQTPWu2fJtl8oJD
gjD/wE48QwfAfOyHG/s5TSpancc1AquSeSzYceE3uFwrCa8wxL4rrWFaHi10bi+T
KksfhX3NQxnZD4o2fJNDgSvRB7804H+CrHzHY1AXYH5m2TAbP/yeBmrd7TvviPNG
P3vcZMlZMgLghb05hfnx+CM81IJ4AdHr2QkFxJiInxX7Kuu+qit1uEVRhB459sPW
4+XX/A10hB5GwVd7RANo08P1sbtDDNkwQwWWuuTTp9DqcEgU7cJIyJMobzYMmrwj
lw47O0zT26u1GWgtax1wEyTNndi1blMLTh48N3tWq50K4+Fnfy0waxDWA2zDu5f7
8Y3MDNvHJPJPrYgY358pTB+kmJPpDBl+2JvRaEtufQqnqFvI0H0ng1QsT0jRzVTu
2CsWHNSNNqZeHbwcrsomBN4M2OpV4mKTPcNOPN0z/Yel7ZdDZi9a7a+CBN25AmTn
ER7PSSyFSCIXttlIio1sYRtEooo3GIUGqH9CHq7uY03kM2fR5BUUmGm4Kx6HMSeg
Sk4wifhVBU/xTUHcoBsoBHXxEZ+Y2tVabTYUf2bvEDBsTSAioq3+Oq9MHkfMfFUU
V5e0A5tTCWXeM6m8YOqmonh4vAPETYkopL8oWNFTS80eC4iSz25h047k7dDqfxnj
VMuq+VfBjWKrBCFEMZxHvlyvQBHQ7hVmqJQjiqxyxjiAp80WLC5uwNL5Q5+tEj5J
XRrXOXdEn2IpOyCYYA6ifkYNYvrlZ2w9mI0eESJNvDeBhe2aTUGO8sp0+04Ho1+D
UMA+0Sqf128ZIs1cJuL9DQfC5wAo8tuiqWDRFZwXkQVoPQjrOYJD62qvPXMSKgwK
ah0AMllH8D79lV9T+d9hRPv9AGclvFXsPy0widNvw8hwAb+l2GoTXmyS0ijjO8lq
3I+/8YVn6GB0eOJILIuv0jVCP2o5K4H2PwG+8LLhY+cu/bE8GvA3nCCImpQHUhi4
oJUq3Q+i10/KgkoCuXoJpnLdC9XkvlzTrUKVLhKrrsD9hAC2Ou+LVsgi8HT6zb3V
T9icchiQrW/DcJCZebpkvTqVzVHA6/t8axqKtxksfHPUXEgqiXFsJ1e0EJY9FIsL
zVd/OxqZ7rJiZtcmdxSdhQbOtIibvI270uGpX9jam0t19NrFt/httS0okl0alJ18
wL0pdINp2h1dtFgUoonZ4l8JJuLXD+SbDcMLsHEzDmsiMVtTy2ayCUfxe+KrrzR5
6W155lnImurHSypqttER6zlK+LbAZRjekhGjamgQK+UlKKJ8r/UddfhMGihIKuqe
/yQHUlSCxKAswc9FLdDc/g1NHeFKKsUdA+vaXJ/Upl9z/Ach+5bqb07BjmQJ0Alh
u5sFe2P+bmeGnLpULq45+ypUz0lsZEf6SWzWRV0H5K0KFfzBVUbHqITyBgT7bHR9
PQAhKkQyK0q57wV7gPNnvoO4nCLTkBClbhLHWl2uVK2y0kzs4aYl8HoWKKAAYSJm
9DeX2xyVmJGlJ2reA+1vSOr/t+/ye0NLAIsVE8evnfEcbS1QuB3dCc5kg2xf+zb4
BSZRaG5d1VpwXDElScFfPmeloKT5ohdyyR1EU3lAnDwqupT7n8HUPv90z88lhiSF
P0uDjlfUnLxPLt8VksiocSA5YR5d02vxf13U1oMIh/sVJDanUSpUsgeGmmRCi+YE
iCuGZQEBAlmd/Nbob6f0eE/iRh7VnEoy+L5wDLwnVKAX1ZIybjOVfTOY/KifvRJB
Qfz/35UDTNOxNFQmixUbFffyLJCiwcFat2LgJrIx4ZDasVap+YuLthRwPmE9sHWm
Rp7Wh0KSeq2+iv3yQQuqhTdy9L3xksute8RqkpFYKYNj2bid6SrkLFCUxXDBYyCE
CLNf99qaq/nV9QU8sBMW6rfAbCSS1o5KuGId10tWZnUka/Etq/hhUyDAtd429LWb
kMR6OyTpNKZ1eMEiBTxxbh2VJTR7LMorXNJh3xBzaoYztWtJ1sVmxuvJGJtMbjPm
iKN265CLu2cG6aVd3EvCDIQQNG7l/Yq7eE2dEmvZKZzq0mrRDjhwVoG45oi/z1vY
ryBM+0V1GbVgmlO+IqBjp90N2BXH28PZqNSM90x8hfRcFV+myEM7LcHww8TOq7+7
gB8W7MMLi4lYwzkmMbwgO8jRMuw3NOZQzUzRP51V3tohwkFlPlNc2ew3pjwBR8uf
kaPS+HPv3Jp7rVwD5AXyigVz21m9616+T1yUQwbygiMuyG7qknCjuIj9LXjOtugd
z32qrSze/dG8tPRKJXWSc+U//J27Hbatp6dVoa3XZ14lqvLDqto6OyRLEPVE+dlj
qTk/eV3rLx7bMcOol35p/P9U4j8mk1gyVZlddKx/TZLX9walsUzjwgqfHbQpzi7S
0iDEnOftdUYpzsQh8DCyUcZ4VUPfjYgwo4qiOHjHse+A8EA/0nNNEtQs9c9vHoqC
3MpDWghs1lWVmhTpAxUYRhhp8e2YphwL1aRGQUKvYZ720DhOp+ilKF1NF9h4FUWV
6tzmz/fKlu20Hy1gpnERApso5R4GPmcYYWmOLem0YZ0ADbro68DUsoyQHKjzDi5v
IF/BUmtdz62Mhw3rXkzsNqBO2eAoWK0v7unDwSFcbw4WISiAw2io0SZTLnCRjCRp
o+rfcav67hhCW2371AibhXegFL8po+kz8sEGR2G28fP32UU8vJ6FDpjJBZecIDmZ
ChXacEyOmALk5G8XuFzbJZaCcUlD5/gc1+p3MkSCNIxFFZCTe+Hc+xkmDNqmjDwy
Y60BLvA0s2/3Y7fA+Nkls0ZIUnpqVy2HJRCcveQH9O4W7hMuVTJwendcmbUu0qOz
Kl4xTZoJs4VvijZW4Ow0sA/snMwwdNku4XfsAaqZnkpzZ49DcOrqCp8y1t5J6Eku
32YxBLqT0N/ELxuJgCsYj+VJKKBiI31D5bWeBObyiIX7Vs0eWSEgS1Gtz+c1TaJP
XkJFWnWtHWdI7cip1NngaBCNM7d7nuO4mGvfrGx0kPdyW42g3yYF5Mkos1N4/F46
z3BdNoOFS60C/AN0vlveJ8/0mVUkwlNLY+7y4n2kIVQXZ52NNkoo06Kpkwsb+pPH
jqaWqw64r8hLhNROJD3CTYpNxpDU6y0y9s6VTU5Jn9dF0oSv61q5SRO3j50zdDtb
2uoPvSe+gElZfDUMrS99ycdQv9rBoND3lShgGk+NHvZgAZ6JxDSKEtFPN0a5wvu1
H5hskrkf0f4yG2HqSjBsaqpqw3zDbUMDkH+VwnyO4O0/L4cRXPZVko04TgIjMmFh
roHTUzen9Ei+2c51nx5m4BoJ3k2BGAMinNsKzM5QZBBrf9CjQ4YYE/jLeVx3WH2A
AVH0UblZPrr/NyavA/rYny4kUH5KEtiv6zSGiDZ9FruE/6aEE9qjnhIPB4D9OFrb
b7z4o+J+ZqZVu9PVehVbcpFUscvfzVNc/8gsbp9kP19sSw6AfQzHGVRtvTaQViqp
jNAz8Hqnwi1PAGttrtT2lZSGNYKFPo/zcmGNQbcZQ1J78dOPp3FUSJPFlRNJDSJu
Un7p8Zv6mpAKuH2VbEyHc9XoaH/9wR3Sd6+YD+nZ9xm/40CKTI/EFIU4nCj09rg+
DRBb/xKGickyip8L2kVB2ZRa4urMSIQYvKIMGyKPo8DwHSXMkX3+dgBf1bz1695l
3OsjoVVrZUvcP9OMFehEow==
`protect END_PROTECTED
