`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yhRbUGtnwRvp6bXf2KDBAzSDswehC0sJBBuKpG+JgY1UNU66NiJ2GST9IEK6uKs9
5qetR/jlyNq6achc0V4rUHXiDca/2Zm1HzSR7vrXCdeWHWNJB0OtMzmjLB16/OK2
GFQNBNFRlnvacAQOg2lST4SJQKbtFgbRn7nsXAo+oXJY8rnXiAgRLCbJn7qLZncE
TOKCDBE7VfCV7f2r/SxYZzC12Ud9kk73M4GCs6RF3N8NkUNgGXqdnZJbcWxFDri3
heYptz5d1iwM0RpcudNmrpke8apHNZHPbAmaQKPRMjFjJppec5PJTbeuaPdmOgfi
ZpNkV1qQEzgu4lkh3UvMoLCHwMAxl/rK2fhCMtYb5ci4PZw/zPREip//3TL2eKCM
7yc5iV7KXaZrOLoUGntBLMCCvWj0u9jw8f0z7Nzu3dBZ2H9LF3VpWLEhdhy44rIJ
tLUslzkk6Ayuu2obR7tU+8OlWy1CBZ54L8vVlpb7PyMkqQJNEULf72920DCBMfv7
BPLLTGAO2a9/q0KXSktJdRNleFgPbMRykw71e1bLky4+XR4Uo6Qa35mjPNYXY0lD
jy60G6BI0HwV2DP6kytTDFUgyJRy/NESA+/6TwHBgnyyE220hcYRkOHnCI+QjBgl
//SGeYizMi7pTS1EnVJfVxLU69e6gkPowVQ9p81Zwo9jmEdAf8207CC9jEbgMl8b
SSP5Nyo1LRw0BFyhYE/k4inasI2NyeCqYA6XQ902O4lNiLpHVvbhdVDy2rkic7Jj
qcY1JZV8xOt5a9u7JvF4a+9wy24AXllAUM8cZVxLojmu7Px/vzmdKRx/qwr0lJBq
aYbluTxZWwNJN6DCgcsVDBYvIgmXCkU7nZdenHa/mek=
`protect END_PROTECTED
