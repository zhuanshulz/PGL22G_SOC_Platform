`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gRADP6D98JJbd0xcE2c7jvxJAt1gMEuvy10rJVImsSDzftjMIB68EEmPfLWX6ue
ko1l/4ptNZY8rSI/Tn+jo+KJKnaSBsXLbNjZAVRBdTBo6NMZJIBKCjbCEMDUM2JH
tENF36XTqqdWTFXPUTK7MAzLllhEDJsYRxSZnTOmI31NCANfPRncNVOg6RsasOWL
iL1Jwv1kp4cVArQaHH5nNga4gPkW0WxLQBp3RLELT4bXHxRSR8kGig3YGKdw8vwI
60rXdBVTDgZST2M3kneZgj0+KFuHU/1fiRJ9ZKffe83SZ/cHnUF8g+NinFK7pQbT
W+O8GHYVliY97GsV6/D8VDk1XivR2Qz4fO0ofmfUoloOagcAa8EKDffS3JjHpW47
qijt4/O3BNj9tLxSDjGbCGk5Eox4oL5tIzynxDKXH+byrPKKDVvQKt3TuHSAjub8
VePuBuzkoba0UawU7sUSGtyGv0YI9a2IoidRDwwK/c0r86SzNOvX0+xfYX2biszr
oilYzhsc2HfeMgzaxsGzlQ==
`protect END_PROTECTED
