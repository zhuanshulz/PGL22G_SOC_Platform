`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
serC9uOtF1FzJo96n5zPCWGneJ9z96qJbaS1t0vuMYTMDcCIotQoZ91Qp899gILE
wGqUbPP5czThZgcLvwbshFTWHO7bDxrt6/eyH1o1w6iIV/CgyyydGbI53qTvvPZo
JqNkm/3egL/Kg5SnEAiLC6nppfOea5V5SGx8p4TeicD6c6NECydKiyTQv6E9vYpy
o7xG4yNeROwL5yqaHCe9Bw4z8YTdE1FcqyabbUjSS/JLR8ptOk02KphiO2EdRoW5
m3dkkKcD3LY96EDQdEvu77K9lmihO62c3MFCFHBjmYitkQ/nyMKn8K+CbBlU1Mf5
BfgLfq9c+cmiFm99D7i1pUhh4ojJKN+Dj1IUsYEH7lz6UNlmCeZ+zmZN5HVBi4o3
ugJ76jaPOwSVFYypSpuFdT4w1VbKHLZQeVT8MugGfyotuRzalaCsGzcRyI74/3vZ
NMzipEp5jxgaZmRaazO7chlkt7Um8oUAthP567YpRZt3P7VJoEvBz2ATzZQ7Ya5d
ytvDNDZB169bj7m01dEfuPJIG4RFXCWqryyBRwUcvz4+ZvL4yDHb47HifMLHvesu
gR5OrsIiUztH7GPqd5B++hzqJKMpqbAyzCCQfYvTqDqUBG3EczVKSspNqGQvlzH+
DXL+O3IBN/3Wl33J3lcK02ve5FRYUkPKyxMZGDz2h63mqNqnqMklQc/Ne36Gi2cM
9fG5J/wLTRgzvrlWU/DPFWv2AU5ApzypVVjdYjIgJ7CIhhBTsHpQwDuyVWh+YnhP
2VKEPchVs/ZNcLGzyvhjf/FW9McfSoYgo64G620yvAQk/rOM8wOlMnirEL+hF9iY
pxgRLm2CWkoMFeFU1a72wMTX2291HrS50/c0qRPivq8kfEEkFMY9SHNMM5gKf3hW
++6VgSUYEEg6b6kj44hDbwt+vy+KKONyY8UJCFSAtUv+IqwvDCuzX4Sw9pOnPiad
i6Ek1T7dWr+YFC7Uw8yzk4v3OjUw4YusTQxi4JSK6MuR+6F5iZu4r1WuYo/i95Mb
LWz7RkwPRaEoRkrpNLXduyeFUg6Xc9L+aaAjCSeTbKTaNc+2ITSmaU2Hb9E2sT47
xG5BH+rYpN78lQW3UZQzkW6uJ+Ksdi9Z+l6UrjkHznbnIPJnwvCdXxsmz325sCys
enzXuw6E52CA/ZOV9mGA89yWpwaS5rd/M0g+uUqfd2Bgm83vtuXAU66mGjM85hhn
/H1Kca5fzxjj0PtIx6ErclPMIw96rYnfj+dVVkzuTGdJs46ZHvDraP2h0kT1KvHt
L4Wvfk8NL1PkaYYBCNamLeDNwenRUhuNKUNH0h5OVAAVp96XxHtbXJistLViPS5Y
7fk2YDQjjA31RAbbRvcAabtlI6p803gqqSTvdSDa7GGSRthtzuZBSiAabHMXDb2z
kL/FKBmJDyFkhQsCGFUFddTffpODYubBWj9VNVtfojYUVASjXe/tkvMLfxE5hoEx
NiJE8hqBHRAeR+1guGHynDeg2jPpT0Jg5lGEGdV86b3FLV8QRhy5QYh9YPGNBp4+
U1AGniiJF3+i1HV/DjIuopG8NnZJCDC5m3Sh9lyog6JDiax4MoDOlGYxke4veqeq
0wT4DBgydclGeUBOATm5BeR2b/jyJC8mtxTqpjXN9lQt6ys4gXBf3sDVMUFAp+Bz
p4u/6ugRNBMLniocsxZ67FJbApDUsWHQapYCKOWrKYQnBGUWVKseowbXNPd4jCH5
bFj996wAuYNNw5gRhKRbcWpLFTqWMyPAOaWk1PWujY92yz0U72PYVMA7zkj0RCoE
OeNEam/9n/bSTFhkNzRdD/aZY5r2wgHL7WnomreYYrax/f4JkNR0ITERfEnnpF9o
TWcmUZWplHwCPfCaa6XKQw0TZo+amkh9VTfyo4CBWp1VAllWIIQGIiw7ucS8V1hH
tJP71otakpi07+htBDQ/xyIojNLNE+Sku/aBwqWGliPj2KDoKj8WfvIsroKMpNdo
8RlQJbgH/Mgr6ro6mkdxWGQxY8LCg5ciHh7PcCNuxHrvFVov+B+gZ5WD288fHsZV
osmWlYqBMBuXQr01iyHm3YXaWAshuk2MQFYaom2SXkQKtSKtvNMQ8iM9ssRr8hCE
eLy8ozvHL852YnF+n0Ud4rY6GCw6P+I+b2NG2hpZKFe4Jdsvy87xZv0/U5qJkgZS
nbKRAs5j0ezwCU97+v7wBM6ZFCFTbrI7+VJcu4Ago0we8RmCp52xMf3Ygm76AAp4
7dSCcN84qxKMvVIBxb9XNZwTUEsi1Q72MFP7OOeSWXySNbHTMSsSuY9njrQCpt3l
r50UxMil+uwQ5wQKxJQAb6jp5p50HjFyNiUw30lnLhRy/NrU3MQNZw9y75N66BAp
Aigy2gkboy89AbZgPibmMyCswxbDTWvVSwKkkriagdITNaNhW2ywCCW/fiyI5aT7
+3EUjs6FvaVZtefim2Q0KCjvmvP38URMp2JYAqlmwilBrmaUwaxd6OaeHPQ3pDNc
p3nOsKfYv3Vj75RXqcdER6isrPLoGoMTn/WFTTTKpr3ECofjgp4mrHeTCMwWN2c9
eaRAt90VgNiUbJ8s1ZDnoAS2z+qnfb9o1w+sdddZWt3mQ3Y6WjMjK6rPiCLoEK2f
aVvE0mPL13M9Pww8ox3LBKVDg5gEOgoLIJ0O7ypc/0xn1J6842GzxITjSNRxtndd
otkPBLw05w4M1XKNBlthX6ueV2/7haskpd1+uvf9M0ZF+y90a+s+AdSNKXvjmPg7
UzPQipsukaZAWL2rfi+tvLt5+vi/NoCE4IbQpkzMctKwDy/LDA8723ZXUEhzzE1I
`protect END_PROTECTED
