`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahLL13Ne+UXHrM5tOJEg9LE14BWGGu5pnP/XEwXvyZBHotSG9y9AHXdVDLJ13ymF
jiOMxQxXWqyv+BICf3kgLB8hhNkG3CAfb/cxHPsq/a/4Dt3rB2lK0xhf3XAQ4ugx
tIVSV9fv3hNlnoh0OBBdWI58MCdnfwBFWKQq+1ke6zjK4L+OLns2C8XbzEnq9JIZ
lpswpEcBYkWfrMZBH1OnuR6R1s0xVq9nzPnsC+wcNg77ClVSvQb5z2P8z0YaP/4S
cVcuFPp0NEa6O2tSMcxZ/6xzZIPf4GcUbqi1WvxaAplUYXBDk+uz0x5/9D+4n0GJ
AVkMULohNcZGPq84JgybJpBHAhDZKkrvIyXTDLHpVCFG4bwY+JX0PyFVj4IME8HD
lFYfJ1Q27xBK955K9/7GSOXWYvPtKyn7/B9YPiFzQ1tELbbUENdFwY6igCgCyZg9
nHJ703hTykDvoH0qg3xcr4ZsUjh6yC4YTKGGXMM6iP1Fe1iRM26pooJdKtIzJloD
iOHakiK/9czpYFQVOFaODmjdL2qpSKT8OCjccbJCgXoawOCvpfFhrnnigXgH2NTT
B9md7+e0Ci/R3NUXQyxEM5LhCm34FJBuHHMsV+9NUuVWDjdd1gkEbqZxaD/Hpvr9
PWwhquz9s64GONgq30VVujmg1D5S+784XQuNqQaM9Mhd5+4GWKx3E0+PMKQp8AzQ
K5OusQs+LEPC3oGwMhhh86EHS2HHN4nKA+GHG1BaPOYlQ54SoyC7h7msV+wWAUYR
JxGghcgMqvi9flXpYm809xG3Ppi7Lczxu5LYXpldXjJZ4i5+gvVn0Le0gd6ldj//
ZuYt/UsuXGYyIOKHxqiMoPLrV7VmiA8CGv3L9EoCMSL8RY4/YZuMN8UtRxFK2Tht
4CxdmhpkEeL8e6Gr9EIFeSxSHrf8rmWIIKvH1lAvhw2wRLZLv1nBd15BjV51ioNG
gAOp60KDOjsfjkiYCNhReNrhYA2yMsrGh/wttkeBXzNfAbSfgb3aemwJiv50g68o
ioZWq10Jb8tsQWqVvymm9H/3Zqnuh/0CCy/qtC8UT/QROGdPmfB/siuxhmHLSZs2
lVriY8e6FVYP7Sx5kR7OMuvRsJP+5k3If12+Dq/7xnAM3e+3UDfYZ9vIeg+QC7oF
JmLI2HFnauYAR8gC52uh8k2zXfPhwUGJmqDPcP14Ka5bK0/nueLhdansS0O1Bc4x
n5lVlMMe8jB4i3IdJWDPfsocjHfNoECXAypqsjVJtVYaQ+5wMGJn2HIi6jVY5ErA
NhMgGpsXy19dmSoNk8G1QaYDv21oeGxiKZ80opeXi77apKhlvo1z3vYerm5TfPxb
axkasms0ij1++nyfaR689RtYCa0PGN/yu4w84oHfz0eJQM0cW1M/AlPjZ0jjfUZ4
mdMQzwoIduI6nqYsl4CwcWMYOeBR29MWO1gBth2uPhtFdiNzd1365abI6tDic7M0
P15J8uvDC0iuy300S8Cx7KIc50p+kEvgi710GP+Etf2MF5Ho52S9mzE4+4X4Lux+
XozP2V172Acdby8QlcuhvqCQ801xhPSMf1xS5Z4s+N7lT92lNe4tDhTJnZnS5w8w
JkSHoYONPIexOZ5jDyki2VC9SY8/U9LEHke8ocj0BQjErOi9xx+4OxWluvuwX2ti
GsBaV3vmunWECAi9rvmcMrKeywJ3ssAR8kfzfyOXZYYT4tnDRruY5Y1WqfvzPfk9
pRZqmN1G18jah2+H3bVwvlzZt1taIVqZ87cXnSiUdn+6mWQD5WOsSKtdg2j5WltN
4WJmrqkDNYr4TV+6WjwWHreLOzwd6xns+7p7+Y1JrtQJI98ZuIVjAKXY4sWWzkaK
4l20/wod0eKBY/nrHdotZw3x4uBFp/fPNwzo+3vKMDwz1eRg/APGzMaIVnFH8FbO
oW7XModIjBp8OxOCaubPmyThYl3KLWY6+SowA5eg79wMWFQQo/tj3xfFQGLCP1iz
3eYGjBmByZaTtYChjcqxMkBz6/twL5AVgijtzBSJl7gv1q1fg4D84Fd0CXW18uKx
X43NXrqF53IUd+cCS6ttvfteM3rDBh65L8Qegy+UzX++/MO3tnv5SI+wiM9hzuGl
q/HbOQY7Q0IOQwIwu5QWh4KMe8KGKQON2iin/ZFHGxBMceP2OHwsAZgDSANdD3Mu
AOHNpOrfkRlO3+ET2uVfN8wx7NQ+ybMqBpsSEgReahYh5f+OUA1SMinnkLD6SmNa
Mxk8Kvz2naud6wt/XhlVkbRcWI0gu7gi70ZJvdLyed9z9oiFxDdOBmI40uP4Vl2j
qtnX1/k0e7U0cp6tKyhVxfsUEL8lc+XycsVtOSpdJnCkaNb+FiYxxVFDDvA3Ixd/
c2FabVFbQtjzUPWzyGoy44I/+6lnVjKRud8BCZzNmMBnQnZtFETLtfPnQXsmpeti
lgcafUrLUq6PflxiKAAKEFFv+L5WDf5Mmq1h5EwjVYexteVpLADbIGhRr9OxCe+l
Q8m0LpOsyb53Z1QIL9rsEAUrtG/kP4X1TWR7LP2kROFQSTjv8xBeuo/QDr6uf/Ie
Us0fGrmsCVoZvqdMGx+IJCj45PxgsrbWPs/ROEpWfZL4KpkjWVcbRPrQqv2vAS6i
PKIrHPCb3yGi69Sj+Agh+90TEQjLArQylBk0m3WXZ0mfaGpQy1im8pLb01XVjquI
5B6XYM29RJnEocMgXtgeoXETpPn16cKJzVe/c+T0DYEfQuFt4Iz3fDf2ibdeO09D
P4CbsOqruOuGC9uCYfjJODrJOtWTSju647YWk4pn25RLvl55UbwOw68/k8JF5T3n
AZNMleQjzDOOHUW0hYQ7yLgCHp9i7qAYp17APDzZ5HnREUSxiW11LKNNFMKQ4qzM
icLFYz5XcqZMqymB+Zz1e93/EmxUiyRNW7PZZaNNxdpvqeT++BZ9MW5eBhWG03Jb
guaUwRV8fRSkUIFV4D+47sQh0t3hEflPmurRZNrFQHH2/ouz7wgMVfVc8paXHKXA
6D6ARkl6qoBtbUTaGf01AIUO5I5eZSqEHD9GYBTTCdBLzoeGuYXs7sfBFrCuAo+8
hHq2g7UB8l6jjD64dr0ao3/2DyJb3FLivqu6os3C7Ho7JfTWaTJZEKkgCPh2P8M0
9Qr9EaCSFsZaHntbp6RqyjdpNlBeyMLnXHpJaiC4MxNsDtWR8EXHGrBk3ZqO0UGP
BHhYiSMp40jnU+4//Dt/ha6UL/Jg9atGwl17s/lkpETwSDDZLRenLPcXg48OKbcq
I448jrzNp/riPdUzw4/cqx6IZOSNwp8+4XprS8PsapUHhipY23yYIAEs8hA2a1+v
a6h0jW7q6R4hIBqg3FFBqah45eyS+b1TMqcif78IgAwryiogN4dA4C44Q5mTUpXF
1jYDtZiqiXlA6qNJyjKYfOMDbgT7WEfIjl0iKv308+76qno5g/CvX9NlgHLAlmtJ
UFhagdt5D2XU+PYpfkONZamH2ezbyPGf7WMuje9zL+TgOSc0r1vQfCzWikA8OuJV
elAXI6ZJkPTkreSF0UtpdMj9ah2olr5VhYdySMqDITszJLKh80SpZHbXP0spy1Qp
fUN4rMHGOjyM6Mgw4YfmUQIfABUGKVd75Qz5udXmBQQt6ckXiZjpTCyG/SRwXRkT
ZWwF9xqx2lw1t+Jz4JeXsNL4/0Avndi6QhJuQuvG9ohpF+1vEwuJNRdBgEZq05DP
NYC85m75S1rAtEK1PlIgEz7HFmAACsKLulqwj17exiqijTGP2ea+KTdHn+iAVZO6
OMEB4LBoOOZCA26nZeYg+Tbm0vZpL9yu7XkPaqqSe1Vx+lVHwMqDTBUAX58JRDMp
49wAyVpV1PG740TF26paU+B6zkD9l+Y+AN+b8CPzkWqGCDuQRYj+0EzeOQWXGl/M
Ro/9zZE3O1mJqIsspGCrVCQiP9d2n/t7aFxyjUKhM5L3IxHDDU5ftbkEaWQnXOUe
s0uECnWVN0PtRxvYYFBbnb4KXhHy1Aqb4jY3JskFkaTUJHpO5SQ6KcWF4nZhr1vq
UiWuZBjXh3SzHObfJCevkKDufBsLCPj3kDefZ/FUlEVMVgHZsE9xRC2enn/1zscu
BWVYFymQBMlD7OyidZGE2lTg2Dwgo5CZWYW3Jt2u/vHd0deDp6U13T3RA2u9W7Pj
aNmgcwY5B0cD8GfLaJ9cFhC0vVmJjl7BNwFb2uaPfOeoxNwqBeTbmz6cFfrg7Ijx
5uSBaUTp+B48jkx0y5ilXLYk5pHfsWZH4DRDaZEiPbhZPqFdSQaRFU2LXwgVDxFB
SCTCqAYTBEqNOfAr/g3O3MZKuZ0tbsCMcQJyhy+txzHBaiKBnsTVzIADv/YKjFUn
mu72pyv7+Jt+Td2Uvk7YVKVfGv48sZsZKTmxPbj0gupPqXQ/y1zLH6XgC5sC4oM+
IKS2VBK7SNzZJgPcA4lWYvxrzx8qnx2lVVIKGS43//dsTs25PZGG6WPFSlI+ojlo
ARm4o6w4t6yeqj5+ikBTW425g5Yq6foezNeRBLfrXB1nx+DnMogYqA9sSWoln9Tf
jBHMJRpSYo5aoM+pZUVjE0GqWFQz5WlTjz9f+wB6g8muXy17JUtWi370iEqykv/b
c0nBsyDaI/Q0tj8tB+DZw5ibUe0RGHh1pwbsaIqtrnBNUIUj2nlOcj0TNWuS32vK
jcE756oIM0U2TIwQgABVtv1OKtBZenC4FWpaL1p4L0Wa9SA2QFLw8f+s8k3w3A3B
KkkTyJW5bMdevxSzUdkLvPZZcycWLC8FVt4b9E49F+/X46aM1zBirj9BmNsK1hIf
F/sMtCV8rDBOgEHPB4ZN4zIdKoGTDilQieGZUsipvSEq93WSHxXoe6H/pzDm4u+C
0DtfR1qOvlNUeMNL3/tXaQVF0WEPvykwC78Jv7lii6WVPovkkEBm/69+P5a9QAOF
xJNSRwkui/rGywgHHcNLGPkGruusZu16Isre+AaUET7qk0Y7nZiEvO56STJixeXQ
RJZxSHBC05nRUNkq5+TNGjWPu3782CW1cwPAN+duvhrPwJPcArv1v4fr+jlRyHx4
qS9f1KuZMOzQyPLkvTF9inYL+49scVK5EgshuaSPK+qaxuO2THGNi4iH/G5Qqfyi
NpcgBzc5A9wCAp7g5jU9pCuXme0SL9WLqRNA3CWvfT0bI2zCQkVmKi6w90tymF9l
qUN8MVTXb22wtA/0vlCzZPKAAztsDLI2JE5XtG7axCC5gWLaH7M8YVDy+nRaPYDF
PkyRn4MCpd5pRuXC+1bZURoOKiqwtsHPAHNf60U0RSUM7QHG8ZvVYwa6TOHb8nzT
xmzjGLs6wlgUx04cH4dE6wDwK/B2qrvzOGAIFRUPAU+Z8Np5VAGU4C8hwM14JCD9
n+SOT9XJsLAc7ANLZrCxkavyFWr3hJ1p9rpzhXY8NVANnut4XHbIRZ5p2oHU8EdH
SY+J7hzAglHAhPXO5R4EzoiJ/mGubBrb3DQYFFXZqEMUyeZpiSRh68tpbb/M85Gi
UgryOO47TS11sWedTbZVR454zPIItOTBRK4mrAzkM3LtXfwHlEFLm6gSBDmUDZV1
qYs/8ScRPCNqUJ6IZVzyfHeg04RtxBfJhyafHMiNcR2buqz9U5G52baC/GXrmpHq
Xv5/HKi4fpnUIVk8zhLDGKOY/+a4JxM4QmZUdKUXCaQbXcfLZZvOF4MzOiy2hHDs
X30XtmjN+tvBCW62nLZgwO+idYu7swoGhVO8a2Pbe7sa/logBJsPVZHobKPTKTgl
jhOW5A67IX05OtmTBuxPDncsyHZf00vQpx4MtqPawYihcoDY8RrlHymyZFtEJMUP
4pxeH5qFgX98lYIdkwjPTYgxzzE7yPIxAjwFw3PGEXfAGFuiDqX07IanZYEQtDq2
pZlWpAs+SxaCel/jwysljh4PI4OuRdHSQKBahGKyWv61nco/r2E3cMAV6qNZzgeU
8G9zzrS3igxj+slKdqmJe9iWKdYIPXg5DlIHpGBN0zg0YNIFjOCtCVLB7tYcQHTE
BBPPhLG4kPr28GKl3VjpSxHvj9sUsWlWSx+foxdUZ+asj/RJPEu5tAV4gUHTOAK5
obQKxc1KdmpgGnBQQDMRmnFr6Helpj5fBVGCH4cNy/Ill2EB1EpV5pCBFCFBVzfM
+Klukqi8lpScyzMHdYqa9Vx4vhvIvRsumHLgkeJOwMMToQdMlqVofrU4uNN1EmUE
6tnwsaZZG0kgV+D9v/kOGPIHQefuara3mS1tE1OJ0d8ICBF4/6LnGyYnYvIsmvTj
yBRKRTQjeqeJntPNw2OyEpVHzAEWAamR48wH5yU2HBH0F2kI90ZtprnXQg+zhCsX
kKwRiPoXHxlmvKN4V+aliH3pb/e9qibUi/jqhyEkyfFhCB9+rtmmJhrUgb12fOPp
O1+dl04ebAjlMvggkRjQJtCd+dHphFsiGuwnNHAdrnFwuAA+H3dFZq+w+ASAdEyK
spOZhY5CihtuPQGX+gnWyxRhF3t6Pcckgor3+c+/kjM2xfFZhgNsQkumqmyAsW7z
tRq6ZIW0CuZWAzrhxNDMrNRRzDAm8eKJgiSG8uCdxSchsNjggtVSkS2TRdJuz1AQ
aV4dCDSBIfRgU2GHKhWoErm7XpFY5gE0t777t5DYdGWig+/8D4yt1FAoYxwUaxNY
/idvkr74sonDKR/DN4oFM+6AqzXF7Ar+VPOSQZqHlOXMGKYaacCzUFNmoojWsd1S
flMBFI1GXPcPz5Jx1u+f1Th0N+9Kvg27d8M5/KatHeDueUfniPB2nnl+rTaxkNz/
gNDIyxehQeapm7WXFtWPxjieltQQm4XJ41MnOJdLp5EtP4N1FJSwzBiCMn9vXNvZ
hCKHjuhUnXCmWCg6KEvdq8EJcD1/FZ4U6rmHyD+nRANb+9SNk3T6WGicvzrZwj1g
RQOWiQZZm8lsPZSffbWWfNd3BYXSSTEyEtRrfDCJZ/L0zaOcdHLN81SNfNJIeaMW
zCAh/XEhNn3gP+ncV78HUbpkShJh13/Asri22+5Kbl8CDdbO7ka0ntrzCyclzAEX
UYc+d9RCaz1+ggESjOG+uNaSbjrC0//HNh6zDkhmA35eG8TGAwG8Z1wrToWVXSFy
InkL06br3ixiCRI7hZnSw7C6+AdQieYM6L70dFEXTWFuyQNO3odbGa28romz3/pC
kV2CDzz6rSM5uYCPkbob8ltekEMbqfGt2YZT7ri+r+MDxO+M2sXsKI4rYv0B+VvC
aU5BabGo/6Sp28CLGCrz6ymv/NJ5yVIaLGQ7jHjyDTPTaUoLC9AZt5T5hRnSz/dl
DIbRSYmxNtu9+eEkrWH0XkzVoPxZEPa8HKCbULBjyBg1ylSGlp1IQKX4M5XktfKZ
tpfdOvRDSRJjiYozivcO4sZy5p37LLOIQBIsrFHjltIoJHY8FcH6wZgV1lF3EZVI
OL3vDouiMmnsja6Hbux8YmSPiSMM29Brfy6WMRT8gzSyuOuxyrGr8snxP+tXNVUJ
RoWuNTeOkCcn9XKMTTMe6xuvDrMxV9Jc4gidp6i1q5ow1Thf+FgcaFQyT/+kHfLD
WSMtk1mdrfkQEbTuOA8SYgcGwSR3nsPdN9wr0dQH6molcbzd2vU2h2OeYMYfyN+2
FTcTnx329HgMEASAd434ZV6kdA5SFcwpT1Oh6OH8yAKJYtthSVPZuF+7OU5hrdKg
0M1w8FmG6Qx9PinjuLCylpEM4VKZGs+tenkNIznXbfQRRLqJcsXmppx1jYLHfdfw
Hjnt2SL53Z0h/FViH+HI1pUJ4VwmZMxfPgRK5rgkXnC2ayVwfuVDbVFnLTv8DhmP
W4PkxoPysOinqJwlmHinpy7ZS8akfS5l1O37GPr896YTL/k4Qq9/SXNORkM5k6yn
QDTf7KcB+90LbPhFk/FLGvjvzmCADlSeNGzo7QaIp1IHtJ0b7DrV/3ls4/LxO2MK
4TqBuWNcuEhCNPF0L4Y9RfhUC/oXxiKR1siV1o3Z8qYUUNnvGvopRcAHpkkKFawW
3Sfx0uUkVzviqZDtT4nP4rG7ucJVO3ZFCq/qOVGgo4OP0SzHizulNR6MorJgrGkN
WF+bjzf4DWXjdeve63dF6hPFmpc/2/dZsgv69gbg+iNHXWsXRBD69vOpHg4CMfcY
moE6C6LnIH6GXzFh569fl8KxbONKrv5indJwkR/nW1lrPG1URrxDrZ8k5OocjDzc
wHsc3F/ivp1CwVQaq5nHxkGfZXj29wUDhnTcL9GbwHIi9hwLeUnlsrn98l3dtXiR
CLjArP5GOoiVsH40ERuJqOM2xbsI5NAYFFRUnQF1DloAvhSpKZaxxmrjbc8UidRr
ig507p5JQueVac6dZ+voBJprYKxRXChQ5QTlrE5Dnvju0gKMvxszu5oVAtGxQY+l
ATRo//P5A8UaK/R4W1O5MHgltya336Ap3lwL/dq8Ru9BtDy0+LSdnFaoULIcRmRd
tIr5jyONNt4tbAlpyfIWoiJ8LCYaMURrR3cuhalfb05H1CdtOmCZlbjYsiADyQLZ
OppZk4Ip/FkHxDBkCuE0TIt8eccbdgmmFiektusOqQc=
`protect END_PROTECTED
