`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KAwWH8xJfI7Y7yU8vaxpWXFSh4CFsyat8Meu/+KL9RP98lcxulUEAmsTeU1H2Zfx
1uaf1uUCbHhjnSjA7FpTDNWg5sxj3OHFLzHDQhnc1yk5q9p5GrGfq/MqyiMhQfgd
V8V0TWVwegHo6iHED9SeQIz9nj9dXOjL4uuSM0v1h0p0YwCphrYkdxs1jw3uhLJE
8wlTIPE2HeOoY2KV7J0cAY0NhW+dEN4MXzkS9y8eRT9u9fJnaALylPoObYhEmf6v
j6TFWWok5rJFggi9VD6AqJHPbnW9+H1wdugiMBLD9BJxrO5CnSbgwyy0Jba4+nLy
aS44g4ooT2+yrtUe8sCzqSw7/STL1I4BMAmRdfPUaIWbSwRcrLVH2e7fGPYtx00Y
EZrzqGSHRgOATcZoKW9xSnskrJtNlLZVMyPQT/orBbJt0meoJl+WNyOrSp56Ramr
H3lvSAEJEVQPQB4BWS0fI2erh1aBMqlNN315K8xrZajrukPaCdzjXRDbX1LNOutc
KNyJIWAf0BMYlVITFQFcL90wFDNSyuY+Nh4ziMIQJuyEK9kX+DpeshqUp9skSKUz
kSIkumqx7+nD0m9WZDYXtb9LCCeTzAXbAn1axLrxS/CbW7gwyMIIeh3RmBFngvIr
rW6WxSKzStyWsj7gR4iSyqoKmwTV0z0uIMz7jZWwaVaFGwfPIPHqhrygzZD1SKTj
rL74FSCcdTJ74ZwbVBqRTIdrfiwqnob3FkzpbKzdySsFlLj9R1/OIMynvBTalwXX
SfNVQwt0IUInMBeNA6kxKIhN6yWe5BdeKkGdHU321nafrPxhz6La8uQ+3B9nAzcA
I5BtLzAEY6DUklUEti223sKhA4dq2yzGyljWoVE6XaAAywOMhqH2tukh+oTUV+4K
yqZOTwMlN97y1jIeX8QixIHL5JyCDCdRPXOP7O8SAIP0KZzrOz9zJ/2VIY9MiJ0b
cBM4jGOACL73MT0vq8xkwlkVYlU3DQKCez1T9lFvczH3I/15IXOUfUDntiCf0R/t
BblJXiOIbvxO+xuci1OZapMeRTvzdg8YsUAu9xB7INGPBGH/KhlmukMjrj+FbTf/
9rIzSszr5wA2nxNdyxLPQLjwPIl9ZyATxpYYEGmjMe4rXr5z8cEG2IOZgoARgHE5
53yiIqYOFnhtbTNModE6nv6tt2PPaACRHO2h6xtnleKrC8/MEGKk6nw1kV/RQff6
14YIZs2xVbTd3Dlf+68yq5rOyCOP7aASaRIb9yCcc/P1Ug5EgJtYLeXGKoqw8fI7
B3gE39pQd09r4IjcNVpkUR7y2Hzx7ZD3j1xNufdUWwgxGpPaqB1OIDJY3KlmpUNc
X90KojJCP5CN9A2JBopZLRLtFEkbawHCgiYOwryf/SHZjcQGBbKIMGYmEFpD1btG
tRvpfxn0agk+AX3ci3lR9wioy5a5HMaGFY0uyb6k1C+Q9vtXAtWOP9dqP8INdUgO
mmPzgLdFAakTNzSwRrLEC1P2PaLFKLsP5ittefINslZiEX0SDjderc995HVEuQBo
6eRMK8YFTCtnkq8o0zHrLO9dLssRriq2J3XhreKPZJpNmUt7I1/1sMlhwM7OFenj
ecc5ufvttyNSRWyU2KDLMwUgn8B7jz5r7w0gp61uHa4rnFEZEjt2e0QDt7QG+D9E
qyWBgpKlCTWGn1H5Crmu3hc8fKx3jQ2tUtLnrBDZ3VTI4WrQoRgqm+43bKLjGAB3
J4cTwqNWi6hc1gKy6U5QE5WQwvi6g8kzRyxwLP0cYrZ2aydTAmAHGbTZ3ykc42Mt
iCxjstYTIXk+anA02mPuaxODV3ODPL4jeMYZyna+9bNj+Vq97FmpbiDAbIYRpA34
FIkpk4Gk5SSvI2GAGBQAc/g/ASWnuTyXJzlfw4b9AUL3I/CIG7I5MWWvZQLh7ESk
iC33BIujY5B2EYKY5fCvFMOBbHsWQIYpmCR4gHU4Co8FYWCr3+F/mZOLF+PqLMJp
8RT7Ghbwa7Ok819F3e99V5A0SGRcPMyCceqLq9/L8aM645JBsF5SlAU6L9CDdFLi
BgFBM/LYQ0r8NsH/6TsEGu26/EvN5uvuUMdnEi6/Ix92jXQ529TmRB00+BGq7oyl
yhm7EekrP66jczpK7MotO3Kg/4ftz7pheOJy/5HfXI6JKW0Ck2afBr2KRzZt76mQ
g1eriNPhn++Lplq9ayEFtQfy57dVNzgDiCU0oi2znQjkC7slJBOIDl3+lKZpbQxJ
0vZYyWIGF0gWE6Yu00J9Ag==
`protect END_PROTECTED
