`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4LTlo2jqwgkjKXWlxfO73o5RGNnpHpTixmeyFx5cdUt9Dr9K7V8G8wAoMRP4hcYk
Og24/Euz6g8KLoT5v6NVgFYyuZaLg24+3XdpxH44u1gGeRn6aoqUMjSL6t1bMcrE
aGn6CgFYwInrRKAxty9fiqF4D1Z+Jb39bn1TbFKjkZ2JlPTZpDLwZjCra5Ut28Dn
BIXr66hENf+iL3A3iRy9K9xALUBNq1knG109UAUiO/R7zUGCCoXtpu6UdAl3WhUv
jXQvEGuzHvJ/vDjNfJZ9sYRoCiAA+2H+m66QEVsqEtEgA3h8xCulIO0TSIuo5sRy
jF2x3cQ+4pPfVrhX5Olx/E2kSAx1pBjxMaSbyXQEIoZVxo4gE2wMe63IJ8Du5nuf
tHivrel10pg7sQMOIQ2o6BhqSp28zCMB41xbClHUs6mXRuKjVJT3pCP5opq0d0RL
orLQdIZgFKQg6zP5low6zLY5AYYWvQY7H+ktVOSZLv2vgyqwf/KyHik92STCWcfX
I9btHu7n8omftfxXXPA4MgY73pgy3473/Bn52heYGPI=
`protect END_PROTECTED
