`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxYod1LB77ws7w1HZfEl+PsGogFQx6g+W6ExtJuPCWJYv6ymfKGafNuqHpfPqHFU
TIsJ5GuRQsmLyNET5jzHR94wx9ijXEtG/a+9EN4XlR/+fGuL6ha7h6ebirZDnBe/
k4E8eS00VjAJ2nJYWAi5+ljyj6eQZfWK67qSkuSfqwpKdD+J29R4ncIXPEifR5Vv
vgiOlV5tBmc4I4jjstOAra+M12a63Rr1DJitOIRI9dnk5BnMl0WBV4yGFArxeOxR
LZ+IcVq/XeHe5hVMzr8p/yYS7q08EV1JpXf4FGBOlliUGlfi5FVsxvrcQEMTdzQI
ergLELurxFbi+NBQml5tibm8MJ+jyv5/NSQfE+inQo20+cucKvRWMZFkAjrP8aFn
P7wnTp9VsbKCsbzmv53tcN4H7A9xaiNnPWxNUzSxI/l1QE0hsrRRYTus8B7tpXOt
kGVxjyRGdtT3R5YzXegn8H78szLrgwIklxv0tbRn30DTFsgGUiiDPKv1DBqwc+2b
FORLD2J8DSHgclhNhTtW24QH1DK/nqNTlZME71sh0VhfiNwwRYsh4ximlegqrnI1
u5Jjpuq2JYuP2zGvzVFftAu8OKnrd/VrZSzJBajGd6cBMSidK/ccZiCgDAYj3YS7
/zgXqFCD4qvpPbNBTerUmRhpmegqtlOk5fZ4qeVB0ZnXnpXtITQ8xOGO9yw1EWEJ
0RY5WnDlPGPATeDTulCF1r4hyAzQmP+yepi+voQH9RH9Vk7BGyeEx66iIc2UD5nT
JedlQ808XyRPnSfGz53YxNbHi4b0g++nuoWKsRwZD07qRQmoCa3fNYzGoVXQREsx
gp+Tt30TJA+2Z6+//T5UtmV/wimGYDmH/RmJJMpSrt/ia5fvSfg3lgh+lZ89Q1Cd
lWSFLlypnjjL81zOOOrI3XLjxMWOGOfZwtJxHGkah8QrnrJXZhcHfnLlxZNhx7oq
mM0eO7JQQyqlgL37C5A7w3WiG2ptNBQsYPRkhOvGTaC55UyORbZ7t1KpePqPpRi+
GLX+vFpDNZRz6SGSfu8J+8vigqJtQNdjmavoXo+Y4X7a8+W9oTplZ5ZQEkuY8yBP
c+PFzETadduCCWEAyw73Xp74KlH4cunj9/x3Btx9tvGUmphBPL/y5oh3RMUzVN5h
g/zUjZlsBookoFM3VtjQCPoqY+Gue1CPFwsvW4/NAp+0I+r4XfiTCWjmuWhSVZn3
BouFTyNEYEg3FVlUKBuh3X4Qheegs/TpW5daB3xTg05IGQGs/IzYmTqsHPtd6F8L
B9YwuFur61K9y2v/+7jqugDGwDmI102wlj78tiMayyNsXhI6h4GlNEMc73j0A7yt
8S7r2za7nNFHcrIUjFVCJu0BffQcysX5OkWVmZlxwWrCYqTmIEQNHk5b2CuY+tzD
n4M+aKyxupfIYNHHYgQcshA0kLCXiyFYt6a4G1jg8OriEBjADwFbP8RiFj5K2TaZ
KsF3VeEnjzgH1rP8NTrTisEPiuLLZXVNf+6mOLsFRBnTJwOth4tly2ZmY1LQp/cw
UTpq/ABV/JCxRAaUrM5VO5pWhgkDZbyjToe+cIcHyzTZ5dWyp2cJVejeZAfZL1PA
mHq4vANkSP/0KngpxrSu/s0S3v7OShqpaKThbtanniQhEsyZEZ6dYTN4g9xMpoiX
shrcNezgVQqNxb6OclC1FKFWSOlcQk0WpirGchvlFp2xxnxCQUEj3KesLKqsDTDQ
aCdV7KHo20utJFOgwfJ1GIOlDKqhnzZonIs66N5J6zB7OfcBrQCHKREPILzw/xKc
KVpm7z9DNEd+aqVy/9y+BjCneaJxDyeDYxQ/aZDLTmFamRdX6lgd9HP7lGkt9NU+
X1yN2Sl3AhRR4hxBhSyTK5RcEW4KK83uUDI6oCJZUTMvi8MoR6Yr9ybBT2PE0qfT
4cnzkArky02tvngzAkYzIbA7/+vd6sXCjyNF1TyXr3jlHcSsF7p5XWwHeBcGL1hY
zJ2tjEpimJj7aEtvf7JJDQ==
`protect END_PROTECTED
