`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kr+SLmbMFKhZ4U8SDdFOSi0guCOLSIPXPx4IzqSg658tcrTe3SFPCS5IH6sIbfgR
MUD+R5aANh1YZKDfBSEEZpjpW99gynhAvwcyzYV4NNfM5D0wH/IqThLiicy15p9i
ACp3GwbN1Z+I5ip9Pqy3qFnHfVz8pYhQGMY9UzCZtvNqmYJtPizHlZU9P05mZnl2
s+JHBIHYBZhYRlpUjWtxAlMmYnRMgDzNxHl7DMfnaS7p6UyZ19xdtcaSy2oqcrLR
iTL58LbreoATSRmVwVkbiQ==
`protect END_PROTECTED
