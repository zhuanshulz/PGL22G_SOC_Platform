`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9Fe9D0qmYYmBOzXCf9MTcLmbO078wwYGM7o7pw3U0h7LfakJTGzruiJ0LHW7u14
cDhiENIJ21UbtBjL6LOsHLZ9nx9DCpXpCwz+4Lk2PQRI1rlq/4rK7ZI/2Q0dssut
jxZvSUDz0jjELPd54P515mmICCh+bD9/5LqU8d6JTvndcsaB4fgyjqS0LD2yRSvr
Rxv6w5s9UdhQvqAMAWO97I9YtvfAB2skN85vCViWSS/5+ygdlKkV8nGEZHWaE4kc
yvRYNJfo0205H9peKag6PBjnnB4UyW86yt9yvmOXy0tx76YX/f1IcOMqX2bB62AP
ksjsI8m4VG/HJMDFILQ7wsKq26TwUZRq5LHHWD402dZfxkQGBBw4znSv8JTyMeU9
GBTSAfNq6N0CdVN7v0P3+SS24BCqzJadou2v4gVWgBxLUSo8h1gu51djkhwTdaqa
VfYrzrU5BWDpIt1+FJbS6F3fF1vDCBNUJPCcsQFQLzsmFuKksCgBc+8Pvp9SlFOF
CoO9gEZreUMMJHImuVkjUeqlJ27orOAgzk4ztwXyB6t+qjTHQ7gCUhmA1yRh+FU4
JRArZtuVeaq9OquPJQ3sEHWs4xTfbF/+z0yUpEbsANtjnJcT4YuJyv9Ab1PQW7lS
RFzvUIORbmGGLweX08f1ZnKtECcvxobt2vNfWHIKOF1gGDgfMUaDiU8kldQJjuT4
RHu7Fr/19dG/oo9xtCuOolEpgd32VBM08R8yeCTo0Uzxoc/GzJQig3/NXmAdyWaI
jI0txa4NQuKmru0XbLB9hxQpN18KTk/8SjNyyo3ulo5ILnTUnXUor+wmHEYs9NjR
biYbOE0f4OfQGHZ7+2pPu/V9WqQ5OW5wUyFNBZxctoHZbtzVAV+qajR4f1IxlGA5
XcYf4V838rHEWN76TBVvTbi9160MfzZAwcVdmG6S1MQ0dCVApEbW9Th5sV+BZRKy
53JtfNH2D3IFtdg8LJnOQ/8PkrYQCpgmE83+TL+YhEKRLl75YNov6J+YkA6oOoeV
wDee5aoKWtbVLYpFcI3/knbLPHjWt21QUYLcl5WfI5ybeGJJZGt7JVvlzrN3mPH8
YyuuReYiX4RUFIO0hpX48SBBktuDCZusRPfZfubOjuMtsWvkop1dBMgbdj/Tj6w5
jthTotzgKLCRgkhgWUOayl7AjwyqN/xXPpMx17CXThfNGldkR6ksiUd3A86+aFfh
igV+OFwA9lXUFtRmmTyDJ05FEB0y8eQbLiLA0o6BINuR0KhTQmQ7ud+fjUQZaHkE
c19Wj0H0HnSCD5w0Ygy73T7ctEZYgwj83a37RFSj/Q10QEZ8zqVXgyXA9CnhVuA+
JRQgXDlPp075cdEmDnTrrLTLHT/H3nPk7c9aOXYQxLMkUW/q6qq6eBhH2+bzoeer
pPGIS5jxCPinjWZhH5b68afBP4aNSmWlVHoSpjRabEufW5xoA2x2nbU82oRQnhsN
+BIRS54tALE3jjhq4czoDQQxHdii9uKi740Bs9ybPIlmAmzkzTibdFjzHphdVaZh
QdAgn39e/pxm8IR2XNA5Wn6SYfApMY6rJox/mmmr4v4pB9DuQrnt75mRQ0Kaez33
5w/IyZTiblsWbzVazRL7fEolZtksDoP9uXmSSC0z+wIcky+NhmcIi6AJvTy0SaLa
bYIRDubVXyvQxNBpUtoYQZaIccxlxD7MiVAMnjCqkwD2dl9+vI/GeNYws4noDMO5
cX1cn1OBawhZ7Lsf85TK1cnb0oVlnBRDDKt+sZqB5g0wU99/HEJzkPuo82EnDyZl
uITrDpBUxqlnFbamwVcZYGE/DQEyCwpcHeAGXVdNorKIIKuqTVsPsJiZyRbcihe8
ClPSzeI/lV5oObWUT5ARq1vwXIBy7NUMz/TEV0Lupp57BYLCz4szKpFhEaKPPsJv
KwzSonZmncs3/wrqk79qZ1hEQovEGFSapMWT2w9CxT+tQ2QArndYXp42uzqmE8l4
EyK/q/gCHAus9NdyeOmnaFb2dVBe3JvWTtmbGN1kWAOhrYN0yMVndZ8wbpbicepp
5ocr0tUh6hKMkbTeXiVFNxPKvthr2eIEdgZ0LWdoE8Ks/uRL2ZtDWT0cVN0Lx8EJ
LIVqHM3/ZgLlwXB+7ucYmwCcSgKBEXH5FB0h1uxTZTihwJuAOeRp23AGEn3T/xwS
5s7GxAk8oIu/3MBaWjGGgy6YOimuB1EhENtk2o7OSY8MWBJy5zy3pbq+xDO1d+C4
hZrEFgbATVv+Mb1FAtOBNeE2xuEowWnKmAWOVlrtzapnm7mdZORcyzkiKIpyH8zu
A9rA91MRj4N9Bo/xltNdPGFhwTJYG/o+NPTIwvnoiJiLoUTZeAlpSMwEzDwvC+pz
emdL+vjjPRUjaCeNUfBHVhyixXA3BULN9NHq07z1RU3Hxq5P8HuTjEjQQyE78PVo
imTvmWakD8CWgJn+/BqOEjIZyKBptUw1WPMvVMHH+/lEzTmRZ8FYTofzEcLsOBsv
GiUuccXXt5j0mLLdmfcbRTjF/BZhwzOvHPLisHZP57iRzl+UShH99Mkih2U1UDxR
yGjIXmUjtlkpYtcnoyUvQ5I4F0CcwigNzEeKq5LNdnLqcIuI6SrERA7Ki3eeUL6W
upgjRUHkckAZkiJBV82kFSSjJURKq+0fehy/Rpd/NPoi5Oepvty4cQ8t9GFcS2z4
jRQl6cUgFUB8wrpryx4g8lmgusQLzDWZwPp16IE70yrk4tE4tzQYdWVvhuvQ8Q3K
fX+ypFNi6ktZimI9Z8BKZfa0wlp2h+taEFNSydTQTSm+0rHmtKQlCPYW3kWWiZ24
GvKROL3JztaE7RrNH/r1L7ZXynqU7Ye7csd2bxy32u8jf8KKE8vxCVIO7TqIK5B3
irVb+VOQ7kC5LH94xPuLN0tdkwzRh8H/l6Pe5v6G/qR/BuIeNsWVSkE4TggvbXct
PpXs0IWEo5/8oG8uDkRTFaBMaHtpofy7wMnEtvJGxB3UMXlop21rqLHX52NNqC/X
55OzKmC0RLozLSNk6nFpUVKvLeNQjTDly9ModqNb/ac6VO/Fuh+M1ebDXggH2nLC
gzbQEKOOoGZMWfWwJZU6uQMSUMhyem7fesOYgNJ6PlN9mw5+BNTrUJnXhtF0tmyi
Wv1YO9u8ady2XUWLylBoe5ufzW1zaqbKOh9H4axle5XGsxdYhJp4AhRmxu7KNYpd
27rJ/RmERIqAOPqTVsbH3YoO6m7l29FH0MIDpF0djmZmTnzzFdg3qgI54M5Co4ab
lfE3zhV0sdloTrmR/hHrLqv3HKxDs+qsGpXlsQ78J0Yg44xbxpOC+gvlOFg4inUO
wppc87yOjAhodhSKrjXkQRidbHTvKdBhmhlILInPEr3hBx9pQ+uRyPxpeAjNhNBg
VAAglOp6bsqolE+tp9QHp51aGYfnuV6vSyhy5RLR8dlLdHdjpPiHxs7SqkP+XCa2
iqvCML3nd9gLRPEkilQ/rTHeAkjnAZpKp0yCDXz67CvkUCWgliev5JRxhjYXkyuo
DqpOzFsF2isjVuylXgyvXKk6CE97Cg/w/Y7YoSlsgYYM+PZ3aEhmD53GGICw1xIw
pLhWL8Y/+4XZg5/P4s7MYfCXuEW4opQ0GGKDKqknXFIKSs3Pdy24r/Pcymq2dSO9
9kGY6q+m3jU0F3LNVX4k7oVDGr1Cohim/wzVcNKjv14I5ozWrRtSfGoxseXePjFO
c2zJUFDXPgGJ1VU9UF01ZrQ71S8mF07walLFUGO14lAh08QKjI39aLGWk0TgXTl5
HfHWprHvdnp7sPSEmhffS+UeqS6A6UwPhqk+xl/P7JhB/mWUHSxwQ1RzmzSTnIvY
/wskM4Di+CUMlhRTKLgzi3fzLuZE5Pf6Ju5UAD4QuRlhIIaAFmXkf0LxVpC06nLn
T8TJsd5LybQrvLN19vJgrQKE8pilippA+EtUoMKeQ5Xsk3aCIvKtya1j3W7E3Bgv
OKemB5ciFLnVnEjTMf18z23fmxwn+xsPD56Oqb1hjW5lyc9DyMfAw937Me0Di7s0
ya7QeTvB6+JQnRhqwtXQfLcPuoQP7/lJesRM58YpW1Mg561+SzHJjobgSf7IdPtH
5Md7Ehz9C8h1aOmJhAWKbAOUWY3oeB5uePnUkPiQiMVFz/CvDo+LqTh3PqLSPqO2
BPFjvHOPCPstvsuX+t013XyycmgKkLkzfNwJlVRGWpSGY0GpYEq/xRGDyzQVkD0P
RKrF3YFPDlG9j3OjCZOwTa3T5T0s+iOkTWpKc2DJ6kckPq6K6JWCl8YkLK8DGN3W
TZCxkJJWorf8nW9jozl0Bdo3R4Fv0qxpOfBW8CsuPu0llap7Qg8wJm6/0z/gj8Pd
Eam0qsPsAP3C7sfX+800MnUnPCVPt2FEWgzTYvWEKbSl7gRSTTIPs+XW8c+VijgH
UkhG7kOolwxWlNWiFRXgHC+RI6qXbGllbwLTkzyP/9SBUiL+1TDpD7/q/BqIqhdL
x1d4pkiN7n8yWqKCobHI2I055tOCkpUk5OEX8F/HNs0O4tYGCCJZTXu5Mrnh580s
Mbr8ZaH29f/kpD6AgSpixXsyYFqsNp/kC0J4NlEcAMbmyB8X9+MP8KRXvzsxVcce
dKODHD5tZPtK1PqXtW9IxIRQsiee+p2AI1BWSbqKembSuVGjnBd7gGzXHjFEuIfj
HQst1jtvDyJRRNq6tHT5px6KxI1sfm2OCBvIASW4ZmdW6KpaWWeJVQ85jOUPqF3x
+6q6WxzJT75SlpEBo9gCNJGYA0QQwSGnwVFe8HL/ukIuE4TbF6FtM5cPqmIfmnXt
4YhX5OO3o0449Gt0LI8Wd8KaX54cW3p3MrieruH93mvXqE8uLhOa12pb7FLJ96xM
2irMbdqmbd+0RvXICf4SMlhe5Y4Lu0lQYw9Iwgk4ooGnuT9f/JK0FtNBTecAahDJ
4iwGJ+ynOUBkv99lpMuWmfaDnsBNJJZFbgGFc+an3XJG5CU130n7oA/Gl6p4gbSm
Kg0HiQ/V9QFO9rCdAqP2WM3Z+4dXybZMjWuPO2JktERm3FiiMEBlpLxoAZfiEU7M
sCOvlVF2bjqZcxmHOuYReWAOQ7iYvw7pq3FoKEG9RB3tYE+uvBUSVXn7V7gQJ0FR
0pDjCpTKCGfILWqmOUiJ4svsRAGduRmhlnKxFMQvQI45B3Jpzq+yA8tETepZ/73j
oyTv/QlMMVlE6LVKbAHo96gcFyReYPlrdjPxxb/+bRL6AC/EskIoI+Ug0v00BNWM
5c9tgifLfff6A14R0yM3rVzPIBiqYzCov2X3fjoJhqDiYMMxMCRA2yRZXOGhJkt7
Y4dr+8Elx8ew2PG3VpHynV8tgQkRMV9AMqgF6r/IuphrKTsgIO3ZGD5wWOYkMBv2
8ElxbnobY4/NHxNfbs7761SBKwu9qmn+hUSAuhA7/rVZh8bqDRotCp2GFSpeoiWC
+kD9ZCPomSBLw5QkS7N/MIS8orldYtc9ZSDelPy80PLiYCE6bsN4/ZMNCaNZSyGQ
oVTHOqfb3loBGO9aXsGmS8+Lns2sVrAd8Xjuzg+Hlr2TXd1o0Uo647Wa/9U2lsUd
ceAErFEkVqZz0UmscVrx8JVIg+oIwV5E7uV+nB7kmS5BTcfTvM13t2vtomZKxfOj
hhCb9/cc6L7mmomFZl1WS06TSIhUcg9736+4kFGb/r8OypOuITPcXc2zU07kFKRf
J8nYb/QWgvzYEg9VvnK7nr9may3qmAc6s9zIwMn8+x59R1EBE2t8JgKDDSG/0tXD
nc4WSQOYMXDxlvPI+5FpuFZ4XWmGQAH7s6lQDtZDNbMXCA2e+naWpDKaXbsYfHh/
oMl1dbX7wiiKiIFDKUGC/z6y1WqjO2H8fny15huHUZgEOvTKHSszrLTCiMsu8PkE
EZ1N3pxdu5q4ReCWn94IRsiSzcsWsltNnywRz3ZqlQKVSIK5YhNsQjEIT7HcA7rC
nKkH9te6vEvEmVu6XiVjqhtOuY4Ll1G0wcAiqdHbatxX9TJ1jGGlVBdgpgi5m6i0
vSKvLQ9Bjx8nLIrwOYazCkmnjsrIXCKDY1nVU845Vw7S1EZR8d7IRdId8oDrm8dl
+TqZPpI2pk0P94U9qlL2s9MdYqWIvqYvsxCyp/4NkkYC4NkxgBsdd2G/BDgSRU5g
eKkFnUV/0hVSra/flpUiwe85BMsFxyC/YSunHJuL21zTG20ZvnU9fNXXUrZDyyPk
ofcNMxgqrb2EP2LiRmpDHl1vXbMRc6z9c2QKU/09yzkaBQKQCUSknNUenAt0BUvl
czyPJ8bCU0SIIS6EZ8hkQw9k/7Fj3lKdHhha+JrKSJFWnIuCg1ODc5emCGkJh72P
yYD4eu06LDqbugYFIDbUyE7slhctvjn/PnARPD0U+rU3dOXM+LGCX5vSG27z+XeC
WX0ON0puudBe70/hYkUIBwfRvGE4FwXUpMXFU78RTa06DqHIqD5/gdyL8ZoHbCHk
GO/9zcsX0TiuwnejKkXzzdJ0L66r0LrD5Ot/SZXtvtDlig5g77nSLV5xWDn1LtuH
Uh5wKo8aPmIwgCbsLQtc9MPfYIonZvJykC/TyhFF8SX5ocqO8DXWVIhSrdyE29pr
GviTmURnqyyEIU5gJQa465p91ahQcjRPlwocsEJl1m4V392gSbFWOjdQae+cWZlc
9ngC+Wt3LhnwLfLNdq4muLksq/VFba3djWXkEvynze49ZeDJ3CodTFXEYae8l1Go
GStMU40HVRp71zc7WglDXgHcNZB+XwiTcb1DNyM3cOoplILjZvaP6+C4KwOQpLuI
2FdssZ+sCXxKObNpJfFHGT9SSsRI6TjhgVjG3GzCg11AVhlc66MpOEIKvkacB+ER
sHO2ndMOH02G7N5UzETMEm6eSMknHIcyMoaI18fMydt6BhZJntuPvC7a4jHdqCGA
rWl0xi79XGxf1S9VPzZlyE+iYnxvOIZ/cgzJDt7YDGXWw4NuFswj1WEKqiXOtZ3l
onTIHv0cPNnAVyZwN0h2cwq/454O+D3LlIuVQp7ZzswS4QJK2XiQHUvJnNoYbPgl
uYS8kQTwABlAzeBevTA4sxF4Qqq8GPCfZgYDkTlBwB7LYaOzX0rSQ+CaJh56zl4J
s6JXUXDm/JBBsDqDorUSIznvS3aFglvSrhjvvFg6BMzPaR/OcQRziJG7oIiVLX4V
6WU/DNkJUMx2SeLeINLUGE82DnVE+r2/3PME346vgSP6N+6FB6MeoDjIGSQXUySu
na6p1Yuefikw+D6u4XW0/jjQaMiyt+qQPiJODI7ObOLFum0z9Ye7Z1NqfOdSHpeq
+k4DMJVIXxx6y2PwA8NhHPi2Htm0qHCMg4+ZlgKOFnaBqzQ1oBQjlpcQSN/EefLG
Xy+em5wq2DA4oIbX8TbY7yvaxaesfpIsJHnNx51CFLKm/JlANW1syVcQP9xtPlqV
di9EKNlxe6YSC3pNuN1Bdu8TuJHEGGNc7kzYyELYoJPbAstObpSYkAJPYDHfck7K
jlUv4wA5RL9LCiBsot25HQrTgwRc/wkq1SNi2dUCynO8NT7oeWF/QhmAHwq6v7NN
q0G08KHiuQOqzitiqZqFkjhiEwlPRjJQcC/t8uazcrevFD7+yj4UT5IQdD+ZW6Lj
LnZsOJqdz+CEjopGXbtqZIzywgjXJ/rq/k5tGuH2kdb89pV1mBTGeaLIB845SsOS
LMWN1NoEZRPVMcVd56gRFc8wZiNr/xCREcmyxfCOSQP3coIATuUol37aoKp+dHPx
Ct0K5b9ilE6mliE7wUbNBoyFd4wAY/IV7L3QVHkKBPbx+U1VJEcv32AUOEpXnYot
R5Y7oqGjdEnJCvHxLA+srQbi+7rcn3EtzcDTBy/H1XAZiGzl0hh3v5I5YQD7yjJd
MaAnl3CJyj1QsXLTfVmrcw7iHHtklUyHvYQ2IexxzhsI1MyAlB2O9z6wqF4Eixtx
7e2HxDBx9p9/Z+cZ09yy/jYc4eAjucfjpymFcPer2rJvIt02dq+tMYO6YZxscKqL
4eH84gOKlKzlgoRUHfI+dpGetmnbyPlZZx+3ilqHvtFyZbeqHCoTlz10IuMSpNGx
V+SVQaX+bxVYpVYjCtYAIFrHCqP6t5MpnXxGUFN1pub+rIBEP1l+u72LTNckhPtN
q7GVRrrYq4tryV72VheUpVGux/HJ/VSqB8BHlQrtzWMQufZZhF6HxzfklAT15vYW
8v/A9rW5RXUADfsNdHXtR2kFL2sPQi89x7lx/Pq+ZoL/bo8BLx+LLBcbNZ1m4mpX
210Ouf9anWCfNpPGmYGkKsn0z5xazx1whTovQcgg472zKmdmEu+o0TCHJyIfBZdu
t/flCyUI/eimLizk+w98y9ABjPN7SsM4VA5NhfdOal/auaxBq3qCEVI4CzwMBuTU
YEsa9Pc6lx6B9NHP3kZwqVC6kblTA/T74unEWj1c9mfSuhL8h107cJBt8XFduT0s
ebkbxVnqcQ1u1/xIxuWbatCA7fbviO2iU6auIKx5mjEb/b0t7w8rBoZlVVHX/YVd
QZ1RY/k8orzOqm89h7aga1YWrREQK+4aUDXTyVy23L0+ivlk1xpKdHCvpYWEzCaW
Vwl3Yhh9Z81dP09XCFMD1wMNjZHh6NYDgoQq3S+O+XPHoB/FyY/u0uCjuxW2X17B
bIj7dxqzKgtiJn6zL8PHAKHxElZ/BTOP3x5G8G7XMKkhh/sgFI37FD1RpWeq+alA
vOCO2EYm+CMDxNtXAcanrOjl6hjv1NbmSfuu9gNrNKIMLIFLbF3VLvDkpL50EWZA
NYyzSD4CGk2z5S2o142O/JbTaE6hbUf/J6bkIyEw7LDfJIUGGP5oTBzRp0/O6jYv
12CtkGH8BTE+ZCbs0RiYhrjnVG6R6nTE+ACqp5xgeZa00s2gzoFlKeg6VQSWHU+P
rjniNY8gTg8v9VsMpb2BthTIjUMxRGcyx/SlD1eFCSPYEUCx/Yl8OotFgdbyOcNQ
uWiAC3LUv2FBAJsnVyf49V6o5O9QHJA0exEHKQzLJz+ECE95etbtFeNXrWFNt5fx
KFJ4SuQhFfHaQxRthLW5VKV1lr5W5s81GKQiHTTjPfAZIiJce66VVLDPhGrCSooh
FMFANZgmRzR9CVstBMNAOdGRNFmU9YrRRnb54OvOc6hkzrHrivAl5OJuLIbKV+Bz
kx96jR57OA6+libOJhMqlEKawlrPp9pTYJUz54zRNKo0ctGhfIRP2M8OuKxc59WG
mWleK3LFLUwUGutwHZ+73h2HnIwsdEjI6bdyrfRARv0rcSLIAmEWgGKLfuVMCFeQ
0RdFsKIHrjRGJlTpPK5ZIlv1iK+M+xvwnSsoj3o3ANbKqcrpo4C2kNHHPJh13d8K
M0RUdu9rbT9Qt8zDBT5zs3ECJjGBFiX0EyGulufuiBgY0TxHkMFGe3IstxdYDQMg
XSxUyZMr37vAxUiypfGaTH67moyzKBQYv+4WxJQ1NxHwPCyCz4c/9NeoAfAKrF66
6Zn0LvLZf61YodohlAKyjavcylXtIN7FWx3MKJts5c4OX12zGz14r+s4ZECopBuh
jmmR4GrYgCNj3Ib2zZ1uKh1BFgnypvRDdNZD0/kOS6pyNafRu6Xc3w1GovLvwlXz
cGeH9vavMrtS4x6CfQOy8+7s7uardl1whwUfPaLA0yuJiJ1GfhCJX7qeA75f/6Tm
6rHqHn73rI56ZpZE/+y8tc0vLc8tT41LrwQtw3j5jUwIb03cl3tR02VDaOPRJIWs
LSTsoRNsbVPuyBpLNx9VyZa3C7+n5ZocvvEl2xlpC8KgWDhjttkn8EzDJ+rdUbj5
riDhkln+HW//7qwqlCRer/frGcxY7S6JFv/ZDJPbltiW996WbsmEU+zswe1mSePS
TwQIZPhjB7UKq65PPnD1bLCfn90dWCrRnMUl15N5G+VDoJOvCqRBlJLVnWqcZtJo
bTzqHgvWHdwugWY0fBGU1b6wf+3FxXh2aU4K4Zn83yQ59QV6Tn9M9PJybLwW1vym
CEKMOf2uurFgvSvDfWMlvl2BDNcjFUJ7j1oozzBJUF1H0vW+zhXZvVG9TdfOH/Tr
j0UIeUgrW3bdPm2cLCmeqvfLLcGvS5ne5FwQ5pQs9hMjRfJnRWHhm77kPaA/6fKc
qyvF9NOoiSM+O9u9ZSxofS2dCC7FBOkB5nAwGD/Klx7/lUvrpIQ8HjuJmMzuqjwU
AaJWY7i+MYatIcu44MQiyBlWX5GFXX9VgflTefHzzhFf7Qjf22jW0BSXrc9z9pgn
8v7DY6929niECN0iECSbtrNgyS4GUA8XZUb47PaMSgDv6DdxwQNhFMrSjMuctLl2
sazCh41Lu5Q+7MfnsGIS8BzNPsATPcURGeMObrzVOaVlDet1AqQlTO+eRwUG48qg
EWGBu09a1WmHDqHv8VoOeW7Fa2sf7pWZYyVE2jZdLAKodcg+Hj7kBcNtm/zWGJ0D
2cZOcPSuGQkeqHKEn/YeSSelzLs+xu6Ib611i7LiiHUq/Um1vPW1Ukm12G9StszI
WgGNbliPzrb2lFERde1tVt23vM+1pCwWjgX9EWFZB2a5lrzNG4wFODEA3xr0ID0e
fPnh8Z9JdiJbackAKNIgYaNZ0aZgBWEni+O7Pix1TIiYOWvOVU0A0AHk05PwW3K+
UGKHVESIhsLT1/NXjxBHKZpM5LK1qRDGQie1NiUt5Ps24tJ57lpYlwLSvlzR6zbD
SNiB2RV8VHj2GjEz7+CpqKPfEcZK9O1KEQbfusICDORJ4BQ3ULW3Sl0X37UPMwFP
K78VVpjpwk+oLcYh6y8uFGKrft6VxvYvSmR/TVKcd/R5miPphiaiZLOY0Ml756B2
gAwNHXg+OpFjphmZKqAp2I7e1Zu8pLwrlEPKpTadyvY1qVACESaelOaIF+Q23TZh
lH63TlLDOmD65ZHGeiaU1aVaBZS8co1B0HZnzbbQ8iToeMkQptgSuvxGUwQ05+li
JncNh3QqqWBJYCWzVrEU2I5q1nad4IuIfB+RpcpJfC/m5+Pk5ASW7+kIHXSwA1hE
jRP3PpCh0NF8GTfaUBSVX6WXv67WnbJHdhNrige8m3EfDJLpikG5zeo6t6gVNU95
hjAuPnEty45bWClWFWe8KU8t03fp246MUwpilhN3eSLJRhiAt1/pBVLiotViKSE6
OIxt5LNGqqe1DhO9HxGbTMoZypd69vXUTRw+FoNv+UUBF7Z6vBkbfA84gOdFFrNe
Q9ITLajPzVfzF4N/pkwWSDdUNkmu4DnvuxEAU7Dwwmss9qjU/6t/OFr8mexGw0fl
tU56VPovIxpC2vbBakPh+ikeXqF0FVzL3oydOIA8xHzvUxZiqlR1WtZzHBRlTpXt
ewqdQqhMCrgOXGXM2G/rIwNK5dQsbONP+Y/zDcly37HWGfuDtD8mN+Dp/1XyrQlG
r0CBGtAdacO3cKAip6PED1cQ4deVqFhZC2jm2TMAmzjc4VyE72/TrzGZRG6dcZDS
yUbt6R7+2k06f5ylqJoLwMY4G3A4zy2OI/t7QFWHDP8Tj6t9lOzTf1EdkOY4h5d2
BHBIoetnfWHjW00Gz67QXLOhU/EsY3qMmV5bHh0MyMcEvtlDJH7WtF1IeHpCZpQ1
zPg1NXo8wUSyt1X5m6TR6/NyLHh8RGvtvhsMjm8t7sRsw7s1ehYEg+OUWffZT7O5
lA29Rx7KlomaFIbXD4ZeZ3UJw9/NdNjrkvUjcKfcQ0IxWMZEyFhKeqzkhq1901vO
1aKBowD8R1OVA67nIgjzj+Z35IlCT0Xm58AlU2cNaiIUEmCqW4qd5NhpVJxPMyps
Fdoc0DczAgeVICRg/WK2BFSSxmNupmrill3aF+HyWW0QupAZfbe0FfyCzE4RbhQd
Hx0p7o/8NTdR4GBIvqtGldZ8HXKkM6ypc+7zswUULAPZUFL0bp3B/8Evc6eQ2lAD
jLfxK/qTWQs0ylalI3FgrYoaYFlT/3QNtm0HoO5Cm6BcKSbUFksNO2PiruaihHTn
QEcpxZDl/FuwkrsL75aiIcvYoXX7i8x81kqr6k2Z6TsCPIDPM2GEapeuR0i88MKV
WhQvkO55ckshlbQFKKfrIUhb/ykdxDqQMlIRILo7bS2u0nr63Qs3mWVs9T8RNuXi
HviVWHTL+lOO878phj1ZehApWBA9GytkTFkbFY7vCq2uk77ClrYo3EV/yp9BvmA8
qPQDTTM2NwVe3JN0oaGzD246pFLCjxvxy5Qy8iv8BJffgUeDhbLc6w4Dz7AP7aRG
G78YFynXy/oZaenAuEAxiBeST9y7mY91DoTLlpCoAyO/iS8TYxP9ykXks7RlfT1O
20E/nzDamkDBxoypqI4ZM/p7RM3PeJlJ+YTKDtcbgm5t8EoHp3UK4TLs8OX011oF
CtyAsNnnSrAttMJtWP6l28GpOr4q8BrWc6TiXOdMaR8/K7QVYhCcZCSH16aMyxsL
qoMeL0pb2PXkcfre97Rn1qYz2Y7TC0bWOwPLEmSYmA76GFA4+R03hHWtHEosG7zY
LpWqY83rZ3mTASwvrr1Q3IV6W+VEm2EYgX+OfIaYBd+B0fTK0w9UBOOt5IJ/pGhQ
wpR/hnv82QZFMEBycYuTWK7dZn4xrPBwquVR9UjXaOhwvgBGpojLQgnv8+G0IjxH
JZ0V7UDnJYBl1OHiOQ5h2MqIvok4wgm0NDgVl9jvAvBR3hFG50c7d0hS7m4sl60Z
oddQnfrKm4mWAUfQNEoBgWBEiBvpUz9h9D+ka/Nw323DIDvrVm55GE7kx2v5dKD5
ejmVzx5M5tSNq8rLFRVnKaN56s0y8xbPMcigBXZcTe4RTRiL2mnyv8Osw0gTmxsk
6GcgGqW/hzufZWqeKYQFawG7uZyoxcWUehK0VIACYtVo6w1iDH5D8mJlMk6Q9z4Z
Wq3lucZ0BBbvc0cQk7+wRSMXLOLfUC5sCkvgmCx0VUR/EY0r+NyBvklqJET1/R0H
3hwSudRHEfmuQiNkoCuIx3/KCk9J6eUetT3AbgY4rN4uTLnuNZsQ5ml1EeAB8CCT
ewqQWfIxel5dUfeTBoz9tc/815+A6hrnzpvDpouavQmi1mhPukPruK6udlJP6op1
qv3Mrli8pcLfl1f31m94MjjmbzI0yR2Vg/SDwPIL9Vbj3E+WBpnwX+zT6odJyhWA
1LF2+oxgSy6Mt73CTK17I0Ax75AEpzW2Zhdp/6vio9z4H6qeIyIzAb6NyVthyKX+
QjQCDGOZ2UncFVD6wpnJrBlwdc1197kcerqgv02+Yob4KlBu7FZ2wviHiprF42Jx
tCFnDFNjCoSm74OpZoykRXHaGBTy7JU1zJYV8Bf/bqe6qnImLfCLWoQPmgT179+7
MgfFSyGSaMzbRLpVrTu/TBQvzNS9AeECzVx6KnwE/wmfl3/qRUjnjN++ILcIgTMc
pjwTHbPWebZBcV81jP+AyOIw44vmvApOGFVZ2YA5X0EzD1CigbFR4EE0aXkZqRse
ZhkGy4PLtzM3QDZU5zef2As1BxzXkd+YNeU7jGqMeekvHaWQ4yBPu4ihLpJP5bcd
dvKJ3jii30LLfonyP/Zb28BNolS2MJSzO5ndCqhGRRy2UmH1jGc3P5zdF7b/uMhP
DM1OdixiFy0iUG2keFyPq7svH07z5BsRtCd6xtYxSV5zF29xPiIvSxR8LUz5vDm0
RwfeYvfHtUd+uO716sfuzhkV9g+2fpKHhtkcyn+X7Iihcp2L+hYjlgGSjW3aACKy
Snb828Mwfwu41yvtvu3tXZmjWSspZ5FpeTM0LrL8dOPDGgIqErHNKIcCvk0KRZTm
1SpUnoKIpJgliUxBYXyK73drB0doXQ6YwvkObotauPA0mfZKmTlbCqXyEpMblyFd
QZxLHFQXfCbpzYppv3u5ASZREw9PK4qNxDatbCI1o43ND4/dwJ2Pb6v+DvAWZN1T
VG+PCMrxLU2CVZHU9Eoc+pOX2uxDEE2sP7E+awkcYbeXe61KZe++y3VWklmMc3iz
l3KiOJ/JLhOcUs4LVcmXpRhQiOnyE9ruUGWPsbJ5YdrykHqyKLmUbanhKL+m2WHb
n6C47jV1tov7ZO8EuQgiFpzJVu11E/FBgmhVQz6LQugw/sTu22h63Pvr6I/CsQ8E
woBArVaK5ZXNTABNJjeXHVGgSpMbFkwOV/PV+BGpgAHKgwwN0Ss7FITtMlLMtaHg
LEnGzSpASMpVyntljtmdzT5hy6LQN4vKx1kXmt9FkUlIlheOJcRzcc63guWJJx5s
R2UazAjbB4X43ECdeinRfsr9E3qQ9NdOhmOa7tVLQezpAPl1eR5v8o51ItJWz4Lv
sKYgC9zyfDdPCqsLzYYdyUx1UMUUd1oFstmiZuDcF/HrG+fqO/P5yEUPkDLF4PfZ
XMkw3YRZZSLEvzpGqHrEhETC3uflLYYoc29yrloZOD8Oz1fSAHVikFxm1vsMu6Me
mzo4QSnj06MDwBrPXI31m5/lib50s72sfWK5/yLyVvJq2/yiaZlM0SOSZ6YtjB79
laSqJnMxB6MtAdKrCLk30nbkLQ+L+SeEgX0DOQ2cInysgF9MIqH6MP4P9+DVQGyo
ZFcO5xuche0I6HuTIHGGYL4pXlyhmrqxoCfcqkYJe/+I0MicIYc/iQ2OWVT6emI3
eJILhUBRnUS0HiRvfl72uTwuBk6WXPAsdkfxv91B3E0pjRWxlVdnrIJjb4TX3nL6
hxzefOuhAc7z/+aqiijJMk22D/YOFf5EVLZgSvZUKTaVSx5EAuolFBlbHkn2O0IS
p4OCKcf8qSY7POykggyVixBNOkdUEQnLqbJuldpGF1elAu3sW9zMOWJxcPXPNhKx
zB+CI/1Ws65VPRf8lDxSte/LLNU+TwGDI0frKbhKOWRD17AkTzESEO0s4iJsAV6u
C+YoTU36T6p/MaTw3pZPgDGPm7XCSquzHVMA9y7Ibs6/HrW3eFJMz3uAH3B9xKnx
6646Ggn7CzqoipQLE0nco5lfqVXhEq2gz0aBlEWhOnY1QLCgjI2cL7n6W87q69h/
YSh3zxXDaZMafAZ4IUarNCCmVpdf6NkiHb3t9OeupbFwvLB1EW7Gw2joF2JyCRvq
cb+C5MCTFxA+Lq2TQlNtjX6q9NbYfM3moJDnFvhP3RPb7GroxLuMZfJJxLevk7VR
1xy0WmfHjQOfskI1seNAt/74WxftvdIpF5sZjSn4q4pEVVzcz9xBUM8+kczA8Hsv
qGHimS7Nsr1ciTXQj1mVZDNrXgpmJUBB38O+NP+j1TmigbvTlmTXmcPUtM8iXroO
FoTD8z++/5LjNG5kaegwjF6WLlj54vNsFCLgiwOJ4ncjgUg5JkgJfiCbzvvNk8EL
FC02f466+uCxmrd5HUnRYARcEgwToVlMQFV7Y0XWERfHiquRCn/azD8yAS7J20i5
5shlMHAAlz0Ij38TFSfP0jN3MC9QoS7DiP2E+ZGUCfOSoLYbtdQnG4Tymy/isroJ
uOH0UMheCDqO/b7tpN2nqfSvq1o9On1NLVrc4UkHOuG0m+5rkQZAxwsuh0dGZGXq
8Osdf0eE1cwVTPSbbVCPHJONkvZDFzT6AJ+srPJEiLpDWuGHmYsitJZ6OvYx0MNB
X6Cf6f7bk9fCpAaI5dVXSsKqAmbRswP9GEosJAM4mWLpemTX1lG9iN4ZPpqsPPzZ
0ZqO7f2tWTJOeFl38O6p9oKrqs8ApoEexJDu0ly71/uUTnRz1DXkbSejYU1ofyxp
wDx8QIG5n5yur1HXJt3uZRsB3sNMc3YL5D8emOiolN3marr8eYlBZButgh45YeIw
1aI+QpO/WB2AmYPXox31/DHEvW+ipjmiwAz2P/VqTf8hjxVTTl9DIjjznZa8hZtT
vyem8JL2OftTR6KTI5C4SWVi917uwH5/PkpBECmygNpS9ylBuOVW51SSkO2e0GP4
ZtcArcBX+5QDpWru/ZNCATU2vgArk7xdCUMNQnFb8JlGfDvlBU80VdkUgPubqcUG
5ewMJdu6jdqrROfKPuN8IVw5G8NnilFPYlsdZ7xnckwxnZyzns5PxcDmL0Lh806S
F7YkOlNYpQC9t4Yjwpe+k0fjQYA1sF3wWD2v6iTBmeRUoeFygC+k+mz5/X2LgmLW
nqi2KnUBHaNHu6ux+CdvZf78DUmKTdhgG9izL6w7CwIXfcgcyNt4SaP8/As0kqEJ
36EP4UoWSy4bWfgnXHbsPEIqFcFWPl0ovEKiPvM4idPTlm1MFWAUbV0Eh0bXZMfr
336/vO6SW309SnnU1BeRHqXYKEWV1KFLpdX78Am1+JHNw7libpHAdIVR+wGv/Kun
1sVOic3Z1b0Jp7Ck8+98cVn/sM+NQ05ZXjWthNqAX1hOO4yu0n47KjOYjLov8VGd
vDJuaskhVAaB0XfJI2mvnino+emJnKCjwxYckKs0zgGJhYy/1dFaazDx+g+s24ul
kjKkDYamJtN3OEbodWt902OXt2WpO2Zjkn6sAjEA8eRz2nAWNgQidilS5RGapwZG
cuRfjrTDmkSu698GRZevd+tyF3FpDe9zyqR8Ondx7KPp9OktlIem2Pepb+y5YF+y
Zyr5RfAXyUll/rGB5JLwKIdnl9xqP3Gkb82304ACN58MEiMpfhqCgNI6Dm50I+fc
ihvY7yQVTE5U1jdR3+DtjmegBxOmKSMCcHDgARrGkSYw92yE6O1ZQ3jODSKbtzdj
9GqCBgMiU1Pj+nNnbmcjyLjWQDJW4zSDaSw4gLM1JZsA9xpHNMwkXPnH1F93UT4K
kDsu1ENam29RwSpADvEO1ENcJYpj2RU5hOPdYo9sKwaYkKM5NtYQQz8jbOWZ1y9T
chEWHY5xcwnvFj74DSFXRRYBX4q6UdT/ZzLEL75VjTyhQPxEtf2WQJUq9ul+JJgD
OGujwc+otZbFAladv/Xl5Ke/18sxC8/Xz3q9aMwZmbqByBvRW7KDEzQLasZOnuod
ZVHdgwv76AcI1d0M5RFqerh1NBh60ImzohpBGKlxXPuN5qrYjzsa0dMxbpF0mLVW
P1xDZz3Iq1ujtw8+yyJjmDfmer+5OWHpzYMk2q/rwXfub096wKjsi6jdCzf42kW2
Vj1ofQBjU1WROxXSS6eB3BFvsjMie2jaSxN8lUHKqdPLEUyPqsYJ6m+yX5AHDErZ
51TjC7OyOPkT3bdMyZjmAIR1k3LfeGpNb1P8lJoOokgNwTFtugE3XoHPAeLfUSkk
ZDWWq62a1uMTM4D03i0OsnPMQappdhBpTIv35FhriE48q9qeLylJkFeqrSKCpmhl
7SOAbAI4X8Snm8+sa7Un+dnQ/FGAnoqp/zyDD68jBXB3CPnaPOJtxm6SF0UglnD4
PHNQe1Wju68NrkErNedr7FTeRR6++AcOTrMlSX8CQ1+u/serQxQcdTgT+XItRl4b
hiW7IPDbfv9nzZ9HvURavHcjcXuu0h3oc0yhZWZzWCLzErFa1SciA/gJL5nYHkCy
LmtwNsSxMDrnPqR16+JyqTPxf5ikDTYzgejCQa9wPvASkrMHYVsmx8xXAR3ci5rf
4ChvV1KSGpx+W4XTTPP9SWMS7qtsyU7/luMnOgYaVSzxrQLsOJkYZpCStw0sqEjI
NiTSeeA71JKZW5S/SxyXLSwRXgRQitiZ26WIHDPViqblmPr48AFAxjFQw5t/OliB
cQmAiDTs7mzAu2en2ze/U+ZcwD1efR6IcazApFZG1NI3My984EKazi1Ob37Fge0g
NDwXl4gf1M/bU2mXPLO2eBp1+HagNV6lC7DuFY8Bvubkzzae/v9CzCQal/4kFq35
41RBAyOgq6fYl5p7Qz1SEsmae4RCm/n2Y/WlfDcJTnf6xR1wzoamOpX0ih4zBYQv
zY/4nI21XNnwFyUVCcs4TvKboJGDRV6c+Lf3pvcH+/TQHf23ths/0LyAZfiQyrSt
A83v4TIliZ9jwwwJOxJ7uj+w2hXUJw+FuB0RzG+0dZ2Ygt+TMqKqFp9zU71sMHoh
cCT3DOR+qVyT16F0VT52qGhmigY6nPXASq4IUOl0RVVaMlbf3gGJRFqjCT4S5Xdz
H2e6YiBk5DISAXBFrkLSy3P2XODmM3jxf1RRy7FfBg7Sl701OQvLV7v54sm//UzQ
W0QTS5g8Ucx2hbIvAwBmOVSSIAPo6uGtKBd9+/w44X5Tp+8vXYR8ULI0sGkD96H5
uxlKr82ijM8UfoL+MRSqnIf8XypzwMUvWisOZjrtxA8d9ZWpX1lBDSlZiCdg45SJ
p8F0z8OzoChrADlaWfspAYkbr1sSV287J+FCFMH4cMHsR4oi6iXA1xgj3InvnVLC
WwWJ6Eyb8OeeTL4AiBPIfMVBsKec+h5NywJ0F17phG2c37rGVKRzDMMoY0d8/Sxu
2EkiuTRPxH8ikzugAilDJbDvxSIYjUE63e+lJEZjczBANOh8GdRSuBl48LhEw3Py
nr0IXapR1rIFRD5j+DZVp6xbGdI7VoMAZewRtnyd+XorzTLUZFk3qTI+IQBqhLvj
bhDxjFWB3QVuyOl7SAlQ15xFqoz4VnG1lfvoeQepfxQpeSCtF8QtONMEMpXNuwiy
Vo7KlQbCBKziCHPEh7LLMeeb+reADwdDGfYoA3Q/e1sMbZoMaNOt7zL9WA4W1S97
5D11OWozpQanC2gCrxRucb0B6bd2JGF3pkgPhzy3Bl24M8Jg5BAGiEtVr3BmZHcK
qsWN01gyLuqYvzGgvwFxfWjRuhfhzXWD6ufWgwmhPpx9SlAfNkUcYl1cpxXNCFQi
8+e9dkiTwBZzQWjQPqoyFXVd/K2qUcHPnF/KQBupPYulkblyjBUbZUg1u82rak99
uFhoyrK8mGGzOb5tyzDJhkBtBlkOfp3/1iBzU+TIezlzLwRHTTZVbY+ljmfEuCsi
wJnXbtvkfeEIvURHeYpUd+GrPtAEy/eRIoacdxHeV6W/ndBj3vav2fZKQ6Ek/pi9
2ikXX4eBocc+8iphRHMEXkPkcQgOJj2hIgDJ3n2X7WWDLxcY14CGtxHlb0M/8t5D
nPrfZPVg8AN8X5iBtnWUi1kiJa+a5TGEwj+dr32LPWWGi98HjM3S82PtSm0PS3yT
W2A4FxlLlbiJiBcZFmqqwV8TanJsUA1yYY8MOHxolwheTbQYdYCCO9Z14+ZRv9IU
ONsgtLMbGX+9mCU9lt8HW2+aZQwl491xtrgJ2WvI/Nos+1IMb7aTfzsMDyLKcnwX
E/xZcbqfpDQmc7OxTifnTXimKF6BDrY7b5YHmJsGlqpe8cWKxqqNGsswVogDcP6F
18MXrZusBXVv2QyRQov6mzULuQwJ4mObIPBEnvrRAuspusr3jnrjCvaE1TO8JHvo
NBNJ7x50oA/UECDFKJc610RTq7wmJqpfr61r52uhF7JHa1A2rkgu5gv3rcfv1WkG
dsMcXwhnTkSMoSaJcpa3e+uRsDUn52vB9RYgdQBr+EZHD5rPSnLGUHSbxz7+LFJx
VAw/Zz/0hVTt8/XtqfJlOWl4goa64XH27EJmq+zkjZ25gg2SCcI9yT2UUZNce8Xv
8Q+zqMqVtIekNtlKM8bcNf8jL1xx6cOPkTLfkYvw1qI/1oTV0XkWLTC4R8aVJ5QY
uq0OnfMRVk8nPo5i2v8aQh0fVtA5c9ltxhpJ6BYg8aR56wDiSuXY6fljH7QwzZK5
loFfFmW2dNU8qQG2ECWm29o0QqHX8YsWrH8qz4MfJx8GuRAweOK78Rx/E5UUejTB
CngoyMO0sClw9FiYC/Ks0WmUajnrbQUDjnEXYEvbhhhqqhckb6eQx1+sMQLIfXcg
ECuvv7rq+WF58WerXr+Q0VR/56bz2LPaFSc+1/w052YnB/xzo48hP8mqLrK4rH2W
1b3qXNx8DxjHB9V1xAh/KmgUQBu6jdRV7PZgtJc5nAfO4KUGwqTQfDA60B6fY0rL
OuZNeWC/3HXpw+2Hdc81QyiOif62qYaoqCIryHrgATBYnxdFa8QW91xe3pok8IoI
ITv4jnJUo011QPT7noOEPoSQxj/atvEY8x7DjSRwHnvzfQCRzNHjp47T/YQ2ylHd
TWTKcjJ3DJTBDhwtp1OcrF7jh+ajDE/KcFI8BM5bd+kIIJP3hOA74Wi9dnuIlQ91
kOl9s+diy8W8rD3GLcFO9s0O5qBrqO3z9VLeBVAzRAdyVjqj5bWgTw8AttIZjjHf
FMOznT9HiqUD+treQVprxNajU47XAuIpAB7L/LMe66ygybFhqwuRTFW5Hx3mVBY1
NYcMcskUjF2HUGpI9Qy3CZLygcH9MbXspfwsF003EBx7+KMF2GHQEvpwx7IzRqRB
jAjcOxpqIrIS21Q4+XSeHN3xPCnHhqgyC1dhcUwOuuccuO4c6rkc4NFSf7xiD+7i
tzAgtJ0MZaqXnJEFsHOPCaUE6pofAJGWN4x+8+mhr1A7qIlfjueTfm0yE/htJQQO
XV8feNEqQtzzHPVwahGf9smGLLRoXgr5+CXFzOWzFLd6lLGt7xoTtE2No/4PdHbn
cGqLeAPSpIg0Kh89I+JtA1R7EkucPLOEuawkxk5dY8635IoB/nxmwFifgWxEYL6a
lGJBYGTakwp2hFmdHA5QeXbM74XHr44LGvXaa6oCxPqU69GDdGA/G3A+r6fMNvqM
qYo3LG/MTHXr1JSCPCb3SxcsFwS1qWoG5faRq6mMBwPcwAUWzJwpqUa1ABIgEHo0
qmbfU3cqe91PYZo2p7kArPbtLRiqxSefoqOJBUcGgA4sg7/ujg9MNrQeYXq5b+pP
ZTrD1NhDBwFYV1W+JQ8t2VoFEPeaT3zvcAVayC72RNsGjXFSV2TBcU+5T4A3AStj
5q9mfilgGEI8P1xCFOV7Icu2QGfHFu6TXNoSUJ0nCdm0xgQlqaL9LjA0UpnuKA5M
A+5UokqoxbPghbduR0nUHp+Ptnp/hZc36NRXF1tn6v9nmSAWlBiqWWW5rYtiJlhX
rFp3IkW+WJoDA6IARZoIXtIFivn0mQZgIO6FbgWkOK60T892aIrnP1hmE/vby5GP
A3vDIgeYZ5QkxF1J7P1NyVV/xKF5gRE0F5Qf7aySeJ33nK79ecVN1XeJq0oRc0g0
Hg/S/GLZcbcG/NPUurQT68JxLK9BP4nX+gmBdorme9uwAO4AXGuJ+GZEipF4At/e
T0eFApw+R3TbxgGreB1oZTv7SWwGA0kdLLDS2rjQYfpCGDJX/KBo07oB5GMkq9AJ
vn2hmWrDUWrdFE2g4k17uKYfhxi+mFRdg4y33AOpFTp8v83Ng1+yLbzzeZkQfxUs
K5mfb1lqE9iv7IqwZ4zb1lEHCjYfHAuJxDxqCdOvDy+09t17JWMaXRusDqD6SqtK
P/loOuGptvmYFTZpaawYBxsCbjU3yDq23XDobGzWpBpZerVOYlkWA2PFBL48nMvK
9ZWcLNd0BLn/ybTrEHLwEcykrxa4wZbq9Ui6TsonaHK9Ytl88aTQvqwCwkMznBgM
xxNEkXp1G5IIZf/Lt7Lyyvqws9/ARcakK7YYnq0h2X4CQ9/KpamBVaL5n4DidcMQ
vUS0UoqMtjYOvTGPcaAfvlqKob8Dsler766aNmHhvbqwmZkxWXROVAW/a3dAUJFt
pjlZItcXEgr/Xe7BU3k5IzjOL7T8t84LSUeuZ5fm8SVmZLVwwVv2CZIf3GdkjmVE
wx109pHSITnuWNdJi8+Tkp8yWzlr1SU6i5U47onbjy88AZBRCQrtiD4ybGzWGbr2
1PaByTnLGsJkXFuHQZi7g8GBqaUWQKr7QFId3CI5/HLcCZ2WZMiQmMfbZydNLmew
4taFuhlaa+JiLsMFCNHuIrkCQjSn1F3zqVgaH+6IsGyaLofKlyXPvn9Q0KBA99X9
/17Rebvycp4PD10rEhqJ2zEPGwpdSbE88PkNXk4VM4NdLzejLDFw3pEFXOool7ce
KfIuWdWNEJ0qjcWyYksNYyvLUWi+A0G0zLRrkv4WEH4Z5vVSAWtsDf/LqOX5WKsW
Swe1vdeEQ+owlCDnIhbS0IvgKINK7IGuh1FcDAgdRc/uk+6k9/jcTtXf8T/dNS+s
RnYrYJmAWWIua1yTDXnSAcze6QlH4F70qwqxBI8ZVMn0bbPUf+ZQzOpdH+9J8xIU
oddPSnGPNrAEBN1FKyxc/VtK0QmGJV+rb5NS5PJOxN67IOtfTAwhp4W4y7Bxro8Y
O81bNyytfnnSA4TlSqxgZUtEJMEwFRf7ClJQje4eaaRx3eYBxOGFHfxjNWVyVMkk
w7U185nHZLUXpH46AYBHPIeAdPdSokCGeTqAew/VF0ex4OF1fODV4Rgozca3nzxs
JBrVNeTJuBsZeJ5zd1Xd0b8bdRayMRR1kZebBclbeOKbZGnMIFhjnrxxiTz6OpR0
9Enql58hbys9gxLxypMRVE3xwGELRw6L/d/R16J/fzWkqxcEMVZqVmwX4YpK1ZS4
va+ZE8HfXwBRTilRZeY4Ca9+r8rG2QXNhigHlwDY2b6d8VF/RWvj5po0F/M+2N+U
yzWKfjDtFektVswOBPEM4undTi4IjwJhrOUrNbrfeC/ja0wbaxzOMVH2Lt+NXY8V
8T2JuQX8FQyQRljWvV4gscPzwW7Wwun8BMG/r/+83HrjBz6prKnhRQfDgFIHQag2
`protect END_PROTECTED
