`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfIv8ewbyo/ye0NJ1G1w/yGTSbU1wpE292blnELz1H1s98euyzHgLc23poFnp2Zc
kBcEazmHb3gtCn0NxNZ6tUyUE90a3IuePOivjHeMHlwQG6L4nm9NxaPUQolavpKO
rU0SEfeOTi+qCkBxIH6eLBU0HbDQn4jFlJYShgGCwoqroVTknw91xm3zysCYIShC
TMbR/e25zFsRBqMrVcvNXYfQP9ZHC4/NKrmwrBhFPeBJbwBjUCbjmDrKBOsB3+DW
`protect END_PROTECTED
