`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ilc+YyB1J1R/o/Ms/bAWN+MPQ41eNNT+F/P2FsJMIwzXRNaxHWE7ghNBYtyQFwkr
W1lF+7XviV+aoyjty6JbsU51kEFm4XrTi9sZ03dB34vcAQVhvHaRsGjg8CmsxAjz
kauzeDpW6HLiwwrahIwT9KqHH+s+rumZppr4jPu/AAvEtJb/mSDIJf7/AIDphze0
BKdtcergmrGzbDo7NMQC/b4VbEpQC4IP4dzSXNKGvKLQM7AzFQwK5H8T5JG95oUR
rf88rQWUZ/PEU7xD90iU6BWIzZ0/C6dkh4h5FODYcEwiDwq0tQOTq96wUrBBlHhv
+ruJMqFeCGa+sWUkHb355SMhh+CYgu1tv9Xq54T8zw+kT3aE14zSc7pkILkuU7Vm
xL1ozn+BQQh7FUAUcYJJHLyP09TgbPRUNVeYWtfsTVFlXNhUbEpw8DoYY3sHx6fz
RBkfQDOWD1L+aaOLqjLXCzdiRF3crlXXYM5YgSw/iSVa5Qi/iwv1+haoQoNj5PcF
6R5nW/7Er9ylnGRgj0zpCJNvimnRQCZfioAEORrRZeC7eSsMe4lJ841VeHavQB7+
pnjK5IBswALriRMLl/QWj1BimHuP/934CdATi3wHsEpiOAv36iEYaUMAzCthg66+
XYd2oPSVzluoHF+WvKb3OVmXiJLm2khRN93I1IXHfcWNuWzCs2Oe0KUUR0TRMu6+
VZ0z8nXeccGRAuOzqL88xEPfPEk8/m/Of9VedKzDnVFzaM/W7R0tJNTUNco7G7xl
7EvLW8PtD9POo/DPyOwrdA5fXG1dHXRGDfyZLJhvYVosprtANSXPxCVporUOUwDz
p0HXbiAdho7PZpawhz1UaXDMrBwq/UolTCzPz7TDlW2ZJEyfrGQ1tP6KuwdKinmk
FXez7sLRWJgusZZFvE5Z2bMwyW+jDH8MT+3q7R1w6JNZ+0VLQeJDdCb4ilybZly1
2b2ozWoK+GUii7etqSA4vE/y8XxhwePXyacHFl18rmOKzrxIrBOsH2kgpvTnc/4T
3QpYNQFjua0xuuKaH4S8GAPh2K78vr1BSxX4b5hwCC5h+tg3sB2SM5pG1ZAr+KnR
JRgbtcx0u/JtA3wR9T8S06E4xEPqeFnE7GKpqMzNl6IPJKplyy8r822x/Pv/od6W
yxcm3wkSnzfeOT8aDgOnRLKWYxUz93SKXsl77XF+j2VtgDe/qrk/YadtBWkxS2pG
wnT+rl9z6GKegRc8lCne/mLRdavBz6gQBt/lsoI7UmqvwD9Zt4hRDhI02Tz2I3ty
sSF4KgMz5uymFaSolNOHoLgvOWwoYQwXrFIL9xeY5LCJTUy/0LeABojtN4fmGc5b
JgjcRyUG5ltLPuAdujAB5MOyPpSAy2Rfa1ZV6YCZeGsqRSJb/GU2mo/dyI6xiX6i
QUKxNO73rVq7LWF5F0ZymlxITK4R1EUFGMrDe9FOLDAnnla/WGnXtGRFSPKH8THV
vmjiUhwnSTMIaW+TSRp9QpoWF/f/+xm6x9ux820ET+QJm0IJLS6FCIRSe7lCXcUE
tUTFVr32gGwkeKgnCtfadV9/T8Zx8oXvkKgJQnOog/n9nF9gTBWZTX+SjnAleTyf
G6PU8o3j7Jmtaj7+2y0UvPK//SN4iFu2I5bZz5YZx1PZVxNWel+8pG6Gg3sXiMXB
4ndGxR1PN8RTbpGZ0jUo7WtZxQotxGmRFiRt+0zE3OH+GqbstS+tvJx4uCF0hwu+
L4lL+uuRiq+HO8eB0mtojcDE8zjkQioLMHNDaH+xFqYBs2HZRi9SV7BifLeRcdxk
bDqMfntp4xbRbEonuonh588TFhNkyOe0DwVmB5ZOPo0ba6xaMKiG3LsEcSBM8KYs
hBKtJmoVXrw6OmWBK8Oq3MLQsUGv+KvZ8sROXBLUJkUlXP2VyoQk+KCt2a9XBAoM
W7XHXQ+txzsKDkmtFd4MLA==
`protect END_PROTECTED
