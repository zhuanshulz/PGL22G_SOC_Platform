`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pTey/RxStbjMtm8B8Mw6e9sW6myVqmT6W0SA+qsSW6IkWbt0zisAy63jb5v6KRxF
g9+iD5mGtPVMUJ4ojJ56pkaTciIJraFWucEOktAwTP0fhohk5NynQSWd1Em3J7PC
gWLWpc4AhWvhtawdBlvM2Ri9PjWQX+lOTF/gCh3Io1ORuCdV8ZR4clydGPaZPPga
NlHVosLfupZQ+g5pKf9M3I66FJOvhZ49vc3oU60R22ZzxtD4KIh7W4fuSPjinzeL
26Z2cEZGcAg5M0N5AyfCD0V7G2/abdNZMki4oZMsMYJxbJ1ZZqgZzwEEtYBc1yw7
LjCC5M/CvP3PT1RD9kHE7d1YBn3LuKszimu/E1adqkcuEwLufOFgT9wSI756+/80
fDJ3MxoqrNh4mSfw4k88xUNGdI0rXTO/ccCGBwCTcoe4XkKmwauXrJ1Bre12R0y5
/vO4llKYvV92cd+J7civYjG5Dbm6A5UWTWFol5XWXvjDX8cnu11T/QZw2aWi1Xxx
bnBrKkgRdXDJ8b4OKZd5QQmN8/VxfCn5xDBrQCzE9w6YA3mMoOPBjiFUqf+YvOeB
B2wD34i0hWH5DKBb8D9Bu/3I0aoQZNQBx32bVyOmD1qsaAvfsd9SDpsjOXYrolgc
pMHFSndAh4QROkE0+v/Ml94jdT6V+Ay2IUtT1gHWQzxjdDJC77qL7/c29OLR07t0
YBJjewOlP3nFtDz831kidac3xDMU8VSZK3p8+4eipnGlQbkOu3tY2F2a07DXJsv0
XFU4eBNWkwccwA5KLdL8UdoED3XoJiKWmUG5UDCGmG91TH79UhD3lMXWPTtrPEh1
hBmZ91sZjhbFtbY5QVrakjI0s2GhMFV3T7UMmuDVvVOdIEeH6891G8fcvI4UqM/T
jS5TAhKDW/xAlWoQ/Nnz5mfttlJ0+tSuNp5ry48KVFtTcQsOQsFIlzsjCaI2xdJQ
gUEaN9TEu4dNc11ntBwLZeROmOZmmaEXu50Jzp3y0d5FpMlSQYE9GjKdnDRMzqER
8eV7fxRnKGGj2Od9IxHMtrnsHslmzLg3vz2lwwfQqbdSwqQ7IVUk5iLmsBWuD07Z
y9LZvUIlkmH2nh4TtMBIBacYfkgr05/ebdfb1NEtwDm2NUUqck1DGYEfE8UlmW9+
9WunaIBpGVnyHyVoWsg45bPmXiTzhizsOsfyOb082Eu0Wcs0HJHnySICbncE5j+j
GX/Y99/RQqkhwp9LMA2NBmiJzhqelQSrMSYIbIzWpWcFf/YtymGTDe9XaHi7csod
YVnl2SOy+cT9rhQcaWxhWQ==
`protect END_PROTECTED
