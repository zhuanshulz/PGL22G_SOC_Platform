`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgLE5ZPemFBhbkOL8rvKxCAEoXrVsg8IsGp5Gu43cSr2q4EXHTbkaHFIwOE924+6
ETO1DQObdUNaJPP5AdcdLIXVI3r9S8CgBkGcNEIZOrH8RSLOqxw0Tg4/plk7W88q
ZDGoeWkLeKpdxLLVZ1LyU4BEDtZ/+1GhfTGoP686EAub4vaAQoyCk87kNS7e7NGA
nhY1E+VRHSAgr1rdPnbN7X5mrZ2DzSRAt+erjAfCbqi1vruiWxnCMun2osGYbSU1
IweN40UrnlcfxcsLPWAeIipbPj36YgFEN70FMHdNaeaDcm7/pmpTYgkt8g6VZ41Y
r0QrkPKyihHbW8h3FPzmX65lNg4vvFEXlRF4NHoTGQzaeAYeFrvwRFApED7FU/1b
`protect END_PROTECTED
