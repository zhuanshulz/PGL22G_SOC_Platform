`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PO5ookkR3yIdpn8JvLnoYuJxm1Jd8F+jj1gLdYL68eMjQBuSICnvu6s1qhynZxT5
zt0kKUJJbzAnjEmmq/7ATjMQQ4DqCBvoaJmFUGi3YemHC38zSm5g/zoAGReacGcr
VLMYSdMGwvpPSv5l9wEAXnqSTCsb4TdB+DH6NsXYYcF7eW2lUPq8J6o3z/NIjco2
anZGZgJ4Cm2m//tnHA+ftrritffHK175c9Td86wnOJ7HcHfBd1Nzo09j3XqSYACu
kLrjpW9INtNkz/SayHQ9cc2VQJp4GpsYSEZWwanLaeQxcDGAwUvVBKQpMYsB2r/3
MwxCu+HdEOj0KPQHkxEKFT/tVZ6DBCWVNdiAVJibmETCYMRcUAi15FZU98cdMTsY
vdcK0IGwZLypyNJZkCVlQLTk3APjMj8N6VQiD94dLOD9iuqd0uXno/NH1djfOyJq
sESIy+IogTRpbQPSxovQWwAkaEdH/QpNSg3dtcO7u49thljmMpMT3JR8As526L7P
NKWGhiEV5Cw86FNBK3DtlZSF9EbNEWmuspLDBHiORja52K3sRrz2IWqj6HSdZGND
Kg+XUOr/x78LERKbEBPDzrgZ1h1QDuZ+P+zDqYd9IljCZtxtbcPfDfD0CZ2USd9y
FExlofDP1HYYDMaKndLCPUsTVcRpHMapfhriAt3s6pkqsSemq8eLFiAyqz49hl6Y
`protect END_PROTECTED
