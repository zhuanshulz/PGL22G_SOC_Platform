`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHJVmFYcS6W2sCTYjVfajE3noV+PcfKw1lgBlJcxrlU6eGGbiqMH8nqDOAEdyLed
/irLlqcxZr5t5mq3npe4ZnBft1rowtKXkhxYEWBNWhhP+ArG4MUEkxruW+UZE563
JNg6952V0TLAPCzkUnFYK5ezeB8eyU9iXKDZGgxE7p0LWAwnvMlVM5VHBZZU8M8U
rF0ISTCUn5Qa+s5LQ+vwXGnAQOQk6RNQGOsfWeyA42S+rxFyawx5MbXK7ZTbm4JT
JHbMpy1QEZJ0AgiLOP0zfmQpMQE8rIeIVJla+iceADdIdkbZWEDrQCpk5M2BhiTc
z5Lhl6acEjCFTCb94qgpZji4zTKabV694Zm9wrneaR81Podud2QKVWSPNpOptew9
eQ0cjRoGg3KLTmSxhgr50WYDk0DXpIy/YiA8ZP+Hn36FQRwFCCWX110VI5se88CP
G5Z/Radio1gF2ChqD2SUHrfYBjPK0pMQHupj27Y4yRzeuThmiicv13wzQSIeQtaS
J+zQSTkp+6K4Bbu+L0+sPNtgoUpVjLlk56wOHWhVno6DWQzuCnsUIK4dHdNUlQ5a
1CiXCf4kn7jC4Jrb4T93lVww+2y72W63nu9lFgv9CVf/1qvoNUfwGdVFazDpZMFJ
DS3XwQPi/8bPqDoRZylNvxah8Sy4IByuX3gk0CdDEs0vNa6cNHkb/bxZnc5YSqxE
s2lG9xi8g8ebbeBTGmUJfwa00nAlXa8G8B64LuLIVpkVIM0tri756tyLOFLsVP4r
dAUDEgL0UML3EIggNqMRz4v4wq4WPGX6fHYfVNx7BzAqQQ4HzNDxpkllffOK5egj
mww0GIwohcTCyKlfhtEHImKl76gNirdKuR0p3guCPKobqXB5huKi1xurE11+pbuH
0sMz1tMd0Q06g7kjE1sZllsLvTwMur2GfbD60ayYr4BGI5Qe5KIGMz3vw22R9aJI
JM1s2uCX89gysPu8UfoLOIaqfbFF+de1LGv88f0txC912nuvF+fZrjZxiVSSErWs
lstJfSSJEC9Vo3zi1g2DnwXLC8VzEgkEFa8irNolpzwRO1HY9at2OD2fQWLn2DxI
Ho7QQSj4zFrXsCrjnp+GAZwKYpo0Nb3GIKZDwbJChFLyxUBuFpOYiCUz2WuJfFu0
HiYqmlub6aGOVsCnPAT6p3coKu0BPjUFTw8tJk+98Ge5ehKisQJ11ThMNz8HJTsu
sAd2NsERjOLU24oDmqRtTtZLbdDvVFH/y5wkbKS+fgxQEtXi7J4oBXlo6OrJxbyv
4ZMRnbxY7K2B8/uiOU3M5a5WSz154q4mNLj+fdRyo7Y0TwMBmz21ubc40GsOasUD
lRoHO7ZpsqhnZ1U2p7LIYov2G6x2T2V/4uBQKPLirYoO7c6Fn3bS1nw7iA80Ni3+
Xyu9wV6t8E1v9PcyZdo6Jh3lYLgYDPloMJ0Y+JWrQixcgYaQ5XOnZzqmyxzXnl3V
tEm9cueJJYB95otrfLgvm8wvnxiFt5L2tIyhhQv36pjMFY9US2+MfB6fyhgiBLMf
5fVnG20jVCds1espo+HzVUWzKHIRsG0W1/EpAxj+5l/ltj3VaigOkIpT8FDvKWaU
WgthR5WQRNdf28Nf5DGzSIAD3NS1pmYdVu0zpiUM/CfFWT8YhgxMA7ZasnSvq0HO
YPGaa0SyUHgzxVMlklGFd2iUN7a1bR72A8BS9uU8KaRNLJ+k9ZFg69EAVnmp0xWK
S1Dq6sBjKshLjdqAT7w9ipAjeNptQ1syp79vXdVqh1Wvcm/fcmZBEFRKX/Ga2T+s
teiI0moqUgDykPM8B5R0RXaRUnLl0mq3FHTfyKGO8rRu3iuq7dImsd2nn+2yL7oA
wudH1EOOcup9Gw8w8qB5Ca1YjVjxpbP7q/xm9R7PVQXfAc7TH9J7RNRwwaC3qXk8
o+8eDf1c0W8zBCCvo6dbsFJ2BMkr77d3JzjAxX6W1jEHMlzoY9tLT+0rUAvDIXcz
mHrGD4hdvjDYZZtq9PHzEjZgMsQwVvqchIFOGNrQr3JYfC7Dc7fj0yJ6G5/vH92m
q2WEencxWpbJvT0+wkvEzfW+krS1EfNte7DXTJeIDbWuA3g03gpj0B0YHldcXoDL
yJmDFsZgi8nOvJWHVLNAwqQZIaCaKPvAa4Sbrq9BE1x4YiG+wHdJQBl93wR0t8W0
iVHLXoVWonTXjfq8oOKinaB6JH64lTK+0h9RsXJasv937fPM+I2rdTBzJIjncLWX
t6UjZdsuyxdaU2uM6EHlDV98nx90aL7dGx3u+Q5E+9tv6EDXpPsvLg1JEurbARzt
wxarVSxmgXCYZKzvviPVQcID1y79hnSLH73rc2o9oIArHtQT8hVsrGcIjZBCdstT
sA7lVYuKrfiTelqJwlOsxPWM5n5DSnA+6CZXjGBSEJEqwU2npIkpX88PowXy6/Tk
kLW3H7rOAmyMXgvVFMf96RD92+LkOEntagpZHHETOAtp6VNJwBbcgeia8tPtwxLP
QckfMKnmOxyuCMu3YKZmS+fwyi42CxhMj+tH0dzTkKVIZ9PBBRVyQN9asPZKu/7w
QuC2+0LRuk5uocxHOV7vXiWMAxGgaWNd1n6vA7f3SyIoKHfGapwVuBzer4MCXKJG
/++S0hxk46gHaxIHgs/t//NtlKKZS7HIDZiI7GJePNVefuwFr6W7Pv+6eTDUUWbP
wEiBclBIUvapf9/djCeRGfrEMJJq5o5WA1jxcyn8ApQRl14FgoQDf27SOdtUPGzT
sY6lZFci8KTseHcfj9zQ0n4hMFFHF1l6GTFgHuKhAwL7v1wbfRuxEZc988xEggcW
uJazyN/UqAou0uaplOsTu/yXq/dOOABp3a9fl/Nh6RNyIFw0lf7dW4Es0UBLusEw
Hy9bBbNziNysNqLaCjabcJap88c0MpXNyZRtiGS2SECT3AfEJ/uAgiroAraWKYUx
KQMXOUlvMjLr71p2DrsLP9sW1y+LD3ku9HnX/dwSF5Fau36N0cF6UPL2rZWVQC8k
AknONhIU1RAqmq9qD9Ii5wjQ+THA3OjFBLOgOuVf9aAa5D4onT4P/JZdcs6dsBqx
ODIJnfGH4Vi0m0kzFS8nKReRF69nIIanF/YCW9sZpGf2iCo6Uosgs5+MRiHSl6+L
BAjcenXH3Hy82QnswMMlqqy7DmreYDusfQQpmha1zY13ixElZ6kFZvJ9iDAZaP8s
47jg+v02MxHoi/vJrZZZDInzADS36DF/rs16E64PbZ5CGDG7TEuT/fK7sm+/yvZE
GBFgZ5cjJJ5IGRPG5feHkswaB9Qush3c9apr4fJbKpAJDGh+HzE+cOEaDbOnywfl
M1PNOuW22m2wfAt0b9/TUM9ZvBthjPMJqDnEb8kpTa0ShBfTgb+Rp8FEpUbbpSyY
YiyHjFCTNTnF26dKfVwXGKbjFjS16h1VOG4SbscnslDbjIb3Zreic0Evk5JhG9zf
Syso6jspX9Fa7/gQvz9SSneSbZrG3D30euofUvwdOSC9+8B7k2bKWnQ6s1+OxLYQ
KwEghzGwu7FxKiawoTGkzTNC49XMDTbyCH0+bOm5DQPq5YhuHi2WYow2qnK7CycO
GLpqOzZS15wEKdXHD5jlK0ueH8Q/GqGJPl2Lepg49m9OzgnFZsZ4s0JGIbZMdvT3
v7FN9g6eGtEU8LFSuTCUKpfevyHACO8K5qVLf3+1hnMkvUj9MeTwgADEWU3qooxA
X/4eIIGot/PxDkyIzI8VdmkjdlzHexRu2AAhipJAAKAmp/+l9eEYs0Qjyr4IJDRU
5/GJ6OAkYw+kUqO0aJ9tuqhFwQhln6Ac4xJT3wxMTdA5HWbu7jgWJxD9hfUJ5EZZ
OfnqaphU9KJCL0a9wm+JG9fMvtwQ/77+6sKKYogd3vuqvd/R9co5Dz3JehXz698E
9nQmNORluqKuINqfiQTiyhFllOZPhxhfXA+ICcTyxOnFFc1V0zXQXXaPqqvAGk2w
cjvvCHHSwt1EQ4T0EBJTNCRbL0x+EzhgUEdEZO/S0j2J96T0SiTdjiApCRmccqCn
69OhD1WHP3wHjXJnr7veTlrybh3Np/TbklyS+C93CgrZFGOHTy6kcaWbkAoPqVYm
EABQdXXPPdyeo2iX2fDZ1jkZPrs1GOEJgsxGvjIihMDzruuxOfB+uLCSP3dN7ruO
K+tK378nXkQF7lwRFHptKWEvOJ3ZS57H08qCRNh3Rfc++SFDlr9FqxiDiOnKdhum
RwZq2gPFyQvjkWjcPrpB9svtXgeTHCNd4yVcleIfQ5LEjkoMaIRP0K/qiacicrg9
R/23uymNEelgkqmSYIbk3hjZYZ/VUFfktCHF00XXsop9JAqRF7UU5lp3Rgl6p1EI
C7WLSU122NM+8cFlFW/fI23wNCljbaUtSL6Em0lui2ORQWCyNXyDPQv2GSc0k2OA
Pi3WGT7bwPZ5/XmDzz6ioygG+YKyVVBHASx5sJY3VJnjLGN748sDVA21d00/tJ+Z
FK5Y3ZOzB9VC+IJ9iJfUGs/GqcnVOl/XW6gYbmujPrlr/3pmmEKealqqwdkK81OY
zpYmPbFb2AMSQw9h44H6cF8+yUZucqa1CK2XnlKTcsxm/ZsGV6/FBT0q+YGDUzyC
`protect END_PROTECTED
