`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqAR2I9J/aHKKLRaPGcNT6zkf8N761nBCfHFHqUNso4H/vPbFlGpO5HlQ819NjGr
eJ6Zhm3ILOHxOKhSrLuUX/K95NnPPe2e4BndVSA54Ed+z7AmKERFWvSjWMUEtfNi
UASwALsCXUn/iExtbKWdIgsZX6AkmCiUFw7KSeXL0AZMR8nDRLDsAG28mUnds5fS
ctuUyFd3J7KNe9Vqc1RjjWu/BBJfP0pElCoXju3oWwQjx+vw4YrvlBLVJwUrhusH
2AMBq4EaqC0VhB7JDsvTaw==
`protect END_PROTECTED
