`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2WeCfzxDdowYUrALIxwuye7pDCmArrhkfs/rcjnBvqOVVwnu/NsozZJiA584Lru9
EWJPnxAK4ISoXXu5GKV0kAAbTtMp86nrxHOynyvwIxKNdYec10grPvG1Ec+bM4Mo
J54/nSgFfYm1iOB6MDzVEm2NrIk82ulMeW8Ooj5XMSb8fX++HnlXX3v6zmqNEjhQ
FDsq0PjDijT5/0TEYeXyVnQmGTt1VZT9XHiEUufmCeQoOsM2zVo73JlHgz0vGGmC
8c5TgDI3G7RalYdJ7pL/W3KDLkCe9OhcWakNIxTQwNptrA4y5Y1R8tmqun7FU2xZ
wQaRm63dwXoub1zhmQ60k7+8dpHImfXE1xCBK09eVUKtjTQBeYxLET5m9kOXewO4
LNyOd3K2nNyfmvVMWwbUKN8cblG3g+JrCGxpffdajaA2ewOefewiXJgYGVSu3fzj
N2G75HcTrhnP2yaFdcy6ihZV8GG7UCXzOswxcIyKp4Wp+vc0bxdlbFG4Y2g0YS+d
42JECZmhIxLvoYzsAASAn/s76bxaKR73+GqgvzoxC8KJTboSGlM+USvH3gsW8ZWZ
oghO8+3MoeqIu/9iZuAcTd5XpKhHOxT3RymkLm+IAi0=
`protect END_PROTECTED
