`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1F4S8fsJwZ/+kVrzUbj7bmozt2JmiK+O4tABl1WW9N9bZOc7KMD1bIE7L9o1C53M
jZIUQROkXf4qGAdinSYhWf4u0uWn9RDlK7OtpyjYfkAEYELB6W+8QOJq00rih5vZ
3Wa28BohsUHEMZScvse3Zpisy+UZqPX96EBAun4cP+wWN4+NzdtHj/IkiSuG4aC8
RjXY0SxtS6su68/uQ1UIu4SUne6qdGjVCB5Lr5DhVFLi3j48n5WaQfreHdgJLwet
rLMVm75fV0QDnin1wIdta8Zo+VVXOoACQT8UtMImLbLOg1Rxv0XeM0PJcxTqn2zD
otDeOB9k7wlPgc/yr8pcqbdOK76aL0R1P8///Az7tF99wqbbkWo4cURWBvT7dvfe
EluCxakI6GFjycHU4KUkf4gb6v48M6c/LU5dVozI1pCoAVR19zv9QBUtCJ/vHAUj
rIzeZxmADR8YkLqMN5A0ylNS360kYUyyfMRzfoh7uS2dZ1cZVUbOjyy2v9yVUwR4
xvjxbP5LFlsacBXuhRr4w2P5oWXuKTTPgRWzsyC1CEphh+9+VqyIdYWGfJi7ULnA
fSE7k/EJsfXC2UfHwN0yaCh1bWm7Y3ZxUI56HXS/8fGKFm/g7wrDpSGQDEDlqkQk
V3ul0WfAPe16bqbRttVwPjg7KSfTH14B0tMsByGu6IhD+4+Jp2WGGje7K5/ief8t
Lb+ZK61ja66rF6UXNxgpqHyqc0MZAcQDDt+M/VBqqneBhVyI/isgvbM3Go/1a5oy
ivlAlqQ0t0B5cqTERR8bi1mcU4BbH0nQ/Ox7SXtkqLyxtsnX9yJboqn32NJpTsoo
JL0RBfohpubhaLapMTs4u2XPaBO0KkBuZFJaF2+3RN7+PZrw2XmqvILabUZ56Z5X
441pIe675UOnTHAytcdEwWiuYzIyodBW0fGqTCGRAlC5YqMGPl7ZapmMsBHGQ42J
1dEGXqF+4PjKqEDHGap3YpHjbXD+Kwh1XahQcQBALDxkvpg0ni2B5x38rZZhYx+l
2yMKEdeeVfPOxYjqpBnAgnshh/9hY0pdSrS9x/G59ALt8qHtsegAfgDOrrCPYw0e
P5daGoLlT8IP99PX7EQmz0voH/d1OXXwAgDnz1kOIlSDxcNo7S0N+RXegbIgDo8q
aGpJcbYIOeOo6wcTDRBvlINz4fOc0+EkBiaSjeEn2AKrQK4aPdm5tRKw3brkyTl/
JDOOYFwzx+GwcZmZyqODZjRzZWE6oKSol9y98gSpm+wkKv2qcGwhfK9WXSYR/4Ad
XhS6c8FJyjYDxkEwC4r8EwUL2XJa3H3nEGCCKJ3+Nk7uGYAneHZ7Kn7MgbSMwAJI
iGrSTWopqxN5SGp1fi/O1QE1whNuiupShWpiRkEZKah9+S6H35k/6U3S7shPnVxr
EOhfOWl5p2hzLArRrGatkhMScZgnSy84od7bV+qaS0icSCzSzUW7v8vPRSLiVc+b
JKioBxO/QRKswmK3o9Wz4C1laJkcj+n2stmiWNNsCIY/LLnhckBAGyVtZjc+tOT9
MUd6+bPgaRrKVDKw2Vborij7sdFeQc0pnjqcFUN4nRgKdRpSLRQsb9aFJzZXIfgB
k1ok/VvOqwpDmizXrRF2dtBESAMlhowEAisBwfSchXeMLZ7NZy98yyTgED6UUEJK
8NE9Vc1DY7+91oncvjMzzkifSaXSX3XNQqAbbyCrtAKSWvOnzlwck1+t8u/J8+Jy
tJMe74FoW+XIOOTJGyP6qC6Kq6fnRD9AFN+IXdVe17wh3VuIjXEl4JopchEYryUS
v7ZZfaXuEeGl2H6vWOjBdMdlzRPWGhbmED42VC6+Fg+fiASX6de6ImdLwP7b0JXf
j0iLE7ul9uZZQO3bodKDQS1jJYdygALVVHR0asiZGHdngcvBATgmOQR7npzLfugE
ckj8VJH+dY8lh2k6gh0Uk3P2ViTKiARBOdBAXtVyPpoT3yAiv748OxVMia4EBhz2
3PJHZiOO4MdF+I28r6XmmqLYfBddwrC0uQdyO4slLDm1MrTImJ8NCcfEwXQDb9Vc
HVfWgADJBE1PU/uAWGyKvEJP/eDhwWIFK2EOjh7OxOBOWaUIzkRjM20QeDD7qHLY
XaERHQhDKFSqK4q1Ro6TVS9/hQ79FRKQ0434SoU3NA+2IqS5ZioImgkwsPQAUzEt
pe80ZEPB26n1+B5yOjKBHRH3+8yjcvxgNXzHLnflaucfJB04WMgR+D+SYz/e2Pz/
kRsO9kWq4MGi6zIB7FOC9h/9qu92vJP2O3oWIJv3UCg5nZTqkdmZRkGhMTVCfYJ8
FVz9VvoWcTFOM9s4xJehy+ZnMeMNPuc2xJlRkqArZmhHaS099HjfPKeT9Ip6S2vp
WK4tb9F36k69CR7uCIqDNGEX+uQwXr4+kV0cXn0ntOm7F13mRsl0vKPiGidVVgKU
DzvGyK0a74VrJ21Y/Pg8+XX5B0NouGS71MbyD+L0jlOuzS3VSe9gSEKq06Zzlxzr
C2Wrc8lX+xu5nMVvK6Q9RqanVIor4geuoBpgVxEeXLuV5gpxb1PdriWEIM4/e3+C
U+E8/hALkp7R6x8OIGUBYDa4Y2H/TLOml5zrmoVj3GJbETcHpqb9dXejGYRw/dW6
8cMsLhhgT3ohShjiqIrbEqkeUvoDWmdblCg/cgRO697XuCVFNXmZ2/CgrvM96plJ
wIwkAxzBkpy7e89hdEaHjAFbNzdCwjfhH0g6btg/kYS1wVwhZdAq1Nb6Rt01hrIw
bTTLt9xsNrRKK2GtIfQOmH8YXqTHV/BKf4SePAAT4KtJx45GhQMhLgzXGT9d8o6E
8MvURiaZjr8DIHvfotTxFAwWTVCzqXRjjUTDwjod+0xiLAhXycThF9G6LdaDVSct
GUFD3bsaB5L/JTSY/AUIyoI3W21bWGg13G1ts6fxPjSaCwb+3PwYFSoJfNiDgmXU
wx/sTjpZ8qJzmG/KOpuo+BBrzK3Oj6h7XK0tEjvhj0/krD+REKSN34TFhrAlK/TQ
z06wKvnwMdCI8jOHyRECSTL63Btt5khqOEP3oVtW1qRT5X6ZyPsvfCpGePRVvz+j
dYQrx8awRJ/t+YyPa6Dl5Szgra5OkuLbWJjiHmJ1Ez7icGJvrijPJyA1XsDcfOeA
6bgtNJfE+A+BkoiSHS9B2XWFM9QiTxEqd3LO6HdK3iG2ua3MGYLMASH+avmPGoNR
om1Tz6MbTJ0vG1l58msGFYSgb1DRWDXBZ1MndyTJrcAAbukLvJgR6tcjMSVDgVie
q8wCryGwhKKGhqqh/QRnBZ+Dz22RAVDT8GwKff468GefdwgYEm3+27AW1PaIN+l8
NOVDlz+LrR8b8uNinmYbbqYJhqysxi2slxFQ8zYjdy5W4jW0+wnoiVBNZoHu7GPr
Zgq2B8mlyMKLVx2SU8AflwEef5j+8dOTBo4lfhscnWT1uK+2qDdOmynqwXAGzvGD
/bGXK4b1m8reIlLFIklaVInOWIOHdh6bS75vvzcvmGZ/k4Url5WqChmm5UeK51T/
lwMdB0qRMqY57MaTqRkCzDHCKYjGUZO1Y82KoQ8FEbw7MHz3+A3dJinbjrVCt1wb
6FC1SDgWMaFQJxxpMF776GM04fH+VXlNOZqD84l3ChuFyUYlKn5u2VDcD1O0BzD2
xMwEmBS8h+8LZrsQbES6iI3gVpALaYpmc3pn3MQWJm93LUkmCA10jHjM4/XPbfY8
MwXwi355LkOffb/vXnF+zUa31xBub/JhmEwLp0olIUrC16Q56NRkdHx/+T+l9r8u
wJyavjEzDlz1OY2z3wRcBw4TNI0YoYIy1PVJTlivDFFxgjhuI5yLg3ftu5Kvk5bI
F3P/IhLpYsy2iEER9EWD2pgRhb2LwijM6u8OH0SVik2KmINj3t/TcyIvgxzr21S/
e7+ZhqtrLYINdW+cB1r8YzH5HNDYJNKQ2lF1ibVl4cv4voG3WsFB8Jkh3Cg0eBVY
YHbUXJR3RqvBSPhNU69VbtUzFXccGVGKT/QMWAzNdQ/p8tSPYf4DbIyvWXbUstjS
1hZMlzaYbkWWJKe04Ym9YZ+kgQOMcNkmV8Z6P8ABl7IYHsX3oGutmpvz/jV7vW6F
enrWIIuwoEisjfNZhNgJvEVidurHG1fjiS7ZVKRudv4p/dIb9pWxBxD5++/h/wiK
jbP2xoqC3eMvqPOqChzLYroaOHMi7fUj87vulr4zWPKeM6vuBGx3BZCTgYUAIewO
/Frs7ZQ0KYzUoPW+2SMvS8oVumLRgfpERb+z69ztdTyQseNGCGUsdNI+Wmes6moe
lITV5LS4bCX5t4vv/UHFAA+SAWdFuhY2T3oJSBtbW/71JP8veLJE6zpYlcQ6TolY
Fk5xluiMJWc1eBXfoUhIS8lLe6gUE502S+Jh3v//hiiL0oByw2gUFRemka7q1G7E
AeUiaqb/3OpiOffY1aqK+fj7DOVcNMvb0UuZ1MNL6M/02en5OsC1SObtbBeYud75
4Mt50TNKACJeww5tjWKhrA==
`protect END_PROTECTED
