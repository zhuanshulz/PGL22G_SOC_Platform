`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kd4unR2+X9yuHxHcd+AmT13hQOg/qSfxRiPGlB0j+CR8ShPlwR0FQ5PP148dueT2
fxzOUm2YZYq2azS2I4gQMFt43yoxmbUPKan7Rc6Qd6hmQtlvGNEr81G4MFvx5BhF
62Z491ns0meVio6wXb2x5Hd8zbTTbfn69lkcEm52fxSJPs9MJpCLs/tBPXriM4pH
/Db3GSAm+vkavJ92kvB3+Ufe4Y3QMpQevFyzCxUILDzeHipgu8AaLGSrkUQFzxKu
kiiGwVt00Ksxn0Lq80+R44SIDaYiSkux+2NQnAUBoQ0NfGmfsgD0WvLA3rrwVH9p
H3tIkipfM9z5l7qmz20NP96X+M6mvoWZ+QhHEijyjEqjN+8tXiVEvRMQioW1tPsO
jMnCw/7T6Tr/LmYbggywD5DytdNxk/jkgSr7DGIhaPNHkHUUgXJImP9o06KJaGV+
qt/nCOyMOW3FvAAbxoCfX/Rmo6c93iGOLmloq8ya2wmRKkLHGE4mah+soRNdiGdK
87PgtKRq3NQJswhEhenyI/COtzLy31tEHAX2bZy7D0WRnWxPpAOmsqMKWg+eB2Zj
2hC69glnYuIU8omF4PjEtoARgpLCtKi9XqTElw335h861hQZ3T0vFtlkHqYnjD3S
yU6tcUNZsJRSFn/NF9EiFzIkX53/sh5Acmd4T0YZitMV+VxvxaG0LqK52MpO1TVq
`protect END_PROTECTED
