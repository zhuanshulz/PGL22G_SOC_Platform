`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8oDuQXsq0D5AMdXXnPGTXTMLmYNoht4DRnI3Sjl02a1CWfVFO6QtW9MdklA0kd0w
ki7lBdMLdNU7b9fezKkLkXK+hkQm/TQu5qSQBaTe0tYZNdDUvDsxhPt0JuBpx68W
46n76ZzlRnbbVux7ri0zOIU13xrZI7UYFkHvwnNzez6pqxOQla3qfqZcY6BBdiD5
HLwo+6h+lZNHGX6hA1YRUaNRWNlHmH49P3IHkAjIuAHvnRX+LW1QXw0MvdAy92a+
ItJKlblI2sHH6cnUzVpIxkHSjYM4uIoMTYrFtQTYc0MJNbiyYCMvqGAl1CEY61KS
skDtg1Q3/8a2IbDLia1o8KXefW3VivKPC/6WATex7dGGzlmhzm9Y5sfsuSWxyX5l
uSzHNoDCIknrBnO1XZKEs0YByoQyhPdsITE69OXwD2lL3ElP95RDPg4BqcrFa8yq
EzN30SY9RN01THMTk2bGl8GBFnd5wJlSVeD80FrNRMTNtm+T3bPkhhquQnQBmpuc
/6vz4e6rC5C3sxWQtcK5Vv0nV8u3kN9DacwycjjSXKDE5JDd0wXJ5UWff3FmxnQK
+ue6TWZZwD/62M3psa0FLnsopH1F115Oe9Y9Gmv9roDrbqmy07ezQbHP0ZonZ11S
4Wu0o2z8XJzaAaZBGP76Fk0+qnDq35+v58P2sbA+kS8SKNTmWMsloWW7hNsq2DnM
+NQBxUsB+LF0upslRMj39X6g3/uJmz+44UQwF22HmOqzznAAj4M8M1nVarSZ3h+x
1n3ATG3QpC5GIYI7piHZ2TUj2YQsU2KTQ3xBgneMudjN5oTvRTtaUKK4woXZuaNj
QBe/qDGDO+WGSeCc7L2hQH32WJZyDXjl3CnaXzuwYWLpALb3u/rulUSUs1SxoMma
5HVNESvEo/5upqAAucwhj+hbaKhCkUIAFyLtNlM/AlSEuSKLgNMgSiHMufJOL1Cc
qUaxapvJpvWVcaNBog4xwTWpaC9BekcOz9F81nzjpKKy889SolXRFO88EPRRHcAu
jGcCuM48wy/eZQiBf4e2eR6ylg2abfoGbQKcEHJDK325qDOrGH4f2tuuD8umEU1p
0QHDIDHIXpk5XFFsBXR7Iks+5Z/4/5dUyCYYKrB2nN3McQcMerIjSh8ZXD/1r/2E
bHH22+xbFkIJVziPKPAcxtqYZwLer0FJw5vHLkPKh4ePbNf4qCAj1YugvqNEn+Dd
BZMy0p8rKPVPmRkGVj7ABUlkPVxM8hteWl1ve14T7PoJYL+o8w1FUNGWaVJsWd69
ZFE8Rlaam5xULK2ek2Xpk1CXN4cTGEhH1kxVLAVZkshQHwPcwJlNIUl8RUi2b94T
aFZH0o91uegGn/J1I7PyOYVldlxicq+h5A7HmTkGF1krFIYgvwA8qTa1bsh4FeE7
34gL3cqF+6t4eQ1DUgdfnVMagOBMIobXNaAjv6ggCMUXsAZQDjE9Zp4C4zXXloxj
QoM4jSG2A+myrsJFJq5UXfpw9Ftzibn+BhngqoncBS+R83bMDLFg6l8w6uhkl5+4
nfjiBEQEbN7Bm9ba18ajuCa1hpSNcAq5N/STGcnfVxYwKdU7v+LwlgF/5sTQIupM
Ky/ctQVLM9JZdJqqNPuVa6vSvFRfiZBQASKx5erxs3Cag8B3hh4mWgz40CpqNZI8
6/JJCT3gYZ2IVMKARYN+wmTPrOQ6eTJNskuXQeIDA/rNBv8xOjtnERbLTDpLJVaV
LKiNzO3abLbxH0MS2icAy+/QDW3dOJIpiYziXPXMkCERHo14k+aXEk50WWE68rEO
ZheukDYGYDaD/kl+dBK+flooHL6MqnhqPgfrKiukLRToIeBL+4/uFf+MX624ujc0
AhE487T2/4JwFiA4exc1jcUV3DFbq5+Ixd5iP1NGeM+9j/OJwZoJo8/WR+TANcru
A5Y2R0+SXjf3fpCmAI9lc2YDjHxRcbGAurehXUI28ZvTJB2ofXgiatQ3G4b/TmZA
jVWkA+4nWVl7ZGGpZTRZYrtCsFsaKTZNdr8BC/8qFZuYcKbSjEulIH2qxOgDvkWv
Oswc1dT3jY3cleUwMTPaZ+YSkeljMHyyJ61H79nhHV4n/UgPJ/iVCF3nBLReFNCh
BA2pSucX9YpPzxc2toOZcJjIOUj0JlX+tEeFTJmbRp2wMLxRzpbP4+ATo2/6NOl8
xw5HAPYFWW7oXW4cliBUuJLQLEvEQWGo+mwXS9tauWJUMQS5LMg0CENLT0StmoDe
H0W3JWghUCBOAC8WV+l4fBf8qTH++TcI+6fbwTTps2I0kxJMGENdX9/DtQwe/f9Z
fLNLXPiObe2VXrN+bPJ5dWQQs0Ccsllp30IGca8pP7pGy0X9wFbIarFIBTYjIPZz
YCKAg9X6J8cCN3ZIg49xxbMsaFdugiacOIYJ6gMfuBV7HzRo6KkutxQrz4oVRrXq
6i4xSvgTEgQ/Camx8PY8PP3D+WbixDJdd/YAJMSwDDxbAsfMDXwyzyR7+i2huoMl
7JIv2SIJLyQnuaFabo802xJG5VOxmWWcvLozADhSjqLick0hKvPB26vMnL7KsqCL
YZcWTqTgdmrqkQSWKhWsB17jAXzeE4YU6ZgmXI5X+glEgfIRzLeJg4d1xs0Vqj3M
TpSqK3/UkvFqhmJkE8X2t1Afehb/HHtc4oEZW5fsWXnrHHJjSMyjxoeKDxvUj5n0
wRYgxGZtLVHPCCigCelqCsNFZp3uvnBjjcDYA6Z4h9Lr5vxtscQlhlyG/rUkNjtn
`protect END_PROTECTED
