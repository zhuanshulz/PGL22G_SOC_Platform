`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPCPjcPuMv8ZorG+Am+abxQb+vg4A54P/Rb6YeJr/dbJ6tsfboD0w7s8PVPqZ+Mi
CEkuBs52z2NzyCko1Qxi9bIWG38yumYkVCFYv25bleudwn7pk/cA05wk1qUn2VcW
6qZX5LsvUPjik1JcicNuJ3IZ8jT/BrVxmQM3YXYnWXt8RqdQqhzwAfgA63Cteyyk
HBuUOfuGbbS3k+LdxelSgb2bObNPsuPextlMBVUuReoZ6uxtGyfCxtI+trh2ZP9Q
v2FK9eSEF2PU48m+t3ubBrBfoDPi9E6S/CWm+Rib8fYAfVKCSml0+ma/7wTpJ/nY
dVUq9Z8pJ2vin+HsmJBF5bk9ZfznXQjz6uLoyeQnxZ8LGfatruoI8299HfmnQ9IG
EBC25dmhqh5HqjsyxtP09A==
`protect END_PROTECTED
