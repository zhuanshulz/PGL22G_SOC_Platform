`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90lmMfGFsBA1i6Yi5/24687NksQiyeViKXDL/KJnp4gpsVF+dOnzFpiI2wcvsPPq
U0ILA/DUg+tlgnju5tv8/QZevzNlY5ufLP7TLO1qskeZiuXMvNLPiR8dHRDlwIfS
15xgRggcjhnpNUa9Ota6Jj2HMKcLzfaM2yPAfOH2sgIbfwRPJj3kZNCaGLr1g1MF
hM4E2/Jttq9pDXVedHbvPC0rlWradQ7EZW5NQs2iZj1qpq6pyKDrz+C85/8/3wpC
osQWmpSbi9tqbndfdHovqJz75Dps7nh5qCdgj0ONJzEXjGfQEdo8MYl3K12xyqeC
AEza8YLRZCmtFefFQCrvHimU7vZot+QB8TEGk4qTPZPUkor9kZ6T9ZWWwc5QxcML
Xk+SD9iRX853IrXZ8QfAtGdjW/ztpIZ5Rjns6rJ/JxkeH5mzIpHoIjyKc39225cp
Qvc2o5eOFVC6FJUHgtCRFZ8yjYr3Q5dOyxxn24650Q3Vu6JKaJ70t6Dj0mOgJaEj
ywB+nx2TX/ncv+7iT+RJ6FzS1dmyRUrf+4idyBZhwxjmkWDTAg7v5UeXUDvOFE4h
mkt9Pno05G/9BeyQl4doZGDD52gHW0UK3QKkcg2q2v07ftR9F83xQaFTMuGf7gle
8yWhNo5B1Jidr3+IkdpPeW3W2TBE/vGAQiAa8FQqLDPCcVRSuOmCbLVo4VvXs5du
pMCaxrZIhCsBnLgvMEDQqgvV1sfUFG7H4jNjs7k0CqkNuBsNpkhsrh6MzrnuMqs9
7Ep+KLpxn8IcvOfM3IYbU7bKz3TM5XMh8lw8OOwJyF/ck9l9DGZfoctB/5Ekuahm
L6H3SAgsMstOdOlV+Vz+fkm7QC76fucLlytpU+KXqPih+J6oaKavnl0/e0z9/wVH
0ajy02f0r1hB+kTs3OwiBzAJH+2b2VZo9ywbDR7NpuZBdJ1MV3oY/61o6vyFB0G+
y1TbJSdT1NIbl6kxb8wBbgSEXtZI23tnThElaPLUY+G+nC+sc28t3tfJCu6whgqV
w9L4X58O6sVwvfrmSaKLgHxzza9UknsR7UiTLT4VGN7RujYg26fbqCDfRyJRN6uK
pFIeSgOMyz+r30E13UvLwAQuGJYAjvf9skBMi9V9GYB6XAoK87L2dTTyeXb5/AwS
j53+vmyEyI+pg40t368hOj8JA5qcOCYo/ssUHww7ss40fvnHIKwwsDO5v56k682y
pQPhphXPDiZS+HHZui1MXTUKL6we9iVmpL5BCH7HcEbr07aZxzi+gscO98Gvhol9
DrtzlX2OGIkUjvBQZUysgtMHk0EmpOkyfr2lPUjel3Q4UOVVarJaO4CPB6jGBu0H
o93cMpzy7I7D8TOHXZNWV/DPucxMCucaNm9uVN2v4plXH2Z/x7B0aA2NJgYIQdEy
q5x3qKip7ZOOOtsu+5zrZfi0cQlxUFNF1XvfG955Wt4oWvmPXomvp/rmiStnoe5X
3mzJWOEkueicoasIX8xZIzKbS4h+c/LLqO+ElYe1IrOG0XdejLDsh9z0TkzjgOv3
BWwJ1lrDZ8v8rLZqe6ep5VsLzz/+jutFifSC7QH3W31ySo2bVndzIrjlhTi2o37E
y79+wYEmA+QDSeZfX4w3SDrhlEjSTC6FC24wtz5tdrUtFEDkyVroS9581Mq+QSY1
lanyz/5omIHsvnfoJXFp9ZrEmRMitYNiCufcuB9K9y2OE4IYcmONfzJTGUAz0vLx
zaF/fQyTOWt69GxVN8igI6aDxzMahyODJjekJ9ngYHtBYOO5XWCdJWQF5vaPAv4k
1Eh710trKw16DMK0kkapr2H+ICY99Zi1C19AoIUsgD806boG5H+Z0B1v5XX3H8rL
5IvJfXJi7VBUHZf2UuhAaa1o0LvHlTPw2LDo74gv0Cp/6pvj/SwJjRxTboT2vyRC
Dk4rsVy1+iLNOtd3ATBKx9mKNCZzRIRxKT0apatndW7S/rjt8Q/+WxHuAVgCjYmD
ua0/c73VkOXag/veIGR/k/xVsS3Olfqm40NZSWvy6iQTtu8s2DBq+7xUKT9Db6Gn
4RIQ/7A2cv0e0h1d8U6wJPscu7/N5kSjLOsEGpqE9HugdJ9u6mBNxhoWiTCC07v2
IhJ50kuYDUL/eFC4SWSY3NkrKy27YC8bButWCWTcRxKYw6wZne0X7Hd5K7Vxg7mX
5Gj5RKs+jJ0HeKj2dOfhi1ZjAAT5NwufGZ/M3GUh2wCViA823e+66gJDe9lkcUcQ
IuaYpwVaog8ezIZyMpba6OXZZB4p+TYd7LT4qCsZTqiNXEQi6DoOPtENL+Cz/N3C
3afMc6i9DPgaIzMAFz4QTAKqEj/mm46MRWQ3vRNCcPl8FcRrCGHgwlGa0iF3rLrf
QI246INubMJDa7OT89YQqJ+e/k5/EPDuCYVOPmp5gIBUJf1W1NBAOIsInDkwvOcq
pYtnDt+DyWFv7T8wX3pgZmhd5KMU95luy4JuCaErCiH8HP6GoQRBqIMoAE6n1ZIR
lRhuMLO2nWk0zqnVdZGGgh7jcZuHpQio9o7XpOMLdPXNL5MMs8RhYbJ1GtyHXrYd
I68VjOaEpKKZc3cAxcwrIxEmWJwDMVAh2Zq8Oc+xZ5dIA7ohk45PCt/UvNsaCwWD
RHfjrKKcxCqyU5kutzX0+ZP2AVOTI/xI+1W6Wnun0F+nve5shsakyl/4GhmybwAd
vGsWQtVzf9XhgSMhVqN8Soad32W4iHIGQ04WmrrVda9wpwdkG5Dx7CnlGoSoGTDn
jS8R9vXB/4WNulpYLMIH9dG/w51nCMkk4yW8ha8h17V7f1CzIPU858FQf5mILvIt
TaRHKa5UdPoeIAIDE7kNW79QWW1RiUwcLPhMfMLvhPFgH2Fjo5s6/d/+tkP0/8Il
bq1IM+L84/7lAnJvIzHVgWAwsvkpB1sOU5hq3nZWR5iD5vEAdJpIYTKBVkw7azLd
rtotbAwldIZ0iNMqXpY4MbipfTS297f5r7tig0H7NLxXh/thjam3XZXkhegHcTmi
zclPOF6mbgDSNYxQw9Ew7e6Y90zRatbopnK3ozzzwzhMIZAeZJZRSCWUjGNUuaS5
+QPjqSkwXiwIHX5Kc5yPyxhs8mJM9RU9ViI0YJ4Dp/pRT8PQrmZ3yBGqjrV3+G7O
LOfDuhpV6ct8f0NZYsrJWInyZhKQ5tpbGhVuTFMgZvo5xGDOYfHltNN8U3H3Zbzf
cHwY+q/LkI17WQ74BLHmcE7yQU1CO8eXDOFTDW5cIKnVeBbcDYlj9NudAd6f2roG
wf6YGysY/g97YWjo2bZ38QwAL8Jtwx4iY+EZudpYFVh2lEFD8IvInBO1JtknQwfU
mQA/NNWJiqyHMAXHnF4LkyLOW4ehKemS9nb3Kyct4EnH5UmEVfsjAn8fxYqY3sI5
OwkUTYpT+j7H35ETsflYVRCnb0VzunZkV1UHHFrvjykD+K2SShbJvZBuctMC3LxW
4vHkvsTYrROmg+7q8c9BUm0Fq5QoMhRNauZ/CUvOhaX3+eNIxlbg7TuEfaAqJaAl
oFB/YCD4lqn2fOwWwJqFc7Upcz17rO71vR6PrT8dzABfrmJ1GUJLH2Nej8Ro7uUG
y49984wlxILDvcaagxoQdAv4oXs1QqH6X15ut3tFYiljRTlXDFftRVddIbQtPTj/
IvPOu8gj1LtKJDnVoSyZYe6hNUXRqY+vClUIZhtWKzxq14g8GgPCxJ6VA8dJM41N
Zl+1sAilnn8a98Sw+Y+XpDq8ASCe0QmbFOEQylVTSCi7469HuZp/Qbzn4EWhfkqB
GL2c1ZxDZreMWz4ThqN1rVLRQkSuDLM3o2EKunAAeZnAj1Z1HwzzuJjv5QE/g2ci
B8XBFCgNCx4tJ36zXGbiK8G8Jzvcm/wjwrRRWT/SRNFRqWtWA9aa0dEiPFP4fD4L
CKXNGy1SCVjojUZB/PW/fOuP4Gf+pZtqnDf0SzVnB80EeP0WxAxei++577iUyuXd
HSoG6nceOmuTJcB8s6c1qKtwWozP7/69jvmttLj1WqBP+p/dvt45MXa5kOfOlqaZ
n8GRYyJFrPyM7ialY2LyVDIzzCAzZ25k80iIMBd1jFH8mO/zVDLKqlUUHWW9i9kY
qhNlODhCTSztWp9TG247zcn/YeklgDxa2M2Lx0R04wDzgf6KqfQiXwahPh/h6S1h
+GGL3P/5DyayoXOeAB1kkrULez7AgXaFllElKnQX14tqiYJreSvxykm0DD6ncIng
tWj66jwSkFjkb6ZUrukYuFNFEimZSf6zXF18LtffpO1n5nE20eUOopg3wSDYs4o+
e7LgBNDBnDFzy7QTsLJV1Yh3LPRlUV6KexLk4Oh7zR86l6ReQYbSORzb2YvuAx1W
1LAP14t31WyppDq+EQdTjX2WhHKoY+docNIgimNhvki0BJ6Mm7t9WkyarBD4qppM
ENyZrY6V8nCb6RzIW668Uf871mha5/NuXQUjZ7t/dQF1MAWqBmaDXumG3AJ+DnSv
MYR0yKCf2SWUtPRqKVUmw2vIYIRnvv1NAntMRuUK8GNVY1ABTcl/10RqHZDwf7wL
Y1MZ4lVbUQ1Xr+IKYq8qj5+pIRj1oal0EuaSMqGEdXo+N45ZP8ePs0HpQsEX89Mu
SDYFQgPQc51vFOWMFBmmIZHvM/dwgaHHfKTGM0HfbwxdvWvBqlJwz2Tfsjj3qbN4
p4yQsaUSVCt5vn4F9h0wPzmnA36JB37ndEsjpMk5NzkdgORt0S1fSIBVIpC1GLR1
LHjKNCVGdgDkvYBNdwHaOLTHTTrgnS6lWLlqN0O/+swFFZlU80vf4hHbFrZMEPd4
x6wWFxXZrYuhY1jkmkgp4KPp0/i1nEgIv8jV9qlQXC7zNlv81KjFaTheTQFeL49o
gMUzqFhizhfkB22IyK8Yn4xa2mvJc8BkMAvDZQ+dlf4oUOVsINAVMBObysiZaURD
saIufgvRpSt62mf3fadL7lDkBTFfP0BeeG7tjArSnwte5zwfHXmkMEBpaGKjrUYv
4VfdRLZSlRxd6FftCsiFqiSoZKuoL8W7IS6V6/jvM71K76ZJ6wBElX5uKg5RRJsU
+U9zc0zscs99QDQpVkt0pQepXrH7c6KCUlCFWwMVA0yvXvOSCLrF/231kkiJ9fQh
IRkGBhancQHE5tBc4BnMl7fPCVMwu1MGMdAtZ5JcUsQs1egp8OrR5c5rEtPR55I6
/qoQJMI7eDGr3TidMlboPeg1TYFX41Tuky5qP7wTnYkHI9fXxbhxTkhyiIRMuo9W
0hM0M+jxByH9PYVRurhX9hNXsTzMftyTrVTvp0Olfcb2PeAQjl96E7X8e+3NilS3
7wGQyL9W5RqaUnP0CSMFsWKvNEqgdE9aWMJBpKGvxdEBaRFi9rP6wQmF5pCNMEq9
OPof86V141Ck/W/YqmLObwV/1Q9R+JjfDxjsziaNyRCREgsmIJC5D+VXG0IPnWG9
hroDNqyLHbKOvHStcs4NMLWkVzy/sVA9yIswPsoWcvkSpwog6TV14VFRDgFPgUL+
87T3UBFRTDOELTREhAlHXSv/1WB+UKEwgY2ySQiHokgqbu2bPNR62/x6UE2bF2ka
+lWAvinuiLnx0FhHdTuNMrRyLLHH8oVaim+gux6R0ojgPpO/NXPH4rJNXngEtavZ
0YomSVwDKseVzYOnIM91Wb+jJxYXj1qXtW3Iu/mbk7IqF4eKQjYdiAQgnI9EDCPa
6TGnhp5CZpc7u1HGZe5Itm5b6xjGJEHIA2OsNAOOSqP7oFHK7ZJdYe3ekWTQ3V6/
dPXy3sh+17yC9pgZdgKAEGRslC6Z8FURJmye1rnjChEtZ8sbrEKlpkQ5G9wXEx7c
zwbR9B0lEZXdZHMK91V/FHZUv4Ig1XouRw1/UWKKA+6fsA2GF/00X+wC07a74V+m
KnS97dmt3VolKPLkaazwjOjVCHouCqmhELqhK65z83XQvPckEfjfRiPeoeb4m+UB
D6TP/ven4uW08uVzSH5/X5RBeOo692H/Gr6h53Zm+jE35L7tu3incs3E1/TJ+pzA
JlZRt2mNjm86BZxqyCw9xUXWe9tbgW1FKS5G2hKxL4MtA1U6RwcAII3hLcs6VB+5
BSiU8qoJveA36yl3dg9BFy2UXVRdMDwwgTxfqRdysLH8gVI2E+a+YXV61Lb6A+Cs
9u+YvXnZ9NCwEgk29yqIeSRLoG2541GMfJuo4PxZBgY2wszq+4gsNoVmex2Tky/9
60IZdT5gLmaV3woduHqD+oNjC76B3qSYmEFleoPbpGYXnFyfitarA3NsA48BkfMO
x1O/yq7ehZHrefxETlM+pVFXBL2xYDvzQPEv5uOjd0Z8VlhaNjf+lUKJhEmB9uTm
pG/HQRcYKgiXPdg48szwmjnV+UrhWDJRrzlhcpC++K3Dc7t5jbcXgE7zzLopdgaN
0mfi87Ky8iqP6W4rQ35mMRnOMHCmypVM0bOR5unzETl3Mz9uMws5fD1WU0iX30SA
iYZ4qbDiTyqDV1FoI48sOFJj2/7koQ408RESdc4pByYGcZvO6/R4ZI+eVpY1P+Kj
x0yZc8F9Jpbspz14niG1qiUbhaPduiUAtTJBMzEVYG6voW/CCW8Bn9yRVrkIMMqX
OK6DL5igqLREMcY26yUJHbWGhLDeaGSTRU+GuM3f02uaA9DxjmE9kkob6Jnej3Z8
P/ACvMUg4VMzBxBO2kEi5u7yVA1bbxctIkKmhhrO9f+fzdEy2hhn46hJ7kqhOvXA
3sL3kdAAztRboU4Qncb5K4OW9jCdgPWz8yd18dFoQL6KpmTI0o32asLRF4jJiOni
hX6l3LrwH6ETbMomAlkRan6whkI1eroDB6WlGxl9ljpBJrQ8ET2+FLm8Kh+6UELW
PRjWe5jOgdNTmHM5Y5VZzTOo6WUTmWqaZ7O7XgmRcVtPFTKZl2DDggms1S6O89XY
G3qzJ+OJaK1o2qfSd6zsfYHvsR75LfVYriJsFTbmvcKfcVokLzq4bTLfQxtw6+E/
l2Kmp+6liuFFCEAbdV9RG3mvOqpc9DssQx2NU5C5eH5LciLgJUMPvdLjcYR9GxyZ
hn8X5JByBqCyJN9WF4r60LiivrAotCwShaGf5nqJ5ix7WxGFAULQxcRx6pxzByXb
1mn/9ITsgulNvQonH8MAo1ki4Qn2usf+cVfqSjTevJvFh8tu/hzaoxmpxDcmLs9I
kiPUALj0s2AV3mgKtqaFGf0Ah6i/W+gLrpYZOibIaoLwZb6727120A+jEYIlSGAT
RbtiZTh9q4CGPKSsPbAJGjNxfK2vSf90rrIzV5WJxJLFO1D+aABlQUcHNe3ytylF
Gpjs9u2JDXY4HqaojlH7DxMzyXoOuiBnGkqmvZVIo+eYZ45IBXNB/a9p1LZ+91wC
ycOmuItkq/ptsqJK6EpDWNb9dRAOsCtmEgPdA9D7VcLPaOcKFZ0y/wu7XE+HQwew
n2lck0qbXJZhMC9btzmtg4q/2mqspQJQX9yfeE0vY+pNRyBESzH6hU5GO0oNmV6m
VTE8AgLEPFxpdA4L4c8CT+9Ru2Idkq1FDqgPhC0Z7u7FPZzcHDDmt4lR8EInAkx5
slYA8wnrfdwpidLpeUfz9FVKBnfKiRvA+MnlWGrj8ADAFr3abz81t8rAjvHOYmBg
ZNlrE/D3VKGGuAb/Usr1sjaBpe8r5I0tZpN36AVeYq+lSh5Z78xdq3grQcXTQ7Ii
yNq2Ff8XmM9vER/lbmWiwW0fhfgPlY9/7H32a5zAWhMS9hr08e4vzht0fvi4KqlT
5v0YvVjEbrhP6noqYnkJtTSS3RtNe1sUTgnu2bvk58Z6aEsG/W51Dz/yLi4/gcAw
BZqj4n2z5Zo3U853TbMVNGpQVr2WqIogjA3+g6cAaI7iZAzb2GvNscDmroP0oXBZ
UbdlaV3JQZihOPSocItyB79Jn22bWoqhutFBN8CDXXKdma4p6aZaHtodceQe0E1u
3qVj64z5haah7s+drBF+gBtXS9mJuIJfv5UHSzq+FQHGRTbdTAUs89EIQoXB5bdx
Oz7U3vGB8ailro4YdLJaFKn9PLR0lId6wsKg6K+wFeNLt9HQM//yGEBP4pklDBxt
Q+86M7twaWMeYGiScEscCcIycw5hEn97CuyKXcr68fTMQkhZdWclIvxnN6WJLdY6
85pPffPnABHoE7Y1Pn5LmIrZZnqXXlN6KLbBQFBVPmMXSl2qGG9yz0Dw45xzouHX
I8YfjALIrsngOCtKmrYY1wv0ATBnq0F2WAoHVqo6ZhwPpnG2aRunwHyi2NFi/5eT
h7hnva2qTetIqDTUqRN2znNfT/Re3fTbiat8LkfBCDs9z8aqO6x5FJckH4URaaj+
lfASGxm1yfpUxpyYGyW91Sd5qyXKlDEqw53TqCpbENI75Gbg2oHaENSidmJ0K5Es
BZtjRFDGug4IOmD8vs9cblby+SgpL92miKOdZ49L9Ehg/kqUuDr9APuvQHtMpplI
mhoHdn8GAB25qdfGR8Me3V16WfcPBp0RMfqEPynOrW7t3aMvfTcRLQN5+xfIlVgW
GnPqUONzLmAOohZ+UkKGTYdl3vCt5XHE1djRB1gPHY0HamxS9sjHgRuGLTv1Dlql
jygnPgP+fmZLjqXSUO5dzhI0/aHCBYwumcCaLmMzFPtHiO1t+DthxWbgsr+M5CPV
Y+cXHQZB2eT7F2/fLKUFGdNFz+ULIjY4Hn9nifZFllx2DRB1AVIibNKHIvnD/FAR
7rj/EGgjzT8fewk0OahtVOOZ6uZubTNVgVjpkW+9ypYovjgIbSz0c6+Ggy21VlRz
suMYzYKjhjumZGOYj4nGAvFZSyQVpopYEBm2hMBJ8jey/PdIKVWb5GNf5sJuntXp
62H7cviHGwQGW7xg9hKoHEz8IoePPr87JSNyGv8WFGQgNn0l+CJTtk8wNJYm8U/L
DeEFvnjwTGUrgoC2tv75XUKgOgdq33e7r51l19T63NkxxyP7tYlxvoWzk4h3wKRV
K2AeikQ+GByfgGE9iip084nIkx4nxzvoupNzXumZ9hnKSP1tmjMH8nOKrEV+Nlct
CR6qhr124KBauMeSqaAET9iWTICxamjGjxU1PQyZkN8hNbfI5Zn9nG0k1E2AYoiG
LXR7KrcthvK32nKrK6jAmWbVo41bxw/7IGmk+8y5sZP9/g2DN8XP7kJUlSTQ1wkr
FtLTdDp3n2FmwBIz4+9cbbU6GT6E0YzcR99drKiRhg7wU5z3GjfkuZh2dvIEHHOh
PJ338mtalvf+UhyBvDpUSNPzxnnutJwpRXc0F6km3gBOuutauc72LQvr7bA9GcHm
xJAAiEdENLV5Si0EN2CVdXyz99XJKooP7WbcGexzT5th2cDs161Puchl9ctsoAKS
0FPLRinsuTHasMTLGbLNKmdUKr/VSmA/ZdMgqzFCVANW7SH6lTjiLI9X+fpGqX6H
HxEdHqsD2QhnsZQIHlBF+1PoUa4b+2A5R242oWEsRAhe6HTp6Hpk83jU07WuD17R
TvFuDBj61NZGXvl9u+YGuGh9cvOvIN/KQXEnJlOkLXJmpQanoz/jA4WiBn7n0Fo2
O6G/3+pRWBIF4Mcg4cRz3Pd829xi42KDlGZaWc8BBqIxvfETETKjQn3oYoZ7GB2+
uvh6TKFBAxYI38vGtIiDDIeretFR5zBeg4IhFlb3xay8tY60Kt2Drsw8hlZNlSQY
ooGzlOywJH4nhsqxQgeX6MrB1/e3UVU7GLbDdtX79OLSqOJhJmQ1BU3Eqvlp7Rom
/QzOif3oeUABfDJIbk1Kmn+WdpUJ1WGcn9lv8PcFmvzMXIATo6Ofsd2RLttHliVV
Nq1yjMIIUvpf470CxRpBKW+niJls5jwFGitxrNvKwm5o9/zr6BcRP2Hb41rzwQzN
kXEgWsk4ed1qKAT6eZ4f/AfEICUo3Lat/G/l4YPhZmrh9gM6Lm+yfuhsViaga00b
PzWkhKFHK+LVgMzVDtieZQmB4DYJwKvZjESztT4zBnSySGz31nneOpUeioJeFtXL
D8Cmu/Z+cvx1U+IsYrmG8UBKmxtvKDf0YTVyUpIK0ltgqvMp+Fapu6wGkPeWppj0
zALUngAUBTFssjDnVjtHRbuNvU0eShqZ2ZrNk5BYWAHmhSgMYfjuXrgPtnb/DjrE
3YVnYgD/QjGNZZB/crI9PISNdINhOUoSq33+aT+5O06i7awm6HesR/3dgO16ZnTf
BQGTwDDco7UwZ4wS8427TxdmzjTtBE+H7uC93JwE5Hx/5e60KGpBdOWI5roltyLH
+oKzw/nkt0Q9nvUg3NYUmrlqwiDtNXggsZAMuD+7W79xMt8cOmj/mQ69Zk1Xh/5V
isJb7F9jDPKjy7yo4KTSGF5+D1PdZGhVAGXMqgYUo0CAWeW1C/r7BFlpWGcrFgce
EAkbIdtlEzRUoAu39HkB/gJF5RlDq4xlYOsenbZU4i23I+UKVLYtZonxJZqTkvFf
G/O3mDMq90xDm0LV/590pjDwTfrvjOt4+IcFzSlKQ2J4uReEiDU0sNcCQxeTqN93
U7SJiPs28bPgqO9p3HCAMhQaAU34bPWmAS+WlfLuuja+xbm2YzEILF2KCMAaX+V8
5p0hp9QWHIGmNLj91Exd6A8K1Tt4ZoPNID3vZmYizMRfl7AHuqFtn4iLVtbO4Phk
+Sq+pYmI0eCMi+TyFe/3OOlQEmYksoZjhmJ2n35ZPAchIeB49T5sExKn08Iz55pL
BGpDwtAurG7Z+0+KYZZaQ5VGHPfxfE8EHHaO8aKtA6iClnDR1T3Wu0t1///vKGFf
8mZ6kyF4jWrgDWUAKEBpSfF6t0YUbRYQE4f2u06V0pKPk9K+4ca4lrAUUbQpuaFQ
sP+ItxdvYtAez7bF91f79mKgx/i9m6LiIlaEBmmHKV1n8LZr3qdAtgTenIsZNIrd
NWnBQ3eueVyRCbTb/OQnt1D6zEXdtvCDPoBnG5mdPiMcz9HfYDVRpTmWOw1CweEN
HCZImBXGm4M9mA5J0uqHfWUbpjlcgf0IeGMthXWqY0FOv4qF20y6/SZcxOe9h88z
S2WveiD8AIyUdyzYZi7JxIjSreQyT+2OSKR2nJ0riiLx5w4tBzeZGGb9ARvXfITX
kwYlOGof+OOLXZHwQ//oF27jXibFQaB05EzXa1y64Ymv4u7fVMiINjbdxVe5KSzN
i+fIlczJNgDmRlZEhpL1lYAg/HG2kf4fZP00PTsClbL3f9vsLoJySN0hpoPQMv0o
4FtxfM+4/EmGUwV5iinVZ4XiL2Yyp6kKH4S1j1tBL8HBK1yUpAhSZavocxeSyxUW
Dc6ToJcv99vEh1JmQ+O9NWtZs6PBKAaOZIhzwwc3ec6W1pyWKuLT9/nzICgt0rle
jdGw6qPNcFb5PbSDAWY0AcnK0YWuvp9YWvNGd4vKiivf5PpRBXPbynYhxVCvP9Fd
TPy+CReTEQMRBAeEUPSrrkvD0uIkOzjKNV7SgzhqAROliWNhhPIpvhStr7EKb3S9
NVcY2Ie3YZzCYm9bq3Ual0PNDvHn7jWuIGRz0RdgzywpJH9XO6Hm7DWJoQd0Lfob
ZRod7QSDC3yj4S/M6frtoEmi+AKp3x7W6drwDTX50iyPWaYiz1Q9Dq0t4pnyql44
W17W9MY2KvEbMn/1BhrnBDTfzP/hva5wn3VUJ9AgIvqBRX2kIKODR3NhXcUfY3ts
Uaq2npmNuTs0fYtgTBDVFbzx/qz9TUKaru14jhSUzHx3pANUbePWisW8QjsNgqQq
vQC+AVcGt7Y9yl4v79VqPZx/txAkkc+bTR1PQmp4Lhc2whDfQFX2Yrdmi3pNMzza
b9wmO28CWeAD3qKXfeXm5/RgH9RWe8EpQIJ3HInu9kX4rdVjeCL0T/7i1icHuYY2
Rq0oPymeKYnfGS1kBG7JQFp26u723PefUCI4ScKyj5XHvB89TavjdKaDy6HTcMcE
ZDrMu3ZSEKYtIvYjqVMhT3eoZb4op4nwDUsWLda21ZMbNQHxUBOZQDjO9+erKb4+
g+aiMg7mnV2rP+NnK4gt0wk+tny9ioBxwH7Rb1kZ1ZltJDZbj8VBN8DNoYzWI6k2
N158EaOJMKI08fVvqZrTvXm9BAFA+fSQOy4H2aqLEX25dTVgIVeOzI1fg7xGd8dI
tM/1GSKSrG+cE2AnghauEXVpjnliDB5Shpiq3r509c9L34dii4LU5g7ejD5xD3g/
vKdzjmSwhU5GoEfwl3GeQ39CcuDT6SkgprbsKxBEu0Lr60wUNtRAQRD2m4i2Xysu
ublcXZ5NdjEyUak9FInGas+HWtIwaOsJwucivH3E08wK2uz82tVZ3UoghDjZewiZ
ih9qKw5nWkJX2OT3vuQdvnOXXa1GOrD7LuwsY74BI/JArv2qWAg0sLlCrGIVOteZ
XKCBeCqOnFh0rcoDUdmJuH9gkBj2d7NKzFITFeW/Y3T313t7fqSSjZgkS6LHI9iq
zZLiwBWEBoJH9W9l5WDRIDjZ+lKFWuOkCqctEhdnHoHQBQrkRc8pEfKXXHDm0mZh
yVLPsgtVu6s9ELpdXDMsq46BPA1qWbOKjLPM4cqMYq206ZmXwlJizi8g9OSAY+/X
uiLBUFjejoHgpjt+LtSENpORmA8IdL+6n6p4NfamwoRaV2q7EOnoLBgv1fnQGzYu
5KrEbMn8D6RF/U+VFUd6eCgSdhtNnRZkZoGcVy6wfb+fR4rNLyQOHCOeFXvYpnu8
E7e0zoYWno9k21HHYWdFlSimVdY+k2wEM5+h6sk2l19d0O3QzpWg3SRLUjJrmXgD
6NFmGL4VON+iP98ah3liCL+1+3gH0QlrrVwdMEPV0v8bWwe62f8yt+I+c69i6MX2
XWBHxp8ZnB2UqYs85gwVaED2LDslsghcP7AFMUUtJ+s38WnLz9LKFJJNPH6SuFNy
8Z5N9D7vKwNaRUOnWxIyj10XlYEU5yTgza0RwiIkgkRKpeEAPxZA2HWtdDyGjXq6
gR9DFrrFSi1lGpmfxGwXFIg9terkW9afjKAwFA2da7s4fLARRPOUjzXOOuigWIV9
prEA/pQ9z7LmT/eFE9tdlp4VSj7XoE1wL8xwfElMlxtPpSbSx/hoKt1szE9wgp+Q
EMcTqJ2bq8pcZ7LQ+n+z2Lgy8X1JD4FByTgrDl0Q+pIBH/Aq+9+GKjV0cFnTYa3B
Tz8fb9J2Q6SubrYUlw8c8rH9h2CUJbLO4CF1SryLbF8h/MjECJz8oSuf7X/o5VY1
+OjpagPjW42cV0gHnv8eqcgwdb3Fh5F/U0hgazUu8LOnR8MiCxziOaE/gIAQQl/r
LAHXMv1MrMxksPvea1DOhgwKzptBqHatccA3kF0ijG9C9n8TOHnewF9uiba9s+s4
eB2ers3QbUGFGzbuhy/AjB5Xxu8D1kuEwDST7YbOLUMses5XXt/01WL1ICneQcEK
NRTcJyRLK5Cv7meqAl2yaCQBbH7SSOwKntgbpWX+1xeW57L3gC15tDh/MIckv9uj
ar8Cut/ez2ckpyoLcuKdDDXhCNMTEmHzCyhOTaRwekqTcXLMIryn9XJUSjADaBNT
gjMYYJ1IC94EOWeb34oCE8FTvGpWgVAnn6zTjure5QxHIVWhEh6RmEoGDqiJkZa4
Tr9lSL7ktTmXAtGw+Bf/9NY1it8F16imMxKBILUZ4dekQYEthslrYLx4wNOSb8ED
z25+AO17xtIGXYL16vCYFMXwQ6VnmnavLnScjjhkBWTXZDEhhngcYpUXID6YYwti
nqNhx5LyUm0jBEv3FEXjF59jok1klY93uv2y6wlo8qSvHg2v2wRfES3o+Jo0xwjm
wn8w6m34Ku4m88R7RkIvIIdZBOoG93P1AlLSRSj0L8ZpozqELkzA5iPW2JsZewTv
muB2LR4+yrDVmGRPLUy2PgrTXVqkoVvDHFlnxM0rF17HdQ6VVLkh7c1GeIubhSDj
Aw8fcl2Z4fvcckoa5P+/K72kXeyPWJsWTPQ+kMVgv435H/AuuW8BmFLYIDh5L9zd
ZldRsy/jEfABSMdEmWMNPBKl/isrUfA3tnlHmvrQialieNRLXJspoflGxSoThGwG
x+0J7Mhcc1vVKJPTNC9mIhOAfFUgRmDiSgn1ubpasRNmIjhXV+qPzooRng9YWYuD
hw0W/cK4gX3z9nAJaSfM53hizAK4lX3ANjbyJvwWqJ8+QxO6NI/qoFhvALV4yNlZ
QwQLp1OOBLep6UlKpP/bRtMWKa/2ORfCp5o8HwD0heQo7CucQL/0zcKNB1YzOZXB
49irsOz3dsRvrvZLMq/53z0oJtwOt82myd7PECSHUVv1Z3V3FHmtWbnqgYGoQ+Hu
sjXraNtP1Lg9pXJ0+DCpM31Sa3wDIkcgCVj2dxe2YWNwkTYkeW3bU7F/7edHLAGb
fSAG9wONagYQ1k+acTwEjHD8XVnZ9qeEA5ue0PKFOBwS/WhPHf4ce2pYtmZhuDFI
wYrIqLDWx1+F9YdRDPp5l7nyq0sdwZTgH04OgcAd36xrMiyVMnPy9h0k0RaEtJm8
zC/KXGwwCTAv5xMczE/GoB8JtxOwpEskrNC6o8MBALMczOppH9r1VYQQjYgFuVPP
FdoXKUlihFwqLiSnJLvtLJMd/J//FoPsSxqe9zLuV69HpQQKCaSsYEUzGcl2lNeM
u1o0IDI93P1IF2aGM1jRn/XdBuq8AGHhiaOxjE3ZH3vVuQVLkcxwm2oDmdjnimSr
rt3DmjcvT0/nhYAt6Bjf9ky9DA7i89vIKufQNQBBTjLn52a8KCnOQiKHFKw1Vz2a
draNlSnL8cE+uPifR44wsFtgW/XZVMr3B5Sczkkcn4AuCp9yWV9+psY/Sy1lFEIr
kJtn+39C4DPUJ8/bP4ujhxr+5s4RjvlPMFHCKRhqG6L9Ln3m9WjY93KLzs/Uk+Jo
cmWM1C9B5V7YCkXlxBOiVTI/19FTifxGEZ6Q2kRlVncrslUI1DFKQX+9lXg9DWsS
O3csFtUE7CODtyXVpNJlLA1K/LjMvvcTjFUFJNhiveyw/+SGJP5+6+1PwsQSoUZC
R3a2yLfZwIk81NdnI4aYhWLf+sRuw5C/5cV+a5//PU6QYSv/iim6OcVXVOLmHmxE
FAv+7sjHKqR8orxGaYRGZ/+D5OlNYPhW9XpRYSGHMeM1bvJKCoVkq9RMO77faRtM
pTtwle4edFDlvf7BwfzZyQ7qLC+Xj2xawfH0haJhiNjFFHcTv50R/WfaJ8jVQYGu
wDMjBl8+jDq70OI6Usqp6vf5u60JMZDjrjGC0CfS2qc1xpWiaLA8EABaxPeIA6TJ
ekIXEgOUe/3o8Hx5PTYow7xSlVzUrXPKEh+AWseVjWg8LsZHgTq/O/BDsg7h/Nu1
QhtBl3ecIeGZJryJgqW6rUNW/hT/eP8JrYPHJoBmNUTkgzdE1L+LiczwM9PMa6WI
405+dOb2JFVquZ0E4fk8rbCgntQV5OMV+7a2U98/L5bfFGCxdOH+7q2rMfu/nPSu
LDlJ11yFT91r3S9D8YOczYFJvOswcEZZ5wlWX6vntxnndMzINzRGWaFojRnjRaqG
gktmNNm8wZ50ximEbf/j9EfRKap7Jkwg4EGM9Q7RgIWCBbqcSjuNEXjuEQTzrp1w
WxcMl5hRYkwHJiJOzyWyPqNvbl9v4SUGLcuIPqgMsGBPuZtEgWA9olK+mZ3paCSK
1zhz/git5wYALGeB35Yy16zmFf6WVei30zsfLpf4yXRyFAqH3u/OFALmpsDQy2+c
UcWcSC7onRjIteLGkhhGLeaClhQN4V1WPd0dBdePFbuKPFU4pJgsT9ueU7hK+jVA
/6E0djx6uOUAVyYgvbwkF+RUmg9kOCZCCYdAwrBIEYlq9ceVIoChyOKMWOQJNYQk
SCgs0xWrq6raGpfGJT77mmvEKeMblfGuexrXO6EMStJOwV2AclCel/XJ8ZNOZ+vA
G2FWjXGUFNdeO2bREjXSRVEy45fwRAAJb1hLYMcVzNL9dI7Ny3flhHZ1g4XgWfdB
1qr2uwhz1n5EmI0XjjI/kRByd4NuQDYldftRfK/H23Udt3uVb6ZtOg78EE+wm8UR
PpNQQHqyUeWDgpZuFOOjHpYWT0boeGvzJoMlwB5+0ba8OUN6oHqodU0RmxXFcsjF
0vSCVpy5OjQW9Z6xkgP36ClCO47bvymem6vM4PwwTAJL+tk6jwY3h0Qr2MqQ+PR7
NwUdc0m0SzQeTnrYvcSsxCsm7r70YuuacDbveVP9b0Z2ysd/JRb1DvL1B4J+R0G6
fkvEeql+X4LsZVXbiim1lkpMB+qFzH81ztmTyJ1MC9S+89B6fT55e+GHJYE9TtcS
qMFrGB7UVhAPDsw6Fkk+wEaF0wUtX6O0ZXtjRGN+HQ5Nst5l2A4CL3g1YuseTn80
MfPN+Go22Iu3H7QF8K78pKk3d+aVMWWe2eV8BS6rt8WYARzP7R6U/kRJZigTovkW
hTLb4aiM4O7Y2F8y2h0OBNmfbtwNmTOESDUGcLUVkmRDDCu9W06tcn2qZKAq1CYZ
X6sYH+IEPuxqaj/BQop8FLccHnBPqmc2EntsdtrjIo8iQh/CWS0Gvm6PdpztgE8+
g91CtDB/j15JZH++zLOtFoWv7cXuT6TYa/+ZX/z2BJPz5Mn7cz2YroapHLp9dput
IDzDfC01ZZ/mhsiRwAg6HT+G3MmLV7qyIeqMkqJr1ooUWhb7t69WnE9PdgZxxOtb
ZuIgpvCIOF5LDoTvN2WOjAqLAE9CxUyo8nEVCcg+T+AO1pqRlFRiNXhlLem3xNeH
mc8l7FFL30sqS/KcZINzPvIjspFoKROy2ArAsQk8g6UQ5IDgukDBf5N9koPy0Sv4
Tt7qjWvVF04Ppcui54WB0fzCQ5LZZfJJeqCfjhV8Vf8AUHSLraCYRrzmeGVEzTEq
S5i26nsF3weOV2Lm98R8YYdQLVXCBOInERuteSaFGgkQtNV+itrTcGWKHoAChZqw
Z8HvvQpZSo1H0fP5bzYYAvYPm1kfh8/GcQKeoSpOVUDoHEzGtLSxfkVACxgBG5xC
xGIFAKMQvHUFVUn7Rk9rlETdgRhvuKP1mKllOOdxMTKsYVSyB2Y3rbg0hSzQ911X
qbyavoLHKck1jb/W6NabSsph3yI5dLZB8c88eRUBxRF/LHdqCeZpOHek1NoJYc+f
BkBjN5j3UE9mL5P4la/ysj8Vci4KRMkVxCHG3/z+bQLe3SU15CVafi+Xz2I+/tch
NUYHiOWnKD3hfv6ca10fF/wIPM+sDlmxE3K1JkUc1zU7TdHmk5hIB/+OhJ6yPN2b
y7x0ZFvUYp87WorvW/JPyHps+hCdUaxz+QWWBRL9HCPlQBLhCIPavfqxDQcfQMq/
tdbwy5QlyzxuyqgJNEOMWiuu8NjoihUA2uGGvcU8YlHbp7GextwxEi2c0SQBMQnC
Lzt3fdHyNo1vV14+EL/B7dMZSSYNqD9tNXnVAJPMRSXNn4x4WIXd2i83t1etw0hQ
0hcpAiQjQQWS8yHhSaBrROSRNmzekFYKE9/tra1B/h3hCOnyZb8b0RWOauCDRBXj
9PDoA1BfFLziaiqkjIr0QKeOyVKWAkJxspEDrqWqUCXDm23GGbukL3kcI3VZ5dtq
xbWyWt+MyqARAjQkUix8UkgWJyU0a8/z24kJlUSS2xE4MAtr6bEXWK6yNTjKvP3d
1159A2mG9NWc2ERpJu7uKMPG/A836EGnaiu0dtXOVyR25zHkhB93TKJKd/hR8KNQ
uHMjLptKWgjWAeHEiWyR8hd/uS9RLqDxzGBx0XT6RdzqEmltv/VJSzQYiNmap/J5
NhBMVk7uYa19FRv5YwXA3GzZ0CLV5ALZYzdybOXdbbqfF0nIKE7g4RziLduWPKsF
C+24abYjdYSyEiUaaS4K74vR14Yk1FzN7uEvFCyoW9Pwhp8O3nmFnAFwWMhJwG3G
1/BNG7emWhFsmzBKODUDfxEvXnQCvupy70NggPz3eq6d04WSOxEOso4o1Z1wsMHp
F843jU/l57CVtWIJj2bJ2VxhgPoKvMAaIdYwTpK6uh+Cjtn0JdcSp9DbpgUjCLHk
pjnw7txDkInnZDW0lBl1sUVTFSPuJATwPhoIiW2yHAZbUYJRja3Ot4WRqXDqQD7f
AYljaJmiORzuqzIXqTNHIZuP2QfUPGrIHqdbZa/1x9urFMklvjA7bS1UWvxyAQxC
3V/AAsbVvChbgmyigm2GkUy9kcDVF2cBCWBCaLXvw0EtoBkO5pW8vVcN6ky/ZWT7
3UKo3KTs7Cg2komDbT6NEJCAUQsu6JYURSiIIoLPPK1ej4Ed2Qms/cTOdK6by/D/
LfilvXgj+wCHQL/Y1w7IUXX5cqm54yFgXIo9u+qf3KWaOLO8wYFELR6Rg4R+0WT8
b2L8F9VcLTBPYQrE4cLDYODuaWAXjnIjWajQH+sNY0LAeVv2B8+Qft2SuCvEhMkW
/v97ex/XxcNdbNQP1Ur525B3pxnkeZZkvpwBlmdzFCE7wdU8FxVqVr0LpZ7k32XX
T/rEKbwJgXiCIHW7dLQQhjJMs80DtrXPeUDb+tDAWwVZz8CCVuvpCXkrZoBftJK2
rPfGxqmNVGaL4sAeT0cgA4eLlatrCpP7dapwKwPBqX1MjcxbXR8Qbg8IllXngZZF
XN4Y+yB6scGn7a9/l1zkABG4/2koVj4ns0bz8OjMd3VI2XlPTK8U4qaA4pYiAp+7
+mTlnK0sz+ZMi796/dJ9fIZlQtdLPhj4/si3l5LCvY/g7J61wqIF4UZx37O89rlc
twYhlfw/xsbK73LVMri3QLqW0LGcxHZawaDE5aglkn7ijgMxCU8uZYzHqrSwKmzH
wNq/HejmbzMeuoCCgVKvfKghhI4ThD+lDLN3Q1r7dl8ntxcF7Hu7Cxzsp2McUfUp
49I9xUQGqaV3HHEJ0MpJe8g07QlHcNEo9eTRn9XjKg8FIFB0vbWm0FdDOeDiugHh
2ulRniE7n9dHav08i6Fb8qsYO1wwzWTTE2hQsY9ArBhDT0JlmRG65g6gQKHN3jEq
Z16YeTOTWsT9fdGOjM745F9MhGGtymwv9ei4iB4rzFkhvJ3eyhCpu2dAYDJ2aJaU
wbeDX0dr7b/z1qwbrVHVMZzfaD8c5g24A8AhIdiuSWcA4AtvltkUyZ1C5b8Ha/MZ
fUCd8Ih9gE/uZtGcwKYrx+TiU/vYJ2WyI6QQqbE9DbvthdjcJKnl5UwPXa2FBCZB
yyFcbE/wgivy5fUkZYRsXTXSOEnLsTN9djSRr1amaiYF44lqRNxNwBoDjAaPeco3
LcwlWeTu0Qv1esUOh0yOcox4REbw7z+UW8h+IqCUHza/8k7YoTuDQ1JRxkOFxNqL
Covly3LAUl/G7EXMJ/qw2A5KKv0QWSxmkapXae+GG/CQLBUzWIufcjZ9SJzqVOcH
wJk0Q4mWuWlpqd7eaDzBVmo+En3+cJwEg49dHLRwyTt3XdqNo7mDw442sXG1W7C7
XiI8fgY5UuAY7AHERe8MRAJuf3hnUaJ3XeRZq0nUVoDje3J+ONwLXhZjsaJntioX
Z85YJGuFBB5igeFH0VWZb3ICYLFGdz7fF0LGVR728oAM4DUALVxxfudQTyUl0I2u
XbsUW+qqvYjltwS3rNBbbQ0oXs4EU7uEsZc28phzCVNfxUpecJKktSX8vpyeDrqV
HykC+0N+ffk2R/ABqBhlkswA6fCXqXw2QZc0uGC2KTG11oTW0UUqWpQkUD4g9Dnq
7lBfnUVVmaOc4H/pUVNJ5aPE78qEU1Avjz4kDfNLw3LgSD55Jmj4Pgd1qxF7xfXl
pDnhYTRUfR1OWN/INuu+7ItNSpx2WXWAGe30paHVn/UC1dvSyPOacw/BOWo/sQfz
ON6q7GPMEX185nIJ1rgcoCT4Fi/WrvfAE6bKf6ILfCBcK2468lZlxHYb+P5IjfgK
Qh+kQiyJ3faauEVgUDKlRZhPZhGsGSiuIGYzEsuo7I/BwgEZowNVuS5UIo1FbibH
8lAJHE3IZfpyuaRtP9FJoPdUDnpt1UJHcxy9KEP8+H3znBIjXJ0t0XYEfAXMgj5s
twxKK8cgdQyEQQgOXnltwNCw462IQTJ7l2mFkAdkSCENwj2FBLJp/Pe7sMmsuSEc
NusY9i0i7GkGVRgqiZfCLjxjsZx+sqrGWCjgyNcByIfH3F1o5HonVaO1CcgHtFGw
jlIoUjEwQgOuxMg9zd8WCA/hNlHNs+m60kEvUS9XekoGNP5LArA6KNqOfcfFQ0tp
RnmcQ0sAxQ+ESEOa3j3GBrO2ACiZatHb24060FKieHQqcdHS4dBYeZUUCYe0NSRt
VpBxbm0Jk8OtkO/lbtYBJ2Gq4kam1oL8aQayC2GINDlytfVVs/XUXxF8zEC2p8ZN
aXh+0DDjNJO1Q99rgKMkZ2bQ5ue7Bos45WQBRevLbGeQoNhbwV6PjUU8igXRWnl2
MEiRR3IZLtl/KKpeGDU7C2fslWEZknUBFLJelLzIvP6BvHhVLmn8d8YJun4A3bnc
Z6sWlx6zJ+PWxahPLP2i8bjJQoCzRTrXSRAvlTz+ZpBiQexWXe7AszLkJzUGmGDW
tBWbRlR81Gv2jEp1Y8crHVYPRsMlI5xGNyZucDmxCEWmR/hnwzk+3pR6gtsPlqgH
e2euWqRmrqb6fv6ih366WIC+LwPiZeuIWlDSO+7v0xV9x2Ms9Zc1vU6HQW4qlQX7
l3Wxy6jJBErvALsL+cc8XBHpmFCfgOVF7Um/UUkwLIB9936EdxrlNVEDldEpUJqi
GNQpka+lXTSmPqyP1g3wnGsU5O8xtajPktrrTPYq97xleI8oTXwGP1rYLnPZ61T7
S9COnlCPAnltUoJXR8y6tOKz6kiZHvJX7KfLznHqYARqtMnYHqImMOTbfPvSgVlS
iBpIntK9X4h9FKIJw8xVDZwi+XzJabzCiuf9PpyZzuHfyv3QQJOYCY96vP9sFWdB
afJTP2fEXPsiSzkKQSeLxnft5/FWmzVjFpnbA+SWBErsel5XK2L0/eERxxAnQXwc
s2JedbER1hAYr54JeMPUhvWD39iq8yXCreJT4KyQtGvo/KWl4HxWJbgM2nhNJNcG
iy91zEqJru+sgN+VjYJKt0ZJVvB3KcvrPZbC7O3mFmNZ4ld5+e2xwLuQVvdG75D6
Y3whBERejmuPcmHH/fqtTx7RzpldVCZXYZgxWrGBz3AXUWyz5O/AaMZVr1mbibls
nDy8eTUmsCp6ZDdzars5OQFzUMoHfArsnzUEtq7jlREHKwwseeiG0Kw5vLX5jtdr
lXVT+XmkhQhpa5ZGWE1LnCBXQrfHIAatfOKkeUVO0CkU0yfoxnpYYGwtTa1xNVX/
JC5cviaj9OsK704YzrmXdsPuYxj/1XVUTuFqlT5aW4JNtQMkAhOc1qrVOsqMngvB
UE+IN3D8jN6eAAErvbG7+hFTLeYdosBm3V1DOpLXxbtrXjs4Gk2jbPlBuEPobHu2
0yIZN8CBSHbDXsEZsdO4EAF1YfKON/jILBrhMW9kEa7alxGU1iEfk5P1k26Qia71
ULuKaF0ocsZnXtCJIy9Bdc4GfBtCZ/zP/rZKqge0Qlb9S9gW0cxxzE99fEiFllvk
B8UDaWgq6Vg4lC4XnMRQ9rqhT1iWAFw2tWC9MWzWOQCX5Gi2zlLsLBD3PujV68pd
YVQiwRmZrFaHKzsoUG67VpMZX3skcOxvsZTMFGS3sF0qOoiL0FRG8Z+WigSBwNjl
onJuG1ER8/Jg1AnRBRbl4KaER2CQVmNOryGSatAtDyFZS35jBEjUmbW+ejNrDYJq
0Ls2j1AiIX2770mxKaFJuRD2MVEbfYOIy/zE2phBDP2DcIGlpwxT/E+uEEC+ySlg
xyCq7kECgiVmoTaM/Kjd4YiTuxuXo8DVu80DSWhRmWVmZeVzWKr+cfGw31JifysQ
h7BT1RblCVVk3YAvAmn36Fu0az61e3wzUsVVifG7xtnUpqzVOWBmByEBs8mPsABT
SiAIhEP+VzQjy7LX1H9qi+qUjEjjDkGyEcArFm863g4gbVF+3TtN682TjQJY2L1z
anDH2Xwgdmx2kh3mdmwkafaHkRQ8SWSsU82RWQ5eJvGh6aVN6Hs6m6dNG50tWVVx
Ho2ES+ijacpB3l/VzDFMX2qLsBTXR23e3OzB1mO1USEr36H2dBcQwCAs4JkQc9Y7
nSWteyAqmBToWiLXRo7mlB9RkH8ev/l5aMbt/9x0D2E0X8bY3hZ7HwOO3opkaJaZ
165K+kM/zS1r3+UdPsnnVdOJB1horuUauTIc9dELu0KFmAFCoToS0ipGfGWPdoCd
Y42akgWpkJ2pCmR0OHCpM/jnjJhinSCYUSc21sUuyu61/yeC1Pwbaih1g3QGlyLz
dFh/9QNu4H//I10y204oBKDG0OLUd437EYRK79SY4pk9dS68TcF6159Sh3twfDlO
adusif5b9+j14iTc0QeoOJ1lxH39/v1sGkKIcpokTkrOuN1WZN0Ucr7Ot5JoPOUd
Uk5JSv2/wfCSYGl3ICp64V94X42UeLXflsUIJCibCbrLMnIEEqT4ImeGM+lFKLJm
xw+AQTNqLM+lDlD5kvVL12nzrK/5iWyVGZW1oU82N6wf63CFEb9n+zIkHfl+P0WY
biW4qg2+RDjCFmNqfh33yXRk/DR7NczMvx6lFP6W3gLUEyB8goo/yXqBvxG069DU
hap4em7O0oqqppn7QCrHenIVkj+JlgFYZnuUhkCYckonFqPZMBiYfy+x44RoTfVe
sGyo6eQIXDf//Ag7AG1ZKtzq2W8bXhfi3Q9rGSrd/F7WWdhTStL1Zr29HPUwJe7A
UZcF3sIGenUGvAMb5W1J8p3F7TDED0syelSeXyftML8U7e14a1vS+JUDGVG+XW43
o2KCi75Y/VBTKUd98WsLdxa2CXt1tknoxtSPXnqCo+CbnQaU7KnaqDm3hWE61+KK
vTfEMCY7A7IX8H4NWheq/QLHAphCB1ZQZZ5rviuVPRrH2piPCdsGP9vhvwTMv0WK
FHKnjHvmvhsi8FHGUsro/ejpknY0nDsGSLahgjkFK+ebIqp6DCdlRdrP9etXYwrd
goEBZqi9c6rCwyroBT+ZsFL7mDYn369oVmZ1h54gN+byJiqlMhOUDN+Sq1bOTjML
MtxHR2949q1ULcPOK9wJk7NkKRNkQnFjQk+jzY5UljBHEJoxhfFV9e4ZcFRDhlUR
Z4hEYwWXIamubtrAIwoEbL2Eyksk8d8LqHysBRXnI8745OtcmQeRLTL1HZkesdfg
Bg0Bb4iJCrfXHVmkk+SNi+JmYaOVmOQl5h+sIh1u32Ttgg7XqZJ8CDFFyEX2QSNk
6LciJNZYyYfWd1hlIV9LyKcqZt1ox4945TyN/wOnj4UXtXeYZ8wqXEb5a+2Gpo+R
txWYcYV4RzKL63CnB7QmXHa5uvS+gr9RiU9azvkMPt52n8bHEKrtNVxkbh3d7Nc8
R0bhfHf9us+jvrTShC8i94sPEziRNpJ0vVU1ja/09dm6OFJCcI2N9oqUe7F0VGmO
VCRgNVXl/Qkd1wPdwXQRgc/5h3R2a/xg8qnxinJYPJlS+tWVtf3jkuYgCYBRynQR
s4NnJsuP4hCsbgGw/jhTxrdLw4FJBOaH42yysfuaAEfD2Kk9wTBMqEfXQ5QLpFIr
ijushHKABxp9HQGPtX33/Mn/7KBw5PKvcPSvG4b/dUzbI249ZM5HpGvzLfB4Qv/+
6/LlS31TunkSyP/I6ALWriU3SzzQxS4qi1UxYeaWRSzvECo94armc/0XqBbc1aQX
BFjOwhM9NZ84knx4p0jKjOKo6r0JHXp02V0pNsLPGiH/Zr9n+5hN/pWmtrR1VASJ
jNBPwhkUwiwM7WRggQUtaY8/JNP9MXsiyaSYjdBmYq9OVO6kzDF5S9HLhlKVjZuk
oNiLC5TwERNlYJ21NcCGFvNgDJriyu8VG8fXQSgkTD0WynHJQwnl+Yi6u+wu9VPu
LHE9MPHQbPvJmiYB2MW0r3WtO2Otiva35y2/j/Fnuod1+lfcwEGk0gdSQ92gYE1A
XTTY7K5li4ZGr57xFmfP6oL2SNNu4XPhqWYzjoebQWVpmw/c94bnFWd3eReUUWk4
3c286Zmw9jltniKsyEBdRbg8MkE+G/N38RXuotS9zpP/ygbKCEDb3FdIGR8jmEWj
TjXs3ITD+Cut7Vh9o8M7+sXPc5eFm/hAbTZSBMiW9mStwnPt4E34UotvmqgSvo1O
lQBEUuhwUn+7mdQ/B7phYoe13iYoQwiNaUGPhQgq2V9FJpDVRTACaar/kUnQxTWl
GKZ4AHq4/vdMTvhj/YKzjjZm87D8uTCyB4p/80cromtMz2R3ViuYZ3DgOKKVsZN2
6uRlJ6VvP7adT4O2ffOe1LN2fQEt28w0/arnsaWstO8NtgQmk1uulXVqV0S9jUL+
jfb/Ue3ZBNPGxCO2fJsNA3V6WLDXeY2i03pjT0YtkXTW4qTUoDxHFy+cAfHYyCDM
Bc2LRIdg0HnYnFyWSrMZMujvFoVSMuLD480NHUwwMyDlLWxBHBSMCH2/MwT/8SbA
DiEKz3895uURyb9RRMczXC6FReizoW49oboAcQg3P34+dnLO/ZEXnqFsJnj9Vr0u
F8865UY3CcSyt6+RnmSmR7pxsCayHkT8HdH0FDLXANuWri27y4JgXIZh+aaEjzXS
grcvD+8UPdt/vG2l1v5WnLIysquZpV4j7C8TkpnYZyLK82GaSo+uQR52KByeB2js
ELHnZgJt4z7T09k1vF/6BZUsLarMguThCmiqBiub+t3LWEE1NkUKOWXxpdzy/X5i
D5ZSWJQt0a0MmoZcBV0JfUTc+rjFr8+xYjsO2F2rJHWhVHAA1bBMCirQ7chFZOBG
s494Ofjj2sQ5cfhNv9qm3V1dhSQ3G7mBldjq7wIKWJE6/qiJoo7L+PEeB3L2WLFM
6bp+Ucr1ThSyAYArSN1uL7aqb3GFh63oEn7OFE0oI+zQVxfy+QA/z7lFQdjOmAvo
GIUtpcIvsoArfoJBHx2nOWfj1FO4GtTnHQTyFpLWrwgWNps6Z8r7FFrwpvSqLO6j
eWmlKlUkiycDAZcSCrASH2MsnXRezHEWlr+qdfMqDqpBhDclOx9Sxh+Fgqf04XNX
A9LxGQwJlom62PXSFUk5yN6LXfM3vpk6WWKbnKOWHrutyD2pyRu5JkUAk0QUsFvd
CQKqLAzXhZv5eKK6RPOpw1UTytrvdOG5NoJdOfeCsTbtVIOz+sizDGdOvKxlnjtD
3thT9n3ILQ1MtLcf8R/mSC7Ssq3BN9LwfPR1uGhZwiPIyP2NHsiFVEb86KeTjmEm
awasq10ymNoCUE36IuAjf6ZiJd67hHFdYN4aLMHKyIeNfhlStfpnIzNRm5KBtsz0
u5pueTCWnvNsIytwX7LgRMAb6wk1AUN839r6HVQ2XS+3FRaSPlxQYLdTdMdOPnJD
iU33ztwpfYdZcXRtvFDX7QEjeAMGdUkiphjTvO07q7W5rC+6h4OaeGXD8pb7OAGD
I1R1tfm1N7Qi6pibc0MsdK/LpDcaJoggaJ+oR75H4O/f2bQLgcbOO/yK55vM4GUl
ucDKa4YmJJmRcHNoVGqimiq8zpPKGMOfTSC5HMLZpA4P8/xc4Y6oq217xnyh13bI
wEUzOLhCNEcOg7vwjggqnUavbFv+XUPNw08ZlNXHS4tkdIkkboGSwtvLR8zhsOtk
3pyOJkJQ8SkiOTm1uzJ8JRtmwp+z/3x/ElS0u4u+LeY0TAipgaf5aNPRgQSW9+u4
H8kv1yLCFkbFwKEjT/3mBW9wHZWHSR8dMhDEVD1Jl6QnaabH5Rkkqksb+OeZK207
RPFa3SC9i+7K5Mh37LKV+G3PTCj3t6IrSKj+Sb7NNQbCOAg1FRMok1CVv4+IoCwL
LCVkiTsz6iw8z0Vlz2horpVWofy+gpBNbPMNxwF94MV1Vc3jm1S081hU+w7sDROu
Y0Eru/pRIZF3GVV3w7g2M3MtuifH+sqQH6KogYPe/IHeFgCX3evWzKJP4GKpR+xO
WsIfg/E4lnYflgMhl7Bt096JwDePKA5f6DaM5OXxpbRjXr6MgNEty9x3BgxN+7x6
C6KCaWlIFxtpzzAjo/zr8qTc0wT/CGKIQvlI18FU/PbT+8KcHugKDh4Xi5WrJ80f
BHJTeTBdEsPwgG8N3B8+qOHXU9xTswJGAZFGLVL//iY00TvXOs9MWhbAeEpDBf+P
UiiR//VaW1YlWp90mjWICCWHu6XLxzxITzpX2B4jGYkHtoC4XtYWEELwcz6Nwzvf
DY2+POMrzWprQr2KxlHfIPqTWOZaQMj2yF/ODjeZAvtgd0o8bBO+ONgutcg3D5oi
Gcc9uQm1q5ir5Ek5Psq31gT5mRlFZ6V2kj+cOd5XMSomOpITvuxSbP5S9L5CVbo6
Csu4ZjauyEFFXrCBQvyhbNCGjU0LjbNG2/++zGvY51gH5upcOwcXxH9f4CLV+Mrq
Q47uFS+UcsT+nJZ1//LF1MNFWspbyopXPH3ZhwQFwx/IK9jcTb3tG4RGYjf3v0IR
LvQteqLw9zHu9mAcX2KaSRLOqXxDU7Ztz5G3CpAAWLCjRJhwHHvZB+vbB+YKtqbL
6OjhDtrE/NNrtFkKHuwxTN/k9+cLqsWN6VFjw0KRwm4208uWQrOMDbiWx06DmZ5M
GHNYeZ97isCsjd5Laru0Bn0++RkS6DgzuoBpStGXE/OWYO8tIfXlAeejw7bJCzp3
f+BmHyLhJmXeWO7P39CZXQd4sKq9KgINWOe7QbhVFsKij/Miv42di4Oz9s45b1O/
Vf7/lrJ+tSXgy2535qY1yM1KnKiEIjBtrnaEtuxr+O8lWz67o9VAi+xMhJz80m7C
0Fb6zSIJE5eM/PE8fwjdZ0Ldh9N6ymlP0zgg29G68fxprm9CdCdzInUvkDtaEUa8
rwCY5xnVC4cSY4mG4RH1GEb0hXy4dYMBw143aQT1K0Ya77ekmzXsTXrYRCS3Rdp8
Tw9dvd58TGYABQOZeXz2cfRX1XP+buBxyTgJBNIu6INy2Isf/WDTvO9+6Jq1zAKQ
lvfGBCso1CZ8IIH6NmRBUMp6PCVNt+cMrUMYFUaeHkKjl0UBJgXZTDuPBUHjxDN5
sA1UfTE7GW/N5wOiqqQUtRTGJN3WQtxORsJtP0I1YDAfSxlKFyIgFImYeusXHzu9
yz9D2XAXxQ7/NGYa4vaA2mP9nFEW2qe/v8uIPVOyR5uEVQVIbDR0wN5oU8uyzv3D
Yg/E2vAEB8pq3vUK8yETO3hYcPcLSDDNh9PxXVbyr3wb9CpFPqoMXcuketEmUPPS
3g95Lcy7BTC5uGOKnz3BOdswHK6+enflOW+WmzWts2yjfJ+r3a0l4iYq398rmAa1
1U4kaGjXFEPLPRnqJ+L7XAT257b9tVX7FMknD9D4T0K9MKe+7yO+d5zk9rCj9x/Z
WQFaN5M1SPnmV5w1QB/th/tK8lqokvnfG3X8HZ5LyPpdB+PWuxR0X/HOrrfzcHhF
5mgwGR4jFGk+m33MVTw8/D0nEM5SqWvHoj6Rjsu1mXHTEeOQVRSOdCxPantbEWK5
7jFk5IJUtNaXr6gDGM3rp3tnpGG+GrZ8NbJtUp54EhSE6xeHwi9pNF2KZabsD5UY
K7jhYsC88OCjXMWxjrC7O4NN2Hikwa/1YrZ3WpsnNrFlog4uSn7LVpPkugg7HjKP
+700dbSYE6FEt8mk0T72Gbt+tIMWA6mZei/BfxnMgT0Hfdn1+CogMOIjhZ/+uflP
y1+pkAdWUz+mn+n9lfgxmrXNX38Pa2pWaK3dI4iA39OyykZNgSbSmG3iZPmRdwfb
v+SUIAFrBtG5JHDpHGfY9mn4qGVuXkXgD481xIqefsWTUHHS8aOOUWvf9+QF1q60
OTGeSaUgKZ/BY7CmQa04SJSnl2BV7ywbkLbT4Kw2KJYmTRZlFSxDP8dK8mgJqdm7
kYqr+KEbSNO4w+9LHl1j457BHl46+ZkmQNmNv42abUl9eLuApwZjOrPm+ihu9GGE
HoldNMRF6xGDZCMAFWGrCuJzvOktJ+yChSSxJWThDe/4efm5oEdaKzL0ylfm5qKz
32/NxG0k/58/eos2W+QbSU4c+/25punAaV0b0DFIunNtv+VER84rrdQR/PmSPGgf
DYrc2ajmRyhwX2O8zcWs415aUV7gBaq9YDblBmdn5qCsM3NZ8263Uz76wyxui0qA
DuCWVy8Z8Hy52dlK8nNEbvWMNyJwYazbcoIGdZZwCVThdileKVYHQ8Crfb6sP9a2
un89QIz9ZBWx1hnHLBYy2H8Z8gkDWGAKpRjH8cCf59g9m7sLbttjErhOPIDHmVGU
pH77/x5IC6RGLeoBsS0yp8RFgxKBbY73Av6OXM+NUxaeMowRVlVULtg3vqSCO/To
7dCzB319rhPn7zOGG2mJKApbIqyUg8XiAuIAvnSv5Tq6ahVqqiKhb0NCOk+5OQ9T
8xmaDWhEPGzvJETrwmCF1X47INEga/hnsBIxf/9txp9GYVpHVPYkElZmCjX3BwS4
Vd4GyjwKs4U8SI/kAXUCBNtP/5kU+Ruo+LWo8bE6a0EV/SW/+hkXtI84VHtheTas
8sVrnpQfqZzjYYcYkS5jJnw53yibCqYuoCPFJzYTJpv6XL2f/Zl4CDpJi5w9oNLI
fll74ZXkSU5hqp5at9wVPcHebvEIjxxg55cbpVMc+H7NtFI7YG0HD4ibwLg/Q76O
dTP/uOR9vDfM7prrdpxinWd7s9Hf071nC3zJUooXNy7Iz1T5DZ5nmKuPO6uq0xa9
6CELqhSz0R9C2h1aR3sY0s3Sv79gPR2A927zpILsoEd7hvIJLy586jmqnAYaF+Y1
MaXyRnVT+4sD9AmGehDGNVjggJByLVOC8i1Nbm0LbUzWx3nvuOnqyZyS0NCd8Yb+
9SoVSJAueoTLKVVHgWM6tInO/t8rcTvAGAoke/VK9Dv1T9PfDzdXY3iLUMiTVVKN
28U8SSVDTT0W3RoaAPPZhWmXwmX4nT3aJPn8VeCG6ItKJ+JIz0ddICHeJcxFzLc3
b3XXpW0OZmECc8oekbFLkFa1tzKpzJWTaio25Ta4DjD159zrmcaF2EHb4pM9d8W0
m/NlwBnuhgpR8tyYWD2IrZAa1ZtG7Nv06TnlR0L+jJ+IDj+fuAmihPFf7/iBAZN9
PsjUcxKQ0/keTaIGu1Iif6GEFFmspggvRERNZq0DB8egi7yPtT60bmHq8sTTIBqv
5KdUmLIOHaUFP0J/uHbMKJR0VmejPGuUkdYGgGBDnWyV0aJAsIvbxt0w7G63rZs1
UgDv+vQpSqhWcGlowIf7FJzFZnGZsfKkJ/TtOb7w9h31T5RhrYdAPXG59RoV7HrF
kOHdIHO6rE7oo6lYeQPE5ioBZmRn0+g9lt/8lRdB6NhH4YPQQl90bsbDdIhXKkIC
Ws7qz52WBBua6hMllM1s2/7gAJmdE8CRRUWVp/MWwNpa2vUHxXebwjBNwh6Rgk0n
/r8NY2rbqKVrixBzJ/3HsWBUYznQZadEnpzUx4x1j6dZwcx3On3Ffg0JQ1qbNVih
8+s80eopcBphOMrYakRGOHtASTLtQ6FfrTuRWPDd9UPgySlD0WBMOvoV5LQ8hBNW
J8eLrzYP4MLz9ppyW29QeCYR1Y+TFVA+THi+zxieynbo1LM/2GFIXvo53rOX0QIH
cRpsnORt6TJLBfYx019E9zVKo7pcBAGtvTPIlmJYJB0dJLw5oB2lewLS4A3zYzEN
U8d8y9OqSMQz95gul6PNOeIQxxV5GiZ2vtgStnJtQn7G+4JKNcpc0sXBBUgdgxxz
ITCNarVJ3M9vEurc/Gnztm89onUG45kpuyKCwSpKriwxkaPUtgkj4YRWcV6HF79K
18BVmkxCR6KCd05TUWf13cFvW+ULVXyTumWdiuelgg5uoigYtUyiTQwADJXs4AIZ
giaW8ycoM8GfwsJwu4Xsk25vQpCgAkaAvkGEClcw1wY4h2DL6jN4vONkjjFlezEM
qmBjJ4w68N1vfCfXXK8z5RUmEhuWcBwtwHWk9mfcvSms+07pezcaK1n6ymXun0N1
35/9rFj6w6IW/szX0b8YEvQFucOUB6hLGnkP/sFSVUHVo1dKzmuDtovDn1v8Tz4b
QFOaiNVIQs6Gnkr95d9HKwsf2F0lp826XTU2VklabnsQ4v+nPEoR4PcOUAmUQYPj
xfzOnDAy9KCh9cN7f3z4G4segQd2AuBny9DrI4MOFyfgnFLcT1oTvwwaveHvHX0B
2WrKdirB2DzQlD9j2nOmYiIdVx45VrGHCTqfViH7DPwfXNXRd9CjMaphCzneDoPT
lBwLDP7rRyQwMa0cBDj/+SOGEl4W0aVaTPg4LBNuXhtAWuLU465LIaJ4qSRyh9zU
i4hOk0ctps6chBUjAFq5XfnE4xQX21CjSKvqitugo2J2WPxFtBOffwsl355oWAZs
OTesZma5y1D37VX4B05KZ7D1LwxI7zXb/hMIIqcP2OfObdr1DgR1WtugxgnF9JF3
cCItgj3WTGSGifSslMfxwQPFBd8MIM0wmyqnoDlM8CTgmirPvz3O9eLzjPY690fz
NkYKu5CZPBEglrWYb8ibEkn1CDaBPGhc0CeRAKDW0DlN1CIhZ7EQYpnu2XutryUM
3IwG3rmvb5qpotJmeeApMp43DZ6ahBBN4uKOy/FUFMEnLXzb6iKrk+wCgJ7xJlxr
ozxRfzNuqTslGIwWae+jjuN0V7fd4yz6q3n4MSU9X+ujEwscbN/uwcfvJtuYCsrW
RbCbz/LpvCoP/ipWbdW50BzfbA2P4ens71nidZXIg7JfrH524kEdkRJeO/Ysk+f/
AfZzqIilXkVohAoUEUZyCRgLTl3Ho/xbBVrY6rsAPhcqGVeJYBlDVl7O0EFQGA1d
XKR04paw26mZV1eihQWRRr+KioJ8OESNvwxmJYbL1kclq8GyD4722+prhxiOiQm8
V1zol6sycEMlevrhg8jdbBw44rs3TwOjeECgi4v9N+STxFbjD+GhwDohFTxFfo4P
iFwMDOvQfy4Gmn1qxqi4ZUYmLKu4cZSt/J0zKKVk2++1s74X3jFusqns8FMS5JKm
Xh9k4st3UK+I2sK42de+bbwQY5r2cQhyW4++njcg1TrXxolJeTf7/0jZ6mmfNPZ1
OP7a+fuJP2P5iDLpcAkz0S9ZGGUPRNslQTwgqvBGf9ezOvHZD0ptYetoLtfawVop
sVQsXDT5zDGqHjDRDtY0rIul0giITbbLlsgAAH6ihc0U5lSgJdh+RPpfsQKy/GG8
ZwbZQWejn8uIead0qW3XHCgp6vGM9lo7UzmdIQKAJNDf0fnVIi6TDtNg4BKV/LdD
LrbuQpRCtiPYFgOIjXPFcd8kDHnIBHKEWP8m5aL9HFCdwBCS5ukHU7aD4gQdba9p
UWEYg7qtz6JJOFmESxdVodyk1GokTCTVryUO5iOXpU91aJV4h/pm6kE3FMicsUwM
A7p2hXPKffaktN3UmuYT9KomyIO3av0IiuXXjVDVlQs6gm0EnfuHY1j2oMkWzsSi
OJCcIwt/dlOiOMCqJM60uCkihn1G5ZDLK3AJdKcYZkdv2Wopga0FwwFZ1DyVFgni
XygRx5hqXj6pTovlv8Md0UOdPCmDFPqrbCEKDFRwdZlX3MsT++alMq5l/b0G5ISN
m2KQlDUGOd4VmX2lxSLDNIrTx0CgnRb2HEcGhwxTjMFFwvnBPDq89LA/G7ww64br
vl4CunqAKGzN6C243QlDXM4N0fl6F1RArqqVsEE7scLRJOb+QlcUlOSOGwdmHFTz
+DVbhS4C0gTPk05VQEDw0FMXplsNE5fhYCZZFBXxOnpjP1ZgzfuT0mkiL5kFNuVI
gTePP0xwfO8VAtewxWIe0PIieyiDVAbr2GyLhk8SveLVkCThrTPmU1xhz27SKwqi
N/xZP3xDZMxiKqVMpa6MMnzV8lnM4+kVvdq5PHo8tfkZUo4ovd/oXlqw4sW9EnnE
uqqqdFlNFHPB8cz85JvbTHIn4QfRr3urOxCuqoL+XIq/fbmCJUlMrey7CGzLc6ti
VF+MG46JFotOCYi2uStdv09IcmJXaSyGsMiQILxllzzosYcdjEL9c+80EAGdPi/m
xd+BDR8T5dTystIDvoB3RxtkcIGhLL/p5GZ73oSgoiTcg4saGzUdTj6QzTIBCVHK
e+mIbtZq9z0MbilSl+mvEj/n+JrqSdKWbG/egKgTICBhUQBY20tNswJIWEnvA+Ou
KXdkLhqqcuPZw0jlDRn5YPq4btyd9zLYH9KGSWRutT6NU9WAo6ameI7LsLkPD+Rt
R3AHHUVPQX9JoaT9Ayoj1B+UBX4WwTYHUDnJROwfBElFs22CfTM1xNVjGEEXDrm7
gRVLn0nA+a45tDo7ev8csGxODQ1Am+qGEuNCU5zkMSBCvGJvjP9/N3q1v7FP0iCJ
OifSt7F2ChVaT3eiMD6ed/984Qcw9HqTvokzPmd58U3WUKJOkiCPI9sJa1TtphpT
uEl0YP/zxwPHtv2WDq+RnDJynKQjWMGndPgEF0aABRDmWMdcAl7OTQn+VQE4cHhT
kbPBOOTrJh15snRQPcuTRIKacygVCAM1aNSwEKgZNQvly0nCcQqPKzpqyjiO4kHU
EbovdpDMm+w4xorEHKdpph4PEjfH+ea0A+bhvNNBVoFkBAyjYbcdgD7YObLwBPJ0
jTGG4WIi1GG/dYPVHzkqxvShfCZUeu2zDlYZws02sudUBM1m4oSJGrP1NnTU+X95
eyoJ+V8EP/RSZkn/zHSAb46UFNqXyWsQdUH47eFm45IjvDIhifycSvwpqOIwKx3o
5h6qLTbkJJFwRzbxwd6TlmOayPyZEcpGJm0kI3l3uN+lz9uPW3h7ujoYKKrTiINS
jWl8z01wHdp3Vs8dMPHFJx6fQquDGo/aab9HU6wMBnEfqkg8mESaPjgqEUsGJLmm
Ce1qFmqt6p0BLHYUTFe+9coTGIawea8e2Y/jLKos5uQY215kaAHRPJ00TiFNSemG
fRVmWSIa4fc5VJC9nEOCavXr/ZouVHJGqiSVhpGISoeW3R2yPOilGc9P6QbSqLo7
b5DcH7SX9VSXF8fzTqZOy7pJ6e5+yoorqX3TN9x8hOTzKTJWi0LJytbbDWWvlfCT
MsSa3qgXyOY1lKCEfT807XQQFi7CrkfwShDmmYvb2FcsQX4DK6JuLFctZ0vuJ0Ox
K0Re4+kSqT379aE/MzdA6IfmsLfmrrKDrQBZRbeA1NmGc5oaZ0mn7wq5wRjrXMlb
CKckl7yj7PUBdGWV9cNfh8mAKBPWkc7JR92uWjUA/QRdTXCDmxxbi/zR9XipFk+/
buRaAQ2G5IsO+4YDbzxtRSh3eRmWg6KplFAIUQKC+df7NanwSmyEkyohCg9ezGPF
ls7ulZiFiimSvGT3/wpaW3WQWQ77uWmVpdKTOT3vKF7yhMn7Krq6sznFEJL/kSzq
9TRpirOp6YDdWDJxULoDuEbccs+PiRAhP1tRyI5FAfizuOeac8ajm5wcpuc5b7Lg
AUyOyUmyg+51hLN/UOOc+FB8tGc7v1h7LbbqrHU5Zngf267w5SK/pKIjs9a+7rwB
PQEgL3VIOvSeXKa0mjNOkFIx/pwnziOVea5kysdhDV/8LQlmkxOmx9r6W6lCAPOm
xTrH7u42ggwdN9lgoZLSXw1BS30t0/Ahj9/tjD1kx1MjkHStEsvssuiOaZSXvTlj
A1/mI63JfDt24i4N6bb10vKK10YsD4RxaDkhlf6WYTK5JVF/eZh1FPV2bet9dGul
cwWQG5JWFXogOS8utNgpnKW6kBIWLKLpCCoSEkqrkovTDIWGNV8GEVeTMil8Qtuw
Jori9mSGxpRO7HvJiCdn5YbnQQBB7Hu1WV+Obb8ntZZa5ZY6HPIB+F64qmwNJavZ
h+8skyO5RbJJ7fJtU/dXMsrYmabkkas1yAdJHSd1H/1uCDvUDp6uDGPEtVAFbOXy
ij3X3WLfLrFAVDD9d74kjFZP/2ZQprT340IDbQ7LqUITuGDhjeqwOYR2KTX4udPD
A96IKQGmEM6GOGPDfPpWBvoF6uGcs8GGXOzFe9J+bnJikFNFJxN30ReoaWyovbb8
eEeUBwpfSNAQBycWmgrpcR+I/jNbAFA42OOEkZuJ96cn9R81Db9jyTT9hoGcJp7j
0IE/c7EXuD+sefyIqvu+QYmAWqQpbK2K/QTj5esXMw0PiAl97s3nM01D6LtHTlMk
m9wJaiJoYsMVX47yYZn3b8x7MjwueuHSfMDqW3d+C3b2krVIi9Vd9VX4CwX2fFBS
ZpF5ha+si5hl3Rqek/nrJvO7uyaC8ntAEr6vM87fZFL6kou03Jh0C4+A1HfWHv8b
W6D+bAonTzK2IcVezx8AVss5G4TuuS9VOD+LnOfv/N45+AxdwrEu4birJS4eS1Bj
Xe/BiMvhNRBdw3eKMETe/aSIbEP/B3U0QHSR0/0tZfH0iPu8wO25k6oiS+iXyJC7
R6cGDsg0eFk4LRz5QPNB3L0m+VReIQUIi3W6AX3zjRs3rpPj7pwDV2//gHnVi4F+
5EBL3L4/OVYKK3m8OEUogt3xy/HToWAtth2pshp0usunmYTxijc7VY1FODUtlqUl
faTnSpYhxCri6JXYVbDk6GMi3PCPznNpE6mTAksJYYleB8dZjPwdnyNrRilPlb1J
FxHrLLQg4Fl1uQvnD5Ws17L+xeZ3y+Jv/QJuYyJdvyJLb/hcVErrPxioWF9pKOqd
DWc9bkhAuc+e1P+yTOzparwCDLbLNUAdBVvCNv9Q38injpPE8Tk3gYVx4c2CJesz
O89srSeLuRgFPASVJ51+CE5QfTrZCfNj9LLW761zoBkk6PXC1jng96f5ZFdXd8TC
O1fXlZIVv4+7CWdjwAG4H1pU6Xe7OhlaFqPWqSKanb4PZeM6RXO2wREtit9W8vzF
9HEAdaSnNaE0RmXmxsnCLdSIorYS6C3yrFJzYKWIVYSwJdp0HAzuyGnomwC5J1cK
oShkou4oJ0tKlUrZUIC8Hrnct/9cor2xKCRzoWzFzOD/H+KhkR8kh3Zjvo0u9lgy
tqHGSxsg8/GLadEMe9ujs0NdeQEp7qqwye7DE0jUOuIbyjPQLUfm7+McT22P82Q3
CGYmWxxPmIkrHj864dz5LstMhFVneCy2aJZwrUkBF904N1oU5Y1+9uMg3V/Au+tH
pkZttPVieT7PvmZfGHKyYqtRV3eeN7IZ+yxIdCGU9aXwE8/Trxn8vdSUPwwwBzQk
j7KzRJgTUFL5OiXjdjrw3JMmd8FZKhrJfPui725XaNCRSnLgeOrVvA1wyW6FwE4o
tjOm5dYk3D/wNemWa+ynH0HI/xWBJGqcjWMZoxJMXSiNEeoEqb9HrmTHPuXIKTg+
sBSezUDyfay2UiruIG3vMee1O3sL6ahvxhQKzIAE1hb7IfPDiRd6/ooCWkgpReJC
5nOei3qh0UOfTBZZ3rmv5dvNWysg1fBrSaHi/tgnm+AH+zX68kmfFhFaX8H4Qu64
2dldJyOravtv9bkEUcDVF1tLJ+yE2c3erwdbOlzQsUWNqRx4ABx9BvnlOzPEWPWv
7e3bZeMpS3Ngw10r/4dKX/lgp4/+GLvSe4DeGoBT6ZkdGH6tUzTxB1vL+nA/6LLe
IM2HbfpX09LmwbPmNfPhUbjfgEej6HBEsqXUjel2prYvMMbfxCE31WwVntNkyDLo
Q67QwZgZ3wU3KKlfu8HmDP4K8nZdfsGTjKc8CYZhEt0jcok3fAPVCY3Bbm/loCkb
wTtODoOOuldZn508SuylyF9Gqwx7RjMLr5HZ+7PJCtB06DyZBIgvzddbOlSXTMhf
f4d2vvQ7m/hdyDXTdo3mKshsySwgqzxr+Krp4KZge4NR+5lUQrQTGgQ0YaNKBBnN
0SccRcUxslgyA5h9zEhHxaAN2rqAtA9+8OEcpXdg5nFP3bFmNMk8WxEKiyKg6ppT
2+rymbp0SEYu1XJAx79eTx+6zAoBz+rvrT85K3DAvr74FFKAVnyLgZRasVAQDqY9
cYE51y0DDjHWXwm6Go+osS4fqpJ0+eJywLr1hrVk3tYAgMlKyMMSHSSOn8uQNzaJ
vJNp3XnxCsYiJj9chBfUGMSqKTKMHto2j+S3BC0alRbTQEv0RdjbMBWkABtz1BjZ
qVCTg8DFeZJeVl6WTpLmvrB2wd2GEhzFq0CvZim26HtZAyEBhJRPNGrzkBg09GQ2
uCHKR/0Wgwngxv8vtSoE389NHfxzdCXMB0m3Bv/1ZwyhBDnjAZNCx08suDrQhuMR
vIhKaNKeraPb09o6AMvSfeCCpWjSAr+r5jYMz7/m1ls=
`protect END_PROTECTED
