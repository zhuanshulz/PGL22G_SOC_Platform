`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2KtzW7sa2M1crC9M4HYl03X09wFcLr0EcHDWNXV6rlwps/cIT7dQE2Frrni3usi
Rdni1TOcTwQ4/DUwcCsc0Ng5bq5OJ+V+UqlkL471rXJWvPNMPTHCV40eGW1Xs4kZ
eAMIng/+yBMGFZa5cE8mo0PUBNdGlle+ufO5GcDuXeFxe1inug91xpZAQYH7TRln
7z8bOEEa4iCcIBqWYOQ5Zf6xoMG579WbMiZIfrkBvSbKIs1HI7UJ5PDAnAgv+MfT
+FgHYkT29HXAfczSA0m5F46w495XlKTQZ8cieDhUomIyn0AY9ylLFr3Vxl2Gy5WE
2Jf889b5wzGJODU1nXVy0Hmh3yB7OtYwV5KotV3dxm17073vR6An3WVxF9dYnkYZ
DsPfNHIug8hpJrsgGmrZxEJszRETXHIR6Vxo5MhoG7qyMjEYZicuD90l8HzS2UF2
YerWl3+/BUGu4Rq5vEs2SJ8aN8aojinjUA4dcCjm1vhCGOlYMnZQZpGDHoIIxkE6
rZ7+c6YW2aCm1Y1zYPK+NcIPhy0PJZdjhkQmS50Oy5IE4uNJapNkHnC2fdMv22iP
bTL8+Qbo7YhGxZUMEz/Zvg5I+xO6LWoFAAWX0NcOTVpJ8vi8E+YI1PQZSujrlGiT
S9c8oPD8wP5kOX+mTTv5qa9tjZ6LkNZLF8kUcrangYxyhBafsC4z6toBuBh9Egot
LMXxr8YEdmuB+fmUmxVecOWp0/NLmHOu+usOIUTpdkfhXex1KaWew+oS9bjw4FXo
AMr6aZGuyKuDmWZcA7He0UDa36aUU2+5/o0TiBTpidHofunqCXHSb8FR8xlH0D1M
tfRI+Wfc6Xy3luqIlK+PBqf3PjCzw/5sOjk9KE3ztMm8MC5IE8wQwYiswEDLdVFO
euSW40KNBoJkF9M10HuYEbvGAzBp/XCqMUdhcFR0XxdulwWnJDe8XmJX5gfCg1G5
VC6w2HpzH3tzv1QAz+zmB9xuEmr2do6ET2HrD2TcRWAgAZpYcGvg+3Voa/a+1SJD
+wwshTZsTYWt1B1e2U7fFjAvWlR5bBLTLCzekE+gHvw=
`protect END_PROTECTED
