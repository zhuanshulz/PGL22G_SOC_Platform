`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wThZqpFalb7lsOB1jxHsWVbVu5NpCDYTkaV64Ox9jYarHNZKfIXGz03bqt0YjTrl
dutrHK/gfGRJ/x1iM+90ED0mXQGbd8VnY/84rYTkO1PY9DQQ0ZST7xh0Us+HUPKj
cr8hiT3oh9ntk4Ov4AQZ+COT0GZ17jrwXHQHLZG0x7N8vWrBe0w6hwQRuz9GqDpj
V+sXh67+dh+fZeVBOrndxNtfOfFwg0S4Xh/ZzSCQ67sDSLDzi8LHrEbpdHmPErVJ
DEZ3KRFulLPNVSxlhFdawjDv7jFmk9l25J4JoHmQDO64wBDI0F4IES1SWe5djwwT
88QT9Gip0vUPCt8yiutQXZSs23kNlCliU1Q+j5dXanVFl8SXyudfiK8a+8V+x9l5
DQ9NCdDJcnyE62209/uTmSg0Gs3BW5bv3xe0NGhS2vS7V1IyvUURpsq4d7pTmCz4
R/PUyXyeJwxX/CeK5vtI0pOT0h02tr/gw3tgdy7isiTmbRJmffkNQDDnZf08KPYY
Pn4qczVTL0Ooec+5Y1s3Vg==
`protect END_PROTECTED
