`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nSz3ptnfi9XxuCHpnBZVE8uU9Sm8gSa5tvhXZm3GOTA8K45uqT5yYp4t+yP/4UCs
gLe5byrXhpr+YDNGlAyj541WtwU6twZJzU+AbgIBgvs3G07+dvYeWDfUxVSLkIgo
O43M3Ncw8mdyh98CHZFY2CrJWWn/X+RAy1kA30SlUYvDoZ9CgnZCrXYqoeBniA6Q
/+fG6EKCV+4SB6gQqXBsG7VNyol0fVpRSVJw4PbkBeqy3ue3nIfgo5faCw82QOrl
pBhIt+FBN6xytY1vjrzXVvxmdp+xHzZnu/+NXK4xWrkU9wzy5elZQa/Cyn19lDkY
MThxnkSJ+iWPgarDApzr3YHbdcEZDry8OhJwpdOEY7CgNgEcZlZmJzp2xM6okJaM
uME84HyCKrujS7+qfFGfqjrB/VnNPQKo+iUhzUxlByIPasiMu0IdCQ++mg3A3ma/
gswrvFTOFyoCZGfYOmWKvOAh83XQ5ylVNlHFtAleaDuLAHpnN7UAf7JF4Q+LrMlZ
EQWyEsgBa/h4Qr/zMjmWd0VBzltoJjlchkMpT+swtJTtG5fV95+GuoIk1TaLAp+5
5kfMP0PMSU5IHNxhj6SAylQN3nHDsUS3PKm4I8JEr3uEMOTosfI0LMGfM9EVqQj8
ObolX5McbYXeLAZg5I2YWVbZKNN9iNSGRvwEIHHmSEWjVo+HU6S//VBCVh7JKFEC
YZp0bhZewnD5pGH/4kf7iTIX/Btx+tqi3Wcu7KK4JiY8NreRvJUQKi5wDJBPn0mu
tLthOeylPTUUeXfKj4xPV+uiDYx9/pO7Msku0hEmIC1xEmY+QOM0SQ/4qA2qpnYv
0XkN5QnHRkqZAQDoFRaLRCwA577jhXrkncF9T/C/yF5++r1AZjg7/RrWYzekSpQn
iV0lQet93nMEeYePnhn3tdpWtuD9CEwOspmK90+cFUowFT+atl0FbGiIPGHxjLZN
xzWWPE00Npf4/rN/3+Y5V9UU+AQpO8X6ie1Y4v3epcogP6iTaoI4R0k3RYIS+8kG
jlpTHKsX9pg0vY16xucFuW8i2ZuEvfWywvf2OUyBUHKUwbJV1hQ1Hh9hXQ+hN/M/
k9rRdqsj/2WZB/ygecDIcGV+IIJ5yuAdKjP/k7O+ABr9d6fTn2tWPxUZUfGnZucW
5UT8QKW8Q6AlrDQQTQP0cmxjOGJB5GKm98l9jHm904URAfVwB/hFgxhGh3NeRI0M
oB1/QAIpiwJ5PTDMddru3BKbbUoToqxd0DKYwrPbwiSiC649d/FdHWNiDqvMVrfP
Y0vWEzq0Wz3kYFbwGis9I+C7TdkNrUVX8QKkCd4afPJ4/Ywh+AC7kJBP04T9YEhO
1DYecq+O2ZqwmmNKNFTg9oBj+5htjY5nL4UhLCUO+prcQRVu4vkzVbBhHioSfriX
8Vfvk5xQ57pWh/9xPLzH4p+eb5hY6sS6+V4XnOe5U0FeCDCMyhu4jv/nPodL6mUJ
nCL9zchjrhzH+G0OCd1bv9vwIzgt03bmvO3afRueCQlY+B3Y8KOCvPm1bdk61+LK
LVKm0pIglnqF1h4PEJD2TmaA90YhTaqFqgj6+jeMjLOBO9s0RoWmYyCi+SySztMB
q5TYnEImPx4Uuycx5+8DO60FXPP/oJdRHCYawsFm638=
`protect END_PROTECTED
