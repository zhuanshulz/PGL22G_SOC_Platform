`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOG4LIsF8Ybf6k8gH7KE+uTg83/a/28/TnMfXKI7ehCRC5ngwUqMckf59MsJmkjp
y/OoWDONSK7BDxf30i1dRogQFDdW3sPRJCrWj+G5Ne1tHgz+lGBLAQPmdDXOdBal
/6DoepNxUeyN22PXvdb1KqmVwToAYZbn9fzUqIw0Onb0uDYH/36RUcvnEet45765
zpnL6W96owc0oYaN5xwn76gXwuLqcD46z7AHZslM4u3Nau3Pv0feBeuycSHgt4s8
eRYKxmeIDqWSWT5LFhDg1wwHoQoprEwmklCMDcb04fQsKadKpZawHrxK/RhPxhcK
pMprrwnERg0z0k0MlBa/xT1PwghsvNaq2ConFkPXFzQweXgyv8Qn2UYkjkPrt3oN
mv7+s4qgxlvrREjmb90FDEzJSgY2OSSgNCtfrfMkBMm2MCgvyQi8BDN1IrYpYaW7
Zlxg/uasY7JEn0Eb5c9zg8JjYc+6ASisu9KgWjUZFEU=
`protect END_PROTECTED
