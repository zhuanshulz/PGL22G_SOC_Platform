`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlpaR4jhWmSWVp/U0AF89KGrE9ETyY/iaGmTW60RaQFjXiHh9SwxyGB+5frTw9J/
iLRjrIJqPgIKK6Nxf1dbZq6HXCdrgmJrxNUc9xNQ9rVQwC+X1cN7fXCsKTzw+les
9NUHnWrUGfMzepepVdWnwzIFZ2rG+CCmzWH3osQl+y39sU1UPY8Ip2+t8OR4svKy
whWVRPx4YPBGhKdkn6SRBRHEqw4J/D4vA4ytiMHqJPHMrJNNqKjZjLGguc3FMk1d
UY+W1fWzUEgNnis0oO3JHzfau5tAjcNVS0+EfeSdFnzChlYptmgitr0og6QMLH5D
/v6X3lSdLMa7/qLk7vD519kfoFzolzOzVstBnqUdukgzvg0NjnC4/Hgr0dxNL67V
OxVHwiZhwjQ78P4Wd/5cuL13feF/cjS8AEGoATOczgvbvi46LRmqjfYG2UYPGms6
oGqaZ2qaxwOS6fgQZARUQ/AlSddabTq7/Tm00eGX9O15sdnLrFJJxsSfJoSjsXOb
iq3fCyBXsbHsWhBZLp820rz90q0/I7OATVPVgGOPMoAJxllVIawbCFtXLhSutr0t
CTAErzksQtv/6J2V4JXAAVd1kL778qprOJLYf28OQVzfhrIjbcllseXetc1YR9rg
KgctSPBbr8Dh0JYlbrwnpNuKF5GEoLId3pn7RwmOs9oLIK/R7k25Dj1AvZC55Wf6
1S13a/6xlkDzzhCgPAwFJQHFe25oYml3fM8Er7f64YdeOpjpr4KV+Mjf3FfC29xu
7pYIf8KQJmk8aiCG8DmKcxCK2MMEBJtlGraTsjVkC2aoTUU+B53vqI7cvRIHLDEJ
4MXnIpftc9AaaJ7A8M/rGSI2guVsbjcuxXjzPGE4cmYs/o8zISQ4yzdtfbmIQdov
k8vdIAzwqO3xJDdZvKPdwIMAwRe+a4tmvcpI0rlWAMSBiIOomJ0pngfbnKOShrvr
RJUKpiuDCcfe4C2JS52Jl/CmGwRmpKzRQ9syqAQAYAKeceWCqJrg40PECncOH204
tUHDjVjOKsWNex9VyqvIOsmqq4XqR4Y9qGWUL0b3RNjRV85rTLbCaTKfg00zHjAm
hMZsB5lAdxurFrQL/l3mU5xplDh3xdoMsmJvaoXwq1Vu33mlKbrhLCDp5OY4jU24
69mz2RW8J/xKM0WC6QoQJlBlBymLicWqoUrnQezx6M4AFvsEoeS0nNwesCObsVpH
YJk0bVUXVkHTEFTCJMCa/cf8CHHIY+SbmZdJVAU2hvoFFUg6ykiX3xqLkqrZGVf8
zbDQFCqUER5QOWS5kJYv/oPwYnsePUCYJN/xgzl6WcgPn5qtAaD2M/2eNA7Y8RbJ
JF5pAzkeAhpEJWYApS5dY+9H5wZW/kFQVuY8M5xLHJ7BaHcKJw2ym3sBUCcze36v
fmfEaelXc3l83CSO4TFKd5rucsUsvd7OVoL7+b8ULS9++Q82hH2561OwHQ7wuqBh
OxLW+yhfjlUW9C1XyFzMrgKah+7OEo92m94k0/wAiO7JbvAMxHpIBEwxMwkm+51r
0RLzIflTp9SSW/Ns/bAkkww0JBW/B2rYqwAgRUAM3wYxseWD7kVHr3NOm74DgMKh
9pseb2lt51WzEmNvXAc+8HRAo1GCmafiwOO3NMc/H6qgTmE7v2Kg38qZubZYH86v
mzVs+5AVt8Pkq7EqbU8T2nsChRzDNPOmdWD/UkmNBGS2UcdOH1MeFhj5hqc9FBl1
MLDatNfR9OjAFYwcuVzyXrm0/uQE5YPZZymiXxJ5NHZduV0QS4jZI78DNX4yycbV
mSGPL4lwThJT/isLQMXXK6Fl9ZZe9e0ExHdJcTQKxD4ytbhIi1jKvqgWb6DQY7OD
n9QRIA6dX3u8bYJdbOyILmGXPGhvUBNt4+vdm4XTZxjBXVOVRYKcYrhW8MICbt4m
35skiMhhoFdQCTEqVmBxQGo17eQbcbrojCCZquGZHQ+n00lRevd8XR1mEBUgvU32
JpYxfn59/E8O4OvAJ3KP3dqk5ZjWlsmD5SchyAn9i1TMba2tRqvdcnXspGJ+uB5b
6Pd2z/RmebOqAF/LmlaaL8F/Vn/N3N07cpj+1evYM7FtaNO37mtjSxkRmcmBxjmL
okQK3rm5aIzKEuCqUhwDDlJBLAKRPOGdoqi5uOBaOXFffR3n+zGAhlkt/0n4Z8D3
0jrHLAahCal99oVvSpI23dpurX+e+sWD8c5pBnlu3hGuRUDwtvF84Olhs6J7fYGh
H7esAYI6cXduSAyHYVIIOraAfshEZs4NozlUY3Kk0xNEJdbDo6OXdhV+o7/N7b3L
n0nQBY1RdGm8HbbiTZ2NEZyRaHDWoKlvvLNmykISpzPYTTOOpOjmuLG1pLWaMfBG
EPB/IA5l7IlavLYEsD4eOo2FfVYDd0XNqdtQ2r/q0uQnrk1chzpse6zLPvtonZmz
EumuIr0QsxuksEFhkN0rLqLILQTLibCw0kTer8QZHZmnohjWbipj7G7JLFax40u8
VVlWPIkCBEqLclPViuFE7rcFDvlFSwXDKrcvmhl0sCuWXE17q+5/ZY/AkQb5hxKI
y8s4FPW1ZywpY0lfNGlg6w==
`protect END_PROTECTED
