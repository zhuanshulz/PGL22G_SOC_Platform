library verilog;
use verilog.vl_types.all;
entity GTP_ADC_E1 is
    generic(
        AVERAGE         : string  := "1";
        CALIB           : string  := "NONE";
        REFERENCE       : string  := "INTERNAL";
        CALIB_REFERENCE : string  := "INTERNAL";
        FULL_SWING      : string  := "0.5V";
        VCM             : string  := "0.8V";
        DIVIDER         : string  := "2";
        ADC_MODE        : string  := "DEFAULT";
        EVENT_DRIVE     : string  := "FALSE";
        ADC_MODE_1MSPS  : string  := "FALSE";
        CLKSWITCH       : string  := "FALSE";
        INTERNAL_VOL_SEL: string  := "VDD33";
        SINGLE_CH_SEL   : string  := "0";
        SINGLE_CH_IN    : string  := "SINGLE_END";
        SEQ_CH11_10_SEL : string  := "NONE";
        SEQ_CH9_8_SEL   : string  := "NONE";
        SEQ_CH7_6_SEL   : string  := "NONE";
        SEQ_CH5_4_SEL   : string  := "NONE";
        SEQ_CH3_2_SEL   : string  := "NONE";
        SEQ_CH1_0_SEL   : string  := "NONE";
        SEQ_CH11_10_IN  : string  := "SINGLE_END";
        SEQ_CH9_8_IN    : string  := "SINGLE_END";
        SEQ_CH7_6_IN    : string  := "SINGLE_END";
        SEQ_CH5_4_IN    : string  := "SINGLE_END";
        SEQ_CH3_2_IN    : string  := "SINGLE_END";
        SEQ_CH1_0_IN    : string  := "SINGLE_END";
        TEMP_SENSOR_HIGH: integer := 0;
        TEMP_SENSOR_LOW : integer := 0;
        ADC_EN_ENABLE   : string  := "FALSE"
    );
    port(
        VAUX            : in     vl_logic_vector(9 downto 0);
        VA              : in     vl_logic_vector(1 downto 0);
        RST_N           : in     vl_logic;
        LOADSC_N        : in     vl_logic;
        DCLK            : in     vl_logic;
        DEN             : in     vl_logic;
        DI              : in     vl_logic_vector(15 downto 0);
        DWE             : in     vl_logic;
        DADDR           : in     vl_logic_vector(7 downto 0);
        CONVST          : in     vl_logic;
        ADC_EN          : in     vl_logic;
        DBUSY           : out    vl_logic;
        DO              : out    vl_logic_vector(15 downto 0);
        DRDY            : out    vl_logic;
        DMODIFIED       : out    vl_logic;
        LOGIC_DONE      : out    vl_logic;
        OVER_TEMP       : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of AVERAGE : constant is 1;
    attribute mti_svvh_generic_type of CALIB : constant is 1;
    attribute mti_svvh_generic_type of REFERENCE : constant is 1;
    attribute mti_svvh_generic_type of CALIB_REFERENCE : constant is 1;
    attribute mti_svvh_generic_type of FULL_SWING : constant is 1;
    attribute mti_svvh_generic_type of VCM : constant is 1;
    attribute mti_svvh_generic_type of DIVIDER : constant is 1;
    attribute mti_svvh_generic_type of ADC_MODE : constant is 1;
    attribute mti_svvh_generic_type of EVENT_DRIVE : constant is 1;
    attribute mti_svvh_generic_type of ADC_MODE_1MSPS : constant is 1;
    attribute mti_svvh_generic_type of CLKSWITCH : constant is 1;
    attribute mti_svvh_generic_type of INTERNAL_VOL_SEL : constant is 1;
    attribute mti_svvh_generic_type of SINGLE_CH_SEL : constant is 1;
    attribute mti_svvh_generic_type of SINGLE_CH_IN : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH11_10_SEL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH9_8_SEL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH7_6_SEL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH5_4_SEL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH3_2_SEL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH1_0_SEL : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH11_10_IN : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH9_8_IN : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH7_6_IN : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH5_4_IN : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH3_2_IN : constant is 1;
    attribute mti_svvh_generic_type of SEQ_CH1_0_IN : constant is 1;
    attribute mti_svvh_generic_type of TEMP_SENSOR_HIGH : constant is 2;
    attribute mti_svvh_generic_type of TEMP_SENSOR_LOW : constant is 2;
    attribute mti_svvh_generic_type of ADC_EN_ENABLE : constant is 1;
end GTP_ADC_E1;
