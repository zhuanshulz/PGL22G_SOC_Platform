`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbuirJuaVhTDjB6av7Rg4AmUvgQY7Pe0FTrvfpfaknU3978wy6ZdHiDk5gBhPNXj
8kW74KBid9H/MHcTO+coVXSMn4L3AeK8UXD1Psg99PVQDTBGluQU9/noXAzBv7In
gkHd2uanlAhBBBfhWgO5nrfpSe/zR75rgARMp9NZJzbrraj8MsSuovKTXqSrw3X0
9ceIupaBumxqtboLI2p/pti5xcupiAqSiuEH+Ml1TZ8Ln209Hr7NV0dom2tYx7r5
uUsjmMp0gWu3bOgPOnJM19HIVvz5KcFEsbh6wQv61r/SDBcg9m2RwscUOVioL+C+
rYlPpPkVAhW9vdwlbfU262aUhSYnuu6dW0BVAecFJFj5595puKEKZQZ/jVniom1m
vkCFpZ71N6ByAeEyfD5n9Cr+5gamqXWcZCUPz1pEJdUzSoasBP+xyP1HMIM/V94J
Mc8IKgv4IzRbaDCfvjhyS/1B85Qy/3e8OgM/5EZ9AZgKMYQS9CN0AUWUAdaDhtE6
OvWC0VzmVNYIHPGgst3K2VLsCYEstOiVAsnKkatQ2Wd9iYR/QVnHIrNRjXNp539n
KsSjgqSi2jCXxj9XBEVRFk2YrfrSIrXR56OOUxt/g2HnPcChX9RRElG/CpcNroQR
455J14BzUo46E/nYnw8IsgCZtUQI+l7fKOrmKQJZ5iLakjNVi8EbHORVWl/aaftd
8PYpLcJGoTPQgfnMKr6NGQk+N7I760s7AS43z6csuXwe2U4Ax6GZpqXxHBl4OtBs
aNfjjQ7GUkyLPF2WXRbYZayYLqULZZdwEoCp4BfCvnDBVOxgbey3+gpjbmkD+UPB
trJtDbsFTl960dpyltSTD4ydXkI3s+iujVhrg33IannBVA9ZI2T20MPpo9MOu/Lc
mMgN7AwRLP7K0hyLoGOLTYooywSjL+5d0yU9Xs1u52MbXBN63YUNqdlqKRGWkN+4
UXKMA89xC3gVjZST12T7npXRsCd0+IUSKJTHNWigh6oXSyz4bwx4XkaKU2kza+RY
d5/sjawK3KZgKQ/hDtVMIvjGerarhHKNPJqSCweXJ/Hd6sr+N7c9qJoMuoXzMBtn
LfwXDNbYahQJxg8f6qVhCyP+uRmLSuMG0C4j91rx4PdItJzssW/aTbbNIvB5Dejl
WPMbjm+X1YEEJ/pMMhHpZWETFMX2EE94rEhPooAZhfRi1ws22Ah9ohJ6cmjHXVEj
jqwB73PUDBTlZqlzfVnNXCsu05Mcoh4J3IwEKZ1fMAhLKnSrX3yBt3jccaqksHaf
ok4FI/IGpG5/OtplnSw/Kirt6d9mc/fIrhTEeNfsAu9Zd27qRoDIJq3vZxDLO9wW
2cXL8yK561esYPRtBsuGYjxzp0w8UZDClBcpAAF00DZuCirqbajDo0JgtUDOx0kk
XmvpvXzWng4SiS9Oy3RboWbDCxy1bom7nubPsTohWvMBWwKTh5TuGoHGAb3eMDLc
Mh/6L/2S1Jrz5WgTvllsezN9xPxwHi1Yw71TQ8uIfoawwRN/3cd3fxXYCc//WBd7
weS7uyat3jCivcg8LnyNa/x4hTEDjWJQLY1/QBfCEI2dznF+ygmbmb1gt5XyWZ4r
1dwoJACpm7wZcj9cMAYo58CiSxrNlNtCDTEiKrDeWeOmo0KlomKkg/VQjOD9GwDK
LM/czw8pBYcEmKeJ2LLWlBTx8lP2gAW0aS4PrRy4xXWZzWFEg+ddaItT0rElRlG0
ZcJxw7ABL3G9LAVnyfUxYqCvzjjxmf9LKvUisvYjI1wbo6Dgi5cCubaznVw0GgQt
ikyhOzEWVBvxzzXR3WJZX6ptgRLIBZ727rz5JWuWFWMMtFevGqXYnG1x5r8Mp2qo
isnVIafcnQW0P9xDwkrRmwWQKjwPyhg2Ym7e9oGnmLu/LMyg5A4TT/Y0Ay0Lk5sa
A5iJdmdj4RsBYscdD5phj8xorQARiVSsnBS9v/O/bKY4GkEvcRCRmo5/iNqieisf
CiCYIXNNdzqK5KENGrGKvapw1yu3vPhAMmr+xvL0YhyGNj8uzpyMtYK4iys+NTep
46r36MktFM1keQkmgC8GI7HWY7wC91WQXFfuKpe0EwMzWe3+6X/xgURtdD3rgMYP
DOe12NB0F8KrlH3iwIiGtuiJYF+Fqekes/zQGJ9RbxfyZHqcwahbbCoBvC6yyVsy
Fhsklw37vhXT068nwbWX98HgNr7L5VQtiFN1v/MzhwRI7iyhulH7RnJM1ZSl0sE4
48vnbmdCDZd4phQe2Xv8o/K8QR1jFrp1uoOKCygKlhC16pKiMKsv1TJ2UVPBKmli
SitiVFCJMVZIX3jvZfXgRhDELV+Dnal7YgXc4VYYA8tOqWaIhVc932egc9lPmsLc
23Kv3Yb+KJms1bpYNwLoxcASaYNwUdaIdcxL0yJJbj7cBBkdn+iWL6CgpQkKnhAf
PvIGGlB6+xkvrYR0KfSPI1Gl4L+wEPXC1zxTQAWZ5z+m7qlGxty5zB9gUCdB38nX
nG11s5+HpNybEB0xWueL6xG3IGOYBdjrq4+lvJk4iRXMh2ERf06wZ6VdRkbYeD/+
zTBbJRhvuFGP6sxsJiuw/+CdlTUYv/x/OhfauWkGn6SdxyE/zaTjyRDmmd5ix7vv
eJ1c4bgYHfYA3pL5iqEH1FtpxOzMyhhvmszzodMfkhOIu1uUkYP9BupVPsGiNdTi
Xm5dms8WOyQjsICYMsKfu2gOtHAG8YaJWEQRUpf2sB4P3uoG9NoAQSYIE48akfF6
X+zQsnzLkc6k/lNSZMbvrbodW4kL6BeCheml8MatKKJA5XCiiy1BseQWa73dQlL7
LNAE1+6r8u12e5vGS8ijaxfUpoe1YPUBW6hEz/Fb+jRlNXA5VrTXLw+8W6vpFI/M
gwfYw4qOP7qmk6yaDAG76YKlmI+is1PHaKtdvNLKTdY0mb/8lFsLlvIeZheQ2WIO
5WaEFmQMkOv/VWfst8IUUUOEDHZ0TgN7Hj9R5xje88FXxgvkL7Av41QDaMBqCZjt
i1JVmPqhQTiumrQPI4iYDK8npVQeEvUi7oo7KVW4jlTu+qsLyakQOcWxRH8mXYyd
5tZtg47kLtx7C9+1LBuVkNYezC45j/3bn2M/IRKvizSIrFuaknkaA0uY7K+hplgL
gItONCjVvsfB6Bsh8noRZitJAgGCyWn6DwELGGeUsEf/vPR/kyPCvsLVLK6VC+9X
bro4hTBmaj6SaHHOTA9okWUwH4smk8tC0sNJo3vfa42F6pd7ah5iL0+cJpHa/4rt
Cjxl8rSq/2/7hwrJLZgy5YCrJ8e5vEendJcakGVMcU726+WNKsBNFY+dAIiFxWb4
vE8YMtgvWqj54JYSj9pcTrAnHSlNB5GiOJy9QEOy/KDOjxTvB+siXsi+etNhM5Mj
QRklqkZJLiOeSG/zFgEiaFDKYXI2/7VvK11+MBwr7t1Qf5eyHh/5D6Ab5lrYJHhr
D+wUwGpMfrM0O3H+iP7VsU4OXk1YaY0s6Y4USe+ddW3vGeIl8DG7R/J+P+1vQG3h
bTZF5a5dcHzxge8MPxhpFJwPijoP4GdPvYkbSfS9zL+KAKyqLMKeRVxaPWKIwMfB
1E8N4P3NKUizHhzSMt1sdIqx29/k2+tIBu09zqVKAhUDFRzrs1X1e6otRombdoXx
tiIzhZCA9m2QBWRZ6HKpGV/B9uvceZx0vjyfb6i4uTxg7VUHwe1n3hQqGYnQGbB+
unhuco0Hkj4BFYXDXc7C56z6Hj19G0bT6XQlA6D2mjcVZ5qOd8tVnh7UYxU4jKDD
naoKYd3HvFelbVkGXTBpX5pv8k+WKw2BU3kbpEh4JLsG5kQVAriNkyVPqc42CFVc
X+/QAtdwlUMXBaIEUFo6StYnakdTzWc759Ws2mzEjlhGj60D24xyhTigJFLYaMLU
DRPixLBoQi8CarMJPPPAHDSJ5ZB5fRl2P+6Cf/F8FktTxUGD9eTulWuMSyr9xBUP
HRCZkqxr6kzroLPTrfXAuLgyCQZyVoqV6spFR4yAR5BO6LkhlSE6kUPaQw4CeyaM
87pvrgHGWflEMjC3ICTrcZQFP02o3c6NKIjgVR7z4BazYyMxKN0FkyeGOwbyqnen
+mQeWP1Qu9sQX+crxap3jRsC4pwLsYaPRROIzDHyzWB+oVKm7xQLYbqxQQAQD3Uu
G1IV6L3POHChL7+bhz5wo/klID4QW/2JT5CPxKrG1olUII408ZQS260eI01fdiER
KRYniKD8mjt1+syC5XLoQ5VcJ38d2mUvicvAaxt1g0X21hA7uR+p7rWIrwiYOb6O
qDZFyYJwWCj2ogkRpfktqut353ZmYkAECVpvZ+fk/auO32Yt7pXI2vsi/wWxPAPH
XuSucJ64rNiT/MtWlioGGfcqIcs08Z7dQnV9PYbw5kX6CU3QkOyO9yc/bquEq7HF
+bRyyl09PpCFWK0mt8l/EOjU2ojq5cBJ1jFILxDxF2h80GVlJ2tz6IjdOw2Z5oCT
rtnGUrV6hXskEOvSrSyARcIXY+1BbI8naJC0jkSoAxYP0U226XYDgGpwlRT6AUyQ
gEKGr1Q5MtQYeNviJyG8FUl27bDr1qUhX2QwopILUKj2AFa9lvRsFay9PZ8xgOR9
hor6iZXAK91l7f6mm1+QfFY1sDup+/pylOIh9Z6vqpezpZPBBFlfBI6z2+UmLqPn
aim3Vw0ut/AACfvlQ+9HJHzxZVM4X1ah3hrEoorLP+XJV9EwtIzeyZljQS/LNEoE
MvW8Ghg+3If05ncaRvZkGyQ4WisQbtHeoT3QwxVbMRB9JZT6jQa2pEc9XizlCIo1
StcdnRLu/3ceZDdcsJY2Hf4C3KVFYQgaAj9dM0f670kWwm1/tyb+4RHc+pu6tal9
7rcLfse56t5KNIYzbhe2jGMDVB300Szd7SUujKOXfViR/UlmyB07e2CqhEhbgNfh
6VlSlxkRhdQ95vrGoddbnfpdR6aD8LhN6cD5Ohxh7TNNMkVzeLERol32tDCnF1cB
oyRXjsLqOaBc1HqrU0zMaQka1lstDi9SSK8kv0Y5R3XSM1gFKoI06i4XZ/G7LIyC
W7ipmrrqIOITi4koxU5GJXuR//Y2KClTK58iaVxR8aSIAWZHA7+7lNzdVKRO3lZB
1DPPd2NlhX0nNITFcg7NCKO13p/OyA5BYgZC1qycCM9xkEG70kKN4s8Zb5gG0y+I
N5u8O4Ozpj+t/I8BLzRi4+NOYGIcAkxM9ec+Pe1wKDAhja8n6/9CwizxXTFrVvcD
IoRm42t856TzjOmjcW8kCiZQaSV8LojD202Lgfr4V3LdPLS8myvIugRvAwzZdins
W40YsKWgpT/D1Wt28QdsMVrJVrijoN8zsvUFivtqwg7syJq0rCwoSYb7Y2bowgyH
TJX9Rdmypt8TxzFLAu5zFnnxkwntrdg+ZNjvZrfOTUk6wAHlC1luk3conZFVtrGf
hXa5E8JncmrMxDDYbC7n6EV0c4HBi6ucgQgyjPb/beV6iZC38evtht3R05GR6a4f
SrKaqaC4UazABP6k4Jy1kFMe0fDqlwKE+QFE9Bqqro50VQY+lxlbapr+iWksBydv
zrq1JLHEJzDmNOXBkDB441OH9BPY0r87Ob/ka6mpeWmpjC7Eu3L4OTjTXy5jKiWo
e9JOpYVxosd+g9RdrWZtzUSIOWnnmScMIk3A0sXmjDEkRWqw4DCqSzeM+IwLijLB
alb/V8b6u4fsXYD6Rs8jO9AqVCcpsdN1PzUlpPeHE9iKhG3dHck70VrWc9aUruEb
Me65gMeGgxWEeJC1awpGz7PMDXOD+UJ3fxx55inzPcIUdxZO2sAW5mYecWcFowZ6
JUbJsg5fLFW9sWklCqiPHuJiL2B6RbX81iaygP2tlndOSCtafPvBb8HOqR2CzrKd
goBjuugSMHKWQ11ILVDbrT0zyY4G/BYZaK+x159SKD0whlSkGtnHRqTmLtez6rsm
6BDQ3dCOeqwbAGsxDZt20RHrZI+fjcihjUv7+lWAnS7XwJTulL2thI+ift3+sQBC
+D6NtvG+5Chlwg2eL5O/nYhgeGM274UoTX0kg88IUq9dCQ7zwW6ecHbBjdn2IFuh
Q3VhveQ2danrfRzQrlYIsbudQH1ye3UTM44goQgEATrPBl/FyyIn0wY19jcLFK6X
oktGDOVPvE2FanxOvtsZuFDU3NlRRcZqxBrVQw+QKnai9TtJr/eco5zY1ZxgrPO5
2DKAf4/Gr9MXh/uLfQsT6K2FHQPrmXXHlLE4TFIrUwROr0CUT5WFQIE7LeIpN9bG
4i9LqaQAexQo3BocyMufTBxn/b5+KsHgIfQpXdFH/LmOSnSMWLxsvbFI+lxWSaMn
MBLWqg5pa/tTVa3cuUAUT6No9hPzvqzIvlQQah+ScjSOjEgCSqcFwVCVGu64sdVe
4ydeAeHVn/NzKcQxbNK5/iCONuF57jT6IpIXZtxCt7vKBU2oNpNruJbRAoLDg1Hz
5wyL6FUalMvDpq1r5UbQDzjbS+VXPddoR7G0Mf8cmCs03tY0QFD1iOsBXjQECeD0
qV5bN+nID5im83q5oJMjYmvxuR4wcRGXfOrc71WAu6dSxa7afneDn/6/Jqn0UFfw
AEoVpCSU4O1Wx2TRd369GYhSp4TKjGtB2I2BHhRmX1ShrTCDNUZ81f2igjR2jvLq
HtFqDo3GWAYMIui4WphitV8pHtosSDpkImzDGdf+CRv0Kqam1r8dooNHfMU62nM1
2H/gYTnWPcsEVt4AiSFEj+GwMy5uZkggvux/qoF1NO+6O3UKVYSTEHdykTyyV6YB
rgn3RUS7KQhhZ/NlMXosrPpRZfnhbbWPfyU44RUQ4ayn9ncuEj7ZtjLbEG0k6YKk
L+f0ddhVd/WsBmBmGAKlTYg/uXNh9yYye5bWGb++SDMtu2+4FfJlbKtFLVjXq2J1
ItaL4Hih3SfVU43NweYltql85UjH6S4uC9aP8kYOeHeKL+bqJcP2NcQCl1bGEn1/
oFe6Ud7GVtDvI48X877W5SvCY57WBi5DkUddyshdNy/w0jbQMlUuAd7I5V6w0M+X
Xx1PvaQWwxXDLEqB0294wF6ZZONW3FaHO59ioWoLBdANs+k84mxUmscvLx3Ngymi
HK+Cqu1v/9jRVgN0gpc/aNwKKNeTilD2C+9+R8eWjXLM3ArQiEf0y47lQuGuckCw
KnS9PbTJhpCFF4Y2QxUFbc7kSbYPuP/e35PvU1GcMYFknGNwOlO6Qz6nv/BYYGGk
H/lQk2gv/o+bm5DHddTM8sWfvkNOTYw/Q0+8VhRTsB0mR/LC3/tPHcNIjr8dRRRC
u089NnpzDxnwzWyLRuq9DTFcPyMpKEN050Ga1fhE3EUtNZoozIG0q1A9enUxsoRe
CEOhWv2J0jQBUFeH7aDo5KLrFezWvLuTMPT6fH/w0DhkflNLE5ItpB/bVFLE1R3l
T7VA4EWLOrzUrp9xMs9516FEd0fPFCN2OjtI+MoWWxRjK9DVkQg9LF/Ty0i4ZOVb
t9lhkcitz5jK6XvGZUmo1zEsi8eKYNo9bdOA3lEz1XeN6K6GDH/lCBAu8AkTYAsr
CkmYSe7USF8l9NXaLcvx0x5/UvpVx7MWdnIuQP/BW027Zjqvj3u6c5686m0e1iIf
HvvGjORAxbVv0sPUqnIPNIBqcGITKPkkiTW27asXOqExi3X5pHvA+5T95jzjJAsp
Kw0arve20FmV1joaEvcfFR+J3QAnJK4jEVM7/cGW2UXq2qY4UCVMc1c1EmMzwDEw
EMPMx2yxVtYjxQEYGb0/CCXP9kSyobDBxICGm8uxk/FSkxsI8CWc7QgQP4fXED2Q
L2o6v5UC0SwRE2Eeq1n1yHHaS3q7AEMqhtzu02Yc5w4oSagFOwiWLZqYsuOFrlvG
oVV+x6dh7dmEJmOZNKH5xBUkhNd9KzCiwWclQ0rV/OTKNl0SyhGDIOypYG4i0+cB
M3lS1FQNEZeoFIIGMarrvkTO2JkU+lwKub8n2fzTpUTqOoWUlGQo74Opjr9mrM2N
cS4hU3bAAG9Eix3wQ9QHLDvtBx8GB0wbVU1WvXDkTKtYpkk4yK6OPRSpxY9QKx9E
js8Hdpv8EwQmABdEnMDRX5ycmisuZYKxgZgVw8ys9lDsB8KGfeInL9Mt3tu5rPN1
RzvNaRNXqj0HtuUduS6BfVCm1R2wlWqKSbB63aG85fzlxhOuUUrn7W0ojNVnkUX1
emGrCZkLpAEjEeG53pV6Y7ZCUVVpOhaPbwR+hDr1nJviY13/evtgCStVNl60M/Nz
QrixVwPRXpaDy8Tc88noFVFO6nJMlTsyBZcPqNDnZXtlqQt2QUONIxv/gDszmIJc
MNCS/zxfb3QdeZ71xk2WrzaDmHb9yzzLm6zZxbEsRV+RPpSboqEJMiJ79nmtFV0l
/fR3C5k0448O5DSU3xHjXqCU9hHD7aJfggEEpDRyZ24sbE8p/0Fo10g9B3urW3LZ
ebaBs5ovfWrLu9vyWJ/DEgKJ9LoRO6JE0RGq1XnAGeNbcad4ctB8mS4Ski1kQdM+
LB+3wc54N4bFdVXJKdtb6NQSESCvfkVactsoyLhRxt0DPGwnRSCCLB91nnRM+RBY
UnGv3WiBE3yKbApgrRZDiC18UUTYaoWctZltI2iW7Ggr1YNLfg1iVD8Zw9llEjok
2ePub19TITzj4wTjXePl8UkPbd9HXx8sEMpSxCWKZ3ag5SZymrBY5s1Gwqj6ZKRY
ofC0InFLrelCmczngMdKXnPEpyIpxOmGWBvxDO9NYAh+73mscmVrFKYKJXtTVDUo
Zs2aL2TEaGk0cQmL+OlzaZWoFeCn9mF1b9/NaRAej5Stx4+W4tV2A8Owmzt0r3xD
U91n2C39LpShow7/dvCup7atcZM9l3QRQ7oqoPKn0J2ozKQ5SrpuPjLp96dHmUce
uOE9BtijafpGHpg50IdVnb+QaH4GJKegxZoTD5tGGDzOjrK2CXfGrzGjVyN//u0P
pp0zvaJQztwJ4fppTEvtE//tKPS2AYHPo5ZFIp6OkZ3kDsmFWbmRKO6xqZAJYo9X
nRe1fWEwgUGxBOMHcb1qmosKsCQrCCfWeOPvml94lPeqP0rdLdiPzBW0QkjmL8u5
Cw6OSouC5tWSVm7bIVed5rlEfoM6yjmfDN9d+26+yvsAbdjLPEYLz7xhgN75u9Gb
YDWieOqyIQCHGx//Nt6Y1JkNgGf1+h9sf9yuXfTiqxg8nlgXsWVoXiz48KaxL12a
p1fLHk99Gy7HQIpMrP73VJlCLsZM4VAmN5ryLX/TYU5MYnKZp70F8PiRTVO9zqvs
/S8zWJoUFM2yJS+zpFXsa9xSS0pf7RmBJLVv1E4fOLk=
`protect END_PROTECTED
