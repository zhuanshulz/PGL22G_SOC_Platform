`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQ5Vo9PDDSDLlXo6o5X7nElMYbTwsP9wWMR5mFZ+m3/XPHXvnq/mnN17QlN3fzwr
zcyu+QftWLdZQYHjDX4Ow0sf3y8iNVaOkEo3IkX1O5BVH/JPEpJCMIl8kV2Rd8+u
I1JZRuPm2TNfZ/xvq5AJY9F/tTX2/vAqMjuLJ7b4rV8N5VnJBTrTOkXXFjW2BQK7
IJCO66A4La0hDEMsQtsEQYv52ZPW+wa3AmyxdsEQGFusxIN9xlXsI8fPY+oUJ692
A+TKSqht66WhVJ3FIxeLk7edoW+vCRTn7XP+lAgz2dVkjv0gHNsR2Fbp8oHXgn+G
rOJ2hpvd/uv30Fc5/3CGBB7STvKtrA0O4u74zp2VW+v3yFp1ZiX2fjMx5ixVOuOL
smZWPqoJQBi1OTzYFQ2Yau82tjSIWw8STb44gGszcUiev1lTjatRg7IQFUi6KGZy
RwURJZTBznETXNiZ7yzIsuI6knGL7xDUK4S0x9Ntjb8KtpWtC2M7P+7DMlGJ7HXB
B3qGIk2R4s3yw6jJ6mIVqLIWsYJuielUMFSXRSnzZp3aPWKtYPGHgcCOEgP+MO7R
l7zj1OCa0iLewZcKl1JlxDoSGz9DsZLIrDCI46Eap0t5h2/E3lsxZwKsB1gHMVh9
3si0dzr6rinJNz6LBLB9tdCJvjHDS017BvGUVN0XrrMOzcLdlIFKWqv74kcuZr3U
uh7T59KB1DNeFcRG9REidOWVv+vkf/t/nZDb62zkmHE8mdrhrq1MfjwMO0l9uRBQ
fAYShGhRAxHueJ4FYwK1xolHsA0u/R0uQNntstkvljA1bEV0XCNzVt/W+KVf2G+5
zlZxvB0Q2kqCAEE1CzTshJp56p+yLLTo0YJYfyJ2nYs7LB+vgge8jRXVWmFZAwN8
S5X7MYuERqVKl8ZI3sf4c0z2jLhaJvmrVhK628KsCUCteVLFz6KomSKIygmSu6ed
Ty2wVXs14PCX3RcfQ6nRI7sj1OEPuSlTfLjsWvjMzE2nB+7U5tCLSSAJVql0ZMTM
Kng25NkXal/VK2MOcTA1S2azztrhMF51x+IIRmzSHWmeBrQ4pYSUz+AMCU0ch/Yb
YGEbPOGGIhnS4No6cTOCCe+cM6Zxi8ia2EHT6gOJcyDQJ+hvChwOml4ECD8NJ1n2
fbAQNSrqH8pzbenTClnkwddnCrlJ8OtGbLoa6nus3AofUUEO+aHz0NfUzO85JzOq
RFlD31NVRycgvfS3Xa5lmy5EeoTDn/vGU8iNJxAm+J8MR4kvseE4uRBvsGM0G9qG
LZxEGspJ95CrAuc5iO+1r0rKu45dB0a5MVPL4JjYK75YweujizD6tPbntahEtA7n
K4dXAws64EsJcV0UVxkYFZPEM6LhYnacLDbbBlbN335qO1Tku2GMy93lG9glbUDf
3MCp8S4YekhN4BEuNgHKg/dXPNYgSnYa0qY5T9VaxUZ9U2P0tYNV57yug4rvdLj0
eWXUG8iJDO/A9NFzP8B3fyNkgEjpNacnXHyrO7z8284OvfN3HY7rGx/AlqpKvVQJ
G5d/RABZFgQ9uTbXPbKJm2PBpnfjYfrG6XTxDwrP3ndZIgi7pFE2Upv48Hfd8W3C
beONhn9crv2kOTfeQQNMWOBxeYP4SznNDb6EjXqkRmLtrMk+V8HNz9e0K4O94Pzm
i40hB9C3vWJJqHbTAKHraEimuz4GhPMMm1NnHZhHrEj+VXnSK2mHTuAVSBY6Rm1/
lgyGyBtkVbybqOXiS3cD/cfAyiJbSvO2cn2bSvdQ/PENr3TNuidqgGlMzfpDu9i2
adewSrEwKKRnn2kr7dRRc4PmeFyS6f0Hg6cFCzoNC3Gvog+BR+ZZvNNZeo5NqecX
IKtR9ll6WLXPNrhO0fiCxA==
`protect END_PROTECTED
