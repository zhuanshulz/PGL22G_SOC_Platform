`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ehwRoiNxQ2XC8ES5dmJyGSBf5Tr0ITrvQ2HcHcjjVXsrAaDTOItBN+YDy2jno8qT
ibhMZMfLxfelBdxI/ufNt5BnfuoU6mrS/v+TAuJFDCHk4SH+Aat9JwHlNMWYM3qO
775cbAGhdZNy8y9Bj6utQz3u+4F/UNGOkH8f9uE79RrQgFw5pFaRCHhNA/vZY2aQ
XTA/relg354jXMJkM2v7W0vxikbllJQ+1F8OgFnvTaNCK4QkrjkFDCo0GtR7Golc
yCnBjR9OciGXTSkl0wBSdwot/idHuN3t6ECv/J8t2F46wiJP2Hv5RlhoSxNj2f52
b4C8ofqPDvxGH4dU9G3I+0xprILQlayEJ5sWLvSMDC+XVvnRBfRummafSD9x/GWF
+cw7CJPh1YWFXkBDs7dxAtWo3JfVDJoogx/DRAB9tMnpdcUk//FId33a3wrWph5+
zEVCM8vsya0BfB8lnmPXig==
`protect END_PROTECTED
