`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CchQElm6z+FCvkx3wFa6dTEP5RbaCAXb5czbiEkBRWZd98CQKh0e92kctQKkfToG
djRCOTWUJ0c0qjBgqKya+z27DutQcsgyFto36/NZnwTjX3Z7eoSXeMLxEv+dZYiE
knsPLCx0pspX0rjUCvMEl1XfO4S4LuWwDtPyAdZtOdu71cHzRjazYFAjP1jKICsg
EVht+cjwDdspf3nBb3jScgTTHklmHrXZ/TCAoC4ZjThUNz0/Edma+MaJd4UY7NjI
o2DXRqsQoOHGdN3vCN3g1IYpmPId6RPDaVbUgZia+dHyjxGUpbgeaBuiAMlPkGqd
lehnDOMGOeQvP/1u6KdjIbdlsowl3T2LbgLfTl79tOYJksXB5leBwx1UYMhxU+l1
vJleOLSm2LXwNGk6NhaojIf1Do9GG3ybfeMP9CCYFYdxmprosxLUn4b1JVzgzwWF
T9wqMxKg/hqUL/dyTO6pFGSNLXC9zjxIueXBNAp25FlNwMnrnEGKXo7Ve7hqUUpL
ztbisrwct2txeF3NSv79jMAWepz8+3TwdBDg88NgWhJEPM4RQmcS7SvU+/WPG5Yg
FsL3lBc31kw0qZhHoBwAzSi4BmZpl8LJDuv1Jjw3w29w4Xv60UPou8rFLNtorSWx
ggiL5G8RTajN3+od7XEvVFsEUqBnKT1N5ilqcln6l9X43zlNzVk+VZ6+hjIzcnSd
Z44/KMq8c05ZnHVoFialIv9DZdUAKwl7mURW184zl4gBjGpQAECQKxPTNV96ZraZ
8netjDYSH3SXUJG1oLw7YzOgXh8M8FZK95yLmEoxX08xi4Oly4e9lGg4nx+Yu3rw
LMJAJCmWKQf9SQAGaAg+xoymZ4HYe+KWSwZPx68kYWEDvHkau/hzLJBvabnX0cOy
07weUzxJCi4oVDo1SJ18Cyq9cyoSv8VHq6A9jGXtVXlOaAvaLqI0BeHdWBsoWIKV
U9D1ihDKUP5Yy+vBnqAKASgrHKujE6egZspmm9hfPJc5tL9GcWMrrbRROUW6YKq7
9TWLF5U0HLt40zrkAxxZ75VnNoHFJu/UmcIsl+4N2kiZnz3AuaLsbntz6hf6ZabO
6R98k+ni9ur5ZsFsTaTPw3jCopnVENEtVvTCqLOrhhlZrEO/82FYBPahzMKHUlQj
VtzBWwuutNzsvhsXvJNNk5VjzGwFsXymfp+/ZCqLbTd6FZQpFt/yuasB7gWd1poK
YDLzfQ2nijjIIv/eAJlXKt7DK9uQ4MNGRv+GmmiCAc/vGas3LjmtzcoqUnKdGMjG
VDX3943Bewmtxm4yGiaeERIgEu/0CJQ1zmt4ws5r1ZV0CQI/AXFPfKzeMlZuRrT6
VroHJV7t3P1BnMhEIuQaWFRKnrBqT0JPWSUK5+OCelhrF9suA8bPTRv8jNQcf6jb
qJFoGZASSn/TrzG5E+rM2zB8PRxzDAio/CVeeLGNXRcxAH5fVgetcj9OhIVWWrCO
8t9h6ssOogGXA7V0GP/Mq5XHYjVXqyx+b1qpMgMCOiQ=
`protect END_PROTECTED
