`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tz9UqCFfJPTEQyiNd829WFXuJLpdpXw5guwnaNbmU2iZ7tlq07QMbNG4I8bbxrdL
gJ7nBWbWmrVeZ47ur71ZSvkhcTNZYLoIhbkqS44SqkRmQdC/TTuAOufl1SjDOirw
itoltonfeerRcAmoRSO/yaGUKFtvHb2fnvFdjnkuF3fPkz4aOQCljnKQeRUAouXj
2nOmslZpfmwBsG4Th0uiullElSVGHBOS6t9DMWIMMaRrr9jeGzSc5cnlRl2PHIDH
eRqSQRFN0w0+/iDh+BL6tpDP4h+dKTL5RH9o0qRXuAp30CGH4x50VI15Wr27/99i
ja2TLGKi9UVjCDXYI5+7DYX5F2Px3PzOO3D5rg4p1esdhIXh1uhjXV8tmGr6YdzA
cCRScYC8md4ZjgtpjG2fJIebXJXYkhCH9e+53Imb656+pWG+iBe6sfhEt1WCwaD6
6pWvTKhwnIjqAlfP8zFJTrvOaIbFfvvSzizQ1sBkuMRg8SoKwPDTTaXMbAP2RAyw
y+GxX/JIrpKNhq8Rs7TLqYi3+EMTXg9aJV3Rf9iCQB9DmkndBlWduR2nL9U+f5LT
tVFshoJG1giiUepQBmhJUbICcn2biG2YDwAT8kWgpt9mSO8p3N+bOMVuae62UJbl
SRZ/wZ9oG862CzPnzydsOarM/RU8LWMImp4iYdvDfdEpOkcZ9e0eme77omzIjEEe
lnSGgMiaUGlu1oxkd/PPLbpxldM0Ah1epAbsWlLlBS52C+iFYK5ONYqIL5GvFEMP
FwwuvK+foRlO/4ZLgvMEHkFKjHBGr0r8qx0R7dup278XrVAFZXYzdM8RzVjOt5lS
prOjaQYrFLhq1EkxEknTz8tSHTU6PAQmVdTQrHx1dvIL1VhfCr92pPtc/O13Q2bA
+GfvBz6gclB8TuF+Nl5VMuuv76oEOH9Ih6BML+EuPVLNKHiwprpQ5Q0ajhvPvIjj
woEvYh1jkrUGMT28B6RBhqozwWwm2CmeacTM3zbhf4ppLkMXeTrYHCMqVatefDK6
Ak/RzqyORcXZW1a3iaeaf9xsrB53Yvf3V2GjWe3urda53fi+6umeVbsusXzFFENL
Xp+q2skLROUG6ftiX5ZmB7QPzPXjFtVmcl54tni9FmhzF+mw2d6HmHo7qKAJJoOq
afNf8MKE0QJCWMSXGJHJzeliBGNu2dBCadPasCDhLnMBzz6OI+OoMqWOBBpDEkRq
+reA+xTq7yw4G6WL/9j2UEYKEJ2t7yNZ7B/dp+W+rCmEo53J2xTQMI29Lq6C8Vu9
V8E0+FBCSaUFuRA73n17RyQ0ep6sQUg5yPMlVX5o6HK3jkswukPZp8aOZCG4USS/
9LRCI5cGGQT+HElO9BaJuEVD/jnw2HBXexCNUvoVBP0J7J+3ebiPyKduVCVpOb5E
nAt0Yd9OYYLJ57x/raoncZ6rkmVp02LulKcBjeBgHaQHY+dT/ml1ApnSILqNGHdC
c2NhPFO6o/b32n+4XM0kujY61LBDA7hUYfoLRwIpfN4AWtFpHxn9FGCuLOl2RDup
/f8DnrUmKrwMZVGcwET5D/oC144CbXayxvkyU4l/mv8Q+zyoVhBfA6URoWeeeP0n
5/ySyr4iBerrvQ7GV4+xtgVWTtPfU41UX6Uytb4qP+oa32wr9UXzd3C/PT4UBjgn
e4S/WXF/nlhwRJ2HMu7Y61Hq9MyzLBsToYMkKeLYJGBix6Thjoq7t906obyDPy0L
ljnq9LsxbSfa6zKN4y/VMn5QOrBJjJRLng3NfD9WOKYV6UykICRfKPd+6DRbh+ZV
aGckPW/bp5mpSEmmv4EJ1xKn8KwiLsUzdY25o7WaKv2+UNZl9CSxFVq05M25s3f+
+ndgtFnYGEo9vmDQc3U+3unwep2G4qzgzL+PoqhctuS3flGtgHmGl1PPjvbF1t9i
Jx0KIM4xPZzMCWmYX0u9PTFOJnxaBwGj7FlzVMjI2Z1eJjGJcQAruWow3oU0oguu
IBvSVizlijhZcNiC1nZjVhPkM/dREAoM+FGvxL40t04PvjkaXzkIbAt4SxPm/G1b
fGDAFtlervwrYuz3khB9BLm0PxV42jYsdqHvpqPS4nBMTShfKrcr85+bDQm9Acwn
DrMfFaGhOHgkjaZiQU8JRIgKwnIm5PhaWqwwq2Ay7bDJLHXhT24u25uhZkPWLk/D
kI9w+cbBUdtwUlGKZ9hTdGVpcUsPXaEiyYR0tUrVFS4Wg/icDXm/F2ovm1JJveq7
wvbdHNdes961tqKzVSbsdB8LCzqnSDD+RV+ROpiYIYlD4jNVo6Tsh/FDXGxiiOPh
+/lBGoVWP0zwSO9Ahuj9tLU1chx3cqswj5ty56i1EvurKfiEVGu1TySOcyo/joMx
0GeOFj8/xOskCU0cSDZ6iXoQH5IYJeEDCIBfNflyLYIVqM+TixHR+qb1sAFWIWib
yoRU3XrEWREJ3CaraN+uckPqd4dGbUYwp/cZyGmCLjwkGG4pzwqharFqsc7uS9dL
jw9So1/qZu7vVvbS69FC8MeEwjHfgw/kvbrv6H0dzS2TvORZt8HkmGt6FV+fOOHH
2rzsn3d5k3SQ8MA4HmANTravqpDNRXikNRA+Rxzoo/wWd8eajbLkuCkuq6nq/+ps
P+33VNS3cSLp1PfMco5Kn8KgZjDRpyfX8bKJwykZ1I62SD36hWgxzNQ5N+MMqXcL
YmPwOs7grXCaicSOdpowNZSYslbLHffJsw/UiQWd2FjXeM2IAJnagtBc+LQ96+Gx
VHtW+pBNmC4f8ojk98+To86fITS8FoOLSRf5CJt9CcwjDhiUGMhxrmBey2mEJuUh
9qIw98I9w9XqX9jiQPZXUMzkYpGpaPImOsIk+ycHYt0q/QqYzZ9nnInqhRgYBkol
IvtbKH70y3iqjFxeTOk8cTGljSRmDgWq2AERtoRFgD5rdI6vLwySwL3A5izxWFi8
q8ya62TTF0K0Tt5YkJhgtVYxtge2jVx0lWc1ZyLnmyxbFyT4ncm3nbxbhabVwzAe
qcE7k/8ow7VHYWOA4a41OgzTeXBL55GtTZtlRcWAIuxhoWchPlYiPBI95e3uQSsG
Lq5GGFA54EHgTsyZAwVJt9EGMwiYkiLMuU4HukG5mN1bFvRT8YwZOGVQJ4CLFpxi
ZzVsy4R/zTOx6//DeSg3eTpq60ZO0A6UVz7VuGSTmXOqgFdIO5iL4zlGZRwpcupm
i+TZVnO06ZIUKE0P0wWR/FsW0jymWbsnovKg22jAtkWv5RMB5GkdHDHXU5/b0rtu
`protect END_PROTECTED
