`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YavbtAfENuZCqqTqmo20Jgpt/kyfQDmR7U0QmUWUprHXijQbAhVZWM4HRoWJRwAt
l4xWYAJvENxWhTtkq7xiUViJ8rOkyv8Dtq6Y7FtEB9CrWQMnJryJUqhXVWLGcnNA
rPwQlh2cSXPAijoJYz98PiStu77ej37A1v3UeROGO/gNEEfDnk19/MNCuECDACx0
WUOA79ZwR1dIDVLtwYsoQ18nq/k33M4u7CgU5LyAeg4x+8GHXqjMXCFJ/fE44lKg
K3F8ie4Sh/C3CZPX3AhtXxZUM6x4xnb+TDTjTSR5OpfmlGRka0O405EPlYd6yWAr
YHPH9PSSaIjsgVYu//2Z83LI3h9KjP5qKRQHDAtmbEovADNfN0xqzzImFB4o97US
G9dx4YgNz19amEzkFEORUvgBGBfFArdw2XUVYsQQJxkfxy8bXtOd0xQ76AUOMxYf
O7AZTKSeDRwATKASuLtvK8vHpS6pDsQJKs0z6ktT92hlT3gAgGVw04nibLk053vT
r8zi3gZwgMpM65hzkQUK276iA1IEoWJig9cqaFum9LDXuLnA3ek16ACl5HH5kh1i
feDcKcX8Ol2X3/vTnblesGththzdfs5M/YRRoFaSMwC5JhL8kwagnhJAkSVuf9bF
NoS8ITg6Nk7SUHOxIh8erBvuUQ9rqEpxGSsJUP6Fb90kdAJCwTKoMj5TNCuYsoqH
VO+UP74JZRYaY0p4eSTG1XG8UP4EN3iYKZZ3le6z7OHUG9JL/Yd1ugQbzSYaFayI
W9YDyhUyM6yofD4MljyUf/l2y1d9qgzPiL+aRilJHcMjWoTNe0kwaQGQdSKres64
rsGKI21FRU1kB01FxDFBiyXTJUmpL/amOrL0U/XQM5z/xmzwJVDIPeJDJzGO44JY
ZticwfwMi4PFk4dFQnpFBaZLesOy4QJ8f3JdXV837Kxv0Ewx89W2AUWg1dfMlcOb
0HoAhkvhMDyHXl04S+0Auca1a8GyKg4pmYrqz1zduZSiZGKizj68ZAhJ6fCrdYY4
M0RW6YAtSZr3ZhGcj0AsqyxSsNlaCX3vD+UsPQzjspDDzd5/OkfVGuQp/Ly+dsx0
tPAA5sFxok03wO/tv5fXkfvSiC3ywzgRY2m5t+Qgy1VpbN3uACkyHnmVC+P71ioa
SNj6iLNO3vvwq2uDwqSN2+L0fxOzgmKxJi5BaJgASTUcnsFBVi/qc46VSH2XT/RR
Onjz+/Ex1q9lqimVBikWH1pkqXFs0Gmx6t3mzWMKW+2LoMUU6f0URuCbhHFGgeOF
gaussHTqVAmkt3Mi6eLGWltiakx66BuAPDpRfPxCB6Q=
`protect END_PROTECTED
