`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gd0ImRJYQMRs3CLwbNkSGY3L+XkMzig8NqqZYrve2jeAWfxFP+kAEcCMG7Mcns1h
5ymQvI6AkkhBLQmjm7uA4Z+J4sij9mr0oMozO8yxHZPiv4cFUTk8iOrRM3zirCnj
xB5a9jCvDVoIT787fZhqYi99TaPfxxoTmoTuKwHDg/9BibYdTkELAxt3QBWLzH6k
3tpCNo+X7uuYetbEdyJ6eL59kRPhRwhHDfOg6K6MO7GdMh2mm04TmxCPGGqpGjMl
yz1XCCASERdwvxYpW0qvBt7J0Fq11ADo9qezKegjyuV5kL45Rto+a5fbga8Epm5b
weT8hvb6Y8u75kHw2sTu+VnQxz7RFxk1w2lT45UsT16Kj0DZOu9AGEbYFd5/C0+p
NZHRC5mlxigWki4ofJaAG0FLSvRmdJT3sIScUmImG72kGafPosLv8ci5TpYAw+hd
WdpR1MM3b4XJmpk2eZHzZLgg3k2LcUCUKVuqqGBnB/FDULJhS+A0X0YMm4VdURxJ
vsbuZMEOkeYSM1yphlMwVAR3icDlEzF2eD2FmUXuPNKQpbg7uoAbfUzB3fWZy/HO
Wh3Jndd5Bs9POMeLgZwszw==
`protect END_PROTECTED
