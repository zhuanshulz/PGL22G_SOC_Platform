`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dX2g3FGhqvBL8LRpLkRKgqGwvrJ3v8mtBPJw1+tb7JeQgowFPSjpPvGsigraadBp
clTL5filT6f8RVFafr907frAT/y7sSzna+CmgtoZAPNf5uRiQeRxJoJ82/hQYXyB
uJj/6xDVS4CMhGHMzXsHUfnFkjIZyidDAmZACn5uv6GQJJBLapE+bmI/w4r91uRu
GczJQEL55KnvS0fJHSEJbkoe4Q4GIdFil0S1Nnpk4n2b3NYI+JCfEoRhu3497r+c
VoyRqnJILqkQmAxgcvPnKd3FXEk8w4TcPWcpeOUzpWwX8LgxHW4m1Oe6cvqIeEMt
pGudP3mFaz3GhnfMuItcbmC+D+eK/NhnoiowBahgs40fwNz3EfMZbZ97019Du4KJ
8pcQajf4r276QJvRCIKaUQ==
`protect END_PROTECTED
