`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yO69J/3UcW6h/DCwdM6mocOzjU+kUXiMjWOq3VKikE/ButOzelVrVoMQJi+ioLFw
OMxG/DicExsgDivi09csc4oaHx+3djuJ+FxSIb5fwrcr/2sx77jMSU6+YyzqdfoB
K9g/zJeofAtIQzMQrU6oqkjEz3psPsVfflS8O2OxtEsaFvdFfWSU6/RDBaCMUp1M
BtscmjkY7JjbX8WBGBsNjbt3kLZEHKvcbz+1BD3nDbMWiR3hxaZWC3kDwiSuKFQo
HBTfonI8UnFwLCJI5pM9FOO+kTClfhT2sgXFqvZzeXrOwnQB5AQqqgpRvLvdF7cr
ivX3s8OsrZ3zZND6xanL7XxS46PYHYYyt4MoTtHjd7JgXuYuyx0Jsl0l2ZFcKznp
9d2cxVGeajM87dVu/Cj8XmrVSekWB3R/1iBKcti3Xn6T2dzNVHBVRiTIXkKSu603
YCtjg5ujr/7f1a4a6CmWL5jtO4W/Io2nmjXFA4JUDCuij3DgMaVza6FuSB7GlAan
liNJeyFn+qE4W9SgRh90F1dsswgjUshs4WW2dtTAcKmwe2qN29q9zq5g2rfSl9zF
9QKoGUYZDaWMybNPLn+IExJDaik3P19VCYKHJvVR/P5kzSWh0viUhPKqw8IN7QoV
NRisB6eK/WKFbmM/xSmBslXD+D4csQUceXgwllbMPKP3RFF14XtBXXor1ZctwWbY
83wL7tgG6JUXSqdFHcw0/1kd0RBbNDnhi/lH0CBdhsUV7XRHoYD4CZjYXzr61dEq
UrR/0Khqb+zrb35uAoLDpbcWCQhz7ahsrdSEB5YIMUw3A5fDgrvdpMCXntRE1AZ+
8t0+SwfDWRyY2UrWpl92BktnN3e/uC8VHoCq3v+pgFDN7u5+8NA6PxBSjWZFlzAa
aLsAh6QMIqn4zMDvR6De4DnS+4uGGJfuzIl7pEJjzLh1xoBxl/XvWkzWMhQ29T9I
bvW4z1d6jI4LW/d21NTiCY8XgldGrbms3JhJBubE4nVy0+IRncZ0xxwHyW6y/0W1
d61D9DJChAT06p3sX1St3K2Q655qOxGQDf5mplnAlihIkS0T4DiyBNxmcyNDSCmy
m+ONOpp3V7Kq0Nv2EgxXKTB6qQwJpgMuzsJpUvVfKCuI6dSmen8PyacGRQKjKarf
YsvskkyZPLIYtmPfoJF4eeK0rpREOqaMIeB1X1SxGXUNoQFVEuMIVKG+2NtDOxAh
Wma1tMqEXpcT7QQnagEpP2wkU7eyP7dnsNyzUlQrVHvRQKSdGfIBOEwQLEVjtWtq
/KoCIII/M8D4dX7FZVYC5bJLzeUwvXhTc2SlNFmtfw4jhRkpCV9CoVawqWYfjpyx
tfOO8s3YIWLGPwza3XJ5uJGI4xDB2BdTbhZWlUBUkeevzgCn3NRtfkUpfken1FpH
nK8FAV+6xSv3Y0lizzRZFyHW1hhK0nQSG2CHRkTf8weqwza9fP9nYu+hE2PcikLQ
VrTXwczgRHQN3iJMZCag+HJA86QREcVHOLDwnOe3IcUKpflQbeWbONTvvLLau5vO
B0MD80zSdM1AnHgYXyk8d3skqHwKzJxyFpcijMjLeR5QVqL2EvtSO941UmeQax7T
u582smCjldsEdzHEuG5CMXItFmvEwSJHMY+YlEfgb4EbPm4WPSu6OzBSQes0Z0FW
c7AH6Q/h7Q4bvCWLlsqjsbPWQGnFGmGtwCTL2a4j27rPJgQwBDlN4SWaO6LlhymR
FY+UOjkj2r0C9MKR1+AM6U2h/I56amcDecA19xUxOeDYaMHZeSsVaHDEyqRP3kwi
CzNKPGaX7xeC6WaohPnGOFek7VlaEAnjKHCwCkVzGJo9QEMRaohpYdxI1kc1COd9
O5xBFQKivYn/m8kEa/JmEyjiPiGMQfOgMnOILhEi+tyajRYw7JKuWLE+uwZJ7/x2
QXLE253SaILSoFQHnqJRed+ySWon5+/DLDjerofCSZnMPRPPC9I99GiLiTzuZZq9
7ID2W+C0hxknX+GpSw1BkW+Dl65Wpu6ZQsgmStH3Oblrmq385ofq8GfeB6jbYAZg
Y+mE+1+eFzDe26O2i8VtV5zPLKqmGGf6mGbERcWgddHd6oVM249sCJLvtF8bRnkA
nogz9H0syBsTroT+B054WmdM3UZ6M1b5XLcKngu15vu7/n5wyRdezU6FCyvEsxF/
qB2O8Rbkfilv+3pD9YFXI3nZ/bP8Nk/9295hj/hjyqirNgJ2lWj6Vmsh08NCxNqK
bAJl6CKOYSJ+7a9pZd4bVWCs1azTno91AV9tVLsf5pimtvVCkxbdkn4vCnr/o+eM
7M+UCLUjPEM6/AljvgbVHFapP8qxv2PH/tUKlKpj9hxDeQltDJghjpIGEh2ZFxYJ
rllqBYK7M+uPatadyWSboferRTkGx0qooeBPpX20pikuAydznbrCgaVo+JRsYkxs
RpEhn9uFSCqiHYKaW+y2e0NoTWXm+ZhxxD09whc3ttsiFB6YNO3a7PN6b9dKicno
8B+oOCI6enXBnVoFuExdTPgO/r0u6VTkx9HecY8W2XJeM0TtJ7U4/YZcuLA3OVOz
krHRSgQsmdIVFwXyuio/WJRpPkiMz+rpFo6Apro6Zc8Q9J2Oa0rp3e114/GEnCuV
at0Aka0YoTGk4mCMbNmpuP5/1dp6jA2q2ByPjmjODIBGt+9MIwtvzK8VToHb2WFF
F0FLyLP/PrcgWlQ+gKRPzdKBtgzbSqREENrLiwBks5BqkYjq2Cf9U+/T3fe+NNXg
3tOdRR1aKOmjjSPxX+N2EfA4CJen22mqh3IN7Fgl8eYvyN/0bmLlMIq1McJL20WW
6mPVilqwAkajnWGYttWVDahW4RT4GfV1c7FQ64vdlk4xv1oXFYdR65ErooqO/u42
LOyRnUp1JIbzEyccDYS4Fqg/dduQ0uDvvpGOkp3mdo525PH1nPxlhXeCaw5QJmHL
ZKrGx3Jtam77Xu1UGzm9brMh3RfrDx8IQFAbwevqS4+w9TKPNCFX0/MlLZpfwRsL
NEBkU+bc6QKNdOH4ALNh/CEUKmHkEgUQplJnsBvTxyTJEMjeqoSh24xDvwDZ+5Jj
UhEJeB30lGqsSOzxLRuwxvZv93R97C6Wfu0IhtP8CQNdliuncvhigv80QTE1gykQ
sJ9pbtAu6odsySM+926sRhXB0wiV3RXartVlQet2JVJUi+e9JKTYFt+5qZM05g9K
1R1afTzFATTWcdxhEbjMXbt6HXYmZRcIQwpUqpIPDk7DBx+YYH9A1uPA6stEupbx
mnUSJ2sn5WZMesG/VvJdOd0dtRTMvdV1p8IsNuO+a4UkPdtua349wheCIqhcXzit
3F8YrZL26bc/41ce2lhflDkCJdsM+p8VmXyhbwIa8P0C9AcDeEJ5xq7d7J6JNiR6
hUyvl8P7Q4RMnVMJHghrjb9NnEHFt8jw1VRGHNn7XNRR8sRsh/yji62d0s3iNV96
/YLvB9M/RpYNPAJDst4BWQ8AQ7cpWei0kyvsICHLtEcMejxYln84FqUBKu4E8EwX
dyyiDwa9iH3Sftf4oCCoIl1+ZbksL+7DFBzHTNkiRP98OzhzwLt8Vddi2zuY9AMG
BdEknd8zNf/SWz2YOXfZ7L4SgiXv1549mfe3+/+2rTeZj/0kX5icNhx482Qee85k
SLt1+jePuMKXMxunka72jTH0hCbfd3HNod5QZcJ9M+zrBpNbdrtalrxzxl/v/409
qF7PCDzjpDU2WtMcpuszXCnqEQHRrQ+H+by76GvTqCF9c4hOl/kBbJXpv5KQHZgW
EWONnhvUxZ/3JbJ50CEmX19WFvD3nS0fb1au10XWm/ldwFyuhK0dhk6l6pZcEDCV
ZOWhbAENaSAJDx/MTohq4wC70wRgB+vojPYMmwwT9YQAdzMmc4GlrHYoBw3fgw7m
LiiSV1uY86Lv8Uq7wHMFY2eA1CgvkDjx/GjC5N7lGvtdrPK0Fb1R3skOBgmYQ3YD
XxDzaLTTLEc3f29wvwIiTDK1K6B4n4/n0mRb9mUJJfsbVnhUK5LgUN40Max5EK1Y
Y0SKrcoemV5cKLlr5dnTBVsh70Vfb4vSkARgEDSBIO8ir2y7wh5nr1yuMzOSYDp4
lAqB5IpLCf/ioUL81QN2n+asOOyte8N6el30UMz/fXtXQdml6AWfsdjhQepOHMfX
kKTy+IOBe3ZBke/Aq2WViapIfXf4/CUO/qsN5rXQ1xjXfvBzee8SMYg6D3T4X0DI
bwD6Ib8gdd/n1hHDTkm7v/cFL2rlO4sP3NyhrAU7h6u63biKyfCYba215noX3L9p
eWii0Xr/jXsLEcaq3Ld9mxfq3Q3DRYzRys07l8rHmLtg4xAIgQGPsYZMXVACJUwX
BkaQ3e9lA0BscX1epzrZz7zZlh1F3cQnZuzrmS3uNCGk9qaHBQDG5osjz9zJ5fzm
yJWvMFGgU5dGkSjnVeVddY3djTX83UP3EVvUvRz3Au92452BjiHLaXrB38aRJffs
eC9B5+bb4tIHfEff8/K30sSaRR03eQQFUpsqP/Ekx4BRfGsQNMsG2moJsW+z7Xgr
RguR49aBv0tCIAZAfu60+vVvHg6Zrjh9E2UdiMKtKrJToOvJ2y7JnksJi8JFzaeE
hnuQbFzqyg0Hf0hV3Pr+sAEvThMIZKGstXj6zaEN+gU1GtBlLW7vI8N1f8quOjEK
LDH/zcW0Hy5zke/Fr18whVEO4D4edIaB4cy5n77evIjYiYI8VX09PP9Dk4YT0wT4
hX7hEQOvlPrUouu3EOHUuhEoniR3cxC33dYRPzjZ96iA0ubltyH+VrCazhiUzs6G
PJtxACIOk3WQfh1iAL9atdWdkTDb6KueiZUngABvwrtchF4JGMaUt7x/fBj6Sq7e
Bd7604D26VIhKZOtecPmfqDLlXzf3zGYhJC6ytBdDFZ8aVsgMbNSLnsXlLWEFGBz
ROS0kL8bV+/G7oEQuZ/hPCYeDoZM9N8NW04xBOpd7O0k7JQTLnbkmZqKQlYEq5Gc
y5I7+jLmmfGHjh+qV27ENm5XqjXXjtzCHqDTDdJZbFW7K8mX7FQAs6uROPefU/O6
6t6CT0aSyIOl9zxC9Yxy6KMOS0n2FLAgmhC7uZPPG5hjKMC15sVf15o9jWt9iIT5
cQbMzW1UYghyFbPo5EkAv+Vmg1CN8OlAyYDXWih+pn+2hy4LYITsXJgcfV1JZroG
J5ZYvidAM/asQxE8M/ViSdqzyY6n0D3QrkQZMZzzrCygyLRkbAGnlw3dQK1gwWgQ
ns0W0iAQyg7kMdMIdY6I9cnl79kvCYYY+dxkaW6cw5EdJyPOh07AuQjZjXpPm20j
6au6Y+kAS8dOZ+9mIwQoU/fyFcoNIucHVIrGWFIeu3hEvJOjbT8hV8FqPMOthdO2
iPJb5iKBGHBWGGnbIbuVQnTKv4+yL2qTYzHvTVFtyHg3lNen2Xd4J6B6rrhqzNak
tFwEv4821Nfpomm1TbY4LRaEe6v3fx9lWS+LbAOs+Cz0Nr9Uy1tCY1CFXYueOz5C
sfFFJD25Zdra75eqGIlRpX3++h01LuQoYrdUQFqOFMTr8YC5cv3YPAhpz3mFtFbn
Noz5dEgDAE56bo+0TVC59gLrYtjcX8L1kjPPEw+0U7/oZI7vAD34EmIFoUcm34QF
+lKflBsdN/PR7pD7ednEflR3ALiv0392XTnE485UdUn+9Y6wBsezkyaS5AEDJHQz
+mfeJ6GsjkAWLps2qNRkOISo4Q9ytqC0Rrwr1O/E280CXz/Qi10RM9jM1Y0++ZFc
ybTGmg7WxOiTRhc5liXdYmO88mRp7Tlz7IIJxm23AmevjNNCE5cRJ05oh5XrDnLJ
QSaNWz+rBwAA1AuvobzlD4WAk14tG6Lrf2wTfFHUiLj3rZAacC02XtbVn6Fvzc6Q
K/6EFsqGWkNOSldPrOuheZ+U8onoWHebaD5xh4GwnqPN8p6z208zyzWyAH0QPcvs
pOkFQw2rYyZmMZTJqoG6vowq1u2YNJSejOLmofo86+wjcwsKKGw/rDpRx50WH6Ko
o/o7wzWJszAxtrkXrlfmDCKswEkqJx8IqWxoonVsd71QyG+HYgKTda8Ih/AlBuwm
1Z5PqzD5tOtzxxGUkCwJCFpXgigayCKO76shqnLdPhKbvfNZrTKx8ROr8GOqZsee
oSTywNPOKdI9HNKslzEu4apNYAUhLk2hGDkf2GONsjckuamCfA/wtUEyCb0AKNMP
vTrqxi7A4H414Ep5EGK7hG0mFHcqf1nN0lOzTmmCM/uBcE+4CT/qyHqOqx1yLkyq
oFKy10TRHs4yuV4bzOCC+w==
`protect END_PROTECTED
