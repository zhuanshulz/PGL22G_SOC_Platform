`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkqZy2G2aag9xwnwCWXdrIkI9+D2HaUoXJYkQgDJkWUESK5Ts3luHK5w3Vat4aNn
0XhhsYK4t62Z3sqTasDpX7fjbP/YwSIADJwrUAdo45HDNT3tSGcS6MdUSS9oStOB
ETPJPe75eOk55JPIAZiwzwPRhd4hsE9dMEuIwqpV8QFSmoUq85OE6IK4ZVPAOVti
+0mUTuEyMH5h+UwV90REDYCaA0y9iFYpM+jI2CVbwLss1uRy2yhUwE4Jt4jIpHun
UOWDa32/D20ZdkMtYKYN7K2boY6suSx1yYvRSr17efRCsMhDki5UaIZdueqZQSoG
M4TAiBeElrsn1pUecT4UXypI3hr0NEWkx4+d3j99MMaZusXvThPpgFz6S6jsjoeg
7E2EfgpCUH6E8Rvy98idQIADuje57bPV53N4lRUz5FD/np19rsInWV+3nycbjDvb
s2+98+FDnP0uiJVkI650JQE1rJ/kofFJ7+qs6zdMIG1Fp7mvICkKIyKzElUZ9y9c
iNn9LVD6a1H5THTB+1i+PQ==
`protect END_PROTECTED
