`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+YvaYRFpic1L3oM4Wm+SBc8xPuI2Oa4g5DbRkQwwZAhIm1fdmYBMCTyz3V8xb3F+
Hs1sOxH1MMMNRoK8NDEJ35L0e+vzQqS2L+e4WY99WR/NSQ8htWZpLfnuo7Uj8HIr
F23rTtylzw664yru1QmoBny9nyHDP+bjpDiDwFRYmAov++N0ix6O4LrkdJqbGg9W
DvmDly/02lTk0lmXTCSi1lRVI7/c8FaQ5j1fRQ+OpiJZiorpDexRfdVVAWn9ScA4
aXReGamfg9UdCFkCnMg8p8wYUu5BmMvAoW0JiNAugEfTENQ46BvSOVDt8LeAAl6G
yXypY0VBATd3FqVFLWb9IoW7nmXRrqSHjpVZKsZKZ/+eH98C46lmOZtz9SvSDE0U
NNLZyz9p6m1tSWmldegbnk4j5EpSX7/c49tRwQBmAh/Oz10WKTIGvw1muuzWpULS
zzmymZqXan8XR4LOP1rcHCr4zTUZPnLdmr7ohSOnxZCmlXe5afmR7nfJTyn0R+Pd
xgNvITsPJifw+h/+14ynHwhH9f/Ww0rImSBnFuO06yLBzTBhlw0NKdCietGtJhO5
qhFhblNDZyfGZyo11DEXdyN5SFNTLmmdhAW2sxhwlpnlz4jLua0wYnExlqZamt6E
QW4cGPPBC6b93nIXiDY1e3WwpLBHDQdy0pDs+mXDsybat8hLawxhGSuJ+E/OoAK7
s/YoC+m9/jOOXFF4j7Er3N8cwc06aRJGURg1uKlLzKmPepJ9E0LG34CqBHT4h5ys
VB2TkFcRlfabb9hrbQEgexum1iDRjDRe8Co/kp2xlS2J5yw4qZonW4duNrlEA61J
5uWZcojcCGjgI6gOxwGTEpYhtiwM9+cVWgS0bxwMYvP8JBMGqPIPuAmMGCMXpyU2
qgoABGL62KLJIDOamxTjhASVDaSNTBfaBadbUt2oRdG+P1ZmfYjawjUy/DZkkCjX
1fISlFyXfK5SQ1TG1CyBTWZQCg83Qe0w4Wc/TPIXoq+jhvDQHM4cZbSAokmmOl5/
yTKXMjlwSvszmoh0vWnLg90l78ZLpXH9LxY4vrj98FNsFy744Dv1oOD5FkrKCzCp
EDJQeI4Kof85dQt7ja4sRzOpsr5aewItFghgtnBJgTEYXvAwRxIZB3c0Eq2BzKY4
DrI/pb6Rqh02xd54JFD/kzuL1tlodShvG3GjU4FX48RQ4ui1dOMtcuI3bUD14sPn
9YFKL0rAFZU6xqbADMnJ2r7JHSQQbChzb+ryKU9ETOHjtMD6IY2BszDu1dKAsToU
YOSR5mq4cyKDNYylbHb/nsH/+cadbSoeTlhcievZ3OyjaBkHQCZ/2dJ9UxzivFeU
jKZ+NRQjx+9lCJnSy/5u9chOGMnFNVLv2gHl4miiRh8v1baQ74gADqjkQbVHtqDY
JcDEwoE7StHvvzEb3oEEhHTXulqtoEV1sgmqPYM6yC8lXObgwz++Z02Tq2IbrQCw
B2uAaNWsZ5rkyJaiKBmOn3jenKSmtB3AvHP0dtwFnhNM4yycPsDQ/wnsjJPGVJ7Z
a95SQhMA9c11I7qMs3h8UziX4xKUPh1lNcz4SQ2dYivF7PnkXx8ulEGT8kNe+Zl1
caRtAKQKOFXbqDrrQYgy16c0/rUJIQ4a7hOAXdECqAjWBXywiF7vysLlAwpPeQNx
b/bKQxNB0309K83ofblNAKVZP/R4lEt6oPoCYSGViGUpbwXeBSTVtlOIadW3ZoW6
iCeBAO/WKamQHZ4QREfauoVKzlDNbJPhf/lnGWdi+skXf+wA2KLyvoT5cKlA46Vu
v9TYwHXHp5wUtK98ZIFV3bkTB/XqZbgn7CE7eRFJDS4CC++b8733Ler7Yc4XM23E
csp1uYhtL3arYObaYpuMd7g6h64qzw45Fy3prYrEw0F9ptdfAAzcxOF6LkKumYOc
KnsWAiFm7hzxlZC55k1sfY9Lnnv/HsK5VR5tRyq0/7zySYqkw6epaasUkxeNekUn
McX/C/4SHb4xXHlLJDgjAL9TngJhpuP/s6BRYN8GYPiVOkc9Jx7Bs9D5T/L4Xw0x
A91/r0+eA4uIBNCpYVtnNfPctu9DRaZ2k7OUdCA4OCM55bTOuZ+NHHxI4vN61UzJ
a2gbxDzEdZvLbJwygBRAc4e+WivpslIy4KFlq4GAosNWEokB7NtA97xONtEx+124
nfvePyc0tzPPEJlNjfs/XQ==
`protect END_PROTECTED
