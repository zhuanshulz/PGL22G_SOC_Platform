`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G7neeJgaa9FSiijo3TVIxdDph676H4pW//1v9Xz6yijzHcaDe8Jxe/eD5i/QTwIE
YsEBcZFqttjQ+CJArkRZUY41LIXKJQjELupLagFUONa+8vE8f2GUMp9xY7UfN+Gd
mneVdvy1jjOucFManOcuqEEJ3DOStLZrC9TzhHhyULhXew3HofHLclknNqnAQKDu
2g7pTrZdiobCVgfIk3O3wBryNFHyPjaOKLBfWGuBfiJkwAHLz+8csjB86hAsPypP
CxFuvbprLs+r4vHDP5PhCnw4aff6INXOMqOjqFgaJMkti4dJHj2gxY7wuY4AIhWt
sL1bRTaTO1JuvPkmTKNl2hZYw0Xaoid6M+dhCWCUzt2ugyWbxQi4jUCIIXMBrrA1
H99uJq8hITX7XDZHZYZMZPgfBODK2o1EHa+fGyjQ7BoeZk8O+evr9Io4gJvRMXoY
5ddA7uS8DI9i3U6VVq8iwFkrL+/eghvS5T/1E7/bOBlkPksTkr0bmHff+gzyBwh/
TmBYTsJkRo8wwG9o/38xdav8Q8/uEAjNmJrMd/JfxZso/13z+OaCE+rW4qITgNiU
0KUcc3DrwZYPxl7HfsN5xVtVAtBzGQw14Fd32ByTdN3infEJ7jVFbyW8Oq8abZzT
kp8Ci/T4vLXekjrLwRMOQeWVbLoHo8j2Mzst9UI78eZWuigc6XcWmxps+dW4/RSw
jd8iBpRuedun83/OzFhOu5krzZwbvyNo29Q4MABnLYtiCDokMke1AFblSmMgS00K
Iy6fDoQG0I6zEZr4I1DI2JWKUVpQOlA8cLhEjUdhHzMb3CAoUQSjPm/j+gslXk16
xfsd8dg+SKtukUBGFU2pgxmA2P/Op/2pbbKGXL3HrlDAfMCU3LIvmArs0Nryr0OY
1HLH56QJ4k6zSYO4UpHMhg==
`protect END_PROTECTED
