`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzN49QS0ObxARjuUyAYhBPJktvp1HwRd0NSTKHGW+RiQCz6IQrtC/iAkXtCmFSop
DkQs78w//j3PWCAo4o/S7I+of9K07AOFmSue1ezsETekUQwEOiuqy/QuAQQefCkn
fT2UO37bJ/IBPzErGRm2ZJXOedUhghU9AmpvqmHN2ZmG1zO5MquuvAx+2GzywE83
BOFpYjFVqEubGZ0+NDnli7tJeB8ElhuDLfpzpK26UGL+Z83YOPpzt/OxmdcAi3Ti
TbY3UgXCh8wpRwwB6iKr0Bvq19m4QdJ1s/i4tTdDd29iNq+ylFeOUG/I6VTJKUm7
RrdsEkIYbcxH1SIEOqbTzO6JrRuTyW7GAF9ShNU1BOTo61ECMwDkXeg3JD/KcakD
i7DR4aK1Nj4df7WfCqpFCTvwdebRRE5RZpHOIKDNnS5g77EmAXyt+EekCXvLjxAx
x2L6uXqmBUkRT0R0lyth8+UaAEue6Q9p4tjd3oGFQm8aHKFDcLSYIUk4SH1zS2a3
Gg84srEL6LN3WLkyx438wvyyJBIKUWmH7rv33ypmAFpvSlmMYFP1/oHCcmhVkI9a
nmAudhhrgBz5C1JgQ1rg1aAUHda30IDy9h+tFKsg4r9Fml9RkcQigAPLyHOzh/f8
nYA2AqK1FmfZVs9Ca8F+MglDXzowzqWWXfh+Jfvg5dayFBtHl/muRCNQK1RlIGdN
BnLZXQ9Q91SnUhkRgeYBcXnvFMGIqTgj/auk9QmJVZvT1OBaCKhbnQLWfbm/aprz
zh8UOYDTuogJ6XK9QroCGvxfyfk7gy/HW5Q5UhGC9XsugqEz9REizP3UyjmiyLga
IIVYX0QLlNmid74+rVGVy1xZcmGANS2XtbWVkyTFgUGD1ilk7imSoWfaaHCRuWbb
UrQ6Hc1mRWAe6CpTuFOF7AAKKXG86BXApZQhWgGJK8NUVLfP8cEhj/aZfHYe9uIw
OL7hOMG5Zq3+0kUcGoZDBJ0J/DMDFK/DqQPGRB/5tYPNZxLE+viG/AR81BnCcP/R
UgrvBMM6SIsLBVN+z7D5HiJOf/iBsRSKWESBYnZPSOuQn46ywP7NwNSy3qO0O5Z2
kohd++/cSHcXYfANS4xIqzz35VRXkAS7eAtw6SsCTfrc2AvKnpnd2/Kvh+fwi227
nKgsY6qca5T4vKmKZa7KXu1iyS16T5vnjit/PIKtekpieXIIGy2GysFgbIOKWf/H
a3WKlSKwt2+/hU37qHia6/ypcRnB+2ALpGkpVVDDm0joBfUiO+mE07Ok1pR2IGP6
w/Pfs+WZFvFhdsVnQqKF/OqTjOqSXOFDyTrlnQryLW4WQPlKQgDGtilUolrgi77n
X1+yarzYyuVVJcYRwohCbmvgR+SWQT8cgyOLKq/xO8C0f9ygbikcFT8WCUtWUx/r
m8KK9kPR9w+JGsAmoQfExojmWwDL2ZZDVI2G+euZgtALJFFr0WbO4rcPTiauUplx
P1DtIPoh5PFaQgRybn8jRucuhU9Euh58OpYfAe0LdA5LMhMVhOPysLRjV3vDpKX2
YpMo5YRHcXdn/YG1ftsKY4KSe57qYpqr2Q9aY9WTrbuNH7QlxE6N9hBoFYfVRTja
0P8hLkmANlJzxQ+0K+c8pm6T8KGTo3NEjSC7AlONndEkXDUsMpx6/yTPjuIq+jv+
kkA9RF4QyMCqa2Qb0WaKF9J5ZI6rGWw1EhqbQcE/g6Twrui2rfQcyFMJ2T26laxX
06vZpcMKALI6jVM00zFvhTOWxmLzKHFgWXIIDLi4+KDPy9q2Bg0uPQmtyytzk/yo
RDwjtZlKkU2INa0/5h4EFbmkyPeWr8VwQY805PUyEA6d1Bru+3LoPVsksJRIpXko
F91T+YnVC8AJa9dHnbUtD38ccXus7I7iGxonzzZF3FMCScUyZFIXjndKQpaB5H+B
mjf9qkc4nkn2/U1jqkxg3+6f9rN+EqaPgACOou+k3+74v46Wp7C1JfUKKt1vAERq
ylJwl5SefsW4QTFhLsGEOAezk1xSLBYd6wcRUxtK5dlD6UV+Tpl0/EbRnHuljZyz
+q71RSV2PFO9lFB5P1/gY5loYedcZFcsG7+eMlsvMm6YhUzDhppgb/ZI+u0nSm7R
f+StgUacPqW0Tur3ImQmW4KLEdWJUrtOXH4X8hhX1WFTgEcLcn3f84BLwGF1AU0O
d+XOYpUTqLoy3VlSleuyNAatQ9yn91/Eze+8wl9Rn6UgL/So/RIKTIfYutwA8Z7e
+9kyPl29Ug2mpZm087nYtX9nqGHfopw3zQM9r/HerBIcSJ/qTMJJG0IxmCX4mbzq
PojE0Zp6Dtm0VcMgHDYbq2jh4AdTSZbehkOLSgczFnO9N0WdKh54wPbO0L1j4K+o
o6a75nM7uIEnQqpDyC/tWyl5jt7GLh/VJd13NBq2Ngg+f3o6kmYc3ZeY4oCTyKgU
x5WPoi259BpnQHYBfhhFt3fKO2F33sKEj829rvXPPnfea7jaCtWxOHWQimR7nkrI
CwKBFiVUn+Dkmr7JKKV+sD0uu7mEKrwdD8HpfNgfR6EYCjGzf5GwNYnoG1UJj1+b
Q0Q6I9Bs7g1WsuI74EKJDeaQWb0xJPgSMzHWwnP0r08hIodJoqaqc3PK0AMR7Zni
S+8jqbrxaCqkqz+MSJIMkNPM1a84z7ua8zLdsxK8Vd7ATeQHaBbX2tjj1eO8FCUZ
/PLrlLFjpjgcxWQ+c+TR843h5DwwftMtkjGzDOVguekfxmKqVmX7GhJE0QVHhQXQ
CWAFPYysqCtJ1dgIVM49uKeAJclN+TD7ZppOprevRCc+aAmX6jWAeOZmc9cOsF4s
Cr9XnOB94u+Vx5mGvyrg+4Di678IWCYjQAsJ5jpcxORg1nH5eHE7oQrwJZqAXC8b
8zw6Ul19BQNwwE7gUlFshdk1nWRXAmzt91PCrD5+mcIgsfL+xR+HEZnfsHO+57Nl
kdaCopb/9XwaDgsmwLKIj/VL/27+48uozXQ7i1xh/bIdN8y/dW2j8LMfRKOxZtLG
EFOz4v7rr6lSHGweyacWIaygKp1dRCLiPqwffMVmUiUET4P5O7XIr+reRsDd68Sn
bBLKfo/wxflHcUPGmZ9/HTs9SOg5Mj06WVZ/eMv4GKGXPQbVHPccabCaO106R1/r
WPEH8YksMfazxN4zgpWNyonV/MRhUicnxLCmsi46N7coxbYHRft1dtceVhtXtDx6
TLDhZqi/qQSR4A/8TA4FpiXoDGkTMbOx/lSDmIcDYXTkr1x0BhNgTL9Lpuay+Mo+
AaVtaFBKwsSiHTdMpv3Nq6/Xn973OPqB7bImqj/dHzt4MCysKsaPXfckMjVA1xRu
+JHUo6ZCG12SpnNT6QwhmkVGXhHgU+krKR/N2+Xgl1+In3Kj+9AEW2rIJHpEKiqy
Q2tQJ5ptlulL+v+rc52TKNZO6INbXDFC95Ci1Ne16YckK6J/YybYtJ8mI5Lc9eM/
NHBoq/ITN/St2RylckQlIqc/0A/NgD+bGAHxvEYpeyTjia6qg6+pk/40GCD+7ZLV
vtvf6Fmr6WiEVdt8EYEdRBNr0gIxnyOQq2KX6041NOyZ3jMCWKyN5PRQyyt8sGkf
6hIZ9NsMdRcbsJ9nQOBfdTWEdvOy45EIb1WUFI1BmzuUAap+dEssKVug1LbQ4eRL
8Jygu5D798HHR0u6NMdPSSqpxmKenpnglTjnuyXvnCGtMCLJNnsuszI59Keq+o1Q
98uwgzwFCMGCojs39fJpunOUs8Sf1kpGfH1j52bu/yCA5OK7tfMjrCnbm6jGXAGo
7M5aSI8Grn8SSSs0CXv6+9bk55yxPlssEbZFdMKMXVJKL7yh5MZkZl0HPe/zU3xc
PUw2MI8pUMYAKi99u+IP3PdBKcENlMbxme+s4kVZMBOHEMsr6RaWDr+G/UVpx71q
VhtCLMlXexZ6Y+UhKrNHtsKF+lnuAhjhcvy1g68nJ2G4qmL/58tbSB0zngrFCAeU
ZTHjpVDa5VbjIFMsInuHlYSmAkR+2v1cMa+seIgPTOfRD1bQAf9BDXUqE1J+oBXV
0HlCnk8y9PJednq/un5soViYpd8hpiA1LzhJcslH+aB+tIBP8J61jUNgVTDfA78O
oLruXsMNx9xGH1OPfkdtigVbXAQ9HqUfMwfzq95rNhPdehf6zeOMZzd7qjagX8JH
qOj0Eiq/TAtKDl7yeMAiVRPhQc7ty54rpzAfpjr6ZSAUEDbDFfKfYXccAkJArs3w
i8HYVUslAtMHLxRdoTL8xnjZrPt82FbP4vMlIx4NG4QqP3APe3fI0VC1gDU80/Uf
tNB6XiydummFZuQu5aYBHW/iiRGzps9GsBnLFUvJwwB5CGfn8WEgzkyTPFAbn3eE
HJG6hWY/r7/WpQRdjXtzqvUOpErOj8XyNDyeyUKD0/osSNfyJa9gPgk3+oiXa2BX
qrDbLOl3SxPCABBOMChv8vlWdUtZ79z47ZHJBakM2+hpN0uXF9PK8/Y8UwWzTZWy
aK3F9Gt5/1REFUO9jrzix75kphkDz4myi45yGJ8FotisjkcyAmmqoOGn1l7C6Wg+
jKMfbTGHz12kY+RCxEjF4dPXrCd1C/PqekdZ9IRANXGx5W4jI6LTp8m93XDS8n67
gbGymHQu4leQp/8XPjEIw8lFvxpOFyA8dykHpgHh8xoLgTawGDC9VxgBO9or46ea
PysPzxQwgHyErTb1096D7X8HtyUEBj8oMPxNQ52KjqFcWy/fCIUGdCzpwUC7ow7U
/eOO8pjXmSdww6Q+QSNEwee5uOge6tZYbAIUVFdc3RXZrLkgKWqCuGhuedBARcR5
iggOGpBgJ++4kQdFL467b5mZwKdjx9POlnijy4sVvM6/0ZQX5gvEsdo1R/2hVHf9
uTjfnQ9jzUyusbz6+fg21JapfX6bUST8lq/iaCw9RB5xJND7TM5r35pOjSdBkS7J
bK+a5bOYb3dQUi+dToQ8bWw3JQ2pHdesSmadgriTYdQ2efboMgM7FYqfGNZp3v8e
jVIim0AKO9h+jqrgt6T8Omw0z0fQbZAF0Wtr8xujtwZ5lJ2mBbsKNZqRNRUNdpqF
ymrJ7czzgj/g0RnFvucsOeogQbW4bFSOea7veZ6fI+/uNx6qUW+xUGQuMWRTe95w
yNZ1rUvuVcklwXEX2U0pCDUlPw/ZvjOwJsBT8PJsGrPWPKXelXVggYCBPC7NUaeJ
vrOuWkFeVW3DkQ9x2yiCAJNqtQQ8M+V3THIpSIGkO4XnSFd8F801EVCvEY9UtVFx
o+cEJskEKAzCCS+bzrCOROXR0fsR8Uk4rwyl88v5r/QH6UcExZ8iK1IuyMllwam7
yjQyqUneB9/oArC8Rua91667e2cSL/rOvb30cKVuOfVB8gf0rgWzIImezQubZCwF
JtSIFov3d/GF7B8VTIzwB9Sy8KYNmTZtjr3lBcCM59sCYHqJJqRT62FHNlBC5pA2
7U9/gh9kyUnpB/w2u6sdY5sCGROBZs7JsjwcipJQx3QDtk+EtrKcsPAmmi7hRjxc
bHqTZlJTpdJGuaiaHm+k2PM/0MUOAQBnzX4KpzG65Q55d1oX0DzGsyhSpAkuc4IN
D+iHxnXOQomwmNWGR8j2BimeFW5D221MEIy5g/geAeqpZBqOSsl9gxAZA1z/THDQ
Ib+NlUL4yynR+BlUHOZjMdShSLeVbDYtH/YIyONafmJ/vR15pEuEjUWxdf/rtW2h
9nyzI0jVqFxEYsE3lJRoaQJgG+2jpnnE5SmTH2n7ikTKbHpDxmCnoEoiwHioCZnx
4zC+q6QzKSVxqaXz2dWW7L+XIhKPfStUs3NvUQKXfzjV6DJiS2FXxlRS6Lna1kE/
FLLkepp6lZli9QEUWSn/zrrtgIlegcyUGIhkGsUAroutxmxHSMLqMrSD6870EKZO
ryyySnJKX6rzTlgy+CHvDN0JpgoiDOWNqVAhmV+GuHzmFifJMES8WjdaWQMNUFea
iXZXbTYkoVyFQKLQyqbR4wpN9Zhny3mL9+Le9RN62RIoT5C3kASHU8AxlsNO3WrQ
zWPuOs/N77N1wdx5id6oOAOoLn5R/chMjf1qa4Ty4roYRWFciNimOrfCFyJrx9d3
Lw4PBPjL9fDM6dPV/+sKzkMAf++ZfgFYysa0WDXNSuvrRkC7uayG4021fbsd1vLq
B6LsCpIr01iywkuTbqsF5+h+nISRdETB0HGRT+xkHukfVHkpZ2HB05hXO4PM2tOH
gPUeuJo2ftUcfWWh8UWVAodU6fdfVqkASR9G1VazU/MQnGmX8MqtAD7be8ACTfW2
YfiebYZN0CQs3VtWHY196YfilQK9n7wxabARyi69QatVPqMC+aYulUN5Mq0uKoLz
3FcZyOWx/lGqJ9mXldihZZxVfe6gEmdaOLNnU6kZ3KxXw+GWOSR3HK5Fj992l3Ax
N8vzLoUoEq6pTC7lgGMCVs8nPOZC5WqUN8rf7Tizqraqtj+mkIfSGhZj0wVVbR35
AokXYgUhmGtIPmSiKJMlk0N+9oJlUoDwM+gyRabKYTwYe7mVkrI/8Sd47ta91llp
iA1ug05jTH+p6HI5QdWwpxxS5iGftD2JB0Gj1MF7empppT1ycqzkU+LDVUs0zc9Z
THFlWqWsppwDQCVvTb6Q27nVGg3BSGNFGWhCZYXF3WNHaJZYGkDbs7m5e1DfdPlM
Bb8Wxj+jG+R3JvmiOYycAxbut805HMCPCWgIDEK0kxkKWr9qIOzJIlGw4JC+AbDu
g1S4iNAX55IE2PSWjT26fiz5py8MHsoYgY3VukkWpjRVH0Dl3vo+th7MROISd+ix
PLCl/scOpkn+KPufCRmBNNdJgEO+luH9XwKLNp/i+eLXr9azlM4c2QEUkSImH0Au
iYAhtT4WfIBOjzFqsB1y2MBeQmi+8bfPKKMV8TIfwdELFxzZ3iBwhnZdzuI09uyM
l8ZURhBmZU4w5bO1Q/Y7O8yECqy9hlYKfCzL0RwbMSbFOJKB299/Lt+sYvsh9rOn
tRxNidvxRHH0yZQrgdFrK0lqb89qcd2DaqRtHegHI0Vw9GGRzRPb38vMndDQvdz5
4ssyu9CeFfYH13gLl56zmavPondzsJ3EAaHw0KJmNy4QWyC95dyJtChUlw7AFiUM
x+dZdeal12Ar3D9DPsJI6LkMVQWjxy++H2JkFV8hVFue2+qrEw+UedOtvHi/7miv
nCckogmr0xZL1Su/h4kqDfZxcpT51eYcOiYBrWjdsdRkbAyCSuMC3lcIx7w1mP2e
cyWTa+CCCBv699EwBNhZ5QhyGw+qS/c7VLPRLtSnNDQRyRIEjFv/wBREiegDcfJ6
Fiw7YlW/alth5c71IBlAz/gLjGHYLRU4TmvVNV0VtmXOrPaJHr4poqKUUYop0qIe
F3SS04ru/+TUmRltUQyV6lOxxgQNK1CD6Dy4YsQ0LqZdb4HMlfY4yH6h5VnVg2ow
8sMTPQMAYfyfCD+e04iy6GNzfNsqwwk2gy8R5W7lbxZgLarP4NUq46EfNn1wSYbM
XWChrvP3B6ABIRNDZZsEwfiZjqB5527AknIXozR8OdQUogJFh96mrguTQk889Auj
0nX9PEYw9SVffPaFkBuHIxgJ0CHvc59CtnfqnNBJap+cPOPFUOxQXJQC5fXb26cD
k/3Jjz2kGOGabadnkBzQCSaSM0OP+bRCJyyjW49TNGDquiv3OFWqs2fxx5N2htNZ
W62kKDQ2OEWnMx6LWeApDAd6xhQdjADPItaZBmdtCYZhdGD2ManThTMQYOYjLQ2w
1zh7jJ2+DxKTMKhiK4vVZXNEI1o+2hL4b97n7IwaqnBZsht9wQGp4V5T1ieP0eoh
YYahIySLunotGZeNBE5gLfQPrP5hs2dOT1qXIqNddp3eAU7tbO4LgSdUW2P+RZP6
3wdWvHsuLhTn6pGWNHc5vW1YTEwdYGPjbrIBts44Wvucb7iEXYt5qoIlT+FpakdO
ovP5T5jA8y27zpji75LlXGYuzV47t5CdOT+tAVF3cBBNdOAIhWHt5MugR68PIVnb
xi2spw/avDPOtVU0t4wJfv5kcv3OAYYWdK0BP3TVS12PtrNLVMdgMsq27KT/Kp5X
3empKLU2GoX8KN/o29MXjqRaxa0th1FiAObukqWQb1sXnue6tUmr/cpGIe19yPim
TmkBThKgkgRKRWWtjz5e4lP9MzxSWZy+ZFICfr/V49Hm4F+lDYZ1N9jqGyz8PX26
+Y2AsGJ519Hjmky//GzH4gUVyic3q+kKYhwV6YFewKiG5ogfUy66iZoskdyzn+ds
g/kHq4ZZk2i2jny/9I5ZlA==
`protect END_PROTECTED
