`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KigKHdS5S7YXXUqR114SoocHnEnHhE0YGfU/uFz4xWMVHo/x9YudbjCqrhAXQCq9
88iFip6RgfttII0oQ/Mb1KCMzCb74mFmdedAKwWI4D72zUNg5WVpZbWrK1KnaQv2
WaC317koycQMZvvU928kXlv7QY1bhTlC7mOcbZzT200NK6F1MFhwpCRnKYgsnoUn
HlOV4h1oDVfvkX1u7yiqOqqFMl7VmPV1gdQQ349t/cgmmfyD0fLKLk2ufBFrH/Cs
apypsn3CgTf59wbspNwWfP118GhpjMTy/aCQufLITEoB+a3oMySyGPaE8ZjtMNXq
vsgdXWai89jg5xNUPBTjNk5mqZ6HfT9LHGa5OPRxytU8JZjKXFFMEskU7dH0Zdol
plIXjQbDc29vvJn+MyPBMsTQ2JWh0QU0Vngu+4iT/aZsuUPP3uhsocpHALZxNp9i
h4hiyxNRiH46OdtvpkCQYjKGKh014gLS3tSGbExk+nojj3FdB/+Vv4mBTBEAATli
R36dsC87FtfflhvlN+kIgeBrK3WzGL5c35KvlDC1QUR3Bb9RCylTEcKfwbuBmUni
Kf5rGYKrzQjGHjmkn0a5eA==
`protect END_PROTECTED
