`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkIUJtobKzvZIiewvL5sfYesJ0iKuBSdI7oOX0ZxZZNiUgRDLMhCmTTgQ85yD7mL
bXTE6v19t+S6B/QFq/dww8Yg6HhqSbAoVem++YFVSM+Qe2pjdu8/16oyoOpqyu0P
wvtmih8Cmt2PUuK6mPVPksTrNkv6tVMdJb06bdbyD8sli6Q/Yf30eu6wXlWK6T3p
e2GPG+AIpPP2WFbeswfPTPw6Xp3NN4u7DbdkQUM01cS93TsDYqZylQpoccSpWY2x
9yUFtTDKMVztOLdQL8fFmPyofr/C5vrsZox5theFzXrnRdugNZ16LLz4uI2f/MZO
McMHSlPfV95yf5JifqEV9CSxU6hbQZD45UeuoYQuyIz73/gzWDtCmr6yC91gjXxq
LwzwfQeummPx/fwmN/c3rDIN8Hga87d4wgOUoXP8BRjJ4sQWr6Tlr2jhQ2N5pa0C
dY2AWICCi2urwYElDldQ/rnlCqyVjGiN5Y0PF58UtMtzjNT+U7WACXMms0TGq/LJ
8gkxxcNGh4fz0wB8oXIoJSycLvXe3RivHB5DkHAUXOi2ofLEyavrw9mBQulvejb2
eMRyunCca1+RH/caRckAhA1CqTDcuIhVXrIsDsp5IC8qVB6/df/I3ucYa32sIt/z
aliZItl6JCsOS7Nvs2FWASqymsVZp1qFReoodE8YUxPqcLJvIapyZ2GCIZpvvZZQ
BUMXfmP8edvU4d/JEY/OKbEkvoPTL9bypFLanaCbS2NylbNP8oLMFY97d1kpUdbB
2J5w8btsZLOvkkeMfldYog6rh/VGc7Senuxz8ow2qIObPyzsHf8U2sBox7uAyM6X
bJdr3pwe9Xb182riNpRjTcBuH7cv/bwllcBkKLwkvMyz3JeNqxnMEnlyRK2SZux5
Kzu5zDuwhH9Om/mJKSlfaMzKRlx8qopvO1bipLdl2KFHWaLkge7TX8ygN3uEmjKV
ZepvfccrTRE2UOcYKms3ROrg/aNeB2HXvVQMmsqDwCSwOz767FmJhwbICQyOs13F
qXVqi9v4nA0Hv9BL800+KXleQ6cDyx+ijseM7HQtCWIjJMOqGueu5roT0QPaJ6R0
2D7ELaBODZoFVhTzpAAbAj9CukfsMQd9SN9idWtcTl7G3/LiSkkjA7YAPg7NL9XK
mLaTQ0xF/HvCiocYsgnoSU2FxRtNASkIN6Z2T6sESM1Wb70GBllgkid1Ewi1gOre
30XF4OXpYMMNFBDB5xhZjPp+/G9yv+2HY1reFARW/KI1dcCvV7My6jRVmKUZ4tEo
LDskC6tUlOOCCmBdWv6N4yGs/4xPta6usPoJTcCfPRn1GSjWXy2RHlRzlgFe7v9M
h0Ywpq6oha5ANz86AOPJgb449UxLBKinNqwy9HDS5yz87fLTfQexazm1lrz8Lac2
CNYuPv52rZfSocfqb9C531Vv7uGr9LJ12gTPFsm2CnHWyy76gM8dNH8NkmnkkmxC
338WIAf2ECeR/PknAWJA6pQZYmMia2RPbyNwwxLj929Yf8HyW5uhIPFHgK1MPrUZ
ZNxDYGnpwWCAkLJdaoWwXtA6O1sZHe/93mEFue5Rb/MtJPAQB0ODpoLA62Zte1cc
5zN7MHVvx7JzSILi68xIpQ==
`protect END_PROTECTED
