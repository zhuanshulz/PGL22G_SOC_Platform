`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ERVe7qAW8FxR92OWQ3GcwJKzBVskCMmvzWktfV18F3WukHBJD7gZB6X9l/rZauAt
f/6RrUd9FskPJ3X/I2D0dx3d4fooh7QkhkApFfdq/hZxTKvQ9hSojxh6ReG9KvHE
8FOH6os6Rt+rrdgvXtpPafNP3tC/VUUGCkGm6jAOH/+WWeF40agjXtXDxL2F0LyE
nQPBklAN8cq/oo5Vz+7oxasa5i3SeNK0quQXiLsqZfOMdo70r4Ei4Qj8MDxkauKC
HqcmOKK6LTiFv51HDKlfs1wZyC9o//HoNTPFsS8rVQu7i1hayhQbKdL2RSQACcbL
8DrVys71FFmf4zCVNOCrseo0gjAOVP2az3/Y+s4aBsPki/1FUTdwqqj4YMIaaotv
9TTZTXeGsIY87BXfjwoRfp+LDDlJXrQFUow4lIV1/BHcaVI7VpCfqLY3F+VhKYot
Rea3if4vt53dRsUCMmMqLGWa16R8PNrMfi0dcqDovXOEe+J/fO3D+ohHlpt3qyd9
bQwcgY7fWh5svQTDCIDl4aiQ0lmTB0h+V2N0pia7UorP1HQgFI/24NK5jJ4ylz9Q
JfrdIpTiYR75uwjAYWrCx2uyIYhnQuooNAIUluFaKZUkQpAFGI+4t05Ar3GSFWgP
kYjHQPZV1QumeayCF+fZKHdbLBThbXtsmHwQn8gj2OiAu2/Cnjc3PIhMply+ehid
6uOq+v5DptWQ+UxO1KP5sAowxB2zZvAOtNv6lD3RHTQ5BmbVuLAsuD7JaHnLvxtl
G86iuqLoZqqhS9ddwFIsCYz9oojbm/pwcC9iVDwl1l8F8zxVdBnSZZZ3vmIXR8YI
2jZbymC3XDk7bxtUkc1pwg7FA5FOTVwGhR+n3W03KzPno5qZw1xApD8bY2Sd0qya
ussaE12KCfoEEfA/g61x4DkCfHNhwVH5uchN8M/lSe6ZPoxPTUz7H8T+bx6s7vMQ
QDoLVLePSyiDhvl+//nfT1v0bGh69Vykzy/RK1EpWIuQCrHDEP51cdk3LHnNeIND
sdlCgbLqBt+P2sg/tnqModMrct3EwMy4refQ+RB3z/K5M1FR3P3RA1G2EW+gqDer
K2g2M1JKR5y/RFPxGC+UqMPBXRzFsPdhB45sH8fRGRLwmWTNWYZ0WTzWOqLWLe5k
QIL8LMkrFtjOL+7OvgnGBYRWkbXGlQ+ifdHI9g+UhrKHYBkyGr30jqlhm4WL5IYN
hKA1SbEm6z2R832O2IfsYHzHD2RAjRP+d1xWGjbsW75YuJRY8lF3/CRnwg0K20Pb
m6xS/MwrHGlX/gYuVANrLTgmbLluUXeR/7ZuEi/1wBeFEAm18kMiak1HXzFREeuz
RsFsHB7O9iResbefFq8uCnJ30oN6Ir4bVseXcrmBVg4YJMVN/EftWAg9DxWbArjT
9GN+2umElrAkTD+wi1Vkcurw/bNYceZcMDMgbfRrFFyaNlR5oMvdKgMH/bFFWxSY
IZZ5thKuVq7AzXGXtTq705ndbFOgSEOm2g5Zx8ijuYZcjazUJQvQpZ23Yus0+sZ5
x2wPHCOMEY6vuZeYD+X74CvX/HO8OpZghTD15DcTpBpclPFhXTfNAVNbNDpwqm57
4AvjoAXjnvFEZm8zzIttlX03FkSk6Z7K9wpoEvh5jYQZo4SJ0VrhxDHoO4newgU+
cbfTaEhYOcz/T0+XBGprhXFrKEpbGL0/d8I2+Tx/5liD+USMRHhu8NLbmOe7XJk+
5gWyzN5z7h2fTJ+3PFiToH97dDk6rTk8fG7V3Y5cibX0P9Gl2Gh6rnLNd30Gr6RX
AA8GxkqbyCZ4PEmisIDFBaDXjO6D+LiwWc7HY0kW9kqrI2CQhKNbG58WqXwGpMb4
`protect END_PROTECTED
