`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3CY8lEbi58745iQsmDDRtLwjcv6pt1ypuo4d8q+4UGTNC8nFOKKVFfdW5p+Tfk2L
DqUGO47Ck5YbqqsYvsqv4jkZjoWGOFI5F2G87hnw9Zr5UWN8XEFP+MY56ina5vHT
UkmZyAmW8uSR2lKDVUwfgbgvksEqJlsupGxBlzjRYY+aMyw944HfsuVpX3NQGOWb
Ybnh7jALpmW8JbWt+k6GWhwk9VQ2JIvzd66+iiWNdQjjRzFnOZ5QxyulmR7ASTKG
pAF+sGm6AXdKCoPsTbomzy1yFEh1LNG3af/lDg0OEO+nNAr720So8B72C8hnJqCo
I9PMlUEpJBhmiUvDeyzi8daujk7gEzu3FBXcHt5UhIr5fOi7OW8/Bg0BBHCx7bUM
9H5hnfNMkjfQQBOSnvM+DVOL8gsI396fgrV7G5wPJO40UFzwm6lTnxn/45EiaDYK
RnVtKNZ8A3s6WblS8siQZkiPFgMD9+AX0mINHXPU2HV5OI7oKNzeJRySI56lp5ra
3GctbHBXyfFf/or9CuUcU/m0AVfrCUvmt/goTs1qnr7rdIjBxKeaD+dH4RAxp+iw
N7tvh/54YPjVNq6kpqXvtiwSS9m3vnfLlgjLgYYY/XhhOTHeTC62mHGUyNIe6DlO
W4/BdpPiQrl1CglkCghpVA2zmH7ixWcW/MKUENe4HMlYU2arD8YUBzS/uKyfQxSt
K8FQ4+/DAgy85+5IOkvDCVNNL25Yl7BFqe5M6ssQssBolt2wMYz52Ovhbr7feQ1z
2L+rprY/fwEwla1fnn6auPIBnNb11maNbvJUWMnW/RFcrt8YZNeno2rM3syw1SSD
8tvtcI/GpJGvMdjjGjkb/od6seyaZ3gAg0bZewtzhF4go2YbPKazQk1Xk23pCkJ0
64pXjoH6liA7LZIy9XnQEAhDEa3XUM6zXFUTjYwz14SJY9bzL2wXgPobWfEWmwfR
eDlXwdLYQ30YX1/tCOVIFLtIG9OaVgSc9U2mwgMmHCNwF2u4/sQT6gHDNUdaN8JQ
pv/DBHd2UIwKv53M+nAp+gZiyHsZ6PLniusynBefgSzzyEEuc/xt3vW16znecMh5
AEseguHyzVsgMZ62+xjPtsJ5CnqZv9qTYYHkvUOEMuyIuUduq9jYWQ846/EH+cA+
9oNW3/Oo+2AQUF9zg3Ks2SkN6hhbL+OmOVIrqbmaqZp6gGgoMvglpHlRPOR58MZS
7Bf4z4VSukZPxd1jZiwGD3uue9vKQaWKUAfmffPZ9i5xU++R1K8S9r+7Gyy8cH3h
FVWtlHp8R0EG452xfAT7o5ZcoKxgjGV3BMz+kCxCM03pwBvKYPCYYKHl2FU+nw00
LjMdiYARPtG7qgEKEXWQXOE5S5S9tjDkHfr+W8buiH3MxFUdvjWvT02oJWUgnB4P
5agGPoNfhSBKeHP2B5DZABICQGQ+9y65rprs+VRZSDf7awovOvFXAuSk7rI3d7tM
u7d7d5eU7ujV6CUVPyK+FYsc/shd5sbFOEYdGEzXz5CvDz4xcgUKhodiqfLBRnWl
4EOF7hxa45eu58Krlbuk/AYsZp+eOaJyNramlj6xEdAov36G8CJAmOBPHUoaUdxc
ZV1wx5DBWeUfM+LU2fVZDc41T3TbMnGz4j08XgeZrREdhWTi1pzP7n8YktCaD3Y3
/2m330CD0SOkhUaCO4Q3IBriluJ5tiIk3mbaOR4LgpijyuwOHibxBW/+wbBD7kz9
41F1tBIceozeK7X8WZMg4MIPTt+YzDxGv1mAGAbGpTMkOuFWgHAat1fNk9JVG2Ts
PLTyfwU7VYyTjHbYBqFjpPYm7pYRVgjWmaX+B5pvRLqQPUvGi73fmYay/ZuHSXdn
4Sfd12MQh2sBGiY8wGoUvrM4spzIB8CbycSiSq6tXg4EQoqm4+aP5yStUljFuYFi
xnz+cOJ1WVqpPoN98+EJOFaT8dkm/wyjprc6b2yXc/Aw/iFK94liZ3Myq7e6QmVO
zUcqxMNnWrcQ1XIaoY8Tto12oHxQLjFp0/KcctirJIonpvwkvKZbI0Ed/d3aGt8Z
uvS5zrvsppPMSREyW2NtSjq+SS5UHOL79OguZvJ8UdPLKux6D4sSXrVrmdE8Dc9h
`protect END_PROTECTED
