`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUNJL6qtwAGXDiqkW7fskuJJPW9Diir0CsBsTaUFa1ajnDdvhxxR61+1mgweq9xK
Q54HBd1ICcmA4/cfNvY1cjbX1sO81H6DmGlYw5sfVeUPdIhQ4v8kfdjkRwrAk16E
VHg+IT93c3LbjCma+Dx0ZI4Ov3GSa3w2l6pLXIbNx0qgMWgrKDmqUHIVoD5Nl6Pd
nEsfs/RWSTdGC6tm699EOj0UVbidPenLYbkj7DroKveMBjdUIwgxSqW61CUElj1T
0lAcNd1DOOCrd8dAeHWnDMNV0779Z7QSvdWQAvR/X8KszuY7oH/ygGRc89sK3oJo
cCFoKhaP8juXqXWZnqJFyLUzavZkVP7pRSwYhuBL5Uih5rv3R0OFqtntvPWqnFmZ
KLVFWm+qeBbWkJa+hR66p5ACSu1J2PEYxgnzUewalokSrQ8jNyRwcpdKV7Fn3wfD
fhkBrs/9YdjtjR64KYg3bVuYWauUgUZ40nmqjOewWzxNxmSZcZX0SEUxE+xjexLv
CqIw1vMb0mZ0EA+BGr5I1vLqCpARMFLjZYB3T09KuRGOQdTSr94claxDXA/Qzs+L
A2Nbf7ICGyRAbfimmhnyDuclIJZac4kHvFXdeQ8ZJQdeHYG6fONIFoIHGOxqZFZa
tXg4ZbwFKZx8u0Tzy9Yj7+sGg6/1xUsmwh+iP+EkDtUy+H7C4c2lf343ZeeZqyAq
KwyfqcZujiiTRG9HVqQ55QkRK70xQT55JxjKpByVnH7Fu3+he2T8dcojbgo2rcrb
KCBpedKjzYU8D28VQ0tpN5EKNXIo9HUmeGI0DeKj6/TF5c6IBZPFUgZ2RyPp+PPc
3z009FlYMHV8MW2D8KQQscihvHcQ3QGMhNekDeNDbZwUPJJkJzPeXnV1ZoEd4tnk
hAi6dudhgYUeWzAzjLbYYJO85M5/MjGfL9dobMBC9e10ix2PCX8xUunt9wxU4CE9
IPFsRfxTTJdVCuH7RsfXnkcoVnWyb3rqDqkUO6p7g9P+RmOsF0c16O/RdL31Fsbk
nnQ0XiE7NgySq5ZKLceYAF6KlwsTRJATe5JJUPzDq7hNLV913vp9rrPr+p9zUIX1
ddu5CsgZkZM6o/VW9ZiOdkVZHpYnSIPrdbKVOWjqtAXuCiXimE/kmf50l+T6O1Ns
//DKEgzcK1zg8RxW1ezj6YlbzwzYFEgvVhCIfThnKBVys2iLkKG8ZSaAHZELvafb
Ld5UbxtQs+btuxtJyeG3ZrkW3wdfZfhu01MN5fKXtxijriChTPE59hx3kCCE4sjn
PcB2n/zb9qbD2sGBdXpBfMObC4r2bl67u8hepejiIaYtdxFLMIdW3Ox/Zx4Npfay
/W0fsnAbPDgn2foDMCzATVsutP2lUtlkdpwQxj8+bpNkbK5/ygjzQgiMIOi0Uirg
7JflpuNVndF9xr/didljgTf5ee56/V9X9/C8XRIGgKNSMWEDx+SvLzEi+hSvMCqF
UD3qVbE5WOm3VKe7zViE6Pq+TtyN7jf1x61j9SC46LjAtgS3t6b6Gdszf3MaQY4b
FDy1fxKKx89mW1WTPFI4d0X3SahyrkHIPoWVA2pMUZ0NSLpl3jTblJZpCJB07tTZ
PVuKgagq8YXpoIafB9sii+qxULWfpvwSLNBNc/oSE0FmQ/9SUoUzbqAhZJe+58rt
KLXvpxFQg38+bBfN6xRbdgKkabp2ukfIxDd+ha/S/ox52RFGGMHy0iJ9bI1rFMU/
W/Re1IQY23yETVKQSutmIvSZpfXuwKf2SQsidZp00Vfmdy5zue4tx4E0HkPHlc1s
F2ATryNN9tJdHH3js5n6Pj7Nd1tsvzkoP0OFt6TTRd73H8ulN2vYWr270ZvMVnz8
uM8oHV5xl1dILD8TnpRUqcqxMDIF0C70gfDDiBO8XLyaY7NJ131TGMY0yUG3Fvb5
CKpUn2L0KsPejYNXdtPjXTqCjm5mo6OzwO80YxlwX7c80QQlLN3ReMnIkLjMLpE/
tnnUHuPwQLU31ru4s43JiUhV0hwPqO9E/vOS3g7CLFeJYM6cV49vrBY7hFraJqFT
sq0XuQ//ZqQv/j54CAsAeSpmiKDq9szKm3l1M29UcHGevon9OyXYVzqsfQUOHXM4
RIEPim1zm98vre7EdCGw51EqLXUFfW5i6NQMthoFzoEsuOr0Nsyx+zOH9umgoZh1
4Ne5NzF28ILQjPESceOFIVxEPpbzim0nZOHv6ireTK4raiQva02ONl1UH50HDfB+
VjLnATwkKH5ZoEqxGHJPgH484DKY64Yrscj9aj0H2eKVAU+FJOB58eEffSpNxmru
HfsuKeGsbnV/30D/H1sM3icVgA/aLrW0QoaJRO294ibohkql9SV4JThW24H+YH6J
3bHMHU9MAADngiq04O/P9q9pspagp0+h3bEdX6vr8h8ELGFp6V+DVm9Y+EoY6Vxm
EEnVcBqHyXCvAFgS5GIssE5JNtHm3ZpJ7/UmvFdwsx1F04DpTWuTBg5Iy1Q4+AFW
aK8MekAJ2hTQS75J24mUQ+5ETt0wg5U9z9UlrwhhPUEBv57y625Bc0jgpcp1+dqi
Hsykmv5HZpenp5SfKzea+Nu+7MgHIu6I3bj1grpJynKAqA/uiGrsgGqjxloUo9P/
l7J6t6CSqPE7d7MVJp6Xk/Z4MSYPByRGF/51HLWeEBgcGtufl/M1R2xHSFJkVvcv
+UyK6kADmrzgg6oJzYPQUYcHPYy9meBXklJRLvHZb4vMQDBV7AFvWbG7n5HOClBh
m+E0sLr1g8B3O7SJPw8pVzvjIvOvor2kRpBgKu7DTxhU1pnek5VoG8eNccHWJIkQ
EWxb+MhaWd7SO/sZKvsGr90FOZBG0lsHe7pKwCMlKk43wj+A7Nv3RAAJx46NCgLd
OxHl33WyVsAV9D5v26dbIZd9crpk0P+JWE9sPKb1XAHtNhaOiIBEmvvcYMeTSH5D
rDlGxvoxmqsOmxgRR03fFBv72QYXH6w6z74vo3N5yVii6cRDi+5YP9/mz3kLXHNh
Ukc6PU76OB3WpUhXtroNXOylFBWDeUz+0JAfnrWlRmrY5izMUFDS8QUI4vArZ/Cz
VcMzfJmNGrJcbtAjRTPs61cEw1qR30S1C31wVwfYxmcfxvX2RSqTkFsCZ4AJ1pO1
Y+GvkBwFZi068V4LYzAl2VXa0CN/QVO6At0qTIOAhsZiCQMZ0OcarRa78MeDRjqU
HxIgL7FEZAnsWryvP8+VzNcABzfjp6v0S8z2QvTMS0DzIcAqtyv853Dg1a1/1JC1
3dd3FvlWFW1Xi555MErt+Ra+dcvhyn7lDC5rsJtYIln8uavDhiBjS6yEq9ZNdUT+
Qy2BO7CxIEYK0LgJr2xEZKi+4tBiz0gyl9Lu8i/FLSoY7QFPklkw2+0nlMm4FyBY
mFP1tgNKhxetBdI19UqeT9meOnNRevC5Yj8C/jirhK91pn3iMbouGlzZ2X1o0V84
B66QSYd7CoKjYxqx+wwb00R6/8Y0TVbPbbpiV7a8qTCQXZ8+V0S5+px2Kce9AC58
r6QwbAl16mQvudlvh2jbxq2ey2QvuAkKx5/inlHfQyKp+d6Yr8L0tSppE004wmDe
4jb7cuhXBqZQAMT45FKS6Dgp8eEznLtntT0fnWNP/szSLDejtxaJNzpf6fJxn0jj
wk7EzmtinofC/g7Z+IHOclPJCdIaEBBatXp4FjHuEmYwf7xmJ5zBrPMVksyfrBKK
yo8xVCv3ZaaFgNPlvgWCxzX7WK2xQvL8kr8C0fClpYmlSRNkbauxuBBMedI2ZPYV
DbfvqCfh4JSPsk2hvRyUZDBicI6Z1zu70gT1cN3ATYLKAYfrTfCJzUkZRFnYhJf7
r9U1DZdeT8asmVkbGvhvJTiP/1BygKYSWywDl6q0lVMu5/2UWaK45ffjMddOfQqE
lafk+gZpZe2r3HiKFUJYuA/YS7d2JWvKEc1uBs1hDZEKA2K/7v3ad00M84v4Xsp9
WX0Gt5H/oFozEkCun/NTCwAW07HgNp8H+FHBviDEgT4icfGcU+B2JlENlNUF2/tt
xD2SImQzwVaqu7lCKNR2w/IZDE/28kNBQkY7JUEo7Pi2P2hXTJkyXsjv/VsO9ybH
Ph/AQnT6g8xmQcnCh0EWF1J456Ifgkl7grvVQQdu5sBR9TJXvtteRwnt0w5MDInO
XoSMVxDv4KnI3tSYkNbW7my0E8lC01DKUHtAr94O5NMkr+oe/leZClX2PnP0j0xp
6DhTJ1lshCmPbP9ErgZL2QvqxEIYOPh6ttblMB/mI+RrdtXcNALidN7jj48EmO/J
uPMB6XS99KWmsAnfDprSrlrRcFt2XHlzrKHICfh4FxcoIg4BQ4ZZWGAuRcdqRsyH
5RawoQDFcHivg9EcKSdcF/7RmLpIHGEzMKR85TcG4AaidV0iSNnhHbgce3YHv/4I
4iSqPhDQxhnWCLN4t/OZHO7B/7t37zfNPDqMjWy8369cdB+n+37E5Gs+BvQNFQkO
hfAdflrxovt/vgCnZrHX8xJHGCRc0LcEhxzWwnX1Uhbsbf81DR6mNEPmxaL90qQc
7yt8MDDIn1qEYwK2nccIvYnQXp+Dml8IEJb6MmiuSZHTDxR2+dASmU21d+x6dm4o
bSzSjCuvc2v+awtkTfwUsJ2EkyAPIv7n0KV+BvaB0htMTrUM2AeZNEZ6x66Ga2qU
3TKQfWoyGk2HVGL3d/KD5r3FJOPD8GUGWlJVCKVOJszYY+XCr4gg4YrjAWVXoxZq
yjwDF7bLJtzeFL5LJIC96tMgqgtlR2E+CHKCKgE2XgtxbhJQetDg8ZaZdS0d4HIz
8Sw82G4va9VEakO45CPfiJmzODSRd3LUN0nd2gV/Z7FQ4aqRzxdiwvrsU1roKtJp
p2arIF9DMVhIxhU8HPlO64qho5ax38x9dulNfkcFZ2JRh+7XQoTaI3kk0BwibLUE
R21ecQFb5fYmBAnuSUIZbqlkFCuMkHupdmHQLswK79gWqTZM16+1mFotzkNxgFbd
R/xZcppAZ4lLBEGseFs/atKFPZ5h6zCurQnx5dUvVskKbAF2Bbi0CMT8Ev/1aWjf
lLtA+LtYrk8AqF1mkRdFIY889t1F8bdt2w1ZIGYwzU/IDDHb/+q9WT9Qkj1GnzFs
YilpkSFAcUDS9W4lrSQrhoiOEj+nWtjCjbVE9X/0kg3FoLajPL0ud0Ah0D4WUSvu
Ep8nYoqKj1KU+57EVcah+ttS/8uGGYoPTNgZD+2EzYqjiRLRU3dA/KPjwMqg/nMw
7SKm+SH74Dov+cu/Vz16d3l2CaGb1RkGx3UJF/YKu63ihb7Kqsv9+KBloAwe36pg
8tUQhjG/uIcjVGSUuykZx0ABpP08weCAmwTxJ7KLXeexmZpJZxSpphNkuDGoy+aB
80P7oisHqORvyr94OaYKDGk735ZeO8IadEH5/MAHSg0e0LzC1XnCTHHTeAK8PpFm
L2bJl25NKhdTtm66SACfD3XH4I1yyaIUV7csat9v4SESAD6ry5n/0hws+LDov72S
1QN34GfzMQXy8T31oRy6/Etyorl4anhe3cZcAFfe072ROrAHV7crutDt9Q9Ki2yV
7I245v//up2Uy1HS8zNOYARMT+f0WkuMqiczPqI3VfGvE7Gx5qoK+PwCkLTvt09I
lWe51EDFxgbgGHQBH67aCkmG/Jjjeze9xRyZprBaWCzW1ShxlMuGPatMm6Ts+B7D
7ZARrLW7SjS/mysJR3tjEkTg4QPDf24FpI0uoW++wlUCmWV+dTPH4+N4jA+ygAQp
dqK4nGRXtHQAZckWJSVdDxyfbXS+kwo1OSp7PB261oFXXWfgy1PIOKrdmoPbtJMw
fb9MVycpvIAh8MXo6xVtMbeM502PIHnsmVLGB0mOebJkIe+5wnp5EewgrHbw0Psl
jT3h1oh2Tv9ochtmfHRqPYwcF7e9JqIBhOyXJgvrsxVR1xnSSLcNZDzEMN+t1bmQ
LCcG517vOYRBpfBnwRy925PcbU7AxSNnN8MOxEV3afJ1cQLX1VZG0vmIg3ElxPXR
4i9dK9uwubv2KOXyF51xKdJNAGQ4LOcP+j/ps582bzaU8qZ0dHaHXOdYPBMyjS13
64mmEoYedPDgSbsV6kx1PHy4oiyi9us5rrfZE4iOKW5t68grzsJOvYpvf5R1K94G
jhrw3NPZO14thtzkJ+JwR4vR1AlVHpEB5z1AYr57OSSMq+ptjP77B5Z0oeU1W484
LI+hbA9UZ9pg3mFb2zRRSV6HP9OuLnYcvRsowo6f+Gqfzrm1jiNpIBgEFGVzZ27E
C/9kf9VxaskLaDzrwWeLd8csaCc5dycCKIm5qNe7adNpeVfv4dQ2D4pDunaeZuE+
kvSOatdh0XE06pDk4KuzS15TGbyrb9EpjMTPmuQPhTLBDc9wk5/qvfvv3VRIPgyT
oWjDXrWL8/kPrS9NJhg9jFtDSyFPSTRne5yFj0Y/8roIzzFBppdvYXA18H7ov410
Y3T1Nl6oLjfGhGzMsKkJbQ25nDpjgJhlwXuoSudX/uOcNTTjg1TcZFZyQznDNQ2s
fCnRK5zRmheJ7dmhLQ/sqCgzE5ZxWtNwXLZfw1uMV+jvOYpHJqeyvnk1WW69MKfW
xazWlZqqxL/oXYDTgIk6mUAzTWRYrxA47r+ee/0wYYXsmxQx/+Mjqkcv0MYFRyZF
11D2y5wfvRenTr4XuGUDiVowQDjMzH1KxLtI+RBM20NtqVHMii3HLbNZsLnCx1/O
c+Ygzp3/PEj8IEMaStsoB2oauAqL5VpHRsllnviT3U3rJwrzwAnvkJ7bieRpOzSZ
mYiYITwm0lXaYLgutvjxxFiYlBbwAfZp+pmQyYNxN27+w8OEjqTIHiXKCNjyh+ZA
PT3O6iyPnM3K8qw8d9/vpYypt5o56tb+3zuvi1aSdqm7O1gvclh0zh4iD1mr/V0t
e0Z3Ln5lX1bQoi1dOb+Ckn5Er1Zn5iCldsK6PTe3mbX53Kt6nb2bsSXAGKnkmyYH
Fa6ODHgKHXqrMqPQKO+D4UHEOcjAfCoNmuxKFPD7KCpu/oftVYNkitpM+H/7FzUK
NiMqmN++zOdd6oyxEoAOuP5XGyG6XoQ/BZjp345z5PZwmPF/uv8LJRhEOCsUwmPY
pflJcc2vFwG+r1aLt18AjbLSVLGGGwEZwiQDi3c/3yyt4mfWM2jKasbT4DRDqHlV
tValcb41YkEwpS2iWYd7ocy2C4+Uv21GgVJn5R8ZCDXtH6tFE6tDH2HfSH1W5gg+
eU5wJzH5R4P3clRYyVEA7sJ17jgccV9h0ivThok/yi2YuTvYWQW5eOshzUS7UBge
HR8lcv7mOWwMqtJvM/+jfksSB5qO89rx4b9Rl1YhE2/84MYOe7V21KU7ZAmSa98W
FcS0Y8hwKrQ1Q3quvK68x7WspARrv9D5Gm6axeaGB3XLlO7AURRrypEloWWo4EYX
Q2Xox4VdoL6ZnW4AIevZR5de7/RLowzdRROI8keB0knBxGZB0LOm78bViF50if+g
mRDDYgfKWgMUgLiclndX0kyGgsTLTMtkkivhq7/xdd+y3tV88UyzOEYX7tGfdFHg
CyiDQzQWpcVjRL9Ez+P6pAapbVEpYrZwl3wIEnde/uYiID0Af4sV7LyZdx4QRDgO
raJ/MMDtta1JSR8eaE0fB/T/XoOYTx3qLUkJeywZY4Vxi9zxL63gtNVmwPjDYWj4
h+dfdhnmmxNMCqmvIk5PDikOFhKmwAFFEbBrDEhwjHrxp42rCFDZ4nTPcz8Ia7Ip
5+G6BIcE0FUZkH0iRgkRpQDlKvw/FzwWz/7NnrxdnT704jA/xpSAzhsbtDHzFRmp
woD6L36ydDQqV646pq0RMALxHwIQfuvHLazhfMKHmK8RRbJrg5uOhtNFVhD3q98l
tUyk8Lv4+1zsyjLdxBehyvTmODGGx64BfgvIHQTRw/OhGD98STls4jL1usBw1AXH
4Y3rCUyR/8qVtmV5oXEbseKNniWKkXFv0DTFMj1aCtn/6GrtEsEpgmXKfwdRUWFA
PBeRdzpaEdbFsdIpZ8wSHDho1Dl3juho+OXtF2liNivZrc6FTzp5i1KNHWL1iqIc
2eh3O7qDRdx19mtRmfPXEFa8EIv8sq5ACJkDw22X5NqDfd5HKi7q7XPnCriEyykt
CwkWmRgMbE3k07FxI/K4j+4gX8kr0D3DEiJ/fxdoROHbkfmQUDXbASKC0DJFRlrG
vuSTuAKpsS12B1dfRfz3qhXlIyGMTuq9SSmpJnQZoyAQkjb8lfU76RRq+pDSqTxm
DarCxN65Oz3DU9MygKf5/gyHqHrmV/NRVee/WigFvc1C3nmymrwudkhc4oOtrY/A
rP3J6U+xQM/0ixJ8fj/8uXAXfdd4qVk1KnFadyVqbSvJ9eqR+CZLzyM/KsI+2mLF
9pmz5pfWk5jfiYTzMS84St8MGxvCQZaIC09eB0oatecYgje8Suey4LTOgLsvjSZA
8zkQcrYo7h89/6mw+c3Me9XTQMrKZ7rOdJAgIcJzlMGsK0Wd3XF8Im7ABDDDZG5y
XGOw2mEAf0W2Zeo8K2ItHYeZE3ellVVq07XtpIKqYh5Stkz0y7hOeo/Di5DlsXYg
3ZbdHlwFKD5pl6FNRvTklxIoHXxHaYVLUea9DcynyW7jlUCWBklA0RwTzCI+GI+U
hrE+mHj2ONXX0eS4m2A6S66y49gVsUOQZfieG9IGJj2QnZX24sIkBsl+MqF8y3WP
r3cTrXtZiqlNqqmdy/fqHiaIX4GbIsc4znWzXLqa2ulyy2eAivUQt4USprcgxFOa
DrxsC0UoWIxJizGAXl+5VCh4RJcnvWBaQ0Xlcnr0fMz9whc5z11cAYvSD10WIy18
uCKqSikS2nHnNv5vYUBPFy6AC+t8hfuEPATmNCkAbqZ4x9u8rznWKr25JL9/x8Dk
tmVW4zSuU0mcuPx0A9dhn5kJ1SfIP5SjhTtkHncIgX0sUoYPfFLFHbAqJAZK0hUC
O4TdVPQnup5XrO5kx7kIo1vcSm0rwedaa8tX/G/a14sMCllUu+g8jg909J6vrOZX
AFCyql+puqSeZBCEc1slFtYMEOpF9x9xCiq/9oU38HqNt6GxIo48S/S85dHek7On
EYhx1h811UJOXUV9FxFDYT85pGu+cbPlzBd9k9Ixzzloy60eH58rX9cyCK2OXfhp
yTUdQaQ7WHd4H/xFckcCw61rYcxWTQimkRbjBvOTAqx+N8siA3e24yh/AjhqFMNz
hXd/kbkix/tHCstDL1+1ucE/PF0RLMu9NTbvT2E0P08PkwtgGzRP6NzOd9ba1hsm
/pPcu9VCSyNkh4OGQKvEWVWFKO7+vbZAnuJcWJSItPmfr3UTa0Ix3OMET/UPLLKH
5mErT/4Pf3yo+KbgnchkZrIH8bzgUJnkqqaUGng4MRMurve3Jufr725NKlUtaUvl
fI3KtbuKbzEAY+fSjZgFZWtv7T15nYjDfuHnb6TvPV/LDh1H5ZXQH4azaiXbc/ZD
ORT1s7FKB9K0vt7v15iyEbQD/UzhLsKrCsmoNIvfz5n3195wKrR7N89WeiLVL/yp
yyIA5zlmA11X0J+gXnXNOEUhudKcG2gVaXhJhQS9jlbLVBHkyjQPSwJcjnM9A83y
x44AGf8o/AeACEv2vqUq3PQA4rIgGZcaM7b/Woh0slobY5hb8IbSs7JeMkzLVq7/
AqbTQTFlREZTcFT/o2OTzbTrMcCbQDyx6PFIewHcVrjahQ4YtatwRL4mJwvfiJpG
ZkfOaNoJAEKQLSXJ4pnNcd7h2VuWO10xMCHKQg20CeBWNw85QsTbfwW65Mc1f9J5
/idf2Jk2nFcaru4k93gN/jR6rYAZuR/2VYDuWmd5QloKNKX7NlKXuBMgSpV+tG3f
zY0Hss876eeWvzi/AYNgwUP1yKCibI4QIFwcGeiVVzxMmtuqOCTmA8Xd4fnpxvcN
Ysk+N0hP58ySFPJuzE+iz9YTQfHPJAl7xme4CyKAJRP7mz6XW6TdvcbomNC5xGWv
TOgft04Dkcn+4Pi0o/bwf3u1VARM9PWZRd4FQu1tr4+iH6hkYs7XkcL4sZd/TZZ5
n0sQU+eK21SXMrmUkP2ceq80cVHJcv8tgAl1yTAuEggZqj/TDLuK3eJgSVlAGsVN
34SPu5pFpjyOodUuHeGRMNBWfMsMa7ZbCZu6FLpleNuFGzfNxHAFMohb2ZtL1zTM
HBRZMtKSa3KL0XVrbJjq2bf56K5Az5CjpvdgkxWUzwp4ITvySqrqabm3Uupr4Ggf
mfiTKWBAVhUelWTXCWvc1csejzfuy/lFiVCJdMKrj4BSbslGEODwKuEiuxy/odFo
rQLqE94VtcxOMdJfT875nJdpsVcneERYErBnoVFT+dUDqurgqjodFvbuoYd5emql
3wqQtrvA08IjbclFYJAqwlJd+O7WwOhJR0Gabq2sPZy9+tGGe6CkeOEPH+9E+JuL
w64NueMS3H1IQYM+uBRDEkO8arRhBBpXRi2DsG7ECa58N7f13pFVMN4wCeeXwBjA
uK2VRhHw5dTU+/QfzQ23J3O5LFAyY0h3/iS74AjVakVfYVhMKvkJ2g6Gs67sEtKX
o3iigidNk0EDuVOWjjg077UPAEVV83AyudgJwTSIVlWuGo7W9hNpCertr11KmP95
g+iu4uQPXWyDyFXuZMJWoYCyTdl2k0WcRrlzS5f5MDRvAf6bdQwW1THqHFdbHqM6
1zaeSZLIj5+cl+MirVmANUOTXi4a9zKAHAr1XMyJhdDHWrMnKwfU0Pve9OjQ4deC
vAi9+kNAPaJ6aUKtroUuFehvUPwMliiykM2k6NKjTcc5j3xttv7eJv8U7pT0VfVL
93EhMl/qZfe7u5TkZY6FnbjSiZvFlkbIsBnIoxNnVB0cSgDaLjb7rwkthI2g8nJT
EQ2uSnq2yxH6rLDCyjTmujEyzCKo7dhLN1+zcKFrtq6MTf/DmD9F6PVN4RZTWEPK
PKebiHSkUGXCYSO/I+4ejp8oG1bZ3pX6843RZCHm4iplzy45aOOn0QPgx7hnFChf
ns2A7YbbKm5gQiP3cWbm0rWHDtx9odHW25Sw11rJyxSUVkqtEF1J2R9ljXxLXJZk
0viZknN/Ium2347ucE5/dil2rZuP8+pKzxLgkuMCRMSua3kf5HadEb6k/yUW16Sf
GHiOw5uT6hHyaDn5nxeVxxUlROz3hAFrnwUZhQEMrDLZVEXUOptOR2OKxGaWLp/g
ZDxsCaqHxZZwbcWH2DhxDYRWFu2HXVNrsqkwcEuGdv+YSOTq7k+Jls4uGPNO77gb
cPdy21yFg8o97xYaJNWF96/td2NHjtCoZ8g5bIjKIpy6sE5Q+axyhhp5gF5zhvuD
jNDtxC/Lo8MhQb5/FNpd9hZeGA19NZhKgdshLDDtyIJvXWhCRMJhTKXLJWn0MmNg
dajnWYs/ensmHoAua/WsmQgnwQAV/sO2qnOIGExJ4anYyp9Tx6ZJKmRiN6Ntj76U
kCxFu4wWbVF0fmEBI3zGqpfcs0fVaqgQg/BJrrBfHp3ECoFi0vPgpt9Np1285Bja
NFZJMtAA+iydYs2olnscXEXC7Jir5PftzZys3EdrIrr3mvWbjVp5hhdXbc9Rxshu
xg+dBxHMNvDvw1RrHpYHtyCc9kpvQH3GiXVssjPOQWyaHhR/IMiox5LUQdZvE9Ri
Gvv7IgNNdkmkSP9RjQVAOncxBmpZK07Ze+l2PG00U4W7LtLnmetPPFjnzux7gySu
2pdDKTNF37LkTITxXU9mWJXs4aXn8AXlrSIygYWO0PxU99FVOZRheLYFKlApAhBA
XsXjrlq2Kz+6MmvVlfNgcp4aVgB6ABQI+6Lthic0abF86tEAUodL5G9yDhaEvvFa
5OB6oFJu0HMv3DkMF5F2a4y7JMDWSa4BB10BGjr6Y1JL3vmBJjoXxxKj163szE0c
LtgaodrFULpRkTzPCL3/dpzpgsViqpz80thGQT8qJGnwhFO68qE+XppUiZ8DhGRV
Mfd8kE1WKuQ7sAaErQyXcFFajVorIZkouTGMFTmCS3k+xHuSLG6qUZF06noEn1gJ
vDoskFEimgbrs4PkpbA84bfIEWrTJKE9CoXFWq6w0NgakxDzByA/voWjf6scx8tN
SCnVhTW6O5eIhnOyKMAaLAsrbrh/LCnBZknrzM1u2lJSyPOOZWtkbBIkmyHE08mx
MBmRRKK2nK2pXrAaGsoSUqoO0OHry4VFdd6wuQouoY1wVlkVM2FbjQBkzEv0tGsk
V7sMPTGsnQV3/AeQqmBhZ4h/e60NMAdxUN45hHQ7yeqw7KPHdnaNrTnW+MtvQde2
FBzs81eYPXLQALxPw3NBVZxqmXIfWYcRYGZ0byG1GIykWTpruO6e9Ig+6FmuqqCk
+7XLha56PYGH52OyeOeonYX64Cma42HULnXVB5xNwlXn6ywFbCgT29dtVmH5YUGc
3AUy8a3nEQkBjchBI6/k+fbOu92djXhLMubf7/czKxZ5acgYNrCD0jeFmwCTiXLd
yvHFwpbv0wrZYvq8qwShf83LnobEcVwFLLOGqhJXCfs+7F5pXOG2zqxOFvGAz8Wc
KTz4G+mA3YXYYC7v3pDNsjlk4LM9rG7d/rrL1YwJjCfBUwzUsj5KCUkLPg4o6Qeb
vDKoc0Ak82fArCuU5a7qNTKKwxxVA/RxAJ90iYYhzwsmETRJ3HuOKWTyIaFUXP9U
WqdML5DPaQcxMGyu1+Jya5sqdVFMhISEFpLkwspBEmHrZqhSEZ4lpytvcyTaXe9v
F+OaMDXhIYCHfBV+M2IXPo39fnxfrv8ME11QdS0jlevw4xclkINdnzj452jB/wes
UR0mpIcV99IHzn697Sp2FD2B/5cNZ1PoYCZHrOhKW3ItrBGMnWzRoGiuVrvWC9n1
tQ7XP/0XILobfMw5Gpaolh52udTBirGwS+m12F1ii6cotxGToI4xZV5PbVJhaRjS
A2Ibj81hO4Xa7JJNH1Aa2/NXcGen9EVfRcmwsnS+lm+VPHiZLshithp+nj2vEzgE
5a9Pr/Xab6EXzpH/8iTObUIVowBYp7JN98xs13p4ag8eiNm5u6UO/xiA0FVTfKlD
QH3s/nLKDgBALmOWCyxOWHXZINDG4SamLkyHpFRgrFPkE/xLcGu3VygxrBePckvc
lw70KJYNh8NG68PH4oGIPsmLH/ONvB/HwesYkI27vSZfE5/NpYpiR00dV31SV5Ij
fc7RgT0kt7wyddpL7/ALIZzMoemKEeqShkaxh+8iGnE3kxxm4/3JQ7Hzg8pubpuA
jZizZv46CASOAexLZWwmIuxTru342qQ4kbqDbUyN37gvVW3ysPBNDipOORX7/P4J
8v64Fvgwb3KpLkbsvhQGzqvWQpa2/WL9KfgWezbxq6/FtddirgpQMB1EaRCW6VQb
yROnnjb/4VCkCWDv0WuFHxE1Ci9n+zWRBpMJ4U1DAlhCtQbJCDg8HAj/47++QG/C
a1WWSr0gyl0swvxJ5PjGXHMgGdmAxlEBMWW7jMBpGmq91HVlhcgdm4Ds5jlOCK6J
85k4jyGvCtAzIDPc1+zwNYFaRQklYJ8qQJng6puJWPS2T71ZMsjN8X/avRJKWtVH
5WC4A390C6aNZVkbkG55hlp8qA3nhYL2s9N3lW5wmIZFM7ZSx+KlJK8NBL83iPbK
pPolZVjDcvzmwxE9pYrSdWDnJS8fD/EioA21/+VGHPaAQ588mHk5aAaLlg9p/lkU
dZneLu7Ht4dWSGFxPUpHlMsXX1Eeww7SQR5WEdyO2cQeBKlfI1rXKm0lr417+Hri
dsTRRzxW6RVwPFrfWjwOH+blcKFfY2nXVt2/3h5pS4wWf5NAgc8HE4Jp6FWxuJRW
rUqWvTD4asIWCxro8Kkppu75en15qlqbqwKVxlwWddNIHl71vIJrHAVh5ArAy8iV
xrYjQrWVWTEFBGTBs0+owWWKAMNeurwBDtbmmWFiaTwwiE6VGkeNJqNklpvZAUHz
V8MItaeatNPSz5iqTyGZo2kvhbpbL+uiYqXBnkRiJIwVcNV3uoIUrA+i8PWX7yf/
+vog0LlXtE4TbqNlB16UnAfDCFdR8KgCIMMvqXr636vGs3n/0o8QwLY2uhGKfTVi
IDFxYo/tY68TSAzMYD8nxb74BbVRV+vuT41Nz2f/Zu4dPHmBi898aesb2NY6Cg1K
2a4YpxaY6J+VM4l8MxO66tw+sU6eNUjgPava05SOwzNykxkOHsUvLNYsWWRKpXM8
4E2HvIXIe2EmX6iWG7jn3200MuW9OrSFqJoH+K6HCSmzk06lt6w7hXda0VhZu5IL
GKefdSiaCoJ/eCaBCkE1QcxWiLVqI0ybnkd954JVM4f5QujJ5fmuzf6t8VueVcFx
ZWC92/6z5zle7PD4WTIqHeU1cDyZc+nj3kYCgbMb7DIbZVASDiEJe6JaWu85HkpU
1aqzC8/gnnnK8iK6LgKwnhiGP3MKvEQpZw6tWzbZX1z08wchAfy3uzXKKUnhDopO
8odoBKA+1X6rdO2qW8+hthXZtYTKRmsNyDp78fIUkKX7mPX0JPHXwBYpruu9uO/3
G7u4kw+w9wz01nOgeBh87cTnzl1srLAFWdLoh+noB8KMCMe1MjxpffkILI9T3hpo
1HhhYd3Uij4rJvU+naVCwbpJRsflPrPW95XFQ125mx8xzREtxqLquGh0+KGqd3pE
EyNQICRL5zyhzUhSS/s+1FSwXP3Af/DTOWwN7fLVg2+xpNf7Pr+9dUSxqAJNMLgD
Sw16aoWVnpAK0xETKoH9qOqJb/78xl5iBKcx8TWmz9B0RT8omCHzPQ3TfBe+Pm0n
qYylmRYXgpIzK4ylzRhbOGf0tbrE3x1EftYXOl98fUshRNLYVeOkVY1lJZ50C9Rn
kGqOM7E8V7jfOnoIp9XHtUZw58jkC1Rgshltur3n8lqzcwly+Enjuf/ScAa565QO
bsIoO30K8wdzpUSlVI9qP4v2DvYQidWEhgWZbd01+42CwZfHnZKohYRZVbhincjY
yx3Z1o2iioszre3/5u8tV5uGNyJBs5QpppG+ETEpb2d9bEu7plvtyO+8Ib/Optcs
2XanLGcwD746ySMAGKrDAetcaQK/N/KD7It44HjlPWACMMFxrjm8Rnl6ADFyvk1/
`protect END_PROTECTED
