`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0VnT5SvtUarSkxy1Dku0o2YJwPf+mWDVUflD9lNG/6WZTmpZb2PdH9mAFHHSAlc
NvYkaSqxMkUVb3roxNAQLjjjn91HpRKXqsX4JGK/nSe/4ld8BX2+CRJ9xAGntBFY
Ew3AYA0zrk/5m43+3mAst99BHnf3aa3nkBEBo3oRbwfZVVW3y0Zx3XAXFUdEnsFC
PItuTuZxIEJS+IDDlr/OEX4HYVIx2bxf+hbhSxlUzSVlJDMF1jVWFg/48+tcXWrc
cEtBgcJx0n9DHlNK1AvfoMgnYL5J3vV4VeoZWjxsLX7lUO930wUg+ljhbZ552W5U
Qri6DWT4GGJQLn+iVGyPpAjMZcLquSU5un+OCe4RLoY=
`protect END_PROTECTED
