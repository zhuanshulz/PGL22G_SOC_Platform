`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9VzWkfpUyYNxnx2SDQV1yFvNJMuok1SlTFQHUSTkKv3vCi27WkBUi51CEkeNIdXf
/MPFPaojaUR34ioy6mY5d1e+NjJJKsQbwJtC67oR66mqOMWkclarJHKo7lhdGnZG
KqUlmYg1RRJAA9cGRhPC2lYa41TgnMdMvpVKfu7Bw3ABdPC7A98Q9YOcPT4xlvGb
YWGnxwKIXXcUrbQtNjuuipYSK6paztXbw8irszXFxeHBtwjF8Y4G+VPk8EImBBF/
ovSePvlb3Z6XQNRPfCeGcvC7GRGJhEmhvXl4U1iXvCRlUv/RXp1sYn8VtSub12o8
Rfqvf/k3xDmVJ49pSDpFNz7cYsXSEsHLyLGUdY/khgBiGooiCxwGnBRIFWTvNPis
aYw2VRCRqB6AJuZAdO50YmSR999sY0dJkydIpzBt6SvkqaYNFhQ8JZsOpLF2bD6C
Cn7GrdbXo203VXaQbqixBTHWKwqLxplHBBNCXyLEgoAzKKwtatHPaJufVG4Fw6rc
vUeNMz6d8sQjJ7EFhrTj0g==
`protect END_PROTECTED
