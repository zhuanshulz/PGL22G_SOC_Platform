`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCiwBw3yW5Ya1W/nDi1zY07PXixksMcgcZgW+3jmcSWMcuMeqezdbjCSC1k6UsGk
R3Kl0fwOLik23xW7B6giLIQS2+2wLqZ1iV24KAtdOnxSLgO0Gw/ZRS46MJ/z4tYo
x4c2+UNN7V9QWXOClXPYFc+nHWSy7uhWq3ZyEHn/0edjs9keE9KZ8zfforpFTMKN
7Fvf/lYHUiHx43xpPsK/oXIDWF6V4zZbEOUW0nv62nL2IaklnQtThWLcE9rdUPih
zEhHmCE5oa7wS3K8ZacvtSYS+8GqjnuybePH2pwk3qclYwnfekgBe68SRr23w4WZ
d8JsfrI1JwteP5JAC96ojWjaD0C2m1piquOQngN41JI+U0hKs0Fu22ywIpYrVNHo
8cg2Dg1B6qPcJ5xKv5l29T3QElzi7FCrUCC2VQRKJxmvIEgxzQJv5vphTZWO3P/O
qPY4sfnIjtBQDLpw8Rtj0pVmsrrTT0NVEc9zYYjcdSvg7v5vKLPPX87faDZkxwNE
aLM8NNVGIS2lTByzK9mJJLaY2mLcDKmyO4w1s0hwRppE7q490vhq9dpBPJoVOJy1
wo6TT6mFsocO7NdIlET/3uXJMgFwDBTRQiyC3hdYzXHK83+mj8OItDsjG+nCg1/P
rNTQx4uh92TS0j3rxgnNAwbAJFElJC7A/HfAynhhA9TkG2qU66FBhTOroPj36wxu
NpmXLTh267KdPRpfObMgcXvL224pQ99ie98x7VuM6yCbbHyuUje0miiszYYlSipw
/CpwYIv+oJjTlHhUXoGP0nFl54SHEu8sqKEhePC0RF+GGKrSROy74nW/9F3m/DUL
HaLQRDL/08fkCJWEOdB+Y2wUSaYltDvDgdrOTXshZnkNEKFWyBDtOnsxzesXZTl/
yC4nYbUV67MnyGdobz/2ZhaofF4LWnDwJYd4fXUIuyvhjbHP7RO4ptycL5HkabWL
w+MwepK5VL/FT7eCVVAJGjONgPEm9MF1BAPmMRrq1vzDG2wnBBNmQXfdm3woyy5N
PbUCbjfqiDOlWqSR2TqAdEAdXRT5ena3UKwi5hjtBpDbV1MQO1n82oi1YZ482FsC
Xrw4ftVM00QMcr6tJCww2AfPeTp2LfCZdYp9A/rCJKeW0tr0ejmGhpYkw4W/aWMY
xOCPY/QRePyyisN4SvBnuD9R0vDFfsyZNQf6Ee62cxemkEcH3sAMtkzstncCcssl
aQfKPBGvsyxHDoo2gf/PVX3KC0Wdr2GNEgmDOok+MI9438mRLYJfzos5cjyzLbWU
KnmK9vV4QAee2KNaNG9b1wmMy8jF57JIstxnhrwozAvRPVp/RooBO/sU3BdEjvzp
+Ue2rh4/WYO59yMfve9/OYxc6uxZVF+pZOIgHhQ0NmPPsKxVSGOJ15ChK29K048y
u9l/3vpCJ6TuNYbwAJwE8wjHkgFkmWIKS6pjnORb17Y=
`protect END_PROTECTED
