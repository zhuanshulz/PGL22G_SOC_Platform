`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jz8dthytYdF63EmHRUse0T8mxIQkdJyrBgvkw19dxNcd+SK1pRNIJECNxs6AmkIR
y66SkrcK1p01+CZM7axKnhppm5cFdYpDXBs+/jTx32gg73nTmXxrjjNxchfmg4ni
IwOqMSexKDI0zQ65M2rIeriAz9p0CZuPG/udSPG6kP8aMc76dyr0Wt9/EUsZySRC
G0cu8T1F+9mjl1PYrJ2sNWMfLV6pcXSZYINq9eT9lMVO02EeuzYeUDoLiAcghxyK
3GxMcwQXh2qUs1ooGYglKEqdkWg/vMWbEBbh8FA6Sx4Rse/Ulvbutzg6YVc+DiL/
+LzL/FPYuX4owztFLihXxUy/nZrp6VUtD2hKQ3CmmhbuI5zfNjTvFsl0J3L5J8ew
BE4OnbTRSLloMAGjwNT6NJ5sr/Ijoiyx3yuP9Wg7qM9fMpaRPdWO7Bc5iQCbiilm
TE9ds/0fHyWPsGT2L/d6rtAaS/A4wds1CSU+oqxYqq5D3Q0jLvgFmW/pF5PDpBSA
2fDjmUKL0F/BUtPdI8gaFa1WTx52NfsFSqXJrs86ikLY9IMsNIff5A7sSKDNBrZ6
Lzil5tdQPI5sqSXM3ZwKWUSz8tOc+nRppEKVtqxvtiiL59JEt0IRw4tennISJHYc
zD9P1K+D6ZPCoyo2p6rAKHeIBPNZGgYris02ZlDEXftinpnE6oXzEpHZwWYriKzQ
dgWuUiWhASP6b4QtDBhQFkL3NJulyIttzDf0tuhAVugrNDxbRd1Tv9D5i6Y/9kOD
h2f13ea+8vukSKZFX4+FeaDCyMXRSRuJ6xf+/b+zuiBg+DHt1pDVjuHsfERG3LsV
`protect END_PROTECTED
