`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CLXiJ6sRpG6ZFpTEqm409NC8OzrVZYQiCogxsgsX7fDGbyrcuVW0wKXodmmsU57H
uktrts+ex+/X3y0Icak+Bw2N3wboaEaF5zTPJRRQ5JuLmo7hcQ3YXt/2mDiW9neR
tJY3Oi9Bi8KdV1M5HhGCjbcipaf0vvTaD6iQerv9tpGCzFwzmBA6y9ZBhrwvBz/y
U5yh6YTf7xSD6mZa1fg6QVtizoHLGtX8X7xK1gcDOI7CmCkPY2+j1ExPS/fyeC8C
j0qHTOkABg05C62GqY7JsuOow9p8eUYuUOazigpzVzNma72AXtm+6j94pjwsPqLp
H2VCL+hmAac+ACOVKUdrMkiycDsVf+kYkcnG2jEjqtukbRax6m5f/t9QtX8FMMyc
soCW3+UGaP8SRpM8iCuRR8t8fEsFHSta2LWwWiYpAKN2bqReTA/G/GCc5XwfVRxQ
OV/kB5SaPLYeLgVspD1rgmSweu2YFrD3aCLOTHG1PiVBMUYmbwuZvnCTnl9Zw3PW
hE+u5ecPcK+xuieNfwfYDV0VtA4x+Gft811gBtjTbXBqIVN6IWDyQx+i8RimEkGj
Dd7JKh/W+g7RrkSNcW8jXmU5nm+S/YsMtdRILNhk5GN0Ie6G16Lw4fGSmvJC0tNT
VbPSKFeuvldh0Di4Kzqe1Jn/rXM8TX+dhfpkR82G0zpJHoYAzmfSkIN9in0IYD5U
khbkPXdpbAkOHB3O+0rdscr7Pua1t/wpXqPrqMXT7oomxaawGnVLN1K60MUZFd4p
+z4Go1jjCN3o1kXuj8wHAJ8bKWgehP53J8481pTaqJoAOYNZnQzimIuiiANxWGh4
pxjqWidKDSfgvKMKe+fYYNmP1Qmte38Mzbyz7btWsCs6Hndcv7U811syUFVsXCCh
ANey43iFUUQX5ZuWX+3cXw==
`protect END_PROTECTED
