`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ov9ABNZRIfFJIaXivE+FgkSU24nHossWPYhZ67Un++xXai5Lk7xqeh/sG4ki6vbW
yHTDj8JdoS/jIxO4hNMx2Q+NQn7qYZy39WnedNUuPgajgaK2ddWqR9GXkLoWl+aH
+yq9NcsNuvsbG//EaIfeN9RQI3LAYO2V1JGxrIrhXA7QgwrA975rvjUwVrmdiLsv
1WRJIs0iluua5eONXq/2dSDdllccC3pOCvjKAG5iXH4fr5hPSSR3uB4m5px7H2mM
D69nlPknw7Jhjlbsd0N5OkIK7pS/+LjdZXJky6vvOG/iB961oeBl/ElOCrK6qhK/
un/teM4lADIFEIE+jEbr6UzlAVZAokxFDENzcKGZprCdS+Wv3eFMjX6emqJdYUUc
zOdR1Dnni70OxsPOaRGFsB+vPqZAK0jIcnPELBe22IsQfXZk2N/YpoPOrECzJACt
XEtfUP2r7++iJ3X2ZlR2vnXYbFsiWWGdm4gA4oeqVgAOhHngWMrm0UnQtr4QQHIz
9JAz7dpA2dQVDp0f7IbxaZGxZ+TXOD0ehE4rgNDQrDWwOA+1fVJLMraQSOFoP8gZ
dKhdwTSZkrDPzPhKiPQ82CXn0PfniCVsg0VmLXc00UPn/qrWWAJaYIZjNg2Xf1KQ
TCiu8+r5yYKcfLcAPRsr09xJ69SegkrxhTZeqLT4pmuFGjtIBdN4cP/XyGmuxlRT
bXE9ftb60PECBaKDguuLOlMudUDyx1evzp7lDm/sTebxmcaDqbClcSK1+etEnRLn
YXtWVO7WqLpzUbXQ23T1cTP0+0CmNG8yegEUmyPUxKRb6ZB4sVc4/jNDyqkzEZU1
kP5ZdoTKKhA10KmB5M1MTReb3yQ7NOYeWQDASqJa3CkhmGGiKUnhMPXqxXpA9mgg
CJghrAqZktkJOqNbhBft3DwVmn+jxVwfe6O7B3rtSX36tfA7DTXoQGVUfhSGV/nt
GxBmQHQY/0/urG+YaEfWD4Pod8mgzlvU6d/HpKZWmorCxZTqwmnWJubQTTfkGAlH
6KUuAS4xTjyv3Qf3cNp37/FElI8fkwhE9JYkkthfW9BbffRaBERPZCNI6qdZro7B
tDfqISLChqy4pRr/4U65uEzZkEwXbcXD4fnRcdKPllv0tcKmmdRtGsv4kTkin1uH
OVotiRZe9SKh1Txf+uPvT/tV0B+eO+95tVpURTkkahluBTUiV3XkEyZ5SgUpu1g5
083JOQCvOIN6Gy1fDCHuyS3hmeUpdb8aFCuaZlHXEpdxvi26vpoYcYbOR834GLul
uJY3ttXVHeriz6Hh5u2rm561YqIdTMewfqyuPfYpP/MDVVqXZFOtbAvGkFYQBElw
WUVasSztNJT4BhX5H3AHiMrWaThLv+mySwesohe2oKSO8zLqtgData41KQxrxQhY
Ea/hFhhCS0ZPcv4cSpWljBHLLOXUHzOPCUqus+p7ob5n9cMKu4L+q4CLpBDqL400
fEVjQ5WgRHeSrUh6AB9lV9TbRPCA7aUvMn302yWczco0rUTCSlOGfL4diw5Mvx8i
TAp+kOBOiv3ZH42C/bEI6lcJ2OcF29GfkwU2BU7c9CEC9m9+Zp8dpo2ED+l0/nmq
d888Mwi7MB70Okhek7JG7tV4L0I3e10ttk15eA98BjwafWZhW5cJEwcxO+4gURaP
U8LAorWMhnVAb7iZZQI7EU+/zsKl38JUfptF+s9gz7fFT1/0ENJ18UR6kKt2VsVh
XSezvG5SIs01DIO8bvqFxS0gMWmom6OvesBHuoLRpa5o+T2884/qo89MAH9aNA8l
qF+4xG8JeFyX2lXPgr55zimiwWRom3C88hGel15mCWJXiilGcU+QP7ZUgn6Obhgk
8YSki9lZI69+aenH76J/+CTg8liZImel+13bVv9SgdTMIELchKlNIxrinESSk5kd
8LdJTjV5ayVLAbzpWjnf5K2NDWlqXwwDjWsG2fC5yM5iJqOFlOIFV9bGS/PKiSlt
DMw8+DG/Pr/fLTkSLoM/rYFhhwZlAdyx730tZn2MctkfErR5DQi1Wxys+JgGd3pP
sE3OxA+a1CQtggaiYzMAfG9B0xjGlZ+0PdmXzRvbvAPJo7UJMmICaJMPyvUCFGuE
fKCDxiwgsm5h36nNUfP/Ixlb9Rizc6w7Cni2oCyrAq2hVF6++QSZsXxrtsbRgNFH
zcbGUjYtCEW2iZUXVdMbpcmvutpye4Qo3v76WYDGPGBVNiPIlVLmdnE9jYR4fUJG
foeL7pWo1XaBy+GJhdD9g1Phr+f6pr6sBac3yWRBjjrfMUMYeGL3rOOq/bPJe7WT
QsVe5O+eNfWHE42++W/+S/ENfedxPV42wUPfCrBLcgylMfmuSpqLHqpgdnnlyvMt
3Qga2Bpjy8NrA7MlEJM53bxYQ7LLD3vFjijXz12pfZrs+tRmQqbJfHSpeexF+ABz
XIemBtd6GZRKzUKMoSzSAaDGdh6MLMvQE9tPJLMAAEsRPGadISaJ8/SZLrnzMrOf
HDSPG4ioGmRLTmkeZd8yM0OIuq6ZoiHQMTRnueUoZK4=
`protect END_PROTECTED
