`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pp+c/muscLAavnK5CuoUcuM1XzOGXnMxWUOKdxwOiqIdVTiuY1vshUdwvE8XUIq8
mrneRdha0NhsiUMAmzp3jjZnnqgANcODsArezrS/Yz1ZHcroe0gyMa7kMJzzK7K/
a9xvgHGNvtbIPFSvFZX6Kl6E+OTjbZ3dFrPTPgss6/SIrnF5uMED+Ob3okmG9UYb
ZlKZ/tR2Wnl7a9YvIOItTyCzMwX2go+9YiKl/3yoSPCWPePEY2IfDwnFodDEcC6m
1nXIdsoVm+tZ2zQS6v8kTdtkyq32T1i1cVZaVxIv3sgybhBJ0X+ERaXiZcX35f/K
t1J2vrY6M/rs8G7BEPNI9EXiYOMOPBoucaCiRYwZ/VkRs+LLl9gpOl+MOHIMuBhT
Ss7ryU8FmsKlk91WMJlsB+dc+pz/MD6kmFLj8kuOtsSkGmJ9W2GOcAcdxRrGd8dG
umuAZ01LSD//m7SzsvRjX/RBBDHaVHScr1tw4ySyWj1rIyPaUuUFQghV1OSLecEc
2n92oe0tatggO6QzDzQsbA==
`protect END_PROTECTED
