`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIDbvJXcJ8422gSQXxYJuPFepM4aWtbHZnRmghZVZRlJu8rLvCJ++HX6vZg/4EQw
h0wrpIENQlapUwkhc0/bd9DrQtop/IkOdT6vebUPOuozWEEVvawB1glwIUP4T+rD
EffrLn7KFJjo9JK5x0euRR/IGM4XwkoSFguYi5hL5hGw43ZWPs3W2Q28NZIzhCE/
9eYs2FF2pvl/wShPgLQFCa93m4SDY+CeAa/WcPWTbL9INm+SEW9+stTM5BKQMYnF
kiYhhmaNEbym84+W4ISIsiXxeArHFRJ+d3l7u4f0ien9/fXCwkvHcWmDdavf/yC0
dV3Wi/09fmCa0e9H63AWlq+5XecSv7StEuEZQu1jLBZ/42RlaxD7b6zuVifIUNoy
VnoQior2Ln9hq+46DgcW7l+1dx1+kTDtQn0iPDgu+gTMkmn6dEJvvO1QLMCibuWx
iCfwt2N7GWsMYm2Hh1Ro9ftWNt0T3v1TpeozYwHa39ocnMWwHLO7gqC7elHKYn96
yr8OPX7LT0Zh7mgmKGZASaGwZMqI+YhjOQ7ZYd+vJaACccVFSlANmCbNsCMOKpMY
AAVQr1loUuB2pZSOd3Wgc/9WRj5eRiRDH59ohIB3IDnODmjOJC7/zi/Wo5U7+DLV
f4KpEhodFKrPznBRddqh1LiHN/RK7Zry6KyTdbV0Vg4KpZ+SFUdI7sNTMdSpWWMk
pSl/vi2zWLYdcjwLFO+KSV1urZvux3Vjg00gbawE8wU7+zaH4dGkcMc2M+zoZBwH
x8Y1Q6jQInvMEL/XCt/cHtzHHOl5pg3CVdBk235c5nIbalmdLl3Bz/ZBRGBkZwNv
9Ejpf9hrITD0yjWOa9uUjgQya0ca5XdnmeFWNSwzUdMXQuMIKOzmfnRT8R9HYWYw
rRMPRNXSWlf41NwGtW5R+RuOQWhLDQ6V6rfbj2LhCnFdjfCvUKaTYyFAi3PZAAJ+
yxoRywh4vWGEd6SgqhYIbiD6dE0m+W9vcUPPOgmJhjNVMhT81FHO+O8kTBuMZsx8
94pcMpcUXpVzM0imonCMAUSngdkEdsKT93ul7LwXmmSJDKs2cx7l6RaszlfqaIK5
oKfHbZoD9xtiMj2Svyh2AANR7BrgcwB8gCW0CmrWCoGoagxNKshFgbnOtOKtfKRP
hSzGSZ2Cr2gVsvCJ/MxcEAmb8aUMeTV0YiMdPMpBm8L5HOdKFS8h1LL5Zf9uDaCi
eKZlD+qai7w6qKD0fVUw8M0G2LXzI+wG/MuzmnfJj5WArHUab/0rjYU2mUA8bnw0
nHpxxch8RzkgTYJjjhMrxHY09Vs1rWHhcwRU4uFPyd2OiXblwdhpYoXpJLnQk3B4
7EjRDTuBhy49xNOqJCGJfCiVTQbJr+4wyyQQjUhTp7OZtRLfg92yHEJpdw/9ynHQ
h9pxA5eh+GS8+gPWFG0xWEBdRX31r0gW7Qri2W5PFrZc3YMpNpDqs67tBdCLhe3N
dI3RhO8TK6zcoUyQSrTy4eAD+CqxWj1GOP0n5uePxHZbpF47qSKNSdFhSCRcdptF
XiopqoRgk0gkT89Z1eJz9/KDND8YtUuSvgaGbEa5zFSjgHViKiFWSu8ogUAtOZNN
yUSL5LGsSu9r42iynjkI0ZhbjAbrKhYp4Yj2oEv31eUkJc7XchgbuermWBjrgimk
ARR5x1nXsaSK0ugXOGcre6+N+sMPZAIxjPajPZ7Z2kSkuTJHWLCQuMmk+C+uUzSQ
0KJDLnTnroQKa9AaTlykeJYKgiT46i7KXenDxgdxo7YefpQcDKejk05UGuxSstOc
DRNfvk9U8RWmHmvBP/dKZ1hCtqyzLokGKo5wZGAhboKC5HU7UeOwOAIZE90RQXP2
Q34EeHxCasljOSKbKRiXpVOFnS8h+ruXLmr1m+mX/yDxXEydItBznJ18mwoQzCwq
6wn8xNde9DbrjYAscPkXPULauEC9T4+QnflQakgp7k8Ud7Q+OSAKbTgnqRYkx4+7
IKzpzil6uIZKK/TTeQ4ZANB3R6dYc02KI0H01iRktaywhnUjVgKH/S4xnnzl1+L3
2OC75lOdT/RJitvx90v6RKvF+Zj8aRxxjfuvbbzZcuP15s6adha1K0vYVTvQlqfV
JwDTRz2A1Mk1kw8uuyAWQAlAagy9/VYxuWamP33e2Q3qQb+OkMk9cGxf1rEYtLjP
Rzo8Oavh9kBrBbjZtiJBeN8JzqOJz6ZQlLLlYbkEticI4xpKjfrD0YQFu28Qosrv
rP00T47o3SZI8JXrLuK8gbtBPBXM22Vd8c0ut76dNTTsQOq6ED16VENBGYtIA7kK
FECc3c/UjDgKZ/jl7DP/s/f+ogFn9c+/J5ljW+uHoz9LLIfVsBzQOQGV3GFx6rW7
rubwUlhilLV89nWRx+FwDK9idz2oMZrT8RgnxH6hL9TF5YG+r+UKGD2XbvLlhgoA
rL6iljfcP0HtU2DpAuRwvhMC+H6rfxgDU7iJ1RIwp8cDjWNNSpQRCPwdhTcwF47G
h1DObrCu5NFElxscKGutnW4wtAaJzF3eIyuH8SDBPOxfu3kjM9bfnrcKSp2Q5Ard
7obugziKw/kfMFrj0DYHRLBFTIeH7fj1SjRRH6aP0PtzSAWW2F10BxAqHAz6LcR1
xxRmHyIt/MO4lvrvER0ckY50woc++ES9+L94kDrZLjbUDmIFKIEDltX0xEh4JTxC
jVT7hHRNtzK8nqiQmBe01fbTLCdXqKs5WZ+xvTqNCH4vYeMuBH/HSjrJBGNpsvZd
RpzzA7SHu17tcKjnQINT0OTKxvHmY3HsK/xjAy0e794qhDEx7YtT7s+K4mpBzwMi
G0mQG6CIRo+AP49RHac0M5pBgy1pcXsp1uOIfJBMDRnr3OfwnrRZOx2+L/LZbUaq
plWASa00SoZdgVBVs7VeHorxkBvhQHH4R1EgpRAWm5VchoQJBcA9X4oiXPAPJp1a
klY27ApuAl4JNKJlq57TDO762380zYEEe3qd4vhlx7OjSCAI6MBSagfbr9Adbl4Y
L0ga7CPN1AQe8jy6izhnnOHt6+8JkjWf0kht2SCpV0/Q4UQgIpsan3luHzL4609m
bqwSvF1JPesc4W108XoAl3pbMMIX7lhPPK7Q1Lp5VmxfxdNR+PrXMbXb082G1d41
KL52cXI/mS+bA6aHB4uDCmqwiorfR+o4grOaATGoqApZJNG0+mXsVe7zSU4LLppR
NBiRCUzECZnxVOocf7nImF97ZhMTssGf6T3tvb9Xisj3D3Q+MOUZ2B0RUyMrCu+U
hP2WheANanpin2fdNGgmRf/20GPvv7FSiw+RBmbLpRLF5Rkt7ehOdnXoklfBkD5m
`protect END_PROTECTED
