`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YoE5neyl0kUrPHjo1+V3m99hT5SyVfQAOuffPcteoF7Uoqtcxwrn9AtceQm1ifvS
NW0VD5B3XOMiO+rsrh9Ncdr/jR7crs93aYvB3ivuoXratNyD/1urhk/xzEmBK1ya
4NqZPUVNjDle2qkrM4GB4rcIXUK1Xm2ad0NzQqyVDfFdIaF3V1LyhPB9rlXW6FL7
e8C4QEsxsoRVW+2xlOoATf7avFakiGXvOw4N7YWGHqjr88BY9O5NH4yY2fILyCRl
GBlXbsiCCVcZTy9pvUZelV5xlWN53E2tJt8bhSXj2EIr906n79Eko5a3vCNHOCKY
3Aj1KbByoOvYGvfmt4FFST6F+hSIfbEJNhYZOOTrXd/067dNPaIXsEJyCoPA0t90
n4lFfBP2Z33nNk6jD1ej1ktQITmqnJvqLS8lubK8hV6nscInS+oYa8NBOVLlM9na
u5FSz6lex1u+ozTEsKYH0q1L36UsZt7l60qmK0/lID1VNb/VBxaBNnJM32JlabVM
DjKjFgCmDoeMICtOlJJjl3wDag/P3igIwLUO2H6+kM3IZ42qeNSCgYFSUGJdMOYH
`protect END_PROTECTED
