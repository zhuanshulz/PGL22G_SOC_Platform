`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnWjvL1T74CKpPVfzArS+7xXFb7WwCLzPLmJoLoWXGYrZRj+NSFkegxdVrddKNRu
FX2aKFzz6c8LGUu40tYKBt6QzsdlxcK6VfPfReVNGG6Qw7ZfrH2S7451AnEmKKBy
Vo24/6pf4c7hPxTos4lwgdrzmZNGgO9ZcZzOCW8VOqdaHrlzah1mFWbO+N1qARVi
G1iHb9HUMHUsFZwsiYRX8nGGJWYMUakzzUD6Xb39qVW7QNZygKXmKM5V1vJqxEJ8
vKZpFnf0vbQcHd66FzCe/QtCaJPWhY46+oiQlPYNjqkwCR1ZHTV4gp3NyZygC5SR
GBNhAATVXSnPhM0GU022hkiDQD3nstDas8FRbud9OXlF5o1SJTVzpB76CAgZDiIc
4aQou0EViMxx1jetmgFLgqw4Zm+jOp9DY68VF/BrbdW/rrXwTbeCHRttHck9I9sl
K/NfETOfC6V1LkTTsfQaR6tmScxSsY5jOv+0OluAoHKH2xiUxNjH56LXm/IX2V9s
X7gRyqwRSR3n9DzTzV1yUGJrFJAy/ILlfPZBSxt+VsMngcs5IbsGAkjTvbuMIVKi
fzMivO5D22WL2Q/wcdOS6TgMWjm9Ou9EjQdchpGRLima1LvtcVY7IvgHxlko3b55
UV1oV1Rg83JZ4ZwWF5rCWOo1WSbkC8EQMBKnCZhvSfmo49WSJWO/BYpyVZV0eqzS
hwi3trPCKRa7HL0DYkJejjGRD9LNF3iPxPz+W25vgK14fKkKzXamv6SMxFQXwMP0
v4cOEns4ZRGFlrRKp2O9F/ntX7drNb+p929fMriSl+hHtvjFX0cuTuTG/EkRu1UK
cVdsmToDQV4mpkSqpbWsAQmL55COdk0OD/0ftnLiU588VIxKcbSSOfAZrzfCkeAU
HpC4936+OLanqBEo2TpVAIBgr4GmVqruBVQxdlc0m7lvjJ3pX/iLVfVIlg4T52fL
tSfA1wdJWGUnw5R4CuEmYwN6yTdSML2qxQ+/wCpdFUjTk4BYI4JNbzCmSCY6sBe5
lHbuxaQc1GDXM4G9f0v1if5XVzn04gLLIxZ2LoZLS59iz9FQomjmZuLF1HDHRcCa
oxWnCCTeMAeuYL2rFVWhuP1nsuAGuTRhJ7rgmMRaP4NUcsNPBmxpEAllUhcozxZR
esU1LjugaDGPLMPx+Nhw3wAPfXyAri0iU9kDp5PTMDnke0inCMJm29NDBgKxSy1V
bYH+ZvDQjCZvInvO7t9CieLs9dLpnagfhekyMgpfg1poiObmxkjBH+80zpO7ZiZq
lcDxtkb07PookmzohHqsd2hfCX/0v2mgDtaGC6f50q7xJy8LTYfghSn2UKbRE4Vk
XTaLcjLWswKuUBgL/eA69wMRuDaHOLWFUygd7rlGljH9U3ecFq4elirHqPlydYiw
1cJXMoFRzx+ePtZq/p0HHZO1Ff3aDIq7QZNGcFeGkTUQubE59B5bKIyShUHPCJOU
cn7MCqj1fLj2rAVMTG7mtivr2L1cOPaYbyWNpVk2xbbY2nVwwJGjmgP4uISRy3PV
uivCQ2bDatImevX7EqPn2/w9/UlQ0DpKoR+LSZhWh5Fz8RlcvQPAdoHzYNkVTi6i
P0HfiYMIMPSIbARpIENfAmiUemkqJCwZ3wW/6YGXXRKlN39vKsI1XEMYIESRI/Wr
GCSKvlV2jtusztlruaGIdZYDXUovgoiLqEkDPtRsfstQPvoc1L/CEPKiv0D8MRD4
8+FN8VkksXGNZEQUzmKMwybuwxnFjK0JUyObyjpzxLponJq57vqoE3skrhgFz9WZ
s37YA5SyHh92CwQ1B80xD4zFk1u8I2TMhAOjLuuGeF/A7dWk0JBKxVtZVbrlyQwO
/TsUHRluXw8nf8u61N7ZTY+mAX7wKpWlq4cST6Cog+iMHww9eFj2pae4UGr7Me2O
gtJq7ln3gVXDypqdBLFMVIjcvNIkMnR3gKSb8P/f7bAwA7l0L6kBe8sWqhir61o/
z62Rk+MXy9Zqr2nWrfu3CxE4YU57RQ30+vzKhosiqT12DrXkj3ULY8nySiGZsbX6
NCBBSGLxNjTCBLlR1u1ZHo6mUqc+rO2ycKkaxM47sXYkXh37wGXGnD6YKQdGs0V2
fc/UG/IbjlMG4mjvvTDQq/ccDYagys6d8L2+t26xKRmWTVwUO3rfhrxqkdWz5nJV
fzumSY7a8bH/T3jtfXWLfQ==
`protect END_PROTECTED
