`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1sEtB6AverdosaT/BoSFpyCMe0AYd6i0LP+u7XVfaeooLW3wk6+AFFr7Kd/78Lmo
/PEspKoIZWz92bwbuDtGdJ6xyIjaPl27o8w/MG/GX9np0ms5ueJtr1ye9oBJsRVV
ibOc+AJjfCfply+Jpz5Ifs8dQarjS9j2iCt/gC1stmKiHoWemaO0DYuLyILKKMr/
FuOseo7Wr2NTGEWYB0kMwg9w2XfWG3z1gXzaes9sGGMoIxDh4w7ywaATy4UTXA9f
9ZAKD60NY78EQvtRLgso+HY5ucOekrH02Mp/kkqFMFqZfSUd2Z8SSt6hMSWDlDV/
Ck/GQ5bQj3RPzi3I9KQI8bgnjJdNBOno151YGLDkxrsBo+96fAE9ZYs6Gxyogh9j
qTNeH2LWJpihAA0UAG3ITDo7mO92WxWQKD2zmTh+m5c2XsOwYekVlDGJi3QwwAMh
e2t/IhoNvxMJq+Sy3ArCyegvY+yFfcKx/QOwqSOlvPF8vn/UJOPVYFlfG+q58MSk
t9RisOED5zXet6j2TgDpKo5Djc34nG6HAM+p0dXXtzIiDDx/bG8SusEj+Qmgd4et
2AvNAJ3XAIwLvn1/zC8P8EooVAY9R930igUh5blzu4Rd0aA9KY4lSghuAghTxMw8
0c2n0Oa5k9O62I9Do1qBWrMCzhB7wXlf5SNs5StFCgu6nCTCZb35cFeZmWeOQo32
`protect END_PROTECTED
