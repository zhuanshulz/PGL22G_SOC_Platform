`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QlxBYungWkkvN8GEfnd5zW2rLVgPQ0bJzPFJVc85drsIr4yAGvMXOtDafzKto6V0
LA2efakdcSijRwgIW8l1PzKMC0kvkCxfUDTmwcHKjJhJvkgdFdDBlXOMqloe34E1
GlOkCvtd4M2URdhvCI5/2rMKpUdelhu5FsQ6n4nSipf5TuMbnbxPc1R6Vd6zTY5O
tFBVmOvEpVigGGGjyHhFhgM4kw7bo52mD0kDuhE231soGeLjN03jBOAtLWVG4ZIZ
RqYOTb4J3LH27haF0RoZuw==
`protect END_PROTECTED
