`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RWrMqx3yYSoRsisevsCbss0M3XNrQQi+3LQdHkejtiWm3/5uN0f3cRobvoLMU9VV
TTc6UONyVPIFndZwjZ8kbtifpzZhfMIQzmuy9TX+KVQJeFHERj2+uR+BhJ52mHfL
qbMDT+bilNmy7dlux2c2NbxdzpvgV/uCauAZhm4LbKNzj8eKziGDjodCRh1DUESz
his/ToNgvM0nZcGGrxI9PCT3YTw1Z37rNhzJWKy0g+7e0s+k8L6nqVgnUrs0JUYF
WzAr2WBgnVI1gC18RcQ1zU0ICtfzHcfV50T+YjFHGF8X0ilgnCTx6qZhSr27a33R
+q0CuAQVZB8w9LwbWaacuyt8RTUIWyJJ3Zm3ceCBshjkxolcJ4iiJXXhbftcrbhE
HwSf4e+ysnZMECVs680CP6wAFp1eRi4+wu1Ob327qjlBqcBim9xm8NyFEDMLlfho
+KCTOluF4jSiToZDfL0/r+D+JN8TQ6ADsVaoF7b/jbC2zzBAj8Abx1msB1pg8ZAc
L58+8SwaMt5YH/JBB/pUKLYxcWNydTAJTHkYQRsUN1fQo8sRSV7gKGIgH86Ylen6
UXVMpUv+z64R3ykaoBj1YLFPtmFi6/8cpoZmfPco4Ci+yFqohTm4Q6Td92rP3Ycf
3wbwUIXsUFAXFlN7OtSllZLdXK7VLWeRUyMMKiby/v1UZnkEeCRxvsT3nWbwVJnY
GU/mOKAN83HfypxUWIqJXaf1u/PbtXYUgNI2z1/0kiiDPzSmKwoRYoDwXZcPiOwi
FWQ/GKIcrxXrcnhxp0HWqTgWMLEcZRz7gSMdRonrNYRlurc6j+4huuewT5s/uGT4
ECJC/KnDUDiK3gKpTFHvvjm/et65GCb1G53eONHs/E+npHux0uEM0CK4qYlWeDhx
GUuuRk6+fSk03w3fiAUT7A==
`protect END_PROTECTED
