`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51ckxFKQJQDnTf149OoGGFy2LEDBTpCpsDwynBq3FfHqOoyN2ZTI4jdf6qn5WIJj
RwttKUjvtRwvFj7QIvF/Tc7fTZH+5gGlYR81DxjN9EzQkFtYz2njIQw66qvAC7/I
7+gXetCHAzjMn/C7WBbg8X8aRK4SWa4fdTxZKA8WXa6FPtVUVU7698cVsJ6OXooe
uSqIhzOmAdHh60lBAEs1QE54CzvsvnxxD9vzreTcCmAcjchEQho3mwz0mUVbOL4t
/EvABQoyCJ6o8ZK+IPU0iiBXG9Kw4zq5r2uClDZ34/pEbWRfIDLV49LC+axmm6IA
WXIMGnNTERrTb8CvCEjcInx+nqR5dHaigYVzIH0MxU/Wrw/m8pddXvITAI322y3G
gKrFkBPOSP8NPwiZ5LCsQOEdL+1osJpdomZTcT5Q3GgJ1gQkxTJQx/Xeco5klIeg
qWGGMVhWCAJW8a4ewHZyqpw35gSr8vcrtHz/NvKs3xGIaItFOoMXh46H9m7DHXaZ
79ZnsXaOKH8+VuvrrCsTneLF6jz6D0bW5DGXep3sEXijSMMRyeBVe3lK68upOgaF
hCgn2F8EO9VqlQa81oXdCQ==
`protect END_PROTECTED
