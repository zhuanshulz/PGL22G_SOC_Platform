`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZCXkI8M7I5W0hJ+d0VEQq8h5XwmoicF9dJmSgA/4jGyalrjyEDHu1LaCYEvWX41
baAf06SWBXffJ9YtI4LzGQi9SYmbKbwLKGRM64ocv2XeO2etQLE4oyhDXyTWRKd8
b1QjiJW2sQ3SVGSRru4s8PQFpQDKsu0Eibe5s6BSyn6hpcONE5BsBu75er6X8im3
gizkNgDi+W4pxF3BE8K19L+TOjaOLNVhXtbZVokijP/ZR/RlgonchcHh9ECzl0lk
yMJdMd5dqsRr3IFW2ixKWf4vGA7bMClKeChbl+MfS85o3mBFBwSd/veH6OnNrXmT
IIx9+PMnD8c3tlL54TLtEZ2fTc3qSgT9BIEcf3cP01Pg4GmiZN4S1z4vcFY0DvOq
G62Opi4xYkU8b9GFu/W7tBK3cbQCc09d777If6UZFYhSGYJVaJNbz3FT7qe9wpNh
H7dFnwEOwA0BZ5HeAKlMDB8G+0ugr5zY5YB6DLV10tqfJoh8VALxpvfg3OETeg9i
f7/fm/AE/QqeZ8qtH21zPTgRsOce5uMRpYO3KG2ZtMJ8rwbu9kX54ap/YaBGBCYe
3hM/yTGKfcW9MENYfkPgE23lLSSKWfcBUevFl9uKMR3AXAIsqZub9Pu906x0azvX
dl4xQ23YxZeDdEkSRGWY7Z1NDYKROn0qDlJ8RBy4V3mB95+6qouI1PfP6hy0DM+m
objedTOkwXZd2HPFnFjbS+K3ZBDpEJgY4sIO1B1DXcyPkpL8rKHNbzXsTinDlavj
IXZovEiSnAYvSODusLSoyYc8A/fYldHSsOg4VXqD1y8DA9khhnMNyBTX5SeTyVYZ
8j8QOdmu0zkFqMeBIhUutR/0+5cAsX6N+9mgfQWkR2avDKAWNM3x16XBAHs3zEyH
/UydFHP0PgBtAiu8ym2ozk/f65LunXzOXX3ZojerMGH6j8qrXBcVgs2k8Eg64GKC
unZSfAJvyH2MmDAZTdRkcmkAqsLVmFJMEYLYGbYv8ooFS1SjkM3yfJTS0Qx5nVFK
aSqXJVH4fw7zQdyOTsRg8PO44yC7DF/loC3xccDAf7GDSebgDanVfycsx0LYm1an
gRtOlvh7B3zhcDc+KO9TdlBrsblOyC5+5ZDV1j3ZyZnwtxsY2gHfF92BwMQ2PCMH
i4eoN3KrWMUVRsiVtYwIXIjXECv2fCnsYdBbNQOB1Oq9B8vJF8mHTNSluHOQu5/U
kSQIQPVTPYczAMpchf/NCfgLQSz+e+kJUxrYDcsZBxKyNuCnTKf4yc0GnMH1wUF0
xnZgzis/+K66b/rLAE42rQGU7rIhmXwrCE7yRU0a0aDjyZnDzJetCm5fYMw1BDM6
SlZzY++CwG2sTacLUir6S3pGp/kK016qP3X5y9QN4Kyr+8DCcMubScgwhhaHaS1g
EGUZmFYflZpqRzbqhZMfYkFON04eKGBPjv2VcRD8MFifOCmmJ7uBLKpvSx7gTTq8
UpM//Q+EHP6a+I4yBuZ332qkI4oSW164fra79dPC+fFA9A2F0HsPL7Msd1NFyZZF
HL7kTvc/1AP5l0Ag87kMgZadFnEOco93hxY0urcbuiWpF25knsiQVuHlGECQEuDu
pgPYHwRJiknPFRMgoRZ62ZtVIGv1MCb/t6vbljnfToK9y43W4UsYwa1tAlfmJU+C
cAtFAP11T97QLeAlFYS4rdoXiVT1AGXKZzXhvwWEFtmHZT2Q1cwnRiIjmgTDCHoV
qaoUKZgVQQF/0HINPthGp0vB6esELPFQQp91G+jWTGuU4QlD4KVo3h2sW8L64cvB
661esGRVc3bEBRTCeM2GZGDH4ILOOcGiJmGSXktBF3c5LmtCLaIytlzlh6Xssxjj
wXMw8MZ35nQNJX7f9SX/i4Fq9YnZVCc6WWe+7C1sWeqyhh46r9EQvsjCtOr821cO
vyjpA2L0HYpVvx/MVbT197JNLue/qfJFYZihrdAXYzi8cFp1o9fItFxg7zKsdhb4
yXoReOu9whG8cZWTciXcDYpNdg7BW/cs5s5HB8n7N9SD9Yg5+MVICM2/XdYyI0Ui
Rw1p2qqAjlkQ3dqfwJkAQw2gllsQggGjvsdcEu6+FvQPpX2m4IiSC6tPVpErO6eA
WdWvc1YxONG4sKI5eHUeV919dRLTC/UvdIBy/aSpAKRAPWeRmOtIdVCkB20l/uj8
5oqU7UiMQ8WfAZJ77zQXNXcjBruEoqPnaLG+iFJYD+s8doA0mASjK7q4v6udqKh1
MqML/YEVcD0dFsybOPmwQVde1fpE/pMnv2ZAZoYPd5OhZs2tjdnT2JcLh3hui23U
KrsNbiTtuz+in5VLMJyb4NNrN9mpaXBsjSLJzakzUGGJQ53U38UXe6gYby0DhhAp
8AnvOgVG0YGV1EqNbfo0r0I1cfbBtJbj/iTpqhA76yCLDt367dsmRy8dFyNa8zeB
swu3TfCzyl5oUH8p8+rYb1LvkXuypBSr7Qlmx8hSGDaE/fPMZx8SkbSBUwLdb8n9
POpadjeUzidOgPm81xN8VjxyG+YnJBiRLPsZKsv9Uilf7T/fL7x3awI2SW8NQxGl
Vf5o2h+W9ZBX0XwekOYioB8S8M2x08/3ehAhPHTezFtDAMG7yWk693p9SrhlffLC
EJCWmb4j7Y1FOwegDVDJKNBOvRpYYC9OsPOollRQLC4+liwKiqyHc3Na0hBPwvqj
sCde9YwW8vtPbP/v+9qXoyVp0c4NVQeq7P2JzZZPDjQOwN2h81LJQNFXt5mbddN7
pe0icZMnkA+e64EyBCQh6lWel8sQBk8EFvSuBcfyYYzEOsZw9/iNvCClgll98MDD
DvaKcZ7STUI58MD3n8fG8ZSbAHcQyuMD4/jkESfBO0lSBBmj/FgiaqzfEIx3IxyB
YKNk5V6UP0jHd9Z3flU9zBo3yXRZv4EzZZy/+AhNpJSfRcUwTeoOini5s8tU+2E8
dBSE5r11VYaleQcfdndp1aJieX2BuaVKX2Op1HX8T1j3afsyrEdzIK6Ld2WKL56h
+bIvWodKlA4snSdy2AkJKA+6xa3TGZt/NStkDc6ae2tO8zctuhdkubmayD2LCTuK
/ctLYpTwSVfivcyoFp72woRoZQl5r/HUfhR2PDNMI8K+tWRNeWUIiil+GGMgQFxa
Sw5bl2EHcaK2bkndBMlwR9mcOj/cdDnjyrISehFONIwbhtSnKub8nGJjkiCKXY6S
jQTyYAIeZyVk8ANsCOQpGxEBZqJRZdamJ/RnpyPrO3MJR5+Bvxgcg4osfFd52XNi
ZJiKvTkXTuSwpVUbl35r1O9MIHKe3iWxmlc9cj+X4yyNy97WYR9lwNBF/RNvkopq
EZ9pgNCHxMSGvrldw5o9cg8/CMk2JqUnoe1YEzldK23pIWAy/iUEBVXF4t2brMBz
0SYhkUaU9Bkg5+onncYCrcZZ36HKe7ZO0bD7JI45sVyQ0Gm783kub9QV3ndbKamO
uLixGyd+Oa6+lhtENDgHj8q5LPqUDNqpUh4hZS6bzhOl8w6RM13C7uZaTBmEKQvA
RapuCdfqb8a4Uysr51abKmE7a+IT4ske6la9hzu3Y9FkMPu7bk07shaztV5HkBH2
NsHkC94MM/kALpf7Ta0R8WOOyj9eERFBemj+BgMjaxnmPT9SqEiNyMMJ0thF7Z/N
r4NFJrkTLKPq++mlCEytBH6F86Lxd7+K07DMrhkvE0Ms4NL2cyDvLRZFWyVMLrW1
NNrbBX7I/GIApDq1LJCadBUMa3RNnq5hbDYaIgJaF88U5/RUdZpUEzdjXICNzN7s
seYksO2IH0OQCAnWYKVE8FZAjzehZ02YHhuS4sMELQUV+20vyVQlAax+1AAOv1c0
0omabl1s+66bpvPYhJ8f0XM9gALkmgunmXIRMzpG1OY0DVRjbq/kktX1oyi4DFWK
ik45vJrFCRuxtC7D3qTvf4nBwP51lk9wlPplNYhq9V6W8K5Yz4aEn6dhBiZS//OB
I6fs0DuvcNMdf9Y0qq/QrPlfP2cNsuqAa5k1kdFVSX3PNkBPT2bhlUslQKzynRmU
lGhlz6aDx5GOvu9x32clZbQTnq0F/wup2ggM/az+AumFv84+TUFmbpcpfnn6QrXr
q2w2UX5JOg2nAQl58Oce26aX0GQj00aEyhHd54VbR0DvNr5iQBUWaHLhJJWNz2uJ
DJjAGejwDPReKQDwIuYYQJmtb8JYjSJWem9cH4vcmVBTrOhuV9OJI+VI198f1Pyn
gJV0m3bh2NXPBjrxNLkrp1yhXP1S0/NtZIIEAuLRkgAfLwglEn7EI20nKmJuO/6e
6VjoBh55OIT/gndJfUZnJO7yIxy7SyvrM4rfzcGUVpVQVDbK8QBJW9ZpeRPtXE95
Qh+4G3xI0+ubyQ0Z7YaKE2QikSkcDFebSNeFjabMVsW5RugtuCWVCppXflxANTTr
YKRKoqyccTWnZJLI5zUz5w9wgNqIdK6C0TaE398vmMEwfjr55IMVn6CUkQlXeCex
xfOcAd0Wc86OpTmB4R3lp3CGCLD3LK6Lhn52zPIQKiaB3UTMJbxMyYCPJzrqbHHp
h3c2RcFUgn277poWQ8vY6s200zHVZlNC/7qpwsCsVs6Ll/3Eb6vfFBJx9EJgXvwd
/rwuz5yWjKRtTPIhYnJe/7c2FQqtiL8YxTY3+NTYL+PvOxAtNh5wWfwWG+oRFfYp
HoINxo+r3JqhLcxL8ho6OWVBppnVwnzLcc1S5UH8BGSfMDlKjWIj7vtRxRCJh101
3py8xyq6xyFZnFx35v22TwDHY2BuBIld2ErJPwVevkA3wQCWUkTUyiNBTxr520Xi
UHSMgLOjja3S9MfHTIM3D92EGOO7LA9JfH118psbeJD45l25hRGYsGshUNxjXBB9
l0que6yCF1qRm4ZkNCo5ObACipIXIWThzm596HV7nT4ev0l9xLKMs6xRso+cy8LP
dcndSH204PM3hlY7SCboWf8PC7xH55+RSJKmrKgyI4ymiz3I6tNm0RQ0ja08Wv5Z
AuTjWFtRE8ZttrjF3FsM0Ytyvh6mKzyZU7nrFiffUC9TxgtlKwHGQ3zwt0sJpcin
rWWxwTpbrfCLA9EkbASkkIC28+NhhFolWBMffMk5tlOl2pFPve98fdZgX31013xE
dzQL1u4dMDJnlGcBEYWVon1UvOzJbn/RIXFno3y0EIoOV6ezY7sy9PWw0oYDy1HQ
HxuX0mv/EXxIYP9bVkj6xADNB3MK1fOXQXWTbC0yv+w5bxfSgpAs8kUJjC7Z3mf5
6o2r94ND/vIkTm5B3+tInBjwz4tzsnYK1ue1wKyXucv6/zKVnI2HZxTmW9eBPgL/
X3TBw3ti15TA7CjiRYrAVkNjhsHCrmQ8DvMd3NUuQwR/XZ8JvEdajjcw6X3h+RUm
iTZpm/ANxKDOldXbFDWFWizGvAXDS/qpd2Na7zLpzJXY6nty1fAbshVm8SbaTvsT
SPoy7zupslof7xXQ3oG3oPdCRPXYuE87MOxjlFL2OwoVu/6HaAMxL2Q0RYPy4UeB
aQv2HNelIYTyqadk1Za7IBk2twA1llzGNuf6TluH7W/IVedYYkL6OAU7wA1KgRGX
pOFzJpOG9FfWZh+b5cwzXi9Pcz+kMpqk6H+vlHuUsMGQNDVAvoR+V6ASWY7uNlZe
UJjj1XWKq5JjsIbusjYkv61yBykIk0XqAElMjeIYcxA5kqjp60U8epsu6raVSmiC
fyvP9AwXZEG/7p0y+aE+Omv2MW42bP7TW5+u9k3WmyqiIpDehJvWnMd3TBL3CLiv
iktG+sWRKR7+CV3kT+MUc32rWaQXQoYeOw7Y+7MxEJGAPUIaXnGJOUuE3qctqZZM
DNxrTC5HGwSo5fRadm7t6oT65lmBxsEGuAwmVdUPtq52uBKXt5H3nmp8Lk7qVbGg
6N85JBER/Ahc6L2wFNMTXRmplTl5Qj0u0bBiqZVAvvVX6kXskr3LJkFTBQGj23l3
g6VUcIVD+ST0MlyibEIdv6zhi0sBCxQk433a0gdIacqWKqqYgvVlyHFncWfgtpfI
9jpMelnIOFwM3gGk6/isBOwyYTyG3P9dMasdbtnoLq3N9nZUzfxLl9vcleP+bDDK
hs/GTEZtSPT9bpFdPOyGdpVwuMQL2tIvDUma9gmVjnciu/r1SrE8DAmegT063dIr
sZCxR3K5cV+xC92yv6l5d9ZSCfSHN5Mu/IjV0Sn4odvV7iwd1bglvYoF/HKXsvCt
JlukRglZHbcmRD8Vap44EIs+YklxnLj86F6uosiDd6RkfRWxiJoEqiBh5Noz3oEn
oIYrfby6T7mZIwaNBUEQ8XWPoT7V6qj/Q0DNJX8VBOZJ77D2DPhv+V1hxnlyi5Tc
l8p29v8f/s4DJqlyE+P+2oTUBfIQ00NM47YEsQR51ba5ZNESCsON4FC/OztUaI/T
lM4Nkp3AWLwAzbfoLpfqLKH6Ds01E8i54o4tEOYtoC+k+LraMIpf620OzhF486K6
eJkoWGmFFA1M3nd7+fm6qnzvIn0tGORwKaBKVrtWX2WEn3z+XtBI1vrUPhCj0mhq
OXsXIBo3BBixajhX49xL9MeN9WJqNdCk2EMiNJ24Zm8ZVYfJQHF/Uy4NmO2Dq3+M
I34MdzESbcjuMQdb+mY65K+2wGX1d40QUaOSBeMI0vcCsAWb6J3BsicMNZvdoFXI
v8KRaFlvJS1HvTrhtPfEtbLr+tjVs4EGlRgdxzCXT/aHCxkEJLt9PbNbgaJ7miQ8
Jxb5ThjA6Tld+N5G5JZrNYhZuQ8rJkSFsny3xfQiqjgLWR2RKRIhfnupPNDqAqye
r+heNoAR3Wgbp0brSRpmhfRG3HxrCHoe6EHTKs8CGypiIAncMWTvz3fOx/l2qn5W
2pRn3HGhlmTM98tVPHeKABeqg1SI/MLOUpnzskSogNGKFXwr7PdWietfUeEPGQ7n
9tdLsyw7Zvk6b5/tjzWQzF7I5n7LyXYt1cg7fgedibATNBAGTTxoXry44VdaEs6Y
MLqdFgAbMibrSpFn3URb58OX8wn18Ltvps6oxDxxbymhiopEuPC9xfXuuGwu/7S/
wNbVS01UIZ4DJnWa62x0LHftKasylngyz1jDweYy+t4Ke7eciv3pFFgDaC89wDYY
Jb5y4uWc0zr75fUNgt915fFbjvKkvsaKxhmijW8r+q1TvKZej+JrIqQZh4IA5FyT
mKnann+KUgmO8HyDtpPEwHMmFoKgjdas2ZpbJEYKSJYdFfkf7qfJwwORiNdGb8ST
2JHfBLYq7wIaiTfOddR6ig6/rSKJ5/8olzg5Ywz2WuW+Fw+yWtXJ16ovYowZOVnM
KLeZQlK+DMiaJ4bRYkIroMk4iBNhYeapNxQduBh2pucGhpF8aJmjhVJIavi+AR8n
RbRYcdXu0LJF19QsQ5PoGUUa2CCD8VST/KLvTAkXRmuzbfhvCCBu0OmsZsO5Ccrj
24UnR4o7nOVKq9TGx8j2KIGlDXaIZuLT9Ksez9j9bob4WGNTxB+Xj5IflMU049OZ
yHAVsxcCZyH2yUkuaPL4fJe0IHBbkYDH78WW7YwPCknXww3ye7LjHeq5jjW1djlg
UpHcWOXL/+mts2sN8Jsl5zwqPtoymANrEVjVJym9/WwicP/nBL2qNcorPc5HumSw
Zh0cHEUiNJ2oh2PKgAPkhMDjhA/LNCYMXGpt29yu9qp7nui8iPiT4KY/nkQPS7lR
ftEDde7I+yFDa0cNejjIDNO7S9lg9CpQhWhIR7Lx4my+W8t1qq6k+6KOMe7GzGXS
vGeQJVp2gowRTex3KmOGFJCQ7IxCN/GhE+iO0ZcNzY3fGw+0ZH+3Sw7wUcG7LQSe
ylwqsYT7A0KJeujD0ltlHl3763GeclgHK2fpPe+jUnItqW3h7rGkddGRf8r7uAO5
1opYSCdqNTzi5ePL6XvzxOToJaRTTyNqBMcHPrpxI4WKT6tTPm2f3bhZDn/TXRa5
hRCwUsZI+WWzxZk04VrTNjqPvbi+moM+ia/pfut32RN08Qf5XSWQ3ldKo1+Yokn4
BkmgzC+1uJwqKY7+dGET5QQY/XwsP9pG2tqohnPWFOHXux9lL15Crr99RwYr8j5o
UTNZX6vayzfBC0oByz16eDoKkxWkWY+hWMnBO6/GWVE8u1geLZbLfIE6egvXStu5
Qgg9DK8E0gOGDFnjcgceqsC9mklBmUfnWYyf6DDX2HAlqbWinuENfDxNj/QJKIB6
kWxmvNonspSaQ6phzsMJoSSI2PytGhHNGuTgNIo1R11W/wUQrdcyoVXqi3ZcocPu
iTbAFCnw+o9Rhc0KcUp1DniBpUlTdsSCrTcMdD1gfbYqW+Op2ims+Qvs0JtmoPdJ
pyAiLAGdZk8pZToBjhU0OcC5y0zmM6xcP0BIPZPZXZL+PxNa2Xh2dCbhwbrjOiH+
K1/pWtMDQGjBFK+w5LDzfUCwXt9AEbwZK8MyPbhUx1wLKQEVjyADGga9+wYurix9
bRSxiLblwf79knj+fw+Dhwn0u6Twy+JOTbjRvPRV04Js3xlVRjhqBd4py5kAXx/T
GLOqSPlVa+vcOl7QWMQyGI/FZkPB2dfzqriSwRxYh3t1udrj2A86w+2MsVLkqTPw
5U2Y0oEWDyfVA911Dfq92SbS2QraoEXcat11EcN9QgAnEmOWpoDfdlW195sDs9n1
yj2/1jF8T/Ie5kN6mQIz+IYwl7HrREgipymvqnjmFuEdKAom85hqujfeSb2AjCjl
4deZia1BLvMHFGp6F2oY+hVkmtJYKeMn1qU2qcYDohZDV9dFrf12w7Um0/SphScU
MrBcaTuiQUjMqQQKXvagA+chLXvf1La08JKU+kkIcCExpkvzD/reBFX2inp3Q2BS
UbDnlJCkZay/UZcauztMW96YWsytsTD6zojjo0G1hnuSHQEcJqJEr+4gQnrscVZ1
sJ0T16/79D5tPtta7xT6HHAT7ZlkTirE34iOauSu9n8Nn+7t2Yav5/lqMzCye5VO
xoLSYp5AhzmraFkQV2+CGKHTUgAWddlmI5Dwl7IhFR2faNzWsC72WRLwoLTiVQmH
fGvsZRhCtJhKNmlKJiA6plUy0vdw1fkCvUqQlNeExY36S3REc6cdueZ82kYrrWaq
1SSlmDVxSs7gWrsYzeWU/bQIRTAmmHSRu9RuyetA8sgP1u4q6okJberf+3iHGrOs
aC7ufnF4qwm7ClGLsiqPlj2aB2hwVDzBencgA/88bmC+GfTZQ/k8Kh993ZKC17rl
FRiTWSLLMfPM/a3b6V6yUxwq/sGcJbrkylPasEEWuDxr290swXUgu1CL+YThuiDo
j2tyPz+qB+s43j2awsnff+PkgeyaokBLjpZlG3MGMVOIOEEO0iGQ2/pKnl9FSHWw
CmAEwyU8mpcoEj+gqg6C5W1ffhWsFxWQ8Na8/nf9rSK83o3rjjzPvjxseFuNw0Cs
cXMajXzYHNN1VSWoemnXyQlg8cLKMwnpaakvQmjSNHmMHq+i+dopw8Tkh7bA4iLx
kYeS/yHdqdsVUV6JvB/uFAVjUUtxAsbLlXvDNG5bJIr3Qe6j8DBa4FmwLhTuPByn
8LRNSYYJ96ok7UMyQsIbm5Aah3DqZQ3WGtyXUFL4HnJcN9RGBPu/6FsPebQIC5Qq
JFZYs+fVvUHymkqbZz5tSZ61OaqeJ8NQOURdorTEP3barDZidGcA4agj7eZMRKWU
Xj8aAHApTp221fijlvYwxI4uVK37VbwVOTKkuiXmPcPxoVmkMfCPLYu5pQVwi5vT
+uIMIp22e68DadDvJIVJ2FS/ySBc+dU1ICLR8LpwJZWIlr/9WoDg68MO55rLef6D
pp8GSKOduPuF/xc0NbFoXAmMhKf95XIudPjEvVRdQjMUUnDkMGM8kyT+orp9L5yB
SWRHDyGWJAfoTYYy5XwgOFZ7HNTbMlzAg500cV/nPTc9NaF+M3RQoVSOcyOot1zZ
LkMoK/ecvSWfDAlC7vx6VebhpzTR/w/1AFUuVkt2lXMABi65cMXAc+QI7kaq+dYZ
HnZpelsM4rKBzRzlklFJbi+5eftPsu1nCmMxeKHf++ZBKtMYYjzGFEzE5iXT2vm5
G3NEGvxaM2ioVuUwJ7NMDCPe/OcDeMlzd0MTp22htrkoVVqc/Tiz1KHdzktahggz
23C9sKdYhLNwmIDr4CJNQrkTIM8Mey28qJH8AeikycHC84Hv3h0CdD4omCsVnG3p
uEOUJ1DbAkSouM1ZJ/zIjlsaOFIa7SZb4dTrvQNIIVQLFzb26YOMqwKBJWu7w58Y
GwDJUR1M1TVIUtmdkCnUS/vhf1Xldn+e8Kl2/O4daRxUEhyShaSvp0PLA01CvzrL
KG8UPOGsvuUgFg1/uO+Amhc5oVfJO0/SxC0IL9/2yMuIdEPP3Ssmv8Xi2sn+lsOn
7/CHztI039FP0VtSQaDl5LctLhybOHs9lgSff6qsvqSj80byc5wz0Pn2RRESnk1l
snhhKeT69Gh8PSPBTjUAA+XtZGTPs6MhPXUvQi/UsT3Fikk+YBwD5SGhmniyLlSk
vuCyMmyc7bEBmlG06KTtC67LVVZNGoijmlYOMzpysEw9phOFtRlNENHrlGXqNkS1
t/3nnIxbw2UzeGPZQLjOe7N5xqq/uhgEiEdOoev51ztbjT+WCORWpn3LHqePwaAd
DSZ6kSQLusmVRLJl3niig8mU1ffqB/40JdIMehQ4xOSN6RrpvJxeZdKj1KM+WkQD
HmvY2g1TYV7ixjmXbsvEA5PBNlLQ3PD/capau3vjZRgsGZocbIzsuf9YvdS4etHh
v4brFqU+mI4JxW3m0o2axlR/8bu4jL6uTNG/PcZ/A2I9uAwxn2F4U4sqbeXWXWrj
DV/0pdWuDu/BSxTtcZ+Xn3osToNPoS8Akgw/i1Nizi4EYAa4TX6sRBfYaIUGxD9Q
xXX58cwz2+nYqQcdAwk6W1NtWnaI51j+q1DnhpT5IqNeCdmZDtZ3nSRlTrs072rs
9JMfocx/xi23HlcJnQxCMPnQQM/fBm/Q4JnKQWsh0dzN5oL9R70ldxNu5Ht4CBs5
M6PhBSw+7meQ8Q9rumC/EfSuNw7SsS2OeOcWZ0Ab0kwpBam82zZg6bmJ1tHRZGVS
ngq88wPXjyDY6uZcppoQhK8EOyujEJBUvpTsEzDNUxKvTvkmyVWYMj0gzlQQ8KsP
FuGnfVJflUo4DB5v7IRD1yUq0y9nIsv5OSq+bn9xoSjryrnVnL73o2t0KYXUlLcR
QApK8G1CnafMHGuE8eVxF5k0z5BnlvlCIHosoQ/y2GAb08mdYSLmi7i27jWrQ8IH
RZrspFyaYUrRg7OclYeRHBUXp+i+bRHKg/bIk9AZd02ffP9K/u2KE4w8heDCfWBu
y17eKMjXvjm+kxxiN2bqFb41eCYJrEibnoekBCCpGdUvTUKOWldQfvDELuiBcxeF
a0pyFtRcCn8k7K9xUTqRer5Gd3qqfo7599soGi9oXJFVi0svxyyqc5zT4dh49jwX
V6CZDGAhFlSrG6aJ9rBIQXllB5m+AjdwCxh8Ohhs0nSe55MEgY/vGf0YoPYU2zmb
leCAIosgomeUW04bp+eOB50VznUOScE6evuyQk/55uvb/QNEQItE18z/U9jfQ5qo
XqyKzCo4ZySbNUsi0mma9wdAvfAhDRxdhQRPFGNthOa32BVybaHYXbGh3vFjm7eS
LZyVCA4Nayo7ygzRGwx/5n7h53aamt1HE3B8/wy+6DyHjmvC9ob5mqgy/olgWqnR
TSJUFpTcKy1L9TT4/yC0PZj5nrhvCSSjbj9PNQHIeZxhpsKhPA8j/zkC5dajH77L
9c5KCgwAQMp7slp389RfDMCIviYo5qsPbKZK5AvxvPsVm5x+ZY8I7nmIPqPyxR2H
RC8Jas0nvEs81OU0YHNI1uEyk7zoOC0lfweXJIFxLmJsYEzGBIpeONyXQ768MNha
TOFx4ppPFrJf4b8rVtlVk4jOLnkv6+4mc7N30czFc0Dt92j/c/lKJjw6zeB+Txcr
Bmf4Eun1Ekld+UXqB6yEAnWBbCghJczRSJ+gN2KBaZPrLNjhTwu2yV7iiCRohFcs
YdSQagUlQcxCVYrfXz3JC3h058TrmRJYHC2H33VDyyJsZmKBAvcP4zMbQXvRbuwH
BbN5Lpi6KzJMwToJRb6mS0mUEzniyIpbkXmpb3KaGqDgR5Rfad/5gjZjqp2rx9Gr
8PzEvrcLOra5/JPiCwCcNUWudiQ1AWk+8nsluv+piPjrkW8CxRjK/gp+o6ycC9dd
yD8brXkfb74UYNy6+f2jC9EQ96R5JhrdokQeoPY/E5Rq7LS0vUl1EzVtK7EYDra1
hdsTjHYb1HIoOQ/UVGcjJ+VbkET9wKjyFbFQ9U2onn09FHlomG6zRTHg7ljdFSPD
qTG1XZ29hLFIQtTGnPbOMTiLGYdhw0OVU0lr89nAETvUCI41g81gXfbXy7s/1Y0u
tRe1Kyy2UxlHR6E/1Bqent9HWXpx3PwQXjfdfc0NwJ/+LE0ypDPKYPPzJrqhcbeT
rmR1dVy8eUao+x+rnDfAvStYo6Q5obLhOKkOUtuHWX08UoRhJ83jDcELO/P/k1PP
6xJaxSDMIgk98cotdL4/zw87S8oHOe+uCBNs8jv5dDSY6zrYSztw+S0e91ZQE3/M
teTDAm6nN84WX4ywaDCfkhnf8WEuuuSTVCWnCZOVt23EyxmmyF/XAKceCWc3lR91
iZ0V9SsTlCJJCC7L8Z6dSDDsmQeDrVfZXLTYu9tsFTLLTnoVnABCRUliLChoj27G
S6WcgN8qWvb9XcbRMqr9tQ8GgBra4AtnNIxkx1bH53Z17HMMTJMCeVsoiWOcLmUV
Y9ueWeoCmMl0wT96dgjZY050TBrInt0dOdoGmDi/uXCUM8AdapiM5vSZgZf5rJ44
W0fQhL09mFDShYxukoPT+8ih4NNNBGlJf3PkzK37R4UT9q+ATbn7/OClbMQTVNLu
/D1tWbjFSaXBZ7yx9vzyTXjL6IiStPZ45Th99XOStLtbHIRu9ZfyvyuTRXzorvcy
oGZ2MoakgRWa1HSO2vK2ZdopLaREvaKf7a+7N+NP2zikLnCo2vsAulLVDB0lN2gs
cqcSsXsNp3aIl7/lMMdrbMVfj9m9frWAYkD0De3JOLN8StlZZw5qpixoeQurGIo6
0vPr+bA3RdIDW7QZB6oSl/Mq111x34R75Vkd0VA43Rw2v/ZivvXGDp8uQMyoTW0A
dWA4iHfA9+7gNisFau5RTmK44UuTbE1pj8JEl6EYgfRl7j6so4SXVVCmBoiPXaSL
3QjaPJXKTUvzGZr05gL388aP+5nBrE2AvAQkinS0G5BVO1LeWoJRHaXLiOlMoDY0
LM43v+ASOFY5Hfcf61rH1y4anOW97qr+409AWme6vZNkLWWM/w6cpN82Ow7qUwNt
TnW1xyYBIBcFMS1GT9bbU4uQxhtDcSsl2rCbKyXxjRGhStcsg/i4vAGjjFHIOp/6
OkXC+DLB42QUMPkCkb+5BU7LnVujcpr/Mbs/uraEvVIWoCSl1HmzRyyh2+8FFIOj
qB/j22C00YyYy4tQ0wXtPlycCeGE3doAMoN5pxrzS78+Fo5xeybv27jdeJ+SRGgw
C+/TA6jLyu0JVaVUeQWZ2bHt3ERT1pZDcD+8ZNRRS4dx2IhRX1YcinaIB11Ixnuv
/q2/V2rxTGNzYRszIKI14Ks6HPGVfKWofjVElLrfS6Ae3sw3mYsFOOfv74PH9Gcu
YENpXakU5Bdak05NwHc/lmRgnb9VvNaXoFBrliMlhWNcHr4oWS8V/NlmdXOznoFq
V16W+6LuHLCUAxb8NpFPfg7fUS23HS+grmwoX8aosUqthbqewrDKKtgCS1u4Xj7y
gyykWf5GGn56DNlBkhT+yuL4FC06DULUjCi5V5pN9njXRLgVHLYTFrWbRYLFKFse
2Zfc4iYUevW8GWXDtONd8OSnwB6KSCNvlHKh35tNm46ClhhQDi5yIgReniPA3jQr
pgHKEz9JLPxyIZs1SP1OFz0Jc+cDv+ke95xJw0XoIuGkMHJ64p1KCGE9JPl21l6G
C6nhFDJdtmfyStqPneEOQvwVCwWBDwWHus9XcEKTaNyAEbnWFix0h7pOaCoDIsXe
wxZPRdm9Uku++HquMaV/RT3AILlbytxYQbSil9M1A1t3fyAJYojunxWzGmLggGEl
p3k+1e+PWuqP88ChxzNo9wMB/SGRytmidFs/X3ShEShUVYkc0Va94WtsA/XmuGZO
8yUBuH7ElUPZIIdBRKU6h9dCt95AmXgOESIgMoDAUBBK0yb/F7Ow9TjcPS1LeGke
59nqIy9QMuf8bXFtPVXQYCot29/6c+uQro2BIgnxm5lykjO9rw5AZzh+KmOdhT7H
/4FLnOcbDyAvHjQkuutvZJMVXK/pQWJ49m3ZUNp4JR6/b59ubL7wS1owkk2r17+5
XEBvSfGRj7rEXc9xkbauPlc7G8zHR0kFjnM6uywsuRZG7lW40DXwB08QYAj2p2Wy
dwhsn9L9MId2bhY7Q4Z48U8kai2QC66o9jd/Db59HqY+jgmOmOT3XCHd3x/sp9t1
bkM7s/252R4wPNp0ZZxuENpQarCBsh6/Vl53PSsU0GKmWXbH7gr2dVjtB70FowDc
np4+zQxRsk1oIwDPtcushHf65M/sPRcMpUOwznIgVoyx0d4PXmklIBJw0PzPIfLU
C6Nnmtfp63NxCAZ/fZ95tQtL1fdVMdm0tL6Prk3RWinjn3Z8g21xoQuWx0QQq97V
144KFDLY/UGCt21Cq0quIqcA8xQXSmqx1vFyGFuiHmw4YrHd3lOws8phRoVUG9wh
ce6ZD0uLh5XnfLX4GMnBX4+jf5z+2zBawg1K8+rWjoOlriqpP5F4zMzuLAyhbWPa
ePOc63WuOilqW+4Kx97T+W1xRNPu1c1xPh1WeTRKPgpVuILEYhjGYrsBPgjPice6
O4Vp+Uv5scxZnST27HKvl+byewE6sU38T4pELliwVbFfqoySPTBqVdKpDUs4fBi9
1e10GrbqDwQDlGPRhtt/PGmEh0MEefA5hnnsCcybr1g5CW0K/ZAoaeOZMlzU0+75
fWx69/kdUKG68qS2PKiDDJyYx5nWHAx8x4tywpjuguxSUVw/lCnDB1pWnFl8wFaH
nT3h5vBKQYdB3w8pH1bMKh80WJ9F1aH6++KqDe7jmD+zjcOBtm7n5VfsFWKde0p5
VzPTsv9sT1nAk2rDzgYiQk58gzv37ApxbfEoHpbl+YJnSX6wlkyYxEXahZ3l0X2q
edGjrLoh3qp31mXEmAQjnb27LHBjBK01auiVAKpyLuL0gnFh5QjDfB2O57b0Td0L
EzgnId7XI4qgjFaC45xaHtg7A/9+UsRTHm87r9dUNbolM+u7GPuE3CqtqJDwMnv0
PZW3KPICZ7NWpUoEB+08k5czZnfljmn2EiYvniFVqp+RD9om4TbLvcy41THFvYqu
TuNgbg9i7vq+xTfniX+FMIfJVi2jN8wobtAtWdzR7ouWx+G8im1mMlB8BFpQJGOj
puLiSdb163jyY623DsGUrWhg3ZaFz54XoqDTTMCxEqx0OQXBzatXV47Eox+aSipN
oO3l/YZeM+1vpAkPU82o4WHyZWzKEwspDmXsgUw/y39bht4sUlIryznjkqmtDdyA
Y+/Tf/jkNbNW+ivnMYMEsN7mMuWKdwhabdTEy/qlyRPKRRzedt0DmQnxrpMyUuU6
BILqTlER95ZcuBiY3spPorpBWLczqS+d32fQClzW2UaiaCD7VFARi5fINc9eJ+/t
Vy4gjz6gIAF9j0r5Mbhsi/NOnq+k73/fhuo6YS8uWLOyJGNA0Bdp4jyVpR06pfQd
yat7fjr523eGj8f0pK24NKweOFvmvXzbfqOg7XD5hatx84nstWCiCpM3xeFSZ9XO
DfmaRjZJU/YTp2Zrw9aCyC6cyrUCKHHNjbXlwHdlOMqOWtqzIKSGsl1g/M+xCR/I
dAN3H+evD37NJBMRMhZ6JUd5WAkJp2Ci4j2KdF0decTsfF8xdqLmiXn4UQA4twtk
JExl9eqhSR7uI5KJ64dbINtpTOB0GC/QHw2tRQtUnvZCX26dxxnud9qmG9lf+c0r
7U/44nC0RFKl+1/a7GeE8/pGuYMbhbaBR0A9n8CrFseqyniXd2+tpH0z57vK/f62
VPAK1UpmLLMcG/dhxI8xH4iamkFJOCX+prqqNitunIGEKyzaAUyNMmEQH2OFqRgh
hX7rGL/tZ8MPgaAFdwqJdahOrhCWRGIFEV4Ggebpl8JQ1Ahmt/mlmRdmd36Sb9v/
gnpGwj00HNSzbwsxAJ7xAP/UEIXNIyTqPLtzWGFAxMFd0HnFhXbOOrTrp8FfIuBx
ORWStkEPBYaI5J1Vnp7PJHk+D8nMDQrcjSaLg05f4SzH+CF7Z8rVmPDG6q6exLEC
lXV/X6cMj2ChfKZC79Yl52r0gACzOZylvFetk4XLGgbDWaXJszg49rXh/Bscp5dn
TKjz91y9c//NYvsWKbPO0qZAP8ldILIs3TCbi/BMoQwlvBJfejKUa/wdsCORXpbB
lv5eZuJy3QEVNqMkyKnX2Keylpe3TDoLSWKWm28/E2Aax0LlfQcXle9YRLkpUODZ
bplwQUYzH9z/eZ2JnnsmzcdYta/RT4uu1Qik/jWBjXLzWrDPka+a7hwv84hI3XxJ
h4jegBHJ25+egUOl6YambItLQwzOOWFXkX14yeOSmv6XFbfPidww8GjKAOD4mWhJ
wagz5GBH7c8pZdNgXjFXnAzctvDUkujljf/cyvMlaypWlt9aFl5AOv7Sdk8NZnaf
Gl4NI6MBmFaL+4cPI7WYKw==
`protect END_PROTECTED
