`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M2pwxrGRm/JE9kD+sILISIW+IQndk8J9Enlnmso/8kPwnUv3BJSyxOXZFXL4qduo
K2f4NNSeFD2LbPLeNUB1f+QPqE/4mdoC7yCkrQQiyca35Le9EVcQ8nveEosHyhnA
yEa0DAfF8qHkYbmtyfGNl5Rh3JsrdqXQFVdjNkM5Pod7RvFIZIAx/pYkhHX0VJsk
NI8xK+F2LugiuUKowQx2wKEYuwN1kufUMs6MqQFu+j76wom4ujogL03U4IK5KIn8
wAVUNaqHz/iFjYaOI5KT8ipMD9iEBSUna1NFFkzrHIrCGdBztJ8fiorEWGUIC/Vg
Omerznx88zfGxD5RLYLM8/wevZaHPJ+LXPxlXh3bB+d99Yhy1x5RvDjDFojILkho
JTM8DP6a06Lu3VneuoNCf/BhLVUIGSTBnonWHvOGAEDjgIbkA70uADkbT1y/dYN6
xUwFVgSSTn1xUmBjPh5bI0ZGOcNeDeJHwT5Cc9utrmumrknxMLVw7BwHEemppOmw
WgD0puPnr/cXOmjVaBxEHldFyih/NKWbVTJtotKugINEp6EVDMiSl9WiBXoTxxB+
V2xb7TM1prJaY3ZhvtWLj+Juhl64XCfgNyKR6/oUoMSFmNIHsFxTYqeD2Fu5msvA
DACE6V7OidxhwyjtMKktlXnChSUdyC84WODm2v4d+VbHCN/0Oa07vAehJ02nocvr
wVlmhocmZWTIloy84legWiblZO5dx1RKNLCCAZkf6Hb2AUd9FeQ7U3aLcTOUlt1K
kDum6VHOcjWRZKLRT2C92wSdN2cvyxWg4arQp2UVINIusuWf48Vsf8LHhC2TOJrz
+GY1Qug2pJHTPEeLXEI+uKgR5+fJAVgx29CfiPhE+gk=
`protect END_PROTECTED
