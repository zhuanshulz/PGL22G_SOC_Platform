`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kUVrj/AugUeHr5BAdJXuGqVc+H6CCkQitheo0Me0BgnZIg5jjp+3GEIE84Zya/p
RaEu4DNmgxwp2cEUcQuf3Jrb5PIF7Oh7SzsuOqfLBQYqVj+FjSEz8T9LnvHQpTy4
hB4P9+3EBl5BKev1+KhATFzgAzGlITl2NzzmwmJGPVKQ5pgELBo03ugi+5vXtHZg
6atQcpsNLKQFxCtLH0Fiajm2Kl5VhkeP72ZvUhiB8CuuaB5xtBRAITurqvsy5Awt
mkD4aFAm1+ttGXOIVRjhyESGpsXu7Tvs3cf4nEjTDsBr0JQK9mjvuWjWngwZ2qhw
uStiGS0z9fgXfi59nLDNfHrcyBsuXt30pJvR530UX3OEFs5RS3254Qf1qv0++/Yp
etZhWcA8ulYfhB8dzQu1oBp0AEJP2Ud36sicprSigleSQRhdBK3G7JzqpGYn/Mjc
8cxeY1y2Cf9qZA/My7CCWNcbK8lU8XQVoMDmszVOQUt/RV2lxaQPlxrW09TcZSJd
ZIKQPdG2Qopqa9D11uo99NW87b9Sx5WB8FdhS1O53GaiSbWZKECUmrOisetxO++h
v7XWeLjVXSRaQbNCxrCYKQdibmvxIfCpzruv++/Z6opYJNAFZ0izFz6hi4OGqdg6
6vdnzW3Klm6/pIIazczHN1pH1Pi9v3rTT6oSO1vOW8nUEsL4fTPFj1dodCCH315u
YDEFQ9iCC8ko4uqbG2dBekmZj3KXrIERm+FXdxmPnASYUbuvpmOV5DmZ2Wu+uqt+
+GCNoLmwQqGZ7pynsyCFDBoh86+yqKNymjc5WYZDFi1P9DPqdceig1GN5A1eJwR3
PXZMXx3kPLaPXK4iEHtQ9SzrAUDObhxfY9Y6Pt5pVWW00aLrJ05w/nrBWlcDwnlr
VwdMOwFYXgbCkPFXX+yUdSY/nYqURaYFwEzWD0c8CWEnrEPE7cpVVcAr8Q9k5cMw
pU0RJ9VKqqjrOw3C/0jUi1RDxmjLa5+ld/Whg7wU+J5FSakXT7ahQjbEplBd66qv
MOR2pyUg1DRAj96O9kw33ZVSTJMnIuBGTr8QJXJj/3w34bJL/DsVdXV+6AorzLTj
aJq8yzRsjHfDriFbpEPfXyqWIYf+bFdrMpav0LjFczrwR7Sw3XtyJmQd/5adkGJ8
Qe9TM1NkO8PgaDCG8FU9Vk8Fe8/zVImdaSsnZR+cGVdC0w8rxfwRuy450qsnx9YH
wKm/MB5Fq83fkIiuBXc229YA7nli4IO62TV4bt75X430CkOJe+p93mNx2tAfQdYn
mZ1LV66Y7JwgeSOJ5vaopnt6Hoxw8TkzS7sTrs+n7iz96B1eckSAnTxrzEdE7hhv
Vop3tPg3AHYarqOAGIddZOJ5zTQyt6YzHtud++0orDQ9QucB7vlSUv48S0afciXv
JkW3f4P7fIAo2iQFJNnvo5zwPI5QsjZdYuPxRqPI2NKNNXLd/Xnmb+Gkbw/YeDxV
jQD1tGiQNzj9CtUOdF2ExbkflN5XKt7PsJyzCC/iDjE8r+DuLopLRzPYl/w/e5g+
1Wp3uzEQOcNqd/hqpBqzj8+ZAy8VBsiXN38bT3ocLm3emhnl7uvbQg95yyfSUC0G
QPVzZJ4Wc+sf79haJ0zlx+44g9cQEzDM7UdECtGTGhehUk56BmJ14pveqkyYiera
6nWl8Xasg4jxDsSOSKpNLGb+zTg2T2cgY0gMmxt1pFn6x5n8sctqzrofBU5VS2/I
Ecc82jfJ17dt8Dh32hXEms0ilgC9oP/NcPI8DWSOw4/tWRKkmAKHXXfquG4xLg50
bd5exO0ooKdBmoP1PdqMicemH5HtUTf6FtWbEhjyfbihpN/mMRfr7BNKpaEXVXO9
009kGqcJkcMrGyzLzMmrOz2np21Pz9vS3jrecrlZMQjyeUDl1TxMGu06iPsghzIj
2OFeDCobVYej/kKf3V4Cccg+eOAzgUVgzdom5sWaTjUqDWAOM3MOc+kec5N5xPYS
6yViiKqKtU8Mgs/Wg60Ja89hbqYtrpf7ZsLeAJHnRI/U2vUiAkoF1qXzvlG6hKWP
S27od5wXMTSGWEPoZ/h+AifIXBMaLpzlTWECWkyuGE4fJU+Hni4kLY1bFieGT9K+
+aZGUfQR2jOKUd9XRokQvyTKe14rpUyS5UrljqDGn8M5HN2vntDsZVkDLikc+079
hCscTNU4n15cNgkQ4zr3AFqnaEQelZjstA8TvfeHsrY3H5BHag++FZM3BZphQG+K
JFsaXcibHKmEk8ouZw1ev3bWooGF747v2EDISxtCz6WPs3B8IqvAhpiSnLbQJNoc
f/NEuNa1LBuCMEsMFyA1sxSTU5/5jXICnzMUTEbmHIu+lHyFjM7OEV6AfWjmsTpj
mlMfmvjwj1ISpPep+itoZYTl0ecxA1fW72E6Jyy2JBXE2mlKb9YL2yfDNf1THJZW
yOov9r4CDEl2ve3ImSxO2jIXHjOGd3Ot+e8BFb7oWV9sOfNqfnyrZF6A1zGUxct/
pCBUqg4yhsqI0w8Cv3Y151Awg1sl/BeqP0PG+XmSbEFlP9S2CXYvB2vxEKcIztRv
F1tFJPPGO+2gO6fz+xFbM5rRzurl1bRBWaHyNG0Enhi9DHdo1i+NH6BFcF8NcY8o
j+fFKjkW0MrKSRPkz3mrgXWNXkaTJRKm7YQTbRmt68QweTJkg1D48Pm0IVRAMXg/
zL6HurN1hlxVTGRj3HF+SllZ5PRviXq0A8zYARFu8hRpWehfO7WOFvkq/2QKmgRU
2mIcdrkZWfAFSfkDgVXj2PS32oYap5c6zOqbHtKFsXOWv7g9oUX82OuMdesjXeak
NQp+5fHYP2mqgf8cK0YiWPNwXzI5xlq1c4IVGVVsR8cU8h2RJ4xkJuQRfMza088P
Fg4u01mhOvqRYkck8xsuMxhI0JxXGUaYI5WFAUwshg3gqHkIfL8n49fFfIMqnDNT
moh5Ld3I4oxB9Kqiw0b2SyPBtfPXqNm/6rNdmhGzqkJLnD/kKZb/q1wvN0tc8OcG
MPDchuoHFIisri6oYHkbpl00qCriEushdsZDd3EbqivXXuidzVS6AJXsu6MCx8rB
HFI4XbYZPMd+9vqDPTPLSL9irde+dOle0Td2nI6ikCstRqEgAm8dsh+Rudy9uR41
8q2lyrOZe2ldFa9RgFkhp436VQYK376ejm3JXB5S85dKJZWcZk+TMcwitfAnNHST
8URRpu+rJzqpgjr0h4+XcoBHmrTQVH5hhFgLlIZ3N/FX7fKX9gGYflqV7lRzruhS
tiXiMG7r8IxdOm9SAWiBTRIQLEqj3YLwXS6lMj4RAVx9u64+diVt5xr8f9IRzd4z
OduLBTaC/43sPZ4QVu4zfjeeINCXL3AlcQguSHHirSMWO3RayD8ZG+DDht9r7k9Q
t5qL1OfiMbKMKBSBY9aiMHBlh6GJI8lvgxXkPOmtbvxIIgEOopf4Y5gmKxuTpAna
KIEGlThg3Ddr0YHGzeoddV8YNrVavyR+jzZc6hnzmUlIVeMakudSQhygZ2/xCwY1
GzsK+PPzrQpzbEyV7ttsoKtW05TDHjmF1Yj4Ik2a59wl/wGQ5VdldCmrCpItct8C
cXy47QtmKuAptk1H/qPqGz3LQ/caKKOZ2wz0etYu9/D7VMxLjXfgbksK7igBW9Cu
zPJAbCM/gzsAvAZtD89qvAwzbZRnpu3bO0SWIHKbo/Px7DYfWP9uOkHzfEqfgWq6
nO35u0Tmo+v6WRqOmeUMUM3bhb5m5Ti5jsAbII/PrFhMpvGDvL7EkLkqOXiQm0DX
doVxPj4l4Ik5leBEpua8mIEry7785eQvEXVmlu/+imiRQORa2RSdxxjIP9lUokzQ
dlw/y9vSU/LP1Bz9CnRQW5GU35j/vfEhimf5KZaAGPBAmwyoQqAiNOcaMI5P2oIX
N0JIQtdW3+ziPF7JHXBTA19gUabbQPoIIu2KlQnwoilDkn8qeHDQtMLDH3Pny5xC
kXsrRSMbiLGij5r0cIT/gcu3IK4S8djoTe6WwpMaXEaOfhsTlSPVLzwm+plqglHI
39S26FYxCkJpnOv4ECAIMAiGvf9zG7DTb9tU9ZaeFmXQwo34APIUDgGhAQ6Jb8QE
lV3PkiVddUJp5EISG5DlWbqdVKrz9Mi7zJqSIOFiI+IqH9mkzTz/NBwQJGd9zbEY
nCLfWEvWIkK2Qja4YyXEx2YatPc3GpFm/IjdIXiL0E2szdLU/oZ1pkA3EnCoDCKK
gHRxnUoZ2QpXiBHOvN7ysCtQXWUqg+y7pAiB+/YrA8PWC4i+g4nC64sewrS3JLEZ
sxtc4Z8EQHBHfnRVBnXU4u95DxgtVl4mAAOr7hQMtlleaBYhCiV8qWOP+CBKGph0
IITG/KsWomqgDV03hl1EZYKZUBPAgj38/7uokbMmoHHpGhrWSh+rvnEXSKb51Yhb
y0SfuiWps40XWyCw6xMJoeUHFuNFxDHNGUEVSW5QHYr460t/4pbqNPSTtaS77SqG
Yw3qva6bwSlKvJrNoHiMYKvg9Wrcgu3y918YLz2MFbrY07YZnMi+fC6Wi91LZgev
UMqcQrjgUMOQeTbIpxeIeUk7Fm+ox4+FcGg3nYUhyTrfhX0oU0BL1+L/9AyRLdzU
JGicq3lNYhgXHxZT3NuOwNny3V202lvlgK+6V35SoVFTZlDsBaXh/u/Qs71tRpjF
EV8BOEqM06iMmUTG+QyL69kSOxdIkKmGRLKNvavztcPI63Uu0/bu2dUQ+3BVW3DE
SXIv39ECX8d+Gz//MwJOQFhqHg8BuKLE+aWa9QDy6TC09sb3GRAniycWaVH3gJHP
VBjzshuQvGYaNwUlqopGQ8LQCDvd9wBWfoTM7ODuHMiW3AN2fpOJ4FPKWmhF9cEX
yvhaOXcp5c6O8raY2lMGU7A0JQC6Sq6gctu2dmZ2g15WOdpgGZwteLI0fmOcRMOQ
Pm+tAbeFfGwndgHMxif4WiQujeFZFw81+fy3BDeiXJeBQAvvvQvexiZE3Nkug4pc
njWu/MOxnhNLDt9nREMfCXs+NUb+QmQ67teIawP+3OX3cfbljo3QbSKVuAY30tNa
i78MwI3NjihHi+Mkf2vLd+3FSmZO7h9WTGSc1q9TRCPYgYlB9Yjso9J8xOKhk6BA
K31M1WZrz02o7LYn3KiM9qktrJdSAozvRpKNfAMoSCCA1ho2fX9dr0+209skRGpI
zVluEdv88HNmMTSWekTm5VzmPfS/ukE05xb6MeVxNHapZTYf5XsC4EinBcwMmG1K
BRSiIJYWNevBhtEUQpGKhbfsnG4rPX/WJ7xnaTAGqxBm/69EQXkLx6DRynGfR4F1
tpGb5Jm31dHcZ3ILGM5pt/+MyWOCAcFOsGA4y8T8u5lsVbRT56pQcJMbz6nZGhWZ
S1QqNfGxciX56CVLWCuEX0xKTyMsjYoIWSavF0gX2kc14KxcxmRJnrfgIy089hBr
3oVTzn7MC/HVcUeQOo1d8Fwo24dVcooKEscwCxtABVyJ/0g8dBwVSotM6KQ3DkWa
1NWo+R+AqzES7EWgGc+BcT7Wlj9Dn1F2brQxTW/UnuBnGRJyI1QKTmlbBykNQqr1
mhSwX88b+bwQRtVZbfLnoPkbF7cOaDi2jOoPl4jBMluZRBJLtt85sCb2y23LUw8a
TqhJ5ZFTj1UVvPlEW8D/c7TS9bswWU/dYglIMKB/0z9x4TqOZCETBJAudXj1SC1o
5K7pQjlZsFVKfleoYF23mYwagRAWVyGcumrOrANurkgVxicWm17FxFizpva6chH/
H0W2jPw3TxZXY3E3ndJsB0xA72+DZJ4BTgTpHCPAvR1xq5MtKSTvaKxrXmfp5k1V
XCp2cwKzYgeCbwuGGi+BjBb3xgq3xMX8flPnq0puAcT1MvAEmUvg0trIzBCpbSO2
yrr8PHhG5uTti3BS7rmYQkITmgxYUkYj8EyeAdOb8cv7rZiOKRD2mFpVyrnwHtRt
Mj5VhmRB7M+82hZ6TogHdN42CxIFXUIpnL/ROaK3vczVEoWYBXpYDaVXf33hoeqW
zAlJ76VSFr0diu/3PMrqopnur7D8jLPZVncrzeqtYH2cMeMKjEsJ7o4DJhhNt1EG
J/rzc+P/f+zKLHkz96xKLdpH2HHaoP9kKaNYfBTG5RJ0xvEgiuhhuIgCZkiDIzjv
Aiiosxt2Vt8Jk3bomz3iCSUf77thREM0ZviOdKwTEAA2nvVnZFhFHrr6UqFdaEfW
lJ5WGO6+9W1PzdHHbYm2jXrRmH09XtPt/P29QFtGBSBhzCWe+xB7lzorH/TL+/HV
3zozzFrX8VI+3C17q0Z7jyRqrboD9Wau3KUrOPPMs+An0clx3oWz+8CaZEUjw+44
zp1AGBpO2xkMJH+PDI9lZ2gnEdiMTGj6W9V2DwuL+i8JnNYz0WArmq+AzD/4WSpi
qHUKZXBE7TfhJlhwa83KFk9PPcEv/SQt8oZu0hV9JeRdeH9o4+hfJN8r++xL/DIf
5fM/Znm8xaGSrGLcHmVOxG/b8liG27ltmSy+J8c3+D2aYy0Ndof3o8jZVzsbBysi
YPtFZsnwLPdLgf+Ok6AGTc9/mrTJGyvyxdXwzGBNvETDrQ/TS+s7U6HiWmmgSgWi
jIV9DC4aM7KkTLW/bNjG9Jde17CKhts/MJSuHj08peXbIchSvAecpUhblIorY0y4
OaL2GdLOxodT1ZfxYgsQzcZYRrxn5+QOvH66BeOD6FPKgriNSZWqAZKjciLsnY2L
bJqv29k9+k2vw0yRG6eIM9lW5PXIcKUqZwNGsrsleR1MLTuLHSuG2PIdkIsOkRB/
8ZMT7cwNxrcK1bhG0uT1B/F7K6dqB4kUcBXlaux+ho6VwkfdO6XWF5Y4rwDVZ5dp
eidYpCzWOB/zkSqyO/Wz+UYAaMmQvABM4s9nyJ74gy79cKdDEadQfw8K4o6rGVSS
6sWFc53ZHbpImkw5u2WMTTCoBYHlvGAx8TZ9rhVF/ULJaFAg1cvjspaeBvUZIF29
0CvzAeaxhQHrKi7ZAvKh/OIOVt7IciJ4/j49gnMAt2+Ra0QtUUU1QCrlCH9buJpJ
gP+zmugkLtXwNKdw/ONqPgW0ZRmUgi3skjGZpP4z4bHdnmumSh2062tjBCDPJNUb
k/8wVTj2MC282JaS3dzGe5XegE6gVH+O781VSxa/g9VMDD1akOEj52N8X8dhwsJb
Kg8jzfy8CjTYhOgu08I4cetnx6nj3oAu5+CldaQ2iXRnRq21cgV+Gj3Wj+TopsBJ
luFcdvfc33aurfehHxJ25CYQFNJo8dgbrE2L0ACNjkb4HOgca+CeRZFGsvXAYK0i
M/aaToFF9Nys7S1MUPwfxKr0eM4kb9gZrYqbvpE0Z9eZb69HN5lMt6tyOateXV+a
ne4HmLjXa43oQK6CgXmoJqpr2MtNVPMpYDMWP6X12NMiuvkyinT9lKZZ8MFP6ziO
7oUSY1VsSjH14Nrvtiq2pi2Vq9+nHL1gqSe8N2o5CTOrANKk6cCXqHgQsa6tH8aN
D9gcMhEUqvb9sBpBgLsax0BDz9DQ62T957qFtzB0FNdWd4qWK0f/8vjea81GXtdo
ZWX6uCWmr4f7aFXaY3c9bvwq80uIN4M5qIbHwErdebv6xDlZvruBMCgvFHJWn9nY
nJzJV99ip/ArtizXL57hmDHQWu4n4qQs2bL7hKs9jLL3XJzmKF9HjpguVY59g3tn
IUt8Rrp/v4HL0TmXouvGw0d1TO+LDQSNae1Q/F1QPJ42PmtWFmaGyNbHrum6LiFb
QiBzUcAfZxldCciFCDyHy3vy0/qpkDhWuTZGfpAwTfedUviZG6EwXDgiWMakzFff
L0OeBHMZYdwStZfE3D9vwLqCI5PQ0P2pVvOcf46BAP1ps4V5t6jQnLM+ABJft8cE
S23/14KArQAVKthHdqlbHa3K9+VVPaHxD9wD9URtuDgxEiowBx8/eGEcV3j0/7Vp
fjQewhhpsVC9W87pOJDWFEAP0xqbRGKCNRt/CrLBVqZn/dESJXfEncoVlK9aTAMC
H1bobeQnLbpTfz+sVv/p5MdLTdjcjBbIFyebIB6T73yaBaGgtdx8uVBwxX09fJhA
qG84V8MFjp7pD6kEYGLg0JFnzyuyo+y5rmsUDXBKqq0lrHwhOlqG8mWviOdLFL6R
kCVRwBdMTNzR2D5Dh22DVXJX0Zj8eE9o5OykwWPLe2URDO7PD+ZjBJ2kypkKkRgv
DEgQmpg5Rc1fYWPXQyOVPku5miajbWOf5urlVbL9YzTrQL/GDNVfdog2+6UfKQxs
kEwqzSF/O7MzhVf0bTkZueVNQ8fjLoyESRXayu3D8rrYOibiq3g5KpDgFx+JQmGW
jZj+g6jvqNnje3QOn+WKnGXT1giFvwzia01pM2HUWMEyKbnjIpE3mkez3ZShhO3V
N5Ge7VGO6VMRPbAWueD+VuUBHxT0Zgj55s47xS4nFGu5hWU28uSKevrE1kYY/os/
mCCEyeyR2a83eXijE6Nm5BfyK9MEyWvDrz0bTJvxYirpnqPdbBOcQ+Wlc/CM/2h+
GbViycIl3fWBANcM0lf18fVkmxvagENZojOfpyh3mYMhlBY+fwgrWmhb5ucTR6g7
chq3JG7GEuvuRGIdF18sw3cVlnW3eUkIBUqUWXR5wgHEKzdwtUicl2Zs5NEKTiTF
00YejHCVbl7FDjhXVenlQbTHsLsB7jB1Rn4RmHcZ/nIDBwGByhwBn6He724lhb3Y
Q6NiYJzO/ycFxkD+jfaRVUZI2f4kE0kvuYL4MuVaetaYPwa3trn44TZPvQkyF9EM
UkVuiHJknI+hq1rImabzFMmsVJdLbX4KLa7E9l7CSAornEZER4UwA+0UUcpvM8UO
bFoyzWCYJuGa5cyyvwcZV8FFHbKDNMsLNzrJbzRjAWW2AcTogp08qm/NuDHIiNtY
W7t5lsevPeTmx0pzje6kUG3Q3HWvmT4zR8GoS+0ztn77JlBKPUy4OvBkL5SQqr8f
wmBTOMurlVdqPoEHhEiNmPiBPCWa5uEKHvFqH+zZb3S9Lj8DgrQoFvaZKspknuJS
RrE7uphHoVTxpjIJElIeMAyoWohUnzyON+ycgLugfTlWyUPhkruB4gD14oJlSigL
o6exJ78ycqgsByLHzmnDpvMfOilZ0JHwIuKm9zlC+vVmlMj1JXeJGQMd39Gpnql4
TPqydKN2vJsrpjju0LfpBNQMkFc141+YuAGQWQmbkrpeKy6moUURktFrZCMFlLF0
fi0ZkXThCwWWC7F8K41IrQ3i8vKQCKBGtP42V22D0LkkU/7d5ABXFsQKBq1CXny3
DGCosQHuWCfiBPYDwQoZBHZu+OHWeVsuU6/Mr/rLEHW9FX6kZDwKg4dwyaqccM6l
piDl5rcVwOWqgs+/TyW+b8FI8wX2GPT3lvVu9y8ji3NJJuoibniu2Sc5pJw3Vo4G
gHlehmqu6zL77/mLVLTRSCiFHxrUYPR+MzutTr6syhnt/fpiZCw7/B6n+zakHmlx
r8Ojb7GpsxvPEadH6O/Ln6HmjW91O8BbMI+syN0wjXF2wL8ZLgM79fq0MPtqW3mB
ALV6qJtgqLzYaHMn2QVmB8Xs3+mLhmWKGIbDQ9W1deS1GLkFpss5qJDCk6SyRjly
eXKFRpAOLLLjXJcfcVLp77HXqIy6T6TkOjHMr4SfBFrxvsGrNCxSPGWVGtpRdqSE
HAasl34yyYb+EWfhT0V0KDHnO4UOBideIP5Z038iA3DNts/CcpMx7GsRBYLkUaHu
Uymk9TyR7qC5QVIBA4bNLPxfRlIafa37WQ9xG9ht0ILyWF0GFx61tnUfGgpR/n7n
5TYXImvve6Mlkfn8WUhSwHWDH8giShuNAfEQ6yN2NcTRdwZFcmElEnVLDXkeJOf/
Yd3k0DNhE3ljine8vfBd/PttGQ027+W84trmW/xt4/kwVtWRGlSwOUhhVVsT6EcZ
P8kr2FWAuAp9f6ahcr7ee+flUfy8F+NCC4DZVtAa0pVfHv3bRKNA93dn638yFVei
UJVmFrL3TC0HUMwxjGJn/3AmYKAovs5Fv1KDP5jFXfGkBo0TgRvDskpmo34DfKx9
ZOR2SGLsycm2N9lYej99xnyCYVQeG3pZB9QbMPjrukCEtGzUVdDKV2bWgoTyFP31
SqPIDs5p14zUKvjDMQHdi9jPuewJTIYdlL5er/lSqyVmFUFrmzPydd61OnDJOtLb
GBozkFbraZ43dhBcxQ5L8PzJwg962MuSH5JkOFs1Rk61rGATCK8OVHKYaBDswYg7
kAT+1lGbprGQqyPXn9eftav/0AqcQbb37DBPKiHZpQn6Zt4m1eVkN4yGmy9ER6Oj
vwiNHALLMRENsosTHBlUG5R1lkLYXtS35p3AYcrwVp8DLM1pITEtLVCM4/aBtW3N
fXJV/hYbO8okD7Caa2aQ+ml+6HlnC/YHxgHDprngYzFkQlnC7z7CekSN5ptGk13Q
KW7KSsktfztU4YWZGcIlKBMozM393UiSGIJ6HFE2waFQIFw4tc8UO/EeNcYvZMSW
qctEDtYeSx4IKi1FH7Q2X+d9xqo1NSD/OImpdhROorb/msshcVMfWkhdSqwAiWxL
KvAUGpuZTyAQIeLdxjjBbk4Q5NvFufOa/ghHnYeouIi5jzxrh1pEjxK4Ajgsk5s9
PPQKPaOlGR5jYWELo/BwU/Doh8u+snwr2y5lWGhXEnJeePdASgKIUFqbJ1vUlkSH
KU5NigLDb8kbRCQxbCD7BELYnT0VkPZ1GU5kJOFBb1W1MkqLBYHj4dP+PHhv1cMK
ohv79EF2LpMDsL6pZISsWiEYgzstfKFr39vtCdCCLdwdx54JcBit7tjVc30986XX
3vL3+ryET6K/uisPoLZDg2I2RVmTreAQ0mo7oEv/C+e4VF8siSgC5eGcWQsxo/Vn
IOyIgQAmBYt0/vy4Ne2JziXGI5grOT4MCvucxIObz8vZLjDVGwMoaSQmCfCR+hQu
l79Gj2z2JO5w5KJfoWwpyAcPVj5r0XS7aiDJP6ZmHpMLFmo5ct4wSUFwz5QjpIhf
jv6wUNK/V0rtohTGIMEYY8LP9/SBtxX5GhSAUVg+zjT55RQh3MrHVyBdZwONa7iP
yDlP+NL9LZ6UB2MxICnCdcx2i6xgBe7hHB+u3Rcwt9tl5PNM8zdcGpI0d1j1o/9L
FnAvHilE8wQ01vQF7DvPMzuka/3Dzs3yiPa3FpHvB063NrGj846duUHV7Hcq5GoI
QnkdFy91JIqIsr9ydKdsHaoDq0zsEM+0yQGvoM94ymPk/zuvaOSyrKN7H2CqxCsq
Eh43JaLlo951Hr6O/JnLMt+eD1x0Mw91ee1CemxgksIzt1HiRuprEf+seIxcsbgN
yZNZfp5WQgg/shRJ1OjL1434SFfecridZII1KX7+ONH8vdCDwBlFeDfPHDwJ2pMr
Iud2akDPrMAUHfk/ZQoCU+SKna1LJzu4pxIhtwk/dxJzjWb5O+GaC/uwk5eZl3eV
ZuLqf/d+q2KR7HOk/ct9/U++u15dTDyP3YUxHOx8h/U9/dKSuPHOZRaOPop39dtz
mb1vkWtfhsaUfHJW38O9ChBLFw0pLzSNiSo9R2fJROJ9/r2dudr9wQu4YTItOxpM
Cp0+rYJ6cX/UfoFo6ff0Ds9AqCczO12SylnrVHxuDVdJbAdZCQE6OL1y+0Jfc0lX
9SNIJMu1Y6yyDE6vgB3hxYWJL1+eTo7WP1HpZPv77+ElFEzuabjOcpm/yAwdTyq7
LXKDxB5drSmCQr1Cs50LH2wJ6aDDA+XZHORP+0uIIEMkRqU/cpoLM4s98oEv69xE
j2lLNkM6JlRer9ujvQ5exJflOaP/EwWnKszYqGPvfHvf+Y7rE3Cvh596DAOLQJRn
s4ZtJ2E8+qd1KLc7ESOZo03kifg136u0o51YVQjqXuSHvU3LVIi13mBWjml23bdp
CRzZ7rTFhA8e2Kpc+xSx22x38Hhe0wuj2wbZhWd/yperiGCBHce08axawQRW9+Va
QFyMjCw9pWY7/TIo1dickQYyBMwFzo0x3QlgOCjlnDlTaWlzMpKwm3NChXh+v3Go
6iEwTIXySaTnYNuTscu0s5CtEwCsbzkhGxyJaVL6PUUVSQNweGXZ54fbORil9cr/
lxYq1G3a4bGcQORHM2fFexh6tK7aNiPt13OpvRiJv9sY6KSynDCTtz4z8xD7XmVW
v+kmGWcKBPAwgf4g2YMazHm0PYDUhr8PiCRdBa/k7Gqu3Hb20T3joWqhFj2/TZ6l
YI9Cd0GGyzcH3+satov/JcELQuwTOV30p4L2RVwBigly56V5TxlmBXDlW1XYDZ2i
5PDVKWuc5z83iWBQf2gCI+4zNjaMceqNX62U7IYsKGUERbNTJJ4qzRmvJe4RTepk
OTk5umAxGKloPNOrNqQ9fFIIRXP9wzv/hHd6EEG/LERsbWRfuA2xXtjLtV1TSF+o
evSj9JpmZ1UlTp+IdDMOsp4jkmrohQ4/mF0Sc/fbmgZRw4Xqz6vP54P0ovhsCEhn
1TP1sHC3XWAxFEEIZrjU4d4Btwzy/52B7HDwsUg4wcCje0y7ocFMTdnyajJ42zoH
MntamHpG8U+vvHDQRwrUlQOjB64/wJFjiA4mQ95T4gLBs/cfX9PMCEL/F9S+TEpG
TCj5Jyw47yzl4DNjZpwOk3hQrL9dlH5TnUi4laJTyIK8srrow0jizXiPj27y/DEF
KHLT4UjObpP/UjegEmu+djJ/HrxkXPCDI1eWtT1vCzGFWt3ooeLZPQWD5woRgb4d
1TYycOkm5wOvPh9hLRm94NXrNB3dUgKoT3JnJv+CHa3Yt4uoLy/ugRTVXosl0ZDq
fr8+ZPmvEpgpNeswBqnpxsVmy81i7S7duK+QQOZLJmmriJr15ZLHSg0s/jQ1Vil8
TxL8VpJMLZ2NDSigxZaoC83/Z3bnRBoWT0SATthGT7kw80yVHqkTmYDc//k5XTET
wBfYOMhfHNevU3uM66WFNauorz3lSyCQ0JdSd+5wr/aMUj9WurZAwnuh8S7FkFul
rxVhtBjWfvcvVi7AmjVxjgq8jSnWnBeK/0pw3kwDaLh1OAm/+tl4oNwd2kYN94jI
v83NOiBHpWtpC6ewdw5n80QaSwrqzN6z52BOpsjH6uOMvCYo891z/5Pg43QqxU5u
jP3diZjpN6aHmopevsnLyntMktwz+NtY2tWrQh6sBJoerlz26yU1eP4HUejePH60
6TT7MgTcTdiQtA2vZ0DyBMqsL/H9YvJib9ker18ZRhMNXPmvz10cRlSJIhbO9yDr
1Qm3w3CM5t0xAfb53ZN7pH2E589qAVu0r1qY9w6a7JP3AqIOQvVAL1hn4QL76qNy
4EZAAFRmKlNSnYbsmQutjmVVX9tOQZ3o4hklbBHQbB1ISbkJy2LU4kEYMg379tIH
Jwa07lpskrEbd4nUL34zn2zKX1GsiTfvXUY1D6aBD8/Qvs2r2Umcx5N2TxHG9PAe
lo55dFVLGXfCC/HcdQPoybbhCRLj/UMN7Z+r8NCbUCACGrzC+AviXT1w6tc6LQ4m
4QCLwOZZB2D4mSNPiWGoAcVrEwGzmD22Yih50eMmJ4gkmLSuU/IA6plSFqYpIADM
ClQLFo/+R/sZ1zYoNVwcxLBir/iuea2Ip8js2JW4J9QsO0/Qn/bJzJtL6PljtAzb
Kg7lQSfAeO0hXShZD2CgmVqZdSOukieJs8pPmLcRdkGFNRo3C9CEP/gN1NPyfNGJ
mq3ovmpkddLzuBOocn+JvdewMVGI1M3E4Yes/zjQLyiM7InnqbUUIB/NPhsF2IOp
09OC8hbXeMs7Tjt93RSLG2hVgug1Ysc8e+HZP3/mR/JCIn3RT9GtwI/XmVb+IBfp
pRATffTtn9J4C1zjQorlsXuK4KuebozIDXjHdTeOM+nFQZp5rGV0PD4WIdmK4xfb
bnXiMyk20MTxHoUgDpYEmLQZr4trrAUfsBLJihZtDl1oNI0Rdyk3pDHBvCViqxUX
bDocBb9aSF7jBWYuUpQ8s7jUggUC+npMXwNH1qSXUzhuzxMQ95zgmkmsbXNCtNnW
03f9uP0NTQbghBsU4jG2f+WnIoAoJVy7RQtGMZmuHn7C+EaVf426kRZLBYFd+Rj/
uLisa75jeZyCN9MOkANQ22YTxthK0qywjUVyFgwifISTLe3pKTKT8/akKeNJ6e8B
TN+32mukc8wHZx+PJutneEj3keY8Gr2iAbbp0gs6gsLl2q7QvnlSDV5+qFs2hYhH
ijjAHhF3fFCnJ5Ip+W4MXusWqmneg2KtBXX6G2WL/Vd946WklQB+tn0s0WNpFODd
AdduxiUhkx2fqrjs+IcHaKoOo1P1x5/6YfrQvWKeQ7qbE2VYSxaY/8X/4K+QJfNp
nZO5GTOwY6gc+QdWBtr+YEIViluWZdy5Z8jFPGv9wUArgDEZ6OT6sbf2sF2zCJa9
Y+fLjgxfCUMO+9DMjXiblHuDDfr5UTlS+TDWLtxdGbHfI2n+mFfubAxb7EalyKtA
2cNno1FeLz6Sb5xuO9W4QrjjY7SgoA5eGD7Jw3qrMMrTeQ+dG7+Qy1EDC8tWs7Yw
ISkYdCCdqvcaXCQtSCtnq9rHQFVtzJJshSCekzW3DwvKc8jF/c4r7VwoZDp0FuOU
sJMdc3ieMMPXdHCe3s0qPOZJc/0EdWLGc+ceI2+/O1tf/Iz2JQaxL4nxgOTIox8X
1/mggP/Pm4NgzdiOw9gHTX0wNezhvkmTeH4hWTzeaqYAW1+lpeP6sefFByaJ9sRU
+QKcY8emWfyLB9ZC9YpXeZGX4wLs2iMRg2yAbqwh51MpX/88N7TcuWFA3Vk/uZ9G
c+3ZjWeV06/D7SUj8JhaZay2suv1OKNRFn7JLFOEmeJ4p+81TgWMg+bguN+ojLui
rjOfmGyzABdjeXjeKiTvO6+2FXsr72EWf7n+h1LZX0o6Qu99OwYIr8yYukw5wVHW
P6ymvrxFR8uUFp5NK15gZkYzZ7KIpOdb/euvgbckT20mDhiPHgWMIjfFrchZeX3/
n+wqZ30S/gwOmhgnraaPUc6xcMgg0lVTMAF/RouUCCFLrSoQ0cSlOTlvwWWBCoTP
vwpo0g6ZqTslNaHKFslNwtLZcQCK0q84aJJtPurDV2D6BmMDarWMIGJJAgwaO1g5
Fpmnvg0zKCPyxSgr65Yhr0d8LqZXov/QIZ44/5w/kwXMqf2Xru0dvvundV09Q31M
iiKjv4oLLJALtBIGt/iExXlNs93nDyrn/vgjs0W26DHGrSW6KdhSLd8mp2MkbZi8
U5iBVfYO77pjztpwsm6vU4mmwTkTTaIpW6G3CQJrVvvQyC/nXWZI2UhmsNNzqnb+
vcw93aaB0ylTqII+JrYsbKbvgm5yJ1uw+nu0Gukvh0A6JLmCilWr4KAxs3XM+tOT
nMc+jgwjM1i7iGI4XHLB8d/IzcxSl59NE/f0VWYShaKOVTwxc4PVpV8OCXLBdhbD
ejO53bZ2P6p1Az4TazUteXv2snQ8mVBaUP+L+DLkFYqhnNf8Zqug/1ZJX4sIJpYZ
FbtSX0bMntJnsV39Z3vRnVMRHyQSuVaed05U9afF5Elh1/+jJN9iGvNJ7lkJzcWG
NVK3XBUdxEHk5c5GgQU+fhAc0MAvqiz7SH0NOhUpHMUzINYirgfOgkk+naRAv1fY
kHroZ4nDqAwhUibtC95WJawHdf5cAJ5R6kYH95rIH9GLgiVuS2VrjbHCwOQO3ZML
8IRHxOU0P4z3JDqqjfLJJv4A9zpsoi7x4nzv1kyDgki9SoGXc7vOAcNW5Ta+8A2/
C20wR+3DCKPp4SfJX+nxi2aWlrMKwu2Tqxq+TZvRlgBuY8vKkRzBymFN5hcwKEpi
s6YX1RjjBk73PaCac1w/WNG+MKxC2wTkzITEYV8Rf/VZXZg0GU+8Tt+o3imJLg4P
2pRTokAVa8X3QtfOgFUXk7fl7jmrmJz33UXJtSkeTOh1a/H7jAKBpV7AxCS2jXBu
z3F00rgtcVnjxRqmWDhwKixF4KEymXCaaiNYZ7hNn8QgR1nYUPN80o/BIDY0HTOG
0HA63DBueeQCGOR9KdO4x6d/i9vY0xrjdpkish/W2SJxZNQNdw1vMVz6VUghzOiu
004ynNiHsUwHDjw6OjvwHChcJYhjuMKfrux9sDoiDW479Sd1sREqCpnAsGUxJwg1
nrC0zLEu3okqfKCFFC8wkM63njCL3vZWqSIdd8RUn1CiiGUU3qRjORkptDCphw1M
aJgHp0fMHWl+JwFQMr6rLW30XHN8JML4gev1TFYkPLpPFWByJf4O056RfMM4Gpc4
7TdBKp5oYrHS3An3MA2Qbj6SERgniayeO4ADNP/uH6Ix9g4pzEcbVOpziMoPpAdJ
pigQIwfHpj7e0Fdm4VKacMAWFfDl38+dhqvNgcmO3yPRY+Ee1OOZHr29ACr8p+/1
vNfpGMgBsRmVwgmRfarqIz8P9ZVnLxO9uOF57uwtgyuLijMalhVcIYigXXUo0tnH
mURBGNb04D+TuaAuJQF0yoGc+wjT/Smq7XetUTv/DLwq9p1Hu4XEQyRC615WK293
sc5SKRwkK8w+RiUNzjwU04OGYu4CbepZzQuNAyI+gXZehX11tUOq6FMV9Gq8B1qq
C1LZuGhdXiSlBnaAACaZMPXrSuMF62toQ6qWdFPj5g5pkVMLrBZ/Y0UbIRPmybc0
xoakQpmOZcwQsuE+tR77uI+95m8HS7wfZzGiAyM1yctiGatbK0afPwZEvSNB22SV
QDXLMCGvUq5XlShHZkpNS3z0MHtgZcLLOHxZ9r673IdThirPsUOPrR6qywLxCjIx
CTuJpgmE8VgJRm+XwEIcZr8/XeqxkqtgoLX13Hu8pigDQWabbjoVybEA4FYdX356
wJ+pXqG/RwbgYwE/x5HNWj5wyUmoAz+shfeDM8eD4GfjwLZJFq0HoNGjyrF0uCy0
NhNilfIDoFPBs9pRs2JRLNn1uQ6tj4kaaEmo0xOcZm9O4waJvNnzgT4JkdhEuueS
GaxcSsbNGbYktf7JvbLJ6sJTtanRs/dSQtY0r4md+zgJwLl5FKEZIy/C10UOjzHr
Th4qy1cfnke4+btSAjR2rYmXQsKsXnr7r44b4id9CmldkL49FrFU3kYNbyLSZ+dD
QiGn/WH558UDZ+Tq1EodMKf6Q1kG0yQvX5xkuquNUKoM77cE7XzOP9alfNcr2HTs
VoTM/E9sJI4JoydY7cfqehBJZz5SdjaHQWY45Jtqe2/JXur1mpq8Gjgszh8fyaiP
jIa1TugtWkmzc8efqTJu64XQtoXU/usDMs4GOVwDO0VwwYdcxLIZPLfBG+rgRWTW
5+PQ9ZDa7OsxtXpe+QhumTxteXDHRAo+OA9R6EJmOPpdte+50Avs2qfXSEQ1+keJ
6vSCOLD7pq4M6/KlarTwGBQfge1rgt6QQCYym/55IIlAJKInGV3PWY72vPxl/YyJ
wv4MyAvEFlp8clidJNTPLG5aHBpM44UX1vsjKZ/fk8OWR4XOVOXbFq4/0c0P/RaB
0h5yJQGRsyXm9Cfr6HVzqkfNKnD22P8rubwOsZhJ2jzrbo1NLNuO22fJUvZZsZJN
m0syBRvXj3nR06pSznEcolHhzeywRxAeUYU2g0Y0rLsgWEMfTmYRdD/gdWEquBwj
5uUrFxcLqfeJBIT8aF6JTZotJDu7UXpTXqHw2K90gNeo0qa8e+FNT486ZkS7Zlcw
2CJ9hK6aljbE8xSHjVp/H0pkDYt6e3WuSnrLxM542diHNAYnNajfy5CF3NCh/tMk
mLhnrboFiYpzzfvssNdyCo0nCVdOORDTHVgUFfDx4i6g7YmwTlea7szxBDvOzgjv
IhEuHzeYtgyZNZKL3u2GIy8k3yi+/Bai3YoVVCGfWECn31yimDw64LXFVxy/73Kg
kRCiRhbafxU8xrxeHIXwzRsg1gRN6jqPR29onETswl+0PksnTehsctwr6B04nBT4
SSC6l4lfpse4Uo7OoZ3EM8MhmMPcXNkgC+Azakgj0sqwAepThH5y9lKJmhdO+woR
QHDrM1lrbgpVEr6yloXDSTH0g48MLkWjBB0F3H2w7QToHJ1Lr/UfvZuoXiSodhCJ
BlvxQQGU8mENvelTcuoSRwD3Q3BTRyKEowEbV8++1fxAACUFX58h/oKujqj1V207
7FjmFslROGpO/O6Ofvu+MdAmyQuWstFE3eX8qDBdjP6Siu5c4DNn6kXDOwRhYRvO
KE1vfhKI/vV5YJBMnpVMX/OSl88/M9mZ1ZqhfVaFacv/FKr/5WVteaB8IYvhzS08
a6L6aMc3uCR4sFLDAJZFT6b/0o35yoRiIshAv0DGo7UO2l5yFxhBul3adMQ9c7fb
C93Sr3BNVyMeNeZJqIGvFhYNeK1oY/WDIxnW6sXEhfhofeOJ287RKBegkBE2zfLq
zMQnoGawix5YQjkyLF4WmS0vkz+tt01jOpa9VyfwIkNtoQTMDPZHRdCJA/nuobLc
paWFORD753SFmm7tvrJOx5VNePXMk2yr5/iij5pBVaRh1jFxEYz6//yfLj3fw29u
aqNsY32f/HlFqaGi8lyY63VkUtXur/R9huRIqgCIrJaFz3rBSaRAE9+e1K8q6FSm
18PvgUMAW6clRn7AiyqIaTOJeCkMHIdQ7I6K1USNZlkft5bE5q55GJZCA8MfV//T
lmej4SjsHBa+u6XRgQIZpWnkksMudBLrTTwNw1OMK7I41we609og2KuGm/L1whOt
aTPzKcQT8/mJnGbV52Smp8myQF9OdyUtix/B0EH5RGPcARTECcAU/WV25vO+wiUE
N2s1JpL9tLjBKpjcyLH1CGs6FXM1b/5NYWSbqMAj/Tbkq3AVawp4Wzp2Mm0eWLP0
KDzApAhGEkyE9U3AmG/qEvMHu1rcyYCR37sf3OkLb2wwBbTCwf5cEMAzeOfiJ2cr
fY9iGUQqLpjtRf9gwp0CJNsGIo/jUs3bcWynJxnLl8lMM/O6EH83t7TJpnkkigj8
GDNG2RY9FABwSFd53s93rwLnlQtlxp56chA9N/MT6DWzvRNZLESgJ9nhDSfcmhaw
lEg+t4+wx+ijxloQIP5QIoCd3whR+FXEPGj+o85oCMkfFISkrS+u3e8UkqBltWCl
RaL9AG635xYfqLeTWd3FXCUjRtbYLZ2NsrOGWRO2Pm6KN87lHNDUSmWkiqDIv9LB
Kr0WImJCByFaQwF1KJi7zkXxVfjUc/HYG1yMJjr1NjCaWyYw94BiLYEXY1mp0NY8
Kyd3MBtpFS+ijUMX6a7gm7vtfzWgB/BVLdOaLt2PSQD88nNabbP2SktcaNIqsvSv
1490ryUM1bPGm73sAU0zlumMjiRgyn/Oe+tRuxcdDPABsTt8FzmiuXpiBgbi5u8x
784fyU6t/aOkgfpwKN6Wl/E5RQ4Zjx78fJz/nJK1uFhoXkbJ6DrIWpXdRx8t2Ch6
MRpKflBWQ70AYdNgnIoMbed1SF+idc8UH8AeSJfUweZB6qCp6LbScE/REEfg3ZGA
Omuc8XaI1I7QB0mgxlQjMqsZ7hbM+xMQW4SzNIjyro4MMnRNaPDBpYuQiiO2GDlF
ECq5z9lGY4r82Ggdaw/S5nAX7syhfXxWyLv90Mlke+B3vWfe+3TKIjn+8f1gpke3
bEbEVEnq/vwF/Ow7MrRMytu2lGiO4G0ydZozMObmceeQG5G2bKrdyefZjtkRJwL5
LN+xajTm3Xrzfg5S8tfrf7GcuoKMYBaYFkLLLyj4hHGZsDrufl4tkOQchkkYPw+w
BLwuOpbFnGBcCIYnNI1kdZ0xxvKez+1tRhkBq2X6SJicXk7hoHowV2te5uTvwQKr
47lx1QjvHijUDKhB2rpOlVMw5b0cjytYuRng9jtO0CDR1pkbzaHelo5MuMzFQzan
vfCEnjrRMXtUumkijtBj4OkG8F5QEAeYooWDcZ45is04FbiDP7P5cOyKl1vUmFrb
7Sy3B6AqnWEJKG21lKE9sPm49PqYJQnbXmunfhB6nD9I8YxGChNnSOVZhf2OKb2y
+RvsO0kHfljNe9wqRBii0xHBwQOYcGskLPNHaPRlJv7scXWQtTeozwszBpuT/C3o
6IDSOrc1USp6cAwF7FIOEhUYmuQ+1/7hvxphmfkpzYYelWaRK9LamIXMAE0bktEY
yOgigSNFqxMny42oftuCE5MQ4VptFTtrE5yYRNksgujHijRDvaJWXVH4ZlEZBTAh
dEX/Ae8lpd3XT5RmvxX6Fbo3p+uyiHF3nAxUqGzcPMo8dnYcGCNPuaLkYaE9J8wa
pDaLkgn7x445zL9sH0vt0XHNlTqsbonNBVXnwhnAL/mTp9psnAdt4nIJewUaCsC2
BskzHmakWyXHg5OIm8ZFZQgq+HGIAW2UKbO6MMThDAnPRClHyOV9ADeYeMaFYwqe
KsEs8t85dwknov8becua1w==
`protect END_PROTECTED
