`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44xefkE8iVlsUkjPqNKDYNb//L8y5MkxKnOm8mGX68XOO6je6SvCz6I5rFaRmFqs
5WpyCTT1c4kWMVRyx959NmSZPsz2Ue0HTgtMoxLdoygI2e3msO3fjodxEOmq/Quo
UG91X21wL7BNYoZD0gnlLkEc7qU/TDpuEs0pyy1FFE9XUql/Nh3jsD5g+CgS/EdR
o5Hn8HvPokRZnsv7nBB/QYjaKKHcWkDomCCZhYL2erW6no1mfbkuHA2opK26/zDp
nS0PM/O2hxdB/FIHHb8hkblEQQ7hdoiczwzny7FV1fBpK2I+zzxdj8Dk+u/hLlC7
N0ZKMPja5ZsfWFiKhH0vRZBS3lvLc34vaGMqHBjvG9rpTvtlNcUpdDV3V0o5J7aH
WOWlHX1t7ubeSUMaua+yVLXaHJFeX44Zojbf21qckaXDz3zT5AuILnXWGtk3HQUr
xPcVMYPNplokxLCAoSZ0hhCPyOPlpT4aaZnTE+d94RdebTW0GkbqsuCAYmLwz+dc
Xah3YxMJmtYkQfK4/YUEuoVJqprd+SjDP5o4vcFXF78QAE9Zjw41/SWlJP3fdgJr
qjnPoPJZ9Qy4DqGd2CzQlymg4Jngmv5LwF09zaM81NUEk4si0xS/MK8xC5UW0WWk
0o0ROy1/tLvMEmRtrKDjzS58SHfu2H8nzUVjgdVrQuSdUin18TOvdyL1xt/2QOGk
iOfY4cM2rbhSlnH4YlxQTfx3UqZSx/SRA4p//A7HyIPFp2PJYOMecHKDgoDz8PrM
thV8oNbAMe0Q+uUenaxShK8wP5Iz3d+vrzHGMRMJ+B2DaXBDFbD/Ty7fCipm7jv2
5H6cWgLcAPvnawtaz3E5nrVhRxa/HOaX0NmOaU2LPQCq9yfrqelWDK089+Y9FaoT
HWRS6bpreaiPILTZX0qjJJO+PlFYHAe7DBNj0LwZS0MSp29DT2cj7Q1+Jjuv5BDH
F8NcPlaIuotFJAs7w8QnpzdCq1NiZppoaovDL9TvIYR2i4qXMiPjqz0wPuhAOOFR
E50kVzkYpDDFJ3Z6jHu+LWZOaXxspRmd/T3qVcSOzQptP2MRhIZTKDUILNfKa3pb
6NWoXlOlJm3GTQ80Ntdc+vIe7/M8kcFV4XCYV8FRoMfoB2ch9mzMXmIMPm6rn6wx
BKlSTsShWe8xp1CEzE6pWnbBaQDUNuMT+HP9gwVEfuS2d/SD9I7bIcDUykIYZ695
feONlmqUAvgdHq0XiBoGjDJcj8qJMqy2A+ElAYfa39IhyrnwUG2nmuI8K2r0HU7m
43xjTyUzvmG5qWUJV4pRArpECYDFtEVfeoDr3ZdaXBGfAHAlmTOFhbCvkyfPDcCw
NkzgUByoGfB/5wG7zL+C72QVPWI0k5NFzasnz7GWeh9M7hgzCzQXudbmalspkQf5
SqBc8/HC8e+oarKWFaPxZ8bUHG4wnt8mdtL3zK8gk10fRMTv3OldVEVQa464LO2F
6t/4nOJRDd6ryJiAw6SNLgosCGmhKfmIy5MHrnRMTeWk4CkmSqQmb/A6PV+3uIfg
Rknr2PoegV7ENqEcZHJZO7NtzIKZI67Az3PybfUBTN+S3RswVUqD1cE0xw8NKhBN
sCp1BMQ8exqngrcyMG7jEubEYTFJ064mn1V/ZFGbLCjoQBTS+w/HnMe9MXG7/5aw
B3nC+FZZVhigkSsDdxEIEPTtz/WS5RlL7cGGnvcaRyLk/89R4QCpRKATGTE5i1WJ
bLHxInQ00hWGuqlWFIR3oQuxvfDLLtBXyktPT7T+6gGUIW9PKVR3+IZRyzXUSa+2
redPjMJYZf88okk5lhP1Tg22PIzjac8Z8kTMM5gx9Za1k2zz0GsNLw8I7+XqOtCX
Lm/379Wen4KeTKFcug5eeyAdBkA6WSW/Lu1Oyh+1Z5HCjs0nlhuhRr2lI5vR6p5T
fbgRi7jF96v8z94XAULu5C7IJ/dn+PqYBk/rUUG3x3WscrFWOR5/VvQVLvlurL6V
M05DIlJXEncTHwqKnCFm6LbtAfAUUocrROosNbcoxqbwsCGE0xf+FMVJ7ojGSlSf
rGpHOEGHmXzF0oniO5Vpd1MErRRyybvNluKs8b0wrgQ2cgfGMuXTXBxS06k8g8fz
P91FcOVzLsmDqhwvuwdMZiG5J86JmAtKJE1Dl/+VQLxqOdioXYzbpNapQx3853Vx
0QY9LfTTqllFutDJQGzRxUJFrRmp8rWvVKPYIrCLt1ndOsldWxGXEQCEtOVkPKus
guGxcokg1ZHGhrPSVEF2cyREvhDJvVyaNTK8XGotmDaH0wuIJViaV7O2TQgd9Agp
fKHwM7QjXs8F3UyKQNn3WhjgGc72V0Xz30OzKNAUIVb2E8bw5jNbyCArs793BnV9
/ipkZTaOuEkZE+7jagT0BIX9O4lNkkg4XU+F9Sy7l/zMMLZZ6Vw5QDnFtr9INBu5
cCJqM/RBx5akuqamrBxNUuSOKAzpWVsrCGctYB8pftPZ6gQNGxTslWM2JzNNcy03
/8LQkCX+StgNo0AnKZwos08dNCbqkJKrbuvFnnFbiKG4GPcee9U7EhDctFxFhpxH
m74UV7ECAC1xDiIAhsa9GK2Po937WvDYbBP6YwHpgo46LFsEnfkVI4Z6qncXwCcE
adSXvlgaAtQQoqv/uTFKqb3SWfoHdEwyeh5pHX81MbCw4a0H+uvRGW1hjcK72gry
6QQ6hGOnXfl9/ATrEDS4+sxVZywN5CP5iYPBi1RQlhDnMtgzlKO32Lp0auqjl9H+
CbNBg72B2T6AJpA9fPiIZNmI4VN7Khd37R1xtZPI/MSDcsaU4BCuZIXNxBcoHqsS
PbJQ25EbkZOmCZwOKWvpU1BDfBh4ggpr+Wm0Atq4ZQoV+aGoLtX80cBD/5FDe4aY
W61JxGn40hjRgStGX2jqxFWoWDJ9C2pv0wAe3n3w1gzrEmg7LmPyTi8GLt5sfSbm
YcsRR3O1MCq7MHDSnQG/PRL2myDYRuIWACz7x14ZAKerkZ0MGfgtRDN/dAnYpQnW
h4Y6m3eRiJKqZ0j2nQtpX9E1xAHnLWFLUSIvSxQ474u+RYldyuzm9nZYamYrmYiO
B3R9EguoTyeQCW+w5T7fWxFUuT12Ud0wJFwhAPkPA5BBDNLvewrTxN9N2mEoAv4t
sAS7VfPG/725v4Fqn+B+UNM9f89/i7SDDppDNYndEn9MrwmoV/xd3MiZO0fA53FM
CExn/9sY6OypHES9gezUPlGzStOQLxXfXNMRCwU96YcE8MnEPdlW1me5GRXG1epK
la+/LmZiwTeWCdUJ2oLVv6XpJAEeI4kNHUBYAexVYooVPWdHnT2PShVEQtiSP0p4
UYZFfcVCbQCWUgS1fnOy6gvmEVF85OrCPDYVRddw4FX6EArlt+ufpQQALR1QM+6N
qxh1ahmQIsi8GZ7CJu66+GyKj+Ka25sNvurPpmR97cbAjpTk0eE3HRTXsCgkf58p
1MYnXNgR9jJcduuL1G4+gEw0/9QGzFicZzx/pQLQQMGR7/L+LHGSh/zOar3M7fC1
MbKVdbJtVb1vqfo2YxzYPZn0n0OTayARTS5L+qZ/IkJKY+fYnpEN6Dn0y6wRW2hi
TYjpiwMKRHNzXFW85WEqrPG2/uVAz2g6Df6utESWSVHOBw3qSzq/+MEWJF/RkkMd
aNtgIhrf2XcyDxGimo3Tazo6CdGJC7T5o7M8lTgFZEZOiJzQZwS6GOJghs6cwqdc
wngNadgZ2KSPbVijSKh4AmLR3DN1cI1wP8+7vO/01IKnZb9EhmPAt3Nx7YtuoiIA
R9bs9KbodaCiGu6WJUSX3kTGhhl/sM2AqBJjktLhSvwc8/cHbDr5Hzk19RFGt8jQ
rLGglZrKrT2ck1iaMGivntaeqVR5Ym1/qohQiADQ2MhEpw1uaYmArbqUBRebsGrx
/jM45iNK4Wm3igvnMtl4AS9vPJy5Nch/h3ui+omz7mtDixyfF2g1rpEWxtIK4PDp
1gvAnAHGPqVwKu4KpEtQ+lNFu7ECFZ9iyF4r9Cnx4GVuEMfp82W0P1kr9P576qAb
9mugmUBcWUwV4iMj8QbvJJbWfkP2F9QtyMSIxuqx/bZzGXxqY3XVmEGKBJVKy1pV
BJM4Q5FwEaKc3z4M2NNd2g==
`protect END_PROTECTED
