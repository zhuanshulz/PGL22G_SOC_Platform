`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYvP2mc1l4+vtLTmiMLBCjZabWZ7PtJwKJ+HlkfFXA82vTjSZONVLItkCMs7LU3t
9O+9aMtduBRvTt4ib9b9epOj/Zw5Q9laSxwSJWeSQZqq9fg2HLNLSxRwUa9gIMjn
FLWQR6W8fyHNDkbzrPXUxRgsHtwK0Hu4CqRCw1pLI3/syeQG7DueT7V5vFbVWiTJ
0tcRI1gEwvkA/X09XOh/FaVTgukel4VbCyHfHwNIRJ1/b5q6vCCtv9pwL6Age5Vf
GMG5/YlGvOkBjunfhFbhB7KUFHN3CV5MCUMoXsgnMH7j8TVkY1sKAsMwv8GCjBrl
beigTaWWQItq6TJDQBhW0PplSfyvlVJ6BDW6zTZX6auI2eUi0v9GSGP+lUj80dBR
wOqf2SfWACs28sjkLCm3zqNMFJUcgP21j1ADfr79SWoeBuAiwVSsMYVgHEkoNzt+
+Q49Xy5a6i5M3s9wwVzAKL0H8x9BdeCmYyc9vIGqxeP82V7IqDls2yfSH1vPgCos
IuGjsQgvnu9a3WIsesl7o01JBhh4B6ynI0Tz7otpujlLaDIrAMKlxp5ZWGBwR/OK
bve7OZINrE7GQXqlSD3LEhLXb0yDmItWIB7iHt860dxIsf0Ofmdsjo5Ct/8N9EtW
wV0+Igyo5ot7RL1yEVL6NE8IYqke62b6XPgfvcCWUGZ9qlKgT+C5jbEuY4CmXvra
Z+m4IrxRfYgzmn0SSH35qlLHg2U9Gz46pICyIzdBnOV/eJUjFabYTSwlhttnVr18
`protect END_PROTECTED
