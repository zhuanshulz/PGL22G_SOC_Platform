`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
162vIiCIvleJ23kKyEp7qGsug0Wg50Z3/uEK9Th+G+EVazg10739XoDSzs8ak8Xf
t1L/004RZ6HeT21pmxqen7c7FE1NZQaeVdchUBvKMsCPbEscxFKY53O9t9q1LBNP
E64Cop5AHvQARyNc2feTcOEfn1foV5tk1LbX2BnP6oieKQtEMwBUexbXq8SfJIOh
nSa6YYihHhEadbJ2ltgqbvp+dRhk7FRXSArFN51TKARWbbPH6nuCDg7ZQbh51OIr
QKtCN8VqswgP8R3Sw8P+hx+84HCkQI9Qk1AaRxBrEl8=
`protect END_PROTECTED
