`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hO+gbrJD49rzokNgtjYiv863u1/yJ8AXn/Uj3mKiFTJdaJztJtGC+zXoe0boitsP
k6IRsFdkcZpO6n6yNjhExazyJpK5irKrzyAi3v4xTs/HaynBeZaAw0RD/cvJiO7w
VdBWFnO2lb05IjSYNDBTNxpcs+tA2H30btzB/r4nBj43yx9sAMKDHcgq1z0K+nyr
LFJ9WpKOcDigVaiI9oai5dnlpAjVQC8JfSB12qECLEeYZ1vbj7a2qjhYIPL4UUeE
f5edPcfbgl4aWUo7GwcwyPL/DG52y76ULxhx5q3E0WJk02kqDdVHt5wA5J0B8g5X
+Tiz1+pwfE6bxKzsqQIToNX8AdBjti7KWECTqBylUDsITe8wCaEvSB4dIGI1zWdc
wyDY8h6ajeoteyokSFv+nYQq2am2SxUyWZP100XM25PgqG9RvMC4gdS3ltfuRux2
OrvfKz0kjhzKwTY2OtTx05AoOh6epgWn9MJ2+KdMei6xUxtFIlxR8HFrXl0RPKwi
reg6pfMzVgXvIHhn0xlok3n5PWjEVGkzUG+vjihZYVwRc4G/x3XiSc7W1rfXqK1I
jKT6D+jEmzdsm+2htl1HF9te5sHSxwWl8tyxw6t6RKS5pmkeFA+bWgDFzlq+cddX
p/fnF7rNNdhFhW015Ei6rTCWGm2FUd6FNio52ytfMk6nf4jWQKDDZ5gj0fBXSqw2
oVjsVPexYe99IIKwIkA2pLVSuQS6mXfPKlfnN8NBkAoPkUNTuq3/Vd2Iq0chl8sK
ISQrwcb0NyHGarPtTrh/GDaSZWK/OhPJ+brqLM92ovJ9NSdhGUZEEVZothJnk8ff
R4O7qxpx9F5RoBymgLIhjWIcywvt1vhMN7M58X56JBGweGS84EHbUM+DdYW7lL3u
1UBjzhilK4HvN+cbGViRUSYzKuFQYDoH0zjpG4r1xBtuHaf25dtSjwUxgqBD09RO
ii2Ati+J3PTgoUJ308DWDXqEZWiPkqKQ7H8lfy85cbxFQHSbaZLnUx5QSP7eaOBF
WzqeCExDASe411D6qmC1E4ZUIfB7IlbuOIF59asbX7tHyHm9OndylIY7Cir5N0Sa
W/uFqXBlrEzHTyWXI7FU9RxwG0ViWBIu3ukN4RyTVUZ9ACtbphlaaQEHoZUm8qyz
hXbUFEr5FslDinNGtlrqM4qQLJJSsLKQz8Djc3sIXkdunoOJ+aS4wX1U5BfZJm87
ZLIAi1Mrwdr21nGrBMp3e3EwyEA7edhXYbW1aWI6oiAfwQ29RAixCRP+J1FjzJ7S
ZzGxKBwB3/sxjLxib9RhDhVy7oca/gpbE+XYlRJoN0W/HTbiu4SCvApd3RGD+AxB
RQHezAfLKXdiXUBskPsGPm8WSrDA1S4LE8NnG9u1vse0lcQGIYfuf0C7dwTKxVXK
0ah1gyOxeioFsJq2pBmEpg/ZP9OUlEry7D3F6pUi0eAouMGaVkQtX0QrK2aRVKJX
8GcuaB1DSgaKDyfP9ANk89cH+3D0JaShIIxTduKVSGko+LZQBjaSWeo8JOWP1ac0
yBIiSe9Fg6Q+ZdUDLH9XSM9/P3eo1U8tX1yUqvD5EJFuf7EEwL3REOmVCaCzORZE
0AJFIG4fmiBM5Z9g0ixym9C8SnXkTGi52VHZGf5S2945kXLEZgST32NminNWZTak
cq/DYUPfSbJ7U8wZO0tXXZxFOTKgjAGooEAkXk0vT6HHX7io0ynHBjpmP6EbJFZY
3fuEXmw8qkKe3idVAkswjhXrGjDokleIPZBIZN7PY+aXQtPkQqunFavZU5PtdD0Z
8POOws8ITohZqzi467qIBvREWkyMi/QiD0WZ+79+jXgnzyZVVE2ikqzsPq9kMyNF
IQqp23+KWYyjAaLCb0/fIms/a7/sN+s6kQdtLdF5HTcD1GaqvgyuWjbaqjSa09Hv
VO7pVm9Y9OcMdtOR8m3+DLJc5HqwKZUfT6EnHvip5kXIDjnhNyyjLdrBB8uMY04Q
DHXlwpSglGz8b599dEDxaZkScy7cZc4I5W/0bkA4d/33y1yZcw6+mHEBDMFlKECs
5GSTZ5ln4ckONfqmUKv3RMSTlf6DUrvFCTnAQI8LqkS1wP+FnWtONOBaohpjX7dg
A+Beqnv2iRDkPoi1mbi9hrjxszF2/OtPoh9k2KLeqS1wqLm/qNlGgUveL3p5xrVY
64vFao+6eZh0+68dpNWhMo1N+EFs0wVJng5C2E4fkSqcXUy/Wwv4nvUAuHE9XOl6
t/4p01EEHHklKQ1D30zljRgx39Z+eOTD/3YEFNQ0ycQjdW/rEJ4//rg5x/Tpxtrk
LzU0Ojq2cmWk1MUQ+BY5BEhuxTYSgoFaPBkxJzkPa6+qTrbH64rIzGZXh+2Uh+l7
GMTEuCdCmkBM+e0Rarp8+zLM08xOLfTdblvP2FTDsjP57OnYjzbYU5iPZ1UdlJf9
XD3FBFX6vYyXmsxE3e+ewgoS8sQ1x2Uz1mDDNEQV2IfZ5/jHLhFmXGP63b+HMtln
zM582/yRnaxFq5uXyCt3X0BgceLn6WTrTUT4Fnw1oTm+pp+0WRMP/VMAgUwhPXQg
fazMc/fWxnE1de4M6PCU3w==
`protect END_PROTECTED
