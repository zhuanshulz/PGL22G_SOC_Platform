`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBpKuefxdzq5q65PmVbUEhwy1nBj5YzM5tN5L5rAZu9ddvKlM1pWNNucnL+8ZFMq
p5XsNS+R8COMWnPo6rxX8KOhtW1iAeKC1QUvTKBlkUB2mFtQMg4wiIRu1t2NSefw
9Uau1QSXogJ43NL3NkOaHzf0xsCYr0VjL/DWO7X/iEx0vrlUCCRa2+J+csaSUREB
F1dXMT0wG5QDD2gJzBMl9YIihESfcMk633i0tCAhiLapj5y8NyPlMEyW8mdj+4jm
Ioy6xn+6oKiR+zVHN7nI7lZEf99J9Ca9W5dHBtgFsBh1UnP5QmUI6Pa4DtmR245O
eChCvQWVZG84ZvD3tHph8q3lDJfO9Wp778IyFaDnJhHcsXkYI8xVeQT95c4l1M8D
RsbtkdJFDHwb1wa6pBnLt3YZUQ27Q0qfzANVo8bG8K94Hi3cjpz7RnJxT8Q13WTZ
8Fn8iD5HGkpEcWmRHuYEvmqASNvSV4igeAFVJ5G+p9bgot9SSPNf4IBvxzTDqC8D
fk57HrDg8m8OuTKyCyH0FVEkLlqeJHQYmmMwrqOVi928GCaLbx3zgTDoM5SMKRKV
aEDi3j5Dy58ALVwYNEYPOBSh63BpDRYAlcmLJFQabBQV2KWRtmDpSs2X1H3t4nkk
j+G13wCEsUYNmzw7+9MkwbAzyzePYVHqWJXDfTYm1j2MJx05lYp0CueiUznVDZZj
8NjgndOX0h/VKx9B0kq5S0sDWxBm+SkYGhj7k7kduSSOQJ19vSs3SZ6n0EO1w9jQ
i2XOKD1XSrGWXnnYp16UR5EVp/LoS3/MiLLnibYrJYlV01cHHJS59EZhjmtZPRBN
AARNPgRDkMIGmkP4+au9t6GbneRuoNII2v2FchzvMdhOn2/f9xUkjEhOXiINrGlh
qnD+3gopeMHDfzQFwjsUE6gNX+N+jpMQvPcqllczFZHwnMe97/YXacW+aq7HPCiI
qbCXqUP6K8yMfR75weaahqGeTH4/yVWSGLPrJ/H8hmYXMenKmvyo9yiYJmq+XeWT
HRRM+J4y8gm1xKz0phtx/+VdZK0Xl9o3HbHBzV3FSHmGqkhHLvrydFE8k81nGc/w
b9+bZMQ469W7VsBbLOjMzcXxpyaQAvHAQ+ilXp4K8ks6CD8HrF55ovDZyywacU6k
8xXGbTxwgXfNcIOI6J+9Zf3eXikZoct0+cj6HBd8uMxa4yJ5wZDvesPRZZaJohi/
5SlK2CHwffouhFQ0WDgYaACi6g8EBuTItbjEmq3NqsnUCe//B4VB8yRfltWJ5PS3
lQGsk07V3o1eDjjDYgKaIXe1wjBMQzGID1IamcXeodGz3xxbiCo38xidRhQiLDHr
86aoHciSAf4rGkwcvy7d/LoZQsS0yBMiTpp+KR6LqRtVxxMHdKKfsAqWPrrxwKj/
zkgY37pXdvDEiHsSyCmzxZm85axnQxU16lMXqiHBnO6G0AuyL9I+ICsSjHrV4VDb
2hMOA1yrzQDZgtqVuv3ei8AMcnwXbtEfmeqXQ/1hk4zQXisSTb65gQT80KXuLcL4
I+/3Ep07/UdIhTwF/B/LtcpnwxgfZMtKByBTS+cPVW3zUNR0b+8+Y3bKYyrFB8AL
ngk1Wl/ihnrouePoNPMe5NRgF3X1SSEnom2ezCFdWAdwzN5jSive1knTiQ2HuLM5
sCxTcmSzTrQyKLt2Q6VMkRQ4ki2nGrEwZ1AI8qbUd8xmpQJgPFKlADDHWCoDbDM2
`protect END_PROTECTED
