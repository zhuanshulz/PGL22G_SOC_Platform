`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX8f3a1CaU+9ZuRsAHK5BTl8iKZWz2HASLAgnAmYzi3ENp9Voxzfb+lktZSFAcUq
hRvza+SexVzpVrOFgYPayGREq/2ygonYRSsoh1VWpiNyffJcbG0d8cxnjc1ie8jP
H5aTQLCfRbHkoZvQ5IA6GKtaEDpLg55bTqGmM7vBJh25MLGeCuc/KWPGmc47qb5o
rIWtdTTOgrGe+//n0BQ3TWUZ9ZdgnYmkSj+rE/v0RyzWC6b89Yhk81PWwRpl+pFe
vVjZ5P1CB3LGx6c4yo1/JzaEHtHPbZtZrkq8ZTS+RWfswUaQL+afhSMbGAFwJBmy
DCH3xdvXD4idRxf80JhHpf+X6w9e6FOmazrvoEsK5ZBcHbkI/7TUh9OyVMbFkCrT
F9vCcOgyV87OiFB3iZ/z1SiJJGD3l0/ylfymEy3wtvU+qawRox1Ky4aRUECYS9TT
35Q3Lcp83AigYNflNnuC3H2zbB3tWGP5+8Jv5n0sDWxbP/s35BbDTRJtho/607zL
boaz0pZsq1nyI1/49CJ3ktRwN9vLiLGoYzb8+7vHdtuTjThxb5Lh/COqW8QVoOWf
Onesrza3lxEs/4TA0B7FDDt11lkx9aALMVTUscG2rOhJondwny71P7tGdCCGhiRF
zNkePUqJaKgpdBDYlwKOdg==
`protect END_PROTECTED
