`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KidfcV4iMYbtoU9sjDdLtlwu5z4gPY6TmcSAUEwgzzsbRHgoCpyv1nttgBLotQge
Dou6rDQg5nwFEe+zTF2F5PnlO+Klj4GzV3CAEjN753Hjya1Y/9cLfcHp6DcZvPtC
Lo8nMS8Dblb/5wqurWZJx5oRG4/hO43PC2Gn3aw6wgDHq3CcOQfu/UBNyCxr0mHV
ePd+7GHEbeyQk3oN7V9TQNiYUGKxOLZ664iBPyFBR0lfOL5FDeKBRqrhro3UErvr
j4vrUawAGxlGqr+Xs1pD1Gu+U/GzZtrFidCW4VLffrCWY4BbFnNMWHhNi/Scgusy
mHbtsdg9Mwp7j9+ScXfDDp+C5zf8Izi8ZVvHq8nGJymWIOi6orduGn+5eq2ryX5J
TWotGPA0b6f4cfaC9UQC+hRqgFXVEcScIlcRcNG+dXHBKgWi5icHFwVIvbcje2JF
u0lbMzKpwFcjPZI4eZEbLzRyItvo5UuTkv1WVWryifsYF9KABCV9EI8iRLoGvafA
Ix5huOrACWyYLP/G85aI3tsCGhmVKKBXI3sWEUaUxJVXjLQkK2ZOytkeEu5R1TUc
lPpiCenp4wKMJmTrpklyNUyapYkZyGJvFNPZElavYIXMjiCy23k6i6OCUGYk/UYH
/ktMwoJs3qJtlDansxXghQBMIO5CeSJUJl3AmYc8I3ltmGu/jK8mpNtc7bYE/fLH
vWIPRq/6h5+Z/XsTPTR1LkOTuJnYjvxSbWGXe5d/eZdjG1pWekTNP7/LbKO230GG
/wfjCBl5NwNiQ9IaGT1IXxiXM3N6Yc4+LPdMyZc+zS089lVtlnkFvBoOV9/RrHQF
PPWtMX8NBTzJ2q5Kns1OGaZ4pYznapnjSmcvo4Hlf5cH+uMlL05zSceFhn3lFcCG
wjsgMl8i6kI0bUAribcNrFmduEULx4Rb11x046NGcHALACtmZVfSyoMtDPKu5ABp
rhkbqbWDZYbaR/WOhNH4F/AtMf+06IS1UtPr/arkVGEM/5VDRMw3YA6DVaMkuCwG
IA3kCsyiuoX7JgRK0/VyrL75eLAP7sLE1uqenwNnCEJLnWmOt1vF66EYB6veZdRG
AcfKFFvX2UGxXMV6plJswk14ShDmaDq6WVPiF+VHIm9+zn38MZPPSy368LGLx3Zz
/p6Wfw4wPeLjVUBZMZXGGNq1wQwAo5KiCNif2KiiZYrpzDXog1sXi63z0DX0ItQx
70PS8BeE3io1/pIPZ/Sc6dvif2+srTQ+YAbQ2GXdomcY6iu3BeHwd4D6AVAZdFrF
nkriLe/vrl3GpbbQ/0Co+0A1XFKOqQf21+NZ4aUy4hB32vM6QUs8KvxO2gavFrRX
GDxmuF4PLpB4ht29uE1J3B7mR1u7iNxgJ1fZ5N1HH/d8kHCYlfccorI9HBvS313l
pdz9rKpkVgXC6tFNbVUI6Ov5wiG01av9Gam0c4QvkzNq4LqP6G1+krKVjWPK1t46
fTzQCjyio+8brLqZlB408oB3yMAhxD4MZEFoji1ISRZ4FV/9+anCvy/Eujqb4Hkf
g8R70P+0l9r/S5jo7g5mpTRplzgimTNWR9No+st2wNE=
`protect END_PROTECTED
