`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zl1Cvgv+jmi/ajctq7dYXtRqZ56HLtahpHqrdzdve3PzR60nOofaGLz5YjR2yZ9c
D/To5cAz9K4jIlRWcxE8Wy48qXuUGPFKoNraw6pqhtqz8+Cd7dVnDWnPaocoJ+f0
WvzP8k0QAfz52WrNuzXAQJM9HgWJpfRh2NAlc/S/TbYMKODe0tjmPrKqqO2j58XX
sHHD6iKY/v8cwQmlwT57BAVUIFfOO7fEDdzH7vbvtLonK1sQ4OFun/a/ygsK9c4s
jyHUN6IWOyRZnPRYVQVgt/K+jVxgGZ1Iv9dicOHvGvohCIYRfuqra7idAWfsCoy8
x5G1l+1YBI0ZEQmJS1reyoGu7ZChBakxGZJfdULO4fo/HZK0/ufrKn6TW0k9AQrk
3GicK2B50JVICl5xX/Q7JlvZHQHV5Ide7X/U0c9PFcei0gpNO3rojaLXV5L5/L5i
765qBkxlPxo+/NOOgGF++dJjpMQ7geM4VLAObfiayZoH6iac/cUMW0vppUspPymz
6LJ/7mSh8tPDuchtFPYppvtjYwOF/sugF3nsxRRwwWWMX2sjsKWqxfNLMGjPIy6V
MvR5WoAF0JlGGuaVN6Nf1kHxbFrG0v9mJZcGcL48B1gjJ0yCMH1aQkffU8NfK0uW
lqtxSFMQSJmUmvb25eppJDuJIIHwbge8Nu8r1hfiHXpByebVYy5Dj/R75C2RUAGT
XpIWFKMQzEMHInD98zt3tR6EDDX5nh+SjtnHC3PaaIgyPvU+Nt1S9yIvEDmSndPV
JA7WDXquaBNmMrAAN04z8fhhakFGB4MMXhiDPPdAeeCknxEhhpiEOjzHQrcDOYY/
IigwLOCMZf5yqmncHaLZvtc1OZXrtHo8SUbXHPgNCUzd4yZqXtyw3onQGTxUYPJd
oRQaKbTWTdqNLRpHm/s6Gbjx52Pa5v4QPZxc08Ss3kNMl7PsdF8RdD47itOeMJIK
ZAbW1vD9BCwF+rNszIZMDAPiDMOoKdVt4DfpIQNLxFW+XThAmL2sNR7snq+gHz5b
ukauOPEBo4MRljTl1Oy689FP4Tfank5TqejP5xeVSRQqAVsCRJlO1xn5sxFzcLKd
TtdOYpETga0VKIXXV7yDrbeYYBgMNWIL6cp4wGZEtgyqn+2n6MzW+Zd1M51Tr4JZ
+dPGSPq9mligCS08Jju6rHYKdyOra9RCb/pM7lFh+L8=
`protect END_PROTECTED
