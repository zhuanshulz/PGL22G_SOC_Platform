`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0jh7cGpfGnu+4ASO0gLO6ZMu+AfpQWmOdddrzoJQefHpCBIKHuHzLIgathsz3K7K
hDRvdvPJZOcFVdcb1FajdwKojki8dFTNt07t7biZtvxbRmYnASngRMH/NqGHMY49
c2eBticidO0/ZBHUl5SGg5RWT+AJZoSm2ndKWXALTrB2nt1uHo65OW6P7oWC9MWp
JohudkLsMz7NAvyiXKWDEnjoBlIW53WtQNHxs1V6NFt4uNKhZLnTSaizP7XT561U
fDboqzooXxv1aMB4sQCw7/obgETR5yzLlqukw9qWmIuODK8TWUXhezoWC62YImhR
ZCWKDNvv+c0QqkqeiKN2Y39/TvOYmNTvkFWnn9gEQa+fw166YmenwRMa8wHvOMIK
K29DG4U4++LuSw3VpIBNPwKHZipjN52ZMxMpXuiZbMHCjYiZr3wZrF86wPLs+mgZ
KOd83GwcZ97Q+dqPJu/lKlIg8LUlEuJyVHmah0lwUPv0qZgmPutiM9KuwsLWg36M
9AyuTx54DzdxC92ZNL12jcH3ner16QNwtAdN0HTtsns=
`protect END_PROTECTED
