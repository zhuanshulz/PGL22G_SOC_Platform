`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMrNFTqcSsc1nELb57KYvGwDQ+bh0bPHLHt7MOnkfBeAXxd7jfHpBvA2j9F5arOa
nlNjECUXgOAhBPvJ7LBPO9OYcX4fRM9TWnAmJv/7SU+xOkKVRL6JfWdxo4iGcD2v
rYDPC9tAFkm724sd9y+TKccRmIXwOjQUxKLHg3IXJUFRe8HucAssj7Dl9vh4oll4
WhxjxgMxDg2pAiwMl01g15lrel3XehbjyTQTvpcjX01NWgjoMkM8G8DXQc9scEUz
FRJHrqZN/aelNhm8pTVdB/cxcIaJzJWCeIrUfRqkZ0KnDPTagT10ntzzEXIUWPzf
l1Z0HYlQA5IdR9tLaRNgJqaj/K27Ks1ZzP3a1Pwf+JRxHbvzWbrtHVduPQf1gOlR
mUgxXKANh80U1uFoUag0L2tvbRTNxD1UEbAfZKVqF7nyNZgND7uUweRyVaq34I/7
BmGQLq4P5Bm7BvG0SwqhS4t3wAa4EWiz+8or6i/Ctr2KcHmDAI+XPYeNrbhqBm7g
odBYwcm4zN4/ozpcU3IDBdoF+MqLZhf7q9he/NtoBvmFhjjuR94v6gHtPVnA31io
1Xwobd277VBE0/WOlrYHiZgBZzW1tcW84x/AtZ3cMoH24hB3kOlYizJJak2eQkUO
iBuYVfgHpjya8rvGVmL5Fu8GcvSzieiz5aqheVMNc0IRH/q7I0Hko16GHBSWCzLM
la61sfq33WnFaGrfXCt3DsDvoX8dKSiYQb+oG0/CzWVQTUKYGOPNbs7UOIz+XF4d
LcGz+5+2oYjyZZqptWYzfjZs9c+Gx7gF4Ywf08Cg463eW8eBqw8WXvwXY9a6kwWn
hlJXrsJgNW49/+GuleWF15hex7bjnWg9HGsQI//AxVsYWueIi0n1XQ9eI8pMrOii
VvbLS7cDX78uhwByn1bk7i4iaBfQE2xdU7uQ3MCR1QwhyL4eXf+Stc3l65Kne7Od
abh94UdunN3JcWey/Ioe0FuucgfICM859PEaesN8EAIpfAny65DC08wJ1jfqqseG
uLu6LpL7j4AbKcCnPKq6gxmuBfoXWXjhWLcW/5rRzOh3sYTjVmU5aRu6KFSI2rwC
jlteWDegYInysNCio+JgnIIMRCiuP3H2800hS/yMwQyr06MOjEiYCMs8MuxW7WWc
hHhmTJCIKHegWyw1FQT2kHDYbE+o4ws046OGnVms3v7byTkw1Vnf7kNz1dOvzkck
zXYcRqvDeeffPqMLicghNcKrT16Zp3yKRN+nUI8KuNGqCcSt8nkuFcP07paT3CZZ
nEBZvIDUeUf+0bEZkr3tTgDUfuV16Yn2l0o5f8MNXWaTAWCQJZ1IgKekAAO95jjB
NyvOHjYZgKf8lc8KMSaEIHeVxfzwUw4yMayD2e+Qb9GLk1da9DNCY2Tz7zBMMyYV
uG1Aee0I1aRmVxA//9aJgU8gXmEkwgjvXDv16hcHp8kqoSbDj9H2cnsi4w2JB0S4
B94Ct+UHWbwT/i8PJ0LGZJInrk63lrSZj55TAFXxhRsm1K5Ck7FuEwQuk6TK6nJQ
yG36/Y7adQYLbtXuftlpJP7CmOyHaItwWN43F7YS6baPcUsHX2Yylb4HXQ8vIkuj
6gWoG1xdWnM3bP5si7h5jOLUukYITKkvD1YNuWTqMSewIRiZb4CG2CIFWXbmvpKT
LylQOZpTe+mHxwYWrkDgGW5DdFGMjr4i050SoHPgI0bb/jQgqmiHjv7cf6hiDp9h
UaFFWZJo+pIW9EfI1PMX3BmIk3aovtugbLDjkntN0MfaE8qt0B3AZzosmpcjWICZ
po1bp/AMFKtpeH0pYfrNA09eFRFzVydDanR4x1/YZGSiSsfkB0Ry9F4t55Yj+eCf
LUL69yldKoy8ji/YibjliTZAOxcWzydRz0UY3S8z6qV9uA1G1lq9246aOPYLNnO4
+r7tgzrZbQNoOwUazene7RKIqKBgHcvYujuZGW/hHeLGqyLNtVx3itugRhSzOMkT
c7HpELcxq79kSA6S4pCCXvZf5K3vhUnsFfEsg/NDIqCvs4qUr1yiDlYOWp/C/0r4
frn/uncURLun+d1x+/jQBkBRckUTuh12UelXam/WAoSyItad7MitBbheCOT9Qho/
/eaE3Cz3q9j907roY1eFefJBavcno0/kTkTHYWTsXNu0kOuDrAMDf+zJ7cUXjVlA
PTkCwztiqvBLk3/oljMrQ7vjaUVFpvq9SJ69MPf/WzHwkMfMx7IZVLdI7OA9sMdU
`protect END_PROTECTED
