`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QAXdLp2YQVEBjTO3jSsf4cdtC2lnFRwfauQFkDSvA1sg3Ol7BZDxGX5GNm1NvS1Z
zUlzFYW2m4wcBnIyyAzqO+sious4NReL9NbK/Y9rlEu3LcZtmmQqyKh6xIoQahri
wBYabv4lC8GpTsSBu7E9jRyi8RrW6mWvTF709CJ2Snz0rxI9VVQkvmz/CK3BI+uZ
aO6MLUn6py8tgh1wRhoIQwNe6Yop2hhRCs3t6oEM65ldbgN4sWv5d3lvujS52Wy+
itjZldRZaQivu+CHyqHGft0l767FmmfkVTBNZyGBJDYZJztsI9wC6QEk1C2nLUe7
wC700k1fJo4js791vsnYHFZNx1r0mXp3FZWfMpOqgNwk8QCntzPGDu8NBg2G34++
3V8wFLlfiL2bOWbszSWpnYtfNicmx+R7kenfUv8K4y2p/p/QtJIyNhzz8PdthVSA
YlHYla/8VeewejDWTh9sal+4A6BSflJ6jGv20c7OkO/r22K36FTvV9F7JUGayGZT
1YQEWuPySwFE0NzrMbJFAqaBGJKYKjcJwtywy6U8L2Em/4ZhRgeNLYEBjydDBNY8
x1qEE1AXIJNrEgbGqoGUD/e+TM+wf1iC+xp5ES/lxAcazRS02hx1+BSBHKtkaKi3
vozx4Nk04Ubyl6GN51X6US+PS6lRUbbIWx56FNThHl777U2mW0SxS0WNsMZt354N
m8jbmWtMxMDNMJIijuIpglPLhLMwTH9+chWHVd9zrwin5FuCGD/a5+jjEBzuDkbN
9JxLGA3uCKi+1aPFy5chjok/YcH7JrOXiraSxIBZ/CZ3ZutH4pV8H+rn4K7ysqhN
VMrdRuF03+Mr1wcObiwG8+mbfpbwXv2fltrZ2Ytah0V82h4maAxho7XKeG5E2fvP
Mq1TlARc9RlIx8RbnNrjppN4bhfm0drMYYjebxr4EWQHmpkdEBqs52XpA3tVDbnX
GF83mxtTmqUuXx/U2npiykJR/51mtCcwn1oLajtxVjC3ukcGfGwS8elUcYrc5Alt
B+RdG+l+jBw0CEGFG+iOl1X1AHD7L774cw8pSnKSqvEVeqofOtusbc0LmY2GMQ4k
n/B+ZAzdleInlxSRufPAMfaVZdhgZZg4kQLSI+bflHylE6omc1MAzU/rp2O5x3f3
8jBrJxPBXT/q4jzyg4GUgE3i0m7irjfMOqWtcxOyGK5J6q/M64pd7KLQ36yyuGNJ
uu2zw1mfVE97HjNT+zaxz5up0x1+W87njgcRX8xb57aku+bmc0i7cgh1ubzGAxSV
ycKeeHjaliJviQSVrJvSci0IRTy/rE2CtbEPEQV/iGMN1+NMa5DY0AUIo16Q34JQ
V/jMSvHSWUODcn4PyY4soE7GxJqRcQ4SfxGxCDkeV40/QXHT+tYFz+YOQZnl2IL1
lYQy9faMNkK6/FdlL4AxPRfgRSA/MouDJ7cE4q8UqX/SrnIOOp0kPz8MlFuzApGV
uHN8huYW77A93CbVQ6EO479Y+qXO6BNjn7r2W/8KCveYaQcQj5SxlwTEY7gGn0IC
jge6mf7wRv9Xg/e7Ea1RdjK4LaiYKlJhaqWguuji1MEDNPx9q7daXQkehViCKNvG
Fvt0EMa3UlSChwixi0jEtfWbkHh+jdL9Epk9QueeokNP2pg0kAtv4v/oDiVSWwVi
vLZfqtaTSUH7uqu1YByK47fl5lLL1U043emdEulPRIbVtZ7mALyrK7a7d6DPqaJ9
8gAGm3HJtF4K2zgHD5KHn8bdgPnP65BrjZRdckjJ3c+cpGWd796T0xGiwkSySF+V
UcxDFaZLibYxL+rWjRvEIYXJTOnQdxFgCmmkDaljngknu7LmNICP9HgOWwVIM1BI
f2OuNx6j4TK4I4AcNW0v2sGqyDRjg1JAct++kXDWCm382YqsuMJwHq0sdHEfX7Zi
PwuIG9fGmRUpNKm9OJzd3fmszKtWk4DFx1Vy8BReTRPii2nbW3rjjonVaPXK+3qI
ZkMjTKRR2FRYhh3Yn2pQU0jOAHYAaSDfMKtp9eftHrIqZwokWtLdz66Uc6YEjgLk
Kz0wnvlD+091ShEJUQYRJVrnuiMqCYpalDkkY4u7f12n33fnvGHc9OGvzzm0ZSLp
auuTl+gMDKd4MT5PDgeukkWEJVLJ5rQWUP55WxKUEbTxCJlZzUqkvnhWxwwNm8g8
`protect END_PROTECTED
