`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L7//kkg/KsQH1DVb7LUeRtnQakN0ohuqO7573SCsel9ZOL3gYeLGxQl2Y4Hl54s1
eRbTttNJnfzqPAmPpLaK4mMQExsI2lclmc0SPk5yuXWxeBRFSO/qlrfDj6vVhAxm
3ObS0tCaaOiscPUA5S+P+te00EjuMdp0Pr8sZkS+SLaQtLkPwjEFHBzYrdaKwERE
NrRDDD5RoLwdeFSFLGozn1IzCJ+OXzRw0O80IZj7VCzjLTo6UTIUNaSlySY0jR2J
FZRYjvvrNH8oCz8OFCc0JUX1FgfM6QB9z0GJ/GO16myyzYR0Xc0JjuFki3M+/fJu
ksAZGZwOzD7mhWus+LmaGhoGTpz/Uko5JK56T/MM4k1Fbo/mCW6aluAQhpkCInE9
NjAGBTXvY9Q1IL7dyt8pZw==
`protect END_PROTECTED
