`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nax8OKxSJQXj5WPi8wDhz+s5nVhBiABz/DuDdU23vHmDhdMtPsp1j0q0o8sM7pfz
AiyEYlhqgAgKAZZBVfsrHxuKiwfWo5wlS9sV3oAVriU61UcDFnGh91rSp0UHGpCs
xQbJZY7/FVUcX5nzjwfOSrGdWD6ot5HZ41lHYsxLjWzrV6yDHRoH+Q0x8O+BPTNY
XJ6AGG75TtGm8ZLDUmHllX9L+GcE3AfYkWFvgXPDPnhOGoB4lxisebKDhaTKopvI
SyWbq4L5/eunmg3Z9Ne74fzZylxFhkCoMBrpIVH++eK/aRqE0Vo4oIPtqc1pyraF
W18ouBPEYxigyO+L76q3RIdomqetaXnF7pYbHG/pQzswzYpIZ4i2U4O6/7BucoJ/
aEhSHlFFx0QsnEr9tF80nXFTzB/MJs7QKwUZVbeN7zObmbvUNH9wztXA7MGl2aC5
RyVgXt1ct4bJgewQmo3+g2DRACJXoJNohxhkRSQ8ifEyEPzZypT4lmbOBwOlWipF
3qZ0RJxwBznnqhnFvB0GrC9cIY8HFn5vSs2lg7wfp9+u491vtoHqLEAQrHoe1cvX
i/DmT0qRNiRN9LfDP95H4NbilClL/A0ffkQ5AvompYl9/92kOSyuH95897Pn3Stb
bfnjCxk/H5fcrxZ1iYmoxH4TKNA2ez0z1CVXx3fGgy/LcpCWB0eN2Rp1kguApJcs
vB4ZaRfdhsWVILXHAscL17Zh6E4EN6VZjf7buUDpru2I8ZOstPNGrKPsz9wQmnTW
Sid4+DlJ2cRfJotVoMtArrzAkGl8FVsu48s9nmpzXnhroo6WjVmWVz4A9ugc4DBh
ODRgr40M2XZsx/UhzqwOogdtSmywxQQRTXHhf/Egr5zDRMC/pxpn+gMaR9lfq9rO
iYLziFrVui3RbrwyXbe+Z41zo7IDt3DLmSlf7ZEQke0UmvI5yT097pTD35e9iFqf
4GhZEYzkpi+Ru//MVwnrl7Zr9aEfeHc5Jo2OjPPCHMWQiH8Qn7brMVaLzt13SG3t
wuLb4l6GifUTwFwxtJngGEbTBjn/6W8vhDPXsrx/zH+PmuXiaBtDMK+Y4NpF+ZJU
Fthiuws2anMYizt0acVDO348nYXn7LcfksIF0ETpuQDRWvr5olWvqhihZpqyJVtG
MzBZu04wVyXQTVrOERGAMKYCry9Xv6FjTq0tQ3VshfRVJZTAi+p0hjNFWMPU/Far
l5HaJ3BRiBK7HQFORKtkKc0dpDDdIrSTeiH4LfTqiPh73QjwwfZKMFum61eP1fOk
yxEGEIOHBc2iuE8xLVe0b0lO2AnVelAr3UoI0gMuclGxTiQuk1q2dH9vr2Db3Sn3
r/wwOjGoKWnfb51wV77oYVY70td+rAC1QiS8B/Ze8l+kgeKzDGPBtY3KUJsGnoAy
CTGkgPN+okyNqm97cwVPJHAbGwRFeK77NH7nR/hQJyJkalb7Uua5+KniheRzabLd
ECfSt2WIYz2krDn1dOXMDAkwOtcsSKV27ofGXJ8AHSphr9o4zjGQ+NHCN2b/usYq
wHk5ybgsoww5EJWC28+pubS/7eA0b99Ztw0XvEuKsEebWA5Fk7YnEXXT4hK00rdM
c8tqfK3hofesXBDkz/QFCFsT1dGVa7PXKjYInMN7AFX8UGP5E5H1+oIouHCcgO3c
JYKFpQutScXLkAB9AhT6EpQ45szdIN4SVx83ZFuB4fDQ/Uee4Fs05vfi8r7CZ6Ga
gdQfLzc+CRamRrSECj6CpWmhwyPTDJ8u4ZL5F9uq35WZvBQ05D1sW+XTa3djlfre
XGJbo18gbk6H9kASK1AM6VQMQCHPEOtcFYK1PvjQmJc11NYrCTuly7XR+11ZGo+9
iqbYJhU2fDIRXoGMWOH1soeHlMMi15cCD2zpgR55ZBY3cpLfZUezS5z3Sh1o1ctK
/Ds/ZhZAO+TYz15iTKHfRYGRynKHsPxgL/9Fx7pLRdq7uhdkYWldPFzIDfYCA9n5
vPEHPNnnkRs3AKSdIhS+smfE+eisQTLxmVS1v5vViKZtTXEZ6PqpUmK7pLPhYmI5
nQAPoQyL4V0+vVMt1p15hZIEhe06X6bHXwqVzq364SPED0YjmnFBS9XdId2aonik
hLOTcgb6iUplstwgCpQ7lv71/C8oiUTIwZfVPHhSKsjXiwTmYMFZRqd+0j7Aa9LQ
GBlAtdq+vRuKNRIbahLvI7J/Zn1+pVISiqn1mYt0kkdkinGloonD3Vqp/39uhxuu
oW5gjd8pVc1iJOTxPCCUwMvFhHg9yhsePeN0OgpQx2DI3RSWSilz+joe0pEd8uNo
GSnaPISpwqD1NZELuuY41Dvgio+XY95TjKYupoVb1ITiqmr6JdsHzo5VswFi906l
vdxJ1785rZZV5Fvsrq6QuN+vcJhXz7U+xOwZmYIdAGcSuG8EHpZAG/no8Y2RYZQI
EXj+zYSWQ6WqmLNKvnNfKjT484U3AYjkBPVt0Xnp5v65HCDx9lmLtoKuJXjhqT7V
jVVkGm2jiMhCldUrrJ5C7DHX+D8o1vF6Qd+gMX6kym4/7LYpaM/fHBSeuoTxcNTj
soibBVxGXmbUtJ0Ns4Y7d1bXuVGgBYKhTJWt2RPAa5AVcJh74d5mtEoxM8UkBGOH
dZA2U0hkS23RmTw9a5eFAFGxKcck1k84TNvUcZerk/E7YBQJWKTalirgGxJ+KjAs
onVfYsQ2Og0U0TFqpZ/yVSj/9ewKM3/18/BIWlHcG44Br0MPRE+huJwRHgqI8Lba
rLmk1AgE+wOadGwXntbuvVG8WRBpP3eW8Rk+D77mSB9Exzlcx80BLEv2XP+Bb0hC
NgyoOb5rPUbQSue9bbSr00WeAlhPMBYRjayqXx3I/y+7lsss/UCiimdVXAHyarGN
+CLH74oiG5zOoqA5oFZByLCVdNhB+v2Hk4f/WxYNPW96iXf0JS5BzttOG4oEq2Wz
VDeBbkU9aNHVdeMDhg77x1vwjqUR4jgB2zh1c6P/AbbFQ1kwBPaiOQoJD+tbay4o
fa29miqHaKRedVthYBzy8+UfvAhEjHEMDMmvE8bBtIFxHo4oi67WuPA2q4vNBzxB
nQaapHzhxiqqPeaqd97cnDl6OpuZ2+pGAm0DRVb0cplA22McuDVVfWI26MQa0C/e
2VjAEPZhiNXPrkXCZj2VUNcviUpLsZNyw9TOhaokQwEwrim3eDArKHivIr7Cyenq
euNE9M+Mi4NTYvd9dxiRaKuSGzWVo39IZBRcjTaWWjQwJTdHxucPma6fRt+6WqnJ
HU6ygeaDsO20Q6wpIdS6stBuRv2YU+agv2CeLU4DRKMsWGQ3RX10/XTIPq0VxGKP
Pf8W7EgyhrmF2Ia+gbtUIg==
`protect END_PROTECTED
