`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/a576VrxtbHqRCeE5HKdCDonzqZo/aUU9lRTe957LplqgHThwrUEYsT6G1uAkLXu
Xgeg/7xcvl6X+HJGzpRPebeDChjhSIvQ7twZc6+HY8ILqLwhjP3r3DsWvUbNiNom
N28fZcOFmGLSDRMf7VQV6kMY5QScdzjQHQafbdiSOgue32a4UcEdwoIwxCSWXFCP
LPBTiy/XuOfKBVA33uN73ED2bTAbSKy8VwFIWsv+S8m03P4pv4RK2BeA8Ca02am1
eK6MC0Xveizg/ogm7CnVSHUn/doCil12z5cxAYqacpgIudLYKh/gD+u4rloHocVe
bsPelobhmxJ13WcB4GlvCJRk/AFJsP5l33F+OfiCOyatyrsjHQ0VNCiM25EmF7Gi
JEOQUbetY7JeT/tqACqVBAUn8t4lxhPgKnF4s8mJ4xSBYCBSFSfxwm8Lv++kZphT
`protect END_PROTECTED
