`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+f8S3iYk5eM8dxBIH9pZLtOwJdqqOvBo0iJhTkNzuJ1XqG/gw8AoFoxlW+nkId8
2ezf0EXJkzhKymZHhpx8LPPq8y5phFDy7UwI3NUV94FtGovoxpMkiH1Pu/gnJfxG
u4Qsw95CjStwtE+OVLsFliLki5Yg19QW/yP+LNHC2uZMZCmupUPBhlj22abErUYT
R8Up/w1CFKmi2ZbnEBBSAgT7EYXECWLjtD//j/289qb4Bqscw9RaTM4ZWlYqZvAK
1qTgetXM0BR1RwjyVOYjh5LvavXqeNoLppS43rBOMrt5Xicjc7PUsmh38jdcAUWg
vFybjlkFgS3cBIu/cwGioycCUnydhcgoNuW7x9Z6vVHBcpQFu2vZy8IL1pRW/UnY
fvkNpgplycFTjdWCX8KrlZfRkiyT1sVPspL2h234qmqdE3rJyL7nIz34LL4Viqxm
LZrxIyPCXfQ+dJ+BXYyMnPOyU8lhXwnYmMZ1mHzIeU21vpTB1fJ6W72hZYrJ6ctJ
SWfyOOtByAumLTQ8d41LJbEqmlChjoRpqSGVDUXOAW4jru3ju7mOh5V/XIasniDH
xu9yoYQjcGY1GhBlbESTs1ng0kbVRpzpqYWj0RgSCeZ2ss3QZQ07TnLKWrLwDmYW
GZoIKqs8RbfH9f6Cmf9QQnApZnTk3h2+5wuVrkbejFA18YvYji7DVj1HjgHqKNpD
8h/+0+NIhKsFrbE+oe3bhuI3SQ45EL9Z7jilJ9/KFdH8HjxQmbpfkUCzXc+JeQwt
yPazs8ZK/CBak6ArgPijHUEHC9W7D+ExYpGeH97t0mnKWSzJ+ahVuwDvjNDT28th
xVsJslZSjovBMOjWVc4iCgEUuWlnKHq56yuYsNQfIqX42U4J8IP938P3N11pLrTg
j0vQHLmax9VXRHlo9NdcP2iENEbFTXT9UnupkuSzmeTnEt935I9gCOUmgsYS51Nh
oi0AiGxfVYP2EIMVxKzAuLoAZAH81wtPX+HQy4v+3WHaAL3E7cDjEo+H6AnQeKsR
pggia163nO0FRzy6tVfz+/w+1QxEeezU/6yS7YKMaWHBY/EdBY6tRI+ZLdg+OWVP
xgFKOO8UUtr/zsBzT7vKgWhcJL1dtw03Z4GQTS+zU4yrLVCTdVa2Rzdjik/v3Vn8
oXP8EStUW82bsw+nKLCzy2JXE31YNZe69HtZ6Ns47uX47IFz8YPVDKMGTnAzROjg
HQD80KFUVMI1S3mwYQ44E5P/9n3ZBX93994kiZQFRIrcNbBXb5xjQMTSIEb2BJZx
BYX1nUtADXhFDKOYJ4OhK+MYm8d4KO238Vpc8VuVAV4vgeNEIvHrf4Lb0djMkivu
7sTnzpSWINcPkFBi24SSTfI3MAkmz9rdRtDQDoEneC+ilLd/Jkm89saRhRrUvvh1
c1vwdxP0s3JovMaOqQhrui9427iyulZUzr1GEyVaUthSn9IYpCi0V4iT+95uNi4w
00Kw5xxq5Tunvevf/dyQPyohkJBX4D7in6Epyg6wmhnusHvKD/gOa5vq/67540VL
Oe931xrT5Pjh5oFKiGWx/1K5YYIIZZccfLjELNYFnrluED7Ogc7gxhwZAtdRpVmk
H3QCVPRZfIRz5LKdTbqrZsWNAN3NUM9X73uFdmz4JbeGldNPszJhKY+nMgWojlxG
vTEO0Rq5ol0/UQHXTyrU2cgmAAKW0OvVljEPZFD8LPA=
`protect END_PROTECTED
