`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dag0om1ap9E8ck9L0XwptTdAIvOd6D5WuUzXLb4w1zXeCUPQjXEbQaLunR7jKdmV
SkXVbfL0cuvhkrcbHiEgeiPG7zEk0pQH+nkey/EXwQfi/LLFGq4VTMufe5aHCQjp
s9hrUhrIuM2W0y+EbZFp+SotUeNdciH+m0Ck31ZPn5SKu7faMZpyMuRqfSFDM+K4
CB7ZwohV90XXhHRHd0OYA/4kBSOoyDGCIxXiu65ekrU30J5HUhjpykfKnBYRxwco
UtHUAWJZnwkr4ImevKpyH35eTRtaGHs0SlDcfZW//89qYU/89dTg1AP5zH6eWky0
MMdkJRl6hHDvT/lwBZqwcpJb/x2U0P1pl7O6Ob0YsERfy11v01WXr1x2MBkymdKz
T7LO56AXPotAF/hANjV8MyaJ/9DTY9eS/Qdzu9Xaxsn/X+CfMFm65SLbl+6YIuXm
vsuJqT0Fn0UuRHDA+2Jbh3csnSdbBDuUHgHzenz5qhxuYWOc8Yyvl+BGq0cB+SGJ
PCeUv1pFKdi8q1ondxfC+xR6AvRwBlCVut8/LxRbPdDKIM8nF0m0cSxd0Sg42LqX
4wYRpL5mpmk2/AMfL8+RRWGeJ6QXIBKEb18I7QuwhP1DcxSEJwOqYvLUuKbGDdC8
thtmd73wMl50mXNwn0GFRGi2pbFjhQWKS6+XDWijrjF3UKhMqmd3jsT5ZEKEeb4A
oIp+1PNq2ErEhICFvaiKbhtFuDBTjZ4swJpLPjOzNY5XThXjPmoEXaBtNapKP2VQ
TT4WKRg9b3E7vRyoOnl8C7acgmfb86SJh9koPIje4KvxOlyPKYb0Ro4Vv+AuP/wL
Fl8N9p2IL4HP2xCVac3JlUVJlkRVttFPFqvnEmPbGmvuuHzvXKvCG5tf7DUSyWzL
H9zCp3Hw5vfgWBuEchR4J08p4rubF8Mqzv1G5mWrkbdTWe0UdnCqzhXzvZ50ndLX
l4FErtC5OfBIxVwXJByMGSav32bDDO+uhzB9QUAt+hxP62haicNQ8P36WxKxGFw8
JL1Kw3OxgH8kCF3Xz9DESyrKLe1MuZfXtK8MNED/hBiL2T9EU6/M1ThVegYJZGBD
TbLd8QlxtP8i63Ke61g71UnrvWh06nrMyR0j+27kYD0FvcsvbJdCjqTBMRzIb5Pb
Ddml4f5f48vDLRnCVkARJ3EW/X0sLykDoP4uBpx+DPikjkk+sM0RMTDzvk4uxDOK
fLpKMCYXDuTu35XOmmiJQir+C+oyGMWF2MhDRdWbh5xiLtRo3mbaf4YIkkWyWaav
u9PCzLsPd6DSB3EA/F3z/MrFE6KOg54Gy2j/VXbzlIybSHNBbQlqJXkaTxsqGXK2
qsaSPmAhEvommVnZs8OCa4NxvhiQB9fAgzGM2eEc13/5hR/xy5t/mGIpizgTAe+d
FtlyHhKTn97oAjiOsCqjCzfQUJB8V4rq/52F8UU2W95T3nPY+xK6N7IPrdHNJHYL
7+2+RtG8675NGmMGZCk7C0HDyZiwakVGogG1TXFyrM2Uy0PLm7CLxx1AB1oZGtn8
T65LAGJzirRFAsphKrqU2VaxTfzv2ENOsH/dPh67bpx6xWuCklmrq2wIFcVxpwu0
CvKn0VjSGQrOCj71AkAiNFroiRaVX1kqb6kNapkNEM+9ZpYADpt3t762L1OiV/+n
ua5tB1jJLOszAVC+TGjy1YdTDU+NklP51pBN7BaYoAL01rccKvSiehfUH5aNDRzf
bF/XQa+CwfayqGa5HdXsREn7AhgAA4Y2xvv1M04hCQ13NhRYctucXywOFjpCDaP+
7DRk60rSEewXbWZPW7HoDH7jAsF8BJgAo324kPuwQU6RIEsGVCMkFxs2r/MQq+St
AlzNO+GgQ8Rqo+9wVmTQSBmXld8akRRTggI3EOvwvN5iSJDpPMoYLKdB6QKsnNUR
8wsVlYn2+IbMSNS3kX63/tb4K8aKHcggoKGcwNd/IP+2Tr+MQ8Up0PRJGKWSfWCC
dSPqJGpWo+8+CibaOb4241yNxEjGQC/AVyQifnFbTCDI65X0cZKs+rrVSFsl+yRM
rfywevxfJktPJYbBsVrK3F8H1ihF4AeDNxHwlNNR5rPl8hknDSVWN+/VYLsSnSkD
kVymre/W4KJ0darMhUAr8qbMwcnT11opgH6pjdwFRSMkA8F/RerMfevd8dUcsVUt
62FoSOhmG1LRUPyysdnzvZLLnvuEUyMfjxQ4USYSE21uyyjjY2XH9xT68lQwnhMi
mnQbTpgw/L5suo7vAfQJ2u52PckhyuOQ+gZ7P0HzdpJM2ZwegjOROYhG97tkEWHj
+HaCg4Zwp9vfmGN7QWh1HA0jf2Q2m96z/L4jUqHivyDnvZQwzEXjs4YW/Ge+V2uG
qdGgbxy3mC8+Lp8TEyryqShWfGcXQzEZpDQEjQJ8bPrID37l1NXR0Qs5lNqLiqUv
vz2koj3vmK5ZCtgJSpfP3Dj/cdU2RknC5RTJ3xzRBQo9ZAEvt4lD3YevAcZ+1sYE
CFGkW2arVdwVx1JFg9m7COn8Gw2Uos9/Vy90b1R6RF6sPnH1nBwWMh+EBPJq+BuG
nLRtUFfhCixsS3Vo2JWcaOSZ9/Hdo8pRmOvRMhyL6sBl0zDFumqVnDKviDR1102S
MaQvVXCiRCgDkoO12sWQQjinGGN8tA/DtvMOJaHOb/qfg727Cgz7S/wpVxrmaeWz
3tE1LnGAor1ctbgQnZzVm/yc2/hHsBJMea5q0+LGRArUjd3aO3xXxyAX5kV0x6Ae
5uADm4XQivTADLtygTHWR9nHVLszKxUHa8XNO+nHouQHJZ/YILlFUpyv9fbLQPhr
oKH+jLz8MP60/NaBIA1jDcIYeYfz4xZpIjNeyKDOGoNuoUm2HB9spQDTH6kiquzg
Uhg+lTWLYVLUGR721gqjR3/tIUBgRQZLOZYCBfbAyWTI3KUyOwXvL8vNNUdl/dnK
jgSRNomTdeLN0+tKBLPMQA83Pi0bLt3DqhL5N2lz7QOs2xw+9EIezrsctK5MAGgT
21NYzYwQTUJqUwy2d2btbzbGXq1obv8fZ7lbxlx64SLpFqJbco6TiF5DKC81/Twg
tOGYq13/OZouSFfXHk6mAQQ1J+gr3zNKvCNaNXgECBLallNTMKl82mb7dLmSZFYH
opXxbH6CB+ikR7DVA0qWtLToqq2ME8YkoPGfFTBFLB4AykVWVJU+F+FXYwLxv8+k
O+PkWL8tNqLxvW/KNvrl1hK8JsYcjR+pq2LcAF/zyYthYpNPvhrwIMIqkfXFFeXO
WI/qRbGyWLQHRMmO8adgkcf13r2aDyAwGEhNzvJ2KSVYYfL4PEUFu0ZguLZbg+kS
Ve6+ClI5n0u6/A8jhAEQGqhkXnEiTrZyDui84c+JgQwTqiHH+RNZ89sYeND3cM8i
IHNMeBBiK3Hu2sfK77nsUQwDJtPAGnFiYZmKT6lxULRQ1Ro6beVu3TEjIAIGtyWs
a6aRlSEtsItqrOxi26nUqh0jk01w0NSc3Cn5updO+tBDR6M7WmwpUpbi866qiD45
ogJGINz+BKlaMhexIPgnRiEjrP+IVTC+D8lsk+m9cAh5gbhJQrtbm6vTw1RmwyjE
O+v4VqmZW5tv3J+r0DX1QflUwYCTMq+GWANZalaMhh8mkXEwLlk40bYPhfA8m9ls
Hxiq0FeImrZ3vvUuvVQnc7LJUCm2yYf5rflOWQ2BnS1zMfYb5j+S2SmquJcMj5ts
1phHUFBfrsNWM3gy6KNPCnLmmBQBgTR4qQxpz4JfiDmhe13LStv3YLTCOOf1gLC4
7MxQKWYwKKyzZUn7onOTWW14FvXndo0AJadk41AZNCPcYTpuvIy7iwRp8mvRGxv3
RRr4vvrvh12vjSrbDM7lqsFFoWcmOZw2IujAWcUVezluDlX5rxtz+1VliWguzrdU
QlYr4QHU6ck4TxSo+Lxh/HYqWxJnWJLRKB+i50KByl9vMcprTaV1ut0XwPfsTW9O
X69TPBqEReyPfXcoricmpYImeRfpnAYAX2+VIofZD4QNWGGV8DTMrDlNsNQQDpSe
DPVwnI2hoji7LkKgSbOjFg==
`protect END_PROTECTED
