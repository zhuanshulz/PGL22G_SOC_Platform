`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZcD6pwipL4q0hI9PgwRJdlWJbX1V6FKjlEUmwWQkS5kVHQeFF72bR+o3cXx7m7pO
w6soff/R4Fu45O1o6sJv66NmrSjyLbH6VQNaZrcrxeZXVd+kpe8hIDtp+pMvnpFi
SyK/4KGOi/DO2SZi0T9+DgcnmcB66to4d7J4BzsJd4heeNVuSM+D+OrVMVu44Klk
RMDbHlqKM9az2NbQNB4RbOkpHrzdBVILFh5xNBZGqyGeKSrmdUNJvUPQM1QS9v34
hLY55F/Lr4cJE73CqSGqgVkyCKwhpcuejbeNxXE/I5NIpVmHj2ISknF4XOQvUjGr
8hrWtzttS4HWsGWMy+q0c+HSPBxA5eWMoPmq/IgyZesya5nIPUXkmoipJi0C7lru
bZbNIxQsCnurQBs0s1srpy5UMK9+t8tenEHJ5wX+ZdRB+D6Qp+xhaLyScFg+jzqP
uCfzOp4ih54pZXIfsIUomICSlma4hB6SWDmsqPZn2iz7mxt8upayGm2LAqB1rylR
9CGnno2M3ZiQZIWFPSVyjA==
`protect END_PROTECTED
