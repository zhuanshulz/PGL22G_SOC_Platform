`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBLoYW6DOF9Zse2nCQvozGUsmJ1e88UA+Qzhzl1m0yeQQizuWhmR76f75p4G4c+j
y5m0rk8CVTBwxXtrcU5aoZxTz9BYFGXLJH2PmfnIgEr+e8ZJsWaxRvZ3hT9HSYBh
saEwW1lFp73vZz8As5kfVJtphFyUlgyv4FKtD/O+33sUnrYVNTDeTnRtm3PaRMYi
mnHcgzBA+sYRWioE1aV+7oG9NkS52IiHveL4NqaNdkAQcZxECik2+bDeFtt8pQyw
r251xzlewHYiMl9qls6c+Xghxm7FaMjws/Gp9B4uvPkRulYm6a1fNiDQV/Ybz+ZZ
lqQrd+vE7A7IpN77AmMEVZDY1IADsaw1FpL0QEhrSSmto16fzeXaTmlTHXVI5FPA
iRI5pOCgBckgt2XrKM3rS2WBLu/iieKc8FAhlQx2kYTPuAKJZHXYf8bx/Qy+NwMh
LPglxfMsjPiOf+QOUbTItQ8HudmSXr/tFoj/0haHYXZHhmIk5nf0AxekE4YXL/GH
I71p5s4keRL9m/uOuV24iN7nriwfwiOIsFbszM+52PunQ3Qy8Np9i2OYyz/w3iTR
0B3DAjU9VOeMe9VT1RZ3mA==
`protect END_PROTECTED
