`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVBkPtfjdp5xKxPi1nHK70nH9+IozLa5OvwdpQmSscwaQv0BmY4noiuMUd/3JV8e
ajhaeoqN2/p/EJDPl84edqi2y0bWvI/xN1JRfj64A04ce1O8DyYq1/oQjw6ALH7I
N21BsHaqy4bIwiDnqhNQJBHrAb/NngF+7IzWly9myP3Yz96XBoE4vDeBgAVccvvF
1EqW2UFKsjFbDL/5MOtT4MaEPiE7pVsSS/SnNL1xzTACeun6f9aXQ+bwkQNI3yGj
i5K8Z5Ss8hl2De0UFkp+Q8XmLAquFw8xBehtoOGSYzkbIg3wj0rvQ8sYNLuTF4Z/
qDHJge30TYU9G+UK91SJv7Ot9aX5jq67K2E7iTXUtZ9bOdCsMNgnUUv7TbUgQaGK
hs0UPA3rMUgm4dBKTrfUxriPmFmBB8Vc4LTdWFjZeLRV21z63TADI9LJUKoD3+va
+ozH3nU8n/9RUiNEZnpxuscshR2hZ0XKfCY24VeHiOXNMLsiKLW+qPVt/FsZ3AQ6
5LJSwmekR50BIS7sv0uw4mHbGBmhM9xWG3Jo4iKGPkxH4Igmuglcpiy2siXCC5qu
AGcK1kILBHq2uIAivdGrYiLlYjv7cq8xakuI591j5RP7FA9cOLfN2c3cBJVQ8IkO
yPYxvSPVH76zdxWHcKfcogeeI88FzHhwDvoPTEbVC0m7aNFRWFoi7WiwftMqj2Zj
`protect END_PROTECTED
