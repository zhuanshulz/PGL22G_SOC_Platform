`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dgM7NCtNen3dK6TYQ9fJxwMMJtX6NW9+VctrChqMzl+f29A473URwBpY9mL6+R5B
qLtVBiBlrIYxg4UPOXKKhlNG9Pp/r4MVTxAcfL43lSfumcf1qnvT0zoQyi7ZJBCf
nDohH70IPqCRFN+d/a7yhznAxgw1+GPBLuNdbfQvPdpkW0HD7imC/crMhrD0NDn0
4idw99FuM9TgvQayGG/3qGObRxQvz1YrbU/9TM/iLNO/+iGf2z38J9eZH0m9poJi
XGok1sOndfHt8OjX1yDfuBNQqs63gvP0hoUnAZ/7ICMsY5gKGu3GOKvYui/Z/ndP
2EcBLe8B7OZ87IKAP5B1F42ZsqNi7SI2e2yrUeBqNl5zNIWjx7G5A26VBB28Ai+z
uiVnTBRe0fWKFxK75nuijWeOpZ6U7VVDhsutcSRqHLATQA/0mLJJq632yfXiIO0i
1cJjEuhZ6eXoz5dWeZYulEhzdKI/ZU8suKeydsP/LdL3rLcHU29XWIdChda+iSvx
kz+BWqvTAMBsbKZxh3GT/4wN9q+AzIxfQYFmx7fFEUTybZyywjWjt41vIJ8VGk65
BdwpVmBiZxXxNJWO05NBxow6vQd8krQrNiZdvViKCEld0WFYgsA3ffI/lSlT6INs
7BD4kFMlHJAbefiXH9PbZgqzvpa8gwEpO8yYnokMxOJSmtWSungsLsOZaAryZIDh
ARtNcAcp4A7ztzuB7Lnfu8pkm7Eg4CoCYzbh0+YlfNSxSKCqPh7J4T/b2PerQyv7
MKYU+wdTjcDx1Av720VCexQbqB/B1cOnaMCBFSfTA7x+S/rgWgnp8a9SHUICA2RQ
E+Dswer3rd1k8+UTUg4BjfYVlO+h4LnGuvQwFXNvqnIu8jNWmmwK4HL9vYTfqC7k
VmzWl7z3ieckB9AYaDmhJvVUAoAsOjrWcwXCCPvBQY5RcZjtotNP9tUl0JKVqTQ8
axSK4GUqD6So64K3JDl02yQpNn0FzoGMII1/TLvZpwPqyBCnlGMhnh0UzxuIKzp5
A6y1y932HslINlfMRcou7ppCdHgwpiOIKcz2IJ9iobRHx1w9/nzREK7tZ3+GEAOT
MgjlahdaErJgZmryzwOnu21E4HPY8+RqP9s62OA1jmBK2e/q2uTsmNcWcCRuzvri
sAeAEoS8EyoHVx71wkNDbjCICySsk4CDsQmP6pN7ELBIoFPmGlhkRI0nlA6cd3KK
imRMCqqcHp8WRpn27WXbo9yRWFLgto1bgF7471c/v6feAa7Kh/O0H5xXa50dAHuv
6OXvjf1guEig7AN3mfDxIAYKMndN6+lWTiVOvZSXvFC0fQYvLzOI2s6MangEtl/8
RWwQ2pJDaN/51HaA11UearGpRujrMAoBDMPHUHx+jzMeVELO/LRsD0kET7tVj4Ju
SxpJHdaHY7hrKexQQ6T2oM6mgTpkfAOdfEZIfmyzkb/pO7SxPdHd72mjT1ZNn/np
tGG8tjkoyruez7zd5bI+RG4jqAKQM+82sBYbrCwTLahpzSuFFBdrPVF+DDXqR1Wp
OWRWVns/PQvMbwfQViQu23ijR+Fs44hgVZdaTuTZEcPHzvEGyyJWLzoF2izHnViF
gYv08XO6Kf4c2sLXgf2IJiB4l+q3FqZxS8aIrSJ75idg32QZEN7cpRlp2tFZjVSI
41wKh1uRMsnsqFapXsCtULibHMjf6fl2D/rQQ9CxNBFw5S22G4EUrR/6WEw+aNke
RRMwJ71PeBYsfGM+dd9g13u9B2zp481emaYyNNyhWYUUt9BiLbDXgoNvfu1uq/gm
VPJ9TVKKBQYl30rCIBz3aBML2N1uWPrw65PKAgao1j0aiH7ongT5hvPXjeTVPZ4n
FvqyOVOLyMrG52dDaVrewjGE5umoZyYdMfgnlNFcmUJnoMJ7ouNwggqF/43MWhCI
SSomLhDyjKLmL1MzTQIbCRd9ZI17xDdZFxhMnOxdBf5ox/oC4p/B39InpPXuQZR7
kKikgcTht7xLk/VM2in6Y5y6QbK+6nXFEapl9k/g7M9H7SYTOvkbK15nrALKf/je
uoRVZq6PDwmggLZSrzcQ9gf5gRz3rL1Kj7QPPNYVlNEhOYrD3EdqssYMIE8HVWg4
HjoGrIYRRNGExDjnt+P8fzSaZaJz1CFq3mzKnGWwU0o=
`protect END_PROTECTED
