`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOFU7JqK+vP4+fS0g7UMRuqjvSF4Pd0xhpm5aYLavw3fEaFX8ICXoyiJ0xPLZUgv
bpWy9QOr32vcMNYXe2Pcd5ly/FteA3gOVloOUuQn1CKiAPLm8sqJm0RtMN64QK7E
PXZ/nt/WXHz5cZ13OKKwLLI1DzkxTFmT1FMuEe6ZmW67s6NURwBCXzdcJQ8IfGEL
IoSMmLX9r7TGf6+5JmM5+wzq+Ssc78IKQCN4D++Zbr8MgMN8fsfPyQQQSRIgAf1Z
o9u+cYFM4z96SrBSBsJ0H+j9N6ZwM/E15fUrVlUVjIyP0PMByMIP87CDI12K+TuA
wsMZZpfztoDtJePE0lNmzQ6HBVhXvOWxHNhFCEvL3thGRtgySkF6IBeRimiYavz7
c0rDoSxWnDi6Q1FsIy/7FaXUqC0k4Mo12bDYHdE8CsPZHOugR76P/V+seUrxHhEw
B+L6yuMkixV3HgdlbFnVhMGl22W5TyYmevIVepI/VGPTUlKXhmyy315wOtyEtsox
UqiwL1cMTzq7jzjGkk3j9XiNylU3eRO5pVdZ2hXm/dpLOO02ygngQ7b3Uhh4+X40
Z73//mW6oJFSc77I/M723A==
`protect END_PROTECTED
