`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rYoRV4NlFIvkMUJHGifr00x5XOFD9WZR0X9nKVmFDF/j6JR6qH7eFpZATqoRsFS
SS3AUNsi65xJPJ6qZLqMdlH1K0FTZm18BWN2AxLn2rLxBwZoW21ueEl6uuVfClY1
CoZ5pslsntOFHU/yeYdM73AYtotJX1NYu74WSTZmkgCsI6f5rnONyAEIofwXDK5Y
oG/4roZqxcGid0DRb1SB5OXjO/Bb3Jg5Efjf5LJ2r0MbjexDaY2P1j/Y4IrF0/Ny
17NYZR6dRy/wycKRP7bj7b6ljwMJ3EM1mQDca8mutWxgfRkehILjHSmrCgCR5PF+
mHNE+7cttUKbpne0cohmxyi0HnhlqrFoEVHiuHim1SAi9d0MBhh3b9uOG4sfcUmP
ywfzX+lzQI3rtGYFOOVHQXkUFQXoS5vLUkJB/ay+ww3XmN7d5nIoZz+CeqafH2G6
lT2EiHciyuBKvtsuuldmeS0pXjUxokBfVNPIoasRgyOmKo/iPpJgctwhnrMqvV04
OmNg0w3+MPPB049wRXO2SajDs+CiY+0hma+U6kgDqx6l1/HQZveNpNyX0k0zwGvm
or+IAnfhgvwkDB0QvUaSLrRRhkpF3sLwmU4wss9xgwZqDDTGtifwsmoVn7GhXJ9H
uzPRAhBwOI2K+ODM0sdA4ubvaGc/d9t93eIIN9YJePX5vo0qy++odc+A75Vfmy7Q
qZyBac+weo1hWd1ILDMDipej473Y9dq6GsoMpbDF6YJJnNGudUZzo3MlCXD4YRcc
1brSE+a0F+o6c40LgZ+8SSDU6gXM91PULOoES03KjTNoI0gavTNBESLtdXaTPYun
uYNwHe1hHhfMCD8Kmy+0hjNosNepxMCTMlb9XXcMmwY=
`protect END_PROTECTED
