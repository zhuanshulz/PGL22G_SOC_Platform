`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/6AVcht5p7ruVXyifeDTjqiamB+tgozvuuu5swTFPhyQHkblHyZqkw9iTN1fYQh
Q0aCgEJc/xiXifFyhohF25QYiMudA0gsKRcq1F2vMfxC85ts3Tp4Hsf3VTLBzGue
Abd2wsKxjAkqOxvPgLFxnAZkvF8NjdH38pK2NmdwobiAK7x716YebcZBrE84yTzm
DwFYTXdxfDpUwCsNMSrzrYtyNLtEIrlKHqGpLjtXsrHqpU6L+8futjZwtLGGEHUO
lh1juy0QCaEafUSU9OYHUgAef1WIJ+UnN6IloSIbOkE9QQXXD/gox3IjfUj79Im1
fv0PzoYKyhkaJSgYn2YZVd789MQBuwuFFX8/YsbgnOT5Bd6acCdJcN7D9sFQcvT9
Kk0aNdNnlrX+99rC9bgUpfMpR73mW5mzjgHjRJasMdYx15mDF4f8sEuqdobLkomm
mYulhFknXn1uczoig7o99oh7NvN6jAcAfZGrLmZTeAERyORkX1YE7tde56m0N6S7
rTLGwoVARXDWyT9dJEEyfKG/ypDM0oreJpm7Q+KCmYveHXRrbiUa2jHJ/qTjI6Em
lpu87nGUEDWzKBC4T/Tv3F9VUSktH9LApNiJ0WvyQKF9TAYrPVuVukgyi/LdAMnS
fVrt8KrxiXs5ygQ11TagSrE427xLkMw1t6tn6ITtl4ByLgeHOD0r8/D9kHG8Ch4E
rqnI/C1Ai0AIPTXlBcKJMhBpEZtXfKa6shVZewzEQt5RdLxLicIVUUtQ4mut5Fyt
PtWI7yhYBgM6c/ZwkEkubSsdfrsfJiPprYU90uvV9a+kLQw/hKp8WgH2d3an81L3
+MV6I7qNgTP3Z5mx4ETLPPb6zzCxFEyp+RowkIx56PTs9wiM6YhHXj8g9Zb8WoTy
dvNnxOoamMvXEFpaRtX8sPWb5B4OVwq+01DWNM0KoMQ2+s3lYnhcPaRkpwpM+e45
+FhwI4Jel3+NZxdrTT4fKS9dlFMcQ6OWBx/XSgVHzgRN+fz9DwLPn8hPcYDSXKZO
z+wwNHAlK6unsQfm1WJ2VAacFgso3lDEBp+0Y6OnmRQ8Kc+fC63HOp+H7jTo9XrO
JAwKcHrbUzB6kQdiGx+qLq93hSHSfmXkrEnDVJVQGD6eIz9ShVenqsTuKI0r3lu+
9evIGpBoCgDt7vr4Q/18rfX35dUQ7EjaVhnp4ekf7HNyXtrbPvcejX/H86xRivEx
ieXOnmDP6j4rPDqQ/w2hldCG00y2+Ieuw/Q1V8lJeFuKqHc7HvLS4+8bbWOPtujh
B/ITXh3SpYTBDMNCv8XxA49rmxEpmoAd0QdIm7osglcp16VdUzQiqXGC86jMZw63
oalpRlRN8HTUs/hKMtDg3AB5y4fgN3lQ9rCprG6RZoa+hpLSPcJw6LLKF3I7EsDW
U9xl9hXkUoBYkhclrj9UKOaA4exSS/ECOXZis6X3hf7ieYTL6y4lXA8UHlOa9Cp5
u4gfCnonpq9oLWFS4nuSBw==
`protect END_PROTECTED
