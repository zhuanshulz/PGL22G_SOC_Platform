`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcwyf89k3hMbqRo2ZrU+Vzs33aeN3/EqyzXVV3SjqwTtLPYRTFlesKVBcfibxoxS
UEQ6W3NDa8RGoVIua0ODEWeljNZCeRkj9s76fmSZGvkC0U/1DXv+SkeOoW9gYthl
w7WzPOZR/yyATyl5s+TYEQOi7rYaZjWa7a3soxmCRPfEpeiqoyebI2kTTdB8obq2
PJhUIzxFKE2MMaI+Fzc8u7ODE6BBQWIAHoWv0DO4A+Te/IMd1eNPp75G0F/9mcjo
0QGL2zLyVfEWmAuRymzuaH5gYs22PCqqsdlvQvb/+tfXR6cQ/OmkN4SCMNmUdxcH
9ULLFtLDDESRBXGuXI8AujLgdfq0wGzgpeZYWV9fvQDVwgdDfdO3lZmMkud7X9R5
Tbeajdhyq1/NFNc23AkOuqB3cTzSyR0VeHK5ExRhDb92NVafyooXQ1B4IK2eQ+VJ
aP+JgnjDLyGrtma+O5oX+HtOpELzQYja9nQywnYMus/8K5h9m2gyI+yGN6myqb4f
lzE1dYmw/hvzTduksBJ5sWbdU97HjXqCmxSqqi26lz9BqCD66LU49kAbLsFXZ1dM
njJzecnLmR1BycFLlh6vVvfh3pJ4iVZjtxfiQlV1Ny98In055k4smL9tr7aInVLA
63iXE0WClaTIyGFvvat0EKOCOGLv4bhk5uFkjYzVIs4p4vpehdU2GCXT1wbxWGn0
mDHOEwD0OOaUI4QtYCEc69E1Kv5phcCUctrZbAxCRgEp+IDA5chdKYqmXBShq/ng
SBWq4+OO31VC/jgKp/9FjVrWYkuVQ/Cpyr+7ZUey75KL9ZwU0egjvV+rpUf7nAd0
`protect END_PROTECTED
