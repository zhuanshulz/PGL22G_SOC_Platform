`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pdq1dZJqYQM4LmKUU5E/yglYfxXA/d+OVKaxz8SxTZXBqLt64/vobsjl2bJxjXfr
IgLP6FxJUnnfxfTYHq0sQ2RtTdcbqGYuvyDZRVEgZlMCM5hKWULlA+XuiycYMJO2
IU8KeskY6H3HhFz0ClYbmJ5JGmYhwYTvPOshG4gvw71uUnw1ufno1+Dd/tcPtw8G
tfE5WHaL0oMCEyUk/r8xuiKx7ycD6dD12Md4v6rvDfsC7sbfTxGCmFEpDAfRxNfA
JT6REKRLcn2GNQn8ibVp6itw3+Vbi/NcmFzmLYvojcRVIybQJd9UW48+/OhCaKRG
5e4DoyW8XjYtVEOksKPdAZAtbZdHrl8z0/gZjNJPoBE6ka8/0t1+AOajkDzv4+CA
RqKwqxXUAZboMgXH/ps12wGW79cwfuA1A2fXU8AgdhLOt44zIZL44bTEKPGeCCUB
UWNTUW4xgos+O/+jywDyOgPaSE5cmtsgGLE7nSI4+eLBZFNob771ihdyvSruBMRu
WuCT2krjQcYmHuTreoZ4JdR9zr2CsRpKwpEflp5wSTKA3Ead1b9x7emzLbFAmeWZ
fyTB4wh2xj1wza3Ed/frr1c7d36kNJfxmEsqPZ0bs6hn8ZxZ9q/jJwBs2LM7dUeh
KMoh/16BaYhai8aJ/ZH+5jK3YbyNeFYrPDG+spuCeiM/cDNBCdzEJbTAzjg/PMCs
uAmABqGMxbldJV6IY3oHuMNH2jyM5oQPjkDzwoufhLnTg+mG4L5uNv8SdRyL+jfA
WZa1kxokvSH3D19PUgIj2jEcbgBnSwWu7G8rXr+r0dl52qF4TugDy+2dtQ3R380f
OdJBUjGjdORHvk3YaUN1fdeavZHJxEPo8hjKlPKIRS8icPiVvrHDSg28+FoyAnEi
iwh2T9FTjOBtt+TZuSI5JqOvC1sP1sU5NMTlIX5jYD6aajZg+aGeUpuPPIB7sGy5
wnLaHm73Fm9jrM81DMou/8JvkTCrZr/vcT/GXzxnH7PoPJ/3xw7PeHsZYHmCKbJq
4S1xWvSAPelWoFs0/Lb96xwHWUuTjOe+wV9JIMSJXK1SRTBN1cz142SJhERYmaOY
U95A7l5rk+UV7zH7lTdjJWHLpx23sTLHBqaC/SCITVQNkpTABNoP8J+tmxvMnS0f
tvlysOSPkntBwAKzmsjjPzsMthwgIsiOCXpjf2YYWy0F+peAJRbnlML5dygQ585m
cunJOPPlbGpQdbftqG1v3QadEhGiY7OmcgZ8Iovjj4CBAYRVEkJuzDPTjkv1NeGG
xTuDdaft1rkzEm3JOorbzo8YXgMyNkMk5s9oyidYErqgrTNMiiEgiR/GBobuyG+6
X8cl53u0xGfl50HcCWx4G84DWBJ1ZTmrULHQLFf+ba7jl9pe9MeoFdXIJ/41klSf
ndDE04n5CmGwkrI7txha2Q4WHOu3H4hocarFhrrfkVY5ZgLxgoRe9G1hJ3yM7hXj
JHdOhMjgK6rXLsX3CGBaxrBl8Vc+0+N8sqdvHSdJHByCA/52YA6Rm6v6QKwnu6n9
XEe3eXDy3Z3oS1zCbS4dh81RWs4m8hgD94/ceRX0dcFUtPupnjZBcyn+ldKL7gwk
1wa+waBwaxb+a8bXYUCJOCeTza1jeyUwE4QvBEFGunFEJAtfwWquF9dugbOafqcb
5FyrViGTklmTAu1RKiuNsAKjcBMnL4qNl9WLz62woHZG4kcpTH8v6Zt8W0SCyqrs
E3qJRNw6yLAhCWVh4N0FJIvDIYrXMRZEK+8797IkIqHrtI6DHc3VEdXzbMhP3cC2
/GsC9oCwTlUG/mA3iHqBc8kdA0keHCosO9sj0BdLRnZrprUbrvPMtyzS9h7SncMv
j71HxMKFMPhEq9Y2/3PmT0aGL2izyBdgPuPZRydnDDvjdC1yoUhKk4Gi5D5cJGn5
BTzgro+WZvOC1azUdXGlPjISQJHYAK7MqUfpVuJEaF6C2AmNE/csopEyDtNvqw8/
Tc6CVgAtkZQwTiwhwD8ZfQhGndJLHTR8bYxf1DYj8BNhR5Nh+MZXTpUJzlKiidkv
mkt0Vb5yfeU6PvH0LBSkR1RunFQ4ZFgthRba1oa5CE4lbotlrUoXrgSBOV0GC5fY
2KaAkJPVja+J64VlJgDQkjJ7buJ7mp+Y5dURo4tlqw2U5AuiwkDwZJzexmF2k1Gt
7g2W2dK1KR9HGJt5VigE+wWZuUiFlYzcG1I1dgLnsGU6zeo6v/K5IcHDdU/4zc3M
VRLT9squu9qcGnjgekY9adLf8tnfYYdKRzI3LK0/RN9U2CSOCGnNYmcYHfj23o62
IbhQF7KPtm0eGkSDpxAix/dB+MItigIIMoQQVdh0s9AjD2a9dYPUfHqm+X/Bu84F
QvI6Nz1KovDu6QqxMaKtc0xl8K7FX/N/g6z0VyAIffh4P/ABPXHt2MBus0on9JDv
FcPDREKAxFkKS3s14d/ZaVXV7LP0TlOI8FXxoumGNkZDqNbDqMsMx13EsrGbTMYB
qCo6Yp+OcOIusoPh+mubHeH0qk6RHAxxJxaQ4/8bYyDakIGFFqLvmvleleTWKLKu
7/0DIx1VO+gPSQJsQEoWx4of/6T4SGYiL7/Dk2xEae+cx1KglsbekcH5ok8m2xK8
spROebm7sbrw8jFGalEkdIYOBy9DM76AD4Rw19wgoaPKK6+6H6S9iluHZiyE7TcC
AwY2cNoEXaLnYIrXIMOn0TVGEFReRa6H8xODv+LI8K32QJIeXAZ0z59TgIUZYCCr
l8i4tlQMYJj9o2FapQ3gATfiNipeGzvRpTDhWZcRIoQ=
`protect END_PROTECTED
