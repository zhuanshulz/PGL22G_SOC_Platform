`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DJzxFLESa0BgT/vEhmbuXcViLI4cGm250VunkmQiQId7auGsLqU0xmrzOe+nhFMG
u2FvDpaqZ0UpN656rs3ddKn9/6U8JkA0aTYRqGlp7IKLtj5SZe3njFX1Dn1bdOFa
UnXJthekVkVTqlJD/VQ5SIvRZExrUG63VzGjLViIfSHvkuJO0EPTp6wDpesgttck
4V1VMhIlf6mTx2kv4gaC+gMrt319aSzHq+LIsAOY6DaFABEX86g9jUloxD8/+dDZ
HFTLLrh5qhp0TG1y21dF3XeDInV7PRuPMYk4/BXHSr3HucRWf5i7wAaxtNuDueaG
O4kudHU3KY1Q5pZu3FYaPe5/L8oJiXVj0DxgsWSEQgG0kcbtxsUUxSwlAG+cFUhv
qOnWxkkp/QyfXvMR6VnGMGCOK0ZeQ7IIkMhmQXfOYXhvbQxf490ng/3vbfeLh4oj
vsNtqbIAXNlT+rJH6Yexk+fhcctx/IiwwzMSK1ddu9alWI+RsTit2+4vKqoNRpNj
F6CgoYY9Rst2uyQzjnWzeGTT2waaHtOcm3ap8WqiH34FwXK0JnVT3Y10wN9xs7rl
+WPWc6NxpXIaa3NC7EoK/6IxJFK/jthlKa9/CjqDh+SWKxsJzNMklLn6WsvUn51f
c/oqRRfaikDLBvaOg6RvqSA/ZMvmAtNCpHd3wcNznsqpNT1fTSXsIpNTqe5rjfrv
PP8c+6as53N5phjEGYuA6VJ2cS3mBVCnrifoyl3do5ZnUL0BPbhBEtBWWHGKb6Gw
rh3scdAN5NAN1vn+1uJb6SzvckRkjUHoiI/xWkhRf0+JncRDXBsH/IIMsWfdxdOi
pK2JzZnTtX8900AZr1utS99SI3+8KR4dvh9inxRykBN6bqDzxt2Vu/uq3uA5NlO1
O+jNVZ0G8MCxaaZ2E+iXykPCFG+fT+f+HpD6+Na7lI8/dh3HphMuBxKaqxlRFr8Z
lJHUZK7GqzBf+74VreqzJ2sOX+VCaiV7kwkkwol/nWtPxFE/BwACYMhSDD/rVRxN
/kALrmQ1+8nraeK9zDMJJOnGT6B7iR7QfTdZv1nJY4CzDh8s8jJpri1xCp9qlLsA
eUtMP76VCCIZ6pGuxP0PqW4jGP1X3+c2BgC2H3LkFQp8hrL/H8MSDecg+OdGHtmg
WxVXhHwxe22ijW4WXPNFQgbGhSj5/66naTAA0FkGkmFC2VyJxxLyIZNtVwjJbumH
QQ0dehAppKVDVHty+XJal/r6ZXAZomEqnIaTjIkm7enfie/39jfhGR1bExYzV8ok
SMOT4RvvwX5LVeDtLlp+YmGqRU+ZEba8S+l1myEV+QOrXoKGN8TufY6q8EoxYxAE
2hTCPx6M0kMaKXDPkLOT4HBbCrjyU6ROvkGKMUhCtUbmZtyJB5vZIX1Lj1ufp6/5
uQkzRVTz9S7JbbmmrfgDdK1+RnQ4+DV3DPbhQcnpEvHfmbXnrLwDooAq034gRaxI
fh3RNrEgdVET8pl/e2BFoSC+xo08aIQ3UeEzhl08jGjDufwKgoNnjt10gYmhn6mM
uJOe05HR0pdIuzcuskhbSRs9Ok3c2Vyrql93U4vj/PL/tWEexz4IaB/bHnKoenBm
qDdap14ZGtnxa+XqpgB9YB5M4oticFtPORLq7GnrjOfEcsBJXhnWyezlcXae4isx
`protect END_PROTECTED
