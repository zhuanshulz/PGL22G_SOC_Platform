`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CcORvtl1+91g1EYRTGywFuF73E97jBSVmwPqP5Hrf7096IOQdq2xT3p0couT3/cm
raTyZh8i9NNCPzqgho6hKoUcsQwKlut7WEM5odoa6NJ9hwo4uIr089DJdl6oluTB
4qk8t0CUj7O5DwdNkp0mzzI/kshTCywSiWFkX0eLP0NhHNWMtHUyY3LzCgnqxW6l
tjian1bbVFuf5RLOqvPvIRaYdZnk62m5r9ClOxgezoLcjs0EqtVNBqkEw0FFioDR
5DhW3L1sRqDG7z6eYRv0qgVR5b65kTW3cSj/p0mGf6VC0GQtN3VIowFBMYbMZ7HU
eKAtBVScCHZfo9GdtaqHAJG9Di/JeInCEERg4YjP7/9tRxJDrcQfl+I6clhf2dX5
`protect END_PROTECTED
