`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cg3YPi6Iijsl7zFfEyxGTfSt8TYl1b9syAPCQdeHiMvkWmee+iORGjoyRfwLM4HD
H/ja6+S4dulYuDVamBdNN2cepqbSmnVkzLpOIxavRf7ZRi3HMze5pqIqEJG+wfDY
j2KD0BreMMFne3wmEvnqpjPuDX2tv5eiqZb/PCQhdB3c3Z+rNuw7vosjbH9uJGMz
LScfqjDCe/bgn12AtXMitDlDe4AOhIKeu+GOBxt3BwDvWjGRICwSMbYEuI+gnvLn
+dhVjQSPdubXRMBTongfs5kQrPUHjLRKJ4Gfzne5djJC0p2nWxN5dwxZh6AtmDVR
2ct/0S7+oBVAxZoIeiOAmn4M7Et4WErRs6l481+Esa+bIva9ktkCBwl/ZApG35C0
ODXVzMqh8ME7yXNaw8O9iy61/vo1FwZ8EEbka/lp7+25uKOnPC/j1FSGmrrs+TlA
b/guanozZBHZnCYHOpRPjJ+SdNaAw1m2vKyTCluy3dQ3zNE/0PIcT3jCiKm4PQ7z
GPOsU3dlp9z3cuqMBSWOUnrQle+OUCS4J+HNTvgPb0AtDuiLr5nCwuG0dav1Tk7o
iKiHy6uSK2pLX4oLUu/Itbgl2wjQdsZki/dFfUzUgCkk9ZPoTIY9XYwBFc2EWAP1
qkQ1Ng1qAuIbuyTIhK5nW5SdRyDXYgisZSRXN3eSQGUGj9UqaXilHDidhNzhNb0X
W/irXwOtdcP2vc1Rt6zIVDrFOYXCjPL2YpWabLdjXrSxmE/KCogS3kqxgnz5j2GL
QrXuyPbfYXZW/XkoQ+YbzZvQWPmARl2ihMs6YloebfTh/mk7xVBcWrdkF26RxRuE
Mt5iL0cbOawOfDjGypjN+Q==
`protect END_PROTECTED
