`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Uwl/p28QXpYYKMJ5966wV/M6V6SE4Tgs9RZaVxv17kGJFA37391wY6db4o/y6Tm
pjdZuUgpHvMLvf29yTuNvXbxInnz5tkiS1rpnaOd+TU/DkDrmEySeYtSioDVG4l+
d/rzSsAdTCz74jccqp+DmX6fqiJdxYIJxQNCZ57xhe+Faur+eBd+1QJXz1Uw68Xo
USuh8OvpFVS+KoDEzCmKVhkDZ2X98kOS+ZQZz2W8pUPCSTQISc/DTtolzVaTyCf/
Dj61gyp0X1u/i8cA4LxxLAc4+JyLc4o9ZVb0AdXNtRny/xn/hX9smdk2BalCgUpv
ItzeHJCuhQkTfMxlVS7eKXdaHM02me6QW8MY4T5srVCVCFC3oA5jvhbj1gZcTU8A
q3rFtsAhpb8fXWgzXwL2imSphIuVGeSk23pjMDZ1/dtFzTomfMyne4DISFwGyHpI
cIqXa5V2S6CyyWHl9/E41fntDgq2O5M724WsQguOX7IlL8krLZSQaMgC0cpTP0fE
2+jcGCCCQ4FDHmuwPmBK6Mvw1qII4ybPuArLrvFsSteOj1PMnQ2ycdjmbJxnw/bB
T/LEu+8GthA6Vo5MJoyiP2SQXgnSTZil055mVPLLpiCVi24ca8XkSDZrG+1ZMSK4
w3oa/OThu9u3wqnBLVsHbC+3TgpQJw+Es7gR6wuA2y1kCX333l6rBnEsdIvYiGyq
z/Iuv2MwfMN1ElXbqLH0hNb0EUpTuzZj2lzpAcTkufM0l7rtyTZ/tPihnQd8gswc
YlBWfWt2yUVzhA2dQ1cn525tyIV7fwr7AtMOd6M7vMKAoNmQDKucQDFPo8xzQsOc
aiisu8yUUEf0rjXrjJ9X/MAhrQVe+pnPH43i3Cba9cttYKvIEnVG9Wmz62+t7ATY
1NSE+N4iCpNL3RTnHJ5heLSPZKIN04ZHkS6UDVmr2BhmSez+gaHm6uuT5A0o7vjo
qDJHg7NhehDu0Bxa3NnNGUiEor0AfU6SfyE4hnkyQ03XTbf4Hge91sdvcktTyP/c
9R2toXSyOjRb7xZ+r+8thP+J/ozRu5kPCWjD4CWI7SyyS+azqBne5ndUSj0+Xj79
k10sVk5jvmjvJUnhvl21SquKuIc4nXOB2YveFpwkvxyOLu8JzgIUe/DM/aXWZ10O
uXv0mrCWpaU3zMOvkcGGH6Fk+Wk7Vut/RZbpDlWupBzKrLneqK8NOwnPPHQew0aC
nzaowIkdOJdereUv2ua0Rq+SZhqzR/QQuc3I0WwpHuDDLbmQKJBXhK32f654RP1y
OgBHXNXwPPnNu9sfgNx+2uintswRlbt2IhRKwIR/p6d9Bqc4a4ygAp8abh6AeN2T
cayVlBRBWOlltu0t9QAV4NtM1dP4y+OQX7FNdFNqx3SdoE0tK99R31q0XC1/v2Mt
JvlAPfEzSNRfh8SOMxeQlTYLAWQtEh21smHR8COLxI46v4SD1GStXS7jVtOXJPCY
p6ipmgkRjWAnv1LX69I+t4uyUcW3raRYu42upOvbxehgwBTJcb9oahjZPsu2nLpB
oJ9DbEgePCB5kYwxuAnckj7xL/NYp/pvIB4EFq5givQdgqQ9TV3u3YDRRHeYmgks
nSNsRPC7XWo6qRLxH16HhZVIAGysCNEkLF+6YsdrGB30qQkp3Ees2Ieam08l9GgM
339NomVk6xaOUHj7JZ7yAexDlx1yAv74RCFMxtsutXNrjE213xPIVTb+S6ZhSnaR
myNeO5gTGkP3FsB882xS3gO+DDrmiZuLGYyH/zkC/xvSSu/yJDdse23jSTpbtRlW
UIXc4wsz2YADZ1Q0jbwOViiH3wS5gMXdeVcFGxVVtt+ns4dCHlgOkAUrGq0+FZbq
JY2QChVRy4xy0s8N8Eb/nR/KQh2iArfPAYS5OJQXiNuk2Q+Q5ju+v5cAy4mSbVe4
+ViOWnhzwOLFQ8bo3xL84NJgnprFqa2MJqRz0/PZadVprJAMJFUHs4GQepwPlURH
+ZPAu3Np53xcsM5tcii2GbDKePoZcJV6/fUmMpEY+LEQbrKTQSFH33C/7S/iSVkz
tiZ9rsHAhOzJxqh+qnimtmAJZuhjsJunOKnXYh0yk19T3AO4b8Zu83pCPi457JIc
bc5/eBI7M3rv905h29b0hfwL6iHrU3FxwZWqb6FlxdFavc0njUvmvvSbn8Ui9xBj
0qyaanroH3TAABT5i9cNF/q1Z54A17x5qSx37CtV7JnUnOa52dAmYIihE613jylJ
i/FKLJll8UDFUkPTemKOobzun0ATKL2i63VCipXoCsemyVYrPkcLsxudwCclHM2F
LewS+o1twG38K8CYzLdDRuyjvF3MvDePlV7v+IzCYhAbfiH1zQ134M1x+kg6lOQ4
/TT+rm7MZ6SOuIDuRjC2EkRDgCzdcsLyK8QaZALCuChF571kF2yjALCnNGwiuH8X
r7VG0EAEOh8is7FgylYi9b2iZubHl2rLj40NHg/rb+U+PaHSgYAoLPvPblpynZoh
UHv7sSLQCPAXs3A26KURngLvhh/F9aooYFrUJhjYKOhZ6X8LujQLEsvhk61ykVhf
/836onOGMpsepryMPqiF6OQ6jDtmicV22xJWLdEJ+pw=
`protect END_PROTECTED
