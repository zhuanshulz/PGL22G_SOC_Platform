`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9Kl8mJVuKIBGSfDaBXRzacsYFG/bjUq9rH6ub7G+W++33h5vMA2ig06rFKO6tuw
DLLxPEsUpd0FhlzDOEH6BJJS6b2eTosfLD6Z8OcBXfc7qVlB/BJpdPZcpYahcC6j
/VqISav2ZalTaqhxW3G9fOhIjAtx/XTPQUCZ4wwXrMcrIN6XMO+SATVO2xRCluz9
5vKX99D8gYnfK5WeGPXQ8oAObs4SFtKGZiq2KYexKYKPs5pfdU85JqV/uQ6GWWI5
v44D/LXH+YIFjNslxXMdeHvpdXW+A1WSbm0KksKCT34Sx+RtvbjH2JJCu4VKjtdc
JAPqkFNNA2dZpp5x5mbF5qBZB2VNep1f4E2YHPQH6SMCpV9owaAaE5vzbgoiBg9M
SDAw/phCp2ie/5TiQ2Krs3byNwSCBel1P6/OQRB1VjCuBTiL6767Vhaatx96mMjy
NiQhAoBxlRnQqmOK6p29blV1nn1bEuBdy88vrwYXjib4ajDdpCMwiwqv6NwzY+2Q
hJ5OE5LJ95aMYjwIIDdwbmhAqRgW6sLGaV19kGkAlGk5rifNSnWq+4YhXG07vuD3
WPInc0oakb5qoqblDw1alg==
`protect END_PROTECTED
