`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Amkqt2UDeWqub8+EMbPKrSDGu5vOu2sx6RWUBTe5svje6QUqoJfTcdK5hSBXZ8cV
b9CTsznjOJnxglZqGBquSmhhvQ11/5z/zjZvoJin/miKHQT8/OQ5NLb7T84LNZDV
jsyM3YxwFEpkTG8tNKj991eOwDkZcMVOJmL4cc/q02LXEJAtS7YgyCnY0DxZBgTg
d/r5yTQoHxnnIF/eXrVrQPCtpavuAND4ALvtN1C67lRarolxoJoOaH+13M02VnFL
Qsdwm938ZBMbC2QdTCen8D716quf8EDheWarUDWcYMjiCbN/RwLIK24ebCwK1kyT
Y2ZruKbetK4reTI2mMZoIm+l2wintfbODu+Hht7KnwtlGUzfh45CCnBwRcXBimS4
GJreERgMMvs35t4A3rpJnxHiXEPJF+H3gADejmAWJbR/aXizRx1TxP4pkTBmHvjR
1xdATcaFhOESg/CC6Si2VXzXdA4Y7OLd0xMeF+3UVdHJgMXEuVUA5uidrmp0edCg
dZDRnt0cmWUQ3Hig32hnIm168GGyKxmxs6RgrcCWeFlRMlgO3ftW+nQyx0EorPKM
gpmpF3feG3hh52BzCwFLT/AFiwuQWfY3X8I9w+9WoJ1QJigtKxe3E0Bbsv599k1r
NfwkjN0KZ0IwNWNj/+UHlXOkeS2jrDRFBvVfU9MGx7gbd0vR4l2xwhyyH4c0sluB
zMjEnw6AtsEMWQz3dqfM2dRDQib7NTOCgg4ptsE0jxQOGJkknX/dqke2IEMPa0K4
7/Zv1PJ8GchxYf68boicC7ZaxmQnf+hN4yz/7m977kCXFJbk7SgWifRQkQ8kJb6o
k0ZXu6bSX5rny+oe+0A3DY6V3mEqXWXWPlFRDQFg5CkBW84bTcNWuwUBioK0su73
Tks9qgGT2DQsoz87s62EZbTSQYdorzhhoNnIwUShK0ogYeUd68xfNBUOR+9EmoLP
Y1H3qb8145zAeUjDABt/bKd2RPfchJG2XJVZ7mUd1+5nRTALbirWm+x/Z+6msTFr
`protect END_PROTECTED
