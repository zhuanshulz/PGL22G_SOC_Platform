`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3cMn4wGOvoln4qtObgYck+Y3nlX6lceq2slAa8p+V2iU1zip5Iap1PNCrnrlEVM
cw7fl8cYsQfiWUCc+XoH4FeOCaTjQKyYSsMgnT39fGQKeGYKat+5pDD8q+avm7RS
cvo7gpxiWENw6vyYuEaE1/SKJuZgH5QrEtBUjsaedaKGEyuClUor5qCPsBfwg8CE
lyFxNmoocQZXje3cZ4/u+zrElBOkiMQy1CZJ588WJvojhxLbWLbYlzvJiaDq7Hfv
CzLeOT1r5PpDoojz+T3YkLgjLi14YAyT+RxFxmzvEGlX5EV2FV9w/aZbCwAHK9N8
4VY73gAP01n46E50q7zXB0LHcRhfnVZc5QUVIzW4ECZZJ/PxDAFC+R8ofO1WnTtJ
NfkZF/DigwFaUv0hk8q3iZ+M+vzDijKnjtoEziD+reJGkzfhu4ugam98YBeWYqMA
J/Wun11/9fLthgiobOpMU6Sv3l9r2gX8ZW+1r5A2ZknlyorL1xiotb/EcSbjZ+tk
70Q7VT0RJ0M5iKHKMVTJEy3XDp4BRaWhtJPxdbI98n0/dh4TK/pcTdOkt8azZupB
0hbTM3Ym3n6Aa0T/d/nGV/rN115Zl3/XXH3nb4f489XqkDvUPQ0UpygzUZqVhDTn
Olculnv54yX0UHiXC90K40jXIpIOcHI3sKkfbR4tx/4Ax1Q4hgnlFpsHIVKAFxjQ
MyF8G152hsMZIc8SA3vZWtULXHYidjczPancGD5PZ5PIzKX9KnTCLXE5cKa63OrM
JucWnL7othagvDfeGWaXBsmPVVnzVf8caUoEETyzxOzZ3+dXF/50qpmbEqZq8grH
/YZJ6+Wm58KmHfXJkNkkH/2u+Wle4fIt1atof9b4Bi12EMYJbf0bBFYBFQJzT72R
h0HdAIKngsMosfKqyA5TI97p4gPBCcdIgpcfg7MLOhF9Y6Ldpx6HHbjfWWdzO1lV
PTGKHD63A3lXb1OGx9KdHt7z9oFoejBtfWwk1FCIxaPN0feyYuC6WJ8MoIjVGcdL
f99PWg6rf+og99Q4YdpUwDRNrrrEXwpVeqfsyphaSbDSvBcNnudQjV+M3dpS86Cr
1y38l5Rw9qHFgZVl9q2a3mDbx0rXMUrl97EMom4MBh22E/EbySXtLN5xniGSCgmb
Py/aAe6HXQK8HznuCSaIgk1wM0t+XNx1pnyfls5eMRAMCcHkKV6vYnTrU3mQuqcy
AZBPN+MfXhhwoeU40XZDnKZeW5yxdLyZIylA+i6nNU1+XvzSSdGYZBEeQN3WkiVB
K4UvqXUUJrHWj7ZvHshxxf6hxwDL21FK9elhq0hFFMG3MOfPbzYrBxK1KFU1Tf3s
9X0spRIz5NKF60tDC6b+9AW8SQUfNZTqWMX51lhk/KZbb1B38y1FDWa8LKFUNoBI
iIZNWS/6s/sucb3aNRDrJaZb5aP9zc/IbtXdCei1K5J/DmqCm3lQmBT2o9DW3vqC
1Y/a3cMNuJ0YpgZGAVF4XlEJA3g546AQAKPOW5sHDsWVvE7J3JpSyY7PjV/52mzI
X59vzIF6HN6ZDTzVKRlFEnVxXO0A011gEBRmKJfeDuKJOK/7+lyXAPlSdMUYVBaH
AZiNKPlGthYklEITH3yWMwN7en6sNNI128RIWM8RLPqFIrHVANnnGbECWI7wLtTx
in9AQM6dN3/bj+nZBaJL2m4d6ULydb7HoJCKYDO3lbEHvr7fRdgFQ9RrBXaAdeFL
B0WjgpEf+TVWVEJNx/rg9xtqAEcPVtRkR4RrkKWy7H8PSFA693j702k23rw8YqUR
VTpSSuRB905VkyUTCXRXH9pOkT2eZZiRLxD5+BGqlZUvoYRoAcuJZvZ3yxTcBIpF
U0I2bzyBlHDJ589336vI7AgyNLESFZLTt2g28786xF+GBhOonbgdioeIwS8IOdUy
hBqSc+OW04W530Ycl5Ub5VoL8eMNJtdIXaigBaiyO5vBLYnP9cl5YRksdKQ4+3Gt
4eZE6cdU2QYXUJh9veNFyf5bf2hGUZ9NpRPmKCJ6uXoVpfDcl00SovXf3bhS0ks2
vP+NK0VH2hz2ecO4W4NzVuKIOK9iSwcMOFahZLDJzdAXjMW6pZ1IpBLbC4kGXWxh
cYTYvLVDOcyZ7ejGF7e15gtydJDypbss7tRf33uQ63iwkrgqT6zYHb45dSiUiIhC
BVXcxk8DIns3IqndwNGrM6YGFpa2o4CjTP2JKuFHD88QGCnrxvXGwGkRolALau0P
xL9dmFjEC6CTr0KMtWex0n5U/e/hc/V9Chxnm0QevYGF+Kxfl8eUOcIFgco1A4oa
AO0Mo6lTqGzxh1d50XD7VIQxlZV1HWN3LqB0651Q+f6W+dI2/KTzabgKXAuLfZs+
pBenBxFpzareVADPeMaejw7eURHcQ7Zgl7UHqtVa9EqNfj8IxFdmc563GCSNtNiu
NWaAj2mMxCY7JQxN3N5zNHxLo+ffdKWxBhLqtF4UeH9Uql2BHd4uuKuYqhDl2TGO
jwP20mYa4v3O4ssB+VNxCCJgL6Ui1d0VBvWGLPSwWCd70wcnrREi9HunaFMtspqs
FGD9sN6w6jsg+cycnXCqcwhiMiqS0rjuEikAO1TUyUIgOmMbzhnGaPZ8cYkvjz81
GdQQTuZp49aBT5UcDNuaXg==
`protect END_PROTECTED
