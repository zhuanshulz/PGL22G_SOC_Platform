`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DyJylK/luX/YjkJE6pvofMnxbe3ON5pOtXxDiOw9ApnOh2ekLsikZJkyjxqKlaXU
3Hxd1YpULe87HF3qdXkT9ZvPVBSuJTcTXqUF6yc7LcSORjzPxR8Jq9zAdGaby4T+
MKat8rYdiGUyrwozP9Eb23cTcPh7qE/dL9udNih4JLDHj8zryYUTDeIF21X85CXP
SPAS9WL6tCBYjpQnz71JeHQFvti/o0CbpMixUYykPLJygyOGjej8fcTqQTNWqbl4
SkPW+dNWtwPiR5fmjjurydh7UAooOyZfWbtI9vzYvIn+QdE2QqutlDDjK4WwlzZ1
1Mc/NjUpyayq21NPp4Yd4DIT++Uw4tjSXjrwPD7DA7QGE+p4AxAGk79L3f7zpfnX
mS6xHtBSDcR7Y6PuYdRxkTSD2j02gvMH29X9KGW+gys7wJ6xR2kOzk5M8GeBjgjM
c/hhD/y3s3MtkTMj/eoYUWVgsflIeKeaqbpHhx4mjbjdYjVFm60I4OYs1MKWluIT
Cfod0hf6M8ZsGa+Geys+a5mj0E+mtOsKEKEADKm2IO0R740b75oUw7+eNB1cIAbj
QmOIxpOSRv+LCl+VkvAuf7qpFH9shJ4ZSvJhs2pqF1tMJw++N6tsNg9Pk1cnzFQH
7kNa+DsjXHqNs5K9Sj5zBeYN4E2nnjl9GYK9tcgvZIJkaCilzYJIPXNhRmLBR4B+
xRTZFhfT0z6HjZh7Ty7Zp0Jp3euwW/iI3FCyJesTDtj2eMh+FuldF+0cQN3XMCY0
PTd0mHitAnS6WLsoq8j4g/qwqZMWMfjztAex6fH14hoAVRIMCq0ucLSsPBR+ic/v
vjqUNwRelHw1nfClm/QsS/6OF7BIWHuh2/eLachFxy1GpiDs9sOmhibehvpKrL5N
enza5X/6ahLNXTet0sDuIuCCvuOJDjxwmFjEJyuV/gYQO/IuHmD6fgh0WlZ1wmbT
IrWzp4MXSMmiUtLmhy5LTfJrAm4vQ8FhXoR+SppcUER9KmdmuQRcpiHaeBN48+ht
4Bukct1lVbkXlEvAdtcUEnX4a2qHoK8BDBGUQcJkip7tYIHXzfg60WX+AzY1d6tc
nFIJr5d3AkPptDJtNREyrIhAjVlBXCuZ7mK4owtwUm6QXvGePLgULA6j3YjA/Btu
uP7RAKmexNA065I5Cw0tC1TnAOZnABNb3i5L/WnLIjEu/hw/TQYE8Q3bfiF/EU6V
1/AAVePhiQBlaHPiXZd/AkR09Afd863WiYVGz2M4HJ81kPm7m2Bg9H/4yCsbJjZO
iimf91lNFsReUbDjIcZvo3kieARkhDNNXph9ui2YxlGtuPPTFXa3bDE/yhaC97nK
igt9jQC/BNOEELDtdOkoYoh4Ob1UTlN2bBp2GpHXOqGdkTBoo24zVAMWzu23noEv
onlnCS1M6hY5ua0FHta0f4XpSu71xSyfQEnulaYu6p5T5Axqet7QWionmGDmBBUj
zHaMq6x6AaqMcgcabaPaWt8jDmbGgCaMKTjTLBh+z6kC6Ff6sy6Ajo3Et2WZWaQP
tJpWqDIhI90WSNDfoS+NyKncG5tlFW+av6WZwzgmP8tO7yXT8pJM1U45WSx+5hOI
v3YDKzjfcSZj4a0SjteK+kIx54fBHB6j5B/yponS4IO++7xx7w3AiOQ1lqqrfwWt
9DvbYgorfYraGYaduoNvh/+fqHvsm5AOjrjboS1+Tsk37tiW9SSA6FhQX4+Waia0
SpW/W/TdkIHtjng1q09Us63HNQMs/EcQ+f3IW4bHMO/92p0eCKBIfkPCzuOggORM
ATma+Agpi2YQ4MusmVo/jWOvA2LN13oDT7vuSIDR4LhDrdcigJGyV2vYWWMwpMVp
0A5cTQQend9UUVxn5xmdvEF9ip+EURmclS9j8So26fmsJ0EyduW6SiEOINKfJNPk
T6nP9eM/80oep6MA2WRSk2O8UG9PJphMfR5+QofIbzq9o0qgYVqC6Ja1b0lc6cPv
yvrK2Bpt4C6LSqJr3ZoWXQ==
`protect END_PROTECTED
