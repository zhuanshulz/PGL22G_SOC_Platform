`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1v6CWxPOPMixtz0+majOTZ03WRSNDCuyXV2ARuJu5Z0JOAqKDdgyocDlTqjqVZsv
XLa1uVBYbyWHVNZBRjQ4ObTGnfF9UFe7erQhz8m+NOa1jQshjTMa521bdjGuo9gw
9E1KtezFYxZjaF8fd4Wcx3UCQzv1FpiYgXG5vX2FglyovPNCJVY2s3Ev22zu7SX1
SJNxKNKNvTcGrpPufhEreSvyOT3seimZBAdbXHy8FnuAbyLk2istkNx88vLpH9eW
vbmZ6gr2976hnJzk0U/Ye3+QDPN5ka1gwelLsP6xCq28Fpevl05SxVLnNA1MEWdz
OJHZP/zuUQSAFIRNsvfdtQ==
`protect END_PROTECTED
