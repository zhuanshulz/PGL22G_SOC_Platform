`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tb1Vumk7db5g8hLfRyIqAV7k4W3zqTKja1SLKyX0RB+QwdIOfVAi3vZUER7Grrie
7JW9IqiIWksziTMTFQ0NLzGdT9L++COzFtUMTWo+CNh9j5CipKuhYiz9UBB1jiFZ
QtSAfYBHgbsk9xsh79woDZxQirOqXHs/SB5JyLdOdE4UM+xlu+7v8SVu8hjryHLw
je5bbixqGgMfbrR9D9DCmF+z5AuPbXEVfRdiB6lkLmOjOeeVR7YyTRyF83GbPHA4
O984PrsxNvQoVmWH1KehtOs1G0mKbJhSumZtxY56HH+FGuy8GNUyJb1US5MgYAaX
FapiKIWKCQDDK5GTCO/myyc+O8QdD4v0OJJrVltOb4uMbE3AWKBY30b/Spfx+b2R
qOHeyI4XMHhPeBC0mmh/n5HdbjH8mGnH00nRTkz1MvRfxJ+BtB+C+nV7b8rQVGj9
zdgageWuTkDp65jvCJZL+Mtgu0ocfMX8tLKU0UGfbx+kfRCfQ4SWSAiQMGIci0OO
Pd/mipWbFqGcqetwHLNyvLHUgDLojJsR1p1N7/95MBJZsj4WpETZvIT8n3VJyqGd
rJFcOgcHOeh1AZq0vepbrjB5FpcosnDZ4K56lhAkA183aiKyMpLCpWRXk3rD7UDn
GuqdXXUZIUIO84W7ttf/ye7RL8UaFb4SwpeQ3rPXEcojoJLOl6narFeaSvCotEsV
kZxvIUneomqNU8LbRRXhxchZo1mXtkgRddSxIy6fWaVOEU2g39djIOgxJKWH0RJl
bJGIryd6UmvRXeORiWpuirLbP7WyyP2a8qcDRUl5Rz+qKt9NCL3byEdMG70Imj+/
vc9AbtDwIgtw4TM0VNdB0R6emWKUQgIDrde3JyH5pkyZkM7/Gtog2lOMwYdP5Z+S
3d6q3rhciqb68iKc/ahRHPKxDLnhQ7s7LHrJa2yIKi8zvodBiP9xpDrs2sPIKJQb
ZR+QLpSVbgmu3f0X4XdY+rBWE8VbuEcl1X9JH/1kvWhrk/Rn2aqAxsS23EOW0IOE
F7ilIxN5NLzONN9Nzm+lMNJzSyBG8x3RFU/qhwRyx9sPY4KXgJnN5/JU/K7RSsb6
0MXY2ZfBZQ5keL5Dc3mkwr5Ual+D1MIOo+j3ODsT4YjMUx2ZhDv76dH0xshZXKQn
P5GIQ2WZh4scRvC34Ot5UJ4sbQ8h9CsYTuoYv7E/I10GCO1/n2mndKkB6RaN6Rku
kl/TAHALpy0W9znc3BXfx2jNYav9YFaBvyXei1mRDKx4YPGfeflYJ3cPUUpmx6ja
WCm2Hj/ATjpYO5m115U5Xe8hReD/3O3Ux8MJPZ8W6uk1Ol4Wp5P+nLEr31ikcAw5
jWBF4mpNgQF2R72/lYBKCgmY6uG6s/G6TKEy6hAlv5fS4JPzge/wR09klxeNCMtz
R/nrHNGhTClEWEwlVrpYKgO3ntTSwO7ShAFMcPAX5HSTLkADs6GmU4BTdeZ0pYLB
UFtEVli6uNwmSa0NE0X4ESFIMXTIJUL6pRH7O5y6TElN4goNYSs7TCQGMujNtJNI
eyJSIoq//VE7BLG0BE/Y8p/wdF4HQ7lOg8SPJ8qaTPmxR7QlP9yQ2VAOKIfQw+YA
K+BNx20zXt7GKH2YceNkkYHgWqU2g6AMT/Xo6TEp1aSpHDFS65uw5PGBeM2UIAXH
pAKngNfOonWgDGIvRjRncP8S1j3efO4TJrTbjIi1Mu9hKWvKVufHDblNF3cpEOsT
B8bYZGBeCTcHU15RONpUg9v+RDRfhLnA3uyfODLD+BSHA2i/RDH1fBolZV/BJ+3y
1niu1o3qIDPQ+NyGZHU+ziz2vLNvnAI389CjmVWTNy9D8mWDM5zFrwq6e+5PzE5H
0imMVTVbaHs0O4fbc1JdwO6OgAzVkEsKAyPtax2MI5/y8QQ2AmknRATIYH5Lj4Rw
Di31QLMJKK7E85Fg0i+GjHR9XnVLcEe3yzdUnjGLDHiIln5ld97LE49AccmXciRH
vmDV4tDnFEELXW7EUp1SprjeRTy4SdAnRZ+GpcVYIhmHjrGzFJzTiSccgK05Tggh
iN9fMbCRtn+9FIOajp+dWsv/nu9o62MPV+9twddJwL9pkiWu3C+2HejgYl2Dkcrb
NrOVIgMdZqWLBsIqi+os/YEhI6r4JQVX82y1CLWIk9jv5UCGrFcHsqif/hIalRwj
dedTeahnKri8jynZZosABS4hrAdbotXwjeJZ7fDowkRVAPiIhaXxbKVu2uakPN1f
5yHUMZA9hfoKh6RCoLDamBbNQhRSLxxMjzSK3WBR2XahbPA/SVR5Mgw18/tk/D7W
UUiTa82Ov+I23ia1/kf0G5bDpMLGhsoTtzFN1Zxnf0e5OdKdXspf5gRQSmeSQBFR
8GKaPnolePKWFxC7xWcdIkeXf5fdb49WZxYjzYCNEBCrQeqFJXrFbUFfVN9Zj5yn
/NvMs7EFCVh/8yWvElP4fH2Y6fiGVZcrxas7k7rY2zy7TpfQ2BzwiEfytZb4IFB6
j8RJ3oPOsmeeGNSoYpGj4ykuLi/bh70wdg10An1RtC4YphJTGkRsxDxQu1hGTDq/
VZa8P6IPX54Rcigbu8NWnx+4uVHcXWledpIi1vqtj+sm6F4GIxnviIUmFhoRoZFH
W8krERAZxlurJkezKGEau0f1W0WgrHcJkGJnst/gJ6PcrpDjwgzn30OSuoz7YkCj
JHXUt7WzbOI4D886rxG43GSZkmr1Nk1Eev3VMjPvsPAp6lKeQ9adPGH+DrStdvyj
PVrtnWCJGHtDb2sc9zMtREVg4V2kqkVlbR4pF6Lp2RzVnTOWFAy3LqOPBprJ/UMi
0V01GPtcNqQeNMJYbyCAXwpDqIc/zwbbcRyyGE80t7LD6MmAkkD68PG18uMYtT/c
2M6SOSjNdzyGyAOxNAYlliQMjZ6XdOXn+2IwQCll9AZSH+6LUVlXFCz0400soe//
tAN1iNKZSy6NHYJlqbRnJEbGlFuGF6VuaLepq//rOL+Q4BQI69DxNvDkXmXm0aDg
4zXsuH9S1ju9IU9OoOIoIg+NUCI+gENXGoWI8p1dMyBkNpNfdBOWstLEhYKisDfz
phoo1nE+IbPq4yV8qWbsISsG9HEEjj3XLd6PVt0stYRTlK+pez1o1+RrzAsPia+E
/01IAghiEnNYB7C2tigVfHjRsaxv21u8ol9gF0rrVn8ZaNHBVJJ9c3j36jPlvLds
tiyjJsXQmuc2eDjBdwEkaJj3ibN72zCzqWHLz8X+vnVyWjWQF2SpTXw69OrNXsgV
ljI9duwvCodSi7pDHlRYl0gOoqr9jslg5TSOyvtA4cWP8Vmt2p80j7YEfqryc0Gf
4PGEHeotUmyQdamn2JgMNLwW4gdyw1ZDCRhH++IF2lkq3BtR03JZjtusqlhdX1lY
bnRQibUx0lp6djVBtfzyl/99pCrElmSvE+1d4XRm7WqP2KCmSDx4MSzCiYx2a8o/
trC/znAICal/snJ1mPdMPNCcz6JXa+LcJtF9ZWxcNLw=
`protect END_PROTECTED
