`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfk1/AgBahsgG3FP5Kc8vgnpIHf+PWmSohsv/DaZ6XWPYNryhMRm/th+C9jGjCRF
UplozG1blCOv9JTm9dUUcYIv6p9C089K+fS9/ggwKFLUkV22VBBFRsGD5sBu0kWV
9H0hURjNX/dOBwYXXRSWfvJqpdqwCty9v3HDDbGR3zU0sS/Uo1NYIHGqMbQ2ATYV
YYYsUworVBHSDjY3hzR8xtKnygVUWpxtTE0zjVTyQXXkuuB+yTx+KgGd31Ktzlep
J4bqkx2H3FHkUEzZfunD0fCmegPjIzG3XjcfMr5Utgju7xS0ygM7zP9f57vKX5kN
qBJMicyVIQ6CGGBsbDgojEuDloXvyPy2mfMHpQZkOqqH/iFFR+8W+L2PXB5rsamz
TK60trket9YnA5TdV2YmpDbNKFket0iMkwTfEH/DrrcNk7YtbHroSj94QMTD/R+J
cWF0IGO7P0b8/yFpr4bdYwtwI2m178IoautLSZYgEciWIuXgH8cGshq1IlttNccO
ksUv9Ri2O8uEyrd32w/kXgZ0cgVE0V8VsazXW8wvrsEgvDwbPy2LGxbPMLE1TRwP
WBgjIOek+MQGBQ4pUPP8j9hXV/zPBzKXUpThmO4N/2Zaa+0q7La2cpQQAHCpH9Gj
iCQLQi6y8CaPqc6GH45nA4rYzpr7rz3KUfkoxN94bTtbUFdLWLem7I6JuLJpw3Ut
u9rjtGq8WzvvFT+VA2FNcKGIpMIwkv7k3DfRhwTt4/8k7Xe0o3LRlNWUZ6/lrQNt
`protect END_PROTECTED
