`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dy65HbgN7X/ZpvD0JxCGPNGjTgzYM7ZeShNXCn5Rn6PBJ1WMEtK5WdqHop2S8srU
aJhUgWHQjCrfIhcVgRx1apZT73P2TZtCi/2w7tyDT4mWmDD4VfhoiLFrjEEkRs1q
zZIunPRDcuJwBAYCDdijTr/3mxulXzrPUXAXc18TfBgRYoS9JmRnObrR1yYJ5fg1
7hLrYd7q+4ADuwcCgIJq6MKZ+kBIUVTZQM0C+EFQC/6c2PQKwnN2r+WO/NbFtRSQ
AXFMNrKWLs7WcKyQmO8yA3hJY0+HjFa3n9T+xOkD0ZEPsOA9S35EhJOuFro1hMwr
q5xJZf6n2Y/1zwdyilXTg2/2eLiYjHr3dKqKOCO7OQrKYFMGjmBF4O4eDRHJIiKw
g7vVTaLd8QHZ7Cndkh8QLUQWr/GIXrKUEl0fo8nUdjc7xbJTrVbnH3FIorp+3NuT
gGIWYujs0/p95zMuHrcvr32a9BQ/YH4rngqOy0AzhH+v60MTJio7aiQayQIfhl2R
kFWtRJub2Ucz0goZtR6abpgCVaR0DhA7uPp+5N3fm5ustm9D8NxC5tvn7109pT3U
RNTiNG5/xnxYeXpwlS27HkUfzY4DvR+aJ7GpfZdJhnTiKhaiNNybsxC2oOIKvbzj
n6YAJySbzwnPdEHZa9cQH/skA+Ne+WMGHFoYIt6LqlQBqLXGm3+3kREMWw+6sD7f
Mn9IzcN53T/qRKFJrW1GU3Wd+SBEbTnwhbd3B6wY6DJnhJBVMP6OoHZ5RZKfF/K4
LgUqPo4byyb0RDypolgPVw7T97bZMJZ9kI1C6rIvA+Cuzmg8gNLftuFP0vSNujZD
batPHr3P9FVCVCodXcoPZx8TrXW61QzPG1zJHE9rbdjy7LPzZ3n4w2XRHezLfvAa
`protect END_PROTECTED
