`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GyAKlITgFM57e01yGoXNHEUhjUkAwwWptbCq3DRzjXmtm0DozUqDS+fRIOzv/WGr
c0WfVlCY6bSX/DRqCsIU5jSI50p0Babr0NsGibmemcfuGJchFrfIJIn3dfRhUq33
BNBYIT+S2w4/kPYNe8QH090+odcPEd0R+3PHdI+/ZDn4uMu3XjVP5s/d2YnTZIr7
rcEMdK2vq9KjbMNKe0y7Ga6lTuTxmlZwyqJZUA4X9X2LNCqRvQwUPDnSoEznBCFs
n3o3ifBsSqS1cfMsLISHmiXp+16ge6wY+0cxc42WbHqL/lr73V2aNsJoBpNeCt0C
oRTjCFS5Hn9/1wS/ZDZ0w1tmX5Futmd7dlTedsMqWAW7amJ9AKCAdE9J0DLebNIh
7ks74xn9CbF6ElxhFMbg4uSTSTPyAxrhnuagVsFoalojUsP6LkZVgiUsKJS5f5H/
dNWfRTs57ciadgUqJJOVERmZmrHcyfdFgnekgAVVl3C0DwCRaTvV1SaPulXu8l0O
TKSWrbw05E1NVnRv7GdwbM5wFLgpxkV2wWaReRtcaYMcqR9Xmli06Q2jb7A+Hhxn
K+N27Qz87YiXDgL75Tnki1b1TN0dQ4990w9O8MkZmXe61qyjSeoXvy9W8z0uQmB3
C+oQRI3iMC6vQWX/IfW9RWT+EkPBzy0CcH8jd7nOLEm6lGWBd26b2Jn9hJaKzjKb
dO3EfLWx2qFyPWhv0g51Ax8nc70qiBbz8FwQkFxcCDR4PwRTCEVmjzdUobcLoz9w
bO27OJ7nmkcpx5L9xpxWju1pehRH7gJvmJJ4m4w3scYjliTw6Ctl5pi29XqMR77G
YbVxPWj+2eyr/ZpIjtgd9Ixz34XYJNervmSz9KLvcvbvCybpJMOoqdYOfXJ1CO5c
jB1WGaF1EWngi09u3gtKJ20c2+RcbRJ8CgCZjpx+TccnViMO69+iFoDc/74CF5lR
yL1zMYyKBly5giY1neHQw29b8OBUfQInkmvN49QeCT96dZiMHmGcvfm9j2cZNRjO
Kg+wUbPmHtqvScNLSqz3dHSMJc3Q857XT6ubrNMvblXizafP5sSUi7WoruyMvQnB
Yc2czGc2ccuAMIUyjO10JZ6fL/os+xTEhZqt+xrV9tFbS6Sh5QuPemLyftxAc7WA
+1oohOxk0DxIRmCKOgd6AbFVXpDoEHfqoQ1B5shUebBHyF8Gtu88Wq3fBMPcuSgq
gIDQ9eLQiY0W7mSrnGM1SgIvkJVz3YDVV/bcCRMcvdhRadWdh6cDmxDnVYHx544a
cTFjdDxtk+neQtC4bl5cNufrYF7wKxPDJcijv4cveMpm356QgrIV5+iKmGcU0Uzo
63JHMb81Xyq6Wi50DzP1z8HvJuewKiY4xQpvl8JwC0GbcNELhoAskRLSdITnWiN0
yPTvcMpxhjc164m/vLA0HBJCfU4d5ym79SyZF1MBatfphsr3z9vJlOsXaYHVBVYa
7VZunCfzGO4mKyLyIwZHuDvthRB8eTFg8OK0+Ld1spLdjUEuwDWjw5dTvpqJNwLg
mxa3LvWUOIdcnEvgMS8WV8onKhacN3ApsHbyDKrKMsHAWqYjpr8wY9i+vwfn59DZ
s6r7WdR7DvEa8hmbxBPPLnyTrarvUuefKHwj0XBTuknDQzS3K3Tri2c0wER+beIC
YsciRVLJTaAYSIBv0kjGYM+Lwv1jEP2JR2/8PXfBtOqTBpu+rVAbbL3WWDrn85oV
M0WlNY1JSXpEiaA7k1fLsACYxmAkdMJRaaGGvZ2GPm30y7bD1/n4bF26X2ZF4R25
RHW7XSX/nvpUDzaTzH8WI99sxHB013wNLsCD32iJHpOEbssqJkHke2M2KuT7zBFd
gtF5/GIgdlLZx0ansXDtFt3YgZvg5IUo+cZFiKWh53nZBWidbR2GgPAtOA9NpTMH
VKbN9FTQu2tI8F6xUnnzoMPr1Mzma1vEZqVZHvo5cioo0gv3abTakCxE3cHfnjfk
jbkIDFIapA8EXmPgB0zAGLit9ux3o421RzqptA7HyZgc2XkYWx/P3/62hP99Ry4S
HlyylZPbyXr/iVhZgmuCCI/W+0KHK9ofhtnwHLyWkCML+k5CKKwYHZXwggDE/otz
4V/zdi5qtuK5wcigPA4cutJ6rGkvSWx5GZywm67rDR8xOpI7wW0JV3VF8wfdowTB
pQrCRpLVilRpanUKjQTKy2aa2zFyDmoGC9YicKx3GXAYZFBCopsfrsgIlmg0YADg
NFeY4wrK2t44IUupAGxwdUNiCIDwV88RT+S9NQUAGtcwLA9cpt03MpfNxCGajgfb
rAfwK+iqYL4dXK+JJ1VJDY8/jZcOR66YHQErvkLb702M2WLA1TtHZupeqT7Jg6JK
FnlLM9W3TDqBZWepud7IOOhycMNF0FXO3fXl8nwKi8Vaxf7Kz5XlBA0qa7RGpkIM
OHbMKgLSjnqZizXI0PIUQgwy6aMrRHZ1kbKzom5Z9PFHwCaO8zZBZHbHKSHP1kNB
f68uKBbmcS5C9f7+Jooi0URW7VHEunRbxrGzfXEIYTxB3D6abNfgQ7zSVj7vUv4f
8tJSgvODG8uP62+yPlaFFXcPNybUDgRHwCX8QSXbZ4sC3/kDq3VVvPO/M3yTb9vF
hhjn7C70QEZwWdoRt8A5mqzH39IGDPOkLK9ZHaYMX1I6QMFMXlPb8OgmYXHL02/6
FM5v3ZjuJO6i+zCuVz0+ucXixio47uiIMsUPdd46nTTiEJTx61Nboo7x/STVauLW
hNyv5K2YNxn7JCLhmkNXummJIVEEG5aGR7Rf+croNTCR2OflnVYTfmObxvxbS/ZZ
JzSOIOy3LbqApvGGzeIyW9PkMqID/rM7oTx/T7oOKy2EyIvJTB2H1xPc9WFxas7h
QR7HAwnZHzTzX8IfuGUgQmXR0Ml14ErNYpOD3aZgW8EFWn/HICxog5rLwt0jtGiz
2NukdinZZ6kiHW6xpOvnWF5rvFy8wwQZ0+jYQHk/lM/DiEmHycX0WN7CIfRQbH80
pyKJInreZnS3bGRk/q+A5ErEZYOx3vGtRcxU3d9g6r2yRGZNuYw7UxsiZ8EfuulT
sO/gzDHgK+eoeIqTzMfsWZY2jKtkCXp6WSgjmhb6N5qWTqSRG2dQn5figFb1aEET
ypUIEczIOf0CSs4CpLzuYytBhrxFcOxbfbFVReMSadeZuqOqNKrL0tPSSImb3orN
oNQUOTufdGLP3ER4WZ7OpHeeMPzKZ7NgkHnRQPffB7G9l/DAndHVMpI2iKu8lUcH
zRvcoOP5c5aV10xuqxm1YfdFBhW3NX2X9/yLlzbU6VtZkOinsj0zKSGXOPGUPOi8
WLDcOxZ3vjo5EPPADyjCwRL5z2CCxoXBSIn60KLJ6PVDCsef1TgSN1nYeEtysODl
1cWRNULk9avSf2B8bZoZTGqEb7CFQf8uUpCm4wG5W35wUqWbGg0vgqKlC7Y+jWty
1Kmu0pCwlzLI3XjJ1fBokyrMljNeMLMHLORRBW0qeMEC1IF/kI5t05rJZC9L017+
YjthSQ8AKfF41Ofv8ADkgQzqFFahuBF9l3OZfAkYdnyMkRuP8GMWk+majsj53AL7
eMbgBjJoP2W/x4lnZswm3nelPtbNqfpCEYPfYJyKi+ffQWJM1FtQ9dVYtR+7rT2p
/8GDiqoNn6qH7TFo2MAVL2zznCrXhvhV2SuKax4/hoPsCxA/+xnA/41fXOHDLSik
KEwoHcbNhrHk1muz/Njah4ZRgKcPz0G+nQ8BQ3I3nRZqoyJLtjCl+wUi6I/y5hF9
d+NzAVDiJPIzCzg3bod0ZV4bqOih6wYWmXY/tR1uIZoaXpr54u9uPZvdrxEKIh3D
OgIdlcAbB4a6eEmi1sG2qDYi/Esw1CtYLK5jE2XszEhZUWxwj2PI1HSU/zXfiNrK
Nc4+qpsoMUKQoCvjOKGBG27kx+EMUD3CUBYic3/r8Ccp4Oh2H+cMnqnaFJ4UrI2x
A5OWNcHnu0PtdA+G4BSsEdjYC2YM2J8ULZnqoAzU3p6/w6MskYiI1NRm7QF/qSQG
ePTdhC9Y5PcaHvZcOy4ZyvirCn6l1Ix0cr5smS1Y7jyntsj7IlbtYOV2NbhXITUD
5t1B9QHAKOQqgc0kyoT8WW4kyqXVGVzR86mb59eMwRy77t41u3betlO4Toe6e+qn
8uc2kulMEUuq0B6RSwmCZBsgsKGUI1ZVRNXabUN4uDEx9VFjm5IV2q5vkYU7kCk5
JxuLRcuGO0WLScXLJMUlPnRYlh/3UGUmHuKUp/WkJgH9gz0TuLYgNzpZPrbenBd7
Xy9lYQ1IhPu/2qPW0kDeD3YSglbNJlrZNujU5OIf42ABh/vlxVTzJ2TQst5ecEpX
yZ1QBcdJ/EAC9+VjtSd7QM3LPg/1qDond+cnRTJA62MH4pPP5x7qp8s79o6by/fv
c6SaqQDM6nfNE1Qt5kGXZ0apOUhdh6O+eVmTpj5eHpHDZg55X10M5hAfeGrQlkZT
S2LRIadozFmokzThFr5BajZw8Pw88VN1aguCxllxmzIc+snUFlpaoi1EMxXishIg
v0Dsc+9SxAYmASznPbj7Ls3GRqfe/fjTF/V7UWNZtMS0Rj+tK9b3Mv16kBiZGmvS
2bnhStfM66hOwF6UfZk+WjHn3rpInxdO2Btwwe5NUZsxvhknrOxc3OYCXhLiUBJe
sgjynjH3SzPJoUkQHdF2w+2GT6sGRGKGaJ2cfQQabipOelwNtK1lltWcZ3CDo8DG
4rZb4Jpk9qNvwQsKQW6EwzZ4dYlPN+U8ui0Bxv49bxBI/KQuwQjdxM6Xf+9Hdn+9
lPVN/e1MDtcD6lIOQZ4ELMzNCa+oBsFsOMBG8mAglkT8E5rRIcDW2A3w6EXwLjQy
XHHwqWJotZpHz90SHjqiqfVoAIJVMEL8FxMiiCJDVzXDK5rYr5M8x+fVrXkZJ4xX
BlFg1wy1c+ZTTG3aYDlK91WGOPKuwboOU1ylV6wqc2gnCr0PVgdEJBPP6fcdd3/d
XgZd4tnyqRjxaDS+xCMcGip8KkppYK+isQsSx4mK+B5CGQiFGbOxjcjMOLPCGhxW
Enjewh1DUGmsliIVueT42I0rZBvTyv0s7w9/0DexW0molKPdNYFZ1DKxDG1upqdd
QSojsrTkI9xjoWJJcszlSFendeMg0ERsDMYXRSVXEEPXyGTtKWR+pluq3wRW+KoL
SWeX2ZFa4YljLSe2/OcA9YqEn+zqXZaDgxzRCLcQknv2HYUuEGEvUIt+DGtuGf53
eaQli9sAaVgk9QmFB4FWNYPfsOqQ03lT/Drmh2yMFszb4CTYVQYq/Jk2BMyeM0bj
T4FAj6x6tqwQ0QWQ7ekmwIFbbf5dDGXtHz4jKfvl/YLncg2JCOc9WalMbOAPvecG
uJJ/nAI457BgNIFYfawoetoFopFb0GCbII2etVhRPGLutP82/Ltfgo8j4RBlDlaL
I9Agn8WiPARZtQ6kpkVKMXHoGz7pED/UiCtCL+eGYTiIlVxJVZXve3LpCv+MizBf
na1gBmLKDYaA/RCHVJLHWCL6L2uoc9/uF6+Y0MdfjzFmjsZ5F9UUHvOaMQ0wznAm
UTdIw5f7jJnuJMjILPTGupT4vVFOtQeEbeV+pwc8gYgAZNoBiqwewGlNIqzSeqcn
KNJ2m1TEqU6tTOr0FRa6Fc/dQbIDrgc0IaIugU7G/4PTN0KifbEwJTQ1V/o6feGF
mrJ3rO9e6i26zIL4y/6l3NFvhtuDijlYqe8zpgrcdQhFYWL2hnWdEmQtWpH32/hU
S/+59S3hyF7nzBMdwLugWMwgGlOyl6YXWSZIiG3PEwl5nr0nVTUyOibnShGHOaiJ
2vHVryiC43zS1nCRozkIvsWQFfdYIryx5VcTT5f3GnB7r/J38VhoNY+UVXIvDaYn
PG6FJX6SeCm7vsrFzo4BZZIRBcdXT4zHBwNlNQlDb5HtuKr4b8rVqFzR0Cr/i1aV
m4zbbRou8w5UmxZjRlb1Cp3cAlf5hyPCrzQ768Dywemt7c38VsIkSf3rpDRFEBeK
0OdSydBPKQhcWeQYKuhR2BaISxLzLqfVo3AtSi2G2wr9VmAaVLJhDP1BVbViIdWT
v7v9lVcrpp1aClzOXw58AWqmQpoN6hsp6lQgPZphA5XC9E2lZw1Tgsfn/2Uyt+2D
geheDiUsAKe4S7dm1wzFSbXXttwCa/CqiVJuY7TSKXJhSXS9OxeJE0Iu2CRhfoPT
tvD2abB1RJabSrotWMIbCX7wOA/7P8++i/cnXtFEIv6E2n8To010r+oeOKWQhVKi
vJgbwezAanUgwIoRkTjSQsdWKIoLzPAAN5gDE4HXIakgpJC1clk0ODAAeioVGzJM
rL3b56e/YhjIw90BIIy6/whnb3ddY/4M9eA2Sx5ACoWiUyTKGvYrdlDVrwoNs2FK
WBzXwr+gzn5BpUJT/sG+ks2HFbuAOS/fPYGJgoZjDQxEiiEk3fayIbafKBLkqczU
optgAB9yvFIFGbUqRF207hmaLnPP7k7/PwchXEWbcaLraieu1yL9YYWcEvqHiXBk
BP9Npsf8jnBkGk5TIojQcvabEG7aoHXCCV9zFRz91VrhEq9VOyrYUYBc+bQJACN5
Kq9iNRd90rSHMR0TfWDMVboj5DkqaQUVspUJfzTDq0RCto7F4fYsmz5wVyXcQcRX
uFK3lepEUvS8sAePMPtbKkzGvZD7lYwNAxFhWIorBCajjvvmHqhRmf7WwKUP5yPo
QEwvuUoE2AssOmqKyPtoZT6HWochvlH/rTvoRJfCAzDIYjxxKlBQShhiEF7TBd/r
xCvqyJNzm98BYx/cH45Vt5CE3cjtfC40B0TIAcyZeuwFAj8a9Igk8MC37OwWS2Wo
blsF4m+QyYMXHKWOX1wkGhxRfuDWf0vkTDwV0H5MroGacG0DDfWtgtDnpy8F5vV0
643Z7dWR6lqgbsPYXW0mlXfdXc5jOvBghNMUsQam8Fk/ylPq+8wYm+JRZYViVqjK
xBLqirVN7qTD7OJPiJxMVCcdtGCBYF0w4HeMUYGRzI+yc/yHoujJcz2Q/DSf5B+n
PV1in4spcEHKH4tKRXCev+G8UtazCLHMSPHux8yDEWyLVaRhJTE5hZwMV2Kzcdef
xaZaPisZy9uyezVFjtr+9AfoDPXhXnss3AuVuIoXKrDEE7sxvQtImmVGcVlI5szX
VfS8RzJQRnuJAebwXpltlToUiiixFPFiePz0b42dpRdgLZddJg7UcG/PImnPs6Um
xvLacEHgDhXN0aVrr+n7e/Z9bp0ev+n6RbmlWrAwenVjfMSR5RL1ZFWQA2ZAXnmJ
VxOktO+9dXEc+lbM+gJYL2BuxUlQaZV3rBxVsHHmcjc85rd7ccix37GafOt/vvRi
Bj15VwQix4UrrSnbUYPxOZwfSRrKTRhvwawAz4876P8e3Bt/znAQT+vGbJapDMHd
HIxSbmU2Y4HPuxzD78BdRIEA9YQfqnBsom1R6u1e1Prm1e0iDONfsPXqWbMXj4DF
RME8LgAT3S76Oe0i0nQk3/Xt8WH488F1XbxGMxIMj8g3Tl5eW6ioS2JOYQWgc6+R
TS+F+UZcolw2GqQ6aX1hyy7jjiL+DdTZgriqjP0qkUZDpw43HoRgwgYo6kj1A7VA
IcbfZnTc4qkZ32vEjU7Ba1lNw5bLSpvP+ysOdVhmsyGRoaoI2GHNaxbMv3yWmcdA
bw/jSKQo5Tvi7J3xfBue1u6RkVyQbnUn4YDCtuA/jQaL4QER4sRS46YRYwV2u5JZ
zsxedMOnE7xJvt3r4oYGEz0s/CDDu0aqT2pmnH6g4u4alAc+3lyUDCjik6MM9AJR
4OS5HCukGAhRiq97ElAj+aBqnBj8+Eojpn7v3mXFPJGyGYSHvuFmsoYWYEJjT9qN
tjnZA/Ci2Q5U8pBDI56VewR/9rw2/lCk5SsuCEd92Ym3KXrhNTC4STAiurtZ1xMJ
fB0EtelDaHsWNWxrfCST1XfXv9EtR4c7IAGyr1O3Y5O+9vlMpnHJLxSSmS5Ipvzu
0uJdb2JCGTbTGKgYrFtdjiCvmer9OOmBRI4rPszs1GBf2lyUKHNkmeiXCezVgiQm
iG2sYavOoA95b0HHI9iLqZ68++Xebo8NPH/QLPUH3e7VfdZB50fQo2ncC31+Ux8M
Pu03z0PEhho2BFgCYQB07YV9+O04fk2cFsdLYZDVwDfBT5bSzjGynvKbYlQKwVha
9D+QF2VOJma2DQq72a053SF0ycXHuhK6icKNUc/8sIAHGO7BGBA3L3Uz1HcZMHUx
elct2OVue93CGQ0mGlde/W9j6RUuiNmo7fKTVqWRkcCmMQNwQdKL9heYPwA5uI22
xobM2JHKWY5pS3TNXXz1GV6sHSRmLI3C2xKOzkbAjtQGHiM8l1HJaPzXCx1DQiGp
8uhdcR1qZxpFCR4G0s1TC48oR/uBjvSlFPrBk5ZzJlNkl4xvVtZTmjGcfkPCBPri
IR8FvCcW4SM8hJ2nDitkZcmqupSnN2H+FwqOxxBVjhYaCsQzXS5DGeGCrOCa1t8M
6s3CUsYe4POU4u3bGqtL56OTLHNGaNN1qxkZYe/e891GYzTjv+q6yHB0cc8f1/4y
yGnSNYgjBH8Z4o9Ai/nKRPNfhfaEeKtb2Ph70H+LzqGwq4XId2jhNOIK3V0+0WX4
XwF+Pcgth7c6JW2++98l18q0YVOjLGIHMS5oL9mB5/Br9WempUkEjE5zOh5aGVs9
wrm4UDw949r6iarMmPNuNP9wuHYGLI7pXCZv9a4MWTWiNttiKduVn5nE5+B1SKeQ
4Ai9Kjw6RgdE4aHu8Nh+inC5vVg6sqtyXAV8LG1aR5zhgazfpuaRiwVTkNTe4eYK
2smR8BkpRkMnGdINLAwjeWIy1Oj1E9bCPkyGlFybzsZAIxdX5ovFP/hddSMT5aeJ
`protect END_PROTECTED
