`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TwlQL4yweUIIBfcF0R313+URYLgL3rOZNKUiauqstVRq1LnDhbg5fPc+vLDugIju
LVsVcKIbK9nN6VPyIeq8xn5wK43yJzP7ruvglCBrx6jicKUoepZ7USwZDyRymc4H
RP4pP6W1NQLzt3RqZKxdONTR+lTrBJQcYltHaAkGURezarQAdoKEfdpD6BHQCYJL
EgX8fSRrM6Gdsa4nTKTTCgiC0V+2q9RI9NuV4G5uAMoaEIUvZ/yKVSbjbiE1F0a1
vHPQpQLEjuH5EYYZyDx/ir8AN0ZxVRiaSZ9QwY09oIkZgimULb8ueTUJQEsR+dfc
aznMOLWwJMb6PAX2lJUe03ljHqe/AJpvfBRrJNHv4MaWocwLHWOexnLjDDaaFVXn
YuqNVkQQt7pGZ8Yv5V0pPqRh/xsUxC6Rb6d4cSWky55tMuR/XKC7N4+fjHRm9dqg
S9fgKcD/HZl3g7KGxg+Lu/kf9QIbmlfxhm8PQNxxtKN2JLQuF48I7YYgdXIS1yIf
4xGb5cak2C/jQEkpuQiDVstvfjsa//Lb73iZCdH/V+VbOc1ocsCTtJI0Gjuh2lss
sufDRFZXv9Bp1lAv1ncvhp3rCG0G0f5IRbw4Cznbf9Q=
`protect END_PROTECTED
