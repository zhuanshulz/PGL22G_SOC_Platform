`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OVM+nFNygRX1KhB5PdU9+DepmOnLL90T+AWLYv6SwzR2ZO+LK9bOyIrmiuGN+fIM
H07D+ytZAcO5znwzEUC04ySAryAGwNDfY3rqgEjo8/dhWa08FRVB58nOX1uj1z/w
y7VhmWikdSwbm6gMHvX6t0c9gUqlVuRYiybL08Kt47hqQrt7/OVCHwZBlsbVIVmY
rM+coxvdR+6qwGrqF0D94RGHwb/OY/H4kiSJ3kue5BLP6xhMmU8JyPapblrZ/MiW
Ho4x5tenz3lO0KeblkcjVt/9vLF+jRXEfjVFhj5dMl/2PozLQGd6EqClKyh4E2Xs
B3YjhDgl2P8nt9UbOd6PPQ==
`protect END_PROTECTED
