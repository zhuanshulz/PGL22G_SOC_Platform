`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0n7Ut6kAquQY7qvBfWzx+qZ8WzVoa2+p/Q8CKZg3UgnJF5NwTypjP7HoNJMQsnbn
bX7f/ae6FDUayaTq0tmtc2R242LBfZ6mR3DJhns5i0DHqX8pQB0YbndOx+awfYO2
L/zKUgT4AXY7ILDvrypPktbIhGkuuetcQrkjsK4in9SxOrMxEPBJZcyt867qhwLZ
RIisGM2eNLeNtSm8MwcU23/5Wm/hOCfo1lE5Dj9FTrpSPZmCvGGvoR8dekBp/qD6
BKaXypHSdwd7B3kpF9zGKpxNEUrbX8RZOentVQMORsMGagBxdcIchJrvJSBILrhw
AT2tZ0pvio9N9pYsoS4tr3Y3OGbKESsWYZYy6kDzOKwankykgZ3TvnBAMwfei7I7
lbhDqaUoOWM/XgMl2qQc/RkTkUvuOXrEzvV+Lmuv8G1XGZ6/hRABmkqLhd/xAVW3
dt/P3OsIQiL3ikADddk/N4T9VeP8hWyXqJBLQlFF6iTrV3d/xXcK4SVcT6HzvU4s
48ky+LGcmF+yQ1amP38TkQoY4aN3ktW2GFT0mlSPnCU2uu/pSNA6ifIDvADHlink
dzkhVG1flPRSE4OccwsDvGN638cA1czgTZn1h88mEHDRUlJaEhxkVw6j0sA58aQ9
g4iI++Hr35FkSJOSU6vQy6fI6Dj6R86awjBTYaePvl3oAxfPWmy9kaMVWnOIm+jD
9sPfvRVK6dfpNyXiaqKfu4Lz/K9rr9i8yXBF9/1aVFaUn9RvybMIvImGYkpNMuhd
mUCk8C/TRsIsZEPRKHZSI2bw3wGC0CeDz+K8CbqcKn2sqn/hECFY0lFAkaHYywkG
hIrg7g9dby5RpcOkTfO4+6SbXkTN6s+hy8z3fymziFXXwTFB+Mzt7F1ZknxuglA2
ZFNAFrFTu0KGH/a9vOuam5UsHrheoCcC+h3Q+pm0fwY=
`protect END_PROTECTED
