`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AUBJn5x98cYD4vczWsngQzGhSooRsjIP2Y/JkdkCTA4gzuNJvm7Oj51m3TTJvRQ7
JZxeoxOt23ZLritIQ5rDmisiDxsxyCwXXPRVOWQfDl+kvPjmswFIc6CovtH3tL/1
ujlAjAXLbXLrmzJwLRGfWl+EgdDwlL0l9tRfxzKwmXxD4XVabgekMS6JdPCq42zI
ZQbzxAxYnf0f80Hl5jahpO77q6AsgRmZmGfkacDoYkQtRCbRuFyQb9U3si/YcdOz
sjrBSCuIdWNEJc1VkVLO5Rdjf62sfgdorbrHNFlshTBXw4ZohH6rGA5ZxYROumJG
vuhCtTx+qW3OlJKhTdByN81SdIUNukRoewUHJyU4fayfuAf6KJLJx+fUf5mn6J59
rBfhb1ISjDCa+egH8Yrc2g==
`protect END_PROTECTED
