`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZvu1KDCXd3LSd/xH8KFvM3sKDXzrWtBoP56wYB1KVC0vmLYTZfu4N2aGWJxeKt7
QEgkVr59Df/VL8wHlJHPLIBUIKWrmjW1h0MuuxLiW62ZcyR5qipMzJTC0vDfWpvz
dvpqzV4+HiohpRFtX7uuChAPENBPNgI9VcLg4WTyYRnqPEGcz02UJy7ojXK13KHv
DU7FF3WlpmBg+pQUEg/tWExMXupF/ofzT5wR5RLAQisIBqDyrED8QK6/l5bapGdr
71YIveHDQ4dy+xI0USZQYWotUnO+mCu43QejevbRnJ5NQLudmSNN0QQwdoGY4kXR
1Zp1cj8W63bFw8d+AKQcXAtj0XqcZq3z4xG2buDL9rllnH/KW/2R8VMTO60lVH5W
JQkYbOmKMopm5kEf2XDhSqR9l5hsW0O9tZeDYqVbp22juSEllu3ZNrNp60ZWGJZh
1ewPKkWHMSeBJCdPh6mnX0H6UH6g7fm98oJ1AbuJc2nbxW5+ucOeWvz4I02RZqkc
atKWG25Dq07ttk8y5FsjETq9ZEQzD9b0qn1Zm5OA9aMwIyd4CTRlVayNwaPw5bJN
UHXbA0vdt+9z4LUbfFmNMkSh8Sph7PvAxK280Wyx/DlQrHZuUkAyEJZ8yMdISzrl
R98gg0KOMHegKxzH/KYbx6t90JCphMOuytcc+OFOgEREbd8KhB1Ud/+SRKjNIwtI
ns8fPyfMv74XAeRa/JO4vEYK28F7o9IPwjqYBGnrmIlrbFz9jVCAiJKKep7ixQQv
WiozqawtuaFwP8QNXCkQ0LwwJ2ctEs0X4JpamfAxEXr/2ytUrcHwwlUeYzMrIh4/
tNnx8Oqq/RPNdNlfbTOpc9Asun+8JPtSVXR2+X/mUn71GOnW6CtGqGFPPHr4szBF
scNHWLWUNShnd+U2UU1DyHaXUAJSeAit904L5QF8UyqY2aSFqCoko7PSq+B9zusO
AkgmOjypOjm/QSGe3zJ9dCzfX5U78djS1aSL5zgo38Qqm77j4jpbO6SOTIKNTcoE
0ah0s/eSvTNlMLud6+snYuxbZRhjSsExdWJxtVD7OjEnhCiu1xfC7xhEcZ/1HE0W
USiTOIS9QFkRMajGFGS1n+54q8/+unf3pYz+qlrUmw3TTyzwJ4QLDg1MPtzRNuyX
Gg8vmI/gPthcPXEjyFYZXfxn2REMa0KsdmBAfi9+MvXhV6FGz5EuhIiTRCCELNaH
KEs06aFL6D4VP+SR8XfiSD6tv+pi1IKXAcgFnVXYLaM8K+m18Vof/mZn9MV+/yb4
caFrd/5Dzh35TSD9ByjKrwmFj4mJD8zEmXvCCw4QEVyfLvzRiAFW3X8A/vK3APsa
dYvZjsYSJfq4iokM3xaBta5l+J4uiftpkXQrM3LvOlQ7gdMWDiyYz+1CWIa5D05E
MT0OhWfzkb8J1QGGfIj0Bxz03dZnPnPLQH/IQD1VNLsgCuDjJleVMDsuQOp6uAVO
idRRfOwAMSEBz8Jbmf9pyqO8MhASlvXbGJYY45DMSPJeC9ouHMqiCifphtMLP5iM
sFIW8+18dCzjQ2pXxTToRC8O0YEv0Bpr+EWa84r9Q1EvhsR+uQnAsE/CIdZ+p7uM
dmEz3t3ZG4uUHoHyfrHRzmG0hqC6oMe2BvM0WXnkIQB5Hy/s/bmVy5SfPswPMdm/
sHgz4tKyOmAk94PuXzxCnLcYoJB+k9lTDcAdHKukQLtKVxSFv2QA8j7i3uZ4zbla
5+umX9v4HAS+6JK9n3xSx3LdNshel5vR72JyTRV2x6NbtZ9osjB63fZH/cfT4vUH
N7gexf9RDX47+/E4JRBx5xgLJxKSEmULchNE2Px1pVKq7xpoVqtX0Nn8oTIAqGHy
IHUBRRzoOVaI8uSiHn1PC+sSOwapG0VGxJbe5OgDFrWkc9fLTvKA/HJ3n8lhJgz7
wxelIS/mKzkAeX0ripr1TFXFN1NleBupEOG8JAgcWIQrpN5yZCbfELxnTx6wZPsN
n4VpaOwfBnyqcvtyiuZG4GWUvOp9mKNBNkCH4vKeRZk5UjRfNAuI00PES5c0XFwI
ojDKCXsxZm/C2rBsfKyRLyzbAK9VCV89+z+W6Z3HS3BVTlrPMrAWHTu3eFm3/NCj
qgOIKa/X6lY6ah1rjmQxaYXvoTkO8kclcJu6ZWbglYdKTuTny2IXM/W4RdkItAwi
i3/VF3UtvDYcixvBthf3WI5aJ1v1mvff0z12PWSmTciHHG4HmH9snQvJ4Y47Jaxc
svZ3Z8sX1jw8+a53Ea7YKF2XuGHGY3+323Saetq3PPu7RsZkyNyFzpOBOvsXgcsZ
r4D9hw+dYoK8Ym0v7jh4k12Ypft/Ghx9hAR/JcVJXf8v+7hX+pBcqgd7BVZV0PSL
SltgnodZvqeftPs7QHCYITgb76Cq1UmUYx+rzLuS0zHHPsMvH9MUhawFKTJLOTdF
qEvbRU1d1rhqoMe6CbHN+U/4HsKNmg4LhUXHgrO/eb7RgTf0f/yTzdzEcMIKJuqY
m7EjrQtMf/zSyyiSGhwNiihMKht25yyc3qSwsaZ7PF0rMM8K5vgDoSDLtCaGxdxN
dMjppVbRsuXNhOcbERcor2XkDBG/pEqgVn1mgNtBJaCuATXo/ObAXVmSL9l1yCG0
4FvgHtpTn2nULvMzczbhUYahZpsXeBZwMsNC3Ezq5rhb+7hPrnQPHsUyVL6dVhI1
dwddxhna0pr6aqS5Cdzly94GfTlRRUCwQ/5cMYB9hlp/4ZLuWk+F0YkwZFRiNV1B
zj+it1YMR7omXv5a1KH/6e69HdkiZ90yM0v9s7MfGu/l+gxixZ+YSNLvFNtrMQiW
hpxLAwiUOujRKQF1nmt67EvhGb421SgLPftxpdwrfU744x3tvWqWxHX6I4VeG4vw
GEXHoUL/BnF47RKHUuJ7DYK164BGP6eMxJTq39OKp3CkzpN0M3E/Qqos0siVmGjz
be/LFC4o2NDCEJW7ws6pv4dLd/m1iDHxiGOa1T5+eUJUR/PESOOpSqQEnNdvFCm2
byeB65oV7wzquscAIl4KEmcDxOTb6udTci0uYXqbE/mVW6tkj++8cN6QFy6eC10G
kY4UmBChSu177fx0LPGpT7fsv5FQ3kqDucu1Qm+Idx6vJHC73aPw3Bb4O7XZWO1t
HT0NKd3JxbR92mROqlqbzED9R4wP24r6MgoxwGBCJOvXlvU4bKmUqIEES+aPagZh
hn1Ky/IXSA1h34oz4oxO+PFklKhWKjxJpfEq0EIAS57pwq2X9DZ5owlxipoHVFLr
voLmyR7VXmbWxCvr9U6lx6h/4AXsPpmWa4PLyoyoXTuggoTAXSIUstDVYImo96LY
/nyDX0/8j7rTxWjz0SlOhpyvcPeEgnI9d2zc+ETl5hLTe4xNjRPk1Plkt7J0TWt2
PCRM1a9uYhOEUV9lWiYR2KRJv91SibdEN7463kg1zyKVxkABuRE6et+yMuEBBg+Q
rOVczaWPf3kVkSel/DGjm2OtfAtzD+Fnx392GdyK7CH0p9AmOPP+nhyCfcqMY52P
BTyBeWqc1m1iEYOlKbKoe9ljVAnyrEOVgQ5CrOUMtqk3A+5fK5oD7Q1GPT97yre0
YFwMV/VphPdSor4zHNdcRs/rag5438FnukfrroNRg+Sy2fRI9I+3TbaIyXjV4IUn
AHgtl82T7+LLkOxe/tlgrVzrX/DoOrn063aaptJ19djT9T7Tg6qexwYEW+RlPIvN
L1EMsvaUm6pp1mtZqxr41/m1fW+SVpVw9mM9Zpq9edAoFFV8IEZ4vcZEK8NbL/6U
gfSRXtFWc9u8jOTnmuRBt9iF2CtXf2Bvl4xTO8bFzYoXRTIj/OMsLOh36SR8P40L
IutoyMg7rEBnkTHkbLdo6UUYLl3ZtNOt4Ehkh8+L+v43x+uwHjp/521YxBdnYZ1/
JwR0YooXOxRPUGZiNWcmI/A6TiWaKQVid6Dt9LI7zC5LnYjF9wSzt9VSm78XSnwN
UlStmVEmsTIDNb1QoiKt29bsoSBamB4Yewb9KFTDieiJ10c0t0LOO6e1bPVCxlYV
A4UZElA2SOHGNwtz9erhgnkNzfzr3W7Tkq26UASCl6f7tYdWbnliaTtpptXdx/yt
613MrXikI4VoT7KmjOcyhajx40bhjqVsHfUC82SHJ8EhIVrLtNa8s5f8zVF0xc/8
b8jjAvxUbxZG2liHLRkGRh6M4IaISKsHA5oTsF3EWjHB+wWVjcX01SzJ1S+6EytM
BYiBO3Gw/9A1zKHVyr6c6YpfDrw2S9vqwdoZF4i1nA+Bq2bznu0dyDAYJHyE+0J6
7eGyufsKtlO25RCuPPCt16QNB6R9VEBA+XCO8xVmae63Y7ujoYK4w7K+BaZzQ4dI
3NksW8/VNZz2iDSELKjDi5j9TVH5HdKk1SAGM+dyOgkysOQk7TucILlgDIalJN/w
whRLr6qW6kIxTvf4/Le+TGyTSP4SYb3GYokhTqBD5kiTxZ3CJQal89p3bEh2zNe/
UAzy1aYqPOMSoEmA4WdOgEdVgYo/lbC6iuTMgp4cV84odNI2mHjG6ahbQBeWeJ4q
oXPYukXkzGcABRimMbpj+JneeO1KAlc2J7R9BS1HxzJ9zyjC2jiCB6CKB9fF1qbY
hp+g5WPmTfH8PRE0C3/a6aCujYNfhnqakGQ7rlWikn9XnH6KK3npyXdDq6dePTfi
MA5TMvBi9eXuDhKWGgr26FJdYkMbMTPkiXfYlVhh2pOJM5ali4hJSlGPc/N0X4xt
kYhtDB3+mk/QOUf2XE0+4N/Z9DlNomVVnMGqCHtQs4RZwAgZApiITqD+gQSlo3Vh
np4LcLF/VgU0ArTktpEi8RdnS1nTQ1vmqog5Qs0z0sTPzUJNqMNK5TinRfU6rBvI
hjn0/iqHczKEh4flxUrpTJBD/smDMW+c767TSChQSzh34tzMEcR2TZgJqkuIbTat
tVXmWYiuq5TsRmWyxhb0K6bx2GqHTx1ZoiRyMgyrH+CofyQ+fCnYMUYNN2OzCdEl
W7cT1RqMs1bliJ2rhSM2AMd40eICjJT8jwE6InEOPf04MFHgvZYSBPk3L22npf9e
czNuk/JlbRKKrK5NqEJUpfLGvjeCQi4ZSLc18ZgvmYOtax1uQ8jbiY3K7H/MBUgP
2baDUSOw09qDDnhtz+qk/MqTwyMHY88AUqnM5EBwxXrrYr+x6uQBEjRPjUemhsHY
fawXTo7Loo31TojLI78QWgQgJnL+TSIe/kmYb3R5+rpeulGZWE5hCV6vkaPSd150
gdwmRGE3tIp+7/92b2WLEVwKA+eZy7Zqeo9g5s7RMaqoiQ8EtmRuBZukK8bZAqPK
XjCdZlCWYPB3PtAwSVVw65OlycxqpilIB0WSykC1nD+xwitqbeHNSUmNq97o29Om
oQPmui0fJQGNNHsjpeEHwr+TzthmoNkQBqWj/GnxO2SOSPoNYuLZuBFdfYR61QeP
ud70ZNOc6rpdZYZRV7Z266oQ8aNywVsi3NwnLsZew2WwiQfy/TYqz3d8F6TW5hi5
YgNIxlvE5nS+SEOkuFZStR8+JwiWN/PArLr0s0tdQYw41PExutOXQMq82wkdWzoq
rsBQzlg76xkJhmDaN6N45LB4ra1JQGBlOCAQtLzzcBzaoLsYr0rRwnm/+EN6U5V6
qX4312/rMHIxEd07YUwLOsxdLmCi7ij4/iuviQovoQIaGdfc2fZly1Gdapy+7qfe
BNC2MdbVZ7Cph7oFo2RESBL4UaZr8xOmmSHUlL/U/16tenXiUyHTgX6KJV4WvNzH
lI34McoI+BLFjdOvFc3f9Fm5Ukg6Y3Wksbn+gDaQupbeXzI+pJG3qlSwv1RTV4tB
12Pk6ysxQGPGH4IWm2gW1sgFhOzeeqeTzdr76AUCWNQo6YS3bppkqkE6fh64quy7
TxM5TqV7JXoqRzByRuYoeLraEKi96eeGl/bT9nr/jBf5Fwe1AocZXlrr55zi/SKL
t5gwITC14DawBS9hlQqertPRijJ+DkKyw9Bs/Rrm9DmJy1rTH9xWAHpEUNtOglRl
rDzphg/KPbhuxVs3qTXxF5knfQXDFIew9mbxIske9DQjjygxxcviiWnWK0CDu8JR
EwslKS0+xC6F/BdxPb6O92AswC/PhKF8a89s/9hOCsXzwbWTDtKspvUEZRn9cwR2
NpRbzaOCSlPqh+Fq3Cq9knMaKdXxQgNoHQtea4akPNSQ2e6metDtuCJEnX8/fT6i
CtVloR1FjfgE+amCczs2FlR5NQlf83vnyLblriAnUHuMvHrWzo4sVYr5WQ/vR5kD
VudZRQhXcTXIkJFXb300NKvCGfWe4WNtzeW49e3+T8f46g9DB6zb/tUY1WnTT4vN
Pd3227WagFKARYscvchkJZiIuRV1kx9D9kjrAjDgDLzazTcWTddRaZRyE8AehE41
Z4NHjPIFB1sxZzNtlcsO9+hBHiOH4Ce4ijidk4XB9bx0VCSdu7WVmCnUHoU0Oo7Z
AxoM50QaQ1S+wBdv03A85hb5pBKMbFXockOCdQzhkfQIKJHKeNMOCzugjvJKL2J6
ZkE4204Ruf4PjZBYUaP5H7NhQR317n9YMBFpLWtw3avrYswaakM+UQBR5P2JGJp5
rq3lJ1lQIKHM4lxJQ7ObvHnLvIVkJVoZS6jsIPKrA5w+FHPNJBPXoiTr2B6AfEd5
XzxThc2xYCXRlTzJTBoblymguS0ccwW+mcfQ2BF9y+VObHWc03mDhz5S2gh5aloR
1+AteIxZQvYXjIGEx/BRrw==
`protect END_PROTECTED
