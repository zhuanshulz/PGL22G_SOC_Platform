`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qwQ8k7trUiScI2KTuIik+gowqZHgzf6mKwAsvJ6sdSoUXWlR6n4g7Ic76x1CWpV
uPWJC5dOrAJHV0+ZQjAhPB+VEhL6pwHzQ4Dyu0qGMgO0QdR/OwR4dVL+XtKV+YDy
yhfo0dehl88mA3ZmW7A7FZhz5tqcfCiJnAf/zM62emOB1IYNzVuy/8FvjQG80NUt
/d2u7KLAabURANzbqvmq/Gh3YcOvGl9HqRKmxSIfBHKCDKzpMgAa5uH7tY1wNDzu
w3y7gaOm6/8NbL0Ohv9wG52dz5gKoLXPrjTU4jRg6q9E8cSPlh8MiyUMXJmM5/VY
hWHmI8+v8y/RZ0Q7Q7TbTT6Jao+JiRAuZkRmXmz9t/Sx8rnb60xIStJu9At1d5ow
dRZoWrtGgqZ8NUY3tQQddFFdZ29DNrUSqR/O3GH89ZKxah4nqZvr0mkrIwAHt2C6
W6Dt44z3RWxb/tK8IW3lQVaJIloejspNAyoUdQ96Bvu7owPlLSCd1eDQZCncA8YN
wy83LbQ5BiEMSf4dS+MzbphJqFgvLuXWNptFgqWPSCFjmyJ7QUsFX8XYZ0Ics7dO
wFOMGY7tyzCTS+eua6l6svnm27tVX7de/UpUpd+d98F7rU+jFxNPWSCKALftUa1L
oGAFAstlTLMan6roTVldtjaJPbXop+Sl4rPI3DdAc09NyeDlgP5oXu1CZDeIGKAt
sW6UF3z2WjzelEaLQQ2sA69aFu6ay4jhdCx7jobxhdR7hTKgAuG/WA2E73wS2t8p
68k4iBdEIaoAsfJwckeDtjBXXrKlmkWAUW3xxb/L6gBYeCZzgSxFmtdCSx9BB1k+
PwrAdQsi7GN6ZbwxJqiJ84BbvjZAtd1mXlDzgrDTB/eJyI550ekR+9HDkpP4MeJY
R2Xam6RmB2RQFQDnid1kgcqV/K4SRjoY//AkLO++rsC9eoUQXRCCx3BYOuXcjtrS
U3HD3/ZuFOZa7q6w/2IgEA==
`protect END_PROTECTED
