`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6dn1Qy4fANvmAU5UwYL19ZQasjlXtCgwpHAptZ/bNUnUC+0/N0qulsPwAK6Yc5I
H/3Mw+PcujAIwHNCxrEHYIPpVDX6qbo+NkSuqiZeptH6pcraXJHRkdCMSOFAF1RK
s2drWRglx7cPKh4HBKxePU0Igv2dN+ZoZIsvdoinh65DMMw+29Vx45XdpySC4fcO
+e8q57Av3xPoBzC+kvDDVtfggajyk6y8E3QnTQhxjgZYsN4gdQmeGVGye1cc6VuZ
BOezoOErWYaYiPPs4rmQN913YVs6ga53hM0gF7xZi3rhrtLL3fVS07vznqWpk8fH
kdCkpHYwjDFMUa2/N0AJRFDWM6ZPllJdP0zJMb69FBQWeYjCIyxAwraI8+KF9c8C
u4I4tLnoBySdkdgIaNvb6A==
`protect END_PROTECTED
