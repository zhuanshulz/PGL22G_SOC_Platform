`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cNxSb1DalaR3gpGrfIckQ5bbjMe0TcoucI0VSwAL5ET74LNz8O5z2mdJgPp/m1ny
QbG35sf+GvwXi4dhocVNathqjamhwX5ptQz9znGwvf51bPO9zVHLR+qTA+UZiZ61
KktZbziCn+jD2awzvNQKal9tDEp+KR4J6WUT3Kj9xb8Hd1B8aYnM9mc5hGY8Z4bI
P/Mo0FxI8ljLi5z4m8s7Jh+hqZNYyMjVxZEMllJtDpmhzUb5nv3N8ttfdinHXIIy
9GeUH6xXjs029WIYP9Ns/oTDx66ed4A5wFiP2TG+RwEUwc0Vf/dtQMqiXjKj7Mbf
2Fkrr1QPzdVXtjO7JIHNgYDMU9XncXFchEM//xE4WhYw96oyhsu9oqYyrPfBNShQ
dg98WBWY74/ukR8R2fPZPZiaUEct+gYjMRELUuxIfEDYPXalzkhE053ezuawJ2nd
or655PNXyZ8EuDLFTV6ghGliexNWUTQMszo1+f2QuF70EDhuSnPHDkI/Fz0s5D2H
OfqODSzPkILu+Fg2F2R9IZ2Lb/651AFtm/UW+REm5ekLUHJaACcbu7rQvKU3WO6G
zvPtfZ/c84lF+tgpYLEIdj/Mq44W04/F6Xu4X6LvWQl5XYF4mdXhV9kISb3/Hunx
cJ/w7tuPqWzZrhDiETHq+khqOTCaH0+LnoSkCSy1uNqOmJapckJOKJg+dj12FM1m
ww+TgGcu9Mx05oimJhEnsoQlWO4j4os9euVw5rtSrGqzTcvuWHf0xK2IRxjgieHw
tf5kGAMF/EPFqEp/gdeOc8O9LkbxZn5G7nslHTra/yw6g7jAdMHV5/5/OVsxf/g1
7JNVFQP5o7qguaXkLvmDKS3Qob6S+S5AHLcoPPG9b6iy2DoQOustBlwGyfU9QGOh
uzpAiS31v7HmXnLumMXqHGfADepZKGE5HsKpf7g818FRi0j2f4XZgbBPZ4F8UUiN
jBL27xGz3QTrZ7k57wV5qZelFCr36mZ3rLQdC71mmhrV9MeFvXfRd1ftUH6Inp8w
UOrOoXFfOOr3Jdcy+IMSoP65cDD5S5lPRdtgS/usUC0kXlUMKuLVBOiVamBvVNrZ
Xq/A+Y9IK/uSbDf+hOaQYGW59GZUibzPI0fuCbRhwEKtJcNgRq3Lo9oszB2iaR7p
Dekh/z6IwobIa5NtiWCRIxMJcIOqoGVYUFSwhRjeJjFUIxPaftzGpPFK9hz/qQpZ
EjeE8SiRDtFrKtQvhP4DGFL87PAWmwwjO4sNJKO6TGF9QgYJoVQ/mjzLx8QLKHbJ
sUu1HspEpHY7O8c8DTVNBz4Inls2HTbwL0TnDfmlRdwBrF5hPygGUDt3TuvT8Xul
OkpteClDFKtDnO4pPc+0VqjLWhZ00zVs34gwNgxFhiaeOxScUuNOyA/wsoDaXfy7
FOeNW7T0Ydt5hUrDyDHadhMKDm8B5d8MesKOlnxmp5wuDW3tnnuhtPCZ6wfo5sH3
rzeFCO0cl7PjXxrtkHVg5u5UY16tnI9OYa1AI6kMAbC1wCNaCboMcobFASrQvLKq
pcWtQow5tQl9v7uiGGDbWOzw0OT/FfrJLuxcrNlEyk8rNNILtOJixjZ9PeU2Tp9t
uUQhDIm+ernT3hlmXtdAXkfHzt0y9l8DBA3Lcenr/onSjiKyI1VIfHcXkq/+nbMQ
`protect END_PROTECTED
