`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F96PmkCrIZG3bXilVRswc60VBFdwTWPr3cZuNvlT0LyNalwuMbdm809c4kMN7tok
1Srzr986PdF7aFcHbOWwf3Rbr+bVxzG5jF0PLFGgROyffxQeVumho312+E/4y0VT
4PNilf4SH8Gyj6El9eNwfMoMnLN1tJh2f+ZRZ2mek8o1O+WFL5bERchC3IEJPFyV
VWVP7fsXfcfr2eFuCu2Q4Ddhcyx4Xym4c77t1Nlr4YDBsXUGwKatjxWSy/OHIAzj
+dwedY8KoLZxv4nf6eGv6X9LrGgrZpOiBwoA2lpaFmAGbOJUKC2mMLVKJlU3oypd
NrIR+cBmlfwaljIc06QDH6exkiwnFOjRTZoOpfrbKE+1RTGlicQBYteaUvRqieXP
7tfIglqwW4qeKyNjXQN2VUzt5L79BONJA5vqSnLcvNo29freppYFC7H3Ged3eHco
v37keerjJKs9nzfJYyoMCWFJ/ToGGUpHNmrfpUjXCCNoO5kcpQc1zsLUZbTcxAbe
AlEhUduvPQZ1poNc2kXV2jGWtoyNiYYBPzGfU+RLJ9mpEBTEH/hYeDEcOn7aYWsl
/5c2OckAHhQOWPmrp7x/WcOt0E+v2Jn8W/aSvt7RZKduGJCfpREr0FmepBddBVdH
90HyrcnMHDa1dnlWdHCjXwFIwnkKr3V8TFmr9Odnkq0aJz2Zhg4+t0IRdwrKlJeE
7bmERJRJcqtb8ryLpk/C5mhKEeGt/e4pCf8ZuRtZfe4sKT6kXUB47QcvjNO8Usol
NchvnUH+9A4qaLeptUdYowtRyTRHLN74MuhEmGhzEwtqpG+WN1KDQVKeA4h/n/Zl
5nOC7VVxRsWm4S6W3ldgegpJawispTfeKGk6hJtslLqV3IQ19Wc0bWmkn7pPjerl
KTxOBMq5G4+0P7Gs8VjbWTBt+1VorlkrP68m/dj2H+p4XuueVb3dWJaX1d+HP9DI
PvzdqdeM+eqeKP3JU69QxIoWMv/xbSjbOxXSbbQrQKTO1uPd3l4J5+leWfGq5PAZ
tnKF/4zlzxbm/Rv5MHCilzOfSlQPb6pq/hm/GDsugiquuoL9z12SvJSBk+fZgaN0
x033IIUb+H9eCanTUSR6XKvrvCAsfU+sqfO+7ZupnsAtSqpHGBy0MWD93AQqwHcu
vzCHwoVcVFM9KL0Ew3CglzjlPqvz8H1axSIxBbJY+5n3Ocn0r1s+KlQDYWn375Jv
/oUBGSbMknxr8/Ikxbr9tlf5OFcqOUzZ79u3n1bZI/JoKgeJJhrTVEL5+uXaeUO5
K3ZNhXRgxhOB6tEXskACEzTlKDEDP4ReeSG22HgnygPnpjGNYGp7beQkaSVhyz4v
1MGeVLWYKFUIC68RhZ3PlGdBHrkfjmRhUQ+B5/8RpmQku7kLZtVCtPLTmN3luFSQ
E9O7rh4gksXl8VxAaa2xCZ2QKBAA3gNz4apgaNa1tQLLuTJNXqgHADSVySW8LxAM
GI3tg5+a2lnsr+dRdRaiGjQyGjeI2OJkSBq97PCMH91YzSbdW1JBF/GsRvwfAk9x
fNaMxf7TrRRhn2++ly8whVH/928ij8JgmgQfbJ7FUxd+qSYUfIPp06Z1cmAWRLG8
FUidV1SVsiQ76iliFyJjfFsIKe9EKqCxOYQSXdymXtdt2Xvy5MqOJz5Wd08HPUb7
BUC3RjKpiycen+uBpy/Bn6CqT5MRQtyiK0eYKuNXfom8B79apUas7Ku0mwSOGqTX
QeejXJ5pwnSX4UpPQZqLIw7R6v9dVq0uBnBOH5rjKhxlSpOvEu9Q9YDxDxe11hYa
ZAQ1ATm+uVApO9alGBmfvMXHTgZmgR24SmbPXDHG/7bG1U+lXirTIvsCYz1+rDpp
cDGtW4S4ZLOIQ/RAvF9EqZ9Qz9e02liE5gyKrrdu10/nWKIrqZelxaE7JivUS7H9
K0wRYitfAbcc7V4jibqdjGZcE5fmmMwQP1ztKgxcdDRZlAhPnO250Izp6BTr5BkB
SfF6l7WQRYhOG+DSPryc2KBdFFPwyipiPcufWCc2kg4+C3PFiUZzEbupfvAGwyNd
Ehit0yOgA4lj+TbPISNZNjZ2DgqPS0IsmPGYJ2+e/3AFQIPWgsH0udlsAu2Ptp31
zDnI7pc0xVoooARhwVzvjH6K0HzkWO6oWm34ZFp4G5PXYt1ktF0+wTk1xMxmNduD
YucvH5NDNlHjzbl3InlqHx6e7sT2Dy/BLT5t+DMmPL4ASWrHAMQGfJoSzscOCVB/
PHjJjsUHmDqPffncyD/+Ih1dkH2pJXZ3OyN7+M4YHBvy8tD+wZa/U2HWkbbn4jP2
Gk2OImT3qISTOQWBAsGUagINWFwLyPI2N8EmPkiajhmBzu3KF2Y7hQqxFlDSnQRk
905sW6nDdAmiV2gDRi/Sx8br3qbTPFSt5zqVlpJT29IGLWWDIaX++fzAcsdlDyJ5
O/avPcc6d6XRAGa/Q6xQdnqungOy96cdfi92APHrYg3wk+P88WNDE9rt+mn4Clsl
xsfK1zlUdOe7uUwFjji+nIRd48pYXMH/3X7eFNRpq61H6nOyMu621DrsOH8vb+qT
97yKcKtBat5hXAk0UXz5gnlzidvOE282AwKIBXX7DZYKgo3VWNF+M68AfBJ9BRzi
msTZMeIK+TsSYY6rMwFnPDYRgDImEarS0wU0gK5IsF4QjKSyFhSE6YQ+znNdmVq1
H2Swovl9Xgh0+9ULpd3MafpSGLBnWZnDtbOW+aJn8TA2Ed9JrTuDHpueQeFOYEo0
gsvlEyy8E5xXffXXEKfJvGHsWk2L/w/pzybsCje2Nlcb4V0SAcw5cO6sT+n8Tp8L
XVDsEliW1tLgMpYrkqhUlZTuj6xPpiRNhTvix7jRVMQJbIzQxnJGAdn4Z2GwVKr1
Ga5b6HW9tVIjtmg0VRJyhWLPgecQz+8K/7E0p4xjexWNLp6gKDVV0HKSx3tquu/o
AS5fgO0evvoNrnqH6Q5CXa3UFMe8OVtxdTEFec2/OKYLcaX2rnWA/0HvtTYbntV/
qQ7SoL/hSonEkKPUvpFHQ4Uk5i8+8B5w9FjSTGFYJtQhe2jCB/4Uyd7eRAB2YJRN
Nao+ZS9pEr9rR13Dq8Z7mIdhl1ZRpDkQBGu3JTxVzPSMBLuJ1WQvg7S3HTz2TK6j
vfBdyxOYTtwovslN3VgAEvJFg4W8dgZoZGXKv9Z+mDC2b8g3c68KXN+RnSg+ZiGX
uVgfR5ft7UmmHmaST+OqQiPPEyTPVHg0R+MA2Vy9QQ6ruOTA1vlIJN8vS58IEoEm
+q+opnQG5GEpIrfLZp7MirmKvf0SOY4o/u2DruAnqwuX4vLjFWfvwEhHtdHecGrw
QMj7s0xDyBJY6XZU4AWTXQXNgYj+qiuJB/1IhbaGskhgPcp+irEs4ZSYaonK/7zv
krtHOKriu8PV3HS2OETxjA0QZTTFC6lmIgAL5gZeSBZy/FeSeUSzyO1zx7pLSwzY
Im6nseoVvvyTW4/ISCrTF9FmMQMVjalmdaucA278nzdAs4APQfZhH9rgnJfOpKe+
kbFrdpJA+FKSjAaHfxI94pLpO6YCb3pT2imIG/iIe/YZmXxMR9VMCJet3RINnyQV
JPQhFpiNqScJUxHev1UdIjOBUEqg6h3zFbJeNzmYQ+BUJcolAFHi6dB1J6ozrfs1
DZOWh8ajuqTOZRP/jLOMOQ==
`protect END_PROTECTED
