`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJ/new5O2k9jnwSijQdkHoTCQb1SfhKiGc1cSzFoERVxuDSiW1rTti68dSkoilr/
erJnrWLE+hfCe5/GVrAGWhs8sv4qqok4hPpKtjYioK0paev3Pn6qluTW88b8mlaP
yf4S+clQmK4rlUnTsgHmqcIZ03i5wMbArnybDFpm6ip9jfQv5YO0Q1wJVNLU4Irf
AuC2XosWfw8gK12NNN7KxNTmy3VMB/NqbODh0w+XeC+qtOZOzIJZEzy3JLUj2ax4
m3vmf4QyYWHM1oy9ClEUrRWPOX+2UD/iG347Mp1Wrbh5jIgi9JxI9a55Ni36ykgF
/kVw0KsExnKqPHcippsUbRxeEsLOljJTFVtgKH5ff5ToTWtiKoTp2Ky/kYB5F3eb
06oKUUNLhKmUq4qXkG7ROrq1Wj0q0rgBgr7iD8Y2AD4DxJDlzdvuI9qLP05ORg2z
aX7cS5DRbtRw/h5ynU1GvNOFcxvm6AWGPygenOOBWLKjrtii2tRKZBq5PEN4b1tW
QwPqQ4YwdQ4pk/j2pxtmvvZhiVUGddAYDWiKUnCJm+aYRZMc7V0J6e9Q/OkZtWAj
QSRzdaKZNCryTY9A/BWkxzZ92bRDOZoVYdLUaV+L+KWVu+WqE1SZr55zXat1nCr1
7w6HS3axGEnBJ3dWhrOXPsD45FxMOH1/s0lyGZHwjGfSL44q9dRksL5CsH9Z3cOG
OvsdPAuGuF9KEXUmWaIZcueCnU8GOpgNV53p5SYRNFWthPa6pY3a9muZVlpsYlJK
O90kdDklnNrTCBjT33Mr8St6yPuqmfieztfipW3hDLqR6/vDm9KcDyfhAjkhSW8Z
b8+OyipkHKD9Tk5OXhdgMvA+ZkHtzPyXFCBP7YZaFx7LiGzIAQ16Ffd4YC3gLYAK
PIU1ZPCC6V79+BO1eOfdM5EZNoYqZo1xFQzXRjIcFH3kLlgQAptJowna4m/Xw5Dv
SxBHNAbEbfe/rFFA6pIhs19CJUzDVyXGL/QHf9VbZ03SqtafCGVvXxGGZX7+9hay
9Q5+xZhiqvTUifaQxp6jDKqf1DgtBWZbF3x8v0j/b50hJc9+LzbulnEG4IIxFJ4I
flXqSAT/EktsIonY997+mfXylaM/O8LI/sITWf4VSsZnmjQi46PLGj0Ypp0h6EyK
Eo1fKhl2xQd89QVR3+wLicfxT8z/GTZuj3w0o1n+sbDgZvcLxb/Gfn5Wggr0NSn5
yo4yO05LZXCt1Iep2vx7BnVYzK8hv+3tGYYn7cwm2ECKXmcrEh1POmp0M4DuMdHG
12jFct5lhrhL+jfhjSNZ+MPr7rlQiPVtcZ4oDt75tVdOMrUReInMcXQjIVJiF7QI
/Wvq8w7jk/3HnJtS7OswCtHDlcjUub8hrpi3Jtcgkj5RPQeWOJlqtdbU1dy9AeJf
1mfRTjIrEJ+d61LZRLg6J6xh+dcvjDrzyxMi+ujMZMzc09jCRYtMix/fMcypkS4W
SgZgQNLG+cctt/Lny+MWPkRi7acXECE8Nnc48s+F/fGeCj4ks8P2tNYd+2ZNl/oF
NdLFOSIegEeGldL9oddHF39cSFNIV2HCqpLfgcl2gNHbpSdsk/ghOG5Yt3p42Q5V
Qa3OKKGES669RWY+jyXT8/kYK7kzezy1FO/ACEEGGNCZj+WajD5J1Q/VepzntlCK
CvY5bLX7DM4nFANio0CF7ZR72zQGGcqlGQ4sRpIfEygh1WUcbX+i3wzPKIhPAblx
PFmeJQ+a4V1mXVzmY+FCLocNaKVB1iDF/gSP42hG/n4gf0+5BjVgksU3NE0srYAI
rTS4T17L1T6v+AhYtCWPJiUR64igjabD+DffriGNGxm05QgUK0Z3lOMQe2G6J/uo
IAj6oiA7kdWfDCAavbfgxm9gji9D8WgdM/HH0zxy3jcaWKFgQcJFWxKS+fX+iFI/
9NybP7iabdsiLY/m8w0ytMM0CzKZ+y5q/+OwgB+yjgI7Z82rsjKuDYNyWnFH3hSc
GOlC5aQs68VKtERLY8LCMo6b+zsAEeH/5dNShGm8aYeeHhcSPxhv0EBNb2FeMWz1
rlyJEezdOSBVDCSMcAIiIgB7gsok8ksNm7IAGcSUAREMEMBF1Xr7iDmvWxzkn8Bv
45I13YzE5PGUo6HscLcmiLNUZeq5cYscY8RfxaOZSiKrHpCm61PqSEg9B87X4Nip
92UGVvn6upWtdggggMf8Ng2EY9shHELK32O9l8wPnHBSTFW9+l6yY/rRqFqcwhC0
5Q4aC+Ix1rCIexMZl9MlQaM/CK2U1xmf+QfGYKOgbgLZh54QDbXWb7yA5f63SS5b
uda1zIvycfpesQEM+4IiYupWpGyALfcRyKEbgmVdgpGJQwoPWoxvUVhtOQPJs86n
TOUpTYd12lMNFOdZHEkUg+yifUcGEi8awTOepN1MzDLfXobiv6crx22tVGhmPciY
oDxnZlHlfN72IZ6hvp7JpcQABhW+kD+6FaxUw7HGK+yfd1sJZsviCVje7g9fBaNc
/MOCSdkG/JlffnK4jNiRZovdC3VtEhtWm0YTlWcgxgauumJ2eZ78R5j3m00OB9x0
46cSjLAWYQM+g7GKYkeUni+KBzWPd0X23uB5zuHCJDRlG2v1Q7tsDoXVnn2rF9pL
g2Huh+PByUUSJY1OZK1WnK/o7aYQkcI1Ac021B7nXSA=
`protect END_PROTECTED
