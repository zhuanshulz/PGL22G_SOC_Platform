`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
poy6cdT7ryGFncH2VJCvUAFPuUXRua6I/IpZfFzmSNDOKFJ7vWSI356YgijTNduw
89BtptZTck/Jj1XLkEO8CM/haeydcsAxVBKjcNrObxUxFACN8wbIRUvEOYe9k01n
pb7tVTeJNzbnQPDXDXfpFH2NF+NC3G1BoNjygrUhKCXuJJ9G+X6AZcR+vcz9BL9i
+/au5sJD5d7vwDydEZ0Q/eo5bqZmgavy9rhr0wlRfrc/GBhhoHEDKV6RhFCpsRc7
zU0ePJZgMeljQ+zGxHl2MnO/vSEJoerCNjNZ+uovIqmtIuknmtHM61dhrIDNyRbp
KOrsJckcs2L4bRLT35Gpj+Elf8dE6CGh2E5XEzFUP6wT6TLPXBsPTMwj2oXJsCW3
0XyO5w/8m2en8W3t0aKxp4rMV807CFNDwuAf2DKna3T0em0ZylxniBaBODwhvxI5
m5cuXbdOBKtk/VJlQS1pkUutKIJmoU81uAeMZrT9OLVjTAxRajUgTfTzpAT89CxU
ry/YxKyGdzXo9pGI2TZiD2VW4zNT4TriDPBhWGn4xq0Kx9GsnJDil+KB2SRlG2NY
ZuQTPjRfSDo4/89JqDCRRbAQH05IHHkGx/Rn3Upq74StJPxn2Wet5c5HuvqOYCLi
XCIHVCMoO/TYb6fZQxcHvbK7ra+68t5OXGC3Ag5eKKImpD0JGkvF0+vVM9Hhbpy7
hEVGm0sHw1+z2qxtqfbBBp4wvcUs0SVYtdogqVxIugJRn3zEL033DlXCU9TFfV96
vVcpX5j/dJ8z1xOD6U5/2eX8Vlkp/zh7sMxnFK+Szt/oJXSQuMSC1mo++kQIhIe/
M6vpteFYJh1q3aOdPP0WZSmZ91LCDiDEz+B1Omnv8rAIzendw/Ho6pd7HR+2kX8W
6zPzv6ITrQJXLfZmtP3+tJlLievX7o+uryoEUZFyW8NbQZ7fTwKPRBa/T5WCpnzQ
BR15zpF++g7VqZKvCnEiLFeivz/SVfhGkk9Ky2IXLMtda8pfaZJe8YQPzZLSuGq1
dPFbTVbLQ2YHQAB8mMkstJfBiSnQhSkRiNp744ATokVbfwKCcvTsya94eCZUIXER
JykJnWHtbiNpMDsxoZtU3QqXECGRsNkbdNbNWxnxHIcFZq/UdRNnXi7qDaOaokcO
VfOVeVmS0RtdkBLPFA0lopTYg2da4iI/dkQsfWQu95M2cNcF4wVfse+iOiDhFB8l
K4uqL66OWH/mDTe8kKUObKrsbtxtkQWdYERWLxo5mWmeWb1v9BDgsFqiz3Ix7LhM
N+8mLMThJlpfjK/7+DiUkB1++6jhhLR+Ys4yrh6bEMFWA9kwVwJgbf29ATkkD3/O
WXrZ41CREN2R4SiH/JZyPhFt8TKJz5Ezl08PXnFvLOlXz9+1fyxx+IgJfYcOlIY0
5pFWtlDkNOLHfZqgnm9qQB6hNz9KtDS+MzanPAucrjQjSo/yWAEoOO3lLHQo76SM
+lMprlCaA8+eFPX25FJczK+wFDWmXppg8hf6FCxHFxKQ/KLLk+7PsFgz9KFBMhnG
90iyYvILLen/SgXHKHHLW1DHI3UxGCPNFdNoufJJIzf8ZlDo/nxWgnnypeyuk2ba
7K88cBEP7sMNs7CRbUE1U9jp+f5XiiwFLBm7ISqXslQ76Ovq+agRQU6pabf2wTMq
Ypqd4rQ83TJrip2gK8iFhaeo9gXwF1NYDgA8GRmDZ7uCEDOJaUnGujYPvYhgxfIF
pao1oFA13hxHRE1NblXJAPaAAoyzuVrofkrlTRdCjRqmD6cywtjXp1MeGQLGRtZk
HgrcUBwkP1OYQD09eeMIb/GKcQjtkLmTppxKBwHcJIPX5SRl9LApbRTU6LBRvqxH
f3i1pKIRBDTnNmaoV68wFxqrwe0ZUkMw+9EZv0/7hWAl/mk8wKgDEYPpsXSueins
OqntZiaKbQuUBxwsZDsJgQam6z0pCqRhJuES+HIdHW6xdwgu0nlRu2EhlwtTqzqI
Dn+wVkusxXgT3N0maZIfvkwpO2w9nx2t60EGNMkkXFyCyeppYHfO1Bq8NxzmUC17
WOfL2g6n7bKzqPSNQ5qRfkvC8Q8MR3fAcdhqQhgk6YPEiWxWKxGr+SP0V+zbT7Nk
qBZZ7b+dWuPryu0yLIGQa3JbTRcA/KA0IJFj1IQi7KP63XtLH9/Dp1TOSYZGyBXy
1iv4SgxrT4lFqzRPhqgU4mOqWn0wK4s/TMBbuoDgC6IM8+HTTnfUVOsUUitEKVtl
PeBzKKkfZQh3oIkJTyuV4/NuafYJRg/SX02Q/J+dJXTE6lsXGFf9jbI4+98n4ne1
ltZyblVOMKNB/lefJkugb/G4JiQZvSeheP7xhDtcSU5Fl0OiSpXiKg5qoRyrtFH1
N/xZTtK5YSkUg3gNUS+AlVDEKR4A1Eo//cNCUnIJOextkRnBPRgBS5N5SzrMdOX/
IVR8Y2LIF/8fETr/Tp3xpiQ6os/TBeJX4486Ew3h4wAdpiAAfOjOyAx26FaP5lp/
q7M35g2eJD0ZzMOF+xVe1PhisXp1v2hu9ryn6Daol8P5mZGYEU2jMugvpU/dxamE
/S/UyPX4cGJRpuwYcxMO+7FNGqIXq6FBPMsXrAKOfoOb7LCF8bIArqTH/t8L6ZAB
RkgtUBHg9VqmiRUascZ/bkxkEHGfSfUPfFSdXE0sa00FyyE/D6MNvGwva+1tt6HL
HsfTqCfgcGT/t5kTdU5o7NO2R6BuxPkhKdipc4zHDHKsNZ9eoXg7LAmZXRuauFyM
B0OgscPnLqf5emGfb/ncyFu77cAnKROenuW4uWZ/mj1Xwox+YGif5Qrv+hG7gQxC
7EkQQhvniRM09yN1OrJxXpB/jfxr9fcvOnjifsLORhiUQQIi67eILKpnZveXAxtl
WhsCQnxnBMJURWCeRCr0KwlUlAsc9/rCMPJWxui7RtdExf6gaOL+U1sul7gHK5rl
zDJUHoD2JzPLOi2iqZ8NU2ePe94b7//Dlsg4bE1Ubq/t3jsCYdJuWZRUM5I+koQu
4cTXoAfP1K+zWEsCoXBZ/HhOmaOcHld/4HZkJvXrb3MB5FO+24/iUDDsWfANji2B
w9NIOGu6crK4piQPNMsIboahG1dHsFx7D07MDaDjovKkXBNb9D8nz/hgIWXuAUjz
wcZOyAKPWPodGSI/8hFnbHXWdtFQZf6KBsjTFebMpFTZsooHImMNCRejYPJWtldV
qKw+KF2Rs9BqCgW9DwLAgtCyDbERGnlRpmnvSh0hbKKNy68iIFmZygsN/xt77mxY
d4ZlnbF3TTeJCmJ1gp/IK4QrR1NPWevCraMH1T7lMapOnJzbY9bxC73C6p4tF6HM
EfnFXGOz8cnDFmpyDLTKcFAqM883NLffOBOGSFapAOe92UMmRBVceZwghMVdwj5a
aIB45KiwQ7HkTz3HNvasbXgsY8ijmiYANi0EoGhE4uRpvzXaY3x0yyotjDpnMZkZ
r/Ve91RmvwAwgCYzuLvd9f+3/zrL4AhCiJE59ZuhJq7sXGPopfkprz02gSgEpZK6
g1/Bu9A/Ayw/O0UUJoDfUffF2YKedxJ+WCiAtKZAjbp4xi7tUrbJCTKOY/GYNsyC
FLOsp4WDpOrfrNbjti8aJcLhFTK8jZrmqDdXV+6KUHhXi7obWXOySH8M6HnoAR7K
s+V9Vl0y+ILCgiP0NhYlGWuA5o093R4j3bWU7aZ/nnHxOOeNGjN4xYLS4VrMJGCR
5X8yGTGHwTto7b77Boh8enBOQjzR4KXn50TC75mi+AI7mOJ+scXaMwcBTrS4QmYk
Tr3nvSxJdgREI9oVzhzCmj77haVyPHh5BDahGVNshCP8qmYKF03W4VYSqtPSlJhQ
ksgXyAxhgoSAtaxetcftDuMoK8owjfnojGOgnm75AuQ22Dd7exqB+JsPJQoOGrth
kZ6Z4c3owWdWSpjRPyqLZU2fJFPqLC3cGlS5XT4NP5vXlYcBFmx9XkuIyddDLkQo
qAIHncx7fyHBcFEQqRcCWfA7K3gZXoWLgXzsfC39LZhivaOd32i4NJjFfoRvKVsQ
w8gw/xmHjN+7UFM1BiYbub45BwJng389a4UdmZRD62UehSZN9DXIIn7mtc7LvSrX
6AchI+cb2XJco6M0LvcSh0WB1eHldvyU60CfqEeX7wOQOiOFw99v0+Y7Ky8twvH/
YNRk8khIgqC1rnlWH/plDIW8Qdi+jcN/PBWEMYNrZNndzczNoLB7ttikHvQXM0Is
l7t9/6TkxCV4fIy/m8XYaSOU1e2sP0027iglJQ1sSWDEu7oZcokP3F61dlMFfXG9
ozYqriWN73xZyG9OL9AotgoF6JRKgGhNyfl2vl4f3hG3b010mh/xICmirX1vMwYS
jTBc+rl8Jzlqg4eP3Y2oipthvUaAEJjK0OhprW1VW3Qgak85Cz2lqqasmt6DwV6S
HWK3hkLdrAatBqJpg2eO7AupxHRr+9w88jBvxhVU6dyv6q0HIBKJ4DzAhNrIErIS
OUVboLY3pXA8T2V/CPVLD96/Q0NuggaP5pjYJ/vM2v98c8EWU+HAP5/ewzyWB5jW
rDmyWwNWWn0wPaddWdcnep4mymGzPCdax+F2vWemx8MBpRM2/Ehqj+H75D88vMA0
h5u/I2N2Bl3caBCUA/vh3zso57UwlR35B8R/wSYOWwVrQaYEeWj7ieYnI1jBJ+u1
q57KoBNtb026zycaFpWsMFzwJTelQcjMv0sS9FXw344/gHUNNk+STcHh3zUvEhhU
CqEDTRLmLQySwbRjW2U0v+B0bqKtLQOTMfrWMJE9TE0SRrWSBgI/qxu4fWFAU3fg
lEnc0maGw5JjZJSQhMm97a8RBM+Qc7I0tYxDxn3eH1ybRHbKa41ITq1oNpQFAUMw
c7JGyAxT2xJOY0RkjNhqEL4zSsD2ejQNEy5lhlU2bGGQyPnR/W26ADnKEMrYMZ5g
SPXmSa+KQ+cyEf1B5Z0lYL2K79rBDrKDyYKBR5Sm/ldv18GIGHKZswbsXmtjunJ+
nkit7LKnn9vgHS/X3QczMXyyM8dffqO1PKJNKohxygO1yBRA/nAxYoGwxmF4ZI48
L0gqfrh+PS1QSNVXejkTjMAt/vM99Gx4ZsEZt8tA7ZSQ1m6AS2clQ/reQRBloRpn
2ga0UfveV7N7xifi3QyjuXwDtnZNBriMxdFU3XwdoZAX1o8LfL/Dcb2P3XBrHbah
Cf6dgV/bduhAqEBCHOcdU/05n/D/nI3gQWZnuQsvCmwOAa4OTfLn8OqNK8WdAOY7
04YHd+DKt38sT39LdDEArc79iul9Zk5QinYLDSSvYvuxoBBOEvi8BDFqan+7oh3Y
128XWbn1NsMqbHRN2GQyXZvKlppNXmjsIHewiWbhsLA9QYO/yh4pS/Hn1SvA5Yif
q6MwjK5rMqhSgSBFKb3oCTzbMqmjp0V+ioiqcwBbYw4jte+xrLSMPPXDpm/mCDyY
o441nl7LY+48+MZBOhoEJIe99hXgO8xVHt0Lqv6ie1ACfO/erOq8Azd2xncos5ks
OLGDRpU+zarvcqE/JsoE25RG2/duHy8oyqr21JPQ0WKGcyVz63vsn4T1pnPHFw7+
IezDOJiAQHmEmMte5VgQWYnCUcmHtT59/y446QHTKzC9ClQBo4PNvREwkUxnEfdz
VYDKpY4Um89f61eOziGudnPVUfskaLU9KDUjs9IB9T6pjUBTJxS0PpRLBSTUQHyF
9oxJoPSQHTEVM++45DJr9uUGLhpzkwSPFfUVd0vvc+Gz3JIk1OdOXNdKqk2+eiAf
YHHQaM9D7DeqA8YcMNxhJ+fe/T2DpsD15HtFPbYl6x2mN8pnCS8CKOFaxUgB/80y
dYeRyeDKxxTGTt5jji/8y15/QYL3ktn8PzVmdjkh5Kssw37Euwdy9ZxKdUStxAbE
KnlMAPROThB0d0+SzEq5p9k+74UCch4fFIP1oqOPbclckOPO/xXNYxnAUbn0An9U
alJc8vwIVf/CKpCnGH6TkmHyH1qofQf7SAanfMgfrhVOJKFUeWi7gI+3cyfjSkgL
utHPaY6oY0HyUPv0xj8tS8vHsZ5hGtavvSqeCtnSFGJ2QCADSw+wayloXyO0QjN/
FoBQMKpag/5LcnFNGUCFY5IeabXxYNeqJf90irAnCKbeADFIpuwPEdi/9R+mtkkY
egyyvgzGUBVJJvLP8LqJw7WF+CW3kpXzogZsqfeqPDHvEleP6WB+SXVZYC6nqtEd
OpwCLaSoZi2zJmDUj/w1zGU/vu5+hdeUXuAxcAAnYxTJGespKnurXI++ZRGdOidJ
b+M55Ph99seeJdmxEjwbps+qnQ3Qri6HuJY1NTdAWHZ54h6MPy/rB/g/90bHOhYT
p9BkIW4mHkhkMQP6ncq2buma99fraIzMwe/eg833BixKdv+ovmTVdOQiMZy+Wxfx
dvzrQWuiiqUuw0XOwyctRTueLyZNIyZKHDPrCvm3iBaVS5OotJao93NSgcfmqJjj
6p5RygboIGS/tqXwItac6RI5m+ZtksICeQxKeUacRPZGApFzzLkcnPiaPKnHKgRl
j7wUKMvdtpwrJig54vnjy92hB+kqVTorCESleFw5/P1j7FiRN9GNj+ik7rxIJVzE
Tpej/z4yKUcnQe3v2fJA4jUs81rNyF7QfGtXLJmC4Ul54U7tD8ApZzOoK+dDrxNs
DNxnHPhQEqgtpMlZ2Vi6+sHoUzLislFsyrb0JvGUOsYW7OHXY/gHJSkqo1w4ea5U
8Gn3wY1P6tZdg7y8ganvZck6oBoNWc3OP/3QMRPOcQv0l1oux0sIoSSpOx9+HX1d
DNmmMG/5RDLPampWb1VoLP8Bgeiyx2whNGxjIz5o8mIyCMo9GzhSyzIHbWwjQM51
EcRz1NVaUamLcQ78xRL4wUXqY4HG3qnC6PqUgUcNQ1SLTDQZ/ofzwFHyCZskefme
J62fJ6YrgNHHjlJKFS3fDTfbSawLqfIS+JDjs4EkBTqf6T91ptMafKshoPjp/gJl
zHvp1UpustU0a/8UobYzA1s0c8OlpEiYxSCCpApGC0rzTcOQqBdxYjrGJUAzFZjn
C8ASLmxpvwDPNENsuEyMJq5EJv8n0nFn8/F1XEN52CYdcIwalq72qGQCB7BfLk/a
ltvWJP1DrS0ZmUIg0ULnEn+z6CK8G4uZTBitOhxq2G8sMDTVqbQMBvAMcLlORNLP
zN0r9s2wzSMbipiUSIX6J+pjjbS6P7tQOsO6WtBKIamIwv3MXls8s1/c9eIH03pt
vJjFX0AXcgFWqaL09WdcNIze6v4vUkY1iRgDSNuMSGEnmJo+fzkDFe25vtVnZIFs
lcnR8B/BkIfP3jmRPvDKdrmighel4VWbNI4gb4BqiDIZMW02H/6LnCZxkOK3TPAZ
JAIRY8tB5ng9MWmLK3gy6EIDxVxHjzod3L+sGKs6cNByn2X7/Z0IvVZnnG+nGE7x
tIkKGdVFyJNZP0Zj3y3lfAwsmI5Qhgul6sO0MMoZaskuc2PUslUYE5TAOZyqxt+0
lc/AldsyWlCp0IhHEQY3Y1w/gegFVgV73hBTog5/uNnio5RgSXgxVd5IdOOVgz2s
lE03c3FdAnKM2YNgsz3KnNU8N9eVGrDu+k7zEfV7vucKTgDfua2Gu7DrKFsP3c+I
lYZzdNHXqGynU2JnjCrMeGZPMNqEQki6WOtoviEyBhNgGetPuj/ZuQWRrbj9xtTy
THNVnrYBuDLJ/GcQAMMZo40jIpy7riEBxdHQrulGjmVbBCdi++9ycE7ghEmiXbEv
3kkcZ00j4FXNUe+nUlSsn49WMGcolWwoyELdaMU7RHd5HhvRR+EaH1wT43xjS2nA
zT8ZfVl4g8rCM6sHj/v44ZkGeLaPUV/0mJXhtIj0l8Mc74sk7qcTcGqvjoR4g92V
ZCC2UoQCWTzQmPotLymybBqQJ7JDLIFfclWW7z+5mBEC00gAAK7RoayQOkrssMJC
EWE2jFPorWLY7jL46h2sJaDtOs6qSIeteriUaJhc7eVr2fipAWAzR2gJB2d3T2V1
G7gMuZO2l4lTtzP3qrIOM6SZrzHUSHhlnD0UoBvtggxBCU6i+mbuQhWFh6Bv8Anr
1QaFiVvVluayOnDDy+dcfTaCCXMfGlZib89n6fnzsolGvt2QngNYaJsK1c0dMovf
+wqWvzHdWZhy0rNgok14dlt7AD5kAxVLKrdxPuH418x1rXZmwvLQ0iDND5Hqp4SP
PJj6iiWVziYerm10CHLaWW2/qbj6PG+UHlrdkFkQEvfOE4CHP+Y5w1hRMO1YGYz+
R2chuTzlR5ypLjYt4Ydf/jlIq3eWYdfILeaZfKmhIx7qDRsdazX7Xv3wBtbiTlhO
Tl27sXpPCNrwrqyiB89quloG/Uj1HoEzF9ma1/k4n29JMbO7xxjIEgiJrx9MVkbI
H88QnxDNY4K8+/caJnaNQPbLeFGtGVtAvo+/+nLGcQh8P2ets6oX7YTohAmyAfKy
dALaHg4CuHNfImbd4H8f7KaGyP5rMqOhWA7S2XmbFawqemJN6sO+jz885NWCvIbh
cJVWpz2xTog+S8P2huZK7XiS7e/iJM1QmQ8m3SZ4Jc5GS/2NDo3x0a73aj2wpp/W
4NZPcJhJNo/jBELePh9okcEwGvZVw6T+mm+zyevt0tflxj5mTCjcFcxOVmakrpoq
h9GO/9Do7Wb7D8AR3YzLnBAiB/56MFSS6KefnKacFfw45lFrYWRbWcCnpuARtxND
aKe4l95OSQT1arWJn+gLoLOiyV1OWJwGZ8Y/JCJlvPoZ0dkL7CcD5uX2aLD5bgh3
DRNzE6DE45MQk7vmUsDEPj3iXmvsBEOT5MMJsrA1huCUxw3RfPOy/uRHSXvv6yFH
snNGhAPjcF+A+JIZbGUH+Syv8FXGG58CkUpABQewI4e9hMxgB8wpud1/JXQqMjYg
3ZlOB02AuphXL1aCmjaexhkAjomRf/ef3/WNpa5UfbaItGwhV/umR1Rnx/whKqZO
Ie7XarwL5tw7XEAjq8sMiQeVR3sYm1d5Y00wJBydAPZ5/KVT6maZjz3Yn0rbFoc6
qxgN4fWjp1h8mNaBaYtQJUmf1OmzLAd3s0ROCoPtuXSNQ2b5UN7+J5IauoxhFY4x
PmfVsAlz+lyyUPEm5b0zE9Xi4EJ65w3jCZf69LuMLSHRGFdp77a4Sr2/BnZpMILk
iP2JeyNg62QkOD98mUGTHvJ39IivAp4YDtfPtqTPO5NheKri5Vafz9sf3CHWZlzz
LBJ7de2eO6B2ZxsBoFholak1xfUuDekOqz0M5rFW782xjElTEGS1ad9Fas8vp5Fg
rHGoAM8AXBt36QVu33umaBUXRuD2MYryAqhbSUuVGRpk754Nqb3HA9vV/ld4n2iU
wRrCR+8lyg3ndacOO/brs6Aw8YVMo6j8C4UDx4wap8LnrfzJ7QHsVQBw2NGW/ryq
uJDV6asZSAgg6f4ScYZkHbMaTR00S3qpYxhLynz1AiJjyll+AdNqrSSmMNp0Yysp
X41K+71VCJYAAs/j3PVd7GG6MpcLfkG09MMjwXPfhN0gsnFYIEJqPxLF16VE1QPn
8bjvLs9Ulyt6a2mKW0EnLKP5vjrTrSdO+4ckXCKtJnHcL5FqtG7c29rx3yN0FKRd
j8WCuYHpXH+uLOfheCYXgFXvh22tcKHUaoyU2fbi5+HR1EazTE4v1hGcgvs1Lrul
+P46PItPC5GymJODYLX+V1bag+qHjKe9AiyM4NPQeDIiGbgIzrc4olMLNHXPRMpc
+H/45OJSVAMQJwEPKpmK/GB7ibr6jTV0Q0kuJbYhY0GRBYiuImTZ71DQOvEW6ytf
q9d0S7/l0kDC3zMI7L/o2MJEfE7F0ShSXZai7sa2qC5UUwoP6ta89fd/3u16jPie
3mnU+P/3uMoBnLGKLF36L3ksEqkZLMNwFZ5Oqi60u8JrBnQheeSu4vtXaqaeNR0+
lQRol2+K5iv4eqlcootP2clnPHR+I9MbgzlqOIsTmBnwBC1ljJeLYKpMhSfzH8jW
46nh2nVesRN4MGOIxquVl5rKfj2cc0MjhWFZe7wSLEwlzsSs6dOfntihtBt4eqhL
tOeMRQWURW6nkizThJfJKYhCNluWfe4FDklTpnjkb3NzIhc6p6FaOU0vnsAs5qNy
Grp92Aymwss2L0YvW2bd5W/mqZiIQLwJ4X7pnxyTXrKAZ99c7h8U1GJmPApytuT9
iP/Sua8y50KnXl1Dd8PfUvKRh5Z+zACxvOgsmJV/M+Th3wwAdD1TdOTsGnmFT5PX
CNsFTXM0lQGe0zAobUen0jrCNfsF9Uq7/yH/vckQP7CNAp+GT4BkJ5LHP+16N8wt
RdAo5+2Mg2B+9qICZcxhUC69evi0+SOMsbISD8ScX4DHG57XxM4xjDEFjXIshJtj
nJwg77NZTS+9FQFV4NkHxE2cl2ksMpONAFoZ5la3If0jaWg7iGePuugknXIN678a
M/8/zvTTx0dHgqpTpZzvfl14gDbvo4BnJBbZZzcP1CFi6N2otDdkfu/90BLO7UzT
7ktjtyKqotix9nGOCVXYO8UhDrQvtftNOcJuv0am4vxP2qH7WOWf5QYrc/igfmb9
YUf6/5R9/PI+rXRJCapW2AwVCiaRsPbSkFlAYrmfxHLYipvhIcCz4vXVx6jWuwQQ
7Bcdr74haasGpDoeO68fDoM5NUo/aajgpjFwo6GCb2aY6LqC8YV6a3xTcXYTY8V+
KlnaeHjpalMHMgt6qzS3EZUcEkbKxV02jozQP0ONx/w5ZN7wLAHEXPW8Y9qZoVAD
oh/FO+ZkZZDMIeSbPI12CRfRFezhMBKWfO6Q7/GA+nNth/QQ1HB+l/LQynG8F5CN
kLFL3s+iN2NYKy5z14d0sycfNt7YJk6fjdnHcdxUoXkgZodoXqgtO8IJnWyE+uOz
EOWGdy5k8KGrLnv5NlZO20ohtk7Nj5iqc6UNzyN9AZQQUjMyB7QoZs6JiLnYQyBv
DQWqx0Rb1SnB8ax94sHy+vjBTEW46QsPDxiUD5FQh55SWrNtpmDuyYTbGcm8I8zU
m1WziUXY0B5/8Ny7Yl+jyT8rXcSApaVlsJAp9LXJ5/8aS7a6ZnteZZV63p1y6aHg
SUEXl+Dvew89attwnswSiV9Nr5M3K/USHxw9XRj2mq1KrAZCYjDGT2xMsAbd8vBY
FFi/r7GQ7ARVGbRycmNeTJxTIJn50gg38XEaE1cnPa48EwhCaijZ+HIu1SP+i9zf
11LkoBoWqhvriAoEn9IBAYJTkRVe/4l8253b3Pam/uzwGM5mRMEwKvtczj1cgTK7
DFrUqNwTZxo+whaRczSO3xrATzdledf2j7tURMo0tCRLg1qh2ENhRZ1KOmh+nc7i
wCWhrR3L+ywSnUXGlx4f7TrBMwvaGxKTLsycsQWKIby6kzJD3pdEZ0LX9iw03+08
YJvZE9rNfe1Ztr/w+sHWrWFkzophXh9g0IHhZD1Ue74O36XOW/zeReeuC4YK1Ku2
wK2q8wvUjF3K6/7S1tUX+3Mzb9Axkv6Molo/qiCnt2AFUeItqIyTXCieiV45t2cB
Gx4bBNwWtK+eaD3u5LBhjctKevkzw0Xy36wV5EHgIPIyrdPD8HCuToZlmRaFAHYw
/Hx+rwlKD/gndo3X7qP7jxcVnPs2tGqbAsWMLk8dhFNvPJV8KJGyCWqT0wMX+XP+
dbcd9aHQmBCRHHKUPgTjr3CtJl34MgBm8cXD/EYfQ5P43m8PBWW2JcPxm4mfffen
DvmTX552sQPK8rGqFocfSeU2Vryfe6z9i+LpEAMojYUe9bK3oD8P7uLoct+n3dQH
CnFXlcEOyU3o5TECnI+ZgyRLPL6BbAO43lPxkst/Ka/GhvKgXRr6GUR81GU6Bj69
jtsK8sE30estbVsCxeq1FgGTDKrL7DVPZ0fNf5OJIANa3/U3xW+A8avvwmlW+Hni
7WCkhojwHXXGYn169sDkbogUkoMzP9pDa+QdOo4/TiEmqIypKKc7Dwe6VRWcCY5O
Zf2Kn5zSj1sp0ySCwgVJ6w3Xzq9CcFQXfozmY6ApamZVbeTwBPAsvJfKXx+JHHdm
dABPB1h+xo8k0znjgw4kHv87iHqmmP6laKKD/cAbZ3BQ/j3jyo8xhZ/+Ld6jnG1/
1ipz+8edXyVFFU/76+mRPWWQh1eWNUiAw9i+OUNBIE7let3yFdWNkqv9v3rxyoBk
qEWInqi2aDsn0ZGOOH3oMeLaGckRLYLjA4HDv2UzR+FbVwuF78KxADKTHTw/NiEW
Y69e+dqXeYbkow4S8QRTDfOvy/N69LEFnS5D9Y+kAZkc6GA7VqXI20felQnuFmmW
q55xAuIw7csmnIIzYNyt5W9PjmK9+K164KVNIW72Tf9wEXN8vcp4yVFU7mLT7e/H
MW78TSm1cl19hwdSgFIUfMk5afL48agfypNNyQmUNUjftyUrvdvu34RQjNQKab0X
WRk7TaKY4F3N3/7lndLC+Wv6GYnw9e099GYUaLHrUWcue44y7pn8zmlVZIeRFDg0
X2sa9VxcBqklNxbREc3C+W95zetQOQ2DPBra7ZrO2PNLw0rP+Mo6i/mBQTnRdsOg
/dXvgRk8JdDHLePo8RtDt9r6fSSg6ytPScdjv+LVY8nZHieBTFSMgAmF2L3MOfk0
kDLnGAefkpZLSkX+vz7uSD5YRBpBHXLpgq8vs9w+NJ9Bi0DANJlunoYqMpkPSZzf
Vqe0clvVMnCPXbD2AaLj651t5tOlG6Bm7OBi+yCf7T1/4OVAxwzKq6rRYb4qi6rH
mPSBYkhapwhZcBvbM8hzIKDVPf8l25R/XmSWMUWKMWqZ2+O+7gm50qr1vGn7pPWo
OJVpAhXLCeA32ekXDsOnc6R1Mip2ZKJTwJ5xFZqUrQOTqNR45mXycH0JfdzLg7eN
9Fo8MINttl84GXbBJMuHMIrDJMTJ5pRktIRGDjwOp/66jD0OmuMihdz7skuoi3WM
w2TMiFV3G3ED46R4WSLC6b+Bb2Ui0cXKLv91LzdxDK3GjT8TyGXlRzARK4Zhwm5o
M/4F8QdzQo3MvSpWge4oG7/8CZr3qpGRnw7NN54+iCjPgbc8NkwDPsCjqCTCprFb
hoQMKnXoH1PkeT/k1Js7LOzLaNcF9KDrsasrHWb7YROXt4U2tuh/EMjT8dolzirO
O2rtmOc8p/NaDVQmACRWT18N9zqk5LAtQthZbuq6xF0qVio8VaNKfU4m1fiF6vvS
eU3bysIs11VGsV+2K+WB9SR2ukxYSE3j4FsC8mJJEdMKp260P1f/hLmR6Pk4/cmX
JDQ6PpEZpRvBih+tIak8a+Y52Q+hc4MRzZFYx4C80F70nMXHT2X8jlpMg5J79N/a
IQRsXe4Zta8bnWaiweULKe4c2aB7V8l3vKKCbnOiSooCR1NSG7adV+IlwzX+kB9G
pNlrqi0bVHGSXF0k26IrciFpiw2Mr0mydruZdZGJoue1q5rBWOIIDsJRiFvIj1OJ
zlZTRmLpveBSz1vDxTud34/qK3WOTuIkw1vH6+8gwGQMJGtI5HCt0SldqWaZoV0B
wgcAeg4FL/KBi53+9toywKxuhUbjzU/kTS5YbexxjiskSHKnP9eJ+lwVbau+x2t1
if4PZQVhlhiy0v+23UpH8poCn6PoJDGfUnpfO2Mw6TpSwzNCZYFgwohbMvo+SQT2
BsAuPAMkmnJekxMpRk8+36x99Y1yMvULAKRkVNwxoJD5FDivy3/Z0R4USDa1z0un
b6l/FDzOeZ7dYrZHZF2XGOUVYmaRfN3bViMSWW0pAnSZ0Se3O6rH1YPsgA3dYysq
vHhq8+Vz7AxAZOh3gsTfNYeMXxmxcwwDfArhjK4bG8ygcKGXWAH/8kueFF/yCmfu
k44TDPN0yv9fhqRcd3KEBP+JgpjZ21347dVdbiA8BiRF1tLohHYkZ8P12M89kVVR
OYovqV39o36yZW/OU8QFrEKK+yks88JL97v/LwwnZCvR7Gd1ct0aA49biC8lkmHW
p0h6m7fbovc/igKVY/O9bcaEI26qg+zY47/Tpnhfr9qfF76ZQ87o5ThjH3/0EQ6p
utCynejWCMqDhrepmgtU17fkpYM41KfAZqtIVnnt3P6vXbX2wrEKachuo9qPAAYo
1BQMNVr9ICs1OQJEa8IKb7r8cPMeuRF6Xxjk4soH5l2V+yd1e/vQOXmEo5OD5eat
hF74Kn5Ps1g21VxWcHmLxdZoQHLYogUQmo015HmIHPD/bFifWD5261UkvcxsEyNB
fDfIOCFwomp7psERoBORfUG+KStKqvVNeS28lnrE0A0cmhf7IzsfvIs/cxCaEZw0
trmW2rWdAG9L5i/kUsPX4GKnNZNlPDywHRoQeH+1KqPwnQeLCav+2begv59QMKTo
3mrKq9tn2U3YmO45CH6Rn3J3fHXr+QTdLbwYqU5XpJuvj2f8EZEsGARM4ABiyZzp
cwWMAz9hQaBG5VDyX9Wncks/9ZD1OyfMaYbk8LkNDFpvXrqCEEr4e9b4mbRiyK1l
XJgRJ7tG7ubI8nDtAnPNkRFLCCKAWzXpeqQvNgT3Zn68h7Vp8R4hG1rBVR6UiGiS
kKnx7iig4renTSFEb3Vf67Wurb1Z4ld33GIX9vzr4Y2+RUxdiKlNDm44fark2XN+
nTc+tOvZki/pvLxFmfJr5/V+WtKl9ePIeArIUZOfv8LSMQ9xkAahSFuioNGcGWEY
8sBwcGgLdd839f0mKJpRQpOJm+sohq2li3TxAEm9Cs/rLl+nCAa+I9loGSpr2fIx
+6EfLEiivLvYNt+e9bxQqTHsT9uznbfxGGzeT3zX4QBYEPm946M1wa8vxIABTJmQ
36wk1+bINYqdKI8gkJ/j3a8P+rnpQRKCq5a3LcXU/WCqPfKxvoljOse5GO+SDTWm
cbbK845Jp2M86IL4Yj0NMKlhJq7vUP9Lk/Z7Z1ighlu8M9faygVbQE/NWivmnBkZ
0QNeNEIcR1UW12o8HfC1iujE9PsFw4XlbdfUSAlKjWWhNMprgfEh0F9NbcOoAdA4
1FTs5b7efXk1iN/I3wMlNnvd5EyyOrTmj+FMs7BOpWsr752ZR5cGoIoBE3PG7baM
bMfBoIOvl1dHbVMOcCU6jXyOh0GMshZr20u4v6tvAKmcbLSgA0rOIQ7py/MPFfqi
mPedUpkY/fumdCCAYGH1MFoazJnAz1CSphKb4tbx0nM1Eo4tGmrM1AzikN5tzxF5
+L8nDEPNDUUXM7CC9FOMERpDbDToYlkU3KrIelPvrMXJDS/R1VkPjvJFo8p0n1aB
F3yCILXWGY6j8Xu4axGq9YuFSBfxo6mmk8Se3ex2YSMBacR/exRflKhlfVGEU1pL
+quMnJb4HEystS+wlLDaKxx4cTYbTC2eVItBUB+8grRU3MpnScWKhSSZ+1SbGBj4
sZVDOfhevTpTLFbphlmlkE/Y7GfSALitpt65N1f94co/+37a+PTO9bFoE1lc2Ge6
bHK+AcfMbEqpO5549eENUCLkNY36E6HE3rJr1jLPLeJTuRJk/AQP/7lOswUqrcWR
S0t1D700L0z1cewzcFvrxj0s6UsIV0BsYk44CH2btYVpe6bProwGWIKOpOWjKwnu
4TRKcn5FioYHqjl09wmRDxo/gbwPRnnYywZ8SZsm40QHgPD9ex1kVu72hk6nVwOK
dYHlE+cvS1kqaKB5hHjIWHQLy8EueuGlj2H/SDj+NGNfuJfCH66+pz+BySBboulo
4ZnsOckuyoctPeoqoCNP7RRYAk1VX/55ojNO/TNRmBTrnaMVUFUWOTm64ueqE3GZ
V50aE1I8J74KaausPXc83TDx9V3GvrMMEWuob5TfOWR1DCOfN0rilmvBlxULaAzj
RB1sjTqMBs54gjPwfYGDSNOrV6DGdQQ7LDP59L+1Eh7+Bq9DNvFmY3UQ7keijFpt
9aurM+bAtgPUAhHUGi87pGCq6Zi4Ky879rMoZ/OUUEiMXSXwdgKM+Tr3pMtGo/0S
ILHxb8xsepkBwIwglxYzEgnQaevwbN2XxXW/5N45iFxldzkmepkARWo/IlJYpWkM
VeuiQKLBtniI1dtgKdiX8hQiUnFJVUVDa25IqgnbyN6TV56pNv3K9/garJa+0nz7
mP4b9aqf30aMJR4db1fiXIN2AO606qND17ni8Tow5PFVIqqPdQIGI3w3Tqwz3jkm
67QFfrJfpZVK8Xg7H2JBFCw/NR4yyVu7OjMIQQDUwzAk64ZFDBev+3JEYQFTyybK
srxdnrCkgK6W/mK1oJ+h82PFHXeLKSxVmYuXx+cVBzTgXlm4GnHqEthXb3fLmqmI
F8MVtOxfRNm00R2OyPBFrhRqdphXlxSggewp5H1g/vELZPmmc1JDEMKDlkMX4njD
9vEdd5SMOAI9Mvh+gXWh+JM5/J0YJthJRFS0an7BPpROPxZyD9YjaMGNJMuGzDCa
7ixirS2IhBLbh9apGSuE/sPc4hCRXGcXaMVY3v4SKNXRbqLjS20b9U2gOMWhxgCo
c+AFYQO3ULHVt03HDwoOf1ugchzELEeFLbKT6FlZGIGRdVL88HHUYFxXHwRRwp7U
kXVo5/RiSjOAf5eM5XOmy87Xr1+s9fOc7T6tXvaJf/u6FHo/YEYkoZepdTUiCLeg
UK6yWl4/H67RIsMII7E8jWcwWOY6lPKE9iHeizmpW6pJ5qdLTS12FwnZJQlpwS2U
3vRHKl/ZFn/DBGKYHk+PziHPF7b3rgXamisseh8Q+fYJQLmug60p2COayj5iEE9z
Eg8C0pVlZHeTM5x+qL4FKTCb5Tn8jlJOEJ3VqtPC/gULb5FNivHufOh8C7Ag6SPd
A9JEFEdB9J0EMG7n2IERkGyg4Firw8mEt8lG3lMtWF9aoB57qUGJWBPhpTCWppt/
1637KDl6umTeKjlTghxFnXb7Ii2cfYRg1hKBXHtF0Iw9HurwMJNiwsphWiE4tm2Z
dSFoc9gMcXn4eD/eZJpEifn7pRZQUCAdzQIgJ+pvtoQqAi9VMaxU57kcGhIcbwsJ
hA2AtHZTYEhD+TYKMSxouLsTQu+2d50qD29YbGeey8YZaL7l0omy7+KzZenMBAfd
2XJCexJlJcDdd+F13/0mOp2//aEqPBBAb4KKi0pgOZZE7HugIVDOrWOxiP6FLCEd
FOe8pqKtqHViAPy0NrN6PUP6LA17EREmsJjWkucc3c3xtfES0HyG6iwQmP4ANSsT
z7sPFw0wPjdPoqT36cv54VoCtLyobos6J1BNo819MGUJYN0MTzS5pSzxAex05b2j
bsetNCOvGJd6CE0cgvu9UNbsM0hbSm2hQDeLVCj+HPkhnGlhUj7Mek0aK/exOepT
mn9LlPeyRTouzlXIAN+trSXcBSkbR54XlsSasPYdNzA7UFbvTXvLn+w1HyaCMD1S
6nd5Jl+SBksY9daWad2MHEz3VDsMMBMpyUT/i03q/6FU6rL2s39IaqHHOZIBV4qG
m0DIB/tfbc862E7VCHL1X+kGkltByF1CLzWbo/C70gJUFn66secBVkOhF2G2gCi5
O+QGiDh0OHG8tvaoKpNQ65XKDKoiGIjxRtVLxej11alhKevlsNeRyO13y1I3L+S8
esgJG+qP96VUSYw130cRnFwbFXfA+k+Bia1CTFFXqgb3/nEFi0npc7I6hj3pTDV1
BMBXOfU1FrmQWhXXJsPrDyZwykcr0QiMoVaLPsK9eBtl+URHf2qAGW+qtZOGsUNK
68/0q+kKIk6p9wUCbwV3YnUdZ6a0XT/Z/SBhpQpzJVS++5YSiY63v7DX7zLeCt6/
zu96XQJc96WdsVpAbdI0BEBnLjVaRmBQ8PHXDqAr8jeZunoB7uUe93CA+CwxZSBV
etxHMx6pkdTtg2uw9UQyzyCKVouDqN/dVlofIm9063NdZRNeteLdnb1+V6aWYFHG
9ONnzDlFMPCcrBuwWqrx6Rt8DssDaimAw2GG4Pf/bRa2OmR33LYnezJX4u94MZzH
`protect END_PROTECTED
