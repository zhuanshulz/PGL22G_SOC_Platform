`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i/hg11O4iR89Rmso11+8txNaTGK2kcBmi6APDXXigiMAD1ilI0GXKQi8Dba1/BB/
GWoNwyPR3uPC74Jw9fnNHfWEtswtPV1IkFhLRjAG9c96Mm+uetfK7pM/fcbO9OmA
lj72Hg09r4dwwgtLyaBNniOof/3sQIzLV+9iiBMgIRyD3sbmDOX5VaG6XLkj8C0X
1fz6i3CA6euyFWNu5cVrRDF7q8tmGF3K2/mJrDQk7+jcC9GK5fYGdh7ADrWPnQPB
R3q9DLkabd50vPwN80aTiD/w4qJpXAuzPmkWmUSxLo3VcWDrGd/2S8DOo28joATX
2lhZLb3vsG4DrLhO9YTEbjX2ZZIOW3d6c2riQMPCwAok4JWo9o18/Xk/0bjii+2U
DgJN4DgW1ml+mTSO/s6O9NL4eQt6b7QMLqStNl0TnyVN9wOk0ccrPVDiBUMRBhnu
6ejDqygYXTFMRNewmavK9Kb6/c3S030RytPCydoA+I8CgFl68RftfycfFGl73art
OCKeR/Pq7OT++Q3tRwGsOD/Z5GUfMRT4kXWzByKtmRls5NNOkwJPluGCKL1/zu/a
03Vi4GaULGipeG90ouJbwkwRKaK7u5kXL8jfTW6e/3M/GYXxl1kGadOr+JqNWzkG
9FQUU4aP3B/zGbyvMb0n9w==
`protect END_PROTECTED
