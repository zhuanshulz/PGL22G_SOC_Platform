`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZ6GRhbUvocfdlKwhj5Qzqewd+VaagK2bceIRxggGmLnLvRGL+8wM9AM14JTi/oY
Ea/gqsAiwzd20Y1Sw9M0EIN/nnDE+ixk7PgyoAKh9MXAg7LYQqAECz+f5DOt/UgT
7SxXYQDnTsZQhJ96jf8CNGCdZkNDVGEw3WiNJgJeCgVEdekt2fOKHUEF4Y+uyZvs
LpUPQxurvxoN186aF92cm9JucZeItT7FuIDm2sk08V1uDDALNg6M8D5VCOD0sGHw
v4sbePVstN/xCwy5n7YLdvatqiV4LU8FEqP74fIpzfWh6Rq5E1Qp3F8QVDB7ni2z
rwWAxRpIZuvDG6458kRJAsEElS/Azt08uj7jZEnib0hcqkQVJ27sD/wNlIrC6ASm
uKKH2P9XrRXSM6md2XGYTFGMXzOEFIHYL1tPwC9r2evn0c9N24PW97fcGaiuTueP
YWUklAlgbq48JYGK0A7dZSL5loJZMH1aWS2yo0DnEcFlAPp6SryAQKaH/vk6qA0a
49OHqjwgMxURzmY2T/2ZaiDnmU3UoQoXja56n7T4QXz4zFdU/mg+hOcljuZZVClB
lgCpc18AjlBW84oI1wj1LCQ6eleTqA8i4hNCxefG5+MfZ6e09Mh7Mi+jC5HcejvR
J1GXAOmoAUS8cH4EU8eVcVIxfy18jkzm9Tez6i8YaPaIDwlSstmb3MhkZ0t2Ffry
/oeS/iWJini//hlfQEQFeF1CyzzRsL4q4XqnvLfMv9XlrWImaeiP536ltBnyJZlO
chs1YHrq+foNVU1Cm4hG+Q==
`protect END_PROTECTED
