`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KrfEn3lcclElB4Ovs20lykt5gxj+hOEzoX0rrwdLRqU/wZCfml5wnNm0JSS7BfK
Yrx/WUZi9OsAJlRG6MDZPK96Qf3YoRHlWQDuW/ly/WrjMWIl19BxMR++Qkp4QFaM
kfO9Oja1qdwEUeZRZkqDCT9QsYW/7n8QlVgkXh0mgKinhAjVdQ2SiV1gBOdbbQDg
iCnVJca5W2yrxybeRtVKzwcFtp9ars+kRoVk/T5ogCRWFc4OQWyLMEFZqKSjgOoB
Dc5TzFghkUyCOTjO9LFKlkWpvI4vrK266N2X8qmvlGEofYav1mSPQy3Em3oQ80lm
t4SSepxep37u3/THE0fe/M7dRACJ9ylGV3p1LuUdfJFeYwqXeBWxmeAf7r1UGmpi
OI69ZLtxWiNYzOEwVxbYPuSgcuzBIlM87BVEY3eHJiK/UZX2nuPEochUdfbmcyHF
yVrZhzmiEtrI1idljrXoMiPN2PbE0IVX5ZI3y2YnS6DWm/Z9TkYNQnhQ577Lje8g
HpXmp6jEIWW2cDzInhOr6qUd13uDCXJilHePRD5ILve+XMZ9Oy78hmtrhNTcccrM
UZb0VAnmQ+D4MkScZpiyoYPFb3+gd4IxTisyd6PziBrD0V3DDyMrIIhlEw/z4SPe
hCmUUnsbdFlONNSmly5vDC95M6iNoRjVofs+QEfE2b6S1jtOFLxm7wp2GAHxHzjw
VK1mqkrVwo94zGWNMBYPRDFhuvClwqSFfRoD7daIp2WsTzGh2NbzQUYqwShjqytQ
4N6s+2CAbgBo38PDV+smdmNoMeHFSYmFuVTEWIT4c9dNF44O/DmtOVyo62BqZiJA
9dA42rbBEoKGijxjnvd2TiTFF8aQa2kfVK4htiXYmOovct/dXEFABt8TUGEGzi6E
RJugGj8+vbsNVxBGXEk7g5AcasDshpPLegR5uf46lwpTTZAyQLhDFoeaMn3t9Wlz
bniScKyhEqLmvMj18FBFyxThDdZMyVTh1ZdO1DHZRFL7q+WJRZsrmhmGNnL5V+jS
5pgBp+w0imvu/YTuvHPxSQwkNVh8xodAgo1jAEvDnzh7auDiV8ERksb315TVFO+f
jQzfH9nveSm3bDqSxQBO3/RhoLTdki3kRJJKyhECAZa+SsmCKmjCMCXSeqYTL0Om
8Nse29Z38PErdgih5yXmD5y+NzwkjlvL5/MuB2NblSURgmYWh95skmaKmTEmkOfF
Zn+9fQqgefr9NJnwL5eiiemLX/Xxu5AjRpHcvutdzcBJ5eDNXKNVpWsnNZJE2EbE
EKDJ24o1oenDcIJzWkuOnaFWIwUUwP+EKnYY1/4A9wuvrxxf052017qop7dUmtkC
nmf2rgNBC5btjoD/IfWVr0iomJHVIcQA+Qq1Wold6WfHIcfs+cU1uPmbh8tpYluV
Yaz7vTtaTRJseroUWiu0iMlPQH2pipimPy6m/SHyDPYtsyYOiyfy4ivkNYN+A4EM
mbBGvppadQh6UJAf8WAVaMIRLgN3/5yrddnVrP/qiyqySU6ANmdzxwhOJrfB46/5
2FiZhflMhrPaaTELXe5FgVsWsKfXA7xBIohKO9oNaq317o1K4YPCthdirGNA68Ir
rw9GRm6kRQ6g1LvdHuxUk+lqq0igxFIzZ+G9MDYPAyS6Ate0CIVdhg4dL+cP2qVv
ND31a/hk6CoypBS9n/KKV8ZRX0psF7GDP1RU7t1kVxt6ZBY+oYPUKHLBEVmdzj5h
9uUCFO4iOXPon9W1UWM0pIttdlAgnI3J5v6dWiP/CXNh/s/HGNhbwrVbK5mOjieq
nYWBnyI20yt1whj6W+Nq9F1NyNNt3gRY2TQ5Wmi5HYZBI0peH/yMJxnFfUxSsQ5r
KC1VK5tKRc0b84NaU6zsJGoYhY3WdsiZHOIdWLuGfnqVVHLLemwNQk94O/NQyO4U
VeC+oMoxk+r5aLwY7LeHPgTsMbWxxowv33G8FJ/2mIcWMmH8RO+BYi/LX2as2i6P
e1I9tSOe1/KlR2h0VUqreoCbRnsQgc+zDRvjNtKKjqLPF+t69o37s7NCC2jdAlaO
a0fl21nkegxn9Fe/A2Ko2C6I86Xo7oIbm1Vp3e2P1gYmKbm2+8/b4E9S31JlPTsR
29t3ksQxIxti7DoT/f1Z1QKbCb0LH9w+6fqc5J6la0NHgtVWLBVxA0OgiHWXUkBI
S8jprQb+Baa5NwzBvRZO9x5NEr2bfinaEPAZkh0+RPcWiTZ8irVMY+NR8T0eTEN2
mvVGidaim+pRscm33BTUK9om4HBDPpUTY1PrGkM5094LLVmc2hyzBu/X7QJI2NM0
0H9Q6Nli4p2gugpipW12nSSs79PaEVdtBLdzxualaju8kzsdhVjgYua5ps26qP0A
BzphBP4AyK5gKN9e8U3qraHllVgQJHNId4HRHOHNjHBqLH/r8jHKu3MDsQ3hltrC
nfF5KoTMoKD2RawMUfD5GhbbPjt2Yim2+AeTOVmq55ATIoIjbRvY0D2A9BJ3jNsA
G8CzsFDlp3Kbxyp0pj3g48GcWVmqJlhqFNwzVCrKf9t0n+daPxPcUH6dyAFy8zzy
n1O6XJHy+q6SRHlh5cY48qNnZ/AnHI7nsrbq6s/MvM95pGQexEJqUczpFZsr/0eD
AABqgUy1VdpMjq3KAd/Cx+mrACXI0edv0RFsIFFpiY7heo2hmzNlTLAFzB2EOUH+
W8J1EGb0pxxk3oOpRCpXmA+C+s5ElAr+Kbly5q0ZIYjhdb8edmch9jGk2ZHrtWbj
tUnjmD8pFqEmJBOHLaEfOP/6HSi/OVeGOE24tT2Jq2GgZD6wvQVUspS6qKdqpbgB
iBIHgKB+GBy6XQF39qWxLzdoc6/gz+lGrPDdCLwjs0UAFZy17KlN7HnlxAcpr0mo
+cC6XDs6XJC3hNWQUWE/ZavYxVeerYltxEfElx8CyfuWfXJXdmn0vcZhywH+asT7
8S43IEHNa4/AP2OqdMvHtBsvNTeXffN/WDyyHtUzEkbtF0OphU8nkkcbGogxRuAp
LfsQD4FzO9fCGJ8GGKpZSQUvbIx1rb9FFG2FZOQ4tlnQsvCXsOe4W5TE24rVAoFY
r3zp09Cq7IkBRQiKoacCFQCoxZVwyQ5VouGxLueHrAWISeBIl9svEuREfTVhtx+A
KLW5K6ToE6+tZqYzlxMO/V59ll52Zxmc07tcWEKlhT3G5btDL5c+SevydErgMZiV
wy0B8MOJUVI3rRjCOPyhgzakvSYodgA41C9HFaJYdcmfwej1L/aET995QOFpVuFJ
WlMMZT/y2qIt7/1D3b6WoNLjSff0UKjsEGiVbgDEGr8rskAbd4sdH3d/PCJKe2yY
VEau7axHo+bf3BxKLvcKBohKDU+/IoQdMzViZF7DX2RdY9exa3dDurjHUICy7a0P
aRANZw5g1BeJeiBzsFXth4D7wsn2ctGZLGuVLxx5i2OzYYHysu6EuJNe5Uai3O01
XbqSe3YXs3s2M+T+rQ/3b1gdMh1KUK/nmjWwKoESUS9+GQYtxQKb0/CcEkcGN8vj
ULetoW2xD2Yi9TwfsVbObYupRGhc/zAqg2ZTTbMAIR0Yv/t1OSTffmKQfvSsKKSf
O6dDntoj7qwmtCyrpMdMVGm8viabPyMUPWbWL9ub0gsC+t0GlBi5L5dLPn5w+1PU
enHDEDeNGLns05d+4+WMjifLW9OTIGBVWKEtbxh44GQsH3lVZRRLA5li1I8fRBTq
z4+rl7VwqRU8rCaq0a3ZDHW1x7RM1JG6NhKAVlrMVAhLL9xAOYIOsDfQtGZ/YdAD
GoH+bEnIw3tOSRwSqQetbooXcPkRGCre6z8gBpuDcMogxGpzjrqMBwSbT+f5ecy9
7xjmMAX47RDKbtYpdloivz11F4xry1niHwtKUPVNc3lAes/9d/1X2+Juej0BguYF
LWLgeFcWRlgMVQJv9bZhXLoOwb5GfZGhKQOKCkdakmFJzAHvqZqgaSFH2ZY/JzWT
uM4aqAVddbsGxTddNPjeXCkeVXanenNfvccS/Z61EKsegQuhaENHqzn+sw3uzie7
B7opYQX0berJMK59KrsnOTkZlw1K6m+vXw10JLQD1rKy30L/uslBz0JM940lBfO5
MXgBUMsVV+8t7Ga9LjFi+/smw/LYTX45KjPRZg2P8zgr9cUyL0sAJAwPNERzqu/g
8zeAo5fAVw1wFDyCgz7CthgJ1WWklAp0hWVBGui+T8kj8GEQxvl8hR0bYIFP59co
W3gRtX2u34U9IbXv/RzI6GjUEeAdNA2x8uy6X6zVztxeFvXQDUYMHEaibYILhc4z
`protect END_PROTECTED
