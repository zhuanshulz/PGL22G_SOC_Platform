`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPzJ3nEnXeHCdwuDWwgEq830q/9Vx16AOskb8AKENLRJ/jWdUnmu18vo3u/jZPuF
Et8h/NwzR6MMpExSoPGmt6XrHO1iDlna+3d9Aid1Zs+TpKyzlqeXkyRk2cWNw/mZ
eGLAue4JsS8QpkmW7n+B+NQa2fjHHbvz4WzD5qt2kNcVX92ajuIptKNkkCnNXjtQ
xlBPW/2Q24LfJ21opnPJ/rzxwlNqNhaDWS36/X6mOxGy5BBt+lO/oeONgB7nuROO
Mmjli6LfskHJn8RRvEzsn2IrE19RLOAlFywisU96NYuegMI72nU+oOk54rZKp736
pL+pH6V0RQ7FGRPrPOBOnHKjxHR9694YwSw9ot/kmpc3g2+RWJkCdFAEp5bf4+j8
HE+BK0T1MDiZBjst6ltyj+y2e++KAdTrr1oepEVpogUTOGdLsHKFDyVC5VtELquQ
QQbPywB8cbJUL/9lztrXomHbo2daCOE+YGV4k8P0lyGYrko3ZVTQ3Sk59gVkpRdb
Iok/DtStgmNink3sbZItlXWF62fPfaW5W63DO47be4fpA/89MSjpaMWlK9lE4UQK
vJ5ka0ORhP1YNAuJ9EbWgSqCT69gsSYLzd75UeVqDdYNiRqcGoXUvcy8v2b1Gu55
c9EdjHUkU8E7utOZEipnGRanAH/1nMSwas2zP3UzeSnrRmSc84ys6/vjRxwWZZ6M
bSmROiy22eWojzcTcK9KcAzEEzZ0uVB8PPZMyMQGMHseNIAKI2Q+0SHVpcY3kRtV
6330we5lL9EA+MX/dpCKIruTuaMhblS/HamLR2OKnZ2JI/2iavPNez4roQ2cqi+p
+qR4bwd83R2kphGG5NYbhYaVg9/4fOKY1bSdkTdGduw5glUr/D3zF4BUi1U+AytX
gj0LDk7HyNCillB2H+Pd+7aSFnxekQsx5k00a5OTyT3SYv59PAF2YBMc3ZZ1gS/P
9HzXz85Q8rPvKBuKkNAHDJCjOc1nNlhzuiMcqB5HBgmwbvTh6e4H1hPfAYKkWuGv
DRuHUo9AnrW95cekfefiCfmBz5nnnwE0Cz77+eTMLPRxD2POS4ITSn+HIcES5okx
`protect END_PROTECTED
