`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JVNPNu/sV6mhOf/89d/nZdj13ZF8qLYApZIMJx5R759wJDscwC369wJI5VCtX68i
HvoLL/lx2yE8hb3Hy9ZZvnMoM6fznmGR3HOrrs3UPnNBggqRSvn2PBCFI3Q4wFzi
d76AnHQ5lqelbp6lxbgQ21kncjyacofMS4vQDsLlv9kDUkZ7lrDP4UepzmrAnQnf
xdACFaePJq/tZAnuDbA4IHpq/CQ6j2+UD+zCXGNTvsjYbStqZbs5bzdgcwR/0h7E
xH4rxQMVM/+d1ZAKJIhMlK7H8/OCmIICBcRwwBm/AGTbyzUOe7irJds6QaKZT0yM
TYjJ+hqBrToupP50PgTjnZDYKEdkrCexYKOztHTVHNCZUuGM3JVJVWFB7QCWTf7j
47rc2buuOfy1myo2oEGIlefR1wNlZoBOpS+yhRa4m+qmD0tEKV04qWX95dC6sQyN
ozGMzHnOffSIANyLRlAQ6t9Z7UHgeM6NJ4djoiQaYLoB5ca+tD43aSLzmeKG8t2o
+5Tt3abU0+I53fW1LtfhlvdpFFD8KwnGsmdzVSbc9iwne0aivvkj9eBKyfTWPWuV
a96NZ1KzbCCjaKKtnCbpSKG8enguN+nvyAXcrI57lKMur7VM5xBXEdUkdHM5Me3d
Eorijf3Lg5Iq3KUcNI3yRjzqWCupv2MY147pmFifSNVWebZU6meMzeC3OGyWAWba
OQt6TjL9kS9eCyh0IdVufNZnFMsSXDxIvkybsnCoY6p+3wtvACrYgwODfIwAOje8
VQ3Dx3z6q9To/jtGFHtfN7ywmxS+KMw8BDXoPD5KssAL+7qBtYfWuZBxM46N5QZC
OJ3YzMGSFVJbzz9KGwK0V6tM1VyfTjIN1SSlT4IAicDJOvFQFAZVTbeZmCzDB+yV
hYFTQfogcFwyoGAgUhAEjSK1VkrkQf1NJmBMDuncea1jS7GzhfVifMmbYA8Yovnz
gu098l/kWzBbDezUtHgGdA==
`protect END_PROTECTED
