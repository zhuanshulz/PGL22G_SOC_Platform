`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M4p9Xh1ld83Oo+HD97qvd6+Nbg93qYMYQUymTchlsj7+FDSofegI1Gq63rqftn8h
MwBJQni/jqmbkVMMDRaTy6GXDM10LPhrmqFVMQPY4osrhtfAFeX6AOLf5gle4naF
juj74qBXHlUC6DEe5xEVYkENwMpXvWBihQm8LmEaElQHyAdjq4IslN9ZQO2zOfVk
iUcG7yehd1IPqe8vgvE+CNx0813Q+X+5+bX9OtmAz9rwxOIgeok3Iqq/OMlFcmaF
Kh+Wm4nYVGjS+8yeXjV1pw==
`protect END_PROTECTED
