`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYGCNWACTS6GcTqW/YUUbysUw8SvkGmRQDJL8LpuwkuWh4+ZB9Gb5xZkN9B8uP0+
pXm4jcZ92HtWYS8lc1jSulDiGPpFlKqDAXLddpfrd1OAXz8hmLAGlyqkW0kJ4iLn
xLSlvuqXk0Zv0pd6B7SPf1PMqARMcOIL1NfrqGEHFYoFMLYcKcCZf3eDy7n0OtNZ
kmh8952he5OORD1IcEKHFHw8CsZy5EFGWeXCZfNjH0RJd9ykibpwkGst4xK2s0ub
v++DIlRYdQYNX4qDPD4V2zs/Xpm23oZxuVG8EYo96cBV6bcbrxOB6HYI8Ewpah9c
pYBuc3rkTvTYy8q5mRfj5B9KcVQrn3uFR3hBgrjQctuqsJkutVZMgD2aaT78g1IY
FaG7PP8s3iT38KYv21l4UHO2QKRkMQV9opZseBH9o38fThyOsM5yGikm12tBKYSB
LIt0o1nC5+32ZWeXg7qtgWtjY9TK3Ly3PRzjWZbAU8rMzbd1Nr9A81OClaHr/BV5
O5uwridNt1t2c/igjdbH3a8YM7iJ9BTWRVUYUpaPu4Si/YxahGVc9C9GSdBJiPYw
+x5X1h3/bsN0JJeX8juAgqeOS2oMFEmpWrDtMR3EzU3dx2r381JXikyIbyXnuOWM
VWR1GOUdSICdqjVxLFCcjWT3GV5N9NCco5rMoCdq1F3RFwQ7cWmFauur4E0BMIlp
XrN0Ovt7JzdzDAFOmE/s3CXRA/UCdOCXGHakiqoxHWaZkCB6D6tJL7FtwQZ60U4m
38cN1BP8gLhf5f3cyszjQr+zH2GJAb0TOCVno8ppT3i3QvWWvtnSFLoR9/gM0qco
KPRpiGnOrcXRsYA7XhUlWbQeAxCwu5+nGTM+DMM4QEYO1nb4qOMf47kTxZpZm6/k
7C93kJu4lRYHoPrvw8INX/h4V6igRud6RAkDGDQD964lkjd95H65lI1NIaS9qXcz
eNw7ql4oXrGPqkVy68XKS6yf63MPcUHJu9Ecbn5jIE7ppZzjZ6REK4TMISiS/zF5
RcbbJEmuI+ShIAn3LvkEUp4ez6iBBdwTdPSbqniZUoxWZrVrxoDxmaZyZih3v6j5
nXTU4iFIXWX7W14070ntI+cVXilwCUiG/ZUrFZey2wCgFPecErwDBv3LJ+7WZUis
X8OanwLZ/Rhkxe3oGLUbBAD4oxcqx60FZYk/4DmtMGWQ3U6BcjUPXOcMP4pNdVgh
`protect END_PROTECTED
