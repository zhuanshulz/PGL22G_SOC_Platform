`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZA+B1j8U3SicMUt1AI7oNHfLwB0cqwMRlyZH2akHeaI+4PbnjV/fIiZ3UX1CfnYT
hzwMsIk9VigFd5nqFnd2EK8FSjDbpqinumBueEUCi1lMrb2ynfvtO4qq1HPoTJlW
jazkEfkaM72psWgw0DYVY5J0LAeFU4jCdNlG8KRoiEKYzcR5oN3q00/OPn1zVHZz
a7GWMYS47D1Tlhbzq3hyclS2C6DJJcLaDErjihkWGV7URNcON3cRGoEmkfpyGelG
kld3vZyim5vXWn7s37epLtfNwQ7A8w10bvtHRAgM9csKQkbhfSUlRRdlzrFMp3NV
OGXQK2i9g6OYbqgAysL8H/Ng3z72OzGvJ3GQ/e/lHgVEjO5vKYnZK1YrQhoL1KRK
hPk7WMQPU7KkiieP6txsC7JSS47I9FEid7Dzsd8PysuLcaYOtEO1NqamqoVvv4mu
5CiYZaXjOxMwQHgEqE/sz/g4EKhK8ZkYWRZ8Ra2suYNWZmxhCTnup7KJKXgqdenH
TICEh8D5p/ovJORhApEvGLypzCLokXTS+sF9b+4xAcqS0jG26BkFNJ9I65994qCX
Q+c7LRvPjkisEBEqtBQRtByHRZo2eNDYhM/fQwunYbRTgBiItlBYpJuPA+76Vo8b
zqeCIoWdq5g8jaeEV2wXkZWw7uEXv/h9akAOMr3oMRJJaJbd6cdf7u7bgDQt0ykP
uniSdC9ZcOO2nrNcPi2yMLpq7zC0abSj06K46mfvXK+Z5067J02CzkOLXzZeSCJX
6hMlRBcvtJfp6LMex1WFiuT9tZEAOmB6yjumpdgPpKOcDueuS64HpR+Uy5BohqL6
EjZXf28N6ofE7shUFjf4jcQGJwp8Rkinxp12A61+L/mNGkJXyaTY2vzNAlTWkiUz
5Ok/LRZKuU2ha4xuiOFr5E7aTUgzDlc5Qf0BUHcuJ+gS5x8hUdWs1OsAEwLoHuf6
uN/NouHiEEMEAV6Ha+/KUaeSRBtOw5BoAmUSxPJBGSjzEKQumuMP325y4a9Pg+br
XpQzI9suCaFeAtsYqX2hRSkHgyAnHSFqzuNRiOZQfLZs2v0lEv8RrDpO6GeMPJfH
EKswyy43g2LybXVjkjQjxJ/DF1WzdEsqIF0GMo2JvNmFJqxDD+ZWf+6JbWwgEwiy
GCVasOgroRGcEwrVReNAgnwyuDVKayFTvM5lxbE8pozRlNoRmlHZt5EF9Z4ASNhb
UK2svERLIvBt9AROBtkUgzy5+6IZKxdQMW2ErFEzaQNMpJSL661AqtLhggYaUI5d
i4Eq99WfDt6otFYRLnm727EvmI3BS90aqRphSmREhTjBvJe4cKeamAhZY8508oV7
ZqH2f0kZOi1tgodHzb5+s+/TCj+MLEhjMMBhx8DkUatUGG/vBf35bZtaXJiKvq4r
yVPz8YCF0iBhN941ZCO6rJp+mcLJ/rNfF89+S5HvVwoPCnN14BPsR7ETQv8s286u
fekVrfKdYXWBy7tsaWO4bonrTY7MqW0EH56/zZChvYBB1jRlUiS/tzGmqQb/Z2p+
x4ZiKvdlYgQSK8NORvgS97JKXqfViGwU2SFcYjOem5iwrHD2iVqQPzF9p2+NFa4F
JoxAq6Sb2Yu799L7Kuk94V8+1mBlAjeVTZ4tgvq8Awk=
`protect END_PROTECTED
