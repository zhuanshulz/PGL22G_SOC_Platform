`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lgc3v1qqe1hy72nQArO4JGe4DEIJlw76fx1fRg/D7no1KZC3OpNOOEHqrzFOaqSw
5nY5op7GiKlzmbuAIcmneNNKJbNItFrB+FD2BKk9O/Zv9x/jBBkaSym/REPK0WvU
bmcdGG7eNTJDw8P6ecCyR25f/s+D8Rzq6tZqwb3yzPSJiSs1WGNV9IWN3KT4jpq6
B9LF3gBdcdEdY/LQxpLz6tcUfItFsC/ZUrqcMzhPfQQDJ5Tb/7iULU9Hk95/BhVy
+n+pGEfVPf6jGyKXo/vmiVIJA0IBJ0P09BlFFcePSE6TcgfVPm/+xsP21zAAM2UP
gHUJj6y46dmw9Ij3m9koGs2ehd1DZjYgM0gbGedjQ2cMJDUaDRmLoZ9EVcjS+JDr
/pphbfmeiJ45pEiEhXhCgA==
`protect END_PROTECTED
