`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7WnSSPm8IIn4bjM4Jl7C8NgneLJkZHJGcodp8PsuETCC48sTTbht2EteRrbUByq
Y43OsBWcScoy93/06B5MVA8ic1AyhD2nmJQ3j9QRXajaehNTm+G/j6HoFAPunXmS
qJ0P91Q1GWeHWOQkffu6d3453U4je+AkRdSlOfIaCqsSV0OsLssYfR7+ZjKFHEP1
g52jOei71uFMbUibpSQ5Tr4iIDPZNDHoTniYkKhLBgPqflDaV6OcmPEHawWyuMDj
h7TypONk4fLgwzgwgI3NK5I+GjLRw367cv8jVdq604Riyp2gr4fU1KEPkc9p8H/G
KgL2gSw3s0ckz6ZocY6L6/d74UrziO8OHtBAYy7LGPwpGDdjnyRm6N/iB39YI2xs
GGpJngURjx5cxNtodn1BNA==
`protect END_PROTECTED
