`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6DVXjT3b9vQNbR2cQVW2NExfoAVK8LE7mFjou/4qn5e6jSjwDysK7cohjOk51Kb
gkB/oEZkVMGoaWjZR9aBioQwXrOynyWBIr3edCjapNCNE7dAPxjj+8IBMtvHY1IG
nsXp21ggfuxM4nb6R2JrwRDB7r+BFOeacO+EAazvZTE4sLx+oh1SRQZZSJYXjABS
aEXu/4HCqlqxEq+AQv6z7xFlaIjdXudb39sQAZAkeFlU51BCFMVqorZ7S2+rHNMw
oPF7in3yYMPooN3RQz2jcwNqGHzgRcjoeBNPvpPkw1jXyD4mrKskChjsTdo1HOeW
rm4ysZmqIkjqtsERi1sFpcYFaZ2W55V8zUXr01wgsgjSaVyCwY0CrecWof3kNYLi
ypM/GG7ANW7AAgv7uBBRkCMsPT1M4cM1mljpQiBzqdflnY8nuSWu56fPBfjx0TRG
febRlMS+1njUG3IZ2FDSDOZXwXOdpJXZVR32iPpkEwNSECKQHFVjDGmFkvO6J2Yj
JzV+IgQdMn7jmGL/6mncHG3Bx5WBvLDptk/ofpQ0hSPEsOKU06vVf6347kR9jjKZ
OCiHkizWNGXnLfE6skILtcsWVR8AvyB/AxVdAVq2tLv5jPnYnZkhKltDBL2fA3V6
yG9j4linrvlsEnutFak0FlqiH7OOu/yQkdI/FSXzNs7OUM0i7edBLVl5W/Ac1t06
kVM4t0CHI2K19oIOOs3lPTzQ37GaLiti6fvaTYXCrZDtOmKEgFuWke8Zo3m2llgq
7LPTGBWzx860bpX6/mYJY/v1ROOADSolC4YohShQOE4t4K2fdlLGBCMfDQvr/QBW
kSWOcGMo/OrFeEgskSk7EsClCQHzwUwUb2tRwaJpjBFBdB1Jnz3dNL23MYxY8J6U
tQMLl+d9mMhdD7t9NGCqHlL6OgHXA7BSe6qEFm1x8JEtDlAaN930dWHCSjfZXzlT
27Hv4srz7M1mqEIeVgb0+QxHykvY+HWfRWOvP/0a7UE9/c3a40FjcUhxnaHNOjED
BkL4Oizb9Aa5LggVL49hlGYMXdpvaxbTKhWyl8z5w8TFc3T82c8p/DslogVCWDxr
pEp9xRfV9YLrv6ifOp6P1Q==
`protect END_PROTECTED
