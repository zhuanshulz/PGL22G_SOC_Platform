`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hmE19p3trhIGCDG35f8tMQAwpZPUbd7a5o8TEAd45XcTbouN04DsSyhO21JxqAb+
3m+QbtfMixHn8sdq5n48vaKLRSclgsxWyC86R8QZpr+h9iPQBZCOF8Sfx4PeanzR
Kd0BVqXaFCjoSWcMc2/lM9sJeQ4nibe0jBmeLQgZTSvwwIOSQr5rPQaLauhpOX1U
FR1iRZu8yreZ1fNLmtlGmKUsDX7g7PExGgwLyfto8ShFC2VDlFG27+N85BO1ujty
UHi96+x/lU4u+O/pGKY6kZDJZqNKpE9GfBi5nAebiscKJ/gpqzGB9+7bqcDvX51U
WXwkMsH7EnxFza6/MX4aKvlvdmKkHSdNVIrvEosYVMjVHQ87Q9ecEbPbw2UtLavX
lbQztgIKEBjXZ/dknqKNZpp/Cqo0mkZ/N5Ft9kNYOIxA7rP0rxT14IB+BTnP5HQ5
2Fd+i5agXJ7Ix/gYE5Ea80ZVQAiecGAHLdqW60IkABVRfVlhPyQfKdVM6eOpih63
s4iVK7yzDxLoyHw+FW75O69PvQOrHygf+KIYHZ5FMTqY3sciqM/V+I4Jow0/hR0G
xqUb3RpYgkVGPdDxXVqG0fUPIL+MslGGsij3mQAf5ymsfNAflnHPfo3o7UeCUYku
`protect END_PROTECTED
