`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7XSGeGlR4fMLKs2rL7/CNwr0Fuin2mQJpgibmXzsDDm2p5c7wmFxuKC7CVJAT+7
9LVG9NWtFP6DnEQxTOYyK2RfxbIlvbmYd0wg8tWz14vzB62Q+F4S+AFkznG8aR+y
o18eujjxXjSLUaSrijL20bpvnSTQuJEuVkXdWUp6bM1+4mOB/8DdvJ8gO5H+juFJ
EuXFOx0JW2y44RZQ0bUJ+6COZbm7AeIUm6ZTt+4+9Bu8EppbhRIVqAd/sLAQ+sno
t2Vi2lUWO7piU3oXtvu9ba+g8e8TR3BKpiWHYwaF2oKfBrkYB0TC5wQq8m9yGe/M
zzH6Et+uz0ljtLzwxILLOm4bNV6+/NFQ1YhjdqvOy7LmSNLD3HSUFQLfjgM7hBJN
ycY/zzCKOadw2vZBztgqbsuEqCfi2F0yn9KIj4MbtoeIX7Vu+khJXwCkn7hQqrjK
h8J2HVZkq4DCXC0j34mB6v8xmYlXhNli9//+/cBUnMQR29w7MJwRqnIz3PonZwdS
RmrPN/4tztvk1aoiI5vJu+H6BTJNn3rBD2VVvAjsbYLYK0pg1dmgsBHP1b0zls1I
491maB4kJkb/aII826ly9CyslFrodFPt/5kI969xoicdD3H+XHKzXtlBoccRdYTw
CyBy5PwZ+jVI4TWp11ABWSmaVlKwcrZe89mfL0lWLZvySTXrtG6dshpJT3P/X9O1
6MjPBsGsOPhY8sBNchoo58y51aAD12VW8Q30wcXzJNMtsa7GJxRWyzlT23wuwnYg
fJmWypbk+//Zs4DkPe6QeYL5nuvur9MdsZnKF7Bp1hVcibepCQrcIFduoVY+apYv
n03ZP8abq1i1Dp1ptUV2j2BJDGaQ5gn3WG4BV+9P2PcMEhKKihkh9Pv6bQUYdTUv
t8P+oq20a8UJHrUNRqGcvLzUeAmUFPAFovxEa2IBpqfkOfCR/K/r5RTxM/hfXQjY
ezaw8cBBU8w1bWXH0+7g4w30kPz0539z/Arww+dzf6er/YdrjyD1Kk8cHVK761TT
iPY7mze1WdirSD3Qjype3dAKLZjC7yeTAVNgCrblEJkWSyRX3e8Dq6tTYOTyELF8
e8xnizKh9p9/QCE5v4s9GbEPltvjHQ2pyXQYASBf/XsBNwtMbrv/MhxuG+Ct8SaM
W/gCHEnwMQO0xjvNCEt5lBK7a6viG6ps0yi+lPYkB8KK+eOrCxACRxbKw4WRWHUS
`protect END_PROTECTED
