`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4U031ZWa9eefzOU2WYGi/u2gWNfYXSrA/yvxK3m0jssm41IzRH1NmRYMg1YrhKU
+hkcVjdnrZhHyD1I6RITeYuhqtF+5+PXM2imLj4amK22zJIqbxKOo0xBphwhj//H
tQck3qkL8qGmWw62f/ufLrdCZUcI+HG8fNT5rEt4vzeYqsYQudWTzOXkyUECgR70
w1+e/JmHsTmqKxAoXyX3Yavw7rM5RyKCfNzx9HeTFNugyRgoMkjCbGTbKzSSM1zy
Fz1hTQwHo4T1TvDS7bFZvtRyfH+gdsb3dCgfp8+ZpVnmgmLw8kXB2SSnyP2kpzD8
zpPts8ciyYlRErgffP6YAJtkV9g7SezLKbOPRpWIWJc=
`protect END_PROTECTED
