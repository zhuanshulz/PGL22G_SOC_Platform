`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPyuBglBXKKlckhQ0sn9LLE5DTCjbW3DF9sj3YCC3HprJsCdJtLoIlbk5/C2wMhE
MpOjznSpBaJ1rgcYkRWSJCGP5Oj12Ni+a23voI1tSYPlaKZ6MpucbW5e8grVK+xY
veShxOnFqjVdWLnN577rP7igNxE5moC7zLRBzOipZZRCYDHTOYYjo7Xgs703RlqI
K3h+Cpsn+sAJ4lTP/2dCJ8TdRg1NGXR1VyBKlFFvy4by/jtRDB/TMhwxQvZoOLJI
FNchAKdQcItcWaPZ1TH/RcY5WM0lXpIyj1E1rSuzylki9PRaEbpdtODMZgIDBlKO
euhdIJvFIY6Afrz2eX86nQ==
`protect END_PROTECTED
