`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lM036+RAgZ2PIxO/jfiNYDuk1CRhVPhoBdvo6BITl/KbXOxIzhooxNejKVN6AC45
pwEAicEWvZe6XLZ3PLprRJhSkdFiZzarhL7oPaEhWgYKtZgENWFC0bJWU/ny3tzz
JkUGv7Dw1gMlGp5IaxHLUXQ6dCfJqQAKrxSG8yIRtkX1Vi0UMl57SQw8Pj0F1R9E
pDI1/JkuF+DNfbbgGN/9+aJI8wdmwevEsrPrFufqdNsh4jwE0LAxzHza3hDbTTeH
1qHF35HsMFvCTr4RtYBeB9ph08B+4jzKy7bavf/on6mpP8l887ZQztuZ5uvu2mx0
Jmz1xOamV1gdFUYwseLbzIzgPNkOBy160XRLc5Knv+d56p2UYXqCV2WwzEqoh8L9
jSlHTjNzZb57HAJYexYKeJ3cYLhAsJOWMRhIMbebaTaMjWEG2zpIYy8cVMyVRXvd
JW8P2iAt0xkk+DqVPo7wTUfeYHnM1u/fxERKDIfIIN562Xevhwszp3vvfKy4eLkz
ul4Gwi6t18dPiYZ5vKsLyyoOmceyVRlsjhUBDma+0ieWLgaNFNH9/VkGQhxrQMMP
wB7Y4n1yHwHe7u+L4rUnkBFrOWbWXHVR996V3DJSQ79HJz5RRzWKexkiEVjXwafu
PN48irG28vCjAxgkqsLDBpxuhpI2bq4kgD0O1AAFxOItFKAS2vVA7dvIdFi/WnIF
6LlG0swi2MoUn4BPYbqepS7F7xpm1Z7P4/Wa4sfBhSYPE/SNkJfM8Xxh8FQLUYmw
kZ9mOM3pc7/ShmDMsSaEtZh6QXbpGADxyh9rfOIK3mTHl6ChM6if3TzFTxfqGN+R
deoqcwwWFtwbt1rIkR1FYW0H+HDgfdT1Uc1UfpYYk2vXh+iCItsplgp7RBLXrNPO
ZvGxl64V6Jy+zGADeeCK8IeRgVMZ7ECE5QFlPsl1C7hEvAmN9w0uWAytgQRZiDIW
KB9UujFmbN1aLDu1MD54UN3dRQ+jUX3Vu27fVvhUJ9uILxgPviFK19StbOq1D/vJ
TEDbzZPkZBuvAFIbVwxowMt6n4A/CnAV+x0D5PECUoyTXkSD/zmQ/Lg0cSprbh0v
58q2RyUOVcE/4xO9MTK1wWTIO9KiaF3wW2FKvvf6JYHizBletq0w9BEAampitP++
Nf+J1rYNFPdtMr2R17MVtGxiqNfnrOIZFv9ZXGqgyEZBmEgQQUeX7n6wS7uhP0xa
+s3OdlqJheJTTckKgmDx/eIYlsKBZGSWgMabBWB5RE7lqm0InLtND7IwxNkrq38U
5D7QOANWBhjTCHE2al0tr5KVsNjpCyhT96RROedLUp6k0Bytneuyb3rZLfPSn9sO
P6VfYaT2FhF6JA//SUeiMMH+QDbQpUFMSVOl2CtRKXEmTwbYhYmYYwr10DR6s/Ai
88+PJ2CxuGAq3KBuUgQw/DwsMI87G+1Wa80pOyd5O+p7e0PkxxXSdNY8m+Vf6DLY
nlkyM4RviO1SxkYC5OcoilGwDaSZ13KnyZvfTM3yXNRkxwcaj8Z+IJ18Zkqzu/Ni
U1hl25ocqCjfSgKvmsjbZAr74FrxUctgeqMJf5ZFf26kB8KScklUbVOUkBUsJ4Gi
2YR5bbuRUPYaJTBCJCIJb2C0qsMAQzLPhPNQqZlTF/X6amp/jSpwu/py+U47iUlM
GAVF/6o6hVrSjST1LP0Sw7xzhsL09ODid+eH2EepZ7Xxbj9UDk6rkW4QvM/IRlez
KyUlG+DSkPHXCnwxKZgNnxnO+gnqsResEqizAHEzAg+vbasj6HWfEqf24KFK0Sz4
dW1zFmQnFg/f6YE/I7xSndxE8aGXw+UjYplzwfYSWtbbNiuVnBvEFSsJtHn/G4ou
sBJr7CAQc3cTEH5888mAx2XP9HijYEGO6dtducrLHSZunWLAKhLqOArIrGqTuQJI
sCDKJM4LxW3+kHSnEEFeSBG5IgperOIF2+K7kWv7XbC3LaaGDp6mJKA+4fHYc1Se
5G4Wx9ngtkqNXoCl/JLCGtPNpagH8MZDUl9n6BG0xa2Zz9z7g6cg1xjlgFP86iVj
LZ0uLdt4t2Y6rIueeRdA2xY+c2UpLdV52gmgIOSRYPkOU+nC0nSDJiXW7Bi9NG1O
0Io385cVxnU5i1ZO6UbT5qfrTIKJqCxJg8zMITEh00C6EzHLW1lqljgu/xs9LtV1
r6FItsqeUq5BOcMV0Gcl/1+iD37Un3aJprVBY98vmZImeTDh/KqK5KKfoYfOwcgB
6gq/9fhGQlNapj5LLQB5/yu3IP3ZH5mEyoKpDuFFfrEsFY0ned+2VAdp3O38o+3W
SbWnd1neyycCWG6hy+T/EZ759BjphLpS0hG8XAR2C/s5wGQeVYta3r3Wwt44/4lj
hF6EV6N08PJLl/TrBaRHO6xZQ/fxDnhcHoBQoFM7O6A=
`protect END_PROTECTED
