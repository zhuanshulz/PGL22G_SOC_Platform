`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KP742Z/fUp4wk14HD1azjAoi6iRaOSFT2SGEwTJnkpiSdYxYxBr+Cdc9rcEcylUU
Rw114cSVZ7cFvBrs7qVP9MY61cUNhVwd+1CTsavtwJrbcXXQ8xd2t5LqM7NGDJj3
9zVywjrUMrbx8WyfHc8hn6Axz6Sq2F+DWl3iaCBhmzwyH0JIrPHPZfj66nEf66Lz
9XYoRbuZKT5Wq24EYkZgDtlKCquagdcGll0954SopeHF8Q2acJuwQSPaGL78MVhS
lvkpY88KgMMxCJevWOMX9vuhX3pCBstIedv+hbGmUBCnNtTcD61o4/9cFrMMpmE2
GedMtNOeYtZ2o8b34KTbVhAHcoCsnSi+sHfaqlQmp66hVesIvewN6hHt0DiTvSKb
gzRAC+qJAB9fv2+kCMPtlIa+KmxxTpzTGCv1ToIUbiWh3v6/JQmYhBRdeoKw3gUT
QDnC7KORSPda1KtZCl6GCAmFtCLjGfxpijL1m60js0vLc2JIui1O4hRpXrpbopMY
Ie83jAMWNAHP1TD4l7jYhDH5JLn5eGh5MvLlHuHIuKDN0s27q786GJBu1oudU1CL
AQUZBnp5mED/r1B1pUIzgLYTYBua/DUiMYcPWkjMILa1PeKUfXcdzeguQBMq7mPO
jZ/yFPYFY8/+fMQW9BEbOzDKysjnEkNGQ+1H8J0XuM2Od65VNckQY4U1EBLsU05W
pNkejM5UU1+FF0EbneqdBrmLBzHLBbhYNAOin2my3mc9pTadN8roK6ybYG7sa6yo
Q7PImCwMkV/BnE+aTjk7drLnAZskwGfaWp4vKe3D41dR0YSBjhNYdh8vwi8SM9ao
Fspm5ph9/LBLb+xSd/EyvGdoR/W0xMEAUYBw6TUz4dPUG2Anw1IZqDo8V6H3EU+D
MAnfiSzBUAVrQJjbXabRboajCPxnAb/1TpvRqvR8jkcCj0UI8SmJZw8F3d8mkezA
9KkQqcPASa/7AN8KHUsETNWxxf0yKSxRJ4E2+J691DGKlqbpW7nuEWjGc4f1XYpq
4h1hMkzzvZl37wTUQk1NCv6Yyy6PhcaWZn3gKszDG0kGXTYPfCHVuJzHGoJ6ePjk
iwEx8QMwFFkliELLAiwJJZXqFVuaNG8CitV0/xFeFRUNf0grFM0NeJx7SFqJ/uHO
XA7nYEY8pTBLyKwN3ADaMpPvUyFSu7CQu85EVOe1JjbByWfSjzvXty7tGn7nu+hw
qZ3zdYHPC0iDHoLaBrnTDsdKf4SiKPa7N0/QW1tOS5jLdZsHA2MH3leqFWDqmO9S
b35YsWak0uewQk252imdZApgZ/syGtiVhpQYd/Ew24qGKIzt3adZ0YWXUXhIRiI0
IYG4qDiFyThYjbvHl6u+6LcbH9R65trO13dMDgahavGg0hI4fuhgMSB0qjQCnWXQ
tCXq74XVUt6YO0mkpBZgiRY4YvfMf2zyZE+pu0U59rSN4QvVaCugJsqJ4woT0sh6
R1lWAqnXyVDp/oP9FMxXK4qcxQFech8LYs5W7OhZ0+g+igsCMq8dk5FE3xGEzsfV
BZxdp9RDEznPxuY7k+++sk7S5Lm1qJqkQ9n11aZkvN6nCZqCg8jdTuzYyM9k6vNj
I1Q9LaYvVBKVt8vUNXlKxACJCJL5yS1x3u+ViRYYVZotb+u2dmKiRgEce9TsJzwd
QwQjR2HgcfpgcAklsKlyPle9v6LzsGcCp1D33YoiErWyMSqGE+FENwy7S60rUNAK
R8Lkuwih5dq8rJkZTfqFEoU3R2ALsCdXK54F8TG2aJkvsXSKxvWMz3C/R2j9ZWTI
UU06Otat8ds468WlM6bDsmt5n2geRSgbF0O84U4FDNQhAzKyvdoQH5n6igedSsfG
Ia9Hf3g6UQiGWONqvXQd3PM0KjJUuUzvXiqoqIZyR6jE8im9ygiU77dEKOpTjpyr
Sqq+kpMwRs81BEqP8Y1xpfzvUGd5J9ueumq4a4HY4pT7hEZeeS/+CRXlO7A3Xq3d
Upr+0cCOPVv3+HwlwqqxMoi2P/yY42LnqSrwu/jk5ZRC/SNwwVItfPbW9osBJJmd
NxGAetJRpagFahtq0Zu34dFlyihkDBcdpxvYruWrxyORd+vX1IIBfWAG0LPQT1ZW
rUwHEmWmgJiWEv+1RUt0y7H86NqirTc8qiMaBqtsWrlCvX3zNowY74sYJvUka7KH
b22iUSO6tPP0rkOIu3LhHI45NSvnvUMj15SkdeQH/Ov59y83QGiLnmWj15PGUTBl
u5v3fu46Txic6FSDMvGljUtEO8X99+WMT8Z/KHky6JSzHsQenVSFfA5HV6dHRxR4
780T3snuqNqD7XkoWRfeQeLChJkcW07yv5sZu/FcnodA9dovDYEIRSHTeEs8PveN
DHgqtdalWaAaM072xMyS00necEaxEYk7mOiYtsdvjBHsuTPtdbQQ3hIN9i8+4aiM
ZPfemv+nR4CotqAeUxdQGTeHXjplQsThIPJjuG1bWWF9NJdOcyAoRaOgtJJf9rHY
pA0WO/54qJlhGzECBfPfrg/YzLgLpKSP4hPj+WFCwT6di+apDgmmTlcX65V/jHrP
Mv/sWsOX1WZ3toJQK5zFK00FBF976TLYrcq+XBnHoGgiJUz3Z8zhMsseXaGUWdHK
CPWIDeXiMCz1U/zN7uku3Rpj6k4S/xK60mMV8+Rxsa7Llz++XeV3FLuRF093axcH
Lx7vbOfpoUi1iLk6X85ibGXlRMpTYzoOnMuR4JYzIQlHWELn7FW7D1K8VfgZBlAm
2WBd4sKG3cQnSSxas4VCViVzrDKfJk8fAY7oMGFMkhRHc6INOR66UpyCYgpwRe0N
H45/PDXLaIJiIbeVlL6aL/xGq5wWFNb+k2sSIrnnwYB66pD+2I58DFVHONoFSoie
UsOj2XOJjZliuXYQljLdFg0ooweYBzjYG+wzT7HsgXHLmsT/RJvIPWHtz+eWqGgc
8EYPALC2wX7yw6oRPsiHejTH4WBRW353ito1sAsm4qYw57fmaLvULVvPy3GD5bYB
xaHcdONWhzMoJKBSIJRQXLsUIuKA4XFy1tpFAntN1nso7iFKZEzb/NyDJigHFaiY
mWDnXQcm0C2qjItu2gtSf3IRSWgf6gHCDMKzlbQX7PjRhQWWQIdGpn7jH3NQT9LC
cL3vfp4ZaXpLcriQuPX7+nqsj5wnHOa0IgoPWZnAuHmgzg5FQQtdo9tp8y2BCaAc
4z5lREDp6FdHHGVX/A9q4o6AEBOT2Wm2ZG6pijIO62xJL9eElQc0v0W4sEAxk3Ii
2h6dz4Qyqrzy5TVXe/3tR82NRppU1Llk/+AgfsZkTNGx+uWJgiqfMNI0iWGQkOTH
nTYoUoBUl//9clX5YqE+NxmQm8FKZDmFDgRANMDJp9wwGDEM/wB3BJ5rfyAMaAD4
ZfkKpVZZ5Ys51rG6NVaP3EEx5PDshcsNueD4GYtzIUhDjLlK5jCGCXEC/iUu56pl
l3nZb+k4udP6Kj4/REFEPI0renPSrqc6lmEEYcvQnJANlVaxJ8KpkAizUVfhlx1b
nYVy5DBHgidC71wHoFWwDJAAD4PSFro7dkM22BoKillfxugxIHSRtPnUVsd0W2FG
sGmgfyXD4msVxjvYQxL17czSLUvW0Vs9Ez8c/MjHe7zUc4bZai1zhkyPM7PhgPf3
nUZj20YcIW6+SpQrkuO26lt7b/HdAeF226xXZ98YJxAijDimn8kkPDfg0jGwPIPe
pSqdxNrAYe+yB6GgAmRdZuLCoOU07D5kswUDNm5uSFekn0HIBRa2bp7vCUGkNNJ4
xbhlbS9yW5cppEj+eWBCDQ9yIOHrMYA33gWhPKwnsZFS0s0X0Wgl60dUIJXQgDIr
a4Z6I5oN4gMe+/o5O5dE/M4NhO5I8DU4fb0jV1W3xkHz1MOKWqgZw1Kl9x/WWLxY
jmRdoE7nXESCuEOvw9hM1fCQ9eCnNJ5S6ydAs4GBLmB9+9TxVwa2Asyeyl//7PIR
FOyMB8TZTr8FBsOEYjFLX6RxDnnPEQmtqGEJ98FGV0dk+qzlyGT+nJn8swBBZl4F
wve48YnpCwSyszMGQVi3voCOMKU446568213c64UTv/0qHUlkya8aOvcDRSz0KUM
OUPlxEIDZq+IeC36VWfqMo9ovRMLRik+BQCYMktJcGestc1lf8KXgrJKmcs5TPzv
LVU6weFucilqGfbxsnxAeoK+iI/DRlhhgVIfql0tAW7eaKq2fjk+GGpXY5u1PyE2
AmcXvvgsZSzvoJ8JP3HVriX5fVV5rU+OSAApsZji34dQ6WqquyuRUBLK80bkTX72
JKIMZ6xErL5IBM8KBTdcjTunfKzViZPV50Xc0itPFA/xh0e/DqAyIlNji31PqHgV
eBpXKaUB4kej8+kAM5fapPK2pEqq+wMndgKR2azaXCFWAgYt1/oqChVoZMXo/t+Q
S3AIRa4RuI+hwUZQvX0kvnhAReWJtlVOdDG0foZk6e4RoXAg5ioffLsdzbA0ZsZM
/NkWQnwovDAO3kfFMH+UtNCOMBBMq18kmclhNh2Ew4ooBXYsIqQjIMEg2D0xMi4z
tVgCNlYSTvG6nd9Cf/3pqZFuAxysecCrQ/38aJLV4PGOVfN8KPtu77bdbLyH2yBi
1wI6JvtAFDXOMWYBE/eQV6NP6cxSUM9yQM2CkR/TSVbXt7khTpWss9ghkDbjUoXA
2Vi8nCKtHZPF3Xq3eizU5e3xg8Z1h9xMEFb3C3O1kuEYqyckgj7BgpS/vbibU6Mp
4JHmvqw0YDESNBB2/4I2B4BzNkJiFS+nKJOou03jSLVBLAIy7rKpU7Q5eNi4KTQy
HeeEFRWvVZhgKn/4Z4sG6PPJ1R21/SQo+FYGqCVEXGe3WE9CqB60nvKsorCdVb9u
VwWyf1lBBtDTv7/j1kbjUBVETUjytOOiDRzkzpMSK9Ik+6T44ihfj+tqf9tzWmjQ
dwoybbuRIy3ekAfDCP8FgTbpxdoKUQdb9JOpiFBS3fhUmHMtUDzqZJMdRPv74EtO
LDGra7YgEYTlBA3OBHigyKuUx8xEPUgLkDKrUuP1ySojJNB0175FGylJ2cGXnEKW
iC8+8oYGtXsQNsQ3rO8DZ8jDE3VA8/mN7o80q5DQIbRopjxr7HccsNcVDvJXbCGc
WA9Gc3PA2thQrKMwUVRIoglp/nzCjgs9O3X8tD4NJZpvOaDyAVtaVy4oDBS+uCBU
FWWZBJDJKkVp7CzXV10qo2ikBTYabWnMBiEMHDBrvW9bMHtBrirUDRmdTIx1FryO
Nz8tsq14vd/KwXEnp13YqiD+YV0e2L5OXjufWZ8E8DOySFZ9Z+h7yT5+sTnwdlOl
S+CVaAc9KnHvztGpRxRqXHcHt97BmtTqCaCocHwoneH4TY3tRPBQblt/PaqNtyzM
vV3pcEXgzQIJMk2V0L83z4BHiE6C4WAbc62Nggo3iTv+Ldsyy8gU6Z18JvhxBIXm
Q8cL/pnBE92hW1vbNZHr4pJJju3yMPXwTvFXQ1WL5eFi5XJ5lcxPiEsBBLl7ETJU
mGSUy4PtSnXog4klcgiqwPBZDDvRL7fur18rf+GanNwqjipacIC4WhuB4kqTNDXr
NXVDb+2rPFbnSS4wgk2am5gK16cLsT6I9SQeYN9FD0BeJhjJCYroMh1mmK1PtG/K
537gCWjCM6+KpWFeAa0mKKfQj1Yju/6L/wDUdLYU+G99m0/fg9Y7BT2ocquxK3MZ
mwOXnnBBqeIj/G0jvJvqc1REyMZ+bN8LIsWp/ftGlN6xF2etSxyzX5Fshszz6+J4
gJl9JAZr0NL3iZOl/VKqpykJt0puc3SlcpRJTgrTi8tAgkEfDgt+DKAoJzUsaJGS
Z1Wzy7K3vhuVkGUp4qYzcOfy3lfNo2Ivx22UeNMq9lSIX802Y+bSGSknFBk++TQp
RjYrLGufkbhN8LAabOUKypVsy35AXAVFRJw7VImQnGTm+zBolEhX9nroP5Aqr0x2
zzTHFuvQFuOzf+/WwCTD/V6fgBTsRpeg2CU2jpGunRcfEr/rfzcZHpwWtwOPlia3
/Kx3R83qODo6cMvjlVWvkPwzQDPH08k10o3ZPU5lMsDoG93YE2NHVJvyIgM0qcom
LfA1i+k7wpf5Z/ZKLlooxY+FImLJeaJ5ghNaWyhwbiLC3/YcEYNZwBwv8QYH+JaV
zPFoo0jLcojW41dYJ/r9tlWbQdqXCh8WE79ukVPtfFRZ7tiBY6lDfOMNYMly3suJ
ELrglP9TtPWB+CxU63Po5TqTjyDYuG18aUtPXnklWgwmqq4d14y4FGm+5h/eZAV7
MevhmZMilvw4m0CgssxIWFnj/TXSo8cVxog17fUyAW2PlfgCLGStAF1RFBCvQoET
8y2cE50aupMdkgIPQ322rEsB315owz4Nr9YPXgZ2D8tugUXH7Ax4frl8bN1RqO+6
f8jpBa7WIgATGhvVl+CYk1guUolppRn1zFPkYYWyy3TL46yM0t1mhHHOCrQbZT3+
zcAVgkWLNP3SWYXf/iEvtIaCR6lNUWBT+muXgSHDRl2+2t0bFM46gq8BW4d1XkY/
SKt/L2qqWvDEHyaGUbJwgVBa7uiBSCPesmYvLRUYDwpOg+yAk7ZZYgvI15b5Aitq
J/yjM2UGgmHzDohvYBtXC5ireBTRLyi9mSnHv7Agq8pqHzLq9QCG6bEFDv/uR786
G6pLqjqo1xY9xLFfPRvu04D9ls6hI/L1/7QwX8Qp9uVzm+BiRDyf9Uu9re5Axsao
h5+aaQo+40hpVdyy/E1CgJeRb+9qbgaf7vsB9hLsNlAdZbpHhkZtik2i/o+qo8Nn
u5IWyaZGuOgJouKBoBlD4dpxiTpHTWfTt1agFplg92q6J+6yRBCUdtFWvknN37k4
DqOcLJa139nJUGLy8y/4B+lyI3yhBjkoSWivN7igY5VggfMx1QDSb6ISMYXl+022
0zi1rs6giCcQa5GrUg8DXCMAjAWdn9oX7+3iFAWnK8RxCiEdIP/YI6ERrQxiystS
lK/UczLYEsA3K3HrY6T00G0odM2kFfC5X8GJlSeY341ZrrIdfT8Sy4XCX1xY+knS
Fuil9+y63CkUk3OsjepLihg4/1RXzcKdH0N3DfOsgi/YaQjA5CoW3qG2NV0zrs+W
HMEnac2O7uWcQ8c2Y2Vff/i92PxVsCoW2j3L6py3hBqnWd17XwxI60/juTYXAsGf
xU2u215d0ntq99B15iPtGGGnHvua87xgRyXk7FGbdCj2z7RET9a/GNpJ1H1Vqtbw
w6taK7+uamfml6OUvyx9d71IgsYEZpT2ZLgLGEOo9XnOl45mzRYiQ+X0HZ8ApLic
/XtvULuThVsMYTjtI67d/9sgzmevXe+mN+TVcJ8XvT0G8MOjMwKERV+DJNVZfhDd
z7Rr/r295JDRbtLcQopuE2SXlKtXvmCW43v+tmL7l+7NXC08DYo4OVrv4++rEU58
MfRJUNM1LBaU1DDcABe5rjw9rbMLS2hmFtWMmXHiYkEwjtjqn4tMID+pdeKoPPy4
lfTzi/p2xpcwDWk4zM/vhlE+Hx61sRpYlhlx3C/XDoncSvqPU+1nPW6fPcC7f7y5
ZRbEn5r6R0/D+iFC1gYNOE2HInCbb5n7PAnI/cHDSXJTCAAhBE2B1QzGk5N4OKLk
A/UyK/UYt7UzoUZdMCYdlxGfWb1QlwYBNytXzHl+xNmpH7+ITduDcsPpesa2L407
rX/M7ARh0Uwd1tqjxVs84WHoo5O6kZATnCN0eC5koSfPmvKOcdgAREd07zi+JYVJ
amiz3GJnw6o86HLgyTTZIuc8XYmcIsyhxQN8YfMN4yb0GL1rLaU8NG2oNUjFewJP
pmyDbIBz/TPcmqDwJTgkFwHr+eQ4EXhgtjLj3IDqKdHvROSiSHEQIFUcGhQdB98p
LwNbtBgdgMasK4ar6+LFfTqoAT2Xui9yNlysvzJEO1Cj0JgxlBhO9uPi8Tk7bYDU
VFl/93JVG0PJllfYALdyNaKK1q7Dg8a5avMyxxujr9R0K3AOIVGEkJ3nsGaVzPiB
tCxyrL3hih5lU3uT0y46ALkFEtQ/ETdnKpK/Sh6szEX1UMXvG7HJSx5ZpnxVJhQJ
LuvcJpF+X5/ZKmzmVRE5ESWJu4FQMbkpsi95hRRiAjwcoWugnFtpSLRbUjSJZ8tO
97aAV0A3DbXdMu+jEhTHO/CmtZkSAS3KEU6gW/v3VgfmBE+7AfkEc2WSZl38vKNV
TGUG59q4zS0UEP9uNULsRFoAGtwqLgp2p37QH7W1sceUdOJQhcZa5UigI3vtFWrw
e9pQUPovLxzvFmcf3Drq4wzHJW7/H07qHGnQPQNxaf9CXg7Lb81Gd3OedQ+uvo5p
Y4gFKzYUTmWQ1WMNaonWv/ceruHnXI/LaXzc5W9L3n0grqSDdeRNWpj0cnpzdUKc
nALR0BTWXEth0zKXbgjEaLNj+LUf3j/IB5O0QvQy6kk/RR0MYy+W45EPkoc6KxO4
EvpXyvbFaqXVDjHn5uxIA+mZliv5CHv4AIJceHE5N8KfoASkorJavCBPOFKrrLIQ
89pUFgQNCwbUMDk9LUqDqXEo4ONHCwGYqXa61zl76CCnwHZaQsMx5bhl6rAz18hA
huv57/yN8PvYYGHuqzhOFdaYqukwqDX+2j1pfJGIY5HlGnBunUWIuqVfGta+8gIp
XEppEnRLhexYqzrIQy3A1T4E2hHqPKLRquK3OdIe8GzOHMa7XKLRGa8XAkSs8Qc0
yCO3nCbIzblLFtuqAdCZrsShhbIvlRm7svMMtP1jczRVB2/eFw038OYXyRTZUjvI
tp2JHQKJb2AYe39u3r8BKac2pfvpvl750b8BFQD7KScYH+tTAwqpVH481A3LhdKT
/75w77UscDVyYkq8IY/z/9nEbGsD3ZxwvaQfxcf6U29Vlq4xTkojkVcwrRc1s5oA
PCavkQ3Y8HbL2wD08uhtjPU/EPgk65wlpSBn+hPdreS0/CF8FZtbiGggLLGZF8kR
O+7XgMFTMyCblMyyBO/0QTd/xWZmY/Ujq0m8NnoCEsCQnZiUz/4wzqlZ9hpzm9g+
4cQ+IFhvSbUC2dS/hPtluw==
`protect END_PROTECTED
