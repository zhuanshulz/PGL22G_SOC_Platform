`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7B6GQx724LvSxeavxS9VBb1UuQuyTYDmtgoHwbGtBEiTidoTNcJz5Q5aXx9lB8Ib
VMndI9nRQ0eR/t/3pasDGAsLNfIpYyQZgLSfUhxDSTbBAIJhiC7/TpjfId3mgjXd
yGBUglWSOlWCLcR9OlWo5MQUaoidg/mhYZ2Gav5QGzmDC4NsbFO3eFwrkCCrnrGl
F2715pTwnPCybfLd2mezHacf4wP09SAzXgx5+6giZtameo7amASfmyO82cqYPmZO
+ss8NnbwvpSCXeOAPCvcbvs01YvMOFoiQr4w2+rE+LjWQ9hEhzxTCde5hPtJ05yh
MgmbqN+vscBsGr0FJ4SR+flaoc3L4A3dLmahqEruQAPBlp2V19TZACTEDMY8F/6Q
zaX7j/agWH3XvFtD3b53zSYy48d+0vuytoOc/EG5od3XHkfMentj61KCPpVZBI0P
cMh/nsMNnIjGc0onAX9ssRlie15Dz0LqmKUSiyCr7BdeWFOJ9ndpqpMLSdlaee10
fisHFicrT2XOf2IPGGezhq3ePAiWpvwRHFoyRsD6DD1UvXJaEgl55MdWs3aVhcrf
08P86p1/TFL3RvxPw7iE4yacb5qH4GAzXJusFXBhatTZF8KV483DoP+sRX6eIkgb
ggKf4acUCGnklX1ILYhOw23jNE9o45+asWQasInMnuEzutrAt42h5ehc6Ehf6QVX
aSCnLR42QS5DbNS8+P1wVWThjpAAj5kDIV5JgKLQcNe+WOrYkji1zGvPW5y5maUH
5YKWnA+vS72rjOqiEcRHY69+7vIlEm5VGKIFqtVp9J8QVZ9C7/f4e/VJ+xuI9UPI
LxGJZ7F2qBasNjtzdgNB9hAuSn/1B1AieElqiXUC+CMtBdImKpCgcqRKDWWg0p6T
/79SXiqVbE9AR1PG2a6Kgr0XfROo+1MFxA2+cZZBeEknjE2MLbPJjpautZ89tIez
MktKy5UfKB0fr3BZ2l4kQtu4cQd4n2jqd2vTdr9QdqxEo8D3//s3rkJwzeTV2uc8
PG+TlryfAtMSA5+bvy+kmcS1x54jdo5lz0BLb+n/qZYtVH/XYVZdJIOOXqzehR3n
A+z8nZtxomDah71MmTZrEcmmgwvlnyyNWAYDU1GMJWtnU5UaZ2HIyq9Y2Z7/j4uD
aQZ/e6RjJHK8399WYgziTia5F7MEFRbRHrgRJcFsnuVcNyHHgP5UGvZ93sNAforW
piLUODkonaKQQ71xxzZuTMUFuVUquiz9s94pcILUZDOWoMj7EJCpsSWxnUFHAXuj
UuDZ4GTzu30xdQNJ/hFF8cJ6JwE4awVtEf3ReE0IrkQP+ovZb7n8okBS3Fy/5ciw
zvkiC4DAqawx8ERU8chY6iwDCaO43qRQxSv4IenmeaQ=
`protect END_PROTECTED
