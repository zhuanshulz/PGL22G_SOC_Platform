library verilog;
use verilog.vl_types.all;
entity V_DDRPHY is
    generic(
        TEST_PATTERN2   : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TEST_PATTERN3   : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        T200US          : integer := 54000;
        MR0_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        MR1_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        MR2_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MR3_DDR3        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MR_DDR2         : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMR1_DDR2       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        EMR2_DDR2       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        EMR3_DDR2       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MR_LPDDR        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        EMR_LPDDR       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TMRD            : integer := 0;
        TMOD            : integer := 0;
        TZQINIT         : integer := 0;
        TXPR            : integer := 0;
        TRP             : integer := 0;
        TRFC            : integer := 0;
        WL_EN           : string  := "FALSE";
        DDR_TYPE        : string  := "DDR3";
        DATA_WIDTH      : string  := "16BIT";
        DQS_GATE_MODE   : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        WRDATA_PATH_ADJ : string  := "FALSE";
        CTRL_PATH_ADJ   : string  := "FALSE";
        WL_MAX_STEP     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WL_MAX_CHECK    : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        MAN_WRLVL_DQS_L : string  := "FALSE";
        MAN_WRLVL_DQS_H : string  := "FALSE";
        WL_CTRL_L       : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        WL_CTRL_H       : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        INIT_READ_CLK_CTRL: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        INIT_READ_CLK_CTRL_H: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        INIT_SLIP_STEP  : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        INIT_SLIP_STEP_H: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        FORCE_READ_CLK_CTRL_L: string  := "FALSE";
        FORCE_READ_CLK_CTRL_H: string  := "FALSE";
        STOP_WITH_ERROR : string  := "TRUE";
        DQGT_DEBUG      : vl_logic := Hi0;
        WRITE_DEBUG     : vl_logic := Hi0;
        RDEL_ADJ_MAX_RANG: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        MIN_DQSI_WIN    : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        INIT_SAMP_POSITION: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_SAMP_POSITION_H: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        FORCE_SAMP_POSITION_L: string  := "FALSE";
        FORCE_SAMP_POSITION_H: string  := "FALSE";
        RDEL_RD_CNT     : vl_logic_vector(18 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        T400NS          : integer := 0;
        T_LPDDR         : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        REF_CNT         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        APB_VLD         : string  := "FALSE";
        TEST_PATTERN1   : vl_logic_vector(127 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        TRAIN_RST_TYPE  : string  := "FALSE";
        TXS             : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        WL_SETTING      : vl_logic := Hi1;
        WCLK_DEL_SEL    : vl_logic := Hi0;
        INIT_WRLVL_STEP_L: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INIT_WRLVL_STEP_H: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        DDRPHY_UPDATE_TYPE: in     vl_logic_vector(1 downto 0);
        DDRPHY_UPDATE_COMP_VAL_L: in     vl_logic_vector(1 downto 0);
        DDRPHY_UPDATE_COMP_DIR_L: in     vl_logic;
        DDRPHY_UPDATE_COMP_VAL_H: in     vl_logic_vector(1 downto 0);
        DDRPHY_UPDATE_COMP_DIR_H: in     vl_logic;
        DDRPHY_CLKIN    : in     vl_logic;
        DDRPHY_RST      : in     vl_logic;
        DDRPHY_RST_REQ  : out    vl_logic;
        DDRPHY_RST_ACK  : in     vl_logic;
        DDRPHY_UPDATE   : in     vl_logic;
        DDRPHY_UPDATE_DONE: out    vl_logic;
        PCLK            : in     vl_logic;
        PRESET          : in     vl_logic;
        PADDR           : in     vl_logic_vector(11 downto 0);
        PWDATA          : in     vl_logic_vector(31 downto 0);
        PWRITE          : in     vl_logic;
        PSEL            : in     vl_logic;
        PENABLE         : in     vl_logic;
        PREADY          : out    vl_logic;
        PRDATA          : out    vl_logic_vector(31 downto 0);
        DDRPHY_GATEI_H  : out    vl_logic;
        DDRPHY_GATEI_L  : out    vl_logic;
        DDRPHY_DQ_L     : in     vl_logic_vector(7 downto 0);
        DDRPHY_DQ_H     : in     vl_logic_vector(7 downto 0);
        DLL_UPDATE_ACK  : in     vl_logic;
        DLL_UPDATE_REQ  : out    vl_logic;
        DDRPHY_WL_STEP_L: out    vl_logic_vector(7 downto 0);
        DDRPHY_WL_CTRL_L: out    vl_logic_vector(2 downto 0);
        DDRPHY_RDQS_STEP_L: out    vl_logic_vector(2 downto 0);
        DDRPHY_DQS_GATE_CTRL_L: out    vl_logic_vector(1 downto 0);
        DDRPHY_READ_CLK_CTRL_L: out    vl_logic_vector(2 downto 0);
        DDRPHY_WL_OV_L  : in     vl_logic;
        DDRPHY_DGTS_L   : in     vl_logic;
        DDRPHY_READ_VALID_L: in     vl_logic;
        DDRPHY_DLL_STEP : in     vl_logic_vector(7 downto 0);
        DDRPHY_RDEL_OV_L: in     vl_logic;
        DDRPHY_RDATA_L  : in     vl_logic_vector(31 downto 0);
        DDRPHY_WEN_L    : out    vl_logic_vector(15 downto 0);
        DDRPHY_WDATA_L  : out    vl_logic_vector(31 downto 0);
        DDRPHY_WDQS_L   : out    vl_logic_vector(3 downto 0);
        DDRPHY_WDQS_EN_L: out    vl_logic_vector(1 downto 0);
        DDRPHY_DM_L     : out    vl_logic_vector(3 downto 0);
        DDRPHY_WL_STEP_H: out    vl_logic_vector(7 downto 0);
        DDRPHY_WL_CTRL_H: out    vl_logic_vector(2 downto 0);
        DDRPHY_RDQS_STEP_H: out    vl_logic_vector(2 downto 0);
        DDRPHY_DQS_GATE_CTRL_H: out    vl_logic_vector(1 downto 0);
        DDRPHY_READ_CLK_CTRL_H: out    vl_logic_vector(2 downto 0);
        DDRPHY_WL_OV_H  : in     vl_logic;
        DDRPHY_DGTS_H   : in     vl_logic;
        DDRPHY_READ_VALID_H: in     vl_logic;
        DDRPHY_RDEL_OV_H: in     vl_logic;
        DDRPHY_WEN_H    : out    vl_logic_vector(15 downto 0);
        DDRPHY_RDATA_H  : in     vl_logic_vector(31 downto 0);
        DDRPHY_WDATA_H  : out    vl_logic_vector(31 downto 0);
        DDRPHY_WDQS_H   : out    vl_logic_vector(3 downto 0);
        DDRPHY_DM_H     : out    vl_logic_vector(3 downto 0);
        DDRPHY_WDQS_EN_H: out    vl_logic_vector(1 downto 0);
        IOL_CE          : out    vl_logic_vector(59 downto 0);
        IOL_CLK_SYS     : out    vl_logic_vector(59 downto 0);
        IOL_LRS         : out    vl_logic_vector(59 downto 0);
        RST_DLL         : out    vl_logic;
        UPDATE_N        : out    vl_logic;
        DLL_CLK_INPUT   : out    vl_logic;
        DLL_FREEZE      : out    vl_logic;
        DQS_RST         : out    vl_logic_vector(4 downto 0);
        DQS_RST_TRAINING_N: out    vl_logic_vector(4 downto 0);
        DQS_CLK_REGIONAL: out    vl_logic_vector(4 downto 0);
        DQS_GATEI       : out    vl_logic_vector(2 downto 0);
        DQS_WL_STEP     : out    vl_logic_vector(23 downto 0);
        DQS_WL_CTRL     : out    vl_logic_vector(8 downto 0);
        DQS_DQS_GATE_CTRL: out    vl_logic_vector(11 downto 0);
        DQS_DQS_GATE_CTRL_TF2: out    vl_logic_vector(3 downto 0);
        DQS_READ_CLK_CTRL: out    vl_logic_vector(8 downto 0);
        DQS_RDEL_CTRL   : out    vl_logic_vector(8 downto 0);
        IOL_TX_DATA_TF8 : out    vl_logic_vector(103 downto 0);
        IOL_TX_DATA_TF4 : out    vl_logic_vector(183 downto 0);
        IOL_TX_DATA_TF7 : out    vl_logic_vector(6 downto 0);
        IOL_IODLY_CTRL  : out    vl_logic_vector(179 downto 0);
        IOL_MIPI_SW_DYN_I: out    vl_logic_vector(59 downto 0);
        IOL_TS_CTRL_TF4 : out    vl_logic_vector(51 downto 0);
        IOL_TS_CTRL_TF2 : out    vl_logic_vector(91 downto 0);
        IOL_TS_CTRL_TF3 : out    vl_logic_vector(2 downto 0);
        MEM_RST_EN      : out    vl_logic;
        SRB_RST_DLL     : in     vl_logic;
        DLL_UPDATE_N    : in     vl_logic;
        SRB_DLL_FREEZE  : in     vl_logic;
        SRB_IOL_RST     : in     vl_logic;
        SRB_DQS_RST     : in     vl_logic;
        SRB_DQS_RST_TRAINING: in     vl_logic;
        DDRPHY_CA_EN    : out    vl_logic_vector(55 downto 0);
        DDRPHY_ADDR     : out    vl_logic_vector(63 downto 0);
        DDRPHY_BA       : out    vl_logic_vector(11 downto 0);
        DDRPHY_CK       : out    vl_logic_vector(3 downto 0);
        DDRPHY_CKE      : out    vl_logic_vector(3 downto 0);
        DDRPHY_CS_N     : out    vl_logic_vector(3 downto 0);
        DDRPHY_RAS_N    : out    vl_logic_vector(3 downto 0);
        DDRPHY_CAS_N    : out    vl_logic_vector(3 downto 0);
        DDRPHY_WE_N     : out    vl_logic_vector(3 downto 0);
        DDRPHY_ODT      : out    vl_logic_vector(3 downto 0);
        DDRPHY_MEM_RST  : out    vl_logic;
        DFI_RDDATA      : out    vl_logic_vector(63 downto 0);
        DFI_RDDATA_VALID: out    vl_logic_vector(3 downto 0);
        DFI_CTRLUPD_ACK : out    vl_logic;
        DFI_INIT_COMPLETE: out    vl_logic;
        DFI_PHYUPD_REQ  : out    vl_logic;
        DFI_PHYUPD_TYPE : out    vl_logic_vector(1 downto 0);
        DFI_LP_ACK      : out    vl_logic;
        DFI_ERROR       : out    vl_logic;
        DFI_ERROR_INFO  : out    vl_logic_vector(2 downto 0);
        DFI_ADDRESS     : in     vl_logic_vector(31 downto 0);
        DFI_BANK        : in     vl_logic_vector(5 downto 0);
        DFI_CAS_N       : in     vl_logic_vector(1 downto 0);
        DFI_RAS_N       : in     vl_logic_vector(1 downto 0);
        DFI_WE_N        : in     vl_logic_vector(1 downto 0);
        DFI_CKE         : in     vl_logic_vector(1 downto 0);
        DFI_CS          : in     vl_logic_vector(1 downto 0);
        DFI_ODT         : in     vl_logic_vector(1 downto 0);
        DFI_RESET_N     : in     vl_logic_vector(1 downto 0);
        DFI_WRDATA      : in     vl_logic_vector(63 downto 0);
        DFI_WRDATA_MASK : in     vl_logic_vector(7 downto 0);
        DFI_WRDATA_EN   : in     vl_logic_vector(3 downto 0);
        DFI_RDDATA_EN   : in     vl_logic_vector(3 downto 0);
        DFI_CTRLUPD_REQ : in     vl_logic;
        DFI_DRAM_CLK_DISABLE: in     vl_logic;
        DFI_INIT_START  : in     vl_logic;
        DFI_FREQUENCY   : in     vl_logic_vector(4 downto 0);
        DFI_PHYUPD_ACK  : in     vl_logic;
        DFI_LP_REQ      : in     vl_logic;
        DFI_LP_WAKEUP   : in     vl_logic_vector(3 downto 0);
        MODE_SEL_DBG    : in     vl_logic;
        DDRPHY_DBG      : out    vl_logic_vector(143 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of TEST_PATTERN2 : constant is 2;
    attribute mti_svvh_generic_type of TEST_PATTERN3 : constant is 2;
    attribute mti_svvh_generic_type of T200US : constant is 2;
    attribute mti_svvh_generic_type of MR0_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR1_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR2_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR3_DDR3 : constant is 2;
    attribute mti_svvh_generic_type of MR_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of EMR1_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of EMR2_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of EMR3_DDR2 : constant is 2;
    attribute mti_svvh_generic_type of MR_LPDDR : constant is 2;
    attribute mti_svvh_generic_type of EMR_LPDDR : constant is 2;
    attribute mti_svvh_generic_type of TMRD : constant is 2;
    attribute mti_svvh_generic_type of TMOD : constant is 2;
    attribute mti_svvh_generic_type of TZQINIT : constant is 2;
    attribute mti_svvh_generic_type of TXPR : constant is 2;
    attribute mti_svvh_generic_type of TRP : constant is 2;
    attribute mti_svvh_generic_type of TRFC : constant is 2;
    attribute mti_svvh_generic_type of WL_EN : constant is 1;
    attribute mti_svvh_generic_type of DDR_TYPE : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of DQS_GATE_MODE : constant is 2;
    attribute mti_svvh_generic_type of WRDATA_PATH_ADJ : constant is 1;
    attribute mti_svvh_generic_type of CTRL_PATH_ADJ : constant is 1;
    attribute mti_svvh_generic_type of WL_MAX_STEP : constant is 2;
    attribute mti_svvh_generic_type of WL_MAX_CHECK : constant is 2;
    attribute mti_svvh_generic_type of MAN_WRLVL_DQS_L : constant is 1;
    attribute mti_svvh_generic_type of MAN_WRLVL_DQS_H : constant is 1;
    attribute mti_svvh_generic_type of WL_CTRL_L : constant is 2;
    attribute mti_svvh_generic_type of WL_CTRL_H : constant is 2;
    attribute mti_svvh_generic_type of INIT_READ_CLK_CTRL : constant is 2;
    attribute mti_svvh_generic_type of INIT_READ_CLK_CTRL_H : constant is 2;
    attribute mti_svvh_generic_type of INIT_SLIP_STEP : constant is 2;
    attribute mti_svvh_generic_type of INIT_SLIP_STEP_H : constant is 2;
    attribute mti_svvh_generic_type of FORCE_READ_CLK_CTRL_L : constant is 1;
    attribute mti_svvh_generic_type of FORCE_READ_CLK_CTRL_H : constant is 1;
    attribute mti_svvh_generic_type of STOP_WITH_ERROR : constant is 1;
    attribute mti_svvh_generic_type of DQGT_DEBUG : constant is 1;
    attribute mti_svvh_generic_type of WRITE_DEBUG : constant is 1;
    attribute mti_svvh_generic_type of RDEL_ADJ_MAX_RANG : constant is 2;
    attribute mti_svvh_generic_type of MIN_DQSI_WIN : constant is 2;
    attribute mti_svvh_generic_type of INIT_SAMP_POSITION : constant is 2;
    attribute mti_svvh_generic_type of INIT_SAMP_POSITION_H : constant is 2;
    attribute mti_svvh_generic_type of FORCE_SAMP_POSITION_L : constant is 1;
    attribute mti_svvh_generic_type of FORCE_SAMP_POSITION_H : constant is 1;
    attribute mti_svvh_generic_type of RDEL_RD_CNT : constant is 2;
    attribute mti_svvh_generic_type of T400NS : constant is 2;
    attribute mti_svvh_generic_type of T_LPDDR : constant is 2;
    attribute mti_svvh_generic_type of REF_CNT : constant is 2;
    attribute mti_svvh_generic_type of APB_VLD : constant is 1;
    attribute mti_svvh_generic_type of TEST_PATTERN1 : constant is 2;
    attribute mti_svvh_generic_type of TRAIN_RST_TYPE : constant is 1;
    attribute mti_svvh_generic_type of TXS : constant is 2;
    attribute mti_svvh_generic_type of WL_SETTING : constant is 1;
    attribute mti_svvh_generic_type of WCLK_DEL_SEL : constant is 1;
    attribute mti_svvh_generic_type of INIT_WRLVL_STEP_L : constant is 2;
    attribute mti_svvh_generic_type of INIT_WRLVL_STEP_H : constant is 2;
end V_DDRPHY;
