`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vaoc8yU2wnOespApi1SyELT8WCWMc+I8JRea0TvMT1kJl8ytuY70lgyu2X/58E5J
TPrnJWvABFAzZPu/M4s8r8tFS4kYYNrsD9F11DYa1Hf0OFZ+kSqAAxI7XGqRCm3R
2+KWKvrI68DIIEsE0uMLOzj/bL5l4WTzQMeaKrPfNL3SHEKr9iOirZJ7qqY6Zin1
jRe6oGzgBgBfPihl5a0ISUUdNtmgG4shmWrPlkFYK6y9fdOLLRv455UPGij4KtAA
Bb5z3nOtIpyOn52IAqOoEsSRl2pXhl2+lg0ISvXh5bGM4AWayf1GMw7zSERlFZJp
3FbQxXK5qAUC4Ese3s+l3JKc8LVn+5vNMYFfyhD40sbz1ttWTLp+DOuhayVebbKy
92JDO3DuHD/FJeWKznI6rIwX7W7ZRtAL7eLDzkO+RfQs1ofqAfQ+So6G9TGQAmi/
klGQamqUdU3wjJWU9ksSBoRxU8XZYI7Tt6enh/macmsWoXaq1o+6JBD/7REik2KV
cJtnDJR2efEccWTyDrm/g0uAJAARJPrIHBOkYWu0Mhk6rDLJXQtihQ4VSN2tML3N
Cp+OpcHYRzR7EpvOo6PUGYG68Gv8WgN1xUOe3NpWmOuBTochHRNVKada2aCHXWd+
thAeWALpBZx68xcyniJtcGsfu+gDLkgBi2H+cE+lZprnMBjReyzs/sh6fJvjDI9w
sV49DuAd8MqNkTPfoCfUtrZt+zuEUpgHIvP/tCrF62jJW0VHDK0LAvoopor55HTp
MgRihxY0PMhdnqNp+h6+l9jSnlUrQ/hqaHI0FO+35vVtA05JLPui8QXj3BMUYNma
`protect END_PROTECTED
