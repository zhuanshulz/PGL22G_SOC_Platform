`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WAzlmn0LdDT6mfg2Q+Cfckzy5YuX88hBqxUwyE6VoWsvWn6EthAq3q3RdjnxFuzt
wZeMmIzio7cExTurLw1KvMoq+PyXQLzwfZvYkkNF7gLciABlWrotyq8WUh4pLZ6k
X9FeOZ2lSorUO4nhqphd56KdoslXAF4tHiNcwrDieMXfGJ1/265AV9tTvrgur5xR
FLHnb+dlw6VTgNmcTL6w66NM6B1ZyX35dkEPpDCTyTi6Fd58jpG513INvU3vYGrz
wyfFG1Um8Xw0HoyRkgCHNgGHLuZ4tCmJOjpPXud0D+skdShHd1OPa0KxvzfConw1
fQipdVYvGByu7lC2uMoOhrm9TI87ghOT9rRosowGNBs5kQ1HqveX0nkCg0//NhBX
0N089Jh+dVfn+0iMrDKpYaFcYVZI9b/iq736qQdOqfM23QOeJneQ+CbSp7L4iXP7
e5utMOlzOF52bxDxV854T0MSpxfn9juZ5W/Pmb1wsvPE3sk0sinSnhNyZ8jpwhZP
r/NEQoGc74lqjfnQRwwwx27pdPDsltCoJlWadSqzWX3QT9GxSFQeIdkryO+yu3F5
bu4tQorlZu+xh3YTxOfoEKJEy5TwGYNoUyikP7x04OVpbwbdvGiDb+bFmT6Ih9Vb
eRjzZKYOr/zKMJcABgLYBd5vY8H8VhKO2Zt+KhxAHI9DL/87Pg7Ef1soRgwro7WX
l8J9KFKrslghpZfhCq6LV+vQjADyVbjJEmsTtKY5zAh36wXGmLfVX6+pQXqx38oW
ndEEHmUxenENszNo3P5RTdiNh3gy9ZDErEWuTwEjC9akrgT+KdAtQ+9+KfDiYWZH
bjYSE8aTWWCSw1+WOgCWXT/fM+T3MnpZwmRvHYrylHXV2KMQDxkp9uZ5+83NMWE5
XaGY7ixEF4HdqAQ9K+v5JYAKQMlTfUysTvL7ahZBlgo/eu9tDOAdzfaTenaI/UGo
VBef/dAr8HwGwBqgIo69Cm400sXxu8ccRWUbaK0Esyz/TdRjKYV/emEH08px7/gU
qrepXNd7lb69FpARXVh8D5v2ccvJaZWckxgedI9w4rTpmh1q/VO1LukzXg60gpni
ROnyDnJjMX62dn7bMzvFatrKJdtp7Q04yXyYwtWjXv6vnaZzfzUx07DWi79/j0aU
6RklHCPToWqMrRVQ1N1V1SAJMu+Eq2YiD53YOl1LYy5DlEgC8Dh7PWav0q9EUX+S
NM6B/nv2wZSfzXA5NkZDwCTHEeNjQ4BJa4Mx8JHX2S66q5niOZX25StF6Kz2u0Ap
PU3MVjpPSG71LU2lqX1uKL8OwBH8Tvyz1PbJC+5dqd3hom7p+pJd+Tsp45n543NZ
rdsYPEG+kaY3uLGhuIcWNWkWH1t01BDNJ+3tKUWOYEzFW8LBVYY5UCjm8IOi4U1f
f8t3e8ALXSNSVpkQ3fvXPzgQ2ax39+COrBwHehLCrDBDnFaFXaXJkljPnxjLr5pP
EmGPTxIh+RXa6ifSce3gNgrnjeCDNWtlGUD9BhPhTATssUOvXfEk5LAXhoBFzo4K
lPyvglTdGC1JujorKDFHodvRqZ6xam7lEKaOeFwrrtQOH8iC+VgwksCi5V6/kubN
NHKtp0Z9o5lHBCn0nrtDycaSO8o0b9U+yPTF/pFZWPqFQiFPgvIHEZfdAr/IEeaA
aRkvWvNjm5LDHuVnN7JUhKTxANAsvkDjjWzU0ykO2hYkyGCh5mYcKQJ5hokSGweV
YCtu5BDnfe59ivc2UbIX1WnmYqr7H109UkMCZN2QJPsMY7D5x8uQoWAZuvsVAbc0
IwESIUbnkaMvOl5UdbFqOtD9y59IL0w74KFh9sngd44YLkI7FooJ9w0BQQMbdtf5
cLeleGOHq8iZqxAE6d/jM2NO3qSTZOF/XEbcKgXnNsByBpWet1w9mRjc0qBXFZGY
FzNQbJm4tV2/FJFI/Z0BDKw5pFrwNYAIGCAFqqezcRGsWJxXp/O2/5RP/1rWDwgf
hWWWiKIBtf/l7xWxmHGPTjrxPhQMYiPW3Lgf4cZCp1iDMGyo5PslbNBV6NfTUE7a
8/mY0jA1KUEi1UQGinScEfhHxRUo5LRON3v0RHiiEMHhA5rCPbyJdLpwcHgnosge
dXQcKzSZ8F44eskXQVSUOVQc0T5j90hALIGFSmI3sF6x3ASpHAWMNrfzIFaD8QFC
XferYbP/q6w0iVnREDnQ3RAaJgsOnc0gtvP2w4HESODJVgY5GSO1HRDjG3j0kfUB
5ziigGtK1etMai1UigG2YxdXkLSHIaITzV4Mhg2HXbVn/eG1caxd5EdUOlDLmcvX
xxMOmvdWdjOIQ90gD+nWrRNdfXSG+m1sb4jXMG/XmKLno1sBphlc8ztwLx0N9Y6z
aKPi4inCT9kwGjSuz/MykvmOy+J1URzptoXs+l255nvM9/2/x9ENU03eCmH113je
veZ3MlwdWQI0B8k6UgvUYgxwOMY6GjtOOTOvVDYBnD0qO8HZWuOt7CzaDWpQoXTz
7Z2u9TdZRFxEkbEOiu28v3hWPyj6GPKzad404SG2oXwTTXT3gPKQUH6HnbR3JKLa
VlabD6omqnln/c3sQM5yATICKlShoC11eCR/Vu5dIrrxD8ZnM61b7ho0Cfz7IgEY
+v+ZxnngUHSefjyCPcncBeDsiMroMP+ATEfGKDzyL6XzyGH038COaENR310liiOA
s4OV4+jwNFHUTkgrYacVacK390kX6PuTDFRIIfBsxXcux/uXXAiAE8SD0/SBchW2
Ky/hTMIp8mq536exa0nHI2zJ+R6zcZqkbVRsYKOmaNwSwA5ZQlhZ3oU7CXn8Ibi0
ho26jHmvOqWEgWsUVqgEwHXGaJTgWFbBr5nPLgfUPj4sfD+LapP7SQqsrr+d6uYd
sVLXRavIj3OSOmFtDbfOSUH76vk3g/GXxI/Q3/emM/MXqCrPdtM0WP0qb3nLWxtB
2XxaqDQOT2USo0HQzdmHOwXIE9H6O022jvcssuOMrOqsO3AISWBVb2pvVVBJD9ZO
iHw9OPXs98pH/S70TSfLt+sQBtriqahN1XtWjXfz+fHOsieWbOwF3j1qrzdR+XMH
E9qZjKypthDzYil/gu4HtjBWLD32q3+K5M9dNS4lZZxX0h2Eg7vhLbP9GsTQiF+m
Vflw+aZBviggNZIkWeC26GMsAVqv/3t4t5zjAHi+XSjSDh6Z7H2SlhkSX9WGUbUi
hV3HkTTzFdo499OKdJsIrn3oMcu06xY+Lyy2UYrFe+UdlLmC0Uo7WnPJJSUWgVyu
OY9pOKRbmjyhCCForuBaqcVaxw+er7yP99qyGfJslPcPp/tYFxC4S7HsX90wQFh5
a3lHGnL0nuTD3k82qVOCmk7dsyMGtDOqPmgKePLEOQyP0kCKWEVoeWOfex+OM/JP
iSEovaY696838KHd+FH4sYabL8Ztr8TWllTPKRnfDjvBn3s8vCTRHPMf5vJP0rRa
w5sxjUwTCgyxQN7zZr1fa341H/ZjU/WLgGu5H/hxySyX5jZuDfNSWwQfXAv8/HdW
3+b6w3EpRj9jeI1jDVYtyhCbG90ofzSlzuP5YMIuyXRp3mbNtR2fLDOOV0ou05iw
j3dMN3gPbwzTE9NoekE47CaTjObLMw6guPJg7yAVuJd0vnf8alUBUOCx3pw1so2c
IQtir8cUgttbzcqC/yrRVM0D5MWQDJzZkiCDdVXtWOTjfWLeL+03YhkS/AVb2u4i
qyOhxWCNuQyjn8Lc0bJRzS8rttpSBpwPHBu84+5ixOKafYxaM3tO3mZ5I0KC2IcH
sn/6H8XqDsL0IuuuX1x5TH7/sZ54lwo2xXHvG5Pf0ssFscUDsMQL/uRpMmti5hAY
4ppxiEdTHFcAfA4VIxx8WTiw3/JdIWB+PixyP4Q2Se19UdvQXwbNAs8C2v8Bbww/
Z2Hkdt19TPYg4Op1lSk6AE6zoEsJFj8D96CzEGxEIPpxrj03D7mC0S1MXttM7BtE
pdRmmm39dAHUuBCydhkATLTyk8WMkbFVnVK0Jv27hCHRAj1QEcpuR575RwwjtdDr
QZAXr92iyIh5Dida/4JnvP8OgKk4MMZeRXwkqjHdBK3WFb9QYpNseuZ/zPiiy5VP
QMoj5OVRhiwue/aLF6jtdpuF3yGWJHypmzyfMDQkS9JqS6o6HSaaSc55ZmmDFaaV
V2Td+p9EOZktzFyBiOOC1/MozvAWpJwPlnEjzDfghp3pX9FBUrmvQubpnEPZkd3G
7q22bddkCe3JtTpfAw8oe4/AVBbmVvwZZ+Uw6/UkvrF+s84kBbspXp+cLgxqSYRe
Nknje9hmbB/G/MKrdLWrW8lNiJZubwtPQkIR7oPV4kkMGpfeLcbt7l2+z2iMYVOd
6XhCYduQg2mabTAluIIVdoU+DCrKbOfZHW1rK7KfWxQmIfVUzvf5n53vTz5vbO5j
8q4gM1fn5HoSte+mCdx7Q3q9kV9/Y5LjyzCwm/jl5FdvwdsQC3xqQhrVgmv9lt12
SUr6VoWZd+Pk9X6V+dm5ibXJ4zXQC/dK7HDuo6vyVCIh73Zs9xd3yYiaYKxztGqY
ZvHpiqw7vyiIBlU8vlH+D/WNcQUH1OeMM2wip7bZroA4cjsd50buL/r2/1BEqkSR
FMCSvjGKtM2B4KlzDVgQqNx1HQD+/bP5Jf2c4/lWZ0WTvSbt12Ieb2KMYZfVpJAg
svbd89vmM85Ceukoj/RigTPtkVltHnfUdzDbnkVu6TJsq0+ahJpI2tZT6IgmbuL0
tzskKveOmRaOJJ2R8MQRNc8v0i9Iik6TXIn0C9V/0GJPrAAFMcX1K44GN9J6zIgO
UXgnG+Gzmeji4Grbd3CiIfP48gvfKeSnBMtLXyaGfmqrpZaxDE9YIV9nVZshcJE8
X1gNYoNbVb/4uqINRG2N5rasm2sbzSN7yhwRqsX4MzHVhqik2hMpFeb21fkah5Bm
/nXR8+TDWWrR9XkvMySgUAPLmbu8NjnVcAU3bJ4o4ZYqz+9xMDt9orECMWoXZ5Jd
zqH+xLbrchA9SG9Zc1FZpp/sr+ADwCl+qPW2E4WiiKFuOIi32GccQPH1QCHkf5Bx
1Ovn3LM2kOrun1X3bVFOeKQ0blAvUoRmMODqzhUsqMRveBh1ggQbqd6rSFqCOpBM
oU/S0hCZB13D4EyONxSTI++u36NPEwIGbpAle6WpNSKw9VfnTBQ1xz3VOUKt/saT
RehgQwbagXK3j5Uk77vmxEXHspOOMyxvdYE9jX4cFZ5fj6+l57BSHm2c0Y2DpC8q
6zph7id14nvCc6+d50PkVhfci8cxIujRi8pwt8ZR1lZGVrwSstqjeTmn4MzPyZf4
tm5tRjWVbBDryKRrPIxMPlIeJ5Y04oGwCDhnUdWjTf/6aIFu7C3c9YjtdHH3Q0di
YiGmImM3eTURRuyPI9vqfY7zUG+XkbKp5mY2b6SgkwDMyJtKg3E2QlY7gp5JkXPc
BchqYXxml6LUdpAP5gq4CHjsvoMcA0wJ3SsXS/EXeGWBEZrc4orllwn1dwUNYep7
4FKUoBMyUCJdO38GVCEJhv9v7DBfGHz+qsyilOZkQ7+6G5g7KJqhxLL011z5D13N
O6wMlIGR8bseg2+mWw7XgkZsCzRCVq7AhnuqjGFiVz6R9YDo+sHtH/nWFQYNkZey
pNr1ShinjmaJwbV99Yb1GbWTLL7y2PGyaE7t892k0NapPj9ozh1QB12iY0gsSH/t
6EMTFleHATTQHKNLUHx/vep3YYxnDQ25WXlfoKA49wTfbp74JLnM0lAZYaGj+yPp
Fb6wD3CsDO2jIktzd5i+9JtcaLAHoWw/y46eCLL0zUZHFiVS6n9+1OvDfCgJmpYd
J93As0L8Yyf4KsGiY4YKGoNocb0ejT0v9wL5+NF7zwDyTuW4rLL+RKIR2Qi9bl75
ZEf86CeyjsUuGARDExygN0cg/OD7zWv2id5D+IDM8ZRTqpcjFIs4WZvnqOBXTPUE
cM1oIxF1de2Hzx7LwBnsFHPvLRvhY8BIVEUaUqLzeEigoxUsnBI0UHPABO37nP32
vpVMHHtu/1q8dIWfpjYiralVpEYsxcnEXD7rW0h49SKq1aB1bqgZSJvAKk+xEFBk
JzmAmVGNtCXDv71K+usqowt2PSjYdgPOHjghHbYUZ99kb9qK20GwUR+t1pdIZFJu
UYgoTLSzXF4LxkzfIntGhu5XZsx5SjUp6yg4thFwcKlo3IgSkeTNyGpZuGP1Xj7W
rNRtozMpTqN4zUF0+zDaz8skfrwzpgydZM5osEI/Ozuy7kQzJAUKEyR/WoOGioQe
DNfj5/QhkIuxm0y17aFuKES4WTM9PW7xfouiYG56CJScdfv7BBU2V4WrrUY51zvb
h2DnHg60K1z30vzWaeZTTFB4XXq7cKzoiTFCaTgNx4w9UhO/lo8PaORPtE6ll+bM
EKzNdYJpusP/t3GrtFx1TKY7E5YhBTDZxPiFUl1LgOdcF7naYd/uAmN8HYh53Lfy
TZTU3KF0K+g4H+qJ0ekG9sk2QTME6ftL31HaH3QYVuN2Ew28brtUIFLYgbf8CwW5
VnkVytcdBOZJYLLU4V7TL35dLhgKPTliZn+zrrGiuw5wdBovAtBc5IDnCPvOtuRU
mPpQLVTmAfqVFlIFYvLDOuERfEJwWM3KKHB7WS2o5c3wxuWg1bVAv6R6YrJXvL+5
IKJHzs1YfuJI63W2G5erUA9jM6zMmKdSYrOnuTuR0sV6s0qzUtAHo+wjTarp2xUc
iteb2JfmlOm/Up3C/lgRvgASiPmtUf9GvjoSuU6bfLFaFohLPZ5wJZID+L6WhifW
41DLUXQBBKvMT1og481aZ1dySneUDiiKnhcrMO2cb+y3VcFQPJaX5+tnd4XuQFp+
5ZDcfPaSx1suae1BV+sQsWkOFDMODDY0KHX9mtfmFcbzM4cbL69DsWDZo/jlRumG
HNKn5NtUtEtWifZgijcL+h3uUiDiMckNeaLIZXvMNNEkbL99SBhIU46pqT/GMX5x
iRDVPcogrxOxWTptm1eqUTjxcMEkz4n3z9/sW+oFsWysh9qdW7MIqaaaKTWzFqx/
dzQJshbCR9lHoWaqaWVHPMlrzRebCL40cIdHHhILAoZ/w7z1BzKkvsJryhD94B45
clrfQf2Nw0BRrl5Hd/QrIOUyIhnhY+qjyxFbkINtnjAhWEhDN6vNTToTgBxV/i/3
`protect END_PROTECTED
