`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5h9Dt0bfOhHMzyC3tzv+sNAUmBwbvXDHJdvmUJ6suDv2erMbJdXS9IX8oBX+/vXa
82m49Iqg+h2rkgaqc9xBiP9i2trG96iorduEEH8Laa6Kh0gdKDFlY0a81R2/Ly0t
luTZ26D5LhVpDz7EPQBO52nLpmGM1tHTsduNq03/9tQPFjpHWJvjuATwCYphne5+
AMjPGEfkJ1VzV2tyVI5FOsXo31c7Tr16NBC7ypmc8rgTBRZrajdXov+elWBdMHNl
3dXV7hRxus0YXO/GqXZ/HqbfkEASLdr30MKUccgoMLAqOrL0WvViM3WawlSJ5v07
QuFopG0j0w7paa9d3D23wixhN9SW0TT8ejQe6b4Kj1TAHo9mrxkggL00r1E+qNAR
5+Zb94F/r18pGBI3SeuZlYhJVDyTS/JzA+1Sm+EB9dlDdkJ8MbyLRjguTA/olxyB
03LJP+pqx/d7vXmXQ/vIwMKjnn5W0T0Gf57IWDOX2EtUBCwQ8tyUIEhdT3S9QeD0
44B560KdlpGvFVU8Y1AGLlM3Jijs3ZOUv/SALIvlSh68G30pDeHTsaDSbNlqZ+3n
G8j0phTp70hOl3xtQ33kT83w6IkRg4aSowa1JCSu+jYFt7R3SlS3kTRTMC5D5Ust
bdlfIE0IpnGlfBUlkX0wKyZDYAw2faW0S7Sfl8B8T98CsP9rzgO3kK7eUsPRHiiR
l8HzFqNaTuo08T3+SsE9QOSqkzfH4CjM4LOTdn8d7VNnellPgeaACqk4TvkPuavs
8a8f0lyGpa5a5xHZ/uTyq4KcsCXcPeNgTWwDmI2X9l2r78ofhvjADhXuk4CPpANb
4iX+3cqiqlmBITSQqaFn0ozbR2e5SLaT1A9FP3/Mmlss4qyY9s6r6y4kkofCC56p
Hup5kxJ4qzVpLN6RtCsDaKnJx9L0RtC4YVzUv9CDheRFQ7NpUgvh6wREX9LQS5cj
3LeuDqs4Gkd/r0sOigzfhDiv/jWKFSNPViAK2oFgNeuKxO3V0fxyZ7s+MkyGh6MS
Eli6FoQxYHzOVcukH4zWHQRvEhwjNM3UbjkDC4xoGXGjhjOb7Udg1WJB1ZYb1qZx
YpGmmTiozhQohsuC9XiR3fBOiVZiseTrNjP0fT0+Mkt/M/8LxhA0czM1hRDl51QK
UwQuDtJjjX+WivNA47IPEIWtcX6FZz319gsFAhlABItkxTNyfVhV5jiR7foIkog1
rmaQELzB+FuZv5vZL/dGjgSoLgIbrbkCpGltmhmqxo4RF2MGgd5/Z5mKPoupltzG
OYaJrVxryeiZ8EQsLNsEZkSxbJx3+KMR32yADIsCE/BpeKQmLdGsqJRq97BmzE+c
TbBDBOdn3/gKrDfC5jLSzjOf0ZAhBx2V3ix8pA2YV5BzVF5mZ3c4SISKFSL1OO4p
r49n6RAnKncGIrk4LeS6m86Oyu5tUoXv8dkUSEL4xNLOVEdHHjKGgtQoM8ie6B+y
TwGm1DX0AMxgJZ6jPnEgY2iulUa3VvL9+soSV/BWEDGkd6qvkariY5EuJbMj7TSz
pfXG0/cQsMyx3JBqTGYb1uUqyFC9NqNmgbAKR3aWil7wG6+rfoVudMWn3BkJ7+O3
+l7ojSC0cim+Lcawdzn7DGPvjn5J02UZan18/351aE1Sj+w+LojUWiEXLlZ24Z/M
GjQfDfjq8C7gr3Drz+wiET6FQ9bfsuhNHsqeXH327z+WWOLlgfopzIUzbLG2UNOg
nD1fQgMG0Z+VlhaRqRz5iujo+rbHrs95JN9EWbM3VtFLwkzw9mnY4zRqpqGC0Zfv
RJh0DroHzOz86MrG8ye84vgbvJTJqJ4s509e7LcEE8h/Wf9Hwlx9tGjRdXkgZIVq
Ad2QELDB8T3EtzDOKL4y5cAUUtA1vn1na8b2hn+BhI0eVWVMON40oNBMjcTWGn3D
CHvg1kXl/xL3tbiEkhfPI2sWar9Gfu6oRPmtTUCoS/SyZSoCdOwRsfGkd5Ht6hk9
Bvtqh/gSH8BIfUwuqtsNLllQkEd/DHt0qe7dAa7ZjtuY4titu1HdzMycYwZzkCba
kGWTrDn7WXhv7ZJE1Hqxo9CwxX8cM94W7ubvRINZ8pJ+zfk+eqUKdj5kRI03Va6K
F4KCjWxOLBahNYJAiQJMqGo9CTY2KXa/ooQpDGgQZxKCw2JLjEM+zJu0pc1vVVey
seOz79ZFNgU1NgibtQ0FPD7m4bFvyNdK9l8+fw94nxMxGBdomU/bOI5XGCO9EkSi
YQxm5Ml1wWcsvInNwKNYbeNJpd6SS+bwnBtekmgAhSjGy5L++2401E7JsGy00QHV
jRf07ggdwka5pLwtfHJrdzROKmUPDZioFQGyPOBlZyu3iBoDSZzlSSUPtMcWTnmc
DdkXgBi1ZVvE4+WFEc3ZFXaCyz+cXLjW8+Rfoj9ihzN4XajKdwhincNMShjQQQKu
YtxR8K+mu+h55viCOu9j0SXFkK+Dv/QHmOOyvudoqfdaQHvb/9JgFqHjoXHy3QiA
vqS5zYO/O9i71Bb7+QYOhn6t1qkgTdJIhYLJYWt552QNwV5iYhf9cCrqL4VvRcmZ
XL5mtlwdM+OIo9pQ0AkunFrCBaZz0ZG/BX00sbb+snOOfAVHHgVF5sXkDO4jM7oT
gLaSvVfBLmb6liMk5YtdCqq7EF8UZlW00oD8RREv6fhganqIha+r/sJjmWKClbxa
6gKoI8XR+dC1sJV1Lda8Q/I8hR/3RbaKIZrcoeEP+gdVYcGxpJZJvAIWE5dyf9t/
nMyj7NTNprxV7W4xP44OKsgnCr0BzOBhOBZB0VonWA7Net8kOxSNyY3Kc/Oo+KkN
ARU3h94PUyUJh+BKa/LOXGAO5sx5FFGdXdLblg/26P+h4b6P7ABofhMjKRhI50fA
GN2k0cgeT0G115fwElLYR1mUK/+6Xd6SFuR0EBErYy0q54P8QpcbuHZpFJgZFZd7
RxA03EjNbejW9RA6IX1Hxl2Fu71QWQbPyfXZxrvfGnToTCVVDWj3ihojO3bfU3pC
j+1iwagIDgb3Vw5zvRrTQQkZdn+NezjMVEv/hL53xA2AU5WHaFFdx8q0/wVurB8B
O0yUrDVPSEoVqPELbmQLwfmYnZmLQEUZHk/rP3oHorTGvs8SKU8kgMZsEffpahwv
wxKXWzvYeCMYqiqq7kIBJESd5b9dGqw02rDG/vfDXtcx4hv1ymBblf6bVB3LSHpP
7VkBuqA0M+xaSLel/v8VMuJGR0ZnkC0wo6HicsNAGG0hU2jTVwvBwX41xxdggV9G
rXS8VzKA1D+7GXINT1+Stt8H5G2FHbT9QPDIzl2IIVPcBJLrkejNSvzfPIyP3C2i
fFmKO9kv8Ig1JHUsWUMQelMcO0fYJCczhIAk8nfu33y1dpYfL0rjvfe0j1Kxzaz3
VMefG18XUimMCGo0hTxBm6VvoVj59jhHSqomyegj44j6M4qSlG3w5VKdbvoLSkY0
wBZn2fDkaMssg/506XVbHUnAlaJLJBBn/k77jiXTwRaoAshXbzy5v+9V3XEdLJXz
MX8SoqbpdGoffUdo6Suq3ozz7J/yQuBU15P5c84hya+2ws0xplhJ7+ocjcyPEJFx
COZWup3Um327jvamnmwwnQPxC8GU/0moCAGxBdqyd9/bGssDhc+lVKOrHEXQS0ph
93GpDFneMWcy0M7Q1mHsIwrdhwUhWRMzxzAg16lQ5ThHGA27OSXh83V7h1K3YXLn
t+m8obIQA9jYZt1sBQRZMTooPd/YhXhiA4/L7fWZoIHCMm8KGrNJwkukTRJimbDV
Pslcf778CAsEtc/Eqrw6FFEahuVo+YPupqusJZ4J7bgc76S0RiRCHsJVjCCCldax
gJBn25zQlnrADSvclTSPLMfXx37E4JXciDAzeZh3yDKJSAuTMdiHbIsNNAvuD1Y/
A+zWKjtHE78+lnnY2OlWQi+bpJVig2J+LSNgfeYdyeC5Y9+5sVnlR7YtrEcuwKjK
J8rvkajGfu2CCZUyR4x9TiFw/iDIfZtCXVTHoejg0N0jE0BNeRhXpRF8C0sDqVFR
VZBOBYlGrmlHR+Q1PZnFeP4bQzxaHFubNB4jzL5tYtejlIV1ctfBZPFlfUwUcOVP
U4hTTxVn2hQ1aRdvwsaUCuGC9AvCEUzxTokBN9o99Iu+ZRcjmUfSUCUNmcfxbmwq
rmXVHV31LFfeuBohIe0TBLlRLCB0N416+QQ8KQjryub13+DyfLNUsF0ohZXV/ViJ
Yu6y8C3v59uM0Kk+h+smjQf2rDeV/DnxalEfGD3kkURk5307CGhGuL+bgw5mRus9
Q2+VPUrTK9V094VGsjl9STywaGYupC2aI7hha/2hOKDKUSv0hMcex3B25Hu6uUcD
1s2UXHRZTL2KWcbl5ycCyYokckbnk6I5DpFw9BbkakvWU4D3T0QjTUL6SCfrA0+K
nmY3pJYTRTNtAIcQZnVXPzhq2/GLUeCc7/bcfY8s9nhr4cpAbI6J+55FZxOcOkEw
kzbwXEN9T4ysS7QftgjzftgNT4awBn94WLFeGDYTlzSk/l4rY5Pur8tdL4PmW7i9
EgRGh+9FPRsLtVDjikGgtoxXZYHvCRoClErUMcyU1hay3JsfKH3hXN/tDisVxLZv
3sftiY/0JdEG9JoE1vWU2KHd2TrT9V7zInZVLHIusziSMKG5dQqePPVLb3Lfg4PQ
mfq+YAGmxiMH6JLUeMDJfEgelDSpaaRF+qW0U/3eoCcstVzvw2+U8JIenz0DcbDT
nT9VLdwq3EEoefJ20knL0AWqJuZMXoBCLHvh2QbBtG/S72O4c9V/GNUc3bI4R6MN
AswF33R+jkE9HWD6vud18i5qAriRxa0OudRL7EUvH1j+SqBez6NyUcY8Mrgvb79j
DqkhyaaFdcvW4ofvb76EggOWLrRYeufnCCttBi7Ugbk9iqwrI4Rzc67NVH53OZI5
OLfabvuwwTqtO+jNe5zdFkjpUmy4aQ4W5cIsXWSKQpAh7nzWi4GsCl6R0ErTRZLs
`protect END_PROTECTED
