`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
txPvH5Oe+LYqYfSMiwmPvX9ViJ/b3wUaZ/A6LV95BMp6ZWs9v3z/OUm4QN7hzGtR
H5m93DkKtFvnyAZeUbM5rnW+BhSCoZqf7emOHTgfwBjhV0EgOm4tY/YPqChcN/IN
mVLVXDkzQNgwuwrLok8e1dKeC3cPOH8pMrB2EcRzEB0ZZjSERMm5CuXjk6imQ/xD
KdY+h/ReLlUfwJQMvFyuRG/vJJqksVBzY6ZTuphZGV7ho16fJlOBGOg1qqrt8n9N
g3hSssHGxhvYQYlTSOSb4zhq4inL2y8XV4CKbG/Zt90/7ULpLIxQy7vnXVyqFqr8
NQokYtU/LWvKHiKMcSklYQ+mM0ajyAo9PZAJzEsdqXE40arfjDUauWWAKcf0hBry
dPBjpeV74qr9/QSwPUhDtHqiw7Ff7vm0ATLBrKeWwjY=
`protect END_PROTECTED
