`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pgTD9xx6bfrQmCuDgxc3T6WMXYS2W6bVgO17I4KlchZcdOHsaocz5ug/rqyHPQGZ
iYRQewIHu+cFebPzygumt+AKQokBi6S2n9/I1m7bL86JmhwKFzkVzouCwQcUxJ1k
RKDpxQ6LS2TQxeX2UOOVf0Jn7Vb5X93y0MY9zOBnzEU/9S96Ylaoh7XMHRK19ryq
Qx/ZJlHpJYBg2B6SWfHzJibA5fIAZbqh7TriNjqnv5k=
`protect END_PROTECTED
