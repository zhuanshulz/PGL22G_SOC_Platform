`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bsyZw/3sD5tcQAram43c853ZAvAmkn1OAt3cXO1LMyBNwb16Q1up2NeYQ+BxsY4J
aJyr/hrNPXrcr1VXGrGUy7pmYFxtSi4cEZu5rivKoq6mXPGsWz09+toFsVkD/ogn
M7nn9DqVSpaGp6QkY1JW58W24BUDZiKJcsFvLk/v0oFwO3Fx4LQSHX3FyznyRIQ+
G6Xj3fsbjMCfpK4fPAf1dV1tO7RmWgxLfaajaxHe5lOaC1TLALLEbShTPEhRQQFN
BEwRfuLVgWtlEQVch8LUuyaPykv9KU2t7h4Z1ftpQp7GBlBlaUuE6y7x/maxQWn7
yf2FdsC1JeM7StpbmqH9G8QsjuQwbaYN/KhDedoHBkQf7VpoT6JG6PTmVsw48cL5
PNg9npVKU+81iJCdKKPabPDFyV+ci66W+MfOvfmiVx4acsOx9F0s8TKSZ8sNq49p
jITs7s14DGAV/DAflOVOAZiCupYcaftv42RHFTSd480cqGhLKrKm33dStDJyhaUq
5qqTAOkFLvzSoEP8x2r7Hj1yqF7strjmuaecHSkufIqkRqisQMn3gamCEI2ovPz+
lP92YzcWTGn7+xyl7Q9IQ0Yhx4lnQ4zXajetSBIZwZDVJPMnGtuxE6DNBf6ovFKs
c3JGfAe2AgO3pKENaDOscBbPKXibWEBWh9qss/roU97bNTo22ydGVNRM40mD9ElE
jLUF+mB129TkwBoQIKvu2STSH83TPK/tVDXk8NaAGqGRnAVbP63dRjwZMyeLYqdr
5CFIlrJdZ5D2VldgMODKUy1Pe3+UZIJxdV/K6nG7/ChsB/Ub04SbHG0T0LlpvkuI
wQ0knDAV0N1s3lmBlqOqbBaazt3qzO33WixhcwIKnBt8qGI6KUr/O50YijweDT0O
+8raXGoZ1jm80P2bHStHeG6Xx3JFL84CGfsQjracdZdYm138kJVTbaA5GSS30HBE
xelAv0rF1JxJE1hHRCX9Cxq3u8/4BWzHtDrUJh9Ev4WDm9aDCUxjfT0vTl/3LKOz
3EczUogQxZ1bLMPBYELIKS2jmKL9Ckx/QvjdTVoiQlsv2CGJj7zx0rIhzTIvhEbu
TgxpIJp2HNOuFQS5qep9UVLkAZCo/TC+aWO6Q61WQlChKzE/8LrUs84ODXXvqEY+
tIFWIT0UHEQIumse6JP4xZBZv5yw4R6CPCvKKj0Q+O9RGfJzZQy+j5d4oM80a7vj
zvLM30aUmBs5CWalcl7vduIbxPwrmM+X1H2s7YavEyEtzKMj2qtY+QoXoT15Zn4e
KB2UCSIlWkS5APdvegbTLBtMFEw9RRFLsPiI10K2uZlpgC4wJu6PzUBMondiGzkB
SuhK7/P1vPdyDYxUNX+Ial9j3Ka/0rZA9mtacaymBxA0LcNrZprdctTYN8mr1ZG+
Tlyy5WOjC5KquNLWSeIhxm+B1F5yzVX0IDx+bCCcmr96Ra31ZIGaF3T9VsCnPjMI
IdKmgiyW5xyFAmRFClLNs8suirID/MzRUj3D8OkwDHfsw4V4nidgnSEaslTC/Cg2
ty7Y7V0QRDDFp/Q94So3foISGeZQRH9wnZmf4XudORQ7AoYunBgisBTGwETkT5XH
jeO5hvqZIajbBUfnsM2oFV2JsIBztDqZz3wEOp4QyS1qcC/HfBwEhsspesTSHseb
P11esOYTJv0jHcl2lKs2FgeI7LNe6Qc+bQ1lpoEkf+hjD7K9XWGdF9IGk37V0vaF
2KrjY4azHfT79ODMByE5+1t3cNfh9bboyMnwvQfl+G0Vve4CT0FrtXuwbWP/lODJ
MMD6vTGODC9ZvuL5LhXbLx35cyjevFEpNm5X9nCZSLQ6ryLyT3AgcYxbN0Ko5jGQ
wTjlU2chfoJq+ZQvc/VrdvaREHAKQ2JrWyt6JNapYlGYCZmQ6Y6XcgQ+ke0vsDGm
bB2zjeiMJmjoXTZKJUpoVZnwr+eljBieTy+FdPKS6pNvNaAd2yOzYiWNz52l+Eo0
lXW46p/RgapgvjWqocEMC+kYtGBaYE0XqSna/KoKqKMQ0EE7CfExQ/CSbznXaTsU
NqutNEqcY7etdjFofM9wyrkYauHfQzPBdeKmLV/zeQ1kpNKMosFQlVhO5ACfLBDm
TpmoBhvTwCKF+hOTtJ4cAsnazjGh6gx+Tx9vF4aoAs+AZelWfVBsVoiTFnSCPWxR
R2bm1ihgQWdqP1HwwX66by4+hp1h0WT9Lv0OMwE5n33xdnEcTadU04FcETTenAMa
MZa9B5Nn0FCXLe3qPk8We2z3G2hR1brfBySzq/AkBx+z5Fc8NHXfD5fz+C+Es8UZ
cbS5telw0N7UZCnY++Q1+qufPvmahuMX8+bKdzAcjxa2QAecHYo3eQaes4+OuMKb
rxhLT5EOl3z7RHbnh4fspcHLkdqI2txk/dEsN5pxarq5TKyodcDopIDuYsr72r7+
UesnfXkol/a29FDeZxnGFaz7H+P3ro63aV8LpgzwZ7y84yhACSW6/Fjr9qt2s9j2
crWcyLo6CC8SyFIyevkUVzDeWv5MJYvOhmrTWdI62Hy9lE+tm58mFIVGs6KXwLNa
IqPrdGGZ3QQni712ouKrzuyMe2NglhuP7XI3yPlRbd/twFFdQCyM2j5YcipLPfcQ
C6hH1Ud6YfUzCsCtSGjbPKg6AMM5/xoS7R1ivTHcWtvRXR7596FrUbYxy/3ICuSf
J45L4tGhnD52vo5Kae2Rh5mvZXDIMX/1OaYT87GjZ7oByZsuEXM1UJ+i3iViu0Qq
fjGTqvc6KllqFvMjlyyFhdOdXk78Y24DRsUl+uT4ebPkbEEdH7p7dRQodnZc2Mb8
mN1s1fSgNZBG3RfgOUXO300g0DHzG/4l0tpGOHygo9l6R0UZcgvoj0ftO62nlQAj
x7E3uAk7xLv3mxiVAq4YltZxdG2qZt7G6i4CMKf82u5LyT0ODIFEXKBo8REgBZ0H
o41rhNVqjRQ5bBMZEBLaawxI8kxihobMon4mvE5OHdQfIYhlX2sx4fOesKrzw+ar
Q9aMLPnXNzYqYYg24I+wjfYMVFZJ2cXSPrkD/MgGCvGXBVCNyE0MwzUnkJ1GW5NS
Ja/CX2kxcN5YuHGamWH6gRCoctEbPHXBDwXVGlbRpFeQEgrewphKU0M+V0A2Hz6W
yIRApun+wR8CBiZPPjntzXuxpdSgqwBoDPhKRxWbIYbxCumxUOa6nBHr6BLD41tI
DU2pdRcSADmBw/+WC7sBBMkgY4e/oR/W21ELTRfqLnbkv4eQs9RY6VeLgFKsFSMr
Ap459+yTZPNVTB6USCUNLdg25Acc5E2jMfFwTXJSOTVEkhesyxY9CZaAkJ355+sg
bcZ25K1buYuch3IereWD0c0mb44WYoBOOfBs25MFgqHGswOE5ywXRQbNeHPuWtto
fMf37jzFnIqLM6YTGTD0SRZhWCjkKaTIn7y2QM1DzXA0JK2rcvh3AuZDiWSYRgNN
hxnIzmddaMmRNP9zEWpSziuO6C57obtjD49QSCksan6hVFkFxnCcmI2EyJL4ER0j
9cH6I+xQ+EzfwK+wLjwlZmfV74XU3bE2n/V1JjBAJXrAi6DNijk8srlg7qXUqo/z
5URLCjOUCvFUiMTVetAWY4qzNcF6gf4fJ/1JFAaxS9dQrbV6aOWPCn7CPINw2I2X
wjn3JN28kR8RRWXGulbE2Lb2NIbRQfaj3r65BdW6o9ARvB0/lUFbHjtWBG7NEhfJ
PfbNThd4HR60Z46ZIkae6shCpXBRQTvATyRhkaK3HaOWyh8LzwiW1iEEAcxd1Fnx
b0XrLz8cwk2YkFXxC7QwaC6TFx8JHkY9xr6lLFsS+ZAbRjTj5ETOyfraiEgk01Ju
TPK/9GhNbF8r+fgfabHqPXeopsvrs2OJ7vm3LWO830oUM+atHfdXt9Pn7TskudpF
YYVr9sBQsEENfpnQopqJNs8AJdfrDn7t81Ta7azuw4q6t61IqEoKuT0B4bA3AGS6
veSvGhc4lrnHIFlARO0b8X3DWJRrMpG1Kausvn/HUS6bYhg2dT/7F/cwuilPN51o
2mBKsDAe6Ks74RN3zW+WaryskLSi6FIK2/VBsaGuSFCT/cl/987b5y3tCFeyJNFw
r/x7stD/ifApQt2nVTAb46cWJ/j15lU/0VBE7w5LSw1zIAqXzZbaahOlnUuAGiWg
UiJXjFrZzdgnGZ5AG4oUJXbGW9TTbgxY4ig13Y0oIftLAE2RfRMrmbuTnSeiqqjx
j64RjxTZf7wx8e1ph2+RiLc7Q6wnqO9Fpxcse1ppU7xapUTi+70c81UBB33LIkuh
F52jPARW2SizoKdrBuLwqvwCgBXRE4s55QeeP7vEx6gySrlPvsbWOoVGiCEIltOr
5ljfBarvGvoD5VhI1g5XlSp0Y6ctb4QJyxMoKVE+iowzeiTX/QnnlWOrcGTyY4e3
xQk86/wm5OsmjQaEaYHukgqnG5f3KcJ9ZjPFLoPlej/oM4ttRDvBtXESyE9AzhL6
od1IFnBFDshwXS5GhjWqbHRKyBxa0pWNmMUx47USc8ysiF00hkbx7u6GMylRGGIE
n5gHS+VoN96X3xopgSqnIfZAHZfwlc7Se9TsEaQv6ITZ5PDadyav+00DXG03Sr3h
p3IGCTFAnrWuoEYASpHJ8Y99n7k9/edAOvfFhH5/wbKtNgYnZuk4Bk/M3U2j2G66
leknDohnvHrUyJoGqj/qYR0arKjBEm/G0TkJlFJtJVhp9+/bvXCIdPIpvveoueB5
CsD/vm0OHXjb1skR9tP5rA0cxisbYlVBx4JHl7dsgqUr5f0mk/disbXFJCOs8zuM
v+qg+pSwVXnTu8LqCaWyrdxmTZeBiAFXtz8xZZG1rG8s0fG7eBYJ+faDc+S8qBMC
ZFTm7jOPe8z369/xmTkYC8Xkk2nz+sYhHThibSEqHz0KMRYh2gZ7NKODxRsaWhZV
SepNsdvSB8FrSL98geBEvIWiLMgZOOTRV5U1AZJAtQgLVrpL4C+sib2idsxrmEd9
OjWzdmzXdKamPnYwR9oFUGhTKj6mq3Mr2sqWar6lbHY2sZW6Cej/3mp7rKHsu8vq
/QgZeziqQDMkeu87rtjYYZ5so21aKdRcki3qVEAyHBUYbKncDb4T1FUNMKG18kvH
74nolyrD9TygmbxbZTasI+P/dLDIVr54G8YXL+b2XV+OjoQIAWJMjLLLv+4YS+XH
fGhx6aL3YrWSFrWR0dk+a3AlKhb5D7izZTUHGVH9HX8pR5EmJ6c/3cYXWR1hkxvo
Zz2NmK5tchgA2VSwbFNORruHoefTeaLTMTr8rp5cv4v4K9LUsLcQ4h0iIOEGQbG/
FmI+TGAmVjKPb9VtieEDhWDzJQcsRMgMh4MDEI4qWVJs+/7ttajx3xPTKk/l519j
1O6Hlsj3dv4nJjq+jSFvN35wvK0hXmg/1nYrxZqhjB7Rphu6qXmIw0CW/z0banEK
M73VWLoijm5ypzSEf6DjmpZmvRy2UN/UrtJ98kZKqDY+5DJAzfDFwLuZAgc5rwtp
jEz+h5qtZ12z6cp4gd1fMswLRLDKeSJTtYlDxoGKm1pV/ph+wpyL5I94WVcaof4m
QzsELMY6TCmUBrXVHEnkWC76vR8N+aeVsfsezvGjNVadCJTMtotmQQd3CHOi4Ga7
bJ6DdHqrVV+8bx6niNUiWSQUDCbpGsTUIyQoNKslD+1wucdup6Hqpoi17wiCuFct
Z8MiZvQyAbQihJ7JZ+4FkdXniFuiApoXbOr9bqZFq3E9el73mvxs8BG7O4T+Jaun
KKFA38DQUj3H152e29djH4BiDs2a1s8akuheZ8XOIAirLXW6kAxCq43raGw1F8CU
+PjRA5nTSWOiuHxnzsqnzfk2haFR5G0dH6ZI7wUFNmQFX+9GEw2cTD0FHdUQzP7e
lca8Q4UQ4e2eR8NPxFymyd/vCzTsl8YKJiz4ffsf+hiTkOqrZOxUHITVKGB5fyuu
HwSEkAO7l3fqWLMGptsw1Q2fqtbl5hqLUmBGQ1I9hWgJv9hYIXxcR7PGodG+4aCz
32h5+mxaG306ct6Wz2CoFJpPfY4lCEfEyAUe+0Wj/g0TEJJlRosmwACyqB2GlxSc
VZerlG1kl2tofMNx+DGUHuXpO6Dlq5uYvbbAMWZLmYfcKRIvrwMjKajRB0FsuweY
DQahErrcDi3gVGDFYNHTym111W51MIJcNH+p/VvGCXDcpBPS/QPm9iGcoCeqwXqn
kIJa7hzmC5MynIqsMqcJmKs+j3LgIEApAPRL7Me5oHPdUEUhCNBeTUv9rmdUM5OF
fiEgx5Fc2+IQn30z9NfXKT3FeSovU27vHh0zbIm8TUb4ruxQPpblyQ2yCn1V/NXs
Ka3zvmnmcalbAEnHHddyUCdatD28IxbbgtRHxbOsFh0YTTzN55JiNs/Gm5tRKOCM
Y0zFJTBIWm3g43o7mA4reE91ihHekGkmSqiDpouSniwzA39bWo5Hif7nYbmZsE/g
HyOGacCmydLBGL01qevev2z/OnyFtJSY0aKtQx29RbxQh9mF4hZ7p7XqVBioFI39
TieS8dd5hAdNKZQI9Fh5bEVjyfLgzPVwD/qi7md8OQhZVBZG3KWJjip2X90ZLfFl
RFWgWuiERuGCtghI1Qfa97yqds7KQXRMQVrgAdCSGBfKI//b+ZS9hgilmbZRXCjW
NgHzjRjZ+inPbNJugoPmu7dsNpLgrLhTziV+vWco+7YueOstueBod8cf7Oejzvu2
IK1u6FsSx/8FA/qvdl0O3kdVt6Lm9hq3SEaeBKofNTVbt+NZn/hpjrm+048Ijy0w
50XaHi0JFGSoNbZMnKV4QnhnMJClzlu9LrGRBpJO+rwZfzJ1F59l5qtJTvPSOuOE
r1d4QRDuxFE3VKHQ1ekezPs0Q7zAIwcGoEd9vXZUAlhp7lBol2o1AXtSk6pNHB4E
BUb7LEnPB/IHPNIoHY+gJDvNnPyj2MQpVbQPDIHQsf6fhQwqzDyCUDCik6b5mvVd
bkgl1MK0U8xGU8vRVwjdiNlTRQhaCy+wKAIiQTxQ4cgTsRGq9oqrwwu9VzTEeJO7
ugaXCCcIysq/Oal/w7SkoFJzkX0W2mWTm/hxPCKarbZktqtVJAbXRVLp8gf+hFnD
fGPfqYtz/QqjF0de0pWr/ScLc+fVpAMSVZom9v3d3ya0zSxExovId00IcYybHawX
lAUOdh4Bzxl5oStmMpeunCOBj8LR+uj7L5lw894/PQJfx7DOxQ218By8Viat62qr
72m1rEqEL2LNwDItGcpbKrm/fajhIeZBDLgGVnr8zV6UqpqfdtWKeZ5V7wkjg7jX
YncbIdxAmhV7OWRMZVmbElXfMXjP5b++qf+RrJd1b46m/aY1L5rFg53wXrGkjnRk
h2XxksWm7ueYz6uraDesw8Mc9wlPE7yzgxCVeH+Usb8Cd5S83GzGX6dF4M/IhMyh
nQg/jOTyoXxlbMcBxlN8+2ARHbeIMUa2V827YJylqiPioq78bhO26GuB7OnvYby3
/FH+9SjT9NLt+CAx+ZIeErt+zpGq74U5JBiec3fnW1mmET0BoN0AAm/ZZCc8eq3o
Ll7qUTkPdHg6lqpEzdwGhRptaKXOxzATe9gOVixtvK6HZFOBxtV6alMYNy4ZJ9Pt
pdcuSq0EgD/0nz4eBO1w9E07PHsc2Nnd+AldN62lT3nXomxKlj33+CTnobcgLIWp
IFSs79/unRi3ad+YtUxjSW6c/llomLF3+BdqomyvB9kn4hFG96oHF9cFTpflAYzE
j8Wbz7OLsKQVdd/nvMpt2GoeprvDEW4WkyFVHu36yINt1lFZ24t8FCjNheBYdllW
K/acYfROj+5Xm6M0NFCNDvBp4//fWvMXNQ3/nX3GKf07JksY7dOtkVyw6Ide5q2K
Mff9QJWFq7SWb93K2MHNkqho/1V3nvwqJ/Ffc3eOnOvQdOUk4TQ9vlnh3ctcWBOV
E70nDPnvwdixWSecbpRgjSMB2VY8GOZrNWzR6DjvK72efO/bmzD9BgXYBbRG6BH9
KYoW4Xmw89ypltYIemRGJLZHuFLH5PyRrCKHRNiTyRE3fIx8HSBgcaGvQZ5P0m+O
xTCsdMniKdbAhs5zysZF7bRszsFpLpoPk2H8kXv0MV0FV8G7mrjT2FYst/Xs4qGk
7EQ/xtWg+K99iZQeOhtobEEaNCJiXGZuaXbOwNx4psKAMV2OOjTibU3B5aH2I1Mv
TZtQ5UhlW8Y6FVfo73ytOCiPKDYOSdzfZIrngUX3sQQsyQM0zC6VbUQ3jbyXQ/KI
5vFBg8OQaVY7haS8FtaFoF1ESZWCEi4NA5h3UlwY8qH6Zgj1lxI51DM13Hkoilbn
Gkdi2RsckDHbUIQq9QaouNrJnJjcu+n+UAWJ80Y2kbYp3w+xKBCBZgYqeFEY8IFC
hT94ipTgzyFrGOwXcvRvdwuWqcfqmGAHazIY3frfMlajj3dbg6iM7WHHcodhkwv/
qsS6V8iW42rJF2hDVVSZ8BEYbz5M0vJv2MGLHqeAsgitApSXSghsLXpo9QPjgdui
9qqxpHreGejFVaYpQ96GxnpSiIsja4IWwE1A86u+Xu27SdvGT/lEbx6W4xSMUQ4i
zKTeBiRzWkbKzcu6LZIvB/ytWtM4KLIuF+j/u9tlyD76Fg+LFv7aSWi0XeIoWYug
gRrwUBlUCl7v/X3GsdWQTYn/kaUo5KsFGBFBJgHVzeZxE3YXtj2JF7Y2+sQJDMEb
Z6PnHfhD82+WGMzxmMzBoudop7CLWfQE5NJoKtUxU7xfsfGhlXnTD8yw8x9ldK2q
gDjFpzSAj/hnC1cnC2REihkilBeq0MlWFrFB2VhKxzWSBgW5EJcX7pA+jnlIg76A
hyoywwUafvF4CMIKlnZnuqJ8OmiIxXKklVbuMgBSDI6WyYexREKY7BIAbk8F4llF
rz2olreWf7ypM2wlEkOtsDECbmQE0q/YPg4jx/hTdWOT6ROLTsxPGW6+Jrhu9Az5
Kq1e+sk5u/U/qjGhoqWSene0vrFmkH57VMRJb4OaIBxVuY7KkYwaxqlAQ6mc37f4
tnMgfHaezj92Y58Vn8JfoEwaX6E5gAp3NRBJYz3hqg+ft3c5MgfP74gSmoJzIXdp
3TFxg/CEFrN433v52SXO16ajThDH/3lDeM93fVyJGnUwaf7YP/cEZEmQA3tiRQrU
Jy9s2/D96Y+1rgjhDw3JRP+T1+H1gb6+jdsw5KTUAehapHiTy8zB/XcbV/rkC1dN
VMYOiD27x5Trv5ZarLcpZmbZGzFR9iD7uCAVYZU86L4gf1fG7OevT2o9yGPHGPSY
QcWgWmWWSyLyfyMeFDaBivIswGjoSCn9JcfSQFPoieYGW5djrb5wT6SNsIHS0O3t
38jbH80W6PJLYVm1DuZasOHI0eHksiFpoMuG6vveFNvtbOODy/KuFP5E1h3+8CT8
Pk++424+brjhpMVFbrYE9AlwoIuF/JJ+dvWB6wD95c5YZq9hjIHKufWcigBOcq6V
mPYVkNajxIYefph5QdbudDNDHZLAK5VAb3cMs7wAkvDbmKgk0rYL7FTtyFb/bem8
/iKoz2gUiYreYBgj/nuFxl1+LgOu2KlXC+RV98OEcGQWdjyCea4nvPDVDSaARvGb
wrNEVXFuqZ38x9DuvUuD1TG5CLj9PZZhmnZ5QJwCTDipGZtVwQX/3+rTrOndLrKo
FF/KcYkGDjh4bhEYez58YmijBprLolkHKShnUuXvKm5MEHusTvobi2BXOmjkPemD
2rYQO3tZMoN7CHT+Lxzf849zj0cWZKww4ESLaexmJ++KNx2QdG/6sgw8XQnt2UPB
GSHG0Udg6ednT6L//T7TonHHeo/7ajFz9xfymU1tpMK2l2zBSP3dhJJH2Da4WCB5
XfT1Q1dyqT8A+taokOd2QHp9lwsWTPX2PHLopThNgqUbmzELGF9r1t0nfU4/BJJi
lOYD0cTgrr/G/4XjCqQDNoHyzVgWZEicXBm/UrX90zEDJpZmDztmjxEbXAUiG8re
Ml1WnUPwpay71MdSu91iqdIiuDScbDmwWdm279ViAsv9w6T7GG7w1G2imvEGd/Hp
S+kqjt6XheHBndeeWp0S4ls11CGqI8iDuW59qeywcI2lWLQyOXSMdHG+5PAfLUAO
dE5+im2sK8IDVe4Sus/ZsEYjzM19xxx80VkbffdRSm0gCwrNz2rV0gZF9dfO/iLH
9Pp5uaNna7mMqJ+3BWWNfUQJg0F0ym3G9a6S4IATAe3lyrevdzKUCyRENPVEEXvk
6/F6RPjod3fEf11LcuY+wLYihntBF9z+qjIgeHQau5yMOAKE8F+LFN3uk+uC7kZd
GQG6rvmj7sudlpWlyUsYDECozywl3ErUopMPwGZLpc5+XKwlCP//eh2pyGXweJgy
gDpnzA/0VRBMR0sEPvSjTfQh5UbPk2/E1ofrDUDt93AWaZ+FFqJYJXwSqZowvZEY
q77RsQR/CcvfKkypGrJ0lrI6eGhBIeuahfYWdflIw2ytq2RSxleYs/paXBSARjGJ
aRnEFYgrDCmZxYcm5inmWFIOKn7l0M0EkO8yfOQlXdE3BDaqjOZS5BiZvhhPPdtg
C1l8YpABmpYHo3H/CFT9MsC1XVC5RBgd+uttPac05arn1B0e1YalLpY7b38wu2BY
Xcwl+e27ZDHP/9CEdraYHhDoiP6gdlWWRJfPo4dHZXIcx/VyWQXjMtmq7lJrgn5I
3ldovxQhIkBH3cq0VhWTNgp5kjH9xREiO3XBluUxBykflLTkvGyFVueJglq2dxkP
JayDMU3B06vls+UIERw+Vp4mbBNf9nf3TqwizsQzNQhcL6dzboN8Cr4LLvS3TArx
OZdb+pbiUYayXRRIOwV11gETjHLUkqT3FL2Ba0vrUc5hZrBNrq0zsTPtl2zG5xPT
CFX6ohb+FVRUqLnDWD6dqMOrlT52h50FgwgTpDN4gE5P+aLTwVQJhRKkpggaH7oP
IIU2MyS19pdufYOe1a/oHGWfZcWhSQjSrCiPh3n9qvPoA/eGbp9MC2wJPHu5NcFH
cN96lAGOFuMRCYB32+OJCM68jvTkCb+WnJFAsiN2lcIaOWbA7qQimA8gcu7JddOG
JI5DQFea1ICunqu0s2qDhwLW9kQkq8Ahe+lu6oILPDozErXTS6b8r0Jnx55Yqvf0
v6gsPlcPogozy1FWd5PhEz1x7g1kAgn728PZbaa+7M/YGeJKl9Dfk/vqxWS8QABA
Hb0OEFVwsyprhzcswRoxbml/66pWt47YHhHpPfFBubLa2Ly4GAldTBwepUJCB56l
RxLrP6v8DJVwk2DCK+BDXyIEAlOemEberqtv3Uee+MSd4L0zZyVYuoSpBcDXVvaE
hK7fDgb8PyaYbXecfVy0Ces08w0H+DfK8286OzFSpcQHXtu4PkVrjLRDH9gUDc2R
lgmgyc8m17TbSNTCHS3Rhrn5WHDpa3Et9D14qDNPvreM5TP1x+yGarFeeEcUrI4P
AjcQdxkixTH5uED2pueFCKgp4HtCkE3sp/nN3yyjEHzV0lsW7KZok0rbQyUMyp38
H7p/tGLuuuQibF+SlHB58tQvsb6mjVwJyZ/TdkTmgEKu5vcMtPEVSo1sSMf5j3JB
AOqM6JAK+ZMRAa/AtE/aOFoo2A2R8OkLCW+47L6NH60R8piIpc1Xjg5ZN1VZy+H/
K63vpFtzk3+hNkQSuO5paqvKA8l5/Y33E/AlE4h/fjJ+Qyai+xgAtd4rcj5jFsqy
YehwG7piCQ5lnYTeANi8ruA56dJRhWJLOCP77vWbAiZk9bOL/HyGnCT9i/lQ4FMg
vcggQyfZa9t0todlmIULJZ1HGaQ0saJkRJSeF95vcPTCdUdr1u5P+TsB+e1XMXao
deqz7F4Y+ZkmCdWDoxs1dzLljncSw59JgvdGxn57EV6PCqcumSl6OWxCtuyel5Vj
QM+whgZN8E0yW8l+m9Uzmo5Vr1bEe4sSuglg8RNdQCDZBN7iEijheD+Hjsml6wMs
Cmf2b8sb/LBy39H0vaEr7nIei37Kwo9lNCkemyse5/3ZdXsHCqJFdcrEkmNNi3+V
iA7ScL8tXGdH8xn1bkDoXU+BAr+TG/AjWme8wOrFoPwm6tHo56MlO1qA//g6CHge
44OqoyEJedGSEsLQeR4Zwv5GLjq3uUSS7bnjIlP0s2gtUwFvRTaHUIPjG+RS+TKC
bKTofgQJEdNXYwatqbcYwAA3/lw+8CfUfnaME32Jo69fJbJcltOKMorzLwmwACe1
5rcu5sWxZqd8tShYWhQs0TUv9tIeeThpWawbxgjQ6DzQTGsn9Y6O34i1xyn5MkLO
EaQ41a0oEvG0VCzDtW/ByZT6ffieFEjVDsPEN+PpRPoF1LLsqQwqi1EgwURMB/Qd
bn9p4N+edmEiYDl/kRAmw+fR0mc8K3cXsyOGXhhrlyMjmoN/zp+FmTrrdY2PzOZi
pephHnP6qmafN5XSOVUt8KEyNjOlOzP9wQ8SvLJHuuRbH8PQfmOn5X9c9JWagJUX
WfkUwY3aDHgN3YopthYL8W8OSTfvdubjSL/2CWZoLVmJwfOzbXLD6RN9/G5+5BnF
eiUzdpBACUIlcTutEoLfQ2+KUVY3p5xJ0J+UBxyRLVZPKN/2+gWkQRmd+KlY4c02
WVRpNUFlEn9HO0Fh44JlOnUPPPzQjIh4adr2qomTC/F0pl1CBaTnjQrAsqozNklM
2/2tyiUWAQ05DLHY5zFGSuqb6aDsvozp7fLIj40HFXLGlVDBNgzbSZLDFcML44Ls
D3oDNFo0qMnlOX/xa4ZO/4LvWM/6QmNVoeR5Sws5R7ynGA2KmO1eqlJqswrYGRDX
fWyitmnuKiyZncAvotmr0WWJCDLh0BEF+0j8WyLBfsWcpcA3Hk+VSx56jDjHrTjB
zpFM6H3e8sfoOocvZ3wP68oeCAysE1UR6q+EXdW37tO/ZG+9B2fZz00Usq4b0bxH
V6+GBL6G6wDjzpobGtIesjQ7AEsVhN0B5Mx4lEnXVTZ+LCI4iIXDuQOeSfucjb+g
KYc5fn9ih8uKXcmG+LXv09qY82Nclv00hpgDQ6B4HmnJfN8WwgDu2ZZyQjGJauID
wR0CUFIVCYpiPt+AtKUnZqj14pUiPSgXyRipXCw1+/Rz/x2kPGYOY84nB5Fg5ilq
pDsx8+jeGOh5wLdFwPDSvRFMPRluRtSL7gHbDVIve2Ff/aam6FM/1BQ0upPX+I/2
qGbFHlBk4w2Gd0jEXRW2CKVVD2sE6cErpiXeSxp2Y8Cmyrt/6CL2DGo9RfMB+DgO
TupZsOHF/pg5zXDTLB9nXSJ8bEWJmb6/h5Mo7BcxmbMjmxCtHBsnlK9lsXsUEjx9
veGqb7MT37oJloRg4HObB2xUmvKsy3Gjpl8sqLQDHhanilpoLu8XRDF24lwvgNIk
+W/08efT7GvYSKyQp3hm7BlM9xCOCaRqai/IK7V6c1heStHDUlAYGL5w6uGCs8Wa
ihHjFsd7Cip0zV2uE56MkoMUhjBlM2d3AUGzVJ2dNJsrRqz8fkcm7N7lpDzpqezo
36eAeMAjfkLUl9Gax9jhImOJmTFa4AKkK/osqMFwBdhpeO/KQEe5EmG2600ND8Et
AxsEhjsJlECZ16boAjz0aiBsm+YIBY3iH4Rh/r8RP+YF2+j9JIBRx3IW+YZ65exu
IGofKvxPrMfOnRAA4jYNV8hgruM8QKZkwTGk7cKlgtCR6TT97gjAaXiouFWMdzT6
uKYRqDiLiNt70aakqvoMvhJHSWmaah9XPKqewMLg67rP1FB2YSBiyf4stdvyVLX9
IktzjfaWyuk3VoREuMzaOqwHBbiFpTm2Q6DKeXDbHJfptLO+fOSMp5Vz8fomJswz
XVudTbRmqjrk87TYz17PoGdZXvyQ/AGvElrqJbFNMoCn4Ilfb0tD1DdhI+V5hoo+
SRclRvhat2EWS2Lwy6ZtSo8MKCPKATq30lIRyvYBg12ehBJjm6X+k7CZ4A08B6uO
J+Jov9rjoIdQJz2xRSXdcBmI0V/h8n0kbIOrJXWck6y4XfFQapSJLxOxi7WqHzSv
QEIjL2NZB5rRjlMqTNuOUqu718lfZV4WM4+FOs7AIfH24ezUKiuB0NFqEHgdQy1c
2EQxZJm5X0dKDTffICgcHegTwKWaEaiw1JvInxg38snMnyH6w20Ov45/2nB80RW7
JE4cB/g1nauK8opV5rk+NXoJa+aQF0sfCt9SYZrNiUoQCcEeLk1HiVX4BFjCCV0t
TZmALlmSpSdFBTjXE/HV5MFBwtny76WfWhGmQ1TeftkzP87nlJdoTLlROSkzKZyD
dEriGm/vzZ0qzOs0d+PKEDSAW0nKpTPbo/FTl4LsXjrlhJGn1gdv7QpHqZMd9563
0/6b+qdpbJCehGGuMA5LPmn/+0GbW1AJjSNYPYpjk5zZgp6hd1xLadSZqMMtVZtq
pJLcmvuHqWXRL4JnBGS6BtiFLXN5nfLbiJBveAKGm4BjRPzYBcAeUOMG7oYvRd2x
i340hTumXhddV1tQ7WstqXrYTQJQB2nonZiaqdqAu7uEKXEPLKE5wfL6KF0VO353
0kTKSy5cBbwCsyxfxLkP4mT7UQAReY/1b3FpGNlRNlCbZX+XuF2PLwBxFTPSN/hs
80e4In9LCNnV8pEOkn1Y4U770ejBTYci/0Iu8et65MNSzFNE0meAclu/DUr9B9rI
Ym3uEuoqaDOXzRKnchsIuAYjgm95O+cPgNGipnwTy34/uNzEmctsbz3SmBzKJd1b
YJZ+uwGpGadFtD07bhGbHrnx+pNfk3WDAKJf7pOfNq40VJ39mpCezjBWsqX2FcHu
7/nSiB4rz6zVdxwp1J4XrTr7qwqHaHM/MKB5O8Q6pf3D2JROQwprmbY/CSJ+m5QD
zv8ux9Kx7zgrSDB6oth8IZrx6mmBnhaaH5IS1VzhGPuLTwSMHEy2aw/1wsKtoN1u
YlPf+whYbqyq192jIIKIZpphAr/h6Pdld7Qgu8r2jR3lheg9yNpZkPcgZTR+ZCCv
eo+1B0fbsxHuOveBmUCMUPjkqwGKjQKatwNw3M6Atxc7sP9d/BXxnMmFfvOGGSb0
C849NprNjsugqNRXCuyiQWI0nchOVAW5iga4c1PzR8L7ENQW7ILZP7wbrvK/kWZg
0PbLBZe9sR38gtTpbhE5KBsctmYVTd3Cvx2oPWrOVUGQIqhrvRRMEEdVrDVpNtF2
Cmxdo3Eq3Oz9XKLPmDTEwut6+qAE91zFm3onajtSqUb/lyOyazckbbM0u70iUXjj
EZHCArFzGfHZyOnT8oNEl9miupEJicziCD5fY7dzrNb7xd28E5VdxCCxbGULv106
MAVDDCtad8pu01SDtY+NnERimJsVIyZ1Md/N3kN35tu22uHE5t7evw1489rtWKcK
thUt7lm8XxFhu6CUe75YPWXKv8tdEH61m6qc6vajounPt5WOkMe+/fPp3FYz8x4J
Fytw3yv5KwKRZIopFlEp3M3Apg5M4W9pQBa0skvk3umflPLNHymYEE12ViPx48yU
Q8XoSLpn0U0ppLKRLoRgyO/2M96jATtsSlMYn7lXkBbVX2VaDJ8G+0II0C/woG3O
xPbyv+i1kZ8OSCdhruq6eXEzLushGFM0r9UznHJ+a5ZXZoB97FNtP347+R/aRxqX
aRLlb+z7iJEgDxT7HUxyGy/n7BU+VHIt2xrfBpX7HVpyrHbjSbRQ4reHwG2C9hMq
YBFA3PZ/LbULNtyF26cT5xsycZvfkBt2Bgb7DQdt/IDmg+5l2MTiT46EkBWxKgMA
4HYV1jtEmWLf+yTTcdBnT++SjOz/aXVJ1Z3NwZDdU85iIIDEqOT56UJ+WmPMn3KK
ctxxozDySAI7o+Ojkb83j12XXeXvhpXNls6Yp9SXDsvsB7mLQLKdnsw9HInzJUqg
EnuV376UxS9q5BP9qD5JvaohQMYf6xlvfVdZOeVLfgxOaEs/E8VyisxsuQfFtXOD
KdFgXO5JLLKU8jClONpj72oP1f8wCPEpqwcdaG9MmxIMjOHTebsTYKHDtmGRIPgd
K9DPSSI02zZef5c0q/Ps/faKF9CQda/djKcT8RE9ZoQxHgpWaU3x0biMWcuso3wD
dvQtGeKiU3h86laZ933C08cCf6CSZYCSQhWZWCBNtvcjljj/rKGTS9OhBIGkYBcN
AYBE2VFPNh6G3G6Rsya3yv6w+pVBjNzIZsfd1J0I5Rgw0H0yk8f0T7qZVSEUJW6X
XxAMclgfiUeV8aq5XRD8fLr3QXl6GJ/ye3gK9FOO1uGjKbVN22uzsNtwFQ3ZP8iW
hCID5DNM5kLd8TbyZQcPqcLJ2NlrwNBatWLkubx4yHermaMaqmNxULBOQO/tZGfn
WCazY9uAM09Y4Tgm2Ot1Jfy2d0N6nyY1mrxIoE67f8oKeoYrF623anjIdS+LsaGu
gdyU8+JIeIH13j7bcQl2niGppy+H124HppW7ZdxKXSFEz03O8OOjrz3D92i7ZDqv
1GCaEd+wDYSbgq4/EXVoPFUUMfTYypwCq2PLVhrVM6doi4XK83jLwxvt0FPnO4fG
DE0qgCpu+vM3OXVg5lTMCTiJSOwTlGiMVepuwZMeyZliBPLRJjF5LN2Z0yn+pwx1
LJivgBVx9PhOIdQ6dTuU34ijPfmNm8Lallt7vxQ3pVdmMHX7hvQt1pJijLmhaT95
2H3EPLF6R2BLW/fGr3lovoUeuczglHOxcSypAInVIOiMuBClORwvIhqHGwo8Lecd
CixdLZ6/D7w27Ok4+s8PMuU0nALz3hRe2JJ5OwJveHOtPCKuwwoDO7JD0DXfSLeI
dl/jPqzARBq2ams40TZCltt8ZZLOjXRZATbrQvFWLKSqJ/640TIRbj0BF2FK4g4V
NRPBVrBaG74KW0ADoYcsWCy4y1MMEY4+vrNYQDYA8f1LDrmWEdHAaRloeiwUHH0V
FG7zJLuPgfmRIgYiCT4mN96mon2LD+RuPp/eBZyqYu7/J7aOVLAPBjm/J2+63W9i
Jl7hcJaGHa/btcZKCJS6PymYEpbTe235+00Byvzr8k6gnP93bqH7gg1mFKyfqRuP
/ngQUuDFUTJy/gDIWiycjW52wQuupOMXnC6Q5YBhrjwBUV5qjBSK/43Y4vsFQiiS
Its0l3QfECKaSGhaKQkM/h4X3lQz/47GhdQIos+R7nkaH1hmAlqfFLkbfJmWJ2c3
JHquCxUVIxLtmN7ufHjHkeGL/EAdlksnZWzQaHp4bnyXmrZIG6jJbUTKWHY2UT6d
91/Ki+cOXfK46FBvAeKHrByki0uWKrIOqBmzzpg2uFTp503OdoXdT4vIXj2uKUXl
SLc/S9glfmilfpqJGp1oOEDWSx/a9sUFk3OBy2rp5T0rhvcyfdUmxUK2kgRqR4bE
lMy472cEvkZbUt1jn04pKvi/8F7D37Ij8GUAeKW+KWIEyVAqHp+Nla6zslJxsK/H
fQudXj3Mqt6KDPgC4XhyPF0RQ7/T0bt7dtObdS9bmVN2MrL7de4GXM6VI9C6Fbnb
aoS/zfId2yF6mnF/Sw9kDpvUMGoDXUYSkKtdpldNCe2DRkUdH9MVDB3rvU2WGQCy
NN+8QXn2JBFr4Ut9JRN8zsjUTogVMkOhlMu0fFyZKEzoIbDj56QelWwGb41yWz60
IOLtf9r1R21MxHPSPM0Aixj/1aFeJRyNc5x1EBDqsZ2qpEMNTpjSR56qUNcGMF4l
YIHQ7VRRV/YQYg69tQxUYUsWTjkHeCOfUwVJXlzuAE2oLCCN1p2mDCnPvyt9Y/TU
bKCT3EA135dwVBgKQNrD5vt6IHK8ysKDW9IYzaMetBiCXcHl2+IR7eYYEMj1tqko
Hh7CQutU2wA9pNpUVarX6mhOUBiXUDyLA0FF5TI21X/0hkh63laZfPYDUKraHJRE
M1zEW6vaTSOPVnznhVHBOe6hPAw+e//QJVnY+bWHZKMx6svdmj0HxercPCFTTse0
L2FKWkRG4HivJSHfYPABLkK8vM8SIMLZ8ZbnDsR7M7S97H+gPP4ZJzQC14UGkw83
T3BTOM1kVurQLPFyb6AzLyhbSkL7oMDaiYZB5np1ECsEfH1v+n4APRF5y1kEFQXn
Xg/apqbRcCV5xGPir0x5RETEelpo/T5+Rf8N3NgVcTUWHGeuIdtBpMqo/75FSZ3M
5pZS1UZ8MfqCXfmbgPwxVJVMSsxzGIWUFA+8jXQtiUD27auN77bvg6peu5IN75RB
KJev55odAtHQnVnh5USnrv2VwWHbuXr7GaRSyUhDxRKk+OPNeXvLHK92K1f1UJgw
iP71qFhPMxYJ1YVnqBk3xRtVxHnErige8+4iyUj5Ws6KV/4oUd1s3xHJZP9JfX4g
gOaNeyAjWRj18XCoiP6SrzqnQxFS7fo+2XWJy704X9OB4LPTdl2NvGa/VczzJKax
BHDVF1Ceez/Px5iXGmZVcplXRP/En/IXz4t45XUDo3LxxVX+kw+v8BW59ayh+kTn
nLvDc/hEgHy8l9sRh1mLm17frnNC6TPql873kq9i/JKsiKard3a18pzCZ7Kk8cX2
+JK52+BWyXzZwYdPvj8GLsF8Cjac1V3aKTPcppQboGBZ+kCz2y34epc6I80Oh/N5
5/0AEPV7MkjUwQAuIxgb9e/Ue8rXNkSm+Wqb72/lYlD1roNJgcWZJfZLDjIBqf7B
6jwMdakBI5vxcr0RAX2PUkldbSs+ZErabGklVatDOlCBQ5id87Npd5DrpqVVUDnD
ODkvE4f0ld8BNL6YP9jETNhAU1Nvq3qaU5ptfM/YoGzZUSFaOtPh1AqVJGxyJjny
Oj8zK3LFqH02blfKsEC5Nylo1KoI8244dIc+GBmfZXP6+PUjYCe53J4OEZa4U/EQ
E+noxSvrlqhf0ujTUJgiqGmnVUkPofKxO2f6kYW1QF2b9RETErnxmtNMJH+pziTq
qnzP27y9TrqHyFlbbdJSw9T9RqpqZjp/Mk/pq6/NvWyiOLkTzR+dzMaDlcorVnCq
qy9c3ER6XyoteHbwXIcicbEK11SBJS3grBjjQsbYwkctC6Po/2MWqrI2VabT7xkv
IuRSDn1dMaT0G/Y0Ro4hCs3CBmMorf7d4s9lQi4AilThdB8ApJpqKJ2vds/eoYmJ
WkGYQH5bnIcAjku4btH095YMQtRZB0uokPoFyxIziiRwI1/p4G5TTxPrTbgL0tt9
i5yIXs523JyRgo+DL3v+Nrqb3Bw5yLQp7oCwM51keHf+F03Emr69OQ7fWpyf4TZJ
s6jH5D6onSg9PIBTta0ckDCjhcSZQBkPJ+DaaO1eFL5Fw7669FDzdupwzA8yY/uS
0MXow9dOg5yWMX4yd4CUAdmhyg+H7kzesO/6TUn6n2BlIyNNot4PrK042Hgrqb8p
ijGrvj5FoHQl3iBoKw46a+w2Kr4J1FWEZ5jdXax+MM6IWhS/R+1NtAxdlUX4PVE2
YhUOpyOKdWfB6gOiW1v7Zre7GKWF+UCFZ/2WFkHn4ZA2wOdXp99oa72mpBFDu1R9
NfGIsQAtOkRshiDTMUmiAlWcz+T3ZCQlM6tiVbSp68+q/U5eVmD3FIf2Sx8xAHXA
FQxvF1dNXQ6NpCDwd2QGUdFPArzCv6Uamid2GsS1icVJOhHWR08ucqvnSEXaLx38
1gVh8uppzfLlvE/rkJC+ksRe+Wj9fVCWHAsfrOgADsEo/Mf/VoMRzdeOdZCi9f0F
HagtpL39JZObwEZQ8X4U3DAxCBkfq2J0yIPKbNHxRbovBpVNlxX/DBWiIRAtHUnk
ReTAG3BZCsTIDiGAnd6LUTL0xZVLdiqa796YH6YZHtxJUqoP38SOOEmY6BWeH2hQ
N+7B0h2wwcyebZ51AuPQEPrGW3UvYzKxgHeNGFI/VNV1gsamMoU8AViOAk+XN2N8
k92YAEwd2nzRvniL7uOU4juq6SHx1R2nDBRm1gGWYOFVa0yo3A3emmvsUFPMVE0u
TgwQesM8v3O/B8A4jg5ifcNeJZYbjMadyBVjflHJMghkhTPPyHFYIZtSrXz/CEvQ
QMjJDilkA1likCD8Ee+/213qJM/FCQp2BLtCeoZp8UCvrnSIGINFJZBMhj3B6sQZ
VbteN7sKozB5MKLSTzSdulljCap7+EqC5swW6NksqyYO4pvM/gWjUvPp9Ys73wC+
2No/5dJRsdSn9xcfjoL0UDgv5QNiwiZRRnonleZ1BIST5vG17nmQO0ftD0aTFoWg
7YBMOyWWGXnVsAwNe6awqosdOsWVL9u+bafKAr50gBzul/S9O79p/e/G9Y4V4/Zm
6HGZQF0lYUqdcF//sj1g5xwt5ymc8Pny0CNeoRtflxkVjc9N+KArrHLUwIpkVCSU
xdeCNrUNtrNsrAn66KuWjb+f24STyj7zwauj4t8caOcVdfBskdRbbIGyrM+Tf0aA
2OI772Sm498CDYon9YFXwZdkYU+BbT40iNaHLZ/xyePaQRMV7qBjWss4/5X93Ey7
aSYsW9iyX37G6mT9bxrB2SUK61lwDvQGP3QovfEnBj0bZBDtJomML31dqmQhB3c3
ySUU8xPopdAd0ku6iqkGMIw34PWUaJP7hkFfT/zzWToFHAbiBl+Pk0vufPeqVMpm
Qg/lj4zLh6atPZc/1EQiD8xQCxIsCidNBhM9wPUppGM9TkzcTyfjwjzOeJdcytqm
qorCZo2rlCDMPZ0+FbkzzCI6+KLXz2+pAjEvnlEdAOgGFmYZB04BVNenlAJLDVCO
9z7ZQsqGHNxyDSX0lc+NyMelya/Q4nq9Tv7RhA1hN/j8hhwUOGVXAR11f0Z57kgx
marvK1W/bv8J9Qz6z3Fv8/scAgmk1e7FJ696BM2Nd2Nu2rFm1vifOQRqph7RnpQ+
eII0MjabAF8cWmqifA7rDngrvF2Qda+EJGAOwGVttlQRkGKMFEdLCFhAOQxVIX8J
eRg9VYLznD02S5cTUVs+3OR95nGnK4u4pw2ioLWEGHNFjTI0pHhIhj/VM0knL3jR
a/zZQZ5SPCaHYhL7siQ/xwOYPsE0GnXmtJjWuaRfq9/I+M8XzmLvBAqcWlwlvWqC
6oZhE2irjWwFaHxcNu59/bwYjhgR0zgx3sr/2iQ0/GqPHZLCzzIcPE5dZ6AzUHAR
yUu9G/qAy1OJ2Mv4A5E0UmoO+HhtgzPQHUP8EZXjSYcasN9/V+i6PBT0CDOGKh/1
U3hnkl7p/ZrUO4VcUyR9OXLxcYklvjuGQTMm4Y/piV6cyMpU4eCpyqZU0XUEezmC
oBaXIFrTSFJa0NBlmh6lD2yH25qGiP7BoUc7hJD7nLQTze2HlWHY6RyDZB30ieza
57Nacu2aaLcprFc1IKMEObLi7eM+2SzHzUoTqOzaSzIYMapzZb/WAivb7xIEp7cG
E5qV1vcRVKcrEXM9xRrUuHcxGV/61XM5SAuhNDjLVulINW1Mvs3P+3KmXMVvVFPE
bSaUzQFdZJSdnoDxy3fl7uInBxO8o41CWFrlyNzNqbzFCOzvcq0XGkVbpbQ5Lh3O
BflYi9TmlarPFZfoCck6fEq/xQFi1GhiY/v2HFR5zuISe2teBZE7aHlvkB350dK7
rtGtSc1ac/KrYVxbPUarBzpr3T97AMeC5l4y82poqJf2rakjtdQydoA+nuxmvjj0
98ITgvZYcvWTrg8/TJYu4SO5ADLOf53MKe8LM46savh1bLpZg0cDdgTb4Zg3PLhi
KrPHn4lTRjNzA/+QQJY6sZBdv1OF7HMf2uAo+PMbxJ87O9+bjjihXhyxE7JO4Bdq
i4dRSXEc2npwkmodX3SnPTBvPOJAfIJ1VxubJCkap7RDSPPHXsoshLI6/8ka18IT
aH1C7o3IdaWATqotL5KYEByd2oJdJq9C3U3nUYVSmqdPOnFCkcsUz8fatcCjrSY6
K1utPU4wwQ9AmBfspJdc40faszhbeM2t5CQxBlwcEwocqwxTcZRxyuRUztDoFAk7
7EJF1re/f2G0EgiT8wF3crVmu5t6lzKSzlENIACqzcwG9zb6Y1mpVDjfZyjRNLVi
ZcxSySefsmD3ysRgGJRISEghnG9jG9Dqozu6okqOUfnkBEG4FMyIViTwMRH8ZIZx
P0uVwL6Tk8R7+JEOF/UXIIHvhjcYk5rmzQP4MXRjHV5KMgCbjsmW1e4ayjfBN75X
aM8Q1OpJgotPFP42DA8qvI4gys8+6iSgaaspmEK54mfo+gKfnAXAX2eDgUWmSqQM
byT9uiCg78X5pEjJ8K1I1dnx5RMlYsT8XKWquEvVxbLakEU8KJyk3BYPwZ+U1Mvx
BKIXm7xIIuEEeq/mkx4TRKqDFS0GUY+gbZKpolyaLKIjRps3CRHIxqeQX95peI/l
o7iMyiGqQ/D7ypkCFZvkPpX+53nWvhLVCT6J6UtAPPSexZd8UqMLPNWdpIvVKTTq
0T88qQfC01GzDAwHsngFeRdC5kQNMMLpvCXBAbI1i0vdAFCR/+oJ6TUsLUYJZqmb
qYPKs+Lkf/wzeYW2hZw++j3CQYruWn1fzzSuCUSFiRlW/POn3HLoFnirOCmjk9rm
eWUMpgfUg40yust9ubt6b4Qj8D0O0yDqBghSB4T0PFXksXB6NRlLLJvn5dKEFOsO
EDmtEnJhuV+5NvqOa042HQqT3kLNkFxtG4wdOzmJ2V9iXH0NPismSAWMKW6Ic0Oo
aHWBZbIJkzRcQZ8661Ch3S9xRxb2yAnQpDhPUNIOBYKmhudcv7jOeICAtzJODWUL
zByCZvLKElyaDjcF1Cd2CRhnGlWnxOpTLAZ0Bh8VxqZ3xdd00fxYyBZqYcT2kt6l
M8TUJdycZMtc+N9JY80J087ncq7J20pPEIR1R1ujt7bHYG6vevlmtFqkta6Mj/FA
3tGTJOTSrruCINkETUQzbEatiBLzj6NBrZORzHJ2UgPsDV19L5fBDZkEebLjff8k
p7lVHLsTP9rOYPaYUT334TX2EKdccWOUuW+0/uhdReDH6VPxudfSJwtHy4g/qN5S
RK85WHQu2FfUvo9N0MzM5qvMXiZU1EPa0HCSbk+yno/xEUkZW04lTuf+3Jws2OQw
HEIJAjyeUTMRBG4yPt1Z/lyCCfVG9jyf0cX92Vf5vg+UySOyaNkKOOT4yVNJNo2I
uoNFpDBpccuKVv+cDAoP8mH778395N5tddBuds5YQMZGjn5xi4T64yZ4AcQRgyVD
37L7AY5NxcSpEyZ6YxADSo45QhTOEq1P4Qwga9sBwb6xZ6zg8syBOUVG+Sy6KdnY
53ndCICJMmd0yzAKO7Q/C5kN2bW1F0m2DEnO+mb9Mv7MLjmk9lI5tN/89nLfREPS
Yne1tY1hTJzwot68V4wTnTBjoqzNES5ItUlsmyfVXbD0ERsDVXxQ+f0qKGTWTcBS
O3ihfA9hb4ISecZEm0vOO7CKMEYT06QfqldlcN3wDrJMZgCjsiG2eR4B0RKZUprK
rlSyoYGMHDbAQT9SvMG9MDKXz4RP8ImAE1W0+zc+42SALrFebL+oWe8N257TnvLq
vYUXBcaXoHCBU2K2s0MmS9CDExwp4O2S2SjGybUkxTkrVbosD1eQ11I6q5tRSXpi
YGbwqwV41sun7fAE491LMPUvKNh8+WlSpX/F2MDmUYmSmvIDdIuWFc5ZqnvvxBdJ
uot8Spszwglso+gEV2V+ub7MkJOe7sbkZjXbmtAKd6RYxtWEZ6QoT/abg6q7fuLb
lnv6kaRDxVRtSyFhO9sEWGIxLrHetjPh3SomZr2we13e3Eu8qpiPVdT0NYjfhQDR
52YkgpudCmVq5yUmytYw5PLYw0OA3gxaw0eubAPXrgwm4NfdDFOFYie5Wqy3dElM
UUf9mi4bv6nNsaEi5bi1AY13+3HoDmucqGnOHzZb4nGoEakccg4Y2kbHTSiavYma
LiR8157QTRywx12A0oCOcLQ905yBRbE40DQ8SCmMsC9PnazieUujDUoejH0Mgxwa
Z0w0KPxSQk3F4yXVEvszI3800EuU/Aq+M6e6ZfPpsaP5kpVidVnONfAqHfpJPTUJ
7ZzF1kBMe8Gi5zlPXZ6IgKWS4SYZlo9qFk71y0o+XnpQDoHHKFSXVAlhfTBDpBJr
nZMiTBh6ThQyIvCCrmgdcB9Vg3D0IJvVk3EaVJeoTDwxPv0as3Vf2h+I97d2Wflt
CZpjT4YToY6zHKWjWCxHlyqwmcmhJko11r1bqWfjIcC3Y0Rp1kI+wAqZ5XzqPAEN
6U2uyVFpd3I2sSCy1qBlp6YVme3/WbUP7OKs+2QYuPEK6wZg+HHvXXg2tjcz8MM2
arE0ED61xA9IP/K7dBjzyCMc0nQg8O41qJY10H0I1Ws0PJvn5KV9qe3v5LrbP9uL
ujPKWNMkyMhyKVtlfzPq/5PIXYIN4TJduuqy8iQNicEqJOk1whkRr3s0gc6cy6xy
wgM8TuylCiihQDYTQHLoeiG9Nciw23nDBTFR0M3Ant8pJHsAfQaMGCCL3oUJ5Qxg
YiADwT8HmSJHqyibbyTGtsYb38Mb/zQfCKo8Mh2HuF/HN+I3ly1yigtWL4DNg2gI
Y3Bx6Shq/hNWbDu4KWj9VnDIDoEW+qN9xoBmp8434OZfksmzrkqNBIgAxShU24Zf
073PU44unrbiQ3hJBWFQq8ysmlpYravgy5WMn8Rz/mTTQUkMWi4mLm2cfGVFtV1n
jNrZmyOp9pUcYSV6bs0BscHsqECfrYBcC344rIHqVBxGl8o50G3TW6BP2dY9xbDO
e89uQLFkJpCN1WymI8oxgoXBzcPG1UEj5+U21xkNemgSjUqR/x9jEHztcPCdTTxH
KWREfW9R1nrPkHA9BnPvxjGPtqfayhareqnvF2cTwydj4J0RGqhkZG9cX+5XLEM8
fFTp+IWU4bt63NK79mpf4kz036YcA8dIIsNJIdIcOLrZds3B3SvLZ7T1OMrGE9uu
EuPRtaV81zcxems/Q/FaaLC49zWa6RnOmt/J6ZPvgBKglLK0zTxgGH3aMgvkYHLt
K9xl7J02lYL9xsVxyWFjzuccD/jcPSWKAXTWSi3LijyGq9B2mpKB1NGZutiuE7a3
khPsFVDWT5YAGmXaS55XEQtSEHWBnLwcSGZe+x23sdRLTvdgiu2tbnf8gT3ryQaw
u/qz7OveyG5wJUjXODGuFsi4z5UNFhf8H1wsCHZKRpyYHu/VfPzF7x4xP7yNmUHu
gc9kr5nr9K3F8UlXtgWbSJGSfb+6f6/QETo94pnluSK/KpJ0Kgb+qpYLtyMCBJu8
S9EspdBsngJsCQ77wpfzkDeZoPo8HELCYxVD38WC6fFXQEhnPEFFR0r84TVoKBov
Q/QzlpnFxcJoMWsUcfbUL6ZeEmFAXUfzq5uqM4MlyGKhm3pznK6lN6ND68BG8zgd
bk5A7C+CDE3knXihtolpenIW8igHffkRXlwJea2/SuEMd/8NIiN8BDYB91SvnjwS
rDlGaAZvkB+cyOVkk3Y/2tiZdrqU7SXW72CTSAcz/IwtVm/2jHw6MmW7msD7jhd9
kIIpqY6YSFO534a22kNLNtQCWuURBSNlaH5Pd65Mxo+g9ImmWU3No0EIJIfRWUyZ
W63k1lPk/cwL2k6C8WI688Nmv5YTrfDBmAruao7yq3fif49rutdG4Z92NIv3gTwt
R1t1vvzfzQm4WqiHI8MUPw+GGJ0ORRUIy5L4tv8GwHbHcFmmUHXWd6Fm1TQSJzT6
cILwaX06nToIXjj98bl43SuE0W2XR8er5ejDSBaIPhiSY6m6oyrXIFhtTST7ktBm
GvLvPqHIosOUnlZRYd7tpC8AlvawpVOd+3+70vm5DkmmE9FZclBOKoc9anxpOxEJ
U0HFO868ZYrDBXddFwQ55joHh1Pc8zYHEzFDdOLZCEYsgNTbOH8goxZ87Bgn+Ljs
4PE3RdThZjX63pCZV12Agl+nZn1+CwpkR2y7gnxex8QKIYJAis8XtS6jyXl3vHeR
XzAKEv05TURb6Fc0cKgSstdE4T0nxhR654b6cpQe+JenzOqivJdofuVdhYgKKzzX
8w3J95GQUTaQ+Zaf6zzJJs8CFSeezPnf3/9ww6HvQ7SWZvX3InnzvarsY1TXu6/R
8ouP9f616kOscPQ1IbGmKHfc+nvf42m4ygY9RaPNQXyHZ+21j5XEcGF9fg1h97AI
j0yORcQ/lSm4bBZndnjnh3fEbYtkxGDbRENhhxs6UEU3T4mv5H8R7EYvvAgaEJ7R
F6B+1u72iw1m3nYYZc55YHON3qMPZfOW7uiLjHsBtQOxXc0JmjrYY+Yx6bkR2zEr
STZ9yCDCeK1Qy170QSzgkmfX/yPYJ34QXSp+lfqAS0pIvT3ZM+MN0Tj1o/B5vf8U
L2x73Jt72LzGM04NRRnpmE9o69J1L6x/LQ6ceHTTajz9jfbGqi1/xOJsWvTFIACb
4IQTwuiTTUFqSoFgZ0aL5X7kgBfQ2mkT8eeacBTUb3cgEOpG7cqHBcAK4OOi0pQr
LD1UhuoIyJo7dwnWiFHwxMpVq663hE83nvAaIE5cZBB6O/05c++bJzRd5BHNmL2r
SAYsRGJ6DayTprSuwMRIT9CEH5UVM83evSXDe+CqppSVa8K7kExjqd/42T00hZQc
cRCKD+rKJ1o2ZI5ydyW2YZabZ09BoLLSFB9RFw1ZiEZnpg4Ucaiz3d92t7j/eS/g
VaZfH9Sql1dSSd4Mfut+b+Nh79cizzX/Zlq1Z1g5NU8U5ZmkX4vVJqE+KBhS855T
Ivii2Ib6/AEjfrNtgai8p2lV6tDfbM50Kp22ktibePiJOr+e/j+oqi3VX6EWx9GO
CxAEeF954fVIVtqPLbmbGLtlu0cnFtvl55V3+KMtNaBIMi5L92+dTa5Vwi7evVMQ
2SgVueuosPEmBETw9TNycsIeBo4yiO/nsIU0Xh0aoVMKTJ0z01S6jfUjTDx9eqK1
og6VAwxF95PVeue9ovalD/I0CjjnxCCKa4gfc+4Xg0Sohh3PDpwWYL+M+O1AemNq
2j87Yzl0o285DIKmt7YIME09F29mNj20YuFyl4nd1f4+GhvFEavwUEORyl+AP27Q
QfMHXMHePpsivZm+r93xyxkGhJUBtCdM0tzII9rPj3GbHMqSBXOEQYSr8TGvPP1H
V8YjkYV30xR2HBmKgqd4qU1kCmGs8d1nnwIAaFBTUK6uEVgajoj0ma6+000+Fapo
LoyJlHha8AJg2yz8o8vBrV2705kkHZ90JjWeIAhqq6PrUVlJHBAwe7nzhFMCd4iO
f7eDH4fLgoqTEOYrUGwLuzcxDio7ElHdk8A9wvdNUd/tYWmEYnmHKkOFPjLgsXP6
N2PKznPChasRur53ZW9u9N28gBE+kEwPQhNesJdUhPwGzSkdqL7WKUbr5vYxxt7n
jaD+XUhcMQ+CD8r3IyMm6FR8Uz0ssGGabGEveV+mBu9p5cQKZo1/8Cd5Tt+v3EJ2
Jt5qENk7qQUUo64dEZAfwnluOmfQmTZ/3ogxsSWubZMBqJSElEBWuappzVnlO1z+
ZXUyOyo5z0FSwMvUadnmKWYTKIo/Og/Xw9PbOA4ezGdVy5f9GWCODnG3z8KVNwDJ
rfMPwfOuz8LQ6S+SRoHj+7QyrSoTpsXDlsnRFQRJePeee7YI57+UapBmNW3Bhepa
M3N0i7GBe1DfIUAdnNnYzZ7fuv2XZutZ+kq9Carkz8a6HW7aG2nUPPLkVNl4A5qL
mK49cigfp4MOhAuAMFT+2PcF714BT1BOveQHej+NpRCyE/syoMYwQcbIBCvS4gfK
ChVBTMM7oq2O+uYg68mR5aOnG29mXnBOSfCQkVBlV1bh98HtsRCdPkEmuseE91PB
MiLxEqtwIXNXEEdjRqMHBmDFdjYLD5DJ1b+9OexrIaLTMEGyXsZ4MDU+azhGLotO
IXMU809vJHUiFUryceOFxA0lKx2Sj3FbUS9OLdqLF5UPdk/qbBy2tv/1xDO+jsjx
WxhL7he7kMyyGSDpCpCJkTSjXJVJvSnfRCdo0c7JinyFZt4sd8fJr66DLMj448MQ
76E0EvPdYYj6jIkgio4t8iRoOYlLkYGr4s5KNlHPjLwqKNdgq/dEZV1JplenXOEu
rG7WuinKAa1QIJrbEFCtBHTytaqodeMjEOjJOJjXnNJ2KSe2uANv9+Jq+kA/BidR
3W94nqsy/b4kYi1OoNJGCtFYNZ0fw5zlS28P39+zUGkSXSFfaLYr4it6uN+I1mwk
lv6l1HMgIpStPySyQX4NXBnR8SD/9j8AlaoNSoyCnDK3Tbk0BpXHci+8/aYB9tu5
HMO2rA/3l1EeZUTEZl9HzcQJ3d4qWPLAw6gVFojvIvKxHGueLoxpvNaL/PkBXhDB
UI5etzp4duKI6CiDh1bsSQoPhSzQcGLSw/c9khGbt/ARjs8fdYr6m3qH/Pt9CNqz
GX1jIKcSM0j+IAeguB7sBTIeMAlCT5KNlxxVtG6fN2vWbG+qPMAs3VAnKdyTidoH
46lKP02ClDzZmUsWVSbpepDdupaP8PjQfsJzYi8wwPUqG0cH7P8orJ676hz0sFZf
pp+mtzsoo8djeof0t7b2e0k1tlLzPrNJW+QY8WHhSKwaQTWiZuk+vQoiw3+SODzK
8rjrsksxVGJtj9qQVwuR/zHLvgxmiS/MEnWFGf0O0BmW8rt72jrYv3XKEz8QIJqE
sqZscQMzG0knTts3PcXtYubzhv2Yl8Ht2Scrl4zrr6EzXm0uVH3DEL1bsBKEPn/3
S4V2E5kIucRolHzawakTdITXRLXFlGxhkLcHk9nrhmTw7SlRst7lBxLaY7bB4JsK
qdqQ1xe5LzzqJfJSXHXqFraPpxzttDrD86zsNrcWaPUa/ZIBPz18NOrL1HkYtDbe
/i7d8n5JnUWgKRPQ2T5ZxLNSho5kr9HDn3Yh/oVEc8Ie4m2+YPF1utRsfg/nEhnr
XOyALRHVVItvlLin6IW/Q36iC6jNEaUeEgFr7qtNli6Qkc4iWwxg9JJ6bNmRQ89e
Nc7v9mmmW5Xd2qk/OhQYUwDB58J1Eh6yIrlRXTLu6G1tMlIzOp+/02CeZgtfvswK
FU557QjLnckWyV3g0OyQm68VWcCOGW/x2yw6rOCdmE4I5GtPEQTOKKTT4EYxrFlj
j/uA9WS+BtFSI4r4JPurqwNBofUDKkInZ4w4LaKtFaYVt1W/gHRZ9Wz0kUTNhaE5
sdGIlsY/+zdhGXJ4cTHEjXHxd5D6NGu3SntrFjU9vwMlepnxPoIPulAyjaALUYtJ
gcqijVlSGIySZ4+F87pnOk29aO3i06tbzwLVuEOsliXnDJokIzz5KjyqBlOhBoCl
GYxCPoMz78tqLOF84fa5BTvuEzLqVbF1Bf4c40g6rEWLOKJmcUeWA32AfayhW90g
JEcORl7G8EfkVY7t7fkwHSxg0V7rFmFw5jsRRhHnDhnf6VNswTIS4M1/sXGA1SOE
6b6ygQ5J8fR68cXWSz1GxFw642vWWStL4ivztfxElWtnLSMkioEdvVTnbVC3x9Kk
CTVFe0mtwQ3V4PAsyaKlnkv4lx72onT/7MisFaZqA4X6KMXkyqIN43OlGqSonrI6
nX5YXQbZtN3vXY0q8dWAFct3QdY1dWlDOJnZIAGHel/plVS9u1aF1Idi5bl8fOPx
xqawKWAOgM8tFnAtXrePMFLsqLR+Zu4dXn9EOSwg07ww/wNVJl9OTJN7eMci5zAC
5qAr+MTNw6J+VcyhXY7/Kot+TpzqVcNftVTjVsbiWQYPXECOcCYjZHYAgGuWtOlq
DKX25vra4cl3YKCd7Hh0yaReByV/1crbc3JpVru668DANSAdteGpxYNVtcwZ97EU
NoVwojOOaX2rG6udwHmysCWi7I+TuRblXnf59qf1Ag3FeVCSEvGTtov5McO6cQVu
JosLrRddmht9KOom6CjW0fRJ7bAOtLlB445n8779iTwklB4xenr7sGzPNVFpM1zY
CUezzq+AqOHH0BORlKRdpcME8A2LMQOMafhYtdVmedjSNrbsLjl+H0G5GOZZWf6t
OjEGk2AijGEi4c0nHgW6d47QXiT2qAmHDE2kbjhPQcRwXP1j87fgH7hRq4ROtqWw
O/Hh75bNZvghs59GUJKZq9FIwAjfvlOVuBUH/4i4ZMvLaXMJBLVolQXmAf1bY6J4
OJv9l194YfkvzCuLjooEuh8hPC3NkHcNSU7SDhonTt8Ny+8GqsH1nC8fAN8QwKWv
ZZ3jsWB3reHxEXnE0a6B9IgSvZrs7vKuSQWahx0VVrQHFcV4RszOmcoh+oEc2WUl
2Kw62Ou/Gk6RcsqzB+tTyYewlwsTALpq89tx0hj1/Aov24ezevKh6Bw8Rs6ijFbR
5goQbK5ktilHeG91rBcalEutXgikKhCgzHqnAyrbFbA4ZG0vD/W2ps1tFwneXNLp
e0oWp8/FqtNLYUOG+an0chATlRfrkMlEtg37vQQYOyGUWLbS2WzqWYnjokocMEZL
`protect END_PROTECTED
