`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ni31Wn8+Q2N+CikyqrcmGOzyYcOl0AqlQdU52/g9qm1Cg2T4WEYQag0Pbxd+MbSW
Yz+7+CCefxLPDRXaKwU3f5eVw42VlOT8W4fG1bIxmiggJgjsJrXv0zYjDhT64+CA
PxfvKC3XU8XW19rJ+tYDjkk3gjYn6MCXmQuZ3M51fJIdUyz6aoS59pfhdr/KBLUu
lvgau+CD6xXlknywSOcZpKPyuuz/Q/5mCQbxL9SPaL0o6XnR4qadYZU29ggtcSFo
w7XjqeBOE5oy3PcrwjfIJWo/md4b6iMG2PZvWA7l1DVG9HhhKyTE7iW50cQAOywi
iSx86SXn8B1IESNpTaN2AqLMkZ0HyZ5R3Eoed14b837B+4HpY97+tvTqSNNt4F5p
sAdR5NceulVP2GgDJ3NMtGWIUmep+Hdwx5me5F9EPyoTXNCL4SEB61+2yIdzQ7nn
kIYCEunEixsGBy3r031Kga3gNRFi1GUfnaxz5MXdEDHRhNs8KXCtIQPw/bAKpvVp
BemmTJVd6bywJcUNrmF6e5l+17QbbTQG27uunQwV1NwsfQlAXD53OFlkwxujBAsi
SQdDJV+NC8c500+DAdfucDabWduxZxJV1NnIJLM5q2ARRMudNjhK5mMCykT54GUI
XSb0dCtuBxR+gmxGjelJBF6mu38M0nLEJOSsgt6KSm3sGr++aF59jcQaYBSEOVI4
wBWi091fvvblZhnT5ocDJqqvqHzlIP86EpTHsdJGKnynAcA3xAvBwjmPZASLUFJF
ZB1v0yfngBKbbGu+LUSGXDPwh99jy8X6E6xLTvSF8O3awfs4WFcKkgUFldOVvSHz
UqugJ0E7FBDLbDZc4bvIwP7BqQmVv9MYLbB5KJ3jNZHNJFaPJGExM9yMq/4bE0Nt
paenm9UvSYnXAxd4EpTD/QzuPG5gDEi50sNuu2C9dAG8uMxsOCUqiOuXfbuPD7/N
SgQsR6Pqj2GDbF+50sRNG7xe9c0BJ1D+a6pg4iDqdujSBTskgiPfBKBNNAyjcPwf
BnGhkuOUwho2z7JkK1EkboDLVVvWeJ9gm4m5ckpOF9DzVBblfYbSh/mtPFNZ+7p1
egRhr8WgR54CRZ0F45RfslmXtF1zYmCi7fK4lZeRwsJtV0Ax0WIbvUju1zNxA3pO
/oD5rRaeYNRMBw1uCC8+RdfI/obIydWCkURpsAZg7s4BF8N/uJdUgS5IiZRw3c4v
PWnaQfVx91iC3/bxwu8HuD97EjO2ggiNxdwkQg+ugdof3HLI8Bf9nJEKxyY4FdEh
MQ3eO+1/7KLnpGSSyR9sDMPiS2xS2SGPaansFMEK+zcim/SIzarbJLVkXcTSfWXT
k4/7DNhFfYN7scc3ivl3cbS/WykdH7n+d4xsK7j+u2BaLmo65SczEi/0W73yXP4r
zKVy0kHvVh4AIOn1B6dk3MGnfR3tJ9K3GP00gY+ZxxFO4YpPnm9N2iF3WVJbBfcp
x5hC2YAutQf98gxNBZ1jfg5IUZXYGhUvdBaY8zRqsuRo9831E4kB+PN3Ux8kV+D+
BwQ7qIVKOSJ88sk0am885MOwTELEQ6uo/rMD5s9P01PAY4QHJVzDX1Tt7gjxcga1
R8RBLUbXVGa7DHYSUugkxMlSuLTiff7Q81k1DXYGZwy/5XkQxLs2HpHLuoUxibun
f7SYCDvwVWVyDaWtnXxMD/7zq2CyMV/ROdd6vjKc62QrRtg/gZfJiUbiZzpfedFJ
npFWi2Mtcd+BNIF5o7wxu2eUnPcWMQwNMT8yfPxqfBMRtprvdokSi2MzY5I95VEU
B5QjMDc3/5XATGVMI9pkrmcqAIe8mu6eQAX/f/GXgQcYCvczjcMCNTjl6cCjQPq8
vZEr0sQFjwG9J7ouAeK7Rmf/Lnnpr/CbvCgHnttC2X9W102NdjO3LMYU+dmioT0Z
0jTUL13ILxSrhziYVgRWau0C+BhfKpTVGfWFaHzQTi37kypPr8kRNsDFKiOcp2AN
+Ccc6aSAe+d3BvtnkqoPW5jeBv7fM6oqmZarRErp49IXbRaOyosw9qb5xyQD1Dg5
CFDTdU5wQ0CMPUYaSRMlzrw9YO71XLLLQEdPeidPrxXwiotcGNjqKGxmeSJRuwt5
Dw51tUM+JPZJjmSPqdfSlGp9IJL5HGtLKlQhoQHoruwVoINB9RHRTtF//p9C6isi
d8StlmrEJv47WYgT6IyWL/gNZQAnhOudN+X2lPWUuG+jrkBLQfHSzLYcGep6lqpl
Y9aFZTqh0u02C07Om9rUGIJFqK08apISWIWJrvme+t7QG+ZH2sxLs1/f9aOAf40B
dBqS8Omts86P4qSCcEH33Pl/iJxAbjAVOSlIOd6XpnKFHqkYW/KWVDaSeHFKfsY5
fM1HTBhMTHeB8ceGz8ImBCddCxQRW1aTlVMfoujbMPfZ7SJfCOx7UBYjKJLe7CnI
s34a0IjoClvgPfq89RHwAPYHkTqSxtjGyzxkI2U07nLn0ACcqCNfmm8CkymDRZMn
K2Qaplm7rYXGv7sH2lIp3k6Lf8431N3ueUv3XeOrdQmyqV1wMT7wgH7mA5UX/JEz
rC0eWBvJzWA5/RtpkimpdP6ZAbZkVJOBIGB9KXa5eZd2CUsS/sRqQTuGKgNlRGhI
SA3CI+tc6DHXqBc6C6886smTlRo0+SF9umvt2T+NV+tuNUyhwGcdg0+rwzi1hubu
5oxuSnfi5g4lAyyfffuz2Naguf+6JChzeVSCsY2Yy1/ahsU/3b4zuD2L76eakmRG
NBSi3NfTOUVSlnSHAkpFPZNp+d/HRS1i84emN5nDH4wDle9+BGPinlLbeoSY2dF1
zuMZ6qAn3sjXzw3I/SVgnY3S6eQ4j29nrrgYHR7ISjIH5BRsxUP6ZJLhOfR3TYda
v3maAJd0QQulbIaeMrBGS8HPvqxGWBC2LjGnwJcNNiLDUznZM2ip8FVjeRfbmMFC
AjgyYYvlv6M0Hl20+3KYtyeIZbj1b8QQdkKUOYjOSP/Y0fx0InhEE0G/e7GFX9HC
B1nwN2Aah4D8P/TXPKXB1xU1iy7EOeFyX9E1d5O1zqFh3yo/tsXqbgiFTn3ZC2/c
IwlCG5QMNH+dUaBl5YxIy0fR9wiaJKr/jzc5E6xnvjni4hIxdEdnKGAUoG4CIOTT
8fToJGyz9h2MKgYdj8wVWHjgCifDRyv9yCv3jXaj7R0w+zuk0UiXYtx8AOEZKEZR
/TnqMoln+Rb0A7WgyiRTsUIhQ5LMmexRPFY6bn5tHV8xXqDqzYtuhv1mvoJKNp68
fD38uCVmLIyNCUtXP6HtzGNF0svyrEcnPmGu323P1qTWIdZjEe4FzmdrxD7ejsM2
NQRYo+AjC1kIsMoIpOraHaNplnOCJwy0417M5tw6bD+dw9QkLS1KHeQzRYSggBCO
8GXvfB3bqXd8+NawtFPd6TSjg7DnE4Xph3P7Xx+O6/AQCAXw3lvWnRT48nnjt7jp
I3HwlJSU6vFFDa2+gCE6/xLql3Z2YtEPg4PSjYLLgJgZdsqDgQ7cvvSN917BXDCk
oF0IdOSAZVTC6txrx04hJZzTA9rCgBbjIQXOT20pDSemI+wFinzzDt3dlaM0FlEF
0Se4bdgj+TeXmeAYxyA4TfvQPZexpmrdSku0a43f+k6VifL1uuc5hyOVcV/tuE5K
KNxePWog93brANtsT565UZB3wCiQR2Q4RhAyPl+dMa/1phB3M3cBIyXhCrzhFn1s
ukpOcbqypfAFrEmkdCKJ1oHYNFNEU/FqjEAT3mXHU/NuZYcM1Kh74GNyVN6B9JBG
AovahsiJj8CGFC3jVO1cjj9xrMbUSJ10nFbkz7jQVMwaYsPbi+qbhmpDw9rQo8Ce
3uVkJdzRBR2wozTe64A8bKHZ7BReq3dSf5EX5iMLWqNsrRt0ZC60kTYFrcFobXhw
CiOdhYeIgR6/x4SncUG9VXy7bcQWhRhVEhK7y7R1dlZUCercIWQyMbBPxxqAIUdS
ueygYUIavVFjr3K10CES4uyMstiZse9VI0QJMAmRa0uZGdcsu9wjB+Q2HA4niGxM
c2XHCVCuP/s3Nuc0O/9wdcBwJUdJfzJyfs1t5M04bWrDGhwxL1fH0OXijtxbnnxO
`protect END_PROTECTED
