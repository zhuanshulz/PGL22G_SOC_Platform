`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNQzYZ3RbDEWEwI985zmRDfP6CO+ywchOOHs8G015+ZvBGTRiDAKLranowJAvn6k
M49yOX/MABx/GGZ5RzcL3ZbYE+5gI8U1+7g8uOSzc7vQ0PI0OOi4lHK8JIK7U19g
28o5EgiDYHonQy08l0QeU1VH0UtqVwBhia/nSPYN5laqf3S5CmRX2VOgtX8QeQKh
OsTZS1QgV/rdWw+Vk9Z14U8zfVwltbGVEkM/hTnjbUe3/FrRwOrQgzpMqlF0ayKJ
aSUefHKfeI3npwH8Mit614D6p3iI7h+fZvOOFP0qYRZMedpxK8iGdiW29K1i5kIp
9zz0WNWLkQjwQ+9d2wZoRrZJa44/XbIo/axz9pF5skWLnR+ieaBj+FZJLAkhOMc9
QxSful92vPhQKiyauHIZcA==
`protect END_PROTECTED
