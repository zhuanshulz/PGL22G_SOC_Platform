`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8sPOtLaXou7HnAE5dPfk8cRGdMgL2RwjYv/vWa8g6saWtKwcwlGfdXkiT51IkFrY
7W+Ta6bxFgXlakcMwFLluvqqKKZEJLuTak3w7RPKNztOhCFQbB/rG8vwvCim5uLv
dIkmVXUzgWh96/v2RO1d5FZXXuMOHs0uRmAUj3L1AD6LNzCIndg8vxAMBT5miAwZ
ooY/gYGIOtX+oH05bl+WajwmIjHEIiVsItR7bq4Zw57LFXXA1tABBhch9mHJ79XP
MiJaqmIhegKiWhzKAyw18XbdY6orO3UcgASkK0T9Sh3lRZ94zW+t4d4jcgxS3VY6
GPY/v8L++V6ypa0G9aFtfLCMSDOgn89zysAZVz/QJf7eSJ55JnCPndsOcaRymZb4
70x4oDXW1Rj2+vfJBmEsnl7zy7hURtgHLkmd7zjejAOwj0/ATJgYIOrOG1B20nhA
6ZOkOslY3bR6j+9Mvopq26Sf8eeOKDpRXS9Tii2bQlEx4tRM6FEizI/xuTtWOGpg
5HJFuYFfj0NhwLu2Gz0fxdeqO1YFrvAKw2LS464e5V4QZTlHfNjEutj8bDRWJTxt
iUuWJ20Gl0U0zYa0UppRyj8Oh/KIN0MTbhEBkaDWp5zX997QaVdttSMowm9/x0/o
mN9i72JE39SQjNe3sNlKmWYrtgoxRXayF4UQzpel85y069Tgy3osHHRRSYTA/gvo
qvYXjnjbA0Ce67LDl5IiUWlVbhOet0eDSYu6Z4yOblkj6SF/E+6Ip+w/ILyZ17GW
BNSN1gHKynXFj0SuaTQTrSle2LiD17nQyWvFHe1NeZ/SJqT1dy89waKqbMyw787T
NgY4ref4g+KOtEmvvn3Yr0+DTQCvIeQf4McfNvD7dGY0IUcy1JrSwLklrdPDGCXs
73pbuUVsLFCaMrk1md7ezA2AmkuBFJjx0cmy438ub/U0FxAHHZt5czOxje52fg97
`protect END_PROTECTED
