`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f7FwuVpHDkuO568HC4HAhZoggSBg2UTEyez2xV4umSvG2nw7/uMzEi1Jb/U/adzh
RmJydf+ZwR0kqMUmxxiKf2dOhZDzD5qcsG1lVquKlwYg8fStYytOYChk5z+Fr0DB
2gCqmczxquyOfq//iVLNrazRUrelIAm4zeHHtHfR7ukPe6Zws16iNocKiq8qryfg
K5jBe0IDKIHIBDmODDT7dTXWNoChfJCjbpl7XHEGkuzCkjbR3Ci34m6S03zwuqB5
7a901Ul5TWpHsHBhCMTAwl6VmS+GNAcuIVFfDH24KBYqSnu8EqrRwHiYGqHP9lj/
EJAHCN8G0D+Yn+/UO2P/PLXufhGu3F14V/ILgPvz2Mt4wM2/mwZ9ExheNh0OBPk/
a404S3kusN43iTbMbmUNJuFn7iGKG28O0VsZh76ZQKPzPnEtA7DuOuVeyCJs3N87
u4XD/urS5w/Lwhj9v9c94dmQdpfWhcTyjOGfa0wANQJq/3HJClSs9BvpXRgpnK6c
YALtkEKsgjkab2kOrDnMkqxhhwsohRzR6FBhocZLyvZ8sELUOBNnxg1b6Vs4EfDm
rz4OySzrwH6Bs9yqVvX92NFzOwkCIPcW+3WWeRTYbK8Dj50FF3Z/y72kMFovFMD6
D3foxt8kgLQ073Ttrz4qUMqQ+iXUoosfq/P4PAW809hi6GAKciO0fEYMzdopG8dg
Kxdvpx8yMKXZW51trt1XXEo/YcMtGGdsu3k+NjCS4ZBIvZ9M7hKk/zXpuJ/8QA3D
o9zrGHFSv8caJfNBRF1yQ8dbBwkz7ewOUs5ffPVQMf3zEtH9+BCUo+n38hyhMT0m
BSAcSAbeH3bOD4QXsmVCaO/ubOdDatWyUc5KUjPaUXxZ2D3QSEU4mt3CEF/yAzqF
DY8Z77CdpQxzGYAGQxBIm6W/aYPtD4S7viOzgTI2GfKlKBIsRo1XpcciCFM26r0X
6lVq7fS5RJM74DMu/Kz5GW84MyWZcj9MHrxf5zvdOQF6ftvirNdZehoDR/IkNb6j
FO8u566p6dJOrIPOn8o20k9CjwBHGwDhVtyPjpW7VyQux/zeM4ENPdj5P7gUYY7W
GAJz2wAGzudM9imWyrOKdoAng1zG1LpiNorCZoS9jcLdrTq3L0mjtr3KxOk8OyXj
vmtJOog210WRlBajjy+pGj9A7ygKlLlGSWo8SeTRhNhj/iF8J/5iT4vSAqWM/ewL
8XOcXk56/nJVcCv5SrTrz5Xc8HAIOKN/62pzqXmoX16tNicllmst64gJTrDRnbKT
DQ8/KrpkOIerSkuEIjbvy8yzlCiAE5HmpIUSjciP2bCeoZ11zCiKS9MBgAJRy0B5
5Fd2z3qmdJsTQmmI16HPGkpr4tdF5sg6aQwfwZWMxv/ishWxpP2fH/s16hIJjSvF
Qzdcv6SKidqQiP5d03kpnW4DSrOgGtNki5Lvu9YivjoRcjTPUnKlSqNEF56WdxQ2
KiG1rlr0kBMszmEed4gzp6mWHegj9+RN9A9/LWI0F5T32gi6a+j47UnBmiXTuAac
nx62xQsDFb+xBvLcvSLeRk9ZZ6/JkgNmeYru0jT15roMz/LhBw7mVAU7eclbPhyb
nKdC7Bx8bxe9u5M2IJPsYFKHMC6wbq4WJrs4YRgyoIedhl940O5DgShnt/fpAbHQ
iWD13E+aysp2bCIhRJLDXF3D9C4nHWAIKGs1IQx+PbmEQtSvQUkskl2Of3RCxfyN
O7gMrKxEk0fXKDrL4z5qIhFxb8dQZIlQEfuNFmofA64Mbl0xRgxzVURYPLSGmcBX
KsyROLzNDhgbGh5AKGwE05QxyT3yyneGt7lq+c/xjkaaNDPeawJO15dxttB7Qni5
E2ispoXiM2tjmG76xqCR+9mVhJCi7tGbvoQXk7Zv1sAJrMhROMtIgHs99/+RFXqm
6WQG1UXSNXRnEvv73sF2N3R3mW7WSmtVAziwEjJ7sPXDHIQTNhekWHiEZGGfwMOu
BiQLjhJJ58jdP/9H2fqiDE89zrc1RQ3ktTy9abiYPs/jZA/0cpnomwRnVYvdDF6J
7QdwRjzeaCbqnShNJflSmlVzStyk9LKJN6twAHRbYrGHDvyEmuJHqGfIzK62c8ja
8y8ryzebpCsMrDhxxIIQS6xdozTMEJOGJ2kcqJqZC+AxVTgGbTjaa+FPgOLnZWho
lifzg0o66WaRVnF8U9aodEF2rHaRb37TEJBQgOid3tChwFjDvMaPmyS7U3CGGio4
etQx/3KWVevClQx1wAawXu7Ob/wLfQh9kPadcckb7QrDF2RgRf7dHbbp9x/T0PWt
pN992ysD3doQ4sNNGtF6JDdiNznNL189OWR/wyOIFTXpwNNAL73HROVkFD3aLA2d
IsZ2ygKUZDBHaIZXqIzIl08iVbm4AjV5FTJmpvqHKKMcFREqmKUYKrYBTuwjXPkZ
gT/XDHn9hmDY5uSNon0E9EHNJ+NrQc3sPeRZr5oht76z5UB+tSLII8hDc5eeqy/P
qEJi0xWboLviyvBvLvLfSH+szBPcQNR5/xxKpO8q5DwcVavIqhpRUl7Askq15IpV
yYrjI2HZMJlI5wDIpsT/plDKMMstx/5D5YGSx1+jiZ7oISS/RNZkW318y8NegUOo
YIjbawT53XCRLk2XLhjuAEnldqcCy0UR/ivmQlV6yZQBjaLCw0tdvGwuvCvdNTii
QS42IC5dP++88RHmC6cQVxoHEBkk17WkgDLU67YZoi5a6o9d3Zo52EciMwoOlTWj
Fm0xKv6PS9fyuYHkHmuaveMsB3f8MINwZwYboA88cz3uQKKJnSGk1pKw5nEY//8Z
tz4ZLrdn0kU1jGVQayb6KmVdLGwnV8m8uClsl/a2kFd/24eGSjqQSCgYRw34NYRF
`protect END_PROTECTED
