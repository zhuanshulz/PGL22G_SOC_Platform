`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YqUf1RPF/sX1vNnc2KEIs4KmtVoxybDSbfKVLA0Zq51svqcUtZiZgQJ3MIPYdpZs
vlEpOCX24U4PIsiSq9N1hjKdWmuBYzBLfdU5uFwCvQC6gavo83BOOE9SmSlvwXvq
02FXHBiesffnZ4hv2o9ohAPA0a8NZO8bRuSvUOTlUGQT93H/PnkyEIYHNlJdLZCk
9NoBjV7beGJKljAKRG5FPfZTP0kiEjZy+YLBLrRdmDHnABPkDolLVjmJoxLoShze
gQuJmgWo60xGEFi5GRIMedrzIUshp7uDjJukhtWFA01bHXMR6pxgC/F9tUkQ3Haf
PJ0E9/TA/NQUSYReBBqkXjJuSoF6Mgqe96xoXcZRJ/V8dxgP1Ia4x31AO8qamrpo
skOybeeLb4mw6AmCc44L0g==
`protect END_PROTECTED
