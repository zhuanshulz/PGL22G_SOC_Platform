`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ua2qNsD+SFV9QyFFqiv9BdgT9XzKRgVm7CAZLdT396nMqtVUWoRVj7jE7ygCleG
Yy1xw0mjMgf9CMTxhQAo9uMcZ2a9Otxod/KY6BBgbtfsCb8IqI5AXDBXMlw67/C+
FNJOrX5Q9mnzrD3HBRjOzajppKyAX3HElSr9fWklKF1WnBBmRvWHQAMDCr2+lnC0
Wij/s755JH7w5SINgXgLV6+YeKak2p+94z8jJYFm4d36z1t74fgryap+rP5JCtjl
DZ5zZQiG92ONU0SreCip/iFv+3+JNchR68lPRl+akT7i+FF3OKT2xmrICj29Iizt
h48lvk/iAM2AWvllrCuYLOIEfv0q70qLrf4R5zvNScBRgsQK5Y4RDtsMx8PvpEca
G3vXg3BL9h7Z7yAgB8PvcIuzVzq5PCdtTwZIvBfBGacOIRbCcNi5gS/E1M8UeplV
jAWKtYUUL+/6tlQFLtFSfOfyK/R358NCOWV5TXtyvswI57XDukH4W/psS1TEeK3/
+ujgb2aCuPGygHqevPAe1t98R1663rFIM0AIEKIkuxAC+qUA400D0VgG9ludqMxo
tMLKsRUg4qme076YYKXXQLmgP7OSbSfnBs7VszbVlnZxit/2/jBM5tAlNSp8JAcS
`protect END_PROTECTED
