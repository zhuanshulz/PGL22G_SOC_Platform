library verilog;
use verilog.vl_types.all;
entity APM_H_UNIT_INPUT is
    generic(
        CLK_IR          : vl_logic_vector(27 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CE_IR           : vl_logic_vector(27 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RST_IR          : vl_logic_vector(27 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SYNC_IR         : vl_logic_vector(13 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        IR_BYP          : vl_logic_vector(13 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        OPCD_BYP        : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CONST_IA0       : vl_logic_vector(18 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CONST_IA1       : vl_logic_vector(18 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SOURCEA         : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        SOURCEB         : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        SOURCEC         : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        IRDSEL_B        : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        IRDSEL_C        : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        DBYP_C          : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        DXIA_SIGNED_POL : vl_logic := Hi0;
        DYIA_SIGNED_POL : vl_logic := Hi0;
        DZIA_SIGNED_POL : vl_logic := Hi0;
        DXIB_SIGNED_POL : vl_logic := Hi0;
        DYIB_SIGNED_POL : vl_logic := Hi0;
        DZIB_SIGNED_POL : vl_logic := Hi0;
        OP_PRAD_A_POL   : vl_logic := Hi0;
        OP_PRAD_B_POL   : vl_logic := Hi0;
        OPCD            : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        OPCD_DYN_SEL    : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        OPCD_DYN_POL    : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_CTIR        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CE_CTIR         : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RST_CTIR        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SYNC_CTIR       : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        CTRL_IRBYP      : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        IRSHF_B_SEL     : vl_logic := Hi0;
        CYSIGNED_SEL    : vl_logic := Hi0;
        IRSHF_C_SEL     : vl_logic := Hi0;
        CZSIGNED_SEL    : vl_logic := Hi0;
        SIGNED_ENA      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        SIGNED_ENB      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        SIGNED_ENC      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        DXIA_PSE        : vl_logic_vector(0 to 16) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DYIA_PSE        : vl_logic_vector(0 to 16) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DZIA_PSE        : integer := 0;
        DXIB_PSE        : vl_logic_vector(0 to 16) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DYIB_PSE        : vl_logic_vector(0 to 16) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DZIB_PSE        : vl_logic_vector(0 to 30) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        GRS             : in     vl_logic;
        CLK             : in     vl_logic_vector(3 downto 0);
        CE              : in     vl_logic_vector(3 downto 0);
        RST             : in     vl_logic_vector(3 downto 0);
        DZIB            : in     vl_logic_vector(31 downto 0);
        DZIB_SIGNED     : in     vl_logic;
        DYIB            : in     vl_logic_vector(17 downto 0);
        DYIB_SIGNED     : in     vl_logic;
        DXIB            : in     vl_logic_vector(17 downto 0);
        DXIB_SIGNED     : in     vl_logic;
        DZIA            : in     vl_logic_vector(31 downto 0);
        DZIA_SIGNED     : in     vl_logic;
        DYIA            : in     vl_logic_vector(17 downto 0);
        DYIA_SIGNED     : in     vl_logic;
        DXIA            : in     vl_logic_vector(17 downto 0);
        DXIA_SIGNED     : in     vl_logic;
        APM_OP_IR       : in     vl_logic_vector(8 downto 0);
        APM_OP_PRAD     : in     vl_logic_vector(1 downto 0);
        APM_OP_POST     : in     vl_logic_vector(10 downto 0);
        CZI             : in     vl_logic_vector(26 downto 0);
        CZI_SIGNED      : in     vl_logic;
        CYI             : in     vl_logic_vector(26 downto 0);
        CYI_SIGNED      : in     vl_logic;
        CYO             : out    vl_logic_vector(26 downto 0);
        CYO_SIGNED      : out    vl_logic;
        CZO             : out    vl_logic_vector(26 downto 0);
        CZO_SIGNED      : out    vl_logic;
        xa              : out    vl_logic_vector(17 downto 0);
        xa_signed       : out    vl_logic;
        xb              : out    vl_logic_vector(17 downto 0);
        xb_signed       : out    vl_logic;
        zb              : out    vl_logic_vector(17 downto 0);
        zb_signed       : out    vl_logic;
        ya              : out    vl_logic_vector(17 downto 0);
        ya_signed       : out    vl_logic;
        yb              : out    vl_logic_vector(17 downto 0);
        yb_signed       : out    vl_logic;
        za              : out    vl_logic_vector(17 downto 0);
        za_signed       : out    vl_logic;
        prad_op         : out    vl_logic_vector(1 downto 0);
        post_op         : out    vl_logic_vector(10 downto 0);
        zia_post        : out    vl_logic_vector(35 downto 0);
        zib_post        : out    vl_logic_vector(35 downto 0);
        zic_post        : out    vl_logic_vector(63 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CLK_IR : constant is 2;
    attribute mti_svvh_generic_type of CE_IR : constant is 2;
    attribute mti_svvh_generic_type of RST_IR : constant is 2;
    attribute mti_svvh_generic_type of SYNC_IR : constant is 2;
    attribute mti_svvh_generic_type of IR_BYP : constant is 2;
    attribute mti_svvh_generic_type of OPCD_BYP : constant is 2;
    attribute mti_svvh_generic_type of CONST_IA0 : constant is 2;
    attribute mti_svvh_generic_type of CONST_IA1 : constant is 2;
    attribute mti_svvh_generic_type of SOURCEA : constant is 2;
    attribute mti_svvh_generic_type of SOURCEB : constant is 2;
    attribute mti_svvh_generic_type of SOURCEC : constant is 2;
    attribute mti_svvh_generic_type of IRDSEL_B : constant is 2;
    attribute mti_svvh_generic_type of IRDSEL_C : constant is 2;
    attribute mti_svvh_generic_type of DBYP_C : constant is 2;
    attribute mti_svvh_generic_type of DXIA_SIGNED_POL : constant is 1;
    attribute mti_svvh_generic_type of DYIA_SIGNED_POL : constant is 1;
    attribute mti_svvh_generic_type of DZIA_SIGNED_POL : constant is 1;
    attribute mti_svvh_generic_type of DXIB_SIGNED_POL : constant is 1;
    attribute mti_svvh_generic_type of DYIB_SIGNED_POL : constant is 1;
    attribute mti_svvh_generic_type of DZIB_SIGNED_POL : constant is 1;
    attribute mti_svvh_generic_type of OP_PRAD_A_POL : constant is 1;
    attribute mti_svvh_generic_type of OP_PRAD_B_POL : constant is 1;
    attribute mti_svvh_generic_type of OPCD : constant is 2;
    attribute mti_svvh_generic_type of OPCD_DYN_SEL : constant is 2;
    attribute mti_svvh_generic_type of OPCD_DYN_POL : constant is 2;
    attribute mti_svvh_generic_type of CLK_CTIR : constant is 2;
    attribute mti_svvh_generic_type of CE_CTIR : constant is 2;
    attribute mti_svvh_generic_type of RST_CTIR : constant is 2;
    attribute mti_svvh_generic_type of SYNC_CTIR : constant is 2;
    attribute mti_svvh_generic_type of CTRL_IRBYP : constant is 2;
    attribute mti_svvh_generic_type of IRSHF_B_SEL : constant is 1;
    attribute mti_svvh_generic_type of CYSIGNED_SEL : constant is 1;
    attribute mti_svvh_generic_type of IRSHF_C_SEL : constant is 1;
    attribute mti_svvh_generic_type of CZSIGNED_SEL : constant is 1;
    attribute mti_svvh_generic_type of SIGNED_ENA : constant is 1;
    attribute mti_svvh_generic_type of SIGNED_ENB : constant is 1;
    attribute mti_svvh_generic_type of SIGNED_ENC : constant is 1;
    attribute mti_svvh_generic_type of DXIA_PSE : constant is 1;
    attribute mti_svvh_generic_type of DYIA_PSE : constant is 1;
    attribute mti_svvh_generic_type of DZIA_PSE : constant is 1;
    attribute mti_svvh_generic_type of DXIB_PSE : constant is 1;
    attribute mti_svvh_generic_type of DYIB_PSE : constant is 1;
    attribute mti_svvh_generic_type of DZIB_PSE : constant is 1;
end APM_H_UNIT_INPUT;
