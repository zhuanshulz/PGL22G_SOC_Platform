`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HulHaG8uu8X0r+GJogXbqqkPYtYoeTqrbeP2KUTQ83MxnJHUx+GW+eHgKFYW4kaq
WVdYfUSx2bvDStDxAjR5M3uHg7/Pv7RkiPo0/p1zyZe6tgfHMLggGHjnd0NX0mS+
jVJ1ZRytNXFcaKF28SofzDM4N9ismnUnnydhMRDycNYcTklDdsGCjzWbTbSotR9F
7Xooidd+dbNaboB71ijVurO7rl8dj4NtHDrJDwPpwQ6fHvdeh7+59QOznbHbgec0
uVnApTBijlj6GS1aBX68YHRG6Y2xi5jdgJczCGWXsvBbHu6nblDHnpQJzwkIQRLL
jGIKV8Rrko7jAtPWKQYRq+ymXvanpD5XXkTVe7wbtQ8NbhWY7Kg3ztFOSS30BT3k
0gqhfA3jQ+dC4zc8DbzOvUWoEusDO4J1cKHF0FMpVbnZS+uI4VyXDsXf01gTcJpm
Gm5YIo03Hs0wB0dDOl0hAMfZlfjnDBX3jR2GORvw6iNgICZGNgmzvN5evmo/Sv5e
Kov4sX7KSw0FgvYlPd1sB4dF1QtXZQljDG5Fb6bQQGk1gLfljvjhDn7NlTcQ/w2s
sYaey16Px0m5d0aqiRS6UCfOeQ82a5D7qRH9XDj6owWlEal/0BjGg9u9w8WKtwTh
cEP9P06tr9h8t3/RUdRSWm1JWA4Af8oKS9v7dEnr7NpTbF5FO3pfFG6BCEXH8y/G
b8G8XQ0NC661ZZdRfAkI/GL5B9DLVkSKRyWyO8lrXHRdNSDwaWjuhJBw5q/Z3wCj
Tk7f4ij3DnEpmIFj72awIvhhNpZHNlJPZVfqRMwmAE8x2dAozfa26aRjtuPjZ3tO
5/4b18xn5MC4HnikKa5LhSoXx3ub8FrLKuURrzf3urzmXWKvawfxgapq0u6+J5kx
HN9Y8N1Qz/5FwaR5/U5zmayu4ribwy4hMXjrSfZOqU7S2V3bSKCMHjG6w4U1AhMU
b15AqVhL6iBoBUloeaYisHf0juORA2ScnsaJdLNlPvw8qVDHgd2oxE/Zkzjp2qHs
uV9OsTqz3iEB5Xl4Ezywb8Olx7Zm92IjmwdUVzdeyEbhMZ3P+RTYr5whujZHacmS
gWn+6rU7OHAcDq77bUrS5I27OkU+xN5+QA9eW9MqLAAGsDCw3tMAJXLgLMb+GYM7
QCo3lktXnlCMHqHlDoT5WA==
`protect END_PROTECTED
