`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxpLhE2YT2kFikJi+AHVE3286I6QSIy1Um9kIoshbS/qURfKP5XtDwEVxzQtI+jG
EnChk1E/uw1lLyz+jrT8roSmBgux8AhYLmLxmWR3BMpl2ObQv2Z6GHax7zggT6yX
i4q93g838+VAFUAvwxnR9RmQstbTEcm5ILtSNxQ5VkscL5D8KQdE7eEpna4Y94RD
SBm5IYPNMiaKzYIHjhWf1TXJe8fFGy1l+y3XnhdudJ0YwDu5nst/X5/rAbggfwtY
/HkckJGuYMn2eV1gnGgnn1NSRlmMwgwtvrxne4f75vHjYTDzPS4RM1aHsJ2GlS0J
biM26XYADoW+FsLskpH3DSayohdhsf7f6hkCXCfWayIP9jPHYhBce/AZAN716YOd
sKMgLmwZ8g6xIiZX04Tb+cOIWk2GQ3pStfx5LfLGqJI7/bMMAhiNSQxX97UFvYYG
3GjMzkOf/Y40RkgZp8w8dNcSCzm0ul554haU5gClbVosStYRL6PpsycwbSxLRC3U
QSvNvIGC5mKoHhUvS8hdMNtZvRACkZ9IgZG3lebSBgHNMtYfH+g7owDBvDjHIJjr
SXoHLtRY8fYlf6iAPgeTYA==
`protect END_PROTECTED
