`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iulda4VSYevvuQkZisSh748dUdBHKGf71YLHspFwWyt0kISfuOPddJpSjWsHEn8N
WBp2Co90DkdZb7NQJEQm/FaPjbQ00+T/Cf6BieuAnpmMLxIkPSGyuLo0OcF64yGV
9mRxkC1t7j+G5fDfYk6moA3tabQcJX+p6OkyvIgfQ/oiDBznw5fxX8DBEt9lXKHT
ZS4Y+F18kHlkiCaKMIENBDx940MxqW6MDkNMkM7Do8SL2eKoRnkKeRHe1+9bZcVk
Lm3eQ/l5MuM/RSodTdXpeMIW8r9dNN4of4g/353pC7l8kXpL4YLnnSGIlTSlpmG3
abPZ2bsYTwVLwFcdicKwsB/pF4bXb+MKyC7apEGWLCREMOJdCcLkn8lTNlCdZ8OR
`protect END_PROTECTED
