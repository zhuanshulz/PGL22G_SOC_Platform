`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7LUSXyNJQJdWyM0WZTMPoGVy3r2fbl3ZnQkuWGvC/0CQvOdz1mGJtllmJba5QF15
bzkxB+T+VcX5H/rRLVXSc5B0CmwlERCIiWFjs8GQiMk/OVENnq2kYAkvH+g/yXZn
bwCXA4O3Typ4upn07yHRbi+zeDpF6eZ3d7FTX3AX+qdpzGGhxKe+i1LU4j0DE7eW
mhZD/jN7hhakwOEozSjFHPdO10GC+GBCEKpferGQJ9AxajcQrlEoiKQR9tXY/rTG
6rnvvdhReDEf1M9kPpqG6cuMV3p3jENH/ltOQtl6WrKn1M67rNPEK1dY5umCPYsb
njLFULhylrRMIFyOgvaYLVyrLz6kOmFzW4ytmjXRf5o=
`protect END_PROTECTED
