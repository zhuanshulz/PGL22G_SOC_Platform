`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r/zuGRykUW+jR379k82xQJmx9F4Tz0TZwXT7BOvp0ohPMDMGwiA6v1+Dj7h4jOyC
EANHvw6x1xdve1VejUZ0zotSHJ5cWix8Emhstlr5Ukd0mpwF4eYrkFgSTTDEbbTb
N9MG+cA2dKQ19LjEo1B92zeE/SRm7c2OZmhM4kXgfcLI+NCWfH8YQwqO0PufnsnU
as3uM3qzCGy9TSX0ZZDJyLm2T4WabExCE6xjXfIf3htvdn89LYB/fY1wdLrac0T5
NXX8Q79QFgfikp9r59yeLWUXlBlCNfPHbcnhvdHyTOkteC/2HN8J6f/42Mcg6tjH
bvzJDZwxyPP/GRUBynjg8Mked6AkkIiBxUJB3avk7rsj71jXkNlyJ2JoI1inVrXm
6mP9Eu++TA6NJPu/RK8bX1aYWadVdVekG4Co/NdgIko5TS4oiIAoF/AeGJ+KJ20j
gdkOpEo4Tw8vlbBSrxpVYHYoFZEib8+gm+CoKM3rhnNd82rNxtRa1L9nc1IvnagO
ap4YCoRMZXaKnAq9a5a+36+VJMTrl0HJ1tOtdkDQLCEv+MgCKx5nV4vg5vrszieE
w/NZDpFbyHOV506IY5awCslcmABasbq6lmTKpZr4ms6WlKv3oLZAkLaSBiP4Hll+
2P3dlSTk2cijTT/NRnjLK/PdaFPYctIz6hCcTO8csSMz18tNyU4Uqy+G6MLL6QFS
EmZ43ERtbpVOPRXvjS+b2w==
`protect END_PROTECTED
