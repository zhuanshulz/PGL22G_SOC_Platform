`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9xQv/nbhEgbu4vzwtYFuNKYCQmnkFFY6+k0snp2avPAMkIAlvbumfrf6xwZ+ofM
TMX5/8GquFIojyL6xpQbzl9+Ucag35vjF7ti6Zraoz01uaAs+4KS7MF2pgvyk+/4
AUBhXxOLzguIEPLgP0Oz97GB5AUiwLr7May6llMmOO7R4q06Q89sw8qa9ZOok1+X
LSN450SjoPldkY3WjdUhUwupPeaUMMIR2EYRnQX+fcUSuX5lVcIAqFlgA2OpsDX8
KOD+QmhOaufRd8VRp5rSaV73vsH6jOrhpfZl+s7GJaQrjBvhU8apZy9sS+fsjSob
utLYwgr2RClGpI44HcBFmuxwG2i+TxCJ0piqEPzM/pu7FeK5hGGpfeRuC77WKqj+
ZouXk882p9CE2OkEeNL8mKiOZfIU9n2ggJ2p0NpyrVzAp/2XC64mgwv7NP1U31F9
6GifyeoHET8wBCQbC2/DpwUXYKGWnUWcFdyDEZJ7MoBVRfSHuAN7LulwH9OvzlyX
86/nLbyTeLrw2b/TAld1dxbF9l370OXwLAsch3TaKFUq82ZK2QLOiwSlu8ORW3Gn
T17grFKK8XsGC9xWgKwHDkURPioTAm8ezhoUkcha92UCGFvqrAIx+xwPNUEJZrn5
KR9DgV96Gf+fepV5QZEcKQxlfoY71i2tbObW6kOXyFn/+jA1gyiLTt7iur7CXrz1
WqgaprGrvLBsqybgq1qm/Uu48lxmrtBxD/faCHqzR4XKFDn/jwaLKANH3WIVOqIZ
OrioKcZj8wkbkzcmN3Hl9uq824Mm2G93KxCYFJFN2gAlcBVQ0Bt/Rws491MnD7xN
4S8boVMrHPj3ZNO9dMoi40AFx2e1mTHtveixFsdbUHI=
`protect END_PROTECTED
