`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yak9LvFzI4JKQbLts6VW/uA/AIX6q4N4sRTRnA/Ssd6hdOszJ4rq0PFfrT/a4L2P
+4ojY15d3RXkoFk8nCjXv9zfhBmk0nQw9vl+HrZC4f5TOJ+6FZLoFDuYG8R0cBUC
lFl1sklhvh2N7tHsJ2YstMtSkc8W5+CIahmJpqJ0pNPAHhbT/PgdkTB5iMLsln6p
tLYwpRSnm8OI1uRYsZpO+rD1wdcmk3GYSUsK3TUFrqRehPBCeeFPaUHhAi+mbdEa
d57cp4WDseI3cLvdmKjwJJkmb1/kt+4Xg0rnT7s4e/W+hhMexeVMbktFqAktOBxr
O+iJWyLcn+8ef7OPqXDrQtLGRABUzVBJPVsMe62fJQCp1H6mJ/Pv+nbnngv60f92
HGMS+oFM5s+qyVm1bCsiLYj4rGbm/E3WVwjy0uDG9UZGxsbdUc4PqQcOQwG9stTb
fxZNz8t2li5t6NjRxL+YSFefRZNV477ZbxqpDixH6o3YpcDLzy1/6FNWHBS0MewK
fV0tlthr/PmimRSxXPOC47/Lb9CGMHBS3Z5Xh1ak5YzGVBRuJ1mn2kofntIx6OyR
+nRHCIle+qrBhvrFyQarP2zna8lZpT+WodzRmzRe98S/l8LeoFOzk/PdpP4w1Psb
vMvTA2buM6RoHWUm2Dag2e73/H2ByleM4FEa8G7G47PTvXNW991j8q/oc7efdQRh
iLZyWteZscXBehtrAlWiwZCx7ZDEOTwC4MmncCgK4/oSTy3QOrXRQ7gjwiOsesfs
s8ow7tDO54jo6hQ0T5d3N/t0uINGurXO4KUnMwBGB+L2R1w+93+mQlaYw/Yruiee
dSzJnOkRxHmbnLFQWx39HcHIke3zqWt4yFB+Sq/YCKSbkhBooQx8cg16K/e1yLie
pLjYfPVpkQFXGFaqMEb8G4q7b4xK6t4vpOilFcoAZzKUhlckgkVPcEE8Erc8x4Ym
YCiqEw4pBWYUTMVy/zOIAWwpY6FTg+J+zulfOkE3IdfvPwjh5PvGD5ySykXdECHp
cJOLsHG4armQaYcCEpk+nxruBHGD8gAFCex8pk+WrJxedK6SDDC0g+5wUBGHhtML
fgHUzlwaVU1E/lclTuhwD0/UVBwlZdclCqzqfz4JzIha1i8RdCLRuJLOEqsKzcc3
vwb9fi410qv6EjRZ6G2SgAmiKy0qB/c6LAFSwVH7cxq9Cve0Cdtxj4S4OAO7yWSY
7QBUgfEXeSOesp0dlsLVa7TQePPyyhHk094u/hs+yu7b5G4NNuKhlMGLYIsqnLCk
gQF9US2hFwxpDEOfVt5F0L6jcvuaZ7eg9xwatxE86QtzA4uHHaq0eOpbW5XOtijm
aMotv+h/97joA/5a15WDwIo/bO9RlYrhoFGpspamOl6bbBwU+3nYOX6kaJmRYN51
afGl0+wdnVG9Q9KNZPzX5OE0RwK9bdz/iHb/q2Vakao/09Bt6zLA8Z63idlicHIg
R8I6MFbctsj+izp69dS+yrvqkpIVq0gkNn0EFlhma+VJ+2VNwmPjAl/q8yLj93kd
AHC5vFeIXE42fRWEOQqC2yUtRYyPY8+yiunoX4cPwNCD+62Hxo3N14/hvkGTVPMQ
yYAEooD3vqqWU2RQk+JEwip2DC7PkGRhgLKFrtrnyFxWa3x4U1b/9OMl+vDchLD2
1B2M4pPqHHWHDbsl5tYXEAHwRClMnc2rJ1e0Fkp1w4Y4hbhXWyGlIdxc0SoyCUd5
Ctfs6kzqGuwIivML24lDJfj6KxmvfbwUQiC3vTc8Kc99vBIp/D7EUUt6Y5AXRXyr
PhZKs9HAIn4kxih/i8WVp3Er4KFV8j7yOETmrJQTLgYv8/chnQyghm1KLy/WaHFZ
l8omd7gF6iizubjmHSnJqCYmFVR1aG28xL891nm1VbthIBHrWSb1gRQpFPov8Qex
zhkuFy2f0RTNK6cG2v8skdY1/QtAVFBFeQMlmgaBvFxVXY6RVlOd5ZMRaB19IR+q
RNZs+1zIkDFJoGD6/tNit1b0HIjn77XqKEr+KnzoT2HgKiU3cmI+T4uys/Quo1E9
VXcO4aBHJzd125zldfNEoaeX/VuPDjiRJvRlc4o5AaoEJnHHBQtPuU0K19t65RxM
hFwhGgWr9ggAmum5OvzlxwQfkHEtHa0odqST4OnnGuZc85FKbMzvSmAiduQgbqTo
SvPAt/gq3mD1IyJNGw7XGwcMMtqLklr+K2TqSPdWcGM3G1KzgEileffaXSW5EX7r
Y3xRQKGtxhwf4itwz1tTRuXv7XHqanJD/QZef5K9gDvjPPyd/tj9UgFIojm/Me95
G8MpzM3psZkDqilM/3QAqvUzsMetKzq86ZefqXGbhOi39pf3lOPWC5j6jVt9V8OG
CcpxQgIYGfnhZGcgS4NumQ8sr6H982bTKXLGzMfjlE7P99WUvnvlqdWJhGNkD5H1
1wPMjDNaiUkF5qMNJCS5YQU3IWJZHa6gzWxto9t0VM/MYn5a1t2QhkpnAJDnEr0B
5tbWMpXQQU+fTOnJOW8mNs9RWznkoOczwRGqi8d3OM8E0S4/D19l2NviCglQK+W5
Qvkh7wSfZKSnXqbpAc2xO/UnzAqTTBTR48BwUrLVId8P1Z1Kxk/bajQTenDV19Um
FFxdCs2MQBE3I1p5XpgOC3LfUJTh649CKD+3om8jiPC95nQ9kibRnZu1cP4QTKDf
PV+EeOE7WE1EXq/CHIbAyrrePfGgUK/LjIJcxDpqeJhzyHfjn+1V9JCaaySdxgU/
r9SOitbIzcTbTyxWiMBvhIaaLoeALdIoFCLORN/5JoEqp8zz0OB7Uud0YhR0jmHN
a9EEnLOWpwhztur+kEDjbkaSPEZugzIBmAutLL8yCkCjRQ/pLS5AEBQhSYfVzo34
S/X+zIKfyyA2aDPNzsZgARUGZe0C23aEjdA9bNIsUkpUbKNBrjdzAf/Wr4UC881S
`protect END_PROTECTED
