`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KYuau6Hv9Iuhozk3Cj1z9e8pXLn0edGE4X/CPLfAiXxXK+W7rIT/7WCnJXoqbyQ
bG7fY4XzOkXKV5RIwUJi3xFGb8SXZvSTNFT/F5tSLy7Yj+WGuC1BK815RFGNh9/n
Fbrze4oE8p24Ske/M13v380TU5iq4oHGfWYS7GN+2Di9GVlQhLm1y9NpyZts07II
Pu5o54+M/aHFPvOQslvFxZFORdrq8SIS/RQCMFcdDhu46UsuNMDsiW+QHET1Rw5L
9/uYDHrd9bVs+RjehV0mCVpEFZCzxhHCpZuaym+TorLF3uZRSjHykU4Cl1yIUtfh
zSy7QopyXNiWKlwC5aLOyW9V7LY0H8hr/7AgIdgneHpS/a0VqFp4p8IljLwNiC4m
Tr1Gx8MRxq2CbbpH9RLjir3rWCvEL/WWHWCehH4Ge03xftrSvLIp/MrrlnGmaneX
exJEQP3nrxKZuJZ/pmCBw7KX1M7lWEP+73FZjzzCT3B1Yx6gHfHS+1J9P/VUUKnf
TzGDjHAewziH3n5PDo5ORjqzBwKXElJYqbYiHm/fvAxlvoQAz66JxqNccVBYI/cS
C70JLUUdWCbaCoiXwBKnGHodn/YWHpiAgRwEUxGWlJkR5rXYXRGSvFnsTjLBjX0B
Ii4suLGUVapJRhGSbVKEZeTtSi+noIO4Jk9vn/YvbQ66aWletolH4R8eZ56kHslr
DOptPuBMSZaOIUZjgl2wmATLeyBVtQ0/jLTVCzZ3rKo5YEC51INWQrkKy3ACIVOl
BHGYqb+oU6ICFWHsKLuiYlrARFzRq9wDvkGN70+8FCG4vXuckc7gYmb3tNI8ZrED
i86+vlcuV2f6Tye0VFQcJpkjegGcV1M68U3pQDodZMMJpEnYeGxrrGUwMgOmAH+w
boS53xSxRY/VG719JGTBGRSWe19XWn2ouw8gS94uuciUIIJqCRdIS3n3gCYsCkiN
6yBpjBPqERu2Vt9YPCllkYAqLdp5O76VOcVk1vlUAlI=
`protect END_PROTECTED
