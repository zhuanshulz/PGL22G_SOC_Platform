`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMQIqCfv5HCs9J0rBcfTd3/38J4GTc9pYA5eHetvTTndqAenKpFLIE+1EcGPCIC9
0RtbppxeuRvgU0akDHj/EUH9Br02Xh5HIqFFbMzBWrrP4okoBDwFgGa14av2yjnj
py+xVavOJ6j6iUmIApMm37wYoerVYx3rYHa3vB5pjACoOqJvK5iziG8JbjWlnlfH
q+RmV3nHYbPjp4NQBDoZbofVeIDA+Nhdvrv15mVceNaOPwCquKFniGxg5DU0OV5L
4s6rOlaN9jftmAgMIOEWIbIbhN4A7es5hBAGafV2FxZfGfLirmJIZM41TP7D1rsy
sXFceC47+xGtZkEZeS6IA4m7033559yvONm1rqKHmq7jeWuRojbSJEJGNKqSyfUU
0ABe0UE9c/EBNpAnIeFZeBTFSX0Pl++L21B17tTk21KYQlMx7VdlKPlHyjO/CmQn
kDDSDCiDXPZA1L0DEBHLI+IBcGEQ8Xt+wMsCj/1+b3453IT4mixIwgGiMjf+j+VL
JyLbq5cvs8Bn+QJOX+5uQrUMunJyJ8utEEQNyinjBUJeWau1YFQwAMChsNBmtbeR
+2jSIFTqSyU32EzQBeSS6Z0rWmBP+e+W7/GCr8ix/Tcl8VtZrcgqqma30za2Xr49
OBhsYcpyrmFOrCHvvVxgaHUo95P+vakf9RuvzivAzbPSN29hwyWEMUkom1VV2s0g
mYDA02l1SOkWoeKsRrKX+qth84LWcCZPSAEWUKi9wY1As69l4kZxSyYsSfme39/G
lUYrEL42XqdbGqu0Jx8flxoMiR5b/RLHFldFga7Kb8kcTbtgk6TwVRlolkYwFblA
N+KQGbHuzNTrSG2N6gDzoc5tS02m8hlWu2j3vUym33dCK2/zTRZNIz+NPJUgXttl
1CTPsGu/923XkyLHlkUh5uMhDOfP4A9w1D1/VkHNC/DhHdMaiqbAwpWN0TyTYG7W
QPZSI+hefhWzIxUU/A50j8gMqgV7ohV7A05kOrz/upFUORVHeRh2f7JGblMVrD3m
oVQN1NTWDPSca23+ImDQP5BWvWOv/Uxokii65ff6ISbsRGSmDYlNwXvq8w2tzajm
4Fu+Y8T8FOpfcGb18XEcGqEOQPZr4Ut13RM3UaYsuWx7cnifNUpme3icBX/Q6Epg
HtFnUncy0bdj5J7i4LsVNSPNN8cx5y9/8tG9iqbH9eaN8/qTJ59Olw1hnFy2j7jA
mXH2aEVEuVZvlQZXkdsbVIM8pvFMBiRQSvZJWTC36CN9+IxGxv1QwMngRXFDnDcG
AQiIItfVFkn5yR/X0AMTWzKu5zG1zoScEu3flB9ct1OBjIIEW8GPhP2aspbYI4E2
2SYBsfMX8Y5HWtO3N3wAYG+1naaLwmZxu33GN5+TUMGqQQ3/nnJXX/CUMG0BURou
fNGIIPXv5xn5f+D38NvN8CbKj5v5U4ZaQmWFhs7xAyogIcrwgq3607QBWaTek1+4
JpUiecN8JhRTYJby8i2PKcypG7ZUCbLGVXtU8/aWcgMIzUUWUbupFj4IFegPNnWw
Fkfzqac4y+1SWBOaK3MAX8iDCYVD8DIAS/VIf1JBdt9GRmCwaEVeauXUiXyiwvIn
2Y/HY8tlgnBXHiS6u62tRYgaaR3RfNytobXd36JRQ4cgtU3uQ+gZ3RyroSwrWB7f
+0hSuJMBoOSaT+G6Jtj069bKVEe3V5PfwQ33x1GH5+Cj+OI+lCSi5zkDUAMz2T8d
UPLMeLO9XvAJwS5tuvKd9uszpB5l70KFtwH/Bnp1MeGNXd5hj6MAtTdPKICa4S58
sBf9ziLti+kBAjtiTCoxr664LfQglkxjFO0WegMZYzLonFx/6Kz12yFWjJot1qER
j1i87fDZJ4FVpvNwlbyefQ89k6EBtps/d6bYUEUioabrI6v300SBB+u/2QOHCLsw
afvWG05Ke8pVET/wDge7EkoI2/sIKHWtofC7vLCAavlS7S60jhBfKXGCi+oX5GIU
`protect END_PROTECTED
