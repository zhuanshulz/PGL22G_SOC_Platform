`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ap5t6W9ymXzsYsHEqJ7sFPqtKEM5DuR/+VcWo6iMcAV2NSJwN4oXiJDc3hZcdNCg
BPD6T4cGKfJ4bJK7hvjy0Bpux+HBS9sy3U4Qi2XXTWNMqEusmI3VrvpYz6TrPF/9
FF52M+cHRA5G9j2IfJ2QtI5KXvGkuZPov4zEo6tb176y68TS6RhoKHOLBcezlfHN
f4KQF0oKLbqfrlRBprVyBFXTgbkTB1tL6nxokE2VN6Om1fblYcX0iaSM4cvEoWMY
zyXZx3BacqspnjYo7pVlQZ3e7TtFVWIM57iAYdEPZjellWXtbXS4pxmEQseQhaf0
8pfFBnGV75aY441TLmy4hYzqG4Hs338FRC9JQ/ikIn2XHgbDJnCGr+zGzhc682/B
jfJ8J2DPF8cX6Yhvd6uBUzc3gbAXPYsVlqZjTMWmFdlTXGSpB2APKOCFgOyAykJ0
q0FGeYofYCA72rE89m2Hi1Lqvihk+bkny7DWfKGO+HeSGAEHiKloapgcVcWbSrUA
MbVmHv4eXj+fkJBURInb++rFHQ6D4cCI3RIWV+RTM15KI3k6pChQSNcRcXlhde1S
9+RxVDkTRJ//QrNHs3kMI0Q7FBuDjeQwa5nzEAigjnXJBzEJDWcsYYfyIS7ao/aB
3N1rNzPT6HtKP8B/+VzOUjWKPv06MKD0as6ERdE/DjnEIeraVvJ2v821I9cOffsJ
pv64gEZXGLxGt71C86TKJg==
`protect END_PROTECTED
