`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZUjYsdntWvJB76BrNLgOo5VikFWqX2Npx5fDbnU/q9ToKZYYElAaPzGjmKjS/UbJ
3VK2GIDjY5Uvr6ALCHgaOKP6kH28Z+PDWPOgICoCoOG/55Xmaj0rAmH5noz4DoBN
qWItcKXhrO8tKJSg5dk8E3drz6cou45/xnxA3Hx1xYEfqCpVe8WfJUSy+i5z0QdX
GbbXWDGcY9m5/HZD4iFWQkLAJonUBrGuwOt/37lWb3IGEFKLMRBGsTK8VS7BDMux
OWjtZveXYW3DY5psWYk5uV0C+mgQKCT9dGnrwf2IG+XOKWi9q4SBDP17lJKgfIYS
hHI4Rg3sBpuh/sclWlUm7uHd1csSiyK00Xj1R2K7Q2H8/A9TtsvBXROFQM36o/8M
40qbB5kMntbDvS2+p/dU0PkIjvXsZXvVEYSuamMX8PiwNtAZ5v+pDHlmKnK23Mlj
4GRkmVUevfTh7b7/L3jUpljwt1fmYoOIwtSKN6UOr/ikvSMsoYvW+A5UVMyoLWm/
HcSrthbug+5ESOCVym7EdD6EvujRhLIojf77ckJBqAVeWblJz3H7cUUtG3RX/sQl
/mR+Q2rNx2+rQ3s9QrarA1Lvxh4y8PUHW1pVFw0SdFQi35Ecj0zHlI7wEp+2UlUT
upyBAoRVCSPQNNrB+6P0a8dnkyc3QSYXLFE0GVpookLVa0kU/LC9+weQKjRbN92s
XQxso1NnuF2ZcFV31V8ySCTAu6P58L3FrWiR2Mg+2aXbKs57JopYLhFh9cxbVAqr
/ploQU5FVyQV3ELAAH9uGXiCBHkdpqQhspAOMZFdY4Ha7afxtVo8Ane76vqoLki4
XIG/QD+y6YjYXFo/8Vyqw+dfBe35uwLI1pHxTx46p4j2zLm+YEsmKpy17oCtOot+
gmu+6j13oXuOTYowa6rtJDOZJDimxPeCZLZ1pFN5MIierb7Q59gS9YtXo4QXJeoK
D9VZrJQgNbmIEgnhSeBHcLkCFnYowSbdKDCpsPtyKrlFc9mw8G57iP0RipMGGaB8
0wVpBMNG70mKQhY5wJeL0ANhuV66g+FeoCVHRKMcDg9Nlq8qMAMzkj7StRDOQiFz
lZvw6xrzPvlm2UVMyU09Cy8jMcg2gvVBdjJ9J6z2gpyfqW55igt0CFCpgufLGa50
WNaSYObnaDN9YYG38r1rpHJjAdfG1tMfmKHkeyFyugDv0Mo5+7LODKuu+Sj8nn2Z
1hm6s6nl27LQvgdhorSg4dL4tXKmPpELTAgPwfP1sfYyVJ0UkP49mTlHfujybSKn
14krigh6s6UPVk21L9lPlOqSWs5lIq/WvdOxpCeR7qtsmRG0vpPxUPMFEuV5LvAj
U+2u9Wg6HsbZIuPCiaa2qGwLgDowJxrMK+gSRitdhr3A8MJTaGRjGvpMvCFPwH3r
QPlihp81jC631uM8weaYKn3wXaaXBgAA5g6R+4ZJUb3cDjqfw3XOZIKJWrdfaXwL
YOOaI2weCcJmA0Cq/Wh5DL41NukfsPfl2EpG4BjyZjuHY+B5kMRv4Dp3ImThlQhy
tGMoGK/Vaysfa9fCvr8PvFSgDJnE4+kh6gJO2F3pygglKze8ccgFX4tHz84UJpLC
rCad6eTgocXgqZjhgWhkP6NLIYoN0XyX/7MLn762eLwF1reYz4hhDJH/zy4aMWYn
oBcJdZzGBS8txs7IdVIYlRzhideMQkA9wqFUBAilreUljhOK7dDOqOfNkSiPUm1I
PGYfgKuwS62r3fY3zi8Nai67gNbP5+8yrePvQe0sCl4W5xyyIznLX10iE+fBV2c1
sdyqooY1l/X4imTQBGFavw==
`protect END_PROTECTED
