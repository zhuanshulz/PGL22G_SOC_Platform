`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FMlT5IXv6nwmx/iubiNfB2+BBwwERjd0jnJWWG9hx4g/dxoPd8J/rD9Ne2ZTkPU6
XxUajzsTfTCAJtXRsHUKfm9LzpVK1cmxGtvk5VRsXrzx71qLNT4aiGgxO0Wp2ONp
+YF3LJv1TpEKdfVNHux7Ub6oLbiI3t6lTjBVOzWx2SlTVjMcBYgcuzhouqNj5Da0
n/oeLyBDFlaxHIFYWWF+pMFItpKYcJTowxEEfI0NBc/DN8pBdnLCpNLqbRzjmiMC
4Nr7MOIcDlMz36IZCcxchSNFxQatKRlxVOFq/8M8ArJtJbFrak0KJ4fe96dVueeC
zWIpp+X2hRelEUZKjWntMET/8rOSYblgMjZqTKFY5UiLiNKSWGsda7aNjq48A26v
vBKP5WKUJOMr3FDCqtfqzH0k7gjjDNsyuedVyQcZEY5Vq2zWT12AHQZ0WxJ3u9Dv
eHKuF0V0n0IcO0wRrDlOV7cIlKDuO7XDVhCi0E+UTeoRjDEuUH/pIgEAK7X6jq5e
P7qg/UmA7ECnyw6ImkCi2KswN1HI/eOu5ox8Cd8eiePY3++TFYYm6wm4m6V6QcQE
KPyLeds1tHUaKzjnOaYSPeiX0O3swAHblAb9qUqZLlX0L3f6lOEmcqtZWBALwuOf
qKekDXBrIXOmjsiBf6DugPq4h4xofCguDITSznVktnFv5Xx8/Oi5mRv0Mbb0RzDQ
2JOTaId4n/vJMFXn1yLxyUKKJefgl+uCYmlXPzDKBdQeF8pagSq3CO2fCiONGwvQ
TbTHk9jgg2cCG4AdtPa/jMEE5gC5llOLp2C+YVvoqmIhzpltM1THwL3DDKRQFVMz
+ceF070KbO4qpEi5gRTr9grBxQW6pa7VIunODDAnDxdkOvwYEhPXmA5PKX2hbL/T
b+xPvi8ZM8B93bEcQWs29NlH7kPy8Da8EML8os7ZJUDxrBynPsgpdi3t6qwZhXFU
KbzgUVm+WEHKF6uHKd/9mV50E0KuLnelIR+Ds4JpoGzlc99xkDVvLVyYOX06+CTl
EJNP/bGx1kQL6At6q6WsPsFzdMJzZKMyW2vmak4LMKPWJp4+3gYgW2+6JpJ/AYGJ
x/+5nT9fdPYgijsod/tIRA3BkBvkMR55zFepVMWzCLNer5qd8r7L+eVfbBoRXpVt
iR6Guy4UCzy/SIJzmR0ejJw2Lv5aizCSgjMZUCw928GwfCltoqvmoopIf2zMpkQu
H3uydxt84j+VaM3iwvS8U5nF/5zcRsGbLvJdnI8nb4DJXbIgTDbxfNb8Mayvejp2
wV9ZoBee5wnNJKo6OF6TRHuoorfGrPIv50/fhtj1GwoUqy8+T/FsKhnGX0eom6w9
C8aqpwzNRGFYQZQ14i+lQgI7A+kctDqAKAMYuUvXJJJY8A07BfZiyFlkdPpoA4o5
cYn43tioX0PYEI5v9aGNlvVrUt7wDPWnW3TBpg6ZYjcc1wo0MaK0YCTh9SlaQLjz
9E6m8sKZn8IX9+D68/rO7mZLHNvJBZ//T2NIP+5CffmNr9cX/9zYKB0uEF1hK0Ku
+Vlc/NPgxLa/SOB5lixO8I/tXa/ZBMTSMCB9YzU+llmwcobTUFRmGlhJCL/bdapS
zdcIQurUJ/NgW7jNv6OZBv4nBjEGUohaNGj/PYjc+Dr2JN0M6A801iIveiXxwg8o
HAfa2lb6KJ349M0UlfjrG9M7dwSrq75Q1iN8+SKNyOK+08AXoWQ13y/8VTqNqdI2
bSx8FiXNhWY09Z2OBAs5CSFYt2nn/O7pfRjWwFobhqIKlhIv/dUD1BK6zsgdZ+pZ
KgCWwPJGxulSwRfhHDmUQs1kgBn8kj9CNCaOvbeItGLQRIKe7WUTr1Hw8YbDMtMy
AmUuFv0n4LYAZjEjTcO72eKz+EvSefRtpRLg9FkfqUV/URT6SJeaP3sm+QAj0zfE
15d5N+BQH5RT4CRITDPM3ZBDmKRW7PJgbKAXPXmxLZXIUHt6YUHEYtGu61kWseyU
uPIuJg3WihP+vQdAhQtMLXhP/pwtZIl3TRosIit+8AO5MaH3QjWVhBo4/KSruadw
pACalDoAipq5SnKuQ8SrD8ORGmzUuzypDSQFn15+TvOhqGqDTb0HEVrQAG/GqE0E
J0GlKebYVGr332QVf5uDV9Vw5gFRAe9gxnwiIZnlnDt2ulaoA+dEhHQp6LiyULcC
TFzicTebF8N+fjT4FGCsaBkB5Bsg+4Mad4fl/6bHVBgciWzPBusAGfS1GjjfOMqp
YRC3AdpTp4cuUhsmb35UIHrF29wr+bwmjnqIXDVD/yLtdTp/60Myd8vRMxvbWdVM
Dti/G68VzIeDP6N5BvdJS1sytHx9LRJllfbToppWCgj98anrr/WtD7o+ttZYnKK4
ylCBkz0KNEY4/V8+XkLE+aOGbkuARhoro/FOqAk0YBaIF51iBFoUc/tWPPHcU9oA
hT5cwz03D+o7z7mLSwtqP5HxJn6nSG42El0sL86dN5R8bSvnXebTXgGvOCL4l1Ea
sbzTJ11RmjN+DSsOwvW1qjtGWxcSU44374dP8+hs7sIBvI58hKguxdAWmNQ5lS70
cpI9Itkii96pcdmZ3nnJ6I+uCNAZBU5CQ57MYgkfqRUJXP7s749TSTYWtszUKfVJ
/irQ1xclbBfD6Vb+Oan/DT12aAFfPnaCmQZg1qXK4qVIwdpxoqt4+q4wlyB2ockI
9CuDrQZ8Oxqq/y9S1+SpJsfHcY6W9ILv1KGgPy2izgimHp0OXc6+m/cU3XEMBhRQ
dPTwLoj+XJt6LCu1X56DOgZ13iQq5pwYQWXviVXrTnaAgzTQnon+DuJO73ZPElS5
Q6eMx540bMVwWd0BG72YMnXHZ6TBbGw3MfHSbnQJdkIYzx/BzJPS/v/4GWcjGLhd
CaAUAj+YTqxmA/cPsHp1ypRP5u0DrW1aMEk3xBe7dADA1wPt9RYxasG/1VDhBZup
kBrWLtBKr5qCm83TGwGLDZ5tof7xthxU01h4IBSX+gZGU1KlK+mxGg0Ihzfpwa8/
hgsijDTIjLxQI4TB4xkucnnEeko6rSWWbM1GEb/h31XdHbCHs8GAKe7Fes8QUtJ7
OOEud55eaR/Ljl348IzycjeBeUp2rUI3AHulrrZrb0xasZUiUCaoq9WZO3dZpDXQ
wMRghqNnbtp5DvK7s1qmvTg7RBCL58wC+ZzyT1c0G2XGZ/Yp7L4ySOAQ0YqnyEy7
88c6l7etwHT2Su2hv+p8pwxtbW7VlHfvQ8eCndQRzELr26BmzN1400Zk38kBrE22
Z4wwmdlDtBqNH5POUDoZxbLQOYbJGiNOOC7+txEcO5UVxgp4U6fv/FWYCxzN5r2F
sYU9S/2KrjGUSWW1VfE3022cun7BF45mRi44gvgq5ctzj6ZG6XHPH0JXj8B/MRZW
K6LvAtm9ZdtRyxFcXqFM03mY3ZTvJHGBsz0NH1Ce3k2iLoSmD5kC/Ackcnos5Blr
zJSvgJSOut5UcKLH2P600jBY0BA8BHKq5VR1EJmR8zLkpoTsJzFlzNp1BgKQSj6o
dpjh2hYj8qysismKvtRWR7ZZ9C+8lQYM0dlTiKB37GETYOylU7+bg32Pxbp/mGRm
uc2dPcN9gd9d4oK2wj7cTy4Gi9FqVQNFwT3W7/3HnMEawbYBDbkxjf0JRuXNcHkR
9jpUSjMvl2shDRObFaYT67Vasf6vnvPqs/I9mhdBZGycXPaRGnHC8NE3+6af+w5R
VWKCHrjpHkxrdoz2YS9UjZwuNvUnN8OjFGfk1tRpn1dISwBzwSO1B/YN937Aheyd
koTetQAxEE07Qf1SGxaXEJ8kmsdaBWoO1QcN+KnTnLWFbUVdrGCBMEgGSe2IG/z/
csCQYBVa0NDPjDfll8o6THnhQ8y7SepRIezb0fpcyqcG2Vwe36aSNkC3tD44nxCS
2Qg+2dDgPO0VnOu2XaTVTG7LrlGeLrPQ3PP9zLdfMVTLxOAJgen2zL82aNbOsRwe
mscUbFgS8Rju/8zjtNCQgw9PZL6bHWlPFE9JoEkFI6ekD52R27nuo8JbZk8xLEl2
W+yaFNnPKMRNGk0HTASEcnHwTLAP085VpxRpAkihkVVdn3rKU31qF+SiwYYPSRq4
rkBfkCHxMkLhBI6gBFIQk1ECFcgNsndKcGkOrhZkz4TNIDx0U2oGsrX+eVsJw3Kl
q2VImLQnSCT+wPBTns7etBFj7dbXx7q9uBoun/0dfMZtut6S3tuIfIc+MsbI4nod
wL3fmpcupscBdUpwA/AlpnkDgEzm9q68eHkAT+3s9TaWNnoxVbdJLzWZJv9AQgzb
E29Bos+bh5vMenk5EIlILWTFyHmufj9GAzs/I0bJaZ+HLBWMyrEatpaIMeenFd3H
iyyieRDzRkw+GIhk/lsfUIYiz2I7hOXXT9S3jn3SghkjLxJ5WM+CSPtkcQR8Ah8h
RnJeqrPcPe59XUwb9WFKVdfkZz0uxhmG+KDRMETm5Od3KxtP9Jb2fciz+xK/RJ9N
V0ykEYUOz73z4XUiLOXG38sQgT6X2gHfxGyih5+km/GjIS1yf+P5lJO75q5j3o+f
u2CmcOyDH+GypKRYSGwkOZDmsXztQ8cNKWzL7qBmydlixPu+yk/GvMbdB6lLfkPD
ohSpKK8lFBX7XekxQu9ol9mM34kwJxnPuklIvR28epmmFGpmHl9PSpwh0BWbdBcq
`protect END_PROTECTED
