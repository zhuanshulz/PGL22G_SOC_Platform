`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NB4/KpYOWNyzdz+6ba7u/JdApir4GoJSi9j5tc5wqbpz77IhjLGFXZCwdTFXG4E2
paU17B5Z3m7pRRapLPz0MawAjFPTxKo9cpYz1BY9/byiF8SwOcFQtKVzDih4k6lN
CR878WvMNsTqiZOqn13Lwn0xqcFly89Pd47DeHEnu8oyhWw1gxGjjdtzg5QZ1SM1
eLg6EYqCzQLDYc5cCQ0hxoxIwiZDe1CpGvG9fKpa0VDX9d5Tfx3QPZ96erDcYvKB
ioBxIRiErzqpt4T3ez8VIdbm/kGMd3dn6dEAKvmHrmhvBMqfiBK9DqEEgbeQzzTe
AEk5X5TKFqgaZM0/1+d2CzpljNi74ikuVveF5sELpEwK0x8HpS6F3NYAh87oxPtl
CvA20kcIYFi/jnBiRIrf4/WS1rUhXumamNoMJgJD23/1a9fpBGaFY+Jc7HIOGNHp
4Mjeq0Iux1EVU+Tz9c1DWa7Sy/ZTifmtNonIwiwDuvW1Hvr0OaPfxlqhDTLKqwx8
4qSUg7fwNXdxDNH2TadJB1urKCKQe8jbb2TSetlhldOB1oc8gt/GjlpvUhHBN9Me
FONPfVkJ6zV3ZjPC3zfKQLkGfMfzmeZMYQ9gA8uetc0s+WuXo61uezZRgRBtb81k
QhzzMMxp/2XMHOUm1Gyy5uB5PVOTtfziTi5QHRtLKx8AsYqfW/ooYyoYLSrdcTFI
jUxW+2gQZlp5xTkJPg5D8mz1Ta15+Up+NNvimrQ9vyg+Q61E0eVuX8v80AuwtqTC
bJQuUUCagcwE01cpLEJiYhBH81sN4alpkCpeux7b+BCIpepUi3sFXPBpmL+Py9Ld
TffSbOWPhAe7hp+SNT9x+sV5J7hY8tbRmIkOju9aBKzqvcUHwiVueRJ/sCqz6De1
3OJHjTqamaQ1RyY8ghpjHskmG+85CdPlSzhtcD2xTozirQWkHIO5se0Uk5Rcjo4N
0EDjQjzEnJVR0zla0hLH+64HkGYHlU1ftCSESf1Qs19co6KD8C0FUOFJgUa1+Cq2
j3XvkuHLrQgpNzTmzy9vIzd4VeXe8G6HT1Izfc+95MdujrINVPLFor1MkWVwduSC
757tIjh88T+Nv83l0ioSOLDeUGuLSBg/8nG2zzCDZkH8+aigcEm86tH8DnuhXV7a
7/szT5LEgDZn0Rz3aUhCbcyJrLp90EU53aRTBbC4+1k83lpicqeFv8zluINRfy1L
DeO7NPIM7rxdg+0VkoV5BseSwUU++a2/WqY0zMja4ZC24TggYWeW8VYSITfysxZN
wHSEjXQ1Hm0wOrjUSijLs3eNsRMKUwmOYLPTet2zN4DflBdchiomL10TCmH+4cYd
PE5Vsd3d6n/cNAvBZLEyU6KshCLnYQkLgtMk6gTlEbTAWGREuCxkBdq2vhe8DU3j
oxRhbdcyheQyPtlIsiYnWjSCj6rAi8K+NVkE1HDBE89LjgVDMSEA8mTdQUYK3aKz
Mj6s51b7QHiyjXYLxXJabGK1/BUhUwTmOMOng/RTcXX2WotuywgkCDYGYFc+L4M/
GTAG7GZ0L5LTexepDhFRpLA3qysb5cOivsGFF4qFgZKBy0B+Bjg4EIOX1WrUbfFa
TxOjfcGM6HHb/WlCQ9cUHqvvzbN66U1k0jSIJCjQ6JLh22aewV3PCD2TEN0Tnsor
YzsSOgHdpY3fX+sA+MRePqsOzuKvYyPsB9Xjh338XOpLMVgcpA8RP2JNdzML/m5S
xmWh/sf5p3FfhNO2fz1UGg4XMLXKH1adM+VUixmv7Z8QrOTLk6uwWH7LjtCQnE/O
vWQ5+UMPlaIEHkHooH2REbGGpjF1DXW+VlUPJm6lWducjiQkwZqmaxEAgZjO0kvS
M+a9Q6zp+pQOafi84FVhKIHzePK3VP9l2kIUzaX4bIIDIucBFo1ilV8qekOhtCwX
FeGLor/2yoAZfSDjP4hWr5uDLeBnc8rwJhR1MH9X0ohoUnYcr0KMUYTES4/FJ9C8
xuvy08FQiSovnW36H8tObJ2U2R64k7tWuiG1biypY8mbQilYzczbjeVxHCBbKsB0
KhkOwzT128m8q8T4pnd5HnxRlXY9oxwjinka4iIukohLGID5JhtxWG3fkaU+iaga
+VVnKDbS4nZEnY/ni+HblpwvhHJa4K/EOgdoDBPqBuKLQFCxX6w8felsq47Qggn1
UD2xUG7wFwBZlaLFujekwIN5L3ohp+6dMcCPpS2QPLcWkBbVFrCAGkNgPEnM3Y8O
T8NETu0GYR7cXqOLIGblY2+AR48yw0NzGCIRG9+gR6s6miNvvaRFmxUbTITDq0MU
OdbWHjSMvjLxeqoEw2lBWMFMrm+qK8MzES43bVhy4JY9dtitL01ptcJjyjNiNb89
4dAMnlslyt4U4uJL3NXq9vQCQTlgrGDeGLwXKUEZorRtBfzwMBGPFsosbVH/UIHh
ie5706CV9Q+Jwgf6oxC+mfheAEjaO41t9giyY/z817hQFa6uUC5W+U3MWDjGXQO3
ltvgwSJyx9OWnwQ6rGMl8S6SrOzM6Rf7AT5mr0beXHp2hrOYh8uayd3d8N1xcwlf
wdGKEudszrsOKwMB1o5zNklYr3A7Vo1sli0LIRS8H7Mcvlaf5Mw7EkrCcbQ49bim
oyGydae+f7LtLF0iv9ql0TA/8jIwMDJFAnb77qgxMnerfyLeN0e2BKlXPKPrKRAy
hun8vU3iyXSRGHNcSRdSyj4Ti2nt7HIXwptZGxVWNo8C+dMAaX9qvgkVniZ6s6em
vFLb+RcAykpWELPSD32O140xRWPPLDPriFIQzwfccEvZ9kYvCIXoP579KK8kbeSc
gwpyNJTtBLLypVEE2A8nYJ/ni/TMfsR39sc0q6YEcbVhCFq3BmSdBPzaq2XrHTIb
C3fFvAO8fiuoJab20HQZ0cnnTnFUUMOMU3HLGANd+LbfxiL2Mzsbs5/Xe8YVLejc
FOwfICWMCbG0L1z8dHjPJ7RRGIP4aZ7bkK/OVcnU6yThaQQSJYcChihivlxK1Wz4
rREmB7NnLY9WU8cHUfJy8XNeFCGeGf8/PyRiQsJVEYplXnpRqIN5rgud2QnztJ2e
FlPN1qq/8h9MN28pU9nKtemfnWPum6++QkQFGPzmNg4Is6+NzpqK9eyuAcMZtRDh
yucaabWbDLwF7Wt8F+x9qAg8pm6Chdv8JFmJcKTdU5DFJiH5PTlZFTM8oo0rhVi5
8YqIIw+7PhiOsccVh9I+/vTO+qybDBtkot9GD175gtpKRHrPZ+lki508KPUvKe6z
9k71JGJG8vJQgGitEVETHX6Ecw09sVt/7PrX68niIrZ1Sv1YjkEZo7SMCAvJHjWc
6Roamojsb1Rp4bkqYVF1ts10TCHE9MJV0wJ99drxnfiofPyRGJERclf5H3mx1VRk
awDXjAieXhcRPdTZ86PV9aVmiTk88NpQE8GAktAC79SaT4oIeNWXNS+Y6MEqm3J8
LP83nFUqgBiJEYRfD8gaVdeXw7DBp/K2TPl33peAlFJ3qTHa4UlfJGHcQjW80xJl
nmzYf8gNwguRQsIaQzP6O08fV88dYVYDHZL6KtRngyNNDDyk74ZnE5jWxMPB14b8
UlpbWwLANPCHDwfSe6FRju9aJVdZk8DRtgLdJY1+u56vPSft2M8FIqTng8nze8oX
kAfLOp0dMy5QLzrO3n5JJUwYnkmj8C+yhu9HLC3IxHJUCNxMgSlXM0YgADP5MjPX
L/HCk7x/XeeV4pdBQ5pDlt75jKCL/XDvmt8VigWgcUFmoJjtWBK4UmkwVPssmL2S
0XrT3IibyOlE2Jj8od8M6+98XEnGW0toZ7EP39Ali9jGwoABW9ZuNvQtlqhbwwKz
EA7cZjqidsO463EypruTRAGftiSw2BWIneA7whDtpqqzifc7gD7GBhUl0GEyrxQ7
ovwxDQsDkOvvncsrpKeUCO7LDJLI/qxBnYsVffRPgRL49GXAiIer6UItpRsG472G
B82eBFxQD87C7r6hjQsj4SU29XLgmifL8SK2wruLJ5RlW72m6a7LLsPh7wQtMO+m
hFX9IAV66BJSVvcDHdo5QTYKconxN75xn8eqBLhncdvG93by6jelx1vFrK+Gv2x7
RFV5aEHLC7NfY8fR+AB4z/fMC+3oAR+FAMNE9NV0sogtAIdzLKNWN1bgLRw0J5ze
7oO2b+4uXtoiZjNN8HdUfDsC0MGb2zyZ7not4DUdD2uoeOL3gXx2v88vXwpriBqo
5uk8SBV46GicHIuE89S7LyMvpbNIleb6m1lL+CmX2SrOWzybSI20bMOTfZmFDf4s
NKs8oGwp43V2wb1Y/Q7EVaunNi1XYowR1xb5kfosQqusybIqKgiP8PaNoQJQw4ao
Xyb8dfaAxwJ0p1KzZpZOVFTdHn2BafzaqiPjabir8A8yALphioFrjqbImQCNi0e0
m9nQzBYdU19GqgQGQvXsdQthDIUR+k4Pv7Kc7Ikbg+8uLYPt6DJoHjVWKX/zdqB/
8/IxMwuhvGima2H009x7WSnNLLVnr/nrzudcGixLn6LsDAcKmlu62Dv6YWYNrAsn
TwOpli9rAcLEG6CLE7f690c2ujzvm/Zmu6mcI/oqqW07jBbgvL4qjUnP+HkEtQLm
RfZZToMV3QOw7PxqP3ojaxaXRTY+DMEV481P8i57Q71BqvdGcih5id1B495KwrEY
kFbiRf4UiqtqdeZawH29jZQyX0hBfT9UNfYFUZ+LaGYPEAfhuKAtTYGnqlevTRYg
AB8tvNrG5x6gO7mpncWgObTfnQdzFzck3l5usyUv6CDMoVx+C/NYD7BazoNOpyU6
Ha6/FGHiXMjRqfkBCqdZ7bQomXITLD7JmhNqiJ3tpz3yv0LpdhIZLiFUVedv/+Un
wo43rodXH1vP8JTG7dM/4yHEJ8Sutr3N1hwBybki0yhGB8uokNY7Zrg/PKLjkO2a
2moVMuJYEQtW3mOEsVPAVmPtOxZN7ItkIQHxvTWStnLHqkKZ24BZH1ihMGvnZa9H
gTYYUC5iFIHSD5/5GNvhMQTwAo+ZiDBfcs425hBelKPEVHdl0vPeeWOlBYRg7KWG
6pnEtHJ9oZ0NJJX54QgWb/GABsbv4CpMVT46bneLqcmKx3gRzotGnOJmv9BPeyIC
AJBXkrYqHcQwlcd6wXxYinuT06ck3LjEJW7pyhdVeuM9sphtfB/F3z+qGuS8Wz3V
uz5QukT3yGEnfabrl62r5ad/tI6RxEuiISSN5lJKpdXRwaFLR6j5BcopvTP6pgej
WMVOM1YxWaZF/yccqHlaR6X4nhW4uaRPTRypaGPO9AgWjjGcodDq2r1rINs0u1hg
ffufAZMCET97GTavVONdm8XeKzMYiPmaNbfA9N8e3VAUW8WdH2VbwvAk0++DgQ/i
vdz1nwItTe/D1ZMprNa+jje3+pKRnT1fvBYKvttkJEfsC7UVT9rLSyZpLXytMc+D
IhclYWXPdjPEtePes1fbm32AzVbFsna2I7MCHkLlT27ZhXPmqHagwOqkaCVMmoMs
cHcXiOiKvfUO1MliNA00wQFpFGmn3E4dQ/XxwqBYHxmaH/A+lJwbQ1Jz5jen0k5p
eMDrdt2Wle7FHABEJo/c+Abm6nOWxqkFW7FPWBdP9Tyi5P3N3xuLYDAiYVIDQsV5
QcByWOH5PLBgm55OVN0t4tmprvnUX4gOFJCkLHdI3wOIeznQu+qlvAw0WhCiEep7
NibYw47UC6eRKEUFYhP3bPq84tRCqFHmzBXwfD9qWozbBWF+1z2ztmqsVoom/tjw
+QubXmf6qMAzwcifEPOM6nGcpjW3BdWd7rlbyeNcotcfNGTdE1XCnLfXgJv1gdaD
xmbSR+KsfEckuB/Dfq3KDN2Ft9Os2Oct3RztkfaBXhIIuFnTCg+qWdz0MoVq9I3T
C5reRMxrli3R9MYMA5xngYKLCpI1QcCbklyyj2YP7FA/n5+c30YYNGDLNbJwL1Y1
d5yfblZ5mFWqsnF9GkeuRq8Tb1JOnhYc6eVIUjF0vL+eQAfZ4F5aGHbzTGrqb/th
fe7gDVYkkiPkwjXFvbyz2J4eJVGE3sQ3P9ECexZi6VFfsylLU9TgcYSCsz+pgJ3n
pP8mgHG6BnqwfuRgrsqW/EQ+YhQ4sb071fMZDP/xyBSgyIPemZlwPjg73ELdpe3N
BvlnlrZPkRNv7EiFq1CPm7fIy2bzbHpdBQywTvGNZdOovin0oRD7REF09+j6pCK3
nGswmmY8Vi0isSv1cyIRUABQpHAbgXyRtZs63yMwj1jy5zmo4iQp8yqnRkZIzSPz
S1QjcmJ3CRzRzcQ0awH6tNxxQzuqefW/tkkYCXoleieRcz2v957s/cupueJ1TH2i
ObLYRY84QZS6yxq4X36q7PDI5mGkk41J0JS88hhfWgFMvLiqgZh1dSBej6yhj0Np
cxWhWAwB5y58/tNKr/b5tkpRmv9gUFzITsQWf04vCCPyTz8l/SvAXMm3pXH3qXWy
iC5gCK8/jXeEoM0WAHvdGjVOEQSoNC3Xl3H2GpZbWMUGSqK4HkahTU2jLkVr6yKc
4PAHk72fNckIz2WOXGhlL/LzWS+S9XnR4xgtIEiP0m0cCI2YCewPwOfR7+VjCcQY
DyH3RcounJc3eHNq2JglXNDCNca6rNw1uruok4aIlYjCDisTBMX6M2INuj/kwoRa
PUFqJQAIjcZa57xvMUpgpRjWRK5Zp95q+HtrZs7+NWXqZ+A2AbqPnVtqp6nMLjUE
ZCPQJDJmvCba+HKL1ulyKi9fG6Qi0YDipAbMN+9HupxUhgLB8/xCKJCUWaoObTxB
Zleq1R/vH8AYMp4FAQK6zBbCkNjqCw5VRECfbMNTwKHJeWmuDkFxnrreNIq5nWcT
0O2djzVduV34oIjFFY1C+b+hMKablRlJox/z1Lt2U062Kv66FaU6kb27z3YhqZZw
QCiCCjJCO+ul6cDa1MN2aZVC2z49RFXDevYNc2FxE8TtQOGOTRrRFOfkAC+mAS43
`protect END_PROTECTED
