`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9IrgpbS2I2dNkxym8al61Fgnp+TsQsYZnQgC+sKfp4/Q62XAN4m6Y7L5lE6j0fqe
1gjdTdXrR3Xwci8kw+iYpJkWUOPKS3WWHsG4l/AsJCrKIO4o63Jf3DJDFY9kqKLM
Q0O2Uc/21k/mQTJ1vQ69nNAdacUqBv0j6ljnRTK9dVkbSMUVHxv7sU3kO7XRgqm8
K5MMfvmE/lPu10DmTYBvNStKC58UpnQtoALoSK1whd8OUNuex14SeB64qAX+HAqp
We5hRqHBykLjV4UcVEl90PlPanA5i/4NkWHn2afjDVD4Jj3vFmxM/f0RkD3CZzLA
uKq79kWXCH97f4WFhS078Qnnr68CyJrayTvaQhdJ0ovB5wPGuoBa9PShasenVag7
PUEsL0f6AhML0A3Q3rMMTBXdJk3gGyO/MBl8zBIrh1h6Q/62IsBSbMZ3Q3L1F2t0
Cjjjc3e9rjdZ3MdbAks89NXPMe0Qly7IFILRJZRF+4NZOsz2gJNvTRrCjsJO0CXT
id3RC+Q+FDM1eJQmuPzfbta66hCF2yp9sE6kEsCZg3ceaqZMHJrxtOqJ1z53keUQ
mY9dWzSFEv3f7Rzf6B+zAb3cYK3xVvzYuxHNRX468aZZOp8Y0JtBbJUsp0d04Irw
WIvZRP3cjL39BONelxi+TpQkjEObTM8oNsd9t2QgXBy+q7ERCwRW0EWgStnMN4Wk
6KbeDJp6SGGMCiWDbgcddOctt8Qa/QXYFytDFzzbZD14H8O7U0DZTYYlmNg50EwE
dYM32ubKsgQWZGFUS52KzrtG1qWlyqxBht9Cyrmc8po/Wa9oD2xOhI6Kkccr4Oih
0hGSmZ7GESlbEN/4xOJssd0ZH0rYClbAeqdtZgK5rumdeqeuKFNrbisfFAD7JYwQ
NJIXl/C25VxKLTHIppvEtw==
`protect END_PROTECTED
