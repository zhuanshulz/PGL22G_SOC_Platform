`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5B9Xa306tpTnEvhWOh5GuKGXL1YKKEh9urfGw0jWN50wV/SbOmz2Bryt/VFIxDVQ
Vy6x55nZ24hD2DU8Iinf2U1HdB1wPMuZhOxsVCz9qSdgeZPfr6XpvBUI2Xs0riXA
n0CIe7XLYPNH9vccYXNxKH4Y/y9T6/iQFolHkmUQTDPwklIuRHWRRJfwB5p87i8J
mPqJgBHYj31SFowV6HMD40i/N3pnR59JYbpwhAiPCtYmjzzJ0Mhq1aYmZyM+IQIO
VDIT6tl4AmL4VvAGtWMfO6gGvtzK4WpKH4b8Rbbc3IBZTS8WAFm2WDbDXBlWoXBw
g8NptMJCM/5k+g/R5gX4E/ZBsinqw24rI/LJP0ydHD1MhUOF3fcDBEW4QhxJjmw1
9goU7Fks2rgdgrkyaMCE6Pc+v4EHiiY2aUv+AN12ExuESereRW6tT+wqfpcr390O
7s5SnPuRprieEuTiKS+xjX2tC+fhGzwxvcRB6RRP7LOLVbq94ebuhspVX7SdMoRG
GEWDEgtNWZm0mheyR33VvQw0IDs7qBUU5nBn4JYWqyQOSulbhqZDhrPpxsQ1WiaF
AnbAAgA/cYKwLg32tarM5CFLFLh4OMAYS/Z09thbLj/JqOeh6HASeoSb9g1vbtv0
VrtsfuG9Su2zM9/2fXQsJECtZtW5BXG+oGksdgy6bLvyqiTC93jy9p0rohF4X48K
nthsOB+BbmdszLEtUEdIgV8aX/sEAXR2A4+hzk3PO5knqcjXO7L9n6ijALcJe/cT
wXRzBO68iJQavYKEaLJJHoXShrLAcdffhVyaWvdwbt/flqe6a5CeE/kFAu6qPk0U
YJu689fFfmQXJxN/t7SH0njpiHTSbkKqdp3dzGi6+47RyWnOm+EuC76brRCo0ibw
10UD5U2V7qXyw4Z/MEE2sZIPkHV96IAxPqD+CdW6fGNK8vEjVfEHYIPkPUbm4y28
gg0AKgy336O0kw94PcgXdZGRfQjohrQK0mJlHD/pRx1I09tdWQtqHTjpXcEu1jy2
J/koJ7h1Y+F5ERj7hmrbPHVNcHyvuhPvSSFEWxj8VvhG37jDCzZCN/xLp8PZRyxU
hTz8mq2k8XwqSgbyyLoR+iRUZU5tCuZ75NlhiTZ3EgaaWkUvFrh88V1YsprmlsTK
Enohe29cAKc0vnBS0nZIas89kUlYxbVqFwK4SJ5d+1KMgpnQSilWDUsSe6Z80YpJ
vnJOPgVkNbHB9vbmn59pWQ==
`protect END_PROTECTED
