`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BgcRDALZRoKz7DFBdMev1/0TVRs+QKPjz6IlOtH464DVXRpWMgV2r3Pl/i70Gzdr
ABaQ8GHx1WFZnXV4OzaCEUP9UBD5AhtMU52F7znBm5OliQDye30N+uUG1iPlgNjk
ZiYzHEmMQB+Awl7tnoGc39rij4t1455Ral1lOvxK153rwbQnK7P6LITJ5TZgBqmE
gQMfEE6DuIrL+qYNIyRrGH1uRsJDjor5RduzzUW28a0CK1Q6+kU9URbBtU3aNauv
SV4jluuQhQbozzbxdFX+Gx7AgjkRnQxEVG0wDAT4Y+cDCtg3SJ50HBRhKgRJbdS7
eeGnblRcW88APokBSCzBF/v7BZ2hFxKQaldp6VW5Qya+7bPA/2+C+w9LJs/8SG1X
DK2l/YpRd+W8C3ZRTFLTh1fEI2QXjKAF7snbco2esGLfVyvTZpnMyPJR8WojGrD5
6sEWAVyEYb2QvAM4ll6cTx7R5rOLQp0Q1Zxaj7vUfPCtTsCKu9n9Tu+Yh7f4To3U
gQt8Bz5dAh8sFVj7d441RNaXPQMRRv27os4J82Tsuvk9Ynv+8bvZ5EWhUGk9/ged
dwlDTij+gp+WjAKoK5JIx5SFdgflkM5SeaW019ZCX2M26aqa/FqqKsnkaR50GVni
R4tnpUfJWW7s/lgcaHH4jDNZIxsjk4nnekGVHVP93t+KqTvan7ylZPKll97AnYkC
aBNRMBj/OzW3qgLnT3XSa7EdgnbDP/AhwZ64OWKUo537mWdbofFxnilFyM5Vvwll
+urlxMIA1wLQylWnkEdnPCmiR7K+4Xy9ztCAMd9Ugu5aqvse7jGBcR/As11E1NZ6
lMlAvrIeaupS7eRPYhz7iH5kiZi0Djh+GanZ4lxUp/xgsz8mMzZmU2m6ISJtPQhF
JIpWXDPs+TfVQwcCqatDjlHzVPo9125G6O2mDFfQ3BGu0nmvjC18UIbt2dCvkd69
c7gzCgm7NHGXWmk/96oB+/6dhC1KOxdNt8wLZp+Bced1oXfsW4NvOI04MNQNZbXI
oVcOVaMxitQuhV6PQtIY2uOQr4ffUe4kJWWYSj2J8vaAbvUGxm8Yj+KYmXAoPD/x
SnEjzLnSueaik96zyTuSTg==
`protect END_PROTECTED
