`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mfMCxTlUHUHDW3Kvq/TKej7vcULnvhq0tjSfNswOABtmQK83ojBBchZbwExsrHtX
A2JyUNVZJbBmjYiP0EP06pxqouVtPrNGCW25/b/XJWadmvHxdVciORd7t949RkEd
I9k2VU/A5ZLH5+NZc9uZphkSJw5uRITaucs1i9wszbS0bdjuRhBfEHc4QUkRb6EO
IJI5+NnmcIgwE96ssBNQJN3xuPi+wd/Kvu9WjUJgXJdj6eimgwYZQnXzdt4RqTUH
yi8oncGI4h1nfoMd6lP70srSd9zy2UsoDEPGJBIrkY4WFBjdSlWgQGaXjHMFiYQi
i2JdtJe/gCWWB55e1ShRQYZCPploHIKR0E5p51nDfo3KCv6ahRolBFERI5VG5OP4
wFRB8cC78UBmqEGY/E7BnWBZtHlx4mAuhfjQMWeGnyG/8voQfBGG2BFaXGj3yWZk
C8OhU22Xfp/J2xVslN2AnVix9nq9TzH+rm7xCLSFIa8Y3fFfj3inR6CGr1VjE0Fk
9a+BaSVxoQcOUY+DBkoxjgO+cR5lvruEx5NS3p/eQcXFouQB16HTZV06eCzxPQJk
Uzcva5wkyx+55zMCXEdQkshVHAUci1KrvfJ3wOYKwWgTybB6hASAoRuyZtns30R1
wv2JPAZwhUi2Am6Ak532xudCBP+XZ60jI6qfBSnlNDVLGeFhxuGJwst54gV81j6H
805xO8kR6NxxMiMUXHcosnJWSatAjLHAUTVU9Nz0KsevFy4BAE52MmTI2LQNjAgc
WBoyIqn4ICQppDtHSRQUSbOlO99y44h7Nc4S7e0/NEKBK7lNmYPD2Z8w46OollAN
SXnneJoS25nAGnRn/KG4nw==
`protect END_PROTECTED
