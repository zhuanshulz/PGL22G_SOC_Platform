`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GR7ktBl/NiCpY82hj78PIaAHNM0BG0B/07bs1P4CJiMr/b8f2bN+lMQxO4kXrWyx
222RNjuQjCtNQJYwRquhQlESczDtRDJ6HyMxrP0+Cx6HFsxCNHkOYxQvm3hrAR2Y
xhVLtfarKkYAf5+A1V2ugozt1MEzUR0p9wpNGF7ZmMmc4lmlNaLPzLBhsgNXMUZC
38IEyekA0URhxKhjkulfq71aXYZauJzLPtdO3MmN259Kt6bwKGqTp6FeLXL0WvcQ
pKlY7Bs07RGl/frgt9CMdxffYL2XFwLcqK9TCrDABQqRRqRg1QJFGxC6iYhPTZFf
C8STYIdy+sYEBc+9K8YlQw==
`protect END_PROTECTED
