`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkc2gG553OVS53T4orH5DKi4PRa56vNrW40WXGGxxHLLqrYVYsAaFYP2mhT8oVaC
w/IY81H80/2cNqpXas1nZc/3WkGvNIhWGdyPlr9RM9kTN7H2I4dWy4R6V/sKjrzV
owvRp9XQCwpXz1E4CIbXFJgDYreudHCDVi88SLB30NCAxxbuY6xUSsWwkad5nZyB
uuHurpXqpSR79OqI5ZIX7gbz9Io4C2bL6WUKPktBg3oSHLHyg+yyjxn7hehHCn/A
VNFDbwP0Q6EG6ukZz/0PoQ+YdAzQiwGrrEH3TS0WqM1hsxsNZIPmsNfa1S835X9m
8nCLLoXuh2Uk+HRupLRpQ2Pnj/hyvggkwrEQ/f8sq2gjqYxOrt++n77qSm35g2ty
pnHrJDxgm2b70SkelQgKMc/CeiayjYw1hdxo2rbyJQc3nYFMP8oI/g35JPTQup0p
p1OdI/JUBn3fOxkAHwYKRJSb5x5eovCMNuAQo5lN1hFVxman+xGyq6E9yw3yMeGN
zJ5LAfjR6j55j5FZZacaMxyWnGJihheNCVWZ6qyw3BVkByOK/4XhycqyVokUFU3a
kRA6Ljo1kD+MlRuWN4zMXyJ1+gKyTSgo+qaabKw7q/VowFaytgwKxK/7dTb064+m
hm06jC8csUXjUj91wrBVT/G+egD3b7pcGz9Ep84werprX0gn9G7GgRhtRlo/+1h0
COmlneZUUFn4rvfh9V6rIfIuZY8FRZIcGaW0G89YDTGQj+mOh0EScpST04V6KE1C
rlHAnj+hdazFkHvqU5M2bkn150y7yyVMmG9bxu+Jyb3t1BrLuliii0W1iOIH5cyc
pfyS81Z/LeH8m6Xn9gyDlVWKAMBC4qW5CcNaFedmfYIoUTq6o/GF0pLqRVHXLZ+B
SU7DzawSp1Pi80YWiEHYvksYSvYDa5lxM7mfiwLX+7h6gS3ciiOIZnhde43CTK1O
vCDKHGLutGLy5LyAWOk4lM6TTBT3sax8QZejWp0yTjfuNEF8AeLqPcw6DMOzq/uD
QgPpsbm5k8vT6ToLJgH7kSMy0SYR5eUZLIyiXOdUaYv0KErjCHkVI1l+UV1CVVCM
lXXaau5ClwV/sVMh9OQ143tjaY91dG8UvWVKPJJb5u2Fr+EGEe2tR26LwEPWD8FW
Riz8kkKPWnIokKg2t839crLAqL8aPRbfbNr/lTiHX2b41o0FUQPlPerapo5bIRsN
mtznb6KFKJABUWjPULwf2nDfaVCKi30akkxq04JMD9tH+DnhYu3BTgsrNKWpEeoU
hqCaIyWaYCSkqd51q7ccC7hxNFv1L8+3gHySinQ3gjGM6XcwGtMBWiXwjagrKNnR
L3gg1UjFmeRiC2XVibRQ+zH9bNF3PfGguoedTaTKbjERXLLbQ2lKfz81996XkHfl
ZgmJvSSumhalt5LWkFXqB7QwY2aqMcZo8ZunVfr1RwLjxK7BNitXEb/BxFe4xh1O
aILqVsmR7huR/dDQ1c/9GtB9Ggeie3I+3+NC6lKQOkOg3T87LV4WDQWxjtXBj1T3
CQW+k9u+v2OGqMfL8S4hPfjaScAdErqIkqZp8Y+QJbIbTP3udlEIE5Bxys778e63
Kuv+hZaG+qKfUvO0TPN23z7ix2iLzn9n0n/xvFmzBxrbRJ7O0hXQMcytzLCBXkV2
liDGcX041MvzUKY7Hfv84ywEJFNrOrOwjpB9/z87KwmU2GfnljQfd1+nKj49vjzp
WO+tatRyd0OlIbmPln72ThgrZbn5Y2wp1G1wblHBIuhXjh4Sw2OEaHFNm3GsOIYR
DV/w42tNBgc/h12u/7EOYgaEKlRDxI/AVsqkJ0a99t2ft1EZLwbhdlJ/5IxhNpqZ
9wgmLGXIdyExht78Uo6zewj+PRj8L8JZwci/7nCpvjCEbIRCMECMHi13sXH7NvkI
kIvClA3PRNyrv3JbrY+NMgsaHIJLvXykhbqUng2JshBZA4Kzn0ewTcM2gqOIBnZs
8LVsGadVUtdCaOb/4XES2gLGcDhBz86p/9kGkhTubqfChyf20Pw5HQD9nUm6C1yJ
rs0HWKDWOoIQ5xocVBB2lm5MRK1KIvMP7qLJ+aHEEvYaNfa4zdS0Rpt5puGeWGhM
idmiOCnrmfLts5uZeVpZMJl2jLEz2KtTU0j5tsXrveq6tuiuG5cQdI1OJoM+kOiI
h6excG0ArgN+OGnTm/ujC8MSw8gGKV/wzwzN6R234GA+oh01030FT/hITHgvGoAr
n2F0N4b5K1+Wr78dT7hCDGBWXRVLCmyvOvupe90Bq6YiQGD82EkmIcp7y1dcnyft
wyiaPa2s8GO2O8DJ4XJ/NQ8I/5i5D0BKkUmsGF21AogNzR+yn47SjphiKgc1vAqO
XlOAPGIcrgn0YARdVkqmNmh+gzVSpiY6J/wcwQ0LphZZbseNONM68KIrf3L8JjQj
tB2n9T/p9UK8tVGz9pTbCbbUm19teQ7CQyj/G/OdxL3YeWVDmzt13m7Zb3ToEohN
hfY70xBkbRxVAxVo8o0CzvwURs/NFKNxSh9sfAsLjVPQQ7SlmQECqIrIPgaQpe2o
JQysrR/OhfW49eM51k37vTH2v71KobxPebf918uMpj9ZVoO/zAr1uBr75qHHXr7j
ad+RFNNYgKgYkBggCuAq/sodhEKw3xJFDOssNi5UsKLViQ2NECqEBPUWMIQQH8EQ
fwmoizcgBlnnoQJV6j89WsEpp+FQq1o61jt77u9h0cUHkKqudZQqvB6KkLq2AIK7
fR+Dcv6eiYoJP1PYADJ3eynz3HRtax6r5WvRRy5pGRSvePn8rlWjunQX1QDJy4Lh
Ajof+kcdykvnopE7Voj4757Ncc4A4F37EmNke77hK2MM3Lm3OLUnaJWGT4YSDaBX
8KZ9Yor+dl4ktXT3xwk+Wj6qL/cZUFjBMhjwSqZgvWmE4E4lkphV400PsCYIgVZh
xLZ5BXz9h3tMjIAr18V6J96gY54bimb2RdgcOthzJe7cJQzZSKlt4Rr8GHFvWMyk
unX/ZsmULHFqhepaANJkXKKXaCdYcAPC/DtMZlvUmpT0CTF6YYuTwP3GnzeYvm2V
rpPirHqwAhhZpSmJD46YV+xrm9iCpfEW4IlIU5QT/iiZpz45/dqtn6nTsLRRwIjX
IhyOrGj6UnCbgPiyc3VftwLSyt96TVispr+8rvwnH84a2lh3TAgZt6fuuj5iZ9I7
tUTbFXh7/8tEoe7YpEjBhls+PuYcysew2r+QH8bWnJ2+jp9JXfyDha/jIRMP9e74
TNcSIsAbreyaHUi/7Ox8iA7Vz1Y2uDrx1cTye/a3B6tnGig/oudMY2OAbcmhAX/E
VErEzMUEImVBhlmmn1uvqgpWrPJsQnYM2rgdtkAxQgIhF8S+3DYi4FmXdK2iybYL
Au0Anj/bn+R/OIlbZplG0cnd5ys5Gt3iXxftk9zCQZcZ6X9m3/EtZfKunf/ri4M/
7xm9ePHebcY/d6K8/jSY1mLShGQxbOkVZpZG+Elenpvf+xJHRNMYFYvb1RKPz3S0
DH5g3W1NHd3nK28IJnQUS98wp/op9yarYRFg5E4nmH6G5zIbt6jqG7wnfd8ioQ7C
gb72pwLBrIsKOhyCsx4WvcHjZdr0JVfIxD2vPvlg9KYgqhFhHDBym+vSyVIiNy85
q0NhWQMvRCHP6Gng+djSqYMUt/heKHu+AKxw/E3xanXDfFpVtLmxr04hMThOMS+i
Y+DZktLedyl8asHqQlJAFuiuRuo+PLJITkcbnB7gsnlgl/BR6xh2/Q7U/TS5rt89
otaQkq3HSX/uHCieQVBFRkUJO3usMUmfJNkqYNUpKTLkOsIQQjIH1ICNI/8+qtLW
OezPMSsle5vmPN5S8Bu5UpNb9jj86dLeGxPggw13hT9Jxht1q+3Iutm4RlUVoyXU
JEnpaiJl0uBe1rg5+SUbebCy9GiW6LqArampkdmSyZVjVmT2aGLWTpuvNwrCbnK+
NAC8+6ASo8w+lDtCSJalLqcT1eQb0bTd/2Kpu6cYGLc7k/U3+lE3xBOkM+I3U0C9
NHeiu54qmClUqdaq4kRNMKSLpfbueHleKiMMXDBmCrn/sh8BMQPqW4okZ8JYdT6H
C/rKaEdNeS+1JzkeI9/mHp7j84qHERiPn79Gh1cpkGJXqt5uHoLlGJJvuJbYUaqb
f6HLIYyPQf6QE/4YywE9HHJUasR3NhcpMfJivI8e0B8vCk5h2DpY1FFrVRH/buIX
L7S2AMdpiY1qXPRNzKwRpdWT+y+vadDa20S1uOQZxcDuuLJREl6HMs/NiCnVNVnp
qzjsrZg9c3SMsyloETOAjCDl6U8Xzpz2TpZJsROxsmHSF1R3riQZRa9j4Iill+Pc
OslkJyg1ogBZGx/Gpog/73TS6yQijt+2ueIX5qjhcArMLe8RBhVBlJ63fLCxvPua
Ur/RK7rjGW7UnD5sp/mTdwO6vzCfZHbL3feky8MLJQhVItJXTAIFq24fLyp4Nt5X
hlJGjGL2mPzt/Kx29z5wmshPp6LbC41lBRJNtMOsBCj5MlFbcG/Vp3CJcOFgHlPc
gFJ7LmBLdVEx3lObMVNOL9YuNlnH8JGyaafd/uFDVsDkqRIqDCC8I6W9Q0xHHhC3
QP/KBNjHk2Z4q047Jo7dUM4d9pBLSxb/emgdfrmwrLY5KsPpKbrGx2gGmE+At6dM
9BFrS7yCrC/b6fZw0jGxSs0mgHMPYuM1cdAT4jpuyFmXJEo94dVTfe1AnfVoh0qW
wAX4dtzTwqijS96+UBsvPR0s1+QyOHfP1OZpQBqs43GlbeZnFPFGFZHTKD9o/VV/
ov6x8P76hgjkD8oN8tKpcrIdq5IjNffi0Kp5iTtb1SjI1nl0e3AFp9lxY4fddZ2Q
62c9nzYW18KMjRMRJe/Zenkq8IfONOKks3zRIZMRllwXjnPufSTwQY/rJideYp/Q
GLTr6cGY6Tk225ZzaXiHNi0RjPqMFDHtCb37kGkRUUjply+Itmg0OXyWUglv6MmF
qUvsuxb3MhGHCT9OvaK4Q+zn6QSz0iXX5KGGPkziJNxOe8Hlkda2PVmGHa9dXVbd
uc+QgPmxn06Pr4B5LL4TSfdLiaFsxCsLqkKUrxVkXrK/jgePmYZNFrRsR7pnpXSM
xnzrTUe2oqH4Pe7RstZPBBu2xq8Jfewtit3n4YIxl6OcCcmVeselTnmw+tugeSs9
9UGvSQrysnLnoScQ/SJeuyaDRDLfeRfCldvh/V8C8vi9K01csRHoUuHWpOk3TKQc
dGTfnYCLq99g2ZSrQYciO2LTbfVEz8c65f0tRKCIgSX/7dnA/tGmr3MjGeUmsZfj
c1T7apEGjhJFRvVj1xamCupxM9fCdNvql4v65bYFLrlHZ5swW6IUeEwPRfCd4SEg
y4bmUJAZ3oa6p3N06ufVLZZxez39StSySEn4nKSoq8wJc9cYJ9kCVq/kBJGIj9bW
KyWfKEshMR8wyLMSIHpysHGZCgATVh0uy2IiauL5DR1YCPq+POf97CfOT2oLN0Gt
BDu0hvdlh7KQQ5C2XjUvn5PHCbQ2iRujKYA4zzYOQQ+DzZTDneo5Jte+ygT2UMhQ
4oF8S45B99IUR6NJtKOPquP/NjbBsd43qYDP+LJXvYBbNbZpXfNGdmEsuXJqUspO
1TqXI1xw30I136BBUQvVWC/iPwmkFZUSRDXZQIGtMcQ1uh3mNuGPP4aWAAr9Citr
iqt/WoPY97RfwX3XucNdnreIo4mL3MHJrP4HDEsS99TlWgMWHXIh/QL4kjgKgm0K
ueETFNKnSUWnEYHiT+mQXOnL9GggHxVPhVZTku6VlMi8zcv4OJHGnI+Yom2fkWga
MJ8Y7/VupsZEsbfEGK5FkFti0OzVDgJzeLqwTbz3R9iwhhzgxZ9zLkIqHBhgZpg+
O4dv95s+9UqqHx+WhW8fST28wE+Vvfcdw2lwv4NGledFnJw/P4nMQKoVS+xIVC+H
4UghZWQg8jNeq6oehmgTOUxJwaeUiIZKU4CfNXPsk7eWt7G0gCKIdO9KdUqQqHxK
Abndid5WnmgSK1f78BM6EgXp9gL6UMOsy/ZCW0A4fvAdqHklYICUp7fBH/62gYZN
GHrg2JuG/6rt0Os+zT3ePQ==
`protect END_PROTECTED
