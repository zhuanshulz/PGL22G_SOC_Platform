`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPQH9mA74DP/8tqPeK+LOy9MIsaOvgHIi46OCsy/bSSwWybtCH5u2mbqR4zx6jwP
9XUTLvAVYXP2xrpE89qhMH+7zCjyFjLoULKWJ/CuEqU3ZMxqBnTs3ZhbRHuNFpzc
tiIXk+cEvaUgKEOAFKlz2Gnc74ITqXUd/MEtlQxQ2DFDMaQ2LOkCJmQxzazjbPlH
1Z61dAidXqaRrsik8Cy7q19zWEvHJRoD+39J5vBNxnSgwrWT3FN3WkBDyqrqVece
yYImH7IGTI0frxbHxF4SA5tPoy/IyOhyEgrnb9EY4ky2LxuBdGOQ7z1LymEtKbV5
R9RWiGtA7R4qZt7kax58jhT1EMhQV4QHGP59BCNsZbrXOvIuDmkAx7udn77pQbxo
ioDJITrNZ2/wV/oRWCm3ovCx7LJN5RTkb1blbkuB5iY8KuNpLRWeC9Pl3Elgudu2
4+cfr67yiEN2abOAPFWFI4sktXUAorT5GlktNPAxuyoRJ9x9dYy+XsA1T7LO71N9
sf7WzrJpx7kCmZbpVPOoJmO/BByzxD9eu6Ti0shcyIATU0wEIJAgXNgMLlPUnoRC
b1lWlJAQCHWVIlFrREtGv//Vosw8xn9QtUEDwwlbKT/YN/6E6B00a2DkIfnUm1E3
Ray9WWa+Gb5iHXYzxKbdoZ6gViiSthRVjqHBVBG4Kn0=
`protect END_PROTECTED
