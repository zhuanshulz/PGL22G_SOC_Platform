`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Q0hzAPvfpnNIPHXK3RxLtgFvXLc7tJMZw2XzJR5QTgxSSwhad+MA+r3av2MS5Se
cRWqhjwXEKDWfgA0UXFs2fej0Yr2keh9uVRrQgFcpissTf6fL5BMH3l8nFUCTZgV
uXStey8MTqoeY7MU+OwL7+JcqxSuFoPwgbBeUW30hfyA7r5yBz0d+nJ+1+iU6/8g
A39lZq/RoONf3/7xksld3IZRkno/rtKpQi9rBAfg6ovrIl1iEUd08mSXD+8dt/ey
xFbVjZINJQgMxSpPYYFw9zh8GMN2gaRKpgF0uzBYrEQph5UljeiJeq54GY+V9vUa
UsmtluTpTtRemz22MF1okHElDfNSqrCicCuBXQjcqfy7eulsMpnxYKv27X+n7asi
off6FKNrzEGJguZXLNdaloWAIlv06InuGZddWd17gZbOQOv4YV/j5MF4RtCO3dMx
el4fUSWAKT5HV3J5dUZwuTxjJwiWK0iHBGrQ7pZHxHk+WSNi56zp1Cr/rO4c1Cko
YObuKvk5hf6gIo1VKVjI4QzEGBWy0jUWeB/XWPqXoYD6kuAsKYwPy3Wj3Hsmr2pH
7PqFUO2Lr5aHVail5Xkzb9mV5Z4SqY100P11V2p6enm30PG0Q2qcTZzAfHx88m+p
gDM2gU6N84Bountj/gw4QRXAaH0//brzQpen0f7NBIQ=
`protect END_PROTECTED
