`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jk/EzeY0I8pnfDhDjtjt7+2yYrk4TzI/ph5fh18OPgZGmgIfsLaJXyPpZMHNS+FI
wTVsGsUC5mvL+TzGv/dVe9kYG+Z9KXxjRmV06WB7GjoZ6bWe1YWY68TXW13UNH0G
xjR09W290dudwLKVxEV7d+DmFIaH7ELL/Rop90qnpfxniCuhB0Zk0cE5TjJYPPbP
02jb+148yM+TtuFa3BHQ5J8Kyzm3M5L7XPz9WZpB76VHf4+0w9iDgYLXILN721vv
UwXNALcom9bY5vop4oeT14Ugpfneh3TndvEiBqnblAySEcuioiv9GlU7HF5laEuu
jPO+lI8FN0DliO4DuAP3ZRYJ9aVcCO2dnhDKQOO8YGYPrkF+5WmWKbju1+b/iiuT
XuLu4m7a7lWJGudZ5NGn2ATRY71HVjO/EGdXGD4IkfjtByanwsz6cXQ+hvjbx+8c
15xoRL1SA72kNRedr6oTTwVM57WWFxlUwAb3IiZV7WrXBpDKrhyqVwh8s9L67nYi
4ijd0hEnbES5umBpbfyedsGubPjcAq9N9cE3LsGnH6mW2BPuVevevdsRzRsjn+ZL
FGEH/Y3LwhXiT1SIsjf2WFkcSzCfUIUKn1+0QRsqU0Sodxtfk4g3R2aUjqfeSGA8
0XIw+X0Kajk4pPg/S1NUboTcnya0JPkpUGWI9q5OkEOUPsMnJ5zgdsOcIpDMeWQD
WtCjUw7m2VI6g+1Eji/NbYKvO6yezpaYyQBV5PBV6RpSoDe4oUMkhAPU6OuH0jTA
teFQYYzcxrFRkOyUMQkMGcBRn9X9FSXWczP9fkiH5xgvxGwh41uh/Tiog8LuZtMR
RGNE8sPoCDS3CbwH+kbxD0YZovEzELtMIyurCY5ZFBsufOsfltxaL+LMowI/VdFd
C+WIt4WGoVp6Wv1iUhKI4Y5O9UL1PnLkCDWruWO2BgYJP52HoAi44xs5aejC/vBQ
MXl3PnXY/dB7W/aPA1PZF9SK8Ezg2n/ysNPaCFxj58ytCfGt6tjyVEkIKvEVSTCk
+4rSeEmD/jh0xxqBEmAUJMl++yaZi01BOVK43E6INkpPx9EEJr/RA9N2Nw85COrv
JXoZj4SmBQMZKapLVgtyXFF6jdqIJmtJMXQD+AYYukSxPhuy5JeBKLadl0PHKNzs
`protect END_PROTECTED
