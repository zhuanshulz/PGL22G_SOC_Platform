`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sa8+NkhEMV6pjWCT0ykYmo9xEnqhFy4AjpD+etSTLjGYvx3skXCNiHI7e5WmCq9
+5Ng3vuaIOMcLqev0rCvR+IFkBt2mizqSVNsja7NDn08KJ6k9WrNvxK31Ezvzby8
xJVeGVuqeBLovmYAQ+v1Ov4iZvMcX46xFFtuHPtGLS9U9Z9oM3wS0G4yOWT2couJ
+TKJrweg/4to4T57XgehBOa+j4wVhXyGwXvs/doi9ECfATDRHnY1O3ruSQTjkSKa
ve5MhPr5McSN3XALwN4vk6aVXAF8XwxDIcK4mM02C9yMe4NjZm7HPFaDcUWMk4Ez
uOU1M0FpqhUqlJVETuPJQPgDGkOgyoyraWqMa1WmkUoGkZzD52PVdspBaDTboRVS
BtQO1rQqKgm0ji7eD5vm3gxIdsBY4pYVb9Z8K23bX6g9fJFc/79OVc1b71pjmA/s
RmIO5YtadiouJz39fLgLLhG6th9R9h5OYxMr/p7QYlfMpURNh2cOEZeIGrEiRxFc
x0Kj22A3mv9wE/YxPeT+YnLxSW0/ZdTdzmZzF/PPpsPWhzUQZjrdn5Kno4LEsSqJ
+tmV8rIe80aRyk+RwRpzXxlYNN7LPX/DviA+uDMFMkM/YKR4Ff8QXb7Xc7acXaMM
2qhWNn03mmamogNBheOFzVlW1ptClNDX1TSZP/jUk4kK99asGiJmarRLjGfVhywn
fzlQU97RmPLim6Z4dZ34dzAqRv1CFo90ZMeTUWSOpHJgadh9mbzksCP4c4l8s1L9
q5s473ZWRTTwYJplDtkWyitGi5efKgtvCJNaXnZy4TC6GGK+QX3uOHTWW2W/FTby
Ng8HpR/kdgkR0HSg0kgHusLIUc+OIpJQ992G5NTwDmcMZGt4EtH/2YBASjflRJOS
Y4KgPfFvtt9xBUC5o9vnFkYGjHvgSs15KhHLX3nbBsvg2wG9cZ8k4+PZRtqy8Hbx
tn+eC8Fbh1tRjkS+ngZOzDMAMNQozMbUlFCFAhcee8fR3u0idVOYROLr4RGr3c2K
7Fowybozk80SvCLGoq7nYiejktJ5yjEsg7VdbckZjQD85IpvCB3nCc2WVh+C4aWI
dFbMYST2Mpf7iYAKgmQ7o5csNyvZaZ7RfGg6wFJKs/rh4FDWB+B4Pq6IWuiFXqCt
4OUmN03UwsXOnEEhrMP2Ai+PWUinqyXjb8qEOiEW6hF/fTMP4b8Cf8vv40mgn8YX
2XJjSLMOQhJBtn1s6EceJeH/4JnhlOYog/q6KS2NILM7NBTJ17dIuFDQZg/ayDat
gW+3OWqTHE9xGmT6FoHDkuW1093HubXlMPYEaUY8Me9W/TPK66RbQoCaqzsoU80c
XznQ0GRu188bRG/n/whEnzIv4MIFP3ycO8mTKpy47QuS1Jvb98qi7Nykz1shCESz
bf/c77Bmt59eIAMQKB4AG0FA5VBG9Wwdgv20ilbO/Q0Bu9c9xDDHSCDxiOsoqGja
fhHNruh6vHr4+6vADfr/sIBC3zvRAxE6WtZ3ejDgWgS2TRbyxNc3W7dyPvrq50xo
qj0TpizZiRBOvwoa41Wz2JTr1CrcObc5YdVB+xp/qvsKxIwxzALTgzlss4SiZulo
aIwpr4kCAPsO1933puCrlwyOxVs1IOS/Efq12qucljG6lOcWfq1wVuEKlRXTaciW
+Xillqr/HoDe1RyHcZjQW6Eiv2LGPwfxs34ySgNtFxzZWGdIKdNOkgA9jIaKRvwO
2wnU1I7yfdTnMHGWosZlzKJQDHt1WrIv8GVKPdU3lJCLEXC/RzCI4nJKpwhhDMf0
/eHDx5J5J2k8XY5rsVLB3y4gbYbL8cXPvBRlob4Yg5OH7r9K7yCumGNZALQsYsdN
HXTc8sDMJetrsmhb6Sp3eA==
`protect END_PROTECTED
