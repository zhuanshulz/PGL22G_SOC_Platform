library verilog;
use verilog.vl_types.all;
entity V_ZERO is
    port(
        Z               : out    vl_logic
    );
end V_ZERO;
