`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJ/H3k4FR9dSqAOUz2AL72bM8XEUF0E2fKEeRBHQ/hs+3ERVVlAD1z8ocplDW2bs
qsb2K1M/55HuqfCd+rl8+JfaQNazlBoidS0yCZVYY5YdiJMLhQE3lbE+aDZ4/DkH
HlvVfgQ1uVtUxah2i8U+S+SSx14xHSAuPyxB/VwsF5nyyf/JIvRtyS5UZyNeGy1A
mfM/9S9YijmkSCcRNjldfhNAT1PZvJtW4lmsLfNvIRwCa1ivqtV8qQRZW4VeYne/
EUuaN60pgeWHFTEndhY6BWN/IUxJ1MCfyTU+DAHpHM1J21sW4Um+KM0Pp9iXsOi3
2mXk5JSLxjyfXlt/ZGnGPuCbw31MgERei+5L/57ypILg4SLmE8E4WbdiVwkJx6mI
0LtPGEXkGk3akhvicaVCE5Whgdx3c0/FAgyeeKSTIG8v0n70flv1UaWR5tmTvbYa
6v43h5lcaR30bGG4LeX6MUC7dxcjxODF4SUyrN/VbmOX5gAPTfvHEO/I3pVkSnoU
OiQDesHRNbsl+gFtO2iT4O9Hi1i2p7ZuD+NovIr8K1tfIiH69Jd+eNqMxiV9BTC5
eeHinCx4IV3FutR6Vk/G+4GK0IwKTpD+GC04RxIvettV86sPiCiAi9PG1H+8l3bf
ECItk7f7EaaimCSss6xeIBq6u+P1v41vn7e20A14+UXYz/uPyAR7bv4zmSdeCJ5x
xfM6iJqpiNq/V6BP6nmU5YXGfrFn1JOl+clSmzbYyB2SNpkRvwWExMSqZKU7ccDk
NtipIe4MPOTTJtt6ytuYLLU/4g6t3hlKEP5LvCIHdUeOyhSRIel7jZIvmwX84gfW
chLECppHUxHnLQ2zzxQ2GDabpTtFdSK6ENm76s2dIbO9r78yjkKCQ/Long+7XAoq
ROLTBHzVDJsEsmd/5XY4Cn2tCiTlneiehGGJ661AT1s7ox6DKrPhQCGwRpCcpmXb
vbRpmYApb2/kfWYstcGjzC21c1wlfdU/ILprCUKqlL7gWYF48KGqCqdGnkqcJXu8
7nxhNlP4CwYLwaF2npPXOMSMsxT4mcmpFrMYdhg3xwj0V44OWPnQJg5apAVziHux
PNseb+xSXNs6aiE+H550HkRdUfU3bfi+RWQWCyvb/4l9j4rWonU7RSBZtXmlq/T3
OHIH29uusjQ0ae9GSLECJEeAb7OcGvWFWvq2QB/ya763kVaZswRAb7oPWU+DQdZZ
P/UtJauDtGSZr/VmBnaM6T9ll8UkqXhfQKTSHDhnwYFrWtLe8XgqgosBx/4aQ4HN
uTi2uQMELXVvO7JgysTcszQEnN22PYCsS93XAAtnYzACqOAz6noey0KnO0HK1RwP
Uxiz3QTlh8lFnmMiHmJGrVMe+Rv3JvoupOZsbjNIRqM9ZBSLLs1Ym4KBJuwsmp6R
cNXxXty9Yp4xaE8WmcXu6RzWuGxALFVW9SQfMgHC59wATjX1HICd072Lkhw4B1wV
8LpmmSdzgQwKgdKWxD7q9nKojKW6MGYbKTzdU9vNx8x3t7DeHLDoP1H5KLaDdaMw
f7fd6INI9YGBml9BkB5E8KsFrWV7xEgUAU617KFc78YnTjGDNiRod+z+kdG/3UW7
DR6R4MFBfRbEZPAs2fxdADfMsiJEykk4n8O6HHYWjGSHTvhNHiZF0MwR56d6AdI4
E1l/NnXePR08c0Xy90ShJrZKCED/FaeZLPwmx/KXpSMwIl2kNSUED1qR/V3BYL6U
6LBt+gEjN+ZqH2T/Gqm8FGmqEtzFSR27/d11dQ4jVpp4yLgJ1Pkz9IjzvJUPQpJY
g/N8hQ0hZX8BVD/HLEcT/NuKuTAdxlXRbQi5sKxd5AkzNC+BFJdLIbdZFqUp0sJL
DxnEh+AFO+Bv7A29Qocdpp9zizTSVQeIcHxdS+aM08yqXw6fO68z42ZkDzVNkyyb
WGoOl9X0+Ab3AGmcDX2FMehYV5mNV9vHzYGsFrSGqjiYSPoEvfXkiLPos+VaknPQ
UKEM2LqTFHa5Ba1yaDPHBe1iukP0pVs7GoEJ4iI0zKlERZMG+5XjYTNqZowPU64s
fu+xpqm4t1gkRvdo20IvP4U8EvdolV/kcqBN/G8p+ByM/6r5+clh7pKqNcBlIiDJ
BxuePSSrb37r+BaJRrAEjTI/wQf0ZQtPreN//xbzdVUh5+1rbATUVk2WZT54t2XE
OhZ1PQMpPBlPzYZPGF7YVguF+Tr9fCUXTrLl5hNGe6+nabXkz2nznnI7gJSplvOK
h5a8QGWdGHRWiMHdvy+O02H/m3CzdoXg8k5ZNNCiEpZiQ9ZA0HV+Ob/X+XPlBAr5
26VI/D57LUHKbNjPlgJUTsJRZ7Wj0BkAlUJ4x51VJDQVAO6qohVQgWdrcLr2+DHd
iijNFYQoOjjXUMkz5yYkLhorx/65BuChsr6qsekwSqE1iR/SCuFyEz+KEWtpdiCC
pDaONMSL3nH71TNL60qY7BVb9gHwBBagvXz3EMNn2/Jtr2vfj5HGS6xPYg1IAIgA
UcYA0r7N+8awtYZymUVpqmtVwpkwZpnY2C02HhcmgqyfuVcHNFyeLhogipIMQuWF
iykATp8LWHKpTOFAaOYEDV0gzXutSS/fRgLSl28P0xBxFQsPXsBNItVbppsxMF9q
jlC4QFTEIH0DUvxbvjpE6jfxnHEfIRshNtez5UsQDpRkyn9JN5+USmlN6JYmMNjQ
cD/9eckyOW96yyIgnySOFGpCqSkzIoPsb25WyV19DXHGU8cTsItpd14VHOR9OE12
PKqEoDNhCbd6QuQ3bajt48CRY4UYI/U3qLfutgEwWGGGOwEKnrjFS6HKxKBNvdcw
zZ2bxzFhfEPRD3AEt6Utm5yQktiWIgIJUuTIvNgUWtuMQANul52gC16hM8fjQSCj
+S2pIHK1MAAejtL/B3Pif0eQyvGK7QvOXuqxf5IdLSPMrI0O8XF2+8FLY9jLMnIW
3IMirMfG7roOMD6Wz7cPQ3yN4FX9/q7iyi9YNrKshnT1BsEOtzi9R/eu3mvW1KtZ
MokTns/I5xSN3D2Bi8iI8VKIYtFqyaxRPPvtFmZ27dfwroqlDkGgbWB+Q0twzdDb
qpfpGJGdx1+p055o7DpL+KTV3z9G+ylvvo2Fn91MQaWYNnilu3DT/lufLwe4lTFH
RcUzwHzyh1JP28puf7xCjONTVAkflQlYsFFk2tKzSW/bePn/vSNOLOY/vvrFmK93
v+ohVr2dnr06dxys+Vb/tPUn5p5+z3DK4I6qSQF/qImVI2boXwlqyIcpEQs4ApkY
yNc078YPjqOXKO4kFP5jRuxHZke1d7qawbkzJ8Vn96ZxxWGZ9muoJZ3uVlOsb6IE
uwaRfiYsnlkxKr+5jSuMe9sn5X5xqdPdutlLMqamBLOscPxqpyX5A5gUIlErntuD
oxbUFqR4BgjtSH+OGsWLTYqOuwTGLy7nDyCRlhbgdonRFeSRTcp4AnHS/m97BXNW
xtmQxU4vZxDRzRgr6UvWDrM5odt3c9w5T/2u9b/WQT1WPpF92MlTRDk6eEiK/887
bbHUhSLTtIRLRWEm36TfclhdY9qTxGyeY+SwU1YpLvdHCMcQTduxArvSY5XWVbR0
9r6c2wCshiRwMslQo/XOkuOeg+Pl1MTLEFLU7OpJuWKHoMLZvlogb2YdTqgoOxWV
GSbRYRyi+vvm6RbPhf3CVoxRCh2L76xsEGoLzFaweOEtAnBMrQR4BmCgoMvbkBqN
vY8Eoc84l93svbJ+syqG65SZ4bbSm6Yencorv9l+y7gk7tD1FnU4yrdu76fhejkf
tWqqv9bRGazWtTLzQ0NPa9zVjf95SXIrBfKT+EE+HFHi9G77KQlfknI37U//2xa7
j2QGsC/C+c+4jN8ra+ssHUA2yCHrDYEaZQh6/JRUbIj4fQwUphV9AfKeGQYBY2cS
BVD4re64k7YEn6IXN7zgrQ2j5lIWcCZluVv+ZeeVnLe0/Yzu4MsDedyEgb+vxnWK
DdKMFIfqkpANxIb7Yq829HqxdlVtxXklGmw6HYPYzaj6s5bSioR6DMi2keTpMSe9
unoi8GPP2zT0HUs5HbHrbezLpystdG7k8OwmBsDqK0NMTjlm5P1aw6P5K1FircKq
c6lHRZNrXTwnrgwO12FnuCaL1lPAf4fzz0DmJGJAv49Mk6BFsHsVnrRDhaZiI31U
gkIzYDEW4WZ2WTxgAWaXYvKQUMaTDYfxwHji11HTGWG8ccwJTMFVSH/AmLmB5BLo
CnWtrvWIjfj4OkGkDl/KAz/HYZyZn893CIrXUx/h3PIsYEplD5CEGR9qR4YGWppo
cxW/aTPK/PhoLVXarQRSqA5g8zIrPeX3e5JpB2+0depBkEgJy8DSwt7vOgtm7ibh
mh1/Kw0eAL8A4wHJFjf9df8yg7L74acu2laiT9efHpKu8F2KmayNC/jbuIEwsqmm
z8qZlP/BR/ItfBNfBd4a0OYYJgXivkBHfNfHAmZBxuOcc6e2twC+EEVHb044F7V9
P3TNtxnf4kwnuQl7ZHndFBiICfJD2cVlYePz+z603WiiOS7vnpObOWgj8vxFTTtL
iSfC+alStgKd7DW4WhaxjBxIvpTPGCdKaPKYf+ee6Y+3bGozXUbCIpdJaoKzNstI
02lDxmzPQZSCvorVd7JLYFPZhL/qhBLAm0xLPPutg68VDQJt8EAawJ/iDw5JvY3b
jaH7ahnXBz1LORjABGyvFiuWjF8d3QlnU99MvV1UGpGNbMxT9TMmohLkAm0ueJSu
vY/oOrDx9gXA/yEebKE+5WSlpncEgN0BMa2+EjJLRqVYvR7caxYRAiwDzDzZhOTo
AxTW+WfGjWCZ4nclGhl28MlVzefCmP2ykE3Hdtpc88pNCIr2Sw7MPr7zfw/0b8uH
MXJVr9yD6t6zAcv3wE+SD77B8yhJMoHrrvIRnGeasaFxKXeZD/QB1wjgW2uew7Ir
ih7ENcCT8mznfaPxXTewimxv0/tRrLBV24vEqQrBkIXSLmaGX5oTGyaQY/yolJNY
ELsO6gGw7zd+oq24k0jkAqjc3YR72+zRuisCm0aH5Xda/ebhcxnhYzs24eMb/pQa
9/n8c55FluzeP8HNG8bq262hXY0igZNOag9lp/2YhPvxy7RhZH8VK/YF4gndK0Ck
sqErX6XkPsx9rFCd2p+bG7tpZjsy7ps8rqAnX5Doy1/NLcmpbUh1u3DvOmDmgU58
2Mpwt62HhXAK4rDLu2sfhpw1grDSsOY5GvawTYr6JmQxYSkSnX1Qb7xgGMehSH0/
ZzLT58hewyL1bvJv6UAr4Tkl4v6DW3N5j2jDCUJCbllEQmMblTUHobdQx9FcjttZ
IWjiwhI4JH8wGI8aeDQGeweqHyN1Looga+sr4v2u/Z7KW3pmpsb9dnnjoxPwIgzZ
9nKfA+TSlLTU5WV+8I+/eBFb1V53gePFHJ85ef0iVu3pr40NBWwwzFDPjWc6S4cG
HfYUmhY7ODtEF7UnRBg0EW3j42sLmK+CXVK9+ifYaw7h1HOmFKLT9ANAQuKx6uRy
G+/thOxy2xG0KO1YOXi1RG3gbYv51p6/2EIuLhysVspiNjRBmWRwvljL08rZvsJD
zZFUbWlprhg5sIeLs0Zx7A==
`protect END_PROTECTED
