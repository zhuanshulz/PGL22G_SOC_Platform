`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kykYRaSjeMWTHxxL2DL7xOjOXm1eO4oaF9rt24zkwFb/7cLnSXPlJ0xCc2I9aNwt
CJgvKCaduSbIafQi9H5ST+vI8BeKRZmTJlbJIo5Gnh7rkLUjrionPl/A2VWan0Zg
hzzN1dhuFkz6zQYqn6+cSleA1x+YWI8Qc4bbE6Pdrmg8cnlxpDvWe+gzrmgHgiDR
zl9Ut+y7oizxXtLDqr08U/MIenWdDKTOuLN09sPHmiKfH1yrKHfkilk7tgJ9FQ/W
KvdGHEDxiILwAsQqhlr2kLjxWXeyZfVrKOPUyK2N2UkpRjNujxOPWBcvf+iHmVAV
IxsS70pf6sK1borr+5UeeA5wpJk3ohzrfvCkGIcWY2ubUacc03STfB6aZxQHXiy0
AEXftsVLcpcFh5ZgJVVR/0o7E/qJRwTM/v4CGMCsHAJTtYAAU5E7PFyioiQduEJc
KqszFrsiWQ0+fK2QZvNTULEyhH+kphGu+SPzHBr9u7IUPidubTce/gahgbGowcC0
+7vR3qKjVeohLRdYIn/gSHp5vo+VZXvr7T5HAT/Kjk68QOJRLTHKo5ibptTR1RhI
Ry+saiXU8QBErOnAlBIJjujbXg3ylL2qOVK6gwq4MHTSySpDQvycLS6I5RhZAo4z
/wfVSPJun56KuAdSVUFJCwNom+6caX/XC0d0VzbadUFJt7TDW2JulEdfImiUEtHD
qXheKMmCWQj25UNbAXfjb1XBeW48qm8H7Il1kCYod9c3z+Tfa39MJn+0H9dDyJdy
`protect END_PROTECTED
