`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VU6/k8MtTW3mRIp/nShqHK8wHyMltF86oyaDYfOw/9PxOTmrzdZwtw5h/OchJVk1
W9IxMkxPoKcPf9YL6oQgnUd4s7e6QlWQdM2XQrVwDXFApg24wDh2n6THTVWnioor
m+ptZBrW/AdlwZKGlJH8hExqRtXPgpIIsqIFB04VgklttqxmjMuz5Gi3dzmN5yaj
2XyGrJ4s6MoSAV97xqm6gLJbY/KCX461DvCZ8Ni/SneHxUfjyW0Rlsfq62fWT9tr
FnsKelab4XMWZTKfp5MaZjbUPPgIk30yoawjwoH6MhlFDrEMus97LMYo3kuF+VLy
b0iAGB6A394OeBIXCALPzvK4KYh3Uxd9H/feWUbSKRPiVqM7kpxTcrMMBy9Oh44M
oBD4e2P3U1dSsRzbDOhhiVf04t2WwWLqlLu9rmNmTSIAocjXFLYMhD3YkLQepw3d
`protect END_PROTECTED
