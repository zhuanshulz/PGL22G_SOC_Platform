`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ewxnjhp6DFDpeom1TbbCN5WNldKB0RH+Pi7k5cJKDVBt3RtcQ7kq1kbThzY2A07
BlNUKabalnYBe98qKIYqW4G2yOZhW+v2J74o5L445aWxFSaDfF+PFgnMyx+0nvX2
8ud96ugVBlh8G1/0FrBOfhz/CfzoamTFx7wiIS0ROGszOb1BbP1wF+R8dFj6ZGPv
YjbMr5qgyPvaytcHxLtqA8AV8Q+VMcfWbROa2WY0O/4EmXd7KG+WFG0BvA/MEsx1
f8DXQmZ2eITlRZOI1jGXMv0QcSboYe5d3tMO3bgjWxsi0RoIU8VcPDk9SsS/pq/z
PUT3KuqwViBokFLEuawNqSZs1UI2NCn432l9JCQ42MzVQcN5Rx0elOr1tTUteIRR
INrSmltui9KyJZH4YP0BNzzqbh37Q2EyweE4WI1uI/RD4keFYGle8KMZYPsHUDjn
BsNmMaACeuuB2zEz+4AGe1ND+w795NSFcX3jmhGtQTb9CPrxpq5yyOiLqMvE53+s
Dl92lZKB8Cm04+Im3cf++1yKvlTXCnyrlJGpDaFFf/ljsvMcTRnytKLe9GP5TO/5
PLYalgP21E8dP0Kp16f18A==
`protect END_PROTECTED
