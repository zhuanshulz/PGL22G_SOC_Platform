`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vaKO59l/A3XkWuId+nS0C1gCwRMK3JcFZ5bljMHAq4S+JC7TLyEo0Tx+jF/hx2OE
8Y7b3qeeLtpO+AtVDlfPdZAIaYUrnPVjP/p7pQRmN+5Nr5ChTih8ZBxfORDmByIg
OmlNKY+HTAckoThF7Bxzx2+8G9w3xcE1U+KH59qvBDClCV0P1VXBfNG7NuhQgUBM
SnvsLVf9GWsQ+SUAJSjiUVhj2+xEoAlDHXX924Onimevz6dmviYmCbsCx7zjfThG
4sWOAV6xxC1iEPm+uisyVY8Ez15mqQFDB4N1FYwhaWemHbun+GA52/wt+Hu/iUoz
7Qb6MIN1KiXu2xvV0NY0h8u7a+4gjndx1pXzJ8qjZN3wQqGcDfaMjF8cVStzYkkC
yRFpVQV3EmUh59kVEq3osJo7HWHd/Y0bdusDlfozRbE=
`protect END_PROTECTED
