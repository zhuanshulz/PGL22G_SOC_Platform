`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dzkRJnbiD0uWaW8dX7BpFNz0RIuBShNpz93p792ZdCsu8dH1W0qmbU3Qvjhwkxjr
tNJ632GGrmaPUB6JLDHf7+ZGAsYeetT+AGMN14aEjp9Ah+xN6L/v4IFtv/eVNMJO
7mynjUznpJ1lkml4kgyH8Hbo8mvEIi7Oxuwr2jR41rDgtOK2wudn8wHhPjbLwJ1B
IY3q3M0WinEN/076qOrLr6yzY+Q4eG63n1SRUnxwA006bKPXfCtGXSaABVH09r0/
aLjZ1zWZbGHXIKqe37UsZfOCebPWmVyCxCzpP3Jg8sPuJ0bHTAct9Cb6hpFlK7Yg
mnm3RBBDO6oC/5Lj/3/EWiTyaLNGbEwaW33RrAq7dS/YlthPGHyFv75IvsTLgemg
maeFDfO5crca2PSTUcgDfpMTKKdBC2xna5++iqSdkJtfPjbynCEc+iUuwDHMYFHb
1V+ZrPHdKivczG17fWe15d6K3FJHEVb7sdDeaK4ofT3PPPBgv35PsrotMk7m2i/F
mbob0pwgWAKTp8JnO5Rl66zld5ZfeyABz4HSb8mDjcvxGkuW7vdPb3zYqwrGaiaz
44n0QyzeGDemogAJqVg/p9QBW25R+lS+AiJ1Y/AslekqKN+YUrGCYaaa4AfBQ5MM
ycssDj8Jo+/wOqxmbc+x2u/bS2QvRREHiij+WdbkO33wIzVIsBl01THnkUyJoscM
39kyeX8hEtUkm0LzWnIKfNEzJnbVF8+9rG5tf0bhSijQwLxfP4qC/J0gmqDew/qI
KPH8qOSf+UyJpOPJ7p4y1kZOHK0jGNx2Kr1AvOyWvG3CjVYFzMhSo/v+AwZFts3A
OuUcOWPoahDhY0DTDh1cFcBLRShVXDY0ZgKWkidhMODsILo27n0BK1ky35KFhKw+
ljpvR/V+RsHBGdypOAlp2bWq7jJBmtkwK6VEU3wIpGMht1K6Oiyfv/NPBx0f5cR7
zZLD2yToHLtciqGH8x/C3HKw4MboQDb00z/FSY3mfHRd3odR9GADDWYH2gsclGyD
IeYRP28vV30c0QghMmQKgTYddGl3vGX+X/3Ru3rn4Or+jB5acZLuv2juXL780jaY
1KdwRQSwIJE5FDB4tx4mcO1tBNBmRSDvHqXb+YYq2YjNSj2bRFOfh3NEJiwHucqJ
kPzDdYKosCDVpDF/fy9WqA==
`protect END_PROTECTED
