`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwCm6YbGztAPZMGWbZBezJcxlebGz9MZwtgOordmEAEuiBRHJ3irEZsh75N/piX0
TSuWltSNpLel5hf3z05ynctgziWvdlf3g+rh6W96bBk/29kT1JuH4XNryFy2KsO1
dRnBNF+YkC2dsL5LWUOEeoEcA/AHk27vUn9DYF0Qdxus5ZQQb1H+hX9r/qrSSqvl
J0I8XhTCHD0KVv0kMq4G5+Gb0QBGh94m9xqvZnJ0/rxF4W8kgQdKeB1pMqmfCAeL
OFmwzeOuUHsmJlvZnPJEwXi3VXasTr4FSKeDdgzYk4gxu4lpANj08DW74qQKuri1
cjyE/ixm29JApNnLYVS/knhQ365aW7me3t56Yr0L1028YbsoHb2vD6cHSBiMJ0G0
5o9GqrbUbloJEWuY5wOeah4i+Lw6lkFg5gZjNJyE2zxM2ryf0iTq43Qq4t5RwpSt
6OieSSIYsyn6Hlb6Ux5GsA==
`protect END_PROTECTED
