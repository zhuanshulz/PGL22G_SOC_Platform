`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tmz+6il8U77ArVkvzf7JCsAXtIQvL7bd0gg3bke1v/aHq0nnQPALdr4M7OCUfhth
YirwnScHUzUuLemzdE3axmJSh80QoCWKCTthfu0/kJZI7AzOQMnyKdvJLgfCC/4o
wAiVDCtKD4mt+NM7Ubqc2sSisuZhdD9djo8o5CekpiR+p2iqCVeJ+R/8fUyDMiNT
CW0FaStdBwAYvGK6W+h9z/tUo7sCTo9ouOCZYa7hFRmGl2fcWsSeQfdoqpb+uqvo
3tCTT85ApPlzur1tu2lLX2X+qQuvjXKR4ls7P/dgSmeasg+jyh3lz8P4Cu/YD4Mp
MncbqByy8o3cqVqZkYEkz7GUsL+H9wXln+VfYfehh7aEXoo+GbiF2ofjzg+gEnbQ
jFF55mK/jJP0KvGTve0LmBNFzm45sjOpGoQTBzUGEAK31W1LoMnGFn+mWJNE6IRa
MTvPLzl7qG6TIVfJAolvv36IW31sLJX8/4yD9zFGENtcmFbS6/YW8Ak4vVb2e9ix
uPUJlZruyHCTda+fJtULrQ==
`protect END_PROTECTED
