`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Xe7iCiWWQEw59SxrUPiNYdYvqSTXjHRe3bpB5VJDur8VDnivDiveJvei9SSb8rh
L9vgjgP8qhbsspl5cAe1dlbxGkAKkL8dM+iCdI6gLQDqjgxaUqJU9ppA0irGBuXd
Cm9inoXOzjGXfMn5yRau8Qxt79Fe49bsiMxNFuVcyG7YtFElZXc7nXuIZ9YPptQI
iKEP+ERXx+hh5BivhjKQX8vkE4md3C5g3skScgnLSyerTYlntaKZ6r1vWI9zLkrp
mF0pnwavKGr7IqFNv35MNea50LNHUbXzOiNxDCdFCJO7OFpf/e7eYJ3Fe3aPoeSB
G8xwUJiJC+479V00ZAYYdDSYc38tlKxFw8GOXcRoA+K931U66OUoG0fwVygLhElO
VEGNI4M5Rwl0vhhODKtYuHkfc/6wgtWp8U451YixW//7EPKrJQiP3qN2/hM9Hrnk
wsJWEogUIjekI7EC7RwXRS//ENoIxb/dIHiXFDDheD8jplo5nJRCIu/d/UQgOIQp
Z4G7lnZ3tiMoOrNHM45q6MYt4/GKj2Rzj+MYEKbkKDfwGMLBx8pRuNJvhjohk6R/
GVmPiEfjmRpKOiSfSWBzNyHJJXstB5HTMP19OezO782CsBj51O36wxKeJJSCNyoN
SpLeI5z7gSC38Z7Hk6a+pMAt1RrkHoy8hV3QHdHGtlrqwgxjXQyyXg+jc39eQrGG
qGQgHmT15ORhMKfbWpQGXFQqf/OSSmyVz8K0SpTxiCmAiabaPqvI5h9HNGWlHcDw
hTNxsldhfBhlCiUBBxom4f1E8m113EJM0so/j74N/FistBxf1cx+v4jaqFVT+bvM
4DNIaSh76z8+JTXUuMYs9DCupPe797ifYa2XoAg9GuRU+TJVAzJ8rpSyo0fiAMLX
`protect END_PROTECTED
