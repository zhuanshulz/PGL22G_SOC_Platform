`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GoA0CMgOoaRSgDHRYj5Eu5BgunFfP/7NtLm+WOzKE68XEcwxUVP6mX2/FWdioDfT
ftgth30A6jHGYR/03m6VVcQbxMT4gcZHjdUuQXNj/QCsLXXcyHz0CMp9Aw57PeHf
pcYu5ACnvAuZcAAoBfgTB/7+UxCqGeB0gooYnCxXVdYkCDMN3oaHAk8EfTfvGYZ1
uU0+MItEjHGaPhWjuYRL6H3lXeh2nYQSuSGNNcVxygnup4SA3NMojY6bDPzRVzYi
4UH5szhPAQtbR1dZTu53JKib4Pl+jOX3xtBDyXD6Jz47wZArTMpZPVyWiHqsIo7r
Q84zp9suj+Hlr5elVtuI6ktV4wGbeiFvMqRs/V3+FFygTqpRmU5Uk9MFAK2ISkrZ
TNeMzqv//wQFbK38d0n+8jRu/PMEo9QvEhTBFDbqqlNO+g80KblCTp5LXj8zoGiF
cnYjHTpVfVMVpXN68Df85RenXGB9Qq1L9rlkloU+Q7cd60qU/TtbguxMcwXs+ing
jW3EMfxcd8zIRScEDAymdi/CWf3eA4w5qtH0KhVStOsC2jtUIoxECsYWJU8FbVNe
fIWzGLgI3B8zqrO9UdyI+ipTPHK7vQ+HyyXglnoLWNQN8QN2yCuj1LNj95pM0MtH
PfOJmvzwUYnMcDoNVrdF7w==
`protect END_PROTECTED
