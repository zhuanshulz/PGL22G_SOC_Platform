`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KlpT9srdQrdmz6grZPJuOTB+yqs5hsRD6ZNuGR5O2Io3Iu8WmxqsmJrs0sRC6q8
4OBKLy+bhso///PzoAx8aFX9PFprAVkvRIIjUu/8kvfS6fGR+j2rervUJcrDcxeD
jEPKi7/cImsGCBUbXK3paZ/H4AUgwl9+gpvPo1mFMqOmgXDHLxYVyrYIfel7uzjF
e/a+j3DpYoC6hl01XQMTSgGTZmvF/xgXrv5QYCigIeXTXBh/WBEyiTILhldwEfLk
7MZjECLEYoLglGtWQnIzmZy25HgPcCLbV+GNM6ONxZtvzgAo0o/m1oJY4Bu2G8Fn
nyedF3QXM/1stk+VDvQToCneBHwdVbeDDIfk/xRBOYk3ORIiozcF/o4pJzBHMIcu
e/BqjEH/7er39l0ud5Ux4MY7UD3rX3cQuV7zgr/6ExgZhQ9T8HINs9cIRxCmM2RL
4k23iHyOEyRppG34qf7Gc+vaIEu6+GvVrMovzsfRiRJuvKWHsSZgsngychqzd8XJ
Brv32Lndhs49nHWFZNhmG8L9Vaen23tzHpMH0M/adOrb1xeKe82b+yroPL7LEt3i
+oYos+L1UbYEn/44Qk+YeQ==
`protect END_PROTECTED
