`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Neg6LNCR7vLB9gRjWWOTDfMMOmRqxxzP8kUeTd/B32d/1+zf7FgeNeSywzqBcrFe
KTXtyz+snr/SNnS8KnZqIJFs0IjDsyHjg5jUmmYNmZtaduIW4/lM87GF+V+Ie0Ok
nraZqHLQN9PWVbIZ4D2e+Tth9egIpnl10cvFDLXqErzZjXkg7QUDtZkbp88JE4uP
qZLJqL2ATLRnC41GsuU67hxgXcnsXRQZ1sCg4vT6Tk1H5u2byG5dl4VNQGn5zDcN
QfSUclVrMB14kVEnqt63eXP4o00o6Yvlz/LByjvQ+V2jYhvK9DXmCYpEu7oEmAuo
EwkP24dUuHC07kQK9STY9d3KBGMX8R/i+I679GUYwr8GKj9jK3yBF3FCDb0fBd0m
JKlHDGBVltYYg73R9TjeQiYNNjQ2dyppD1moRnFo4AK6HBelcCxmF36NMNtWLIPw
/hMESOzaHZC7Zp7zaSNBdNq4ejyZw0oyfgIIhIIfJ4AeEefJKUauthg29xqmIx3/
UTr3y8JlsFGT673nKgCRWrFNo9lu7pcPhf4hVt2NHYo8M3woJImY1UZ6v42p9+Ly
rTU0vJnc0tXlmispFkfOsQ==
`protect END_PROTECTED
