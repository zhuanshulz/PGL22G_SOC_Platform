`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rliiydUdKUqxbcD9OwyK0h0iQgx7d6nxgN+Tf7TVKw57rXkqKYECYP69QBO70sir
y+6BTn0mrUkpCTKEC3atAOg7bD+ujpGXWtfnEelks7eCq1SIm5tpjb+1OnKLpaZh
skD4ZaTYXW4xafSd4CkGkpYCRjizX8tG6oqCJKz1wRpO6OoPh0o3u8JwN+9j/9Zx
dLruso4Frs9Hugf9tua96zdLYTpmUqnTm0KrpVkxUO5SL4Ijr9NTckPkYlwp4m0m
HlVYs4gppS+HWPlaQekenByuxTtfF0MZJi4fa51MlS0kjc7HwiB3py1oiba6Q1dQ
wvUv5LKQ8K6tD26p14234NaZ4nUQ0wx1P8USNRWz2sCRR6sy1hv8hoMuQK0ZQol2
FZofdxDn0ZTbP8e9jQwAPSdW5KQ1/bfTXJNLUOrl6PA7D9XejwNCptzNBySqCqIJ
BYF9XVmzIASs2VptQeWxCRW8G+Qn33CNHDqI0jSzWD7jZxSj2HB2oF6dH8BMwMrH
SmWw/hmsIZu8bNh6izqIceLt7BwVK2BZ4qeEZ8rJQtoDyNHPfVZMp/8FgUKtNOvI
KLbU5fGzEIGeHg4oxrWm0r9anUL99gJFw/NWPpVQ023VgW6rOpZ4aef+EQmN8cdQ
gskLmrp1crt8HbsZxW9BLTvD69c04vOxS7uu1hGz8tf7DDVm+kHYQthgsvqcYChq
q8Mw421PicEaZOqsDfW+KWo4iRgdGU9LhwTRQOhtRjPXVlNey5uOcsW2VL+/0BBv
qpFsJiFfDiHR3oujwFo5mQRI9DMXNyd0whexTcuRENvFZVzuM+yMbYoPs2+IdEs7
+cuOIWy6+hDool++SJ8sUzsZQHxIFl/iyimJO6Cma1du7OfWvFIEkweyJqAJkrv2
IJ+2/9C2H51WcukxwXLkG2JJe236zZDvRrPQqya7LOmkskKkvjI0Cgg59o2j2owy
qc/HOa60FUiaHIYJmt0O4EOXj14F1J8Qbr28G61/I3gkk93VwA5wP4LhuNIPUaJ2
3/wFFX0InynfsbwICAo4tkfloBexP4FnQq4goJNSjCfx6cwubjdHOhigejIkARFz
JSrhKXlYWjo+22pOBprPkGX/f+vfwkjomVBtld4p+UNE716dlSg24cWTqojbv7x7
mCLiQJ9DlY8UxLBOiq2U0dQkmV51RByDp1yoRYDuVGJpO8G0MzHa69WVo4JewAyd
+vsboM+970ac0epMPjw2Nx/KHmY8sn9bw4gxD34Y2lIs0EaS+zBw2osAL9OsfCAu
atGBd+3xa11dMaQ81WlLa1WZBtvrHia05gQnLMHpVxs0bkceo5B19WribO9WU1yL
dik/dOsNCKyk52ECWNNg45AHc0PKBBIzQ4cx466Q9Y2sXiarI1A/ZWGf7M7DAzvj
ojfiSt7coI81UCNqrUaRSMr0z8TRhEj+AHG7r+3t+wgvLTRqbPSUPEBhTj1bI8RB
M+6yzhx4NBqEfBGs4pwgO8pqGumDFeRfHtxKjzAngvDvSD71CRSFDQUdTqI8d7sj
WEX6ACqMt6Py2wtm95AbYYPyEEQUWUxglIxs9gEaLyi5XFa8QfzlSvDcGdtB0i/t
NGyyx1SWl+ARGIJBj3B9ylxaNEN0KxBBvLZB4/ZwDdz/E8aKPG2D/DTEP74TL1rx
rwhgk02WM01CljBLmPW8grB5S4Q/qama/Z39LY9zSt0iU0nF6Bv8m3qX8/xyT9Dh
G9FNg1YEw23lRWvj2hSYkxtmsa7rWRWCyHM5xadj+rvoDgPRWueNo3e7/pjf/HZ8
MFDhERFWldxq1fZppss3WhRSgwH/xcsBnbbmjJpkiSUZzHVwrQOPFYQh65g3hJFw
b9QJ1eQ2s/4ADBnqyVMbtapuIXvn+Cgnd53nxqXvi3IVmZGUvBOZVDuKUzK7dISd
e4kidGLFq/KpeH7m6iEKuJJ0WHRXnLNY2O6CVoVfm4DHzMiqJSH5+01kJyFHixrN
111Owlp33W98f8JNMoJtpE9OuN2jQX5ZzvMdiR46lDVLMXe1amCWUh4AO2ZJnrB8
CRVRqQ72+TmE7+lu6mJO4vw3qamTufEEoyWjWgpUpq5zUXMtbrvCKEx5JMVmk01t
CY8+GpB0yU6ER/ErzSDHN2zXjw7gN1zvd/V8jJfIWkCCmA7HSalBsIzofoskT4YY
eVe5pMSpUUaWWvViV3XuLCKKNMJIPCTMTvEsbkh+zoGkhOMcjvUdNVQoS5xYF2MO
YOzOif5r2kvrsK4im0YbU4xOylacUL04WYYC8rJ97V1JZ0usM5K53pFyT1EISn3/
vA2rxFmvsFsW6lk6rj0arM+Y5u/hcW8f6ggqzuu3uSF6MjkEkcFb2XVLhga4uN1h
r3YgYqJdfg19+D+ScSRCyzoIvulzpIn3LB/YaRVAgczcNTH1XSefx3/Fdyywyz5f
PILn2jIFyh6AiQL01aJCArVTfGryvPQ8jAuUiZxfTtXJFcT6pggCDVkpI4NqfBxZ
wpDqpD8pSZQx3jfxfzqD6/f0eFH10QpygmnTVFo+y7N4W1FbBnJWdal9v95ROH6Z
nbDS3gRzHWs58lBkgFdkPSuZ09MYdb4MRqlu40K1YDL50Ot5i2sYDacBAZ5vKYxt
uKoz/iE2wf/tq3ij1T4eu7sjlS2ji85ZWgj3CGcw9g9mqxdb7iHCey1o4/IOYuKD
ugbZUza6491KMZvK5NzT1trmk4AWq/NsMDnCV6fFZsFzvVUZzgbwmVudwoLh7jOH
1yfmkrK8HDif1vOqiAUptjkP0mKXaJNT6uabpPf6V+s5/wUMmLr2/G1UgMSEPJAW
8QTk+6l9Q1PIjU2BVmMffG2ytjd+xIaOWAwoDIPVDLPGq+G4+C4hw3Kg0tW9fF//
FjcNVqWB47sgIXGytVjmCB7w0LrlMFW6bcy36Kh7wFCRWMkchYeOmvb6+v9x0Hxq
Ao7ksZfO58W/Y9nGUYyLMt3dTdjU5dNejxGhxiv0kMqDnWMH4J1KfXIZ9wsoTo05
GslA3hUjG/E6QKRzIiHMSsmqYrbuet+ueAyTxxHhoehFsE5NAd7Mx9ZnDZdY+ZQy
mT/+QbqYH/p/79kUElCM2qcqYT8XWcW/Y7lRhpPOx9NQgOYKPfxajDA0IC6OB/3f
y6UCerJOgNWufv5BLFp6fim3lF4xmC2hR3L37aGrpQs/KZvZLS0QbgLRy9o4FHDP
TUClyskR6E0rjuh1hkObrQHYm2PEHxdjY4AF2ixb3cKH4oEos7+DIADOEAod0jPx
mMjo5oBp/wM4RUYqBt74tc1Wo+xDckmkLaiTuymH0LMJvanDvG6G8Ody1cT58hjg
enTRCl9VMJLcWUbEyZDuK5sCyZQqRejKR71BYTr46BRF3Daf/bAUdVcroPM5hAGo
5P6rXm9p7L09AOG2AWZbstb8lOVDP/cRSeFzhkSK16H5TfHqzN8mmNQh1hC/rGHA
hLE1G2XlHemkMAJp+hclfd3t2o6nEh0vCfCjYlDBcdgvohRKl+jdGrOCokXJIKoJ
q4yPJX8vC6PUmMW5wqmKRyEl7H8tE14N9zilmfls6TrAOmwm4BuB5kg8um0hEexi
WeZpwIxaP8hzRqyfeZzjtSEz19PS6+XgnfCb4qKNDr3C94hGbMs9E+8jYcMhUxYW
gi8QLzHU82jikancIaHfrjWyclCmOUiXFYhtkO3M8D0dq9PBLTz+YGJvubd3aXHj
Lte5075uuUH4BCEKlNheaucYGiMSnKAOptYqwWgXVFBogx+6mOnDVxNSy6ftEKPD
OeHc4CaKykQTbpXg1Lrp7HZt4aZx1PcraUN0JtZopfQCMcBmxmA5ucI2k/bzCKPy
mNLDHEaHtXHWegu0hWOAkzEDY6FJ7BKcLB1M1OFQBWJVfii0o5RFez6XsZp2UiQ9
NfC7iI/mjkxDitauA0FTaaycb/0N3a7a8Rsj2nzzWK6iwRsEki1+xElt+Jjj2PMy
8Owq7kpQsViDqkmBA1P5uwFsLNjTocdegibbetSxHeOaHmisBVy16M4BORFF70jH
BBqqtNgmzfpQsTyVHyTQMKoBHUQ4o78wnjCjZZQ1AFiKemyoGuIp7bRBSdiqsTdJ
3NIkaUUAh7q+II6KZlaMxQrwYSVsGtafJjTJEu+9h0O9/wSeWpVyfwOIHpMFNyBp
gelVbK1fCSUDKxaLY965OdHf3co2uohCJYx0oEb1iT4bLLZU1x6m2Ja3KlfKlKoa
05b7BLDUkLH1ff+GnAhHX4pXR01tiW39rndrqF+dMQZqxgNxt2hKi3Krxe4LfLxX
9YQyhdWJJ7MpcbzaKbCqYwZD7XaFjyEV4fcwY8nsSNOxwuRT5uPjtbM3U742cO76
UoqTaUAXKsJ59tlnNdQ+YYf96qLqrgacmaFgActAJtCLKVXPEXted5Ac9qwKwMEv
y4D/3Id454olCicPymyqnraWtdunRtuBQbo6qqNwOlabNohLg4WKeF7H1kHRVKFi
N06m/kKcHkRwdqJDETdv0S8ybl77MXLTcnvlgSwqfXE618cMuU837eH1Lo/UN3V7
MelSVLn0nng0Yv7V6fMGdLtccI6BkF4LwdsL909pPOU6bwlUuyDs93k7CjDFcnIr
2yjHCn/vDHO+oat2mgcd+IiQzQ7wDODr4U23stnQJSM/lECeK8GVXumels1jhwOl
FMEJY6ILhyVoO3yFiYR49xBWsKGMt0JdwLM+pl/EnlkHx000lP3uNjeTFwBmQj6l
Cwmx+dPGqQYFiDyfLaKBX1xpoyG7KiRHc6zFvoi9zfTx01eTcVkMX2j8Z0ED48VA
w7JmPEZOc7dsm2T5mDw+kZ8B8jw9q6+3vcRjqukHYzskFdvwJYdRnqTtUNWwM0NN
n9SCThUonXpaCs10/vSniboDBDrEF30IkOBvM5+exrGVungj06dKjFEc/7WzKcl1
ONVWuy2tvXLcyWxY43PItukyDfNuZHXm+tkbjePZ1qL52UTaLU5kr2ukJsibuntq
/pjftQcJt4TrJ114h26G6JMnUAHw5BWhGDEDMbFZDqOH0iROUepEn8diZwcDY6ny
b1C1g4efKDUxt1d7QOnL24ADPLrG2E2hUHZIsjCgG6gKocqzcyPbHLlrjBr6qYk2
5NsVABKzpE3fM4uFfNmcDedGPlIucTnw1OpGVwVcF29qcni8wCqkxnTTouDGhwoD
MRS99K9ktpD5dUyENc9bdXJ7ikN7SmSL88alfJ83TuO9lxMx2eDTbeUxBHx9uEOl
+73BK3OemhBWVUTuPbc5/YAxlPJYSieSvc00CFoQJS6k/qkWdxMWXvMK1lhsHUim
hap0ii1oRUccfl5ahYEJUkFWwyPxKfy3BDC1HX9n1XV41daE3rgvZ+30EBQrXs8G
aySC9CJ4vN0aoTm2MzqFWOSk0uet8j/f2iin4F71wf1NHZ84rdvBE59wMilLQJtA
rmyBewAwxl1ttih6mH4jdWAT/JcM4g24wbTHrzYV8yM4iUif5KXlnvO4bgyho/De
fGDKon4V8tCGDzITp2Zt8QEdVRk6j+eGvVMg/dq2M2fXex4eocvmGqMic3m/x1Ph
uh0hKWzEJBZmokPkBrxfuPwXjuuRXZyV9hsH64wfRKsfpJZ9f292/lN9+0ZNuasT
FsAS+M6V+htsB7e2gJia1+Zy/CDwnAEFJdHsSwjx0lxim/cDv5IYMKMe6Ufta0T3
E3g56Gr4p+b4VVjnqhQYqqWNTpQqVK1h/yloZcK9xk+v+5ubWnYbfCos8jLYHtUI
23p5VVgiy3GWXCNj2BBwOZp4TWxWP0DO5aRxBtCQ1y78Hdbtp6GTmIXgzFXmhTie
+5cR0goEdV8yA0DNZmsKNkr/d7TLCi4MWFnzIBcDXIVJzQEJ8DPSrmHiUJhTnx7t
HjAQe83jLSl0GEJgRP1C4ChVOes5ogyyRFTCnRCXR4w4DtCpywrvKoa1Bko7VWdt
0p7AfPapy/Kr5rnR2Fx9tHdqXtz0SNKJZKYcIOryHyEHs1MOptoJwT+/H7THOpBa
mNinzmfn2uLqW0O3QEXZtwVu4r2tzygurVY2+N0k3yRTLHnVMnq2H8FZS+fC5Ytm
s17MqW/z8h5+cKCM9nTqkqgoaBUMF5K0VHEsAi5o3yRjmdULFKImk6RXKj+qJgva
3l/NOow4AmyFE9SdWhlcb2SJafL2ZJWWWzaVzQu8OAZxJA6v+ZWCvOtjDXz8vxz6
mGJx/HVqCazztw5rS1cKLqDlNK5M2GbxLnscUTJVX82fJlj6SzuW+XbzWzXKKKpi
jdBslARzLQi2cLSGNO/VfIygcPTf1VVrWcpndOVbnAlyKTu7mnjY7hpJ5LrPQ6Ok
g7+hrpeCJJHgtTXAjuQmudczKdQWb+sG91L2mu30iO8SQPYyDmrzBaC2WG8sFfif
uznaPsqmfU7mV9KXmowD9I1kEo7eVthzTU4d2AhB5YaisLN+gOVDq+QK5/ywuo2X
blVBaXYg1FfRFP7ngEID9BISVPiJv5+Nqs4p8aXfZcMsfazT8Pf6uo7Ji5Jz/C9o
ihLAlWgbCmEMh7d4KRvr/zzU+8GBsgxYOvUpEubdIgkB+7RYVMFwLXW0rAFFyQLi
34TY3zmhpQMkgM1ZntMN0rvLjjS4ElqmI57t+1RB6PiRacYMgafgL+3TcoZoK7bc
WgQ1RbUATvJHq/ZsMfdC0b2pkKY0WytOODK19c0/pceBL3+/R3z8luo70+F5Da6Z
n2EFz48ytFrZh5pbfIHJjAq+RO6Hq93NxwntzdOHiCjI+MW2QwK6pEjxNeb6rO8K
NoyagXwQiHkL3yL8ZCjy7STXf/bCH+0gXuVM68EiLBhi4cpj3afgc/eksdwo9LLN
UDuSPNWPr6bHJ6gK0uCsfHqERPY2uSu2IMEPHvzLHmelEMyK4LZpTJ3XsmTlKNlv
wJRt8obxrJxwrtRtNvIz2/37ylmEGeTBVnsceVtvsTq0TCkp6P3/r39Vmddpbuee
QG+8dzKaKTgaovTBLEWuWuBsRZrIcTu/aD3KFv7zcD0WCZB8CqUkm+bhWEaBk03s
g0LFy7wcRscyrDoJLO0r02aqGIHvZZR4C27+do3D4G1QK6Lw5INJmAIUfbadpmPa
nz28TLQuQHZaIdZ8l1c6jF+OEzaPISccBURR+Kb4ODLJAJ8bKx5hXYZPI53qv5Zo
G9THwrByijjdV1MtUmRMOUwXaWxzE8oI7DryfkKQDCaTuN0hTbkR4s+z531CE80j
MCq8QGzCnr3nSDT/KFjLUDnA8Ot0pua+e+V8yZmb0ZuPWhOIF87xicykboKiyoic
QTh0Eqyd9nHpUoSzP1DkCakZeFBX7ixJHeI10CUyNIS6KV4xjVPAHx4J7Ab7FqdE
VTyh8CjYlWvuUsyzuQyBXv9U7N6m466v2wvgP8ACjwjEh6I7EPqad1jhawozHNzA
qXFINIl9+P9DHA9AdshR75+5VzLxhkSv9XB/7jzCTJt0XNWCKxgafRXR3NBJkdzI
KFAPm4sxoq2kYkG8+J2qakoqxDZIrCHz0PBBDvBbAWtAtn7ACoR0eeNFyw5Y4mbf
zh4lvoiuL/SU+axDB+Iv4AiwKSkPLnqnINW3zNh5I+wgMHt6c/UaZaKc0L4eMw+2
sPR04bGXsiyaE0OGOE53jEANq69PQJsljx7ttxWGgEaNS/Rbjio2MP1RdTrrhoKu
BwiHF0C5TEvrWa22zN3jZ94n4z0OarzU83TxWluh/q5Oj0k+BWJfGdQywN1BPLbM
RfZw5MBBfr9ikzuARe+jYLC7xPE1QyehIhDKq6SAAzlfWhpYNEQ1h4Jy5HcTCwmh
NE1YxbO8TeAgSZTVFpWXksWFWrBLmeVkGf5pQhYBtNwUOlWsaBFS29CkZwXkZvgi
6wFxtcrPsOCqY+BEWeaP3LSHr6vfl2AK+QlKEvTIIM4AiYMiFGZqi4HiyOAq+V+8
CFYap55Nz7hYP6TzQqlRQEvmtQ8B8blu2SJNsVFGp68MIZdnCxooMoMgV+84rIc/
MZ1zxehKGEEBzUTrS6eyI1nR2eZCXA6fBpZtA+ccjiuY/FyKgzXwDGH6YBCzw2Bt
893q8mmYiV41t/yvXPLOFW5Gy8oJVKAOzchu00IdD7BNjxNtnGQj7pXyX2OiYIAN
nl1dsh85lNREgBQ81DFhP/tuqDMluzpH6cfHr/XcuP9zspOG8HzzU2ilDGc8K76i
k5NDhPJYZU/n5fvMA/+l3UmMxiCGU/cKesvEfi3ZjU9MCgr3A7MiwwuF7UV0JpWi
/l5/k1Hnec9LIEgizvidNsA5GOCiYTGWwc/ID6M/PXD2cpCbgGCxImdR7Gdd3P7R
lERbt4lRZLjGXTcPhcs8k2woPIdoD3tGpe5wVWpRUXW46vZOm4StC1HNn2FubgE8
MecVb9bd1HhJSwKgKh8TkfMar0BYGSEPUU713gWRBhEOqBATA8xD4eHhM7XWoBur
fZzcO10JIx2JPEsPuoW5n1QeVoVKrymiNHGhBf+QgQY3LfaSR0D6Oll2yg4C1wFO
e/yFisHxhHE2lj+Xgebohp64UdenNTtqlmUtnJoh2CNIZcT7kxvcAP30MFE8lVj+
5cY3ten8wdfhqAsGRLnBJM2Bt0Fx9/R6AATVIy+JS8jTksVRe94XQmXbIOj+khA8
mJ3OSuujfxLTyE3Bxv7ZCwZfqA3rpTWzTyVzB3i/eEH/DyMGvnKoAXraeEZ7Fs/5
6sPmyRBR2/p8ME82ISNQq/bB5yCQi9uOUL3/3Nv8LdFwcN7WUt+SDVWFnsqmkFyO
VI6H7Kjhp4i3JJ4xYAQ+d5KBdKmR8razAkRxd8vdATMryB7X9kVWCHXsc9AtZUPV
3AgSx4LqvxhN7jJfkY+SFRscetglC6HYlv7zWEdp5PzX0sCw9n9acNWXy2s/l49m
RBzhzjbKwJllJmf16iAiTKN3JVSicYMKjmFqW/Y5T7bE8ffBcogBqFxwtF7qaDnf
8qiLgxHazkhbaQCjv6I8O6hwGxQJ4VrRhvX6m+k5EtU9mP/8pt8LWqXpid/3PqVa
go1fVbQghpiF6MxlR8sYLAmh64AvRoG+8mHAgSmhEqbtJy96OxPJ3ZBVAXTAnf0y
NbV87NgrylILox+0hyTlQzLRf3gCHtNDbCsdjhTViMw1EV73mf2AZCqoLMaYMyCG
2oDIKugv8CN/MQznRE1mfmK2h3/RAfw3ENG2dUaLFOTqmgKThsmrc+oguD3CkJ8c
CqTEHRmqU+Y205cBB5P/YzTr6xo25pBAwGhgi3ZL6DYgTd6LQ3Be+86Dw2hLnwTt
ap/OPbNJChe9l0V/3XckEaqdTwuDeZPiVxsBDK9iTG6cvcZkPNpZc1GK5Xc4J3wQ
3MLw6ZxJm4QsXqzPnA4HlxWxubk2aNkBwqra3RiVp5CNk90v7ad6XxhAymmLpVvz
E16bR1qvwHL1ILXetxndG03sBTo2yrPVmfkuo2+EvnCNzJcCr9CnR1obylPigEPf
qIttfL1fSePtbVo1uiykjbWG9s4Wzx9SpgEhzbPHRvuD1Bm+KVtNMUJUom+ERXZc
MqxfTK2RCt1ZA/VmFY4KW56nLiUdCIdaC66kY8J8pIz8J6i9k45Koi6G5A6RHz/E
Qoh0zqwNKy9SsQjYuqlTnwcxVAqorPSAeBV0aQs7GQvh3frqO5rhX357WFBf9jkX
czyY06Y01CdpPl09BG8LLefjCzr9Zi8x6xQ46ovVvshYLJaWU8ht1Rqfd5RsVWAn
HPX0tY+kZAVMMWiOjmqxYWYLgwDg3MxGrbxZzFhaocT3L+2hX3o+5Hv0PrPHChss
mn1a23eDMm7eyv0BBOWIufPOXhlNV5iBS2xz8QRjGBe4sNQgyaa72OLfSBt3ZMY6
H3g4hIXxllrYhn/RvlA706EihTNufcVs45QV3lPbEpY7zjlCX2s3Q7egIT9umfh9
v/zoYqkF6w8yqFvg7ZxJqpA5sFGuvmaNMK/EzhoOd9U7eHbe4VD/wuow8WqIGKBk
OeyFe7W8mQiKN1HR7pY9kU3IylCmDDYbU647sflmOlYXznTs7ri+VNRaSX0ZTWdr
YUTdPPAz87B5IaN285ewa7Ma2r2e3VnE5U1E3dysDJwjsCmVg4wOc0sJDacAzO7A
KTKEwuagVg0sHHU2vBxah8aryNZjpsmf9pmzkN9k+X2D/uLjXhhwOGn7xe31noCV
o2TWpZ0G7D9oyPsXXuP3k+pd3a5y4WAJ5ow5BDI61d7HvQbmSoa5BVOFSLyXADOq
qsSbhvf3AGBCkgVjCAtr54v7Zp3br+2EBgRiRKD6g5o3gmPRbn2EIIOsxgrjD9rn
duqpVqF1+CYWvuJa7z/nYKEzhOOva9oZT511TJtOx8prhkxzIzaLYu9KWKs27aYu
plFYNA3zOmKZy8Koae4rKvCG1Ase4bGIVIt+uaQ4/srFEsGujKPVHX5qY1NSKwdB
dIbqwDw+8jGt1nxzDc0sEAkz7Cs018+866Tai112ykqevEK9WNIYYI+lfrKlj/Gr
UN1mraygmyIFG/S8lBo2CeK7VQJIQOLwwhUA5QeXTpyenzo3aHDp8FVg4JtJW2KT
tfylJakjOTwMBtFQt6O6xdnS+bGXAWw+BY0QmDMH7iTxXYsL9StHkuIyU+kR1Be9
rMlXPp0uGLC3yJZiUm+mo8J+3/0Jfiy3bp3wQABGysnUudtkDPvtdafb4BTdiX8b
UavPIZbn//JOufgDyQ2IC1s1y4j6Vi2ag/MA+g6tMwkglenh9fTdDMwHriZ9cZnV
pid/Q2F627Ar0/4eQZgiGrHQwcM3J32ncvbIXChRZt1nsgQ5lPzCkk1WaTOL5YCW
65I6LYr7VofswpPYzZGChVUH5p8YhIK4UvqlD2IGfCd4aOGWtE0tds5/Vwhh+VS5
c0GQwBgZ+XuFafpEQPm21LrXvB6V9FRVJbCICCAmQoda51Q35TxPTZb1LBBsDhy/
Jnx74oOPUz/Fvwd8CXHG20aEmFOMdeDBOnz1MzPwvlILvBv3g/yLJEivQCP9MDlA
8s4UaJChc9X6vOupDVKurr+uUrzYxxtfN4zN9WDLkIZQASZrj7XUg3Pf2fQoPwTE
6w3cPLdy6EhEKVww0TFrSD4LSxHXPA+WqHShb1ictT47mfp9huI/iDaHN8DRXuUY
Gap+fdKDnbHJ0xeDiUDqzOhmEcdcivTLDE7OohCzipC3zGHE8yTMxyndQ9nGheir
WZpFKWCh917X88XtcOnaD1WmWyKscSdR56hSz6nI6Kf3Or/GX36SyF0k7Mo6d7xO
K0cdPcIarI7itYc0T9yvicHeHGY9ybOlTgIwmsTE/NYY7IfdkcHDATIgnAcUoNmC
NQun2Fkm/R094cyj1BULW6WOle3lwDhplYmdLSdJrnC6aQcC45O4t8adzxx/8an5
piO6ZBVl/RZ4HZMMaM1UCiJ57pSpzx/QbZUeXa92A+etiDFwCkLHnsXebWSvp+S2
qa1dc0TgFJPfU3YFwaMGP+kmU+OQPrWysZm3Y6m0EcEUjYeI3u9AIxhJnHc7K1Km
H5UUwhOhkVKVnKHCxMra2qpj8m04PaVkcieiRSBixyzDdFsaAeIkM51v06zdMz9r
Kujm68Q9uCPFZw4WqdXF6lVc/V1EpIQQqzkiFQW8DaDRY9QUpHBMdHCD/VRPa0ZF
RYMkUt2+vVNBxPDho3SC/Rndvm/9fEHtx1kRAS+Gey28yXUPnPUFUlEwNIGWf43J
6JtwOCDbIF9MOjm3MU6DUMbKn/++HRh0G4h50G15oMsTptU5sJqJxM8b0vDLB03n
3pzpH6pLovmnPGhAqz3vIV4yfLHyI84zHvRiBPyTSOGYu4rZBT3mL9AwD/PvKdsl
l9X0ypvKhZVY2ES5NNUL9twcHK5TTfYJBqd/Je9fdy2lYJe/zaMEM8v3nUYk1FOL
EpxOBWbAgYqAwn+VGVYQhBkce+UCaVBg9zm0QiibJgaJONDRmGZmvnrxAWu9tJBn
Zx0xFPSMDzlOafP4/uh1OlKJe7tVzlTsio91qOXTgXp+OAA24SJl7RdImZEVMTSH
RXbPhJW3g/HOIzTYfYW2NuTrnosMvKKWNRx/R7kE4NVk0aah3PNnnv4PW/BqREwO
NKSNPxuadzHvWMoxV64dyXkdGxTQaO5kRQQ6cbe+AHSuRnJqdpLrvkr1mKbK4BQD
iPNvseFYAdvyHYoQPF52urbWzNcjvrM3yVlugTHvvKcp+HsX1bV06pwh2iCSqLZZ
IT4GWdPTIBmrYF06gdLnM7qX2OkXHMmpqK1dSSkUuUlEipaABlHK6URu/luGlPZ9
QLbUc/m1ntOypoTpaXl80nBDpMbP7H9ESihr0atM2f8GmZYs7Sow9fSn9NUQ0qGX
GQMF7knYcR+ZAT/E4MNk8yy6SrUpvMrMCavhu7NhwGY7NV1zCD3JdlyUlg/QIl3V
KTV6QYyRtuENKnUAwEOJOiQyiQ3yK7CcwA4Sdt6FRxbcjg98zZCP3mVYG/h5gn6h
nd5IrAFDTNKCt14WJgCWOPIAVyfjupldMoad8OBuNmnOgDKCSCapmPc9dIE2hqgP
RS0cZGAGeVV+oqGw0PspzJtOcLIMiHEL9heW36msx71WYVoDg70ZOVYbwQxcEKbe
Q9TbRnYEbm6ebXdtvDHWrXWkCkZbQkaA7qjUjEacw9cwzK2KRPQukqUI4Op7pI7B
b4Jago1lUsgs4tlu12GG/of+RO5uZg/0rpUYHvm7656LuBrywc6bexSGBEHGoAVU
hR0k97LiIWZRKiDROUbMD6zPo5K63kmmtGs1UzSXuazrdpsByZSExxJ3pLeEXL7f
A1h4QkvP+1hQXcmuGgrhOww4Gkke1JOLHphLNYKsITXqdvfsghBl42qf0dKrqLwc
4BtFS3P3H10zp4wojrBKCgvFWsJ3LoMkPbMDf46tJjYULS0Ix94YqU0d2oV0ovqJ
9nVyp6+jmyY4onFx6ACR8QjSgZk6kFvuIDgpRgCOA0uyM6qusdJVvmfGvEH7Qrov
ZohM8NqZTLnJHhhO5QWYGVjUzA5yIiDP8e+Bf0AKUaTUZ6k/lNDHv8trSN0zXrN2
f72nro48LyHKu4ZIYIrZ+L51kKydL+yd2S1mAV9MBOUjAbw4YVoK+wPk8g/AywMR
RihNeoeS+RzKyNj1uHkQjbRmxRGPv3/Yz+2bKfruA1oqMP/JiW/onY5IR2/29zw4
VQFEpHYkXGp4pZs0HMlEVJfEPdJl8/ctl7cpyVg2QJmEiLxhcNS1vcH1WvxU3vmg
9O0w3U39kDajO/Fs/r7DjuooKlqLSuprPc1lgvI+5W9PgmlVf0n/qmOa0giLsJqo
rVlk3UzLbqyMZBNdLT1Vvf7yBhCOG3jFvnBAzSpDYJYH+ntDRpvNticZ0EY28THV
9V/v6Tv27jgoXwBeMAv9JxhyXgQh5eaV3tCNGYPBiul6QFdxsVQkCKHlIiQ3SkKp
QuRsxRBz5MEJdpK3dl2sfzVJ3U7qj5ZZDEKurh+kSPRNG/1ymcAgFrl61DM1QaRo
PY3GFR0kaMRD5fAhpmNzEO9EdlQnDey6FAETcDixBRrK6A5FWFP7Rk17VeY9WXDR
Qt7RxHgaVKp8PrbqdlmB+KmEpIU8nhxdGXkA2BxO9nGsNIO/dbLe/Mc1DrzxdAP1
Jpr4OrnaGumtLZ1desPdUZnp8LeaPVf2vz5ulX1P/6xKfD0fZNosl/68U7HBDaMQ
CUbRavOpkWdeTVnoDn8Q2Fwsh7f29NBAvIuAsMFhXd0NCp+JUwUlfQAS8ROJEbwz
BAzIcnYE3uVHlq/u00WGHb2Ym8Gf5NucPBaXT/TmAvQKBibVLnKghy9MknIdEO9b
F/TDaM0hzDCydM5PFltIoTke+3TJsRRGd/5cjuMILor2K91o+PpCDFAr5VJNc3gW
NrVytZtZ+AEWMTfqvJqZGjiyR+67t+x+EEL7wJrOu/Yd56QNyIxTL1+9NBOcGrDm
hW1/COLlxQ+RqfK3NKhGR0GGJ7GvCcOMGgamModPKyi783CTWMgARyLTa4/ePg2j
ZagF7ILJwOQ86I5HI6H56nqVUQod7T3D3Tg+An8JwimV2og/Xw9DPxnXjuymzKQg
FvX3F4xSVWynaIstiOf6X71lw/6rCbEK47YhjI6AK0XCqOuxKbZlZwK/O8M3aQhH
2kSSP//5+q1JCt192xXrvZyv2rggvnuKLvujKuFH4ew2HhDxdX3YMevJ8imSCbB0
8InUkI9mNoZTbNeAac/tA1zZiMRhKUkeNJUfw/i16UlfZmZTEXuxoxRN2VSwG2tk
d/EWy2RreOlItECMLLR7IoFYPMsZSd8qQsM3HsTmqjTzdQFOMfxi3cL+F5S+puLs
6HfzxxgeVZ23OFN+tLgA9ZCld8Be7T6sj1kSa93eW43lFWeE87pNUICWIS3fM88+
hDWQhOCLLudOh+uNCWQS90lDVSQlXNPKD5x+htlryAOeQP6MWKvO1BmRhGbSFZKd
XXbQFXpbHkKtHkSpoNSAvSeyUlcYiwDVV7fNEoml6jqxIZmAwSiqg1RD9iK6HsXQ
RWQmmyrLVZvmz6xIQU3Br2PZ1B20cFd6vykPVFbkYmuBPKioN6ppIXQPq1sUeFw1
ItLwyPUVH2j/roHGNmdtANQA2093vSIAblJQv/3zqpw/WV93BlwTwbMOBFhlkakR
JEfXsdwITLJU949F2slcShdyJetwnSYLJZ2OLIklulxK0vC7z1Cd5n6D1k5nPUPW
uh50SRLF1iv0HchTgcqtwbZ0jYlczpapJxYQaBybeK1Nvs8bo10LSEchvz5rKz5g
x0mVvHW+Wny1u3LNsHGhrbUKPkP4Tc1iff9w2QZc8FFjyffTk8IcMy40+fiMcpf0
9Ca1LVi16tIrQm0Pcv9fb4NpuhCxc0sd2ADQ+bX8tkIojh1N/bV+g0+pQ8MUuct5
e0uKyDLkPHjM+pHOs7meyAMiJPxEtlzTqtHMhdnPwwF/C2+GJLi9r3ynHg7PfmIT
BwfzHukqG3pAs2y9El9uyzzeHl0vl9E6eyWkeIVxqDLyKW7kKdzAN4NqwNK3dbuz
AH3OQfD+fsIUEkBEDWW/KuVVuzp5hJccEY72keWTFZo1+HE8qZQcUR7spiMOmB91
a8fndRex/RT1l4/DEDp7OOKBNn6c1zuUZJ7JVGRsOQFChf7QzEJzUTzO9pAiiGB5
bXiYQP+x8Nfe+d2elATR/KPppCj+ZOF5IqlEVPyLqthFrmunkyRDGqfwIdkW6946
xW2bKOiAHjG2Sb7sCFKWq5LokUnVWQtx/gY13S1Zi1/vB2GJ0TWqOmOTsQAs/MX7
MlPKOSmFBe83JQj0eM0azJsXDPxrHWFogKJdebO4kIz/MbFsb1r2vts4dCgqeCR5
zulpW6PznGhUnqq6lri0YwWXjLtHVrfPxYF6T7UG+lePUpKV37yGYFJNIJN6fsiF
tUOJ/5k+VvdG/a6pPCYTcriDI5LWuywbpbuSRjFu6SCqRd1oLi4CyCMWU19CZR/w
zi6UjmnCCAOfZUZFGMVl6jVadAc4AYQwxz4kZMWvlnOWk0ZSzgmKf3VO7WET3NRt
OF3PyBea66YUtZS2GM6bMaiCfwhKz02R9vdyx9wdrAFrxnBGAn0Ukz3YLtDnLBzc
ym6gvv6SJWZXmcMn9aRQUC5fMVpOld9ZmQWqxg0D7Np+WohNLLQxaONkkioGrA5R
YP1CtTdJIO5Ir4O1a7RCdWNi6Ryeg79RKjHI3JRx4ENZcYtnEWxsPGw+LlCLygeY
vH0E3meVAmt+Kk6WQas9fTId9LIVldsM69xlJgRoD+TSVRTkCpSOAXoQxvCxt68R
7DyLNtcyrF4EvrNziYWUophizKc0FjatSWR50e9w1B1uaSviCa0kocPMjWiaB8iv
mebMkIA+3NEEhsU74BcRIclnIohpVrwEghbwvVQy3hNK3JmIVfNAgqC1C4A2iUoQ
1t2DvYCWX91SJsy3541rkyjt32K6xHeAGJFGKV5Q2r45CG/dlA5/XPb2LNtce4Wo
7+3Vu7HQqxj2mFs+G6+i3aCra53e9F6cpD6DWBkIAWMUxTN3qEFOlLUeDWFdCh9K
RFnhRXgjcbxBaIfi94kji1s1fmbcVKFhUTLQxzAAEnhuec7aeSY8QikP2oKNj7PW
K/X/G4VnX/jDz79y4N2Fn9ywGC7nx44koQ9B6pAIQzu9doCiYsHXAB1ZOLtrSdzR
kC8fRXliRZpO2vJ24gzoD9fL2LoswfIAZAnaTOyYR8IdGCflK3xc0GfjrDgQnEC3
b47SzHsC2Gf+tMaJhFdgi1AGgABoOTWT4L9rvSV4u/lyrD1e3WebjnIQ6AMrGCvC
e5JvpooXdETMLdIEFK1YJxgUSWXOVgxr/T61E02gCtG+SFSnJYZsD732LrI0J9FN
xuFO3rTw/I+WNoJDYL1JEMK8IJfr3UnS/1q/JEC6QolX+oC4lm9V3GIzX+cZ1HMT
tZ5RINspsRTfbSjevoVP7C+5nq39sKkdxiojsqolkr20pKvk94+oqml8hy5sjiSh
6aV80qmtl2enDRiwtvcDNIkVRpEhaL2GT647drAXds0zFVnHpF05I1QWpHB5qAO1
2kaSD2t2UgqNxzqqdF9qN1iti346lzOgOM4fcLZmmG0i7f4hjOny5ikQkDPNJa8+
hE1IbOcyiZLlBsXMoXvsi4U1cU6Nav51sO74wnUACL4ilTptOb5qIPy0GYPLY4D3
YKV3aYkW7rcIlrg+PsH/sa/2Skrx/14cJWwf81d/ya2QTPO7Qor3o7yPp/kMtlFf
EGZQ0r8KT5H/RDfdb4gu7MO+mEphDcLy/JmGz3foNMVyBC+BZeqrL7HoRRT/gGlv
prWDwTFrJuoKmasPMVgk5ssv15lq4fNhfB7OXxHCU4MrWa7gw9Cj/oNUjMq4hDIf
Iq7K1iQm3t8hWHsiQtc3Coi4A44tcw8kI2uFWvLSx5S0rrm69MZpV0ZqsnyPJNLo
852n1wvJeRPQO2GQoSYbrTcy/Fo3iTo8cbaYvlyZlN2iqZAxXJzMNDbKs0J3RCiC
vR9tVK5ru1XlNJKFh9v2YzL916lfb/96ATdhb4ZzR62AuDD80VmSAATf+76v87lb
1Rd2h4C1f/URvFEVkySVsNaPcMg1xkTsrNTVL/ngysr1EsegZkhFI0HV9JBcxT7Y
3wIN5fTSVPFa7by8X+shRZxCMONcl2ldpFgZrepPMJMk8wcIuCHJc9ustaNMCYQj
wsp+fiMm1pfPQwcrRnzefZuTX2hbSAD1skpjLE/s0lYr5lpNO5deKZuOWP6YWP6I
LVGwLVkY6/zNR7ePkGqDEs+SUXXmnFDNfDfvI3rwUnJSuH5lv5JdGi/c2thl8yef
6RwxshtQ4T9m7X8vKtlCIZlGdGlxXgySceIoS7jCwMu1yx2ak6tv34KY2N0AyaPL
Lb9GcXDYtAkOQk3D5zBHVkKRtGfwxwipde7jWt57MCfJSTeSIVaFCh+lZceinYD4
dq082cowpEVFC1lXKpAOeAdRt8ZrFYqb+cYAR1PIgBd5WZW6NToVqIGo0UHTBDuH
fUHhEUo2tYbQROKwZ9U1Qda1lxogz9HYslNZ9MW481H1FABDG/Bf00PlHlbwtMAd
wj0sAaWRL+HDXDMgddN+YDVULBlYevHL0PmPrkj+oQj2V6A3wWGEJnL7VzfHaCu/
TxfYreWsCRI/z1HsDKIOlyfC0UGoot9D3Ga/SSMDV8sXJH5N6QElTF4SRlXmeLAL
uWEXUTdi14To5qHiwOouXUH8Lh5ovtLFHFOKFFsIPLU/dI9/IOWBenLhKcIhjpxr
K1ViusjDx0D3fSWvy9Fxy2KiFR/i/kgWxKPzM+yd14SRbeT4SkkKVet7ddNugDtE
RwU81sYhUGC6iwwGRjEzdRpdT/JI5aOTi8eBT7oFNz2UtXoiZxAb4qRMEerbCyoE
7aH8x362YpOw3K4oCTtKfNpRQ4QOuH/4Ewdphrnsl9hejWBB86Yzsi+2pZM1t/S7
mhvJKx2u0d2y6k4xXpbeCN1M6Xq4MYeq2W1zLoZuq8Ekk4cDYYCvx/8hgqe4CMbS
c1LkWMSIaruO+4GJMd+pTc5uLbIlHayQJha/pZQURammyRa/8FXRVi3nVOw237h9
GUHg1gTqSL4LAWn46HR9UfD+8E4GMBGu6QaSo/sxdzODyYykYmqJVNldrUvzVlCa
UZYnyKa3A0YKur96pZqQx/XmGa48l9yR3iE31RF2huYXhkhyW4WHOg6yyFzHnAV/
rjagzSLEzuyRCbj1CtfeN0LsuHG5i0xhFydSVLm1sapGd2gn7XcW8ElLqr3H2XvB
THbDU2KGlQ0+Vc7n+EOAsBW3e1qPfa4sMrTR2RqCbzio1hDfcdZJuY+SNUNXcZ+Q
MGQpLAb99pfvZqjN1w5l4GXIZ5Th3+N/oKiU/jgIkVDHTn+qixGryPE5b8Kwb0kg
+npC6Mk9VL38LYLsjCSAhhdmjYRj5rsUGKhDVSay+2ok6E9Ez0qG7rQrbBDgv4Cy
0fCY2OM9c2L+gqc0NPdid2oX4WfberszxV4/qj9HW46nMXyoIi29RhcAZcSmSOMn
5XX3VDdtyh8uDKwjIB4V81wJu03RGKmJJiOr7Nf5v7MmqXMSjbFk+gaP6pENacq0
eCyX7YN4hFME6hXOkl549iRwC0icSoKZFrZ1AwSkpOFXNLiggRtMsS+ueNhAXlUn
erGp5Uz1ntt1weo6twlpbX98QzOl2/GVgwhuHTbN9vqjogGH1vcM5jfL7HAT7d06
2tgZPsd/MfUmdyrVmQraoxvWBLrRi69rTI5+Dt5SJWbkyCRoKq5w2HydrjDTr+rN
DiiN22aCdWxuaN8mc2Vap5J2k3iFMz6v2g2+014OyJl6h0GkoelJTEF+gj8OwccX
M/caLgzryRpdsfNQx979T9F1vYjDStKCuJ3Q34EsTvNThQQQkvSkiruhtsmMfV/9
fRqsg9PhxJol6VHWbm/8ecOCan51P0KEKCb0/iGqw3e5nva7SVU3l1oVzqaDRr6T
PdOpA2vlt7qr3S2YVTd44Gp54dJtc2rVp69gXyXbdXen0vgVts3HdmcGmMurbHPW
WsRDNWbIdhSxU6rhXzq/GdxKOQFrjcy0Nr9KWQ/IBG7fG6VVc7R/Qf5zSuxrz+79
nCR6jn3EBhJsdd4hzycOXrVy4RRqd0yWzd1cELaC6hwkPuu5S4q8rixbJlC/TlWI
qprw1/1gaI6AU9isyRWmcBh0sBx4hE5/iXh6GWjilbzRNn/pYIdpRv+9a405kL2T
P16ascxrR4fWluZ5R2Q6afe3OrrD3y4rrHUdhl/KnvKfVfqNwaGYjYSd4Yr/JWUs
DmNJYlPLh2r9Qi9+lW4XDhKQuXXcaBXHss6rFGQV9+xWDV92Ws75frXwCcHjZPIU
93EY9799Qg+eCWV4Or1Yrc7BzE7zqxb91Kln4tb5fOdKmXL81bY7nosEjhQF+/tv
+2URyGNvo8W8KtxpR55R4x0EVdmQBuVVjrLDR69Pk6L21A1EHFUUjqo72FTz6F5J
ciQViVRx+S7IMbPFTngDz6mwrIzJkQAk2lxYeC3K0QIB0J8KPCx0aq9NVeNO22+Q
cvHwytd2AU1MV9f0BuVbMik0TB3X0wBaMVo1JANW8idvBP6mc0Oe81IJB2Z7UUeE
JnWg9xp/o+TfBETChsXGFwpjZvnQSpj1GtCysW62wUJGr5qw43g6o0tIHNyOzMas
X1ctcBXwlT0NA32FlLeh0zPkFwrs+yZCQD2sd4DPT/Ib0xe+b3NqDqrYWDws4kT+
D90+rA43hN2Wekj7EGwqwiuJI87ctpzPGZAcyWt5MgaUU5nqrN46xTGSj1qGb23O
ifYoT3o3w8ZEH9ZTZyzw9tgiokV6fvcbUJ8OD308ggzdepMZT3+MGZeix+R/oo4F
hgslMIoCclbgeBds9bmVltHIVTd2HSlvYiXuTo8H7UjTeZtmpRPtP+rjQIQyALJk
eQdHPHTkRFsf+mOxSIeq1rPypdh1UZdG+ft8l4Y096bjeHSxtWydz+H3IwZUsBAH
sVxe24LhM7xR9R5BfmoGdiAvuuJDbOYKFRJ0mGTRrpZAGApSKTp2qilXNiwonS+E
1iRbnIvWDZ+geRN3VOGP8NO0JCzlIynoJti7AGBKRzw1njL9kplwiNHZUoymKyPc
tmsWV84eA1JEZBkMim0dWvLx4MyWBAi6J52TrOoX7Lze0vBpf+H+O4ZOHWjS8WVI
zszFnzPjPJbjuGLZ6EkmklM2VO+/YeqvlcxHqKRZntknERTk9VfdeX2WlntlYbE6
SL2QIiRoccBqXfun/pr2Q/46atqNLNn1kQGpU334eP24fpOJwVb37izPh/N0kVbQ
YzTP1KALtpPqS6hJOW2SzuAX5bCep+0VkusJKLk7bhNgOq8arPlmMbu5miO0tvRP
2HZLdbGiJK3ttN8EmL3O8Dnl2nFiRFszkFotNbQHFejmKiFiOJGggkG0eqI80nCb
kb8AjtTne5H96s7v85Y6mKmpJ9VWDenl8Xk9K4AtoCY0uA/bxMlGXifP6wddi5oF
zcFX+siNtOTQFoSEqu3/UYsW9/kep01D4m6Aqya1HL2ZVUYirPRD1Cj1BARrAbCC
5kLXT1DyVeDQ/STeBnt8o19z/XZ3FoI/gl6UNui+zN6A1B6CsVcdXBS+sMy8fcHC
n7q326tkNjiPydl/04/Q+Sf3jkqFUiAA2RTCFNizHSBKEzKGHRg1g2s5jO4Gh7u7
OBTelAJH4XAJ8XSPD2akI/LWA0yRmOK4K4pFw35uqbpZ/pw61c8BPLRD9DrelmgL
3DvAtvimglCkf8Z5WMZYT9pAQ6jd4zZVZoZFYKrjGgTO020N7A28D8ftCgwxyoBf
IHMNA3DLf9AUXYYZiq9fevhR7THf0A8kXo1dXh/+VGxOIRPzFil27jQMrqXZvcI0
49cskndW5BK26hdOIJ+wW3Y4Y5+qP+pdRBdU5jego+lqFQN4UOsLHcwCs5I3zxL+
kapvRwGqcyZznFem2od54KS4VsUn6TqtkEEgBe+R4wz7rH3KLEVvTAHpDjHHcFEt
F6AzFbRFeFWoOJR0x3KF8JFUNLF6nOdmQrmLfk9x7C+1sniTqctd4HP4hZMhH7AM
1O0vhc/k64YdYtPUWDVPwUpJSq5cDRCsbnZeMMWkyLA29si9oB5St2GFwiAiYZIz
zkcQSLqhiR5OvIoN2iG8f8uFakmr7AVdQfEq3mHle/7gIozC4XyU+kOxdzkMeuhW
kNEUGwqd4YsZWWqncczNR0dcz+qfT24iXTMChcIL82Ix4fGZxrFYJC+9TCRO+EE6
28teRk63DCV8LUrHwXN1c/7oCLdOMz4TO54U9cMvxDaS7VHeGE9yd1pvU8iuctrx
BqPD/0yMb15LQSoHH8sZd7wCVX04DiaqgfIZ6JYrisSBKAkOd6uAnyYcOlTA2Mdn
BDJXQLN9FP9/SnH0HXSpu5Po01D5egDgIPU8MGiA926azbduS9rdYOAYD5QI/bFn
4FvGrHmNpVNxifAQ72X6Zy3jzt1R0s7X5uxjmJs60+AAosma6+WO0DQMNfV93dT4
GuunuJoQrvDz/Tq51Fd9F10+ZU3UjvwZaUdxgyoNU0A5lgseE0gpNL96mjs6MvoL
CrvG81TH/RsyO93qNGq7xUF9ZJMYK4GJpdcXQPh9vw8dD6IwE8lFAB/O+hn+ftnc
ppa/GDqvxCejCKV6wZikQzk8xr4KrpCYp8j78vh0zb0hY531jMA3pI2OyRs3n5iU
n9ChJcuqXHz/Nix1494zQvvvCHbLGf2NOLcZ7IB2iGJ3nlfmUCRCi0mWrJ1gP1GY
hCln6Qoj/QAM9AnZYsiIryr9ytLYbDnmUNZUx/p4NcHUCTC0OX+94zYIX+xKVdLK
zrtExkLJzOachNGfXSLFLM1hhZTa8D7bRPRq4FCJRv1VaVWhzNhfqvlqQW6jtkTb
20JE7PeRBKHpsLZdMTlGvcRHsNTLmmewukdBkaYauuzWjfIx3BKeb3RfxT73Wt7Q
bxg55VVUJuMczYp5VPiaYzKMXwRLfDLvDUNn7Omza8RS+0PSpk4Ob0G3btNpJzxe
WlrZBk5qNFtaLg6aviIEsUfvrprI3CZcJJ2RFV5jlJsLJYiwqql+ZYUagsdis51S
KNIXR6cG7QJ5t5PaL2lPPmSGM48r97RwttWtmpv2Bw40w1AWtvZtmGBRUaEyRGTR
CUSo2lIXE3MI7x9tbzBsrInPOCQ3O1LlS7us5IhOJ0p4i2uCvEZGCQkokuclfj3t
JhVLSpEG9IX1xjswga/mEXEndPU2IgEC8o9vNWeVbLjVDwhXJA9KehQ0gUeaDwyk
6Aj3hT1iepeUedJA5MTEcrqaii78ljrbEUX3mfum5UI6+MwtwDUwCBPL3D1Kg5Y6
t2snHMiZMmfnXCsLrHUv4+KhIQKlpJRqGEt+mGiSRvmpWwUpRuqD6oWrsutqsJ4J
CwVzCJm+zX69iAvaEfg/kCUzbgts0BDrgsLaJv2cyQeVrcy5Gyy7Du9EN4YxvdOZ
05JQZ1gF46Kr0GV5B62ebYMkpoBFBXpn5J8fXUO4p3CasYQM51zpldDxiFh+9QqF
dtlnmIXuFa54xzpJqcrXiG6ZcFuQKuxbyYAjgvzhNmRo4KMaeDeqR8ySAik4D98S
bB6jb6MfAKwc9dP22TI9ivCLB0jDlhEV21NtWjuUEIZcE9Mpu+dWoGJEBu6BuGwz
s9UKwvD1gOWbAgsj1vWPnfNqTBvUW987Eeqy3RgYcdJ0oziJtNJ+hIVD00Mo8+cv
2pmJqCow08MZmsbbTzlCfaXMjlV9irUbXrvFVZcsEC47Z2n9ALz5jOhMHbTkaPvI
eoLMbkVmxcEu5qZ1gxaPtY1DS5fteASNcqZ1w8WUnNzlkTlk8bt/stRlyo2xXK2s
Lk/uz2Xg7YFyS6dk9wGiQY9ahA+KR0HfZaEbrOn8UIDzjsbK9U6922DHJTaCEv0o
+AVPSfkXXVIWZV7dwpJan9VDtTazJXp39tosMNRf2s2lYesS1MhQ0ahgnxfO6jIO
2fHBbfFh5L3rNG8laYjByX0y5djQZXTp86motxRW2Zb+OSUjZwscUYUgPH587HiO
IfZLUZs98+OgAu2VEgOK2cdxX9aOLQF1POGsd6XBfNRcFq6iIcQsxNSZxbkDT0TU
h/5POU+7YaGTvH7Lkr7WQi5abXz5VIxUeUnLuGn6pkCsmow+G6oAvWvzPTlJfL+k
SYMyuBP6wh02uGpAhmkRKUoMd7MVGWTw46KMRf14BXAHlxfAtE7hB/7jNwN4lLKS
MzI+NWgeKcuSes7KK82I9sFRTnAoZHjKWAqlpKx9sSuUO4nW1Ojndg57J5Wy1Ztt
WRqKkzwdprgLpMlThW2ftgoQEj4kwpy/kLFri3SyQOdd+4WZ/nfeZxrng2Xb+I9V
3G6qnGzWltEyG1hrS6d6Tuy8Nz3z/kU0BVDclzomNe07FBICQH/i97i16HLwSKwA
1lbCd1Rs7F4cvhJoBDKsI4M717sXPUZXc8OeJdbnFoEi7mwF7dLQRhjGrAZpNVXZ
bpAprdAEM6dGrwiuiwQVt5iRNED6f0lk/nCqzu5dvsoGxM7G/xyYf8U9TbqUuoMt
30WxuxyZ/q3W6nsJDTe6uQS3mQN7/x/1OsQ3XpcYpYRpHLCJ1U07FnfYbUfo368J
4OBUMJwE7Xgk0CClCV7Z4bvkblwCrell1Wi4m1h4nCw+i8HQW7AbwK1CrS15ehU+
a9MTdQcEZR5zC7iNE0L85R3uNqcs6U4VoGCjjqoeAXDPgC6vDDN+RriooKXpfbzq
D+YFtkkUlzRLmjM+Xv/bmEkF3K2eVZUtsrFt0wJnXrXoH2n11Nq7M0XEv9vKwt/2
mM03goD4ICNeU0YBcCXkiHhSclQjY5lutq9DKRihjL0z74YTD/29daMjlICJSeFY
mB4+qmimb1b/y0mcbA4u2eINQG6Psk4saljvPDOErZV4WBrBhNYFCaTQNla56yHq
Rs052Bd3K6jo2QbFvLovUSPlqJXK6+p/TFsQ7XQGImNB00dNAzurU8kMsQ3IlKp3
rwupgjHDTTq1zWJl+mO2e/fSpPbFdVLVUVjFfui4zVvRI9gZgPLLTJBFhWQjcL7e
+XEOSgMWVlg0HfWoMKA/Jxx6hRjxdcNp6nQmZC9zQKGjYdqaXnEp4cZMEje5RQlX
qWvtpkfFVAKdPynrzfTcZbp7SR+bPk7Oqxm2vLPnkPbjBwleY2beRTNzD93eUEIL
Ba/CjcZzwXwsq+evfCsgNZPrbGe414Svb7hiUZwSDbIypZAeadJn/LLrqXapUh9I
ex8wVLy3wyAR1fn/s1t/ChP5+N0/qQl0EQlg5UVeJLjaqjM9QHBV5MSW2cs0rOqz
GzJmWuBXreHU0ybuV4OM5H7Nxz7CLSirA/XSIE2tcB8lc/GSrD1d3LZBN1LPeblZ
2eCaTt7qwekdmcdSet/WF7N0BswPRONVXpS3+py+X/RG+s4F2q7Vuv81a59rlqIG
HsR4jk3DuDngB9U7alFWOWc80BQ835HzL9TqFWxyJS+/GDsEJ+3OWybRkUL+wCtn
xouLf3/QtFyYbRnIFp61jN9lCHoTDNuDPseBY5onSBS7DNgE7LuN1z+4XhhcdA6n
zoHGNvhj4lrjxSFqmMghmBkQb0V3iFIKpUeJJh/4IRdJJxdYj52Pvz6Ra9MsKCUE
0jGlSaqWUvkz/+nTO2xcOFShcySF3s1ip2da30Vr12S4dl7vB6I5b054dwXIEaGW
OoydlM5zyLo5Ydr7x+SkypS4Zdp0RNZXvz5dDpON6ZkzlAhSKtYqAbrnGb81jWG3
UD1NcZ3HhAU6Zjb8wqgrNHxYp9TFjQAPBvYdeNTKlbBuyE3He5i+L3hKuCMyC2ML
UohpqE8ZS9ekML7pzOhdyV9DSPLiA52F5TZFMuGeIr2hckJ5HGnnPoElAvZmpo7x
V34puIIB4RBW6n1KaNnY8ptiu8bsfr2FBIs+Ln2VAdoZfmiz8UQGDSQflkcqkiMx
TG4PkxTO9Nd3PFQoKKN5jDkBGV00VVpLmsMnv/yDR4ejuAQhE7A4sdCIESWLFAS/
1aKLAFPDfL66CedGOp94AbHcQgpQQoKyZd54o0h4ou9qKCz4GW7JR8Ix55LGzWtF
uw1xFs7RhmTlRX3y0p99UaSD9wQM/kIkcn4W4mViQ/W9pxczKogTQcN8vZ3OeG07
caZbqEDOyfvWinirIn6yLQgRNv/W7xF15Zv/sdS9N7NqrQuHXGrGWw76NyHTVa5/
/XaZ68LWB7PmqV+22Ds/mcaZne4AUFji4BX4FKciiLMGUf1l7lrkJ8p2MccWMJsC
7r7rYq/RGJLUG+lNWRbhhv2nKxuQ45OfhArTPRxq6CT2esWsCtcwKExq8/kfLpw/
89Z8OJfXBI/2Hb/1Prp7uC48kzw4jU1K3DkvLpWJziwm0LlKUxX5cJDZiq7Nl8+Z
lcLti6xJSV58+yoJqV/iuW21DXWsoitXllvhdjG8qI4WoQj2Xebu854ZFjSN5NKR
UJosIXuNMBFPE4mF5d66X0eZoxm+syF261cuLBqgEMlS4OdDLs9hYoql10h50r7/
rd0Fc1hMXKrimNSoTlMu79DNp2SyHIa84PfZe+7jQLoTpmo/4dSV3IdkCR9Ft89L
YL/q64Z34RzZd37Q392AxOUkQJCqhoNdnUxCEDTAMyhgM9FpjdX3WmKbsZOzAoCT
aJ/RTr8iCumt9PYIwOlgH7WkWi65rpUajreNMwwyxsw3b9dBfsawqMv0CwPttiPy
uvxpSCJTAI8PFzKZEqgnydyQvVc/FYR74c/wyuSfTuLvjWD0NREb3Z7I8kxdpUaL
xGPC1wF29rRimxRsFwJdGMVkkn+BChtHPVoXPdvLTYkB6GN6WZPCEq5rBJBrezB6
UUjnwym44hyac5QlFD6aXao6b7WBzAFRDVu8Mf5flC6mfLhhApCwy9CnX0aMa2yK
GlJ8pC0AoqKaKjz+HCEbAFIkSwpP/VXnEP/uAZbJHQbQNN3AOmlkw3Rz2wp205Fi
51qgL9mn9BJnyUlaHY0EURooZke19KLut5sws7ly7+E+nHzlfeMT/G5dmBmCjlmZ
Dk4ntF5u/6KUHch5yVAyhSAdMrNdnJxwQvqe9Y3TOtQR+vLamYHgaoB9uM2rDBsS
Mjn7IB4V14aREUkY452IE3rLvAeXb+ZZOdBKxN6rT0Lab3auJL1oYkCWPWc/dxU7
QH/IDCqFrj12CWkDhvbMdSphAxtSaE7xuzQtYCSvBnR7ev+7vFaPckUVq4sReI6E
4GdfRDoz8QN3tisxEMoNqJqfKK6ZjzoDx/C7MaAaCCO0ZawPTS1adfUN4OVKVeCL
YoMBYSGVtq/KkR3XoE0ZQvi+uv1TGP++JbR567wYlCrdZBS0dRBnDLpNy50ODqVH
Y2vod+oG9QnMkp1oEKVVgyDqU+0mvVvjx8Cr4VHSizBpZpV/Kdjp7PRMk6DY1NvO
WpcjjLES/GQjYjHKSMufgnjzd9q1Ei5AY1MjgG7eSEQMAE+Z08yHXGJaoXbDT3pV
EI34fQbiOpNCCSWvJ8bBZkhB6gaPl6iha1GWMK55tgEMKlxB7PVL3QHA+mU5/vMR
yKy0QT5o28pKyZQx0XAsJqOelTL3IbMWrQ6axedNOjgb9CENwPeafuVf4JsFH1Ds
8VYJDStBszKTrHigu924/YiP0Pl6JSkpLOXNEwavwFc2bAtP1sIphLiVlweHHFgr
B/t0lLOca3ffFgcIwoTk/7Gn4IkUXO8rzi22CKkglPy76vMPSmoE4vybl1xD5AvS
TL3972vSyMon76muygOZ+GDiEE03//b7Q4kf+V+IsMATzMLR/3duwCnaszAuVTXt
STJRWr9NlXOvKt9gidg6Jytomu8KCUQtfLO0Md00kZIZjMOxGJuBfTI9VHRd2uI2
xmHgFKFYrqLw2250MLFJ3BAOvs39HDoZy5u7Tv1CFeSF7MCUD+q+eodvqrES7vVZ
itrjFIMt37BT/IVV1uspsSlUUm1HLSS+Z0apGvdrOZ2XQ6990jgll4IPq/TR3pCJ
PGSQ4+Q5/0Q1n2KJGfNdPaTZCGKlw8v2joOgWsvsNGZTsg3VEDPios4/3jm5BO7T
jR4dImz60ZeJpPWG8wZXvJBJpN2gKlJOi+WLpOdJ1CUmmaNiwGho06ahLOKkY5JN
OF776dFjv2QsYH9VXOuPNm5X3GkIAl6LgmiUuLquNgLTHKpUw0TDl5HbG9+Pv206
dGJ5lGS9Q2faxD4jNq5Fy2fQRKbeAhfSSdE39dOzhAzoze7WFr0Rew16IL8/kOgA
9MvrjwkwDWUdGa84+wwvx/LSoXMpvyoQISQDgyi9asrrIpv9dTXvFk/E458OQ1ZO
br7ib9+KF9OcuppNwkfoIIW36Gvkv7JKsvcZQCcbZx2cZ2sQH91TnPBzStCbSbaf
mYGtpzDacBzzlrDCjHbBkJkRLlM0od0OjfwsBTzxBpXMN9xsxFFg3VYFUCPML8yI
V8T1rWCBZLmfC6PW67CemrjpsWJ9/CvMNFHtBQZlcvvJXzwRIG/1vrTbGjiYMQrQ
0+5tO8hTsD1klZB2tQne2lg/tBM4TXgHMDaWSwwycfG0kwDUhgeJXUdFA64mrIp0
e6BMgvXnnaeyy1foA/eXIHn1GqSBSojbVKvhQBJrg7xY+LTiLteSDegUI5331EGE
c6dRd6OhkGVnrg4kzQ6TYOkTOGZ/q0rflmtHNqFG+3bmPKybK7A5aSrVQJcEj1iS
3i+gVzxrhceN7jb+M43+MEq3LaElQ6f0ZIh6109biGBLdTJds3veQ6QBEjtC2FA2
/neS8wYjGCQORP4hI8a9npPOt+rPE7mPUjh/luM21kj3om4uRBN7FnzsBJWqANf/
afV6Lw8LgAM2S8pIK7aBzicXUHVaF1hFIuw7wIG1KLbs2FYq6R8ATNK2/aIcHBJM
1Oo93WuyIT/Cc+NyGu8n+KQNTo+vr9H5LxEvFKq92VHaxyZEBR0O4747LINBvvUN
uvc6sn4Fjfzc7INfSMnsyWP9EBFGRJ9nrN1b90rlyQzT9RLO7FpgL2p+gCicxnB9
/Tbk1Sp0ytYu+DPeJ2XwC+ublbcuv/wJzZykf/gHoo4+pHK240BOr1eK5i0Dvo6y
EpVvRV0oYjlsEXnJdqdQXX4AVVGH8kYLWB684yurRziNAteU7SCuC5eK1yccRrXY
pVoOgP1HuhXlpWyzuKHuAqpZ1iNzHRFBCFp7YyVojHpfWWV8c+ps8854SElWLnwg
bKfTsD2JRevxrywHMCgXyC8SV2XncOw19FrCn8iqq/Goh1GiNmVshdOJDpyIEo0+
dUBKwb7L8MBcWBp39hlMA/t/79B64Tx4okb7e7gf8AhOnqPAq1g+J21FiqTLh6yQ
s5rbj6Ylj627SQ4xso4bF2QNv2HwGQTBenQuFZnKUT8=
`protect END_PROTECTED
