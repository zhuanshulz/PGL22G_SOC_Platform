`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SzOiu+es3gjT9iBIvZXdJOukhgymCTMJA61nJVF0XNFKM5Kgzh7UOcF0PlUv2Syh
Mnbgoat32MJLBARyr3N6Q0k31kG55KXR6mRXx+oi8BKoL96dmYGFdAVRySdKpgJ9
Vdh6huUAzuFJ5KKIMwDCtfh91BaU2qBN7yFH2q7Gz+d8/DcManaB9l/z+s1hU1JG
r4GVP/Q2NV/rWSWYEUC3ot3XOqN9Bvr0/GuM32/nJy87m2S1opnskUubuNJ8Q0Se
Hh4LSjSYWS5e1crTO72U+g==
`protect END_PROTECTED
