`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFBVyqkW65os9pQHTfg3xLEWqSP9HJ0rDx0cz7zEe/AhINzeeXty2WIcVr3KNcgv
k6MsqS7QJbruSlMW5gO4qQ6wi/ql7a2L5xMn6/qETXrHUh9zEfPfOo23RhGA9RJx
bIxV/wojT5TjxDWhysJY1ENl9PyzHpLdQdkN7gLWJbcQ6aCFITG2TYr9Dt8M56de
HaziQ7d5nRwSJlY/OzvppWlrum58NB8t0UGSc6sGtUbhXoSp5n+y2bSZUkOe7Pyc
M/V5Qw+cjlAQIWGwEpviDgkrYVLAisM8Heq8mzYCBSlYVTia3INsblOr1SUfyf0f
aCu4swoUIS7xt7WW+KHpuDPnQOjzGAhBQCrdiJ6W6fFJ10cvsL3mXy7jhS/prYy6
mPqB2L7ZE4xwVf36U//wt+Eb+iqbqVwtbpbX2iVqrZ4DLIVhZJSOrCGbyKjL/DW6
XhkPgo5zb0HiIia6n2xwP+dlTBmFA/NENyvCCaE/sRVYGkE06WupB+de8wb1iv/k
LwMJW5QjM/X19nZ/v/hqvcqUKnXNrb3iSJQIENrUtiGswOyL0yh/RbyHXFDLvwqm
jHIX1lz3dJucw/UyaEc63W9tn2BK8sRK/oaC0fUDEj3qrV0qK2dZ4WxgHkVMfYz5
c/RsBIli3KZVcqDouFiifEcpsHpOLVMBPC3bk85LV3Yogu9QodbvLflAxQzbo2/2
1XowVLJWEva1nPbZaCR1MXHIOK5xhSP+6nrpcRNFKzT/HzVSFyS1fOdbY5hssc7r
9f20XiaKuJAMlar2K42l00fa/cXhWz1xdtQfgtt8F8/9I+Mb+//U/I/vQdh6eI1I
q4jW3QfhrCJN+ppzW4SC+c4SPBvWRnEHM2hhgwSutw9QTM2LQdCxAy07R+C6q24m
ds1mF4GCCWFX9Tr2kAoQrDnEiDgDQl33tYI6Qceu1S8wsHSFb+9zvH1oYlQ2Blap
JIphP4+04tCTcb/VcquRfMGwK5REVXdrJRTzKvDSFZ6PvWCgzi3HKnDxxLeeLb1/
SI3oMSkVyNbmHD+TTcdHjL/IaxtTROzlF/D93Pb/Ite2pVulthoPU+M1O2zNfW6S
7JIP+urk5kvubcBDHCXOXZ/7fBJviezj4upydyR5vNRntUs1/LpbWUFps5mDtmZL
iCvHz+Go7r2uJYkUBn/rdacfPOgZzFf16WMH9grCd7ht3p/zXvtG0SCKSYS2KpdM
NJPfHKSiyIurN4NvVlnbXN4oTqbAMK6QG5c+VpLqQcjlrL/Dwo83c+bsAoRhGuZr
pjB/H+Io8w/qyavmiBteShycHpXcgTI3RJ8LEBvPc9pPS6C6BcGyBHkfNSpR9jbc
C62EyvgPM7/IlbQnHmgpOH+EAP2dsftaFPRJx2Yj1frhT5j5CmsjaORax3xGk8Y1
pQvBxOmwQORP8JILq8Te4kEOcy30dIixTBBOfVpBjSeN9qptLZp2mdMvtqGR/hst
TT1VrTJTyGP2ohzG+yd4yQ1IoXzU5xgNMA4U+F/X/nWzpA8ZQoFc9tlOMp+TXZrn
d3gmvVdXusN7u+0/PdVdQefbY5oh0xsLBVBDswjPhtINkSSZTXmFuMSJiG9Q7xhr
x8Pd2rS4oOSJmS81U7PzqkrHAeHHeXmMbxclrgM6WYVRG8d2bOZQ178XXAMxDw1p
DYdOOituCaOPYvrBH9ytvyo6kMvNhLxOuW75AkCgMr3FXUTdkEDnoqy6U1MGvnpP
TWMfzjDNfRKvHZ7GBCr+whUaH43O4MZjdwzbMNdBYiF39zBTrvdP2P4kRaGuNQEt
bcTE8Na0DPPW8hzeAM5I56vjvR+vqp9JZ/gMfesG49URmOF3JRSYg4nhx4KTbLl+
+uY0oz52Jc2qXN5QoTkotm5mYc7+mvApo1Kz+qGRe0UHSZJOcmDV/oYBjM8kGB79
v3f0cPn3DMoIxgLtU5re296yNa1Qm0V/dPreDQoTrUalqeKJGURjaqFs7cLwsQG2
omA2n3p+262VwRIs18AIL0bYMLHpF8Z3h2eCAlnDVCVqfYvASIarcfzWJR7XYn3O
tx5Fb3kwWjXtsP3/Ppufb7taxELOdGI3spgJoBJvIiT5W1CPLigwz7ZbKpHgv2Eh
MdrCrmtebGKEKiNsOxMYXaa4DwM5Vl60zdcpARHwSufOa0wdaqikTs4gO1xC3e2I
+4ttUdI+7MVS8RGiZSOkNrab6JqWHxUMR9/Mi7X8v8UyBenRBI4OFyoeDBiwl0Qm
d0QQn8yzsuz7QJKXXbwnFsv6QwgJJ1PhVIenZ7eWgQOP6wMu55aASYK24l2XNhB6
mq+Q6VfHKEVAZmsNAcBmQKhZLl7l9th9YCcjkJWqGOl71yPbAyWRLyq805ZB7z19
g94InjR1GiuzS6obFIIPqOguA8HXDlYDrjhYV4CywYzzlECGYvA4hCMCDAk0YKZJ
17qiRyAKqZXOn5XYc/hoJ2faZkblFbTADVyxGUImfU9eJrpsj04+XxKbDsetcHYs
TUrEP3cq2uVB0Rxf6DGxXzxablsydPwxfCY8ye31zIPslueNsiBj8QMLiFHYF8TR
UUL6hZlbsQXHlt7RClOqB/yqhILX1dpS2VITwMR1OfFAJ3e+g+E5e+ywGeLlSL47
KD606ix6DPyIOWY3BUbZTV45oAqlaVJLQsWEBY+JzJXCvlwPl7ntXvXnI6hE38Tv
gzTZN+WtCD18lDsp5vP6FAck14TZmNMVU2sVQHGvQraBrpwiN7Qay+C6vNIFhEAL
FUoo7GbrLfGxRQWM01ihFrRXFz5jtgnlX2Ild7dKQDf+ph8+r743OS87oNWrpMhq
GkPB6krpOfH80axZWjAIp144GGWjhw9XiB8Rx8XpUqi5HwIU+O4JEonNJsOzOgz7
g1vd0moBVPxnbSQ3Q45vxojQbJRZp9T1KwUntk4l311ogPmYYzWWdPFey8piPkE3
kqld20YjKkiVeJj6XWbTfuMA+BrqLkM1nQdhdq7YRx99SRIxtD2RSvAJhaUVAIMB
DYxIZZ6kwQRDbYLtnTxavuDSafRKgV88Sl0Wfw7jeA7ha4LJL5+ZFhEeGa8hiF1z
kKALk02g+SIC+HcnDfSwYMet1J+iTqgYezqpT4pOlkki0/6uQNyc/3ahMAIggiUi
lskv++vqFf30uszGeWsltz+ksISQXhxO1+SRxP8+YKE0mPOh0wvrLmY2nQSiOPh1
EV7yPnJWJ89Jp+2XAN+a525YncExCGHXHYiPgEroZxTeG9l7Y3iDl0umOf21Iasz
N7viT/jG7lwHFQjDwAKUfallTNDOTjeY1AXFcegG054W2fhTgLqFvlDz5eIuw88f
GyYdBAojVTwm0TyPxIynPuKd/RScwhsLCLKXvh37gWVYzeingywLtC0v9ijUvLyv
uiDl30BszFDyiasJdrPS5+bso0KnzVRzrk5rk2BXU2g=
`protect END_PROTECTED
