`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuVvcqqdYqEHZ9AWqHVtwiFPzb6E2FTiuwxBjtSiSe7tSW97Q2QcLz1T0cYUrqw+
F060/ZUGk6j1n81a3uqyWLDdqS7Ep+WDSbkgZauG/K3Yl9675kaGUcfLmfUvRnAC
xfIQqvxePLxlw8IObK+M38Tzr2utXjWPVaMCQ/D5yrrcFONT30Ue/IeGaKi+bECl
CkEWhW0fyYv2saGkyMiRJjEr7X3Pz5AKKV6Z6ooWYcGXMgZp5+wNaOWKxWvq2q3/
AyHwpzL347c+P0adNgVwXn2YVIFsmqlDnyf2uZRypKMeB1gznIBO4yuZbrbnzNeT
1OHCd16S+/HT1ex8swdIx+xKvJ/RuOHhahymrRY4QkGsZzGjo8qnkqlsDm9uSS66
MkV/wj0VDIzX95S6rPi4UTWpGby0Xupl2Y/dQJOfC/HTsw9k9it3IWlojdxP2S8U
epEGsKLqO3wOH9nulNAEjSkkkyf9pVITsH4aW0yj1NWp8yHb9au+Y3EZ0MTKWmMw
P263vn4EDBMHZ5Ktp5HYuc7dDT/wHqCKGEKZt/txpUjaDWQklzByFpH59XQ5cdoR
`protect END_PROTECTED
