`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/uzw0N31/lIAOGK7UQSER9wTJMg9SbPmx9HvxofcsEbNJvI58RZFOzA1Ae5JRH0
UX7iLcWI8C5T9BypWiU3c6HjBp/g1qh/c286kFDqzePTE0CdOrZf3ckS+owdwYIB
+5jMJmL1T99Cm5c9zfk0xft89AWOqlzKlC3ezq1PC+d3+BIK2oZIjG7p8Qp6UMnK
UhRnrXhdZER5uT9n0at+utSIwhDwacd+TREQcDSeaQIdHc/JnnIReEEgikcQsaHK
sHDvriJJlq+5ko9FGNGiYJmc12Ln8+FDmoSHPv+a2HswQ0TPy8A6XFDjuHix09p2
hbBXDmhGR4pwH3mJ02EW5obdS5x/QSHCNyWe7H0UN/luAIBJ689SlRC6RqqUtaB2
G5ck3uYuMXUpQV4ykXyYXFvtctaOQaaIde9V3HTw9W0SN/iM3JcpkGLuTfCSewIN
in1w4grgvUu1u6NJGNRFGqXTDBK9Yw1amam2RRtSVAp7FuCfuK1bW3C/D8SHcMRC
/cAn8L0TqBQEizDyhg7vIHkTlPvnyh4a99A5+GuOstRcoHA8sZNxmdwZV64jXhBP
3c1K5198ie7tJuF+1l7rqpDYH5Ny+5rllXY4bmQlMW69TWJF+y+IJzM65lCzJ+Oc
5fMJZ6BMDlJ3dhlw9Yr27I4jvgs4o6mAcTfaCgmkUB/SdFX5vLmTI9T6/KOuUHXA
1fFo3nL7tCpafDtnUpwxs/WqNcDLz2sp/65uYmCYayJAp+Rtdz7Ws/6rrlqyJfbK
8Cik0RUQhYRGl8//z7m4TvhzVOua937BhgJOhVIUSD3+rDRb+ADfpBsxeqoamewk
JabbM+xIdG9WrNt1eU+StC0d4YC5Ij6aCSPRFpQzQlxH3hpxQ/HxKttsVNsHPh6Q
0U7L2P+YuvU94u3Wm8BvOeIHa8NIwqPHbVGmH4rLsTV/T8m2g+vp/UBnZ1gSb0eY
QhpjmO8kB1TR72U+cx29Nv0g9zOaW4DC5R4nvd5XNt7CJt8xR7ueMxM1BYn3+nO8
/uT1tMCmdYQTCJT+L5BemzQBB8jIyqZPFGSLmrdSteFLdjYli5khHoD7Qk2k7kSU
OHTXOqevhIP0extTlpDXGorFvuhnutRx+OYrVi8gCaeC0HyOONGf8mBw0TP1eZxi
1p6jmzj+wRHAN9Z/PzH5CEV8tSxb/vUgtCJ0hNTpwYhuRqRA9KdGVjYp6FSYgCH+
0OxCeJS60adBZyBj23lH3BJVbqXMG2Qvl45P7O5rP8jKFTCKS4BQYc1XgKXIMdl7
T0r59TK26IdBcZB5ygkIUB2s1BjmTMh2VPJvc5X7Bjpu58zvLdHP5pefRv4EYCef
Kd/s8kH5DxZNLo+ARyQleoaxzNdAS9xUNWz/+RH9Bmg7Ak/K16poc0r5ICUZGU8h
aQ02yr4080QoSRPB58pArnIPUFK7SHhA2d3o0cvGLCH964vTTRAdUtzm/TrSVLC8
rGS8kbRrtJ95x+XoR8Jem9LEpQhR5QxYLoF3T2Xyz5Ojxf9HxblB4wKDOKNK+thz
egI8H9OqVvOgL8p5BALcmijcyM24Z/B2+B6ZnVX1wKyZV3NqaW9Szswpane+Q3zq
GI7f59CIkZ3WbQm7LYEQIwXPKmHv4qExZD2d3rhKAYDhtjSbakyyHS1VE+Ghcs2T
TGKxM+eqsGp4/HVlmjl7kE/sIS+mKtCRHT7LDOg64eP5nunPHI0TPH0LGoUt0mrt
tj3ShpTGzqMIZBTy2BxtCeGEARce1erEraPD6cRv6Vpr7hF+GjrkEd4hsb45QDPx
cGHz2nFo99xdUJsxAPuEVrQMwbA/D50t8uJWZFmykLWA+QvS5gtszIo8wXndMftk
SrAi3GE22Ve5XX/u8ADO2yS2t+Y6hzff+OGp5LgH1oQjGqLt8Oyr+bDI0nOw+o/s
IPV/F1Gp1h3cKe8WwJu3tTbVkmHmfDt5uxbKyRlhdq1dDMkUp4GIpd2X0hoV9JNs
xjzhlsRE4WSKd0pwTfJ3PHBFQj7M1Meq7OY4IcstVS1F5ONcbQJN6cZpgpX/y35i
TfuNqH5o/IrWEYWYAU5McbW442COxVESSZdDuxhZH9S4X8+dbyAuAtf9uvvOjXk3
xo8G3myr89rHGwpLh4OqPn80SnTIkJ7ZlEuEGaG4ExwR6zMw6l9IzQ+TaRSjtwek
FZKS6brSu59bEp79GBBMyKkQZDIbAAeAOYLD4CezX/x8/pY/YgjsDQ5Y9k0ehAep
SgSEk6TZ/upUXY3Ymm5vV9OcoJ2DSUE/KaAT8XiHHQB8nUrk/Jr88tJlyA0X9F1S
Mn7BRnbj8hQS51w51Xy87Y1RJrISLul2OQPcWeAfw3kHEexSoNvweF1SYfh0XXGp
g2Ui5JeM15YUHVMPh/Gpqgst0Tl0rSOyQDWYDxTgvN+StR/JzCuqvL0pgrpUFgL3
MGOVN7ZVaAwbU7yGeLl8r95lcmbesq48y/o6Omoh8IGjyLT2UGuBJ4zK3r3r9n9I
uTy52SGnfNdJmbpdPSme8xPQ401R1zRpzpEWvoAuAPbVKu8CiSP0MD73hX+m6KGt
01MZYGdlCQnolq47nEUzV7D5c3GS6wqdWuoUYYUtccsBMXx/wqM9hGHNIbjQDpBw
8dG/9+jpf33+qAbezdPdh1QqLjz9o+Oy5iiVikZFSh062lvmU7SpartmMeFqAkX4
THBxBPUheaoO/R+MV+nDTeOIqE4KiLsvluiPXJEMNdOBcbtNS4xoIFK5Okg5NP/K
oibxobelY/e2GLT44VtYfMgNPQh4VsLWidQtF1E38rqas8bQF0uMfjQHek0D6KJO
wZhwHdKYtgK4yFz79nkV8UmVLz4usecX0KfpOiUZwO1dOlUt9u7u3JZcMfW0k6Hz
5dqJHiavTqc0HxRmuhGJXjEtpWxz58ucCj+aC+B50tmCxvtb8d9mydv+tMDP84A1
WwfV0q4Ux8A2dwcQaenXs0z/lo2aF9TuavQify43cL3SKFCcw0SjqNkfVi0nNhw2
UEah+iFRutE1Noe0qB+PV4T5JTbbfFkvmlqm+xs/hCNKwaJzN25GTog6LiCwEoQI
2PvfGZ0iWDDVl7ztaggK13B3673+Z03LEkDnq9zgLm//q+wL39v9i9wAZa/i4p+c
/rjJG1eC3UEoqDKBm7hU4Oiz7N4W5UrNcLtzYD7OzAkWBwi1cRt+HvLiM/teOn4O
F8J3jC/wI4Xo2/jY/LoVS9wzfQulc66IMseP0n1yDJRHvXFR67YK1HY8Op+TVk6Y
Gtbt/kIBCEKR6ewQsPEEraaM8zbU1/RG/FhnyAaxhMjM1D0ktGJiRF7332MoSWoN
O+YXq8fCcqIXfyDNFhQKb/EsUta6yCOR0Fu6/0wpjutMdWzMKLb1KAccc1rZDi4P
8KMcOYJ1/FPmyto75qIJgNjdDug4GxfyDGH8ta96avAcSpW1ASWwcjTp+1/FNnPk
awxcwJBW1KBLdI7h2MfBLTvsL5HN9hd33V3l7Z9DW2YSzo3jUDJ+saqygtkgtuha
eCAIm0trkAkNMzjCeZkwe0p3/THcPXvIChwW6M586xN3MuHY0TsdOJsNenr2s7j7
Sm7tQ8s+H/0/S4sfH7hT8gb7GVYqNiBIA6QD9n+0DeSPyth1VKmlxleZ9+9Ebn7Q
rF+x2o/G0gggnq1DrbYdpibAPzSm3+IUz1yPLazf9DC2wpR+nYxNMdevUUdHDUcH
mP2Qn8J3l1oyTgwcvTBX+YXrQm8xNTRdV5aZIs03mpV/340dpOfiWOeYIHeZH+DM
YaOqgI+eoDWoxrlMzXtAozDqEa4+zyJLmUCc+dYGjvNRj4PlZks8Z3z4W4DOg8Uq
+FhhJdchShcZHu1QbWI4rHuEFKqQoGvuTEgPEpzu8ynvPTbxPlKLstfEq70kPcde
WD4T4zXNZ3937g9pLfTxiW/445kHAL0cf0MRO1se5Q1wKowWCqnuToGEcl3LTA/7
MyTJV6lYueGKBPYCNG25VgwHT1bN9esXwuhREh4ttrBZP1ghn5fD9jFc1r0OX4GD
G8W+81PQit5CXThgaCfK6ZoKDXM21MzHqzHGLbr2VF4Iil8yCTooU7aypNhK3tzw
odsPl088TWisno9R1kErG6bxsRwWK6KhKY/elfXAD58V29O0unsppQY19OPgwBSL
A5ffA3ELY5chyZDKk63cGZq1yj/hs5WcORfEn/x0wsEUUF6b4ZBYDKdpXW6hhkXG
A9iGn5EbLwrnZHldkJUetTgMgM9PlWY1unjma0tyR7fsbCSnLg0asx8SfrMrE9E+
/QAolZATBJ9LHiE3Jk3Qc76GA5Ycgu7JmNNQzlMEDw/8eLawFi8tUaNtZCamoRPN
qj4lE8Lt/M728vHi0/TB0+4fgUtBgQSYF2Ewt3Fn6/NUSa6nrpXsNCxPSBnrLqbe
e9pxnwZf9P+kqrV9mnS6gvGbMAZ9ze7kKMTAZTE5seK36DMbAzn4n9Z9z91OFZJE
zQA+rxdckahkQ6f9DP/niqkA0zjFpo3XfVR0os6Sp2XZdrENwp0FXeLAu6bk9Cwj
c4PJJumDNerzgZN86ybfAyk2iwiz4Ovh9tO/2H6f9IuFMeofXRlruoIwZvt7RCrL
aZvVasI+YjT+L1/1xAIziHsrEb1zf1r7E8T+eNAwIaQ2fdN9B8UVy8ETC6NozR/8
IU1EWJKzRJZDUM+hfG8udaWkppNnHsk7GoupYnffHVT9rGeoOilED5nWzhQtMLvg
8eg7xZyuppNki8xugo6MhA8xepeXI4ig5eGIoAHra0tzMwBnmSPd9D6YVpjVSrg7
+XWDWwEe/PvjVB6g3QvPec+IKGNvK85ENG0mJCCbetl4DQW4mRXrpQVz6uggyYBN
M24DdhzHll5zxHrqxlmTwMnNE7NUjZEGUPgnW0W4FYSHlcZVrGl+4ZyXo/BIaJ6V
y1XktrcBL5V5QPC9c8X4QI/xLfNXYuaMxQ1NmwQ8WzDWt3QDEEapVhqq6Z/TRGw3
h+ekjiLGVnUrz7B1o9NEsWfQQ35O2IC7a4TZiXVpG5O/KPFxwc36+gMdP6IVqSzE
vAA8sbeyoYo0whkz1ToxNIDBAF4jg2+ATacXcqLXXXl3crghVoejuofe/lf+EzH1
R/TrBVWrUC8ySRNz/TaVxVopRc5q93z8/r+61aLNN1dtV36u8vVhacZIdPV4CeIQ
rbaVL5HUf+hARY4qssbhI1UdkwWeXSlAcv6QzXbe8F2uKhOLxnOggM7SUD5/BOpW
5f6i4zYoi4Cc7cbf1I0Gndpv08xmXu75UPE2IGAnToIKgTMTEpAnft7Eu2mm12AE
CKKH9MpGBpNoUg7gpMDUrHxQsToDd7cMITYfREYtt/QtrVBhntCUZPZHzDiFUYcP
sIsWuEX3W6oyLfu+T1g1vuu4YX7RGBVykvpGPtjdS8md0dfWv2AD6OjydnQBPL8/
gyYolOreluQBXEwrHv4gItcPqsguAqAl50a5M5rZKpmgjVD1ECfcN7A7qzsVVjmK
HuSTH89VUHlfpOSqjlLFYULVtwnWIu8FMPbHjid6ikZA9hibWlDEGYuPxjHGaAeQ
we6Hb6hQy1mNGgo5aPMGyp7FeRWdT+WQ4NWxvoPn8OiMrJKUFUAVRcLzRpy8gohf
zhfFFZz3cLK9pPAejrD1nmuYTZVOyXuWTLwMtIoIyiSkjaT9rprVWGHSy9qE15FR
7Mvbts6y3tj5ouoZ3jNoCubWvprqWC7g+CuVK5s13DfA6bDMsQdEaXWneDo2j3YM
++RJzXuhEdkcqTwAqMF5Nv7PFrx56oAVR0evIolyLWoJeW29ZPnFQIasLJSEJKW+
eVUW4laKgChjP0TQPVOZA7sqRuAiF8M6na6fA1pM90nkVjHbPEAa2kDyUsB54dZM
0NuIqEQKt+DA9O2mXp4nM6iR24dhjGzKuKHj53lDtGOAlUBlvGlQ5znLjJG1f1L4
RGYMmKkdgVE/LWfeSW1IZYsxzAFT7BZk2ZeWVgJfvP7cLmSuPgZbKgwhbs1TfCiE
dze0K86G8iOUk7wDC8GwWyTXdXethFxxqlr87/FUehCEZMgAgBOmomQMVGD1MzDc
LByWPhGh9vDJG6TRHVD8Gzv6G0UFD1yLDn2NrJJI7h1u99pBz+mVqlYoYP+sNJJ/
pBScQaPaUTR2Nz0BwGen6pfkRAEOuB1vpaEbesuBdsIADOda1mTduKLJyxYBGZtj
wBzf03TskzqtV3QhHyVCYuns1XNSjx8pYAQC+W6fNGRu24z8fyF3IivbPJwri3wq
Alx5zVEWAAsQiC4dOWpvGbN+OBhtqV4qb4/oduq5CnHLpYt49mNnocjMUZQEOA80
6KyWvOxjMuaq4duKkygO0afSOQ6RU1IM5eFDE3AxNZRUfAgijSKDUWKqCU4DEpk/
snTZoPpoNOKBvbk6j3GGr6ef9Qu0c8yWQXACCllH+Nr+Vu6fueDGFo9R0dBXjJSl
Ar0zmvoUhREfVVu9SJKpjnxKuO2h/IuKJ3wSQ4zGMjKkeQ8Nq4J5C7avA4e7OQwJ
D2AP1hAVLvKK8b495bd3dNF1jakJL7/FGY1kQ/7GEJqNSHUXw09oBuUocgeuFiAn
xN69VmCKcOBdTYlPtGTv42BcqsXCxqZvTj3KXp0QoyqKcXTjBzR1dwEKBiX+OWDx
xNrtfHxeROtR0Muw+ZpP5LtZNhPGyF2PHSNpdy0sRG01dHz6e9KYBizouWBbGNpf
+tfMMXyYJvyKZg0ux/D6N0xxkzNXU7GzlU3Cz1qM+HYBmMd/9Dd8uqqyyk0zqMoJ
hlt+wUJ6UE6kFRpzLRDyntqpLWHQLifBI0gzVGkV8kX9jpGFWgQFPUKAlELVnKiy
OovGHNdrsvcLzDUkGcHY1Lo98tT4/SWQ+2P03mtL9Srf/kx/gl24LpgKHc4cJ34c
4L2bqGyixH1i8D6IPyeOfIErw7LVrB07ojOBZLAM7dwKTLTW3FaI5ebrsN0HZkqk
XoIfQAnERJClPJrlCSfY5qfSmHrMU58009vG+E++3XG14mVWt//yraLYvVnk9oQa
jxSHJrDygYoyOU7UmCXkDCERghl/QsuI0KPXQkUO4+CFJaYdWJbehtfTHf0AxLwq
eHnRyN6x4GpxsacLk5qU3VBE/xvP7B5Zm3yKHX5fvpI9zlCyG9LhWMxQs9d6uNJI
i8IKpcrCAkndIig/9aecn4d9NNihaFrcymiGaItRdpZWChFsa2XBxUFyGd9zBVT9
/8hhtS0JSi+AWqauiv/BYzgKmvoCqhHZ8YueULgD4JB8RvvhjH0IJlrP4+I/HTUF
JjI1HPohp+k4kmp7KNCA4JG6/L88UXAOopq1NuWRUdzE+4NW8IXEBddhDYwUom05
Ldx5xmg5wUwmd0BzfuzPfkNqtXAna70wxbhAWvgkbhtlCIMpWHrfQ0m4O2FDYF46
R3PjaFuiP4UhMDsdYQUMY0Km1NpsB3zzn/iAWQWWP5DE5bXez/GTULtU4Svb+6DV
qaH8P6rd1zWW4wDx2dfRYmuntHgXtP+Ow4DlqNWeNxak/53knmRdo6p3C1xtlne/
FV6MhUCMSrNCcDUYiqgWcUivQmw/lM+oKssxZfSSZzEmFgW7fVojC9TWJuUTo8fO
xnLCHZY65++wMbHBm2zjtTApItGx/xmgOcaJq+oCfGYROhEK1IOUIfS+gt06yaPv
6ytHFyNxqtIYTn9T45uGuJYWV1ovMIQkeViVtVzfLhSPMvMMidZlqx7HPDtUakh/
YABz4D57swoCRWM5c+kVMUa1iLv5gOJ2oQKdIdeMPys3dsKjTE/rea2RgGW4LzoC
wbUjadVIH4YKcXQd7wg2x/QApJazzIPOZDPfMahD3/1ZreiBe6YdiiYjpaQyIeyH
2zHZZaEhfHcmuRhO7Hzix0mSCphyHItTK1jpJqLhreXaR/KkM99E1lXhdgAiivrd
wJleJwwoQMxAvwKxQpFWyio9asZmUJwCu712DVAn15dOZvZ8/bvaLopzn/PSLTGG
B7o5vfiPb3wdYAXaZ6w9rYQp/X9ekzFrDPdG/qPYty4qLMSa3tMW2bmXXuLlDLOZ
EHpj9v2eyMNFDaXCZd0q7dd/sBJlqJWp+VLIJnKKXvWdjkoCPngbbABy/rxza7r5
3qsuMCL2n86Y629/vYct/bqX4FDX6UlCg1kNnpPbG9M1gWIfVucqLPhnUADdKv/o
NsqF/ufEe1Su9V5fKNixSaPxHKsVttHd9ucYoNCzGPuc53piPiMr+EBmON7wX++J
S0UikVqBM2x1a/eMqqnZ3rMqhHexDsiENnY2LuqDPU9Gh+MzfEfTwuYbDtlVZo4A
ht3g1WyRtx1HdLqW57tS3dnxH5K8xzxxAs/wURNbcLUPOhd3gCsEzqMz9Pp49mEE
V7Za2AYGzNhvP3L5vP18P4TGaSTa1CIeazdLOZ858JTCArqqebm+IZfEgPJdryaE
Dq+6rfmR3FMiI0fon0K41fyZ61th7bkJssL0hfPkN1hcOL8EUyngGx1b1nkNYRcO
VLcKKOdYfaj8c9T/Ka2NrEqd66XaHfCVuBH3TxnDW/F75afozRJ1SXSmnn9jM0W2
thj0PVTMOw23TkEiyaAWfblgUC7WTcoKntMT7HlZJaprk7UqvU7CL1WGs7ngfzPE
C9pR952hCnpqC8phGsOASfAi17n6F6NqghXpQEoPT5AxY58Oxhz9GFDsq2qIasHE
UET9SIWNKQMwd5v0e/ft6ZcpHVxIfzk7Jy6Dub5Ghhy8VgKHBfEow0f3lD+GZPY3
2e4pJMkXUFP4qBO/p3s5VkVAuJoLgw4LAQuzB+yegTbUUKftoKn5jJVPnnjCDKtb
w+yJF+vrwbSK+18bWl4GEQgx6GPTM8STEK3EMhO4m7gKhaKcygJ1GLSm6lZlWWyB
Fu+6EUDKGqY5MBwVilVOx9XvDIHUaFWvzYzdXO481mc03snYiaILVvlAB+fpwS7Z
644QHXsaJ1pzTUpsBCTK9HoiXn4lp49Wrlmyu2Dc0i+op4i9sgPDnxaRj/YyQ9LO
/yGz+L9oYXn0D5x8qXePhq1LM+iTk63VDtFQ0dcbNSj5g1x/Be81DNILqeVFQGrV
e3Pk4w6oBMYsVfv857ogpnIVEmH6XMhZzzDxYbFGjnU1MgfDO+jGwLhKouKvJo/A
JlrjUUd3WcQ1VE9XEznc1E5e1SMrxSoiQACIxGb6j5Z+wy2AOU75ij7lM/NS922S
FHVyOzjvVdosbA8SsB5LcJAwsPjznUBOoXf22n2+rIWvMESbQchK/NdJvu+HoYF+
rLwlL1euly1p07qQT71tyi1bI8ELEvQrfynYtU1Xf7/qWrahHmnf1UKPxXhCQgtg
l0RQdW4+4yFct+nDzl2Fs0sZF/ShSTfEhVf5dJaRzxoX/1FLo/GQxQuW+ioaZzOv
vX92JcRLxvAZuSj+K6fYHG2jJQOFK+xuA62eMEI/prBwXEAFlhlOrt8w82skNHHe
kCNbHQMQjHy/vZKnR8nl3TFNZm8IlsZIuJz6ZbXnf8fTLiwq6CUDVC+BnMLNLQwO
plHWkQSSFFgx0EBXQvLy6LyodQcFyFu/SnGQyk1hKvKptd7j32x74vfya26jmHE7
1T/HHeuzSfLZmvHMJrj/Oo1H8drC0DM+HXu3q5pBJddzxsQeErhg9rnXNpUZo5wh
Foq3AQyiE4ByQqz07OUIBhZPdUuVn3zgxdd9D8bDpkus+XXaYtEy0JD1XNHxht/c
RRaCRdhN3alGDzMkNzfcmv4MWcy5sgfUaR788/cs04hQV3Ue2giyqxSwnDilRtjr
drYeG2jvWMVt5k63XgUOgaocBcE2XuPmYkYWgRWGPa/4QcpSGLCAFfuPlW6/dtgV
VaM5yRND6enJrHNIY7bO3vCyQyg5o1tTFH9mIH36PFgdz+raav5TEzmMfsVeY8IQ
fMZY80mvy9cgZrDA7ITuhthKa2SZfhDfFCa7xayJjUJAQARzAd7qFlUFRMxONpm9
b80N+9egx6dJykeVyaXjYzldQ6Db3QUtFvcNm5HMu7zgOb/3GE+7cFi+pg0Dxv8U
pTR08XQR7vpdCievUdhU4xiOtj9d3381L6k/Uaa0J8MvkpBGdwW+HnwcnhFE1RnC
Kf6VP+xTnpCXqBsqPwVmW9J3qQJ8siqs+uof2UFalbz+OBdPo7w3w9F0NzJ+NG9y
Q0NRRt3reXImW0ZIjQiY+NZWMq9bizK18eRJAwUfxbuA3DjeTOFLsZFvHq3yDSdK
jK//IjS+LVdhPk1hk8Rkp9q/KvEPDH29tgcePDLB4RrqQvAdbEIt62/rHg9kMX7R
NL9n2K5oMc32KRVYlCOAczgccwPbUuz98LjjOSdbRyKJiyjs/ZnxvIxsdM4RtvCG
Cl512INdPmByfB9Ci07RYgPQBhRl/r+BAtAmzHM/87hFWl20xKzT55Xh46zufN3x
nijBlbJSYK8msaz0gy4omwLSl2qm7jwQ8xrsBpaDtZ2E73ojMguw+6kT/+luORbH
eaRob7TWk85F0T3TtMkDbGJVhUXkmz/D55cLRYq4s9N3S28LOXnSYdbCxilBunTu
q7wVxDv2zbM9L4kO+27Ne1zRivj2qD3SlM2hvCTk4XuYM1LopA+k21EG/ZZuvyca
eAYsG8FKE7F0SI+CtQXEcA4mtV8J2W5MGeWHQjuC2r4UwKxl+02eXwM05wOTbZSD
QGIBwSbAGPJDnrv5jHXCyQuRWHB02AYuZ1fcMpnJmDbCxFs6/jIlZRp0QOn64yPK
nyOlIXUtpK6H7dUrRTQqao+SVG/3nDi26MNtswXeSFBtBKX9LCQCraQUYg5pdZ5/
2tpngBGhUbgq2B3DFuK8wUhFQdJH8T6O0jfhEhEifFB7p61gpjoukshlHjrcvhQx
CUElVvLL9yzSoFRSGrNphFXYq9N2ZuiBTmjVpem9hE5NuYBzHfaa5Zv1UbMzZUmC
3qhqo6J9tyxsOND5vnqFvxx7aOBw3hYt1h59BbdclVT/hB6Fg9WlaeF9fAu+dzLN
XyIqt0knbMHG6Zj7L7b3Rc4AtByRbU7Tu276i8aQqn/9e5fMn4WJid/HQz6MApDD
`protect END_PROTECTED
