`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbFjyw+Ck69ZUEJuWEfXCjhhyK8ObRyybRqbJTQVUOF4ql0Z9Ex78YHsG0tGi66r
JaSOyqPINSB4wTtCWvXPeUv5JkPcplbdQg6xA7UZm5fhC0M9Y5FpxZP1bME3n0js
4nmFh7K29YCc+lgIFEsCVyP1dUocvG5OChwN7BFgzpdn6STRgR3QuHTFSuiVZyu9
2RIeJ78YX2gVLsiJax6p++hhSNIcelY+EmIeps5WDCwO5Ug2ZDfrGzxqzgORFzXw
lga4Nh5cIJ6P2N/9LOU0RNAnuS5yfn6MpxG5pc/ZDzpUZ5EFgOu9UzsF5nykLwBB
pwH9C2ZGidx786D57JRmvwTayJLKzmG6UzqFp3gLGS86ASXGbG2o4Q0+d0TMKgCd
2MeBfABaVmXc+3QKeCioyohf2B7NBqQswpan6KBNbnHAF7nNCfr692C4mqg0MJTX
84X8PtWZXdNLkvU+g2bzgmThpNy3ljI/eFMtVA4NP36eBZNUb+9h7Ofqf9YPxNBi
`protect END_PROTECTED
