`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28CrTTnj0NLHbIDVowVjP4PmPHFuVtwntcM+UEjrRSBenv6U4KRTiYOyXrUm3mcA
7FLLxOgU7GN/sAzGnOvsoCVaZdQCb2R5sEmpXpmRx9FdKrD8Xgawi+GjOAGfbJ54
lJmyFWu/YHlPHgFi1lGjTb3mL/qbWwJogDYk4LoZcVOUbOqQm2NNovdKqwVTuy1w
k3umaw7kBPFtp8NEeSsak77/M2T76LnOS+nNDPFNF3mP4cW0dZgO7Xt1aqNCtkCB
LLqfGFz2cOQDCUrvWuMWNxtct9f00Mti7FyNd7Oxzg9mGxXIORfJ4Mgl2B4y2+Wr
q5TzJN7zy2pAYXloVFI/pbHFxdZ16aZQHhzXjc2pVznIFjH+Qr4hnsezdm771Vtm
ro9zwU4jfdCLpVkT7NO0fTUO2/+q8sqdtsYgbi4aLihXd9aqT+UG/jK3M5Ya8n9/
jnh5DHj3q/fsVlmsQVdskwRLrbQe2p2BU6VxaDfW9YowGq8IeC2yRj4NcyyeD6KL
8JPYm0gT9Ybi/fUATOF2GAwLdtpW9eJSI32dGB0tB8oS31+28npALnOaiJ4R4BE2
ZQ7py1smbxZj8rPWNsj/ZJWj0JJRw5qMQ+tR0+AqkTCNrgru+ZWXVroqwdLprbUj
ZKREwTxH5N+viOBhjTm0uDhtluiNjso5JvYp91Va1sTIgzdP/Ma3z3pIQSuoJp1q
B4YnOS+tojmiBcGgav2bxrcwDe6PYHkMM3o+qb8d/WlysVKRJS9LuFRHA6A0WCLP
70hSAGUfKnivHfSVOyQi8jC05iE03AAzTZaQWlCoVpbmH79Dl4rkvlXhxn/pn9XX
/C75pG16SduF/NixyGDOdTAc2GQx/KU9zgeHn1bIeEEAf/0U1v84m94knshK+LQR
oYGHcPZ5O+7LDDlEW2e+r+zSp6lO8SZbd6uDy8Not3uJnZHH+ePBc/9l1wIVyRnZ
bRTZEalPdQ5Kt+hAFVxBX1B/3UVm92xh+xFRauVReBspBlT1KlPH8SgL+ZAAi4K4
YSrABzLX43hH48KZvkJPJJQHz2UzuqI663Uxm9Jlvvkdf536G52dI8ryFVpHzC96
wxcwDptsXTeMvF3ZBN2mQ0uPkWoVCaUj/fxCaBG6NiW1MVY7JmNTtD5ZRB3XMiNQ
wWbZUFYwy4yXVY28LU8lR83g9Rb/oy+q/aooutq/654l1qUDU9AaCAQ5wpZybA7T
xVzsQJeDxZLf/nWfG5AoWLhu98TCzlR6j0FqDC/DpUye8qLz0zgKXk+5TUNBGUlj
BkLgGKGBA/q+d2bqKBQzVTU0SjWTiAi9gtU6p0RjqY5Ry0ovNOS/Yfp7ZAuaJLyU
tJMxZgU7VUdcDinPJ/9SoWXvJsz26kEBzrAbN/mY96UOCy11RIefvmwTclP9TCKG
NjWX2NZScTmV57LSOfTgOc0Y1ZDkJhr9YEjUk/qRh1xBR4OdRKKP9SAnEE6HFxbI
nAxEey2OSTSA5sw+rnhubmwANZ6zdLDbblKYH9YMt5aiNerqDQmmIaLukDwsKqlD
205aK0JuyRqYniIqHrzYr9P3+YZN7nznkNwmlciHvrn5QPH7sOHRRSMCCehLhFRL
3V9jiVe4vexAcbQdZhX0r0fWGWi6YuY5fHzYuHcsGQjcq1iNgfbdprhU78nEl9qW
hbaTGquR/bvfvr2TOzqc1HFLJJFK8hOUiGeILnDZkeubB+XXmwJfkb3AtdCj6uhM
OvM6pm5gA5CkYGon8uBjHKOIGiUlMfF4K6aTxg1zknGA8Ei8XVO4x3NHA+UWyX4g
J0mgHOUYJFI4ym4ZuYSVx58xRRxZKH4cYbOs18b+LAluqs09Uyz5OWGPmChfIlL7
ygER9i+K/y3JOtb2fZBVt8wGwSj5LSuXDTX4q9UiI73bG2wYzzcM5wXldfATfXz8
/d7+9Oen6vU/AoRWsSEpIj9+xFDux7SPdhUpZ9d6NJuxpaONtqI7wpzS95d5v+nO
W8CddWseeUOTkHUkDSgyDvcuFSgd0k4qhpsvbIX5b8CZbOMMQ6okhnvxS2r2rhAt
Rg7DdOIIFSV3h6ZqP+P5zQhGPqqtVmID0+/SrtfiV0FkENz55JsA/lUe+uvczN9c
wstlsnuW7wOd5edZh9jZPafzUs+GNdao1LQqxwZTqSn6K0eehJ60AGYf5epAE6xc
mIaZHO8i1EKlXejm/cOmt6MSF/iFPB0BI4RZpFFX0LD3lR7uqtyPstmDGmwO5g1h
BsLJrQ9rZDU3CbIjgpD8dytwLxaQ7PwtRbkJdGu38zWy3fjCeB9iN8LJ5yCk7Tq3
8g++yzSeB6dtnIzpwMURAgOtV7Ai4HDMQEDQjmGodjQU+EMAfOVb8VPde2LlHHPH
/6Wwc9pwtL21E3CELYStit55x/3YfSlOXrzPAOmShBC1k/gk+MhlIhiIMpAvm+ZO
qNqjpxf8gR9HSmRaNt3SOYUOyXVlFOye01ysP/S++P3fbVo4CfMaf/y5k5+iMuRx
O4Nd1jJNB0V4I6W9EpYCuE1TJ56swiifrIB6D08CYGPYxohFROFfIx0QZ9neQsMq
8dXPvTdxjELp/lTVJfeD4DQr/tRnyTgEotxwBloGtNhQE3h72G+0QULqvQ0VpLPS
7b1U9sE2XLkV3MHSsELgMACm1R49D6J6ypR8hGXkUd+K5Rez48ULXINLvdJDzEOz
0LaTl0Lmy4JEY5I/g4TjqKxTZgUiGJWuzK9f4qdAIZfVeAv9AKyynvYahXyiRLgg
gZ4Kr+1Qt7GnvcjPW/Un7x8YN866QjwLzQTYxY68cUykAMJMfzCVbOzLkjsFM5Ep
lXCJjXm8hF0StG5iictR0FYUIkyJYOi2i4Pp3YQG6wMlSW1IVcO5m4ODUHz4YWX/
N9TQXgcYNyq03//kch9w3AgsOIBUY890hfq+5egxZFEHu5E4b4OVKCC2nOlu5+KY
uf4dwY5Og3fjfANIDnuHa73qnRQ35S6An/a+iAJMuR9DIZJL1aQ+H+7qjzw8ekvh
UTXRFiC0/IIZKZkx4dRcCBAlW6ZDc/cozK8jC5hiEcUMy+R6DexJ9o6V0NQ+PP9a
0bZJ9t63u7llkY8lfKCIH6cdgHRzOL/YtjF0fpVCkYffipuhSHWTtJNTZdy7MfkD
HJNmBq5kspD60lmWtj5b1yvJWI4//xtW62WzNM04JsAMtN1FD+59UzqXeFRhr7hv
IA2ZmU2hdQpseBQ9xdRvZhtHyRMoGvzwP4ERRnJ2JKB92XPWLQhTtDQXKwbat7Zt
+kMabFbeQs1ZXWRwr7vSIKsVtbnKiF2w+R75xF8Pm1bhOP0EIysb8YdIAeeDBMcn
Zm/9B1jW25ewrzsYqNonN2bJfhd3m8zDlt3IENQyagHJQEJPcUkDWeJ2ZNPsXOuf
XAidDQ68E2Bugdr8qzDz1OqLFAJKpRqQt98caiRh2bSKIIWziXYa1cUdBpS9j35k
zYqjEu6w+aJeAuluJFSEVBjk1/C4GEOlyuVoQWNnkIwg9YwozrSiIIni4GdsClTn
ANXTf1w7ONDZm94zXUV6h4ofg+W0hG8bYhV7OJ9sHqrt8C2JCRAL45WRtcc+3sET
qkdpoi9R2COqbJJri7YU+pDIr9MuSGczebZBeh9jQvvQANgSbTQPk6BE7npDDY5m
Osxe/AK+kbJKvOj3/oE0kVHtwGst/tzzJVCS1SZF9+xVS2nIFeA9+7GYVraJCi17
9Y17Dut5iR3y7TR3iu7UznOrQltS1mxpn2zLoouRzuqHZpLbH1YA/49TGhy4TTBH
cHkL6i/w8QjRB2Dmmr8G0bO123wDCuaCPI1hOKmZyHypz10E9YXrteN0RW/ariW7
Syb+M6e8vQzFjxbuA/DTK94K5je08V4P7M1LtsuCas26KE8dUqtp9A+3L2QaKDJ/
ye38AkDYOADPTR9h3jxMorB5t5iemTxjUp3NyeIBCkiDCkwvFx6hlB8XsV1jnROL
b8e3t+RTSeTWU8PCN3NhIA1QL82SwE9ovOqMaIsViSNl9W9akCEy5iLr0YNCtisx
cw7MmRdsHPkM4Lyu/KHKk7KE1f4D8+atuD1kvvg7EOG7qmyc2mluNpyka2U1GANR
liZXCgyCp89wFSS7q7iEHVpD+BBfQkXRpS/MT4EBKHsMxaDAHRuC96ik56HRTy4k
p3zYSFDoPa6dxJcF2oxhlE3D3NDEVJ8elLYVc4ZNTn1MM+p1RGi0VNtrtwP2T7Gh
XlwBkBzAKzUZP5u74URNISS9D9Odoek7aOc21PnpAIzNTtCGkWM0jFQhuvNw4WOY
/B94sWwPPjn6/s+e8ZGWN+1SfPfMM6pvkTvXBRYMPwh1mbe7W1BvqDlrlvsUaFmh
OSiPepHhiB7KPCc6EbVE0kFZYwMDzeWO6/0ZudOx3pCnmvc0qZwGxHhRoJlixQM7
WFkBrVTLKnD0NiC9nz8uTHaIwz2u1PJ53hywT/oTfKXcpOgZiJXaso3+Ekh11hTg
78hGB3ZKZxg18ALFou41RQG4P0o9RZ2904dYotEsk47n0J9EOi7tamCYQS5FYYIz
kZqpd3xpPeiXv6MmF7zolap/IONinUNUV0DmMVwJpVYnYcELXstdZRoyvGYtpryd
HFavqvXYF164Hnx65rcdt9Fmi9GQfNiVwKZn2zPjA8LwDZeTFhBKs3qJ33Mj7l4s
fIu35KHFepCeka7GhOqvzpE8QdYBELMOP+24Ygn4qpOIqX8RgZEh4U4S/HGZ2s7f
F6xy5zZaAYE50diI/RLekWE+KGMsME/nshe+KVNdf5dBPywcqVhBHmEePPWcOiTa
XUxYhZ74KrblY2KfXow5UMwSh2RAodOyDWkkJl8Y+Tb6Slt+v9Fu0DCV8RccyR3q
D8DiIClc/bvTHmJBV6ch85kocSKxMNah31x4D9/L+xQ1lorbig9UGozDc7Ot3dMK
92dGNg+nQrjFQvP2Wx3D0Hq96VC/1xCYXBTZydVxaoOE5Xi3c/SpCEGneaVd30Zq
SMEQJdyrJzxZxvEMajipa37MlLz2MOHeyPqrPMB2lKSC7WmL76pYZU9mlXuPNg6C
Vtqa4CJ03Csgn9UrbY+lPfIDZwX9WAwTmTFlwa7MywUOLRTZ/sJavpPhaDbmj9uQ
/g8wskumVdgl8EZYihr0mg==
`protect END_PROTECTED
