`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cesmPbHUBOCz6WDj4rbuCMlxUTStQ/2Vrll2EaBO3UXDuk4ZE5w489U5IfhgxLsH
xEHuiOZ8SS4yD2j/8xj/LZ1S8OJpUil3y9sgWaGWsrc4OZ27t+tWg8Qh6CzFQh68
zFUNsuwj90yatBdCxsbCAPd9eshk1chMda3Ib1jpiSb/+oyyhzlQxmkHYZ+UqL4z
SzxCgupI2eVt7FxrnuqEoEcKLQGXWFmJPrAcEDPO0iDPTBWcW/5/8PffNHX+sqcJ
yu1whBS7debuLL9IpJOkakW7r4cTMi4ArfrcQ5ZbeAm6i4q2BfMyYEH0FAHVCKY0
WrqUyjbO5yEIzLs7mDb4QENPh4Y02/YTsupvdPTzpXDb5afO7TPJe58XXovN3qe9
vAS/3SWA32T4qjPpVzmkdQ==
`protect END_PROTECTED
