`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbJKp/44X+t/NF/COMBZr8DI3CJ1GZsd5b1PAYJoZn3hFp1dU2GuZu35EyltCJip
kPUhRRl60dqmn4Mr3n0dNdFEMz6Hjvwc26xgaeXDNzT6zAFjUpwFkP3g3hv74iuF
Tz0DlrgNGq91dAeDohJcfAKRmubkp2agCfb40HjcLGKxd49iQdlDyP1sne6ZKJBh
m+lQcbPtmWZP4pY8ez7ykBsP8qMErg02Wqrc1lPS8gioPylEv8PjM4igbd4NBYwn
PJs2SuPZbScZjXOhoonh6Lrn/P8oSiC6HDwPj2J4xOtvCUvWSmACmzzGPwzs2dMD
vobLDFyA3bHJ+begn7fcF6rJu4/g1e1SNUPfcznOGbsIP9kevFLCX/uInc7SMm2f
KRJwbelj+HCEmodPWAZMNY0/8+jbXWLjDY/zu6TwLuiLvcpz+0ojHGU+NSIRNbqs
Qq9dvdzVUsl+P4gX139NDBASMpkc873JdqwKyaTEPYBAz6Spzl/VekHA+TaAIsRY
Htq6/fYO114Ofek/aYxn0qK02HZakDFOQsgIQQ6lmsK07s4NwBT9sZGPgO4IdQHq
ZZqGKQgGyZ4+k4kTAjU+WdFUBrEoAdelO05T6p5s6hhATy/ZkHW6Qq6aizm9x7U4
ReJWtH50O0HJK3KQNapHLbvRj/YXwvIL2XDxGz0hro91Z2gMANSJ1u2Rtb2RQgJy
s0KWizv4tn5/2i3flodTorTdw/hEEVP9KmwSK3nqy45eS7aXLNbY7JCZ4mgATDuf
1qRQ+qgS46OmZ6IcNMBaMFrL7ARKlaBtmUt0oXnToKDYyN/B98yKZ57yOlwMaMcW
1DDNPp9OI17SqkURCo0jcWaTC4AJYclXsuBidEBAhFn1Et8/xlirUb9zBq3cH/dc
1hHhy4VjQy+hjTXkCk1ftXDOadEZ2GBzCiKYDqaa71Pi4PwXE7Ar97qb7gIosE9w
o9VEFDYScilw5y8o/U+ZevLvbDhGAqEG3c0uHIUU8p3DWKt/KoRRw11EWnPrcnCu
VAZ28X0qb7zgp+mYsmsP/Dzhys+smVl3CnLW8JK5y4WSBqV1ZoI4C1MBtEYGSVwC
foJKxn3KF6G/08xQK49cAulZwrazejGAYnyUQSBsaOn5Q4/zJtotDfY1TbRvyo55
Xxwai/bc+hxMISbafdQmAMB8xlAoxxRFYBllBSIDnij4SyYLdvUmvqh4X9PQIOH1
aN46/Oo2HMF7HBLm4lmEFr/6SZtm3rO4uPy1XRkwBa6jqDhMmxgomf7IqB2YCLMD
fLW89hT25N0EWS2amoiBrNQBE6qGDLfI1jsciFeXCghiPtv3YiKL/ikrbxt7KbdV
Cvur9a0FTU/gNXRK4NFJ0iU5zmiQfpjLCCjMQLTtegg=
`protect END_PROTECTED
