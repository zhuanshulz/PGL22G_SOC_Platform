`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/9XqBPVS53LX/chVr4E5mbMEd8Urc1It+z7ooEx8XD1MNRADiZnxsn2DrEXDGxex
/78GpthrqmV4BCyXKi0iTNOWwmCJIJQH+zZtm3faEV0Idto7ow/lPwedoHUcEtVG
cnQ1KOS/tjR9Tt6UZ8Jl60u0BXRleg1/JWsDV4+4d8fY2pjkEL3mBUXFDW8KmXEY
I45W8bNNpj0pjZEqZRZUA4nbNInQeQL4l7Dh4GuzA5QdXoICuO6TrNPoCKd7Uebz
dA7bZryO1+gK5ihYr/fPHXBXsdaBa9oPPhlqOw3NaK+Hz954IQhhP3/kVsr9ddiz
7w0l2d4cJ6gYPR0FrJwUfMTmv2Jn8fflrcoJSVv/99hw194teM25bz/sxc7IffeH
3wNxh0+PPaXj+xSmhEqi7AjDyHxj+SQRQv/hg8lIsuCRWgQpDvd+7QUvVzYpqAJn
sP31uWBP7Zv+Vo/2XhqLpa8PSuZwsoCsM6uOmAPRo7dLvjNGoECWQtsipxWXAw6I
JoHOcexJDmqarSbWU+ck9/1/OKOhxTlqmidlLZzp4uD7bJEAiKamcaioL1/7VLKh
oSdXMAWBRaVVzCK+LMesNvGHdBKa6OP1iAevDkZwnhERslA+GRTSR3vwlC5gQ9LX
M4TgW13aOFN6xANP7S0Kt0/rO1dg3c22NEJPaD9XaCM/xTm9l8NQkrrgHSqZotC7
TQWtAilCbJMWqB+S1nlcsnkPN0rfl1O4GsWIkB1glCxttHj+qy8Jg+yd5BERcF1b
pV+RGwdcUEQuqMMtIpN8Qaid/2g0w7JDQGNgerJqm/Q76k8qkte2dI0eDdildUhM
d1ZWnWw1ojbodCzqKpid23n626uQvwn+7yoUaew08cWMntZdJq3OelBytcTzgcAU
z2JmlL5NbhRAy0vMaSy4hIo5NpJ6Xis21n0A08gprFO6Z4t9o7+Rt/SZWYMHC/08
QOcTvWLhiFB5Cua2M9izsqnHwG3/CxzV697wKb414b4R3O4TWw3248jmYS8HUqbL
zqg9BOB9woOQPsfZG0LHXeF/HsbtrlvQTa1bw/F/HbpgILfAJGe3OWmYgJwp6ZHY
VHH18mOL09tjo+8UJ9aiohMaEoBPd1K9Osnobc+jyC7qinZhZXnLEnu3SNS8mQi4
nFeOKThqEcYSOpgkQA4LhZTXGjDbAue2dGpBfICXjMHiCAj52sM2QpmdaxfdbbLp
MX2st31dSqdkxSdeok1n8dAH/hCh+ZsENuQ20dAoIjQ3YopaKt7dbSUtphUkRd/L
E1Xr/cznLhFvi3Pctexm2TYIzU9F7JrluQAfHOVZEZpXcYbvRmNRkRlbbBl5JcXi
vDu0kSnYymAUCjQyvNrDBwboABX4vaCmx8iLlGUVkBBDjIANDsgQPDnm7PfD3WoK
oCQLS6C/pGQyWT5UaNQTvaDhrO8YlJ0fLNEMpinBdgInHNtHgZeIiFwSRTivdig0
ZVWl+67SLKRq2/+5i2syP+yKfchDLkK8MFA1S7iNsNjVHK1VcXYtXKgFmZd760mk
F+LhuIfR3pauCanlHlT0tamAiol0aAOipFm52BudoEiQCd/cQJNDGPh/Ls/atLoE
aXj3evZ73Uog2Vgn8aiy5Z1gwdaEpKlwCCkwvTeBSW8g6PggLd5z/iLnNV5umMDt
Nvy0L4sRJzCFnKnrIeNexeY6e3/NEyLOfai7bOIHpEPG90CrnUAkOIUnj+EpFWJn
v6g8MHSv5cRZnW6WFAuQwysRawNY+r9vqva3/7FsBqSod7GnMtAC1aNMysZ4Bd2/
u6XH7ErdW5y5UwvRaDLtj/xZHT2yB1JyNlAbF5+tDqKZdRK08upQmclT7AVEA6or
9ZzEsuF3wWYiNuz5jdhqYsLkWFxVmi/TS3i6V1DFqkQ776wIHcx1o0g6oCst7p8b
MXihYxzCLI9HUz/MeCuHinU903x9VhkJ5047VXhMkBzx0qYTctwTQfmjhDvujPJL
WGWNlDZD8zn1XHpHLB5FcUek+7upZHqCkbpdJGiPxGBs8UIJSjQEqn+1qxubybK/
/ZDgj585SASmT+4AsCMbe+kbS2lELOZ9pLt/+OlPSLJFkYIK9tBeaEIo2XfQd/4W
wAV8TYlMOuoOmqHCbi3HV5d+tfa4Lv4BlkrjpQMWqmhTw5U9OlgqE/O18UMg4x95
pErkL+qc9ijAfBeg6yskAZCQhQkHX3bLwVYI8VV4Jc4VrskgVdusFq+Qp2CNf1VE
H6t1DlIWi5wKNq+T8sW82aA2WVyqSeDnlS7hSL+MNxg4pqUiwqdPkFw5gPSqtw7v
tskR7o4xGsAGr9l1ELOytfoAMZZslQwlBllIlj9uwnBgLveRMwvRj5b3IjmOdHK3
WostXcKYzOD5IqEJAkhuL/Bkyh9WfadqUdmF5C4SwnDsFhl9WxoJ/KNgsKPOMHDc
MkEh2KO20c8athdpNe4KNMfT8hFDp7CTdJPTQd9ubiN9guSVN3Zkqcp69YpkG3YZ
3slG7r708camqAREFx2vyKQEx+dpd4lkurhO0laPUNMnuYkeKni/y36VHZFjW7Sk
/zpDAe+7/E/Pq39pN5MwsLYiKwRLqo8B/5Nh+R3OLT76C9bGOh5ZJD6tjT5pg/Q4
9EjfiwtTR4SZFGGV1+NYgh9vM/AGZmhDs7ZlJLR4vKPf2LzluKxb1pjIEbOo72lT
Gp/a4XzXG7PE+0esqp5/Bb2Ay74qR8NmM5NUCGwnF3bp6jL2BRWa544Z8b7hPKP8
383v/piYk5urrGxk4A6sXaHacdUAGPG5bDXz/Q+hCPT2cRDu1msXpUfWmWXY64AW
iacQrs8SppP5Q3G4NA+GZ8NAZMcTs+wg4C8Yq7b/NZ62q7evY8E1s+QVOtZOkkEx
x/tOvTRHtRnSr+YucnLiCA==
`protect END_PROTECTED
