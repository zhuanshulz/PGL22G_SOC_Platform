`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JfabrPmwPi7Q5LfEtJimZrETaBe7P3rpy+LofcHGFG7Tb5wcqkcJIgZtPSbgw82P
C+FpcWfBjNHSDdis4aD590nlNFyZ/Od4rdt143DMlPDq+dzfDNGrYFJvKSYMqgjy
v1Gnl6SBH2Suqgpieg7fP44lOVT8X7KSaDRx+toWBZrrAdWnsysMbAd7h+qCGiRk
7UXP/Teo40+0azaRP8ZNPOdjimJRvcm7VNzf2IYmQvTB+Y+4LjrvjdUsLqJrG2DW
Ya5gDGyDaURpU5d0lCDoKlFvIlGhOsAAEIjekuRFULvAyQNqv7GyKrIi12gxzi7q
pGhDuRs+OCRbenLeYAjmOKL7jEU1zFivd2EAqT+6aAof1DZySs8CkjdgwhWo0HYp
q+zkQDtZeva5sv6Q8CjyCCMKlGDBIQJZNP7WQda/aXuKJ5Nuql/5ArHmvJ/Ep86M
OD4c2qSiY+FffA23e4WZKexjAAR3N051nFRLFXILr/DNwZw5q56xlQ9OMT2wrozT
MRBPWKdWkvs92G6A/ITfPGO2VMLMwgE5stf64YEhZgS0GzfpvBWfBxhaoK6H0Ubu
V9HQJY4X1Nj4ifI6g3ZVwg==
`protect END_PROTECTED
