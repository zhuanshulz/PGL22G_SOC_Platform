`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E9DvFBhFgnvtTjUB0lc02nfgJctG+GYMDaf37JvA1v/zwSZFz0ypO22FXSQQXQQk
HfcXMlLGIo2EiGxSccQtsM1h8hhyXKE5s7AzG2+HnTBeZpGG6X6MlW355iAXYchN
/4rJ72k+N6PiF8nVYvokU4YIKacZ/Dui+yUKs6MNJxsjGJV354MSw+lbmtxaxuIS
5hAlWuSEXPRNB21U9pfzcZBRX5/X+Hdlk/wYtoX42xPM8JSLuoi4J7cFikRJBKnO
svU5FQsJ17QDb9aT5KJ3G4wh2ONqiQjmuODYEAantNGZ/kds1pPcGe4HDaeC6mYc
95NRMDHFLpRBt6QDQEgcCgB1N8u0UlLjgfhLITzpn7Yo+BeaGPOv+4ocvFhwwqJX
Myo/8eWFGINNwlgUX5d05kYNHv71NzxjlOG41NpYCytRJz0fxhazjL/8ZbDe9pOP
zupQemlzPr2R6zPDG0Jup3jnqOTnnFiZH/Tdk/TvhWgJrECaDM4qGm1MZ5pJeikt
vBUwFq4JGw3fQ2nfxk+yJHn4pT/6Sb6NMJ+pbmuBHzTyasnVtO/ztdoM3jPj3OOI
2Jcv8bAMGfE/mIDQ1Gleb9ZMz7GzKlQ8ZS8GtNR9QlweVLZ9oAn4zGVWJsKbTaph
Fwrz4uax3Kx2rc2vYMfXCg==
`protect END_PROTECTED
