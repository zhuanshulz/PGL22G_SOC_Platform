`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhzJYymJgrmEaS6oOyaNArkHkmLrAW2e3it2QhxP0N3atHHtCi9Go+DIkU0gDXF7
yc/33vsu3x29tn2c2d9mnqTxsEuiggUVkPxfrrhxPZHm/vPs5loop6lzx87Y9Z7G
wdd1qjxJ81zyUMKsFLsUZ9hsdhx3zLdqbxI2sDpJjhc1rzURafrLecagna1jJwsu
0fPLAhNugyVJTY0EcGRTjJXQhdw/kq2295G09Pg8u1HRV4qkoelaSQys+FKzYI96
PBmzB6A+EveEcuKbqn9cZWlEFFZ68A1bgndFdb36Crh3PXZ1SOi44Cc9l7SdsS/X
gIJba1OQeVoBNPIVOQe5qui2ph4cQYqg9ZocsTU1VPLm71mxiJ0doTbYi0KUnqEd
WWrNgfr1NZCt6/AsKzEl/HWuW3ffW4C1i3NlFa7O6oYsNWqW6FH6Y5sR10pdu1/1
JYpt1TaOqIAbPVYI/ks8Redhq+4NUo58gt8Ntkeb+iLGTsSYa2eNeUiQ/gj7z1C7
0+r5MQHt6LYVaSafsKI1GiSw2CiUWintoRs+r5bpZqE3ZslRsdQsDCwdr12rNjJV
vtSdLlwf0t+weAJYtK1pTwkXr4WlfTA1dxtS3YLvF+ODu8N35JXQ0cBoiTqXKRZP
9EowPbi7DYtUCA0d0Cmb3OrDLdVm0D4++zxx8xoFgeExt4rf+EIcNfA1UoFQw5hm
vXgs7z3KPTjrfxEtta155sKidtYYKLU8Yn1O5xX2SGIoqmk7aJsnCDE7gFYuxyHd
PUOYP8OPntmW3wKOnlhptD5gquMe4kx2HdGHat7DzUBkx1VA/oHJ2EVXFCuO9lj1
RWzohEfC+EwbIJvF6PEZ5LYTc/Tnl1vitvU5jxBMpsNHYx/z3uOj0QzbLndyk/c3
4obZsDE8riJw9JVOmm5e8R5/08vmRmhUMomwSXmKmtnkQEBsrgVQtw1G36pvsoxf
DUtfx15rl+h5cgXzYN34VhM29kIEIKQzMDHvvHGdGJXewvDq6a9a+nXz65BJwz6u
dym+7sqrAP0obve+S5iS19Csofi4YWadT1vxxEVyLMD/Ev9vjps6B2vMEFofSwKO
nhgOOgUtTBq5lo6TpeK7+KrornsH11avDIZnoBQE0YUvKgmw0ruXT+hqKIXeszZk
4805J5M5Lu/rwtjyAlmLBBN3nPsOpoNKBUY3KNY3gKNyab5D7QQb2BtbEsPhJ8pe
`protect END_PROTECTED
