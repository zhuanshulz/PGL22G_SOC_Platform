`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fotJH4ACQ+lm5BLNhyEfHgt7lYfF/+aDrQhBbMr3VXiZOZ0QxrY9cr3ENNzyq10G
ldtIsJ01g6FeGKA/yCEWOnWlo4Cs1iJOjnrSbCxFa4I3/310V37YZJLaxgTy1KrD
CNH5ivGTO4itDSGbx4q6jgNQVcClQNWpQXwnWby/WuA8IkJXdOAyCwjqFc1m53+q
l7/vS6cLbdTegR0Hir9ewmDveQQYLKsHyUUMNZH4EdnVXw+dTLL6AMvLbJlm8nI+
+Kpnep5wHOsJDNDEIowq/EaxunB4zt/b3WJkY1sSOB5vWOJdlYy3s9ImKXz/9V8d
fBfJ1kPqzYvw0WDSwKb4ZtFx6LkKduDYGJLLg5Oxd5vFgDU8HGO02ZhwkaFAHMHw
n1pxYjP3Eoym0teHaFVA5frclm2xeUbLXvcnlj6EoKOYSBafxzvwI+ZSvqtys8Rp
JflRKD76+hmxnhRZA0wTrQ==
`protect END_PROTECTED
