`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BN+EHVf8X3Pf8jfyKAGlGfrNYR4F4eqgTcw5GVvFz7uA/AO/o6d8CkjKRB68939v
xedm4cmF2UTntnRe+LPl7ExDan7KdivBKkCws+Ccn9IUqqoKYp9vQ+8bPFyL9Ip5
LUduTpoPKqqkr89eV+X17nGYrp53V2Ye8bnnr+Wj2YlOp0sk21rdzrfTDDMAAnEe
Ejs0mHM8ghaL1vXyWHLGwESBOStgaG/upZcQ2oclVljiJb5kAWTCQFip5UYoaGCL
KsELVwv5juxHrBCet4MVM3DYHwNHkoM/3QioJCPcuGeiF/uYJDN9dfysHUgOiHXd
4wkz3I5/2QtdTiQv1kVzHwWkt7I2KU/0zxM/8paYErGZqnSbzOFl/OhOPe7ScPAQ
dn6/xoVXP6Iaw7W9zdCFenYJ3vipVYeoWjT9eTj9ZwwTzfWSyaV5ue2yW0ecXH/h
QYcF5IXxHkuPPmFYeHcmXdxvgr8an25xJ6LOAPdUhUb7rGBaJ2lVJdpdsTTqDYZp
M5sNLLJyzrp0vEvaRXFGLiLKkLMbQ5zb38/r82AB8qCdq1yZNYNxJyNfoF1xomiw
u1SQgmrN8XjtgdgNHDGNGvk2ZoE8SJ5kdLe4swxT+melCF9QN+Hgrx0X9aTMyADm
4OdC4nniOvu8ls6JODM/KdrWq4B+WcPO7fGq7CLQHWEqNqb/SNSzpLRZVMWQn7Fb
of6B25FBP0j0V85Xkpk+mltNqeTKz9/JABep8Ix0Tgubx6FQF1p4u2yIbv4VOVQv
eLV5yJPHd1RvQCXhbXuqgbcjeDkcocfJgBzUfGWQTMQeh00UOWjMgk8NYl08Ngw6
mpLby6qecbJ/Rb3OVyct648jLlOeg2VPAOOGS9Ucdm1raIRq95LqL6bTpYPpKr2g
XMl7QRlqMhcQMfKuf9GbBUGwqrwQy+lU7TBklCJkkykZZ3NJ9nbGuDbwUC6wNXuY
aSOZ+khdk6WOvVWIAIr597Yj1v3LyPW+Y+neMIvshLyyPiW+xbOoDlspitHr3/eL
BGg1aqTFYKhrRUVRlxB4famGA5loLrI32C9vjfpgOfBa8thKU+Vi/fHcoaTtHq8O
F7lOcNc3k9vW8e5jV2MG9V/3SZ2A90F226jVX3u+NaPMoF+I2tgMiLJQ0xpuS35I
3D1B31dIc5TtXgddu7Dp/uLu/OHqTLCsfsIqxI6n1MOFfmNeWmZ+jzEEcpMQx94j
tUP5i1Jy+SWwnKNjDx95kJdCj0YVstDtGCExQtXr6eXDwX4dqfBs3M1AT3o2LDK6
6x6UKfNOm4ZkWKBW0ERmQYDVKA0lTqJ9OHu7tVZ4MsYIACKA7pcopMSnw7LWyWaA
8i9e1VPTVqZM4To62hUBMOAZo84Lda1w9MHl5Hpcb8fJ+AgqNa6/Qi8pwpfRar4Q
e0HiGmSXNNGhV5kMFYsl7MWEvm6UjshDmAOS/VpLzrAK4UYrCWPbUAUYjcS2sMkG
+tcBL7d9CHqi1LoSmC9Z/cx4T7i3xxoAv5kA0siq2G2leDA3iXgxHmVy7aRhhymn
`protect END_PROTECTED
