`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGU9yp4viJ1Fcl3BIlK1ZpzZ/CQ1Pp0OhguCKrTIgeT8Qml/o35zVsGLVFa/EyOD
Za7Fnvh+Oo7Hoz/5vjMXsA+C/TqY34RV5P/RDPxGWuy8SCJ2rA5MlP+XGYWHn5Xq
K5UIIJ5UMErfo+tJkYDgJFQD6BUnivDmYu/XFjXoMtciultYZTG3+SyR/RNUdELU
BAFzLZBwoohztRJMs5VtFze6W6mCRvHA97QZixJFzlK5QLZsk78iJidoveWiJFwn
HUyvAYGJoc3UhjSlMeQKuVycx3uBj/TtzqDMvMbChJLjivBZ/0G4SsWEYVts0egl
MSIXbFxch8ZPiQ6u3Lz+ufODwtDTkve2vvey4xMH56U/eLoC2agC4ZcffdUW3UkJ
A2TxAAQsoy2bEFYEzjJ7WtNGI5D55bOTnuOMQUx7aqzLU/kXkFOUie7cjECuqrWW
`protect END_PROTECTED
