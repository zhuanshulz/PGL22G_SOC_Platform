`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WlGTOudAi8nIP+1H0WLwMdsevlCYv6hnD7343r7pcX3G10oqEs0kdMzay61oRm5n
ocsRTx2KV3Re32J3r9JyYrt1175T+AcOhWzgDO7iZdrcjUTYXURmXZdZV3eza4Ay
EFaVU1UbZFpzIRYuTe5ST0dBfe6Rq+v6grhaaRP1rkFGpPu1XBmq7eHk0uAggaKk
wPPtrLXVaN+FEiAPYbKdunUgQvFJ/51wd24cP0c+U0V2cZliEmEN5bLn/rL06aOd
ufidwwnHAzruKP9Q4gAJv7MIzfqWbQS3a+ZBtBmGcweLvrEauhrnegnAJ0A0WYJy
8Ajz8HsDoEhpFgsaDcYXYwl23p/DyOHZomfNBmWXZ5fps3EwpYCt+BkN1ebEADgK
5Bj4SpKXqWhPv8Wt0Q4C4qCN5taWrUQKRbuG8h2qYkYKM2VUl2Ow2gQeKs4km94p
QaKZlKlTzmdVT0e/8Ny6OV2kYDVAUhxT/TTCsjudS3ZpTFymFttrRSJZQ8Z8xI5O
5RSIsGrpLDyeN2gV7rwr/FN3RhAd11UIXBIVBKmsRvMMSuuczQDWpcuNQsbmlbld
i8nCENkDlc88eyDhgaMscDo3GtPoQjqZUV+q+qWZs9N2RMWRdED/KV1pymNJ+XSm
Ws1axmaHF0EwagyaVfCopf9EDM6BB4d308BE7WghqBkA0y48xCcnPJQ9rvI5axEU
C853OGLDK+AR7FT6uSdF18VE9NYrj8Zb9yGWRtVo38K9Aic3sx13bn4fA8qOiPN3
fT6HjT5KS2W8YM1s6CDuTweaXhW0btDhGn6H9xLoIC7KYfhfGVQNaaW4iIKf+mUy
gQv3i2d6KwtRLbkGLtqhiUjGS0JMqE9NvqEYaHAJuOBTZqdcxCFrVpa1r3uXBDVS
2APIFTtuOFtRw6j+zxEhoACtKRhq1D979a63C5ne/xPmuYnbmHnJWc6bisFBAeME
i2YmGjZlu2bVwNxpdnABxOOI4S9hCK9GcONyMKvvO5bRbFEGsd8C5kZObahD3+rv
Vgb8Kqc/lbBC+K/WXVvAVg==
`protect END_PROTECTED
