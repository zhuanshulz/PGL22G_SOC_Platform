`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPLhenzSzTRU0Psj7hyen1VlN4afARl+g+CN6zlfrNwqFrwB1UnSGvG8fsCkLIFs
3Esao6sQzwyOpXsceyQJx13C2JBbKDVzvA6Ah41+n4SV+U7q3/uSOmBKoI9gj8oD
kZa1v6XuntXWV+EYeckEqGenx8n120oAYa5VwlZ4CBM92j9LsXmZYQTZcX1dnTne
GeOBj2oOsQ8TSP42bbAnjZxl3XLnpxtha2E57u3EieRiaRuEKnuIDXON/A8kQjMH
JQEfuv1AjaM8CcHeLM+dQLOWsihtr7XB4oj3Jb95Jm12BhI4+ApIaNo/cFq7ImKO
+RkgfPAiZ0zNaun6iK4WIGHgepesDof7ybO4i6EKpt4JTQhl68HpQ0yz68WPjQXo
8jTpJw4ErxKzjCU7w838frCLnwLbcA14g6Zv9+CVB7ZN6KV0YHJlKv2T54aUUIy/
m64GqSXATwReTELAPYC3xz7Gk2OuKqDE3UBA9gHEBsyQwkVeI8AdwhWRarE7dN/K
6oLkVgZ+8O7Mk27fL8hPjfCS9wX4TtU2RJMzuQQTfSiIA+fCKo21KZ5Ne8K+fB4o
uZW/noQGhh6fU2GCWvIxWwssgzjEgHIO42LRgrjv6J+j9fhsYL9VuFtjno4StVlw
pBGutmHQfjgawh5X6VqEMtBCrXvL2MlhQgWhsNmINXKdKTOOiz6CXKjK4pKGSaKc
I4tZYcWaVaGiLg58peeIJKqTrTvpeo3fDrCSrzKviIQ77CdVjOHAWip7pr6+frtO
PX3rMJEFcwO7/xQxmw77vb/mUbxqXVtxfPGNtsw2FBo+qg8Lz41R7OiHEncumXsn
SbgGmJ0AXvW5lsS14Dh4nnAfSD/m5I4ea0RKFboOPH2qQVq5bvlekrwD8t99HYcA
XI93kL5FwnXbuBPXpPqt/W0o+E0izCJLNjFRBffolLwdaCnf9R4FRSulxldOCOKX
JNav4TlLxZWCuiEfzizdaxYgwHH0Akc1y0kgEakjRG7Hxdf2bWfHJwNSBRmf/QRV
HMyKkBU6oXuKH9xnibKvb6sDABhFSBOFIyDUqPk1hq9CrlXoDR4x7wFdnR6UwWgH
Ie8Ffm0YcbLxRLr5NHzEL2p9VKjllkoW8dj1f0LC9nGijKgskgHorqfzUbhcuiZf
VqDdaqPWVv3XNawTsaKw0ipWw3ov4rADuwHPp2h3kcTJuW5iZewPPPv/FwIfzAe1
cZvOPr1qQB3JniQ+S3lcbTU0ie1u8kmNS+g9hm0KrGC7PQCbxBZ/lNGOPSCWe1rC
ddFvBGyoJsMwjeyG3JOudUkRcZ1NSRtqZOJvdsK6Si6AE8Uz82MS4DSiUCkM8Exq
765GtnNOjcdszx+w1MT0CY9dcgY0EsP79Dz1O7kqnT5udUwgS/C8fkjLqrhMkVmC
JXBPBpqVlu1ZAEx+f24f2OdExziKR76btZ5cSJ0SIaDhJmD1uKuzgVyax6LVyVT6
k3GQNvpY8smIYJjswEgRiPobqWH29B787LLmp+KWPWEZMl9hjDupCoT7ad8U1kgs
gDI9vbsgMrc/hEvqTzytsbZn6LZIeq48AhUzq8oXYAiJEJVDoAt6smjXIIO/47rz
DLA/f96gGnfZD20fQLwZJClBXNv7nx9hXTRsHaAVB1geYR4TQpvRnZ9aIv//458O
8+/xO31Bh129kNiKu+uj7SkjwqOVAZADm2A15FwEeXF9l4iUSnqVmf90Qh5A+Csh
J3J6fz/LouSbcRix8hx6k2Ref2FWsmfG/DqFY5/CMjCLTX1Z48O8mj65P/Hmilb4
AYDuV0dKasBEY00XaFJndcnsxhwAK/nkmazAItQuDuqL69hc2vwYl6xbsJc8iJWQ
VoBpKpzgeb/FE9kbJZwsEO12LJUMtbk7S/ZwPbbU52RXCsrSrEE5Z2L6cQvMXnT2
xVi1g/XLjOVPvoX2AeVWBJTixbPJLzC3LSufCqVYF8b3A6fxhni2KfP1Zm7Dmvlo
vkTKDndyUj9r3Jas6mwJcxmq/ZjuR93vsx5LGkBLCTzn0gbuZD0XhIiLSIRiVpRx
nrK+/mKgyhBbYrxMdvjmYSUCyi2+bissivE737Wv7UdEQLFMX+OQHLqLXOzjg9g/
Vc7uJRFsQRnGcwWymlzFW4e4CWDkxgMEcLVd/kgVzDTcS7GP3J5zpIbI6uOIntIi
ZOnAJNFmnxfJNfRte8PYxMgTbCGLQtF6MhbLUA09uIXuPBWHKLg93OeM8k34poqS
kJUiNFWM5I2aabzt0tzoE+7xhUrG3Oiqj6SldZsIM5zAUa0MpFFvmEreS3AKjx07
Gjka1Vh0NlVmFe4sbaZ8994HCvNHLutM5IX1NUM/N8YI5y4i8V1EFpQ2FEfnbGMP
LbmBdgS3cVpi9KWgofdnk6YM0dB15RlHoPMljzUWMOPIqhB5jYnm7zeBIIY+ukXr
QOX+PJMZWZRBE8WEKdgxxxd4cH/8ynVRI0jUURsCgan8ruhLJrM8Oz+HscfZEOB7
+E8tZHONluiZ4fM0bSWQmxCzcByG/g/mbF9gcJvcF/JLFuivrXOJkrUuaKfhDk5D
2y6cO87oCyX2dNKpwiqBgre3ZXDsSgzo8e7MCVOtjUMjHMIJLdHN6rPVM+qlQl54
dxvO+5n5iXXk8z7sqDjYmkkUF2cLKYyE23+jvSKeaiWx68DUarpz6yF2VFG3+ZHe
SednYqRH8HPx9Q+hw03CBqYBKnAcAX92vc91ADpShS5TldaO55DGjtYkze+zAj1U
lgXskG0hJF7cBcwZ0bC3YY4SNvwgWuL9Z+5g0ZyOp3pAD+Z6QcMKHkw5TTOJwBSj
MJCydqIbvLeQH7Vprfxj4hpmwbH10gHMxzEHkWrxHRmUAdjAiEr63OzvV+NyIbUK
JpwQhXczEsofhLQyQF1PLg+nX/kZhf9QWUjCGqtOtPv5amdyi5lpvf0dbkDTk6UM
PWy/bzLEfbDipFYa845Qk+9qtDVzhc2iQF3y4JcP8/gRUHnCt8Kk2545IDizM3fH
9RtzZbcS2ZYRkvOlFJfSGXfeq1MQzbxUvEFQA2lX7RYUh2yQlrr8X2bbrovCE8GZ
zLkj5SKciHIOr4dho1+3S2rPLQz0S5GMescSDZNQ12G4pTMlgbtk1h9/VOoz7/2I
IcCucypSS1f+mD8QUVixV9eHS7AUwABOyeStj77NF4VawYDt50XAwVRv9Au3lbrp
kn3XhCXeNNgL9IOHiii96NrsDIFmVq18XNaaNL5wN3tDHMX3b24R06HH4EkLdYIy
uf/+S257kncN3QGmXOxQ37yFUSxEnZxAgBpp5Wpe5NNtV8LyxZiG6upTBkTrxQm4
j9N1mVk9FPvLBoZ/huVeRRCxlpNXZhdJ9vaZjXQfuKJM28zXGst8W/u/KQCWGTIK
f1vL1WH+651rDMCF6frr0FbF/op9XvQC9/UV4JMZIoJxLyOFZJrac9iEW7FlrCq6
3dhGIChtHufnmxagAysM2bz5DZbI6y3aSILOE142OdI71DVYtuQUEgvfrOm+hf6D
IZ1MmWmS+f7rbDmArAkytFdcEMBoJvDSGoJ1kfvdv0VBUN5BzCF9rpoj6t+1vNve
5eFtXBWnw5sDLtZFy0ULCSN2OTM70J+HEADNNLu7tU4fxp82jB7R87Nn27C/IdzO
PVdW+V6s1vlxWo68J6Oz1sQ2DdhE8JO+g0RcoI8JmLjdUD6eEmY+J7LsBA92qwH/
03k8u3smh0qpYt555F2vPWU7zSbpwW3b0ivAPR3wXxdjYi2g2U9h1jSIMKd0EIqF
+73c5zii0h8+cS83cNeOzMaiP8lxs3qVjFkoyTNyjutLz8WIok/wJydiIsyWIodF
gI5Zikv4uQz91GjFuca99CCrlGRiv7Fm9rjmLXwf7BAnYXecolOvA5kHZ2a/x3SI
XEUg5Gm3KQzNIQMpMy8NqDdGpYlaFdgC5cK0P0+C4+hxDcSoeAfrsxOK2nKnOwX7
5aFgeYqGQJkzJVtPEj5PWFhQ2zNv5pXV+dx601lcFAQHtVfwF70803ByaKg2EpwN
FSkYG2lDlPWEi46oplf80Mv5n2aayNlOBJfwc/0FWMvS3RaTK/HeCM+kg2g56lfr
AiQ11XThyGZDxoRqsH2ntrnC+GsSLEi/hsa4VHRBQj2NmNvOMkNbY80QBZkzg3Bq
gjPg1wPdrR3cpQKtZWCsoK+7ZPW7xsRMoQvp6jv4WC785Oo6qPj9x9ImFetav7X5
A4tBYrfzqBDEk2DZ7b8/SmO398yNdShexJFxcqrgllQH4uOkyO6DDC6PI03C3V0q
pg4Smej7oKC6LziCCQqwFftlBlpv/QLX9m2BElKGioXCKW3biWRq6mrGoGOBpviV
3fq3fo9UpaGZUzjK6BrTyzhnb44S66wL1fbowpcZubKw2Ddflaz8a2YxHKKLxmfX
jNmyyovrt/tR+ho0hlIpn5AIZs4GlaqFzvvColinJtgO5Q7V/uUzOIAKKbzeYE/6
Nr9jSTt6MWqgQ5RGRjQdn90TZhxQfzzYJqcEPPAHAqK8Xk5kRo3b7PcEP20VtwH+
9174+1bf6v8Gk+eZVyc/65VEoIvuy/YjpKwo2Cx5owbE2xUYgvMCpVx3TrlMwT6R
THLMBnjUddXzkDsJbxD/hMhPwTBNzVXaNC5/4Yj3acXrJ8gr6uwnjZZyC6/8SDfc
umCRdHl4zVBF4iog8PlvdiuwH3v5Q/nwr1wsc8SdnHimFlFX4YM8q4BdteTteWyW
XTtFT9QRD4YSHRVow/IR6ZkboOREcj+WrE7L++fnjMesowUbyXR7NcrCycygjT42
Ws6FVp3bUQa8OmXyjsFc2M6aQYzgcJ0a1ZFzKjFfh6BvubBQIFiu+oHIKdH+7Cr/
aONRwJnRSBKhjabgmwLsHxU9CQbYZBlIL/55UPY7el5F/FZZmnSHz2KQTvvQiukZ
VoeSJjnrwe92Bb3wa2J9f5r4Ff6CMFLqk7A+ME8PFNOkgwItVFPuwKAMg8KpYvDF
`protect END_PROTECTED
