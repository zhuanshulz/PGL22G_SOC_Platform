`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGdKqEbHxoJNSWDPirifF0JSHKs0ZcNz+l6h1AA01Z4ZMKu3uM3JbZ6t/w9yvyyL
FoVP6KQ0uK/PmJHlDz1SyKai5NEFOilX7fJEKKs/Pr5+3iqZoTGWgJnfVfc/h7iE
8WOxTcq6uDukG7ehgU+xbRz3vrQ8HcDwHFQSnqa2yYX4ePNuM24VeFMJcXTbUJcP
3THRZf6icZ34cZbBhIDGBNZHhBdxvh/Jxhr9sjI/Lug8IPJ5PsddhqcYF/iY8+MH
8jHrQuqik/3XKRAsdTYgWAPSQues5bUGBNu1/khbZXuDVhnQVeBvrjpmjaHewSue
1/6fMXKtCFREV+3jAH6RDIYuLHN5Op4D1b+2YYqtH8j9T59plYrowwUz7ktOgSPY
cJ+mQbH5ONCmkP06S7JCNaPeJlVxFjecNvqoT4qHuWQP91pevhJbhxaWroCHmWyR
KUjCryTJIBL+bv9mZI70IN9w+yJ9tMJ8lf4oAO1EGtR3VPxqi0M1WqjrRBD3uLoe
tu1chuz5QyhlEEX5g5qfTuJxHiXl6yGbP6mlGsTmNBLlAMDC8dezjvB1qdufRSeR
v62xwOnY6M+vc4fWap9gN5jSwNvRpgAGYB2wdwLQwp4HhearQySr+4/ZJjpfbTdy
ok/h7G50FPRbZGCHvWOesBbOXCfFtWHnVCTQAcuTBj7BOMRaUEAoLg1fi0oZvTKN
gvCYfCw+ppl7q1USfIj94uCll+K8D8TOsUH5L1CBaUXFDeXifIYc5fiDtQI13wIO
O4u+NNfyrug1mFKlbH4v1kFxXKrJwLZiAUf1PGaccn09N4nPvgTgThjBJ6lSx3z5
dflpN/TtUEnUvyIHjpLwEOBzLRwT4gstb5tZJiiQwVdS15woa8DEfxXePeSI5u3u
8dsK30glzvCCTS3+eVjKZtkK5l0buSobPPswV0T+GBtNpVvcT/etUIj/HhknZUp7
HXgZMihrvOCPFyTNcwP/fap0OdWB8bytN+Mazs9xgoP/ZE/3ntY1desYyJucGqPP
i3y0vOO/NFiJkZaY/KWeH//XwhHiEkjfGkSwd9VQCCAkJ078T2gnoc1zQj11DNP+
3mS6rP1ic5ecZ+WWXQj+4nZ+z5YgjSQEgLOWZzvRcT9CAy77OONHFIvv5ORw+4YQ
pResdicht32sFzyx2U1cYjn+cXfnjZ+hfJIWzNgo4xqaz5qTYA/NlNlkIt/Oifpc
fvNFpitHL43Hr/06hN0wAtpHLKoAO7Mo1aZcHbNe4UBG8rVlCmiaSHhxpeiwb4Nv
LzydneRVMuUsn+mzP3Jdz+VX0l0QfEfC+Nf2BTmbCSAwuY9rP1C+hW14E3XuXKQK
O0DnL5LjvqvAUWSzC1fMvYy2h2Kt/BG86nu/ZQHba3CS0u1aYl5BfQ7Vbc5mXXBM
oBT5S0tp2+idZjOIB1MHbey49TFJ+bBeE34F3EYrHkjW7g9A1YA1wPjNa+YEmN+n
7NbN9TpO9boUgP/HzX8HY7rhocss4zYfmzscpIpZ5ZYpFCxEkXFTUxaNzQ4Xpdwm
z0FQ0g2RvdGMe6Wf5RtKX2QIz4qK2h/tosfWfHdDNFqRCLE88Ly487cEoYvNXz/f
qFpOYl9StynagBzrON7dUrjLGYBRS2rqHRfsbiYsuG6upQuapALluaNLrozz+Iv7
yyjpOLs3j/nQE9FdXq/0uD/loKV4n9s0kr2//nkK+ii7SdPcv2Sc7e+qhg/iwNuv
mJ3Vbkl+vWW4t2BQjw6Lf3P5u9gXaFRIVe+gMIL1A4IjPplnsMg8Bb/+Tyfr5/uH
uN2Wd1xbfNEK6+tEbsA+XgxaaPZ3ICzjetSmDqriebMnLob7+EwNwtX5f2dxDW2f
gaMIjC8r/FbsRiPPxuAF/rdKK/EoJ3P6OjqY8/N3KX/41CKSBHbRcYWV+sNYx9nr
hSUxt/hYYEENy14963RrkEeD3im/riZz06FbFbdTBLw=
`protect END_PROTECTED
