`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dge9HlZGiHc3FxouQvalkOCBD0va3vvAL6BK0ZHuHG2pLGGZ3y7/zh/jrC6DSG7d
n6aWJZi8h0vOQC99iZBNkfTTWortC1cVv9CUUxA7UpKdb5Hcz1VvyopoOA4Z2kr3
T166+fyDBoBfWIj5aeG7iuGSxVKrkk5RWsuzrJVuo+0Q95Xw9zoxt3KgFzYRhkp0
WcHTnEGoNbz6CTeHpReuLSBLKLsvTfowMCak1lmP2F5Br4gnDMTiBw3RRyjw1l4h
Y6rNbX0JWJGS+0u79U5dD314M617RPWrrHTR0sF3dFaur5ekmlcZJtAtOsh2kF5r
941Wm3Ev+5YLASLWjtLQ91hL/Ua8ngtsZION0ZNnpme/mxnqmC/38/KizHCLedIA
c1YAL7IWMDZ5iyvjymk1be+c5R8nB3fX6JDDaSfs8tG9IZRMJTbD/7lD3KT/Y8wq
Q9CQTOTu8uN703gkrS2/VhTgYxz1GvFVOeGaqOsq1FdL6yhafz1wO8Y9SIBLBSRv
Jbg8y/5R5MgXMApGy7cWhiD6dHiqUFLmWqtwPq8jbrSwK7z2HRnuBAHwlBCd1CW/
2rJswcVKC3AN1Gb6k9Bo7a+LplXnXj2Y6W5KTCWH/CnQ+ATHZFmkWBt/9w+W02BS
VR9FLFPYScxCtMlAdsWAwj9nmBV3muTpW9smX2pbbuDnWTkS+N8jzTLLlGIn/hhU
9xaphDJrQrZ1yW8fuocNXZ/fe5K1LPWXi49Jf48cLppkDYvovHS/0GPyjm/DCvN7
eXRviKT5P5/dx7gyUOnm8m+U43rjTRuDWPAKENu8itK1tIpSyWwKfqC78Wz57YqN
RPugfmda0OOl83XgvPIA8ZwV0dluRoZZUutJPMI/t8xZmUqG0ZvMEbMCqTsPzR6J
fxThPFgjzjo1+hBy2q+sxoO+AmCrcV02JPXyX2dwqIA249ZQpVfiEfK59t9ocMFs
u5dQKgQ7hHueAA2IVqHh5Lagw1kc4jBcJ5JEyr/NH3qiG2Ya4wBkyQhgSB6juVyf
JGd/s8Lfj0Qm5FWdoMxx1fixHCxlNJ53BlXb6vitLcscLeAtGbPJWUt8teTbNVyd
CPccPbnXnB4GIkySwdMJlxKU4Usj0MvAJW5eDCzBxO8y68U1QUEZId3rDI8y6Vxi
N8c93yylh3RlT7reICqtmBxt4YsGj5r33sk6/gIf331AogxbzWa07gJ5cPMg2GKI
t0bLYyKYN+j03qcX+5a0Nw84h2PPYBkPrHRfwN2iFE76bmSguVTBO6F9ttgYHoPy
SeY7Jqrea0H/3frQbQUdeBBxyk+Gbf3UnrDLYVEVGE2MqU2WnjneLIxnu30EkKOC
5Z5QuxOXWuOlbuudXMcu3GUerqAsk5LMFQwdB4LdHWMaKpUBeqKq7gNlvUANgGAl
DyL1CBVEwUQcOWVym6WQ5QCRlYCCbyfoLjTg0px6gM+pWg0TexL4sucgLiXpHXTy
8LuyD040zWMKGRLWKVVBknpi1wgxkRQgCmsY65A4/Gx/8d2O6iS9ULT9xwpjRPOR
6x/zjJaYpEGfpbMbCyHxTfPLElkx2jfWQqlS0VVKL4LOIfE/VWSlw135tWOVC+nq
+dY2CZsH5imvaBCYGcwCL8OtFO0RBrOEJWT93TJ725tLO/8yYxPVf9F0Zo+h9pS1
`protect END_PROTECTED
