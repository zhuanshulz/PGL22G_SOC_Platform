`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z+pGww9a6e1nFFMnzL8TqDLsfo0jIAK9mguXGjN3O7lFH9pY9QKu92FpnI7oD8mK
GKXGnh8xLAKQ0yAJoyo/HBL9A8pYLXaVupu/72dF5o2Ao6nehV7tr51+qWm+NUCk
SU53h/prqETBKG2XuhdA5VfDJmjwFbo7VL9eR02L6Wq3EkRrhleDkDCoTsxXtnyL
zTWiMimncGnc9FI/4JPJnW0z0UzK6xVLnu6bUANfQBLFxV3Qteby1uQUL+ByVUuu
jctWO0OIRJWWZCbUNcG1jhP1sdzt2QInarZSi5v215TvXPNZypleqtPsrg0m4hlB
UHoCuxfTry3gTAabY45ZZ7md/Khgl4xeVJhTIWZLclncAZ+lQGrRXWLosrO5xjF0
ZdR5ZmVTcQkAHxOYy6xc3XRuRB9Itid0sM1IqzjNhcDXfMRI5FMXuMCU3Sl9P4/O
oMIL2fI6BM1JAEZ9X13qL2ZN2GCoyAot6V9K3v7PJD9WTcsTTnTjaWP/7qJnP1Kp
vSHkws3DU6Bo7ZVuULbTNpBnVPQI8XMFity2wdPSlWnj6GqdzSHgNidJK0eJxEmT
BCZQr0ZX80DEDbRI8mBI6mr7e8gN6GvJOCf5sEYgZDdWT79faf2tO8mSXqvzWORw
DtQ8LU/Jjf4+YLodxQTKtFAza4x57vveEOpxXNk+wUk=
`protect END_PROTECTED
