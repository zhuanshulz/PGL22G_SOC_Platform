`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kSxkhz0r/j4fKaxi2Z8MyGQ5Di3caV4DxlU25bY6o9TWJzTPtYsmrjt0N57kV6VP
KHTq4s8Li3a4fOLxe+c7Epp/jTaASpws6ho2R8pvyh4xNmpYiBGWRtkEfvKhGCLC
9hvt0KEbXMfHKAYdXRHbujiVfLpr0mppgdnDSUSM/UUmJ3RzRO1KedQnK3aNtaIc
GcY46Ey3sx2RtqWShsGwLPuia63QC3WH/6ghtElQ4YIa3mOcFNElZHE1B9xBt5k9
IiSchWrP4ZTHhItEX6/6686xbzPWLW3Srec1fWgMw1TFr1Kh3IcQt3VFaAXFkBlR
zX8McwWe9PZn3a5UAlSyl6DyT1t1pOpueHWWqzi97oNG0zVg7o+SVzaOT7aN7siU
yLPPt6unoF1QiIPu/ZP2NG6/LB6zRM9YpwMTHC6BgvF5oPpBSixZSmkGhMGCdjCM
TAZSCVhqC1NbX5urn2V/gvwrhHmHdpdGbGoTsXIWUWEkdXWK5hq9C2RPTId/ITBQ
rxRzLn9R7xEh5KjiEnn21TqdpxRzDzRXr3LTdpmALH8BwFTzOnruL1K/gGItdSzz
mlTcaDETDg1C5pZzLTvZYTgT68rE/LZZpB2CVCA7UmerzZRA2Zci85yyTs2k1lWZ
CAyRkd7bAiOFP4zE/g3Pt1fJL+l5PwmRr5NKUVbh3POiwitVcHLGuWMMCykxFHpi
bdlnmKIfD9FGLFd9MeSivQivM1Au1eEi3oKxWaRj8LhFKE0JOrBuB7L0OWjMvxEc
OucuDFtQz8OvePLywgWG1j/oQv4ElNpEzbfqQrFZ9rst93oGsCYLyI89oYob4kVT
d5xG929jHq3c+iFAos49LRqpy+39BMA6TLSfPf0PRyo=
`protect END_PROTECTED
