`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
au67UmkjiWJ6MStCQgpcuv8rTEjUWyhlotlOvbXeeeQyv0ostzrbXxTm9JBNfSKK
AB4izN64akTuMBZz4Tss4pruL5eJamHumrGNYoTxZ5LGgiVQss+ECtO9mLC/PgOK
rmWdejt8VaLMvPxAkmtdURIknAVEERLeE5gy3qBMIDcd8qe5ISCtjkYAxL1LRYc3
UfdL+v2zf9sd5d9S20C/8HHKCN+z3jhUK8YnnSvX83VR4BQ7IM98a+7SjpqQqo/m
5bUV+3fp+xhFy/13sXE1QeVVtWX19C+Ohn7eW5iH0vofELY8Oxpga6CpFd/R+cHV
KAy5ayjVM+gAJMO/YMhh4r3rnMRRT7tDdJGC4oqJv9wRrHMkzRMEupyJqjsK/B0r
1HGL3L3jPEYs8DrEIVnOncMzImlkXQ/fZlRKc2QlcWrYgregLh4eweZe0nNJ7kEh
yQhf0QBGl5TiErpWuP4Sx60/KK6Gnz/VrBnA4uPbASe13NIC4nCs+AiSBxc0f1nt
OA9iLPbDrvTjOdjCFJKXZZnrfrydNd84DYpdgjwiIasv91TxxkHHaCZNhrV17CHW
e1Ttvrm65MkIw41UqP6J5d1+OqvuWmlZK/nHNhUbimYaLxCw1Aq+TTAHE2G7XRmw
vvrISgdFGnOGWmpZyNVK3w5CikRO3Uw4EsrTvZEOJwNJ8FVzRMKzx6PaFriTKo9n
rHPGwDuAdy22FFTNjwBTf+fW+ujCBEz1TaY/1aom8m3hOFWxSuXpoonEHTSxdj+Q
88ocMFCpv8wW5U9UGbt0kRIGO9e6U+W9MEUT7eTEDVEl7Kz3lkLO9QS3qMNanAxI
/RyHboevhZmgBu/srX46CPTz8CsDdM/gAfrJqB9UuBDb+mmj4R5iGGJ5HDtaDCej
7qa35a9vJKONl5xYWeSL1P8NQTUw3r7LU1SVXX3ypTF+cHfSAkWebvWFSk4W1nFR
EXVOgrOMaqeZaC7X2Ofbk2BmiW1NIz2J681NLVhTrvOKIFYQPUzkCNK5cHW/FhJb
AFRsCAM/T67cmik9I3IBRUYxNhFX2QI6IRGJO1UiWKfov1XmlqeLL+RDivNbt76t
uNPXHr3+Uw/suxyGVcexefGJ4HbGP79fpjpVSoEVQAgkiCvJ+sXQWxEB+NWEz+O3
Y6xPSOAyhA3hPBngydquxqgpjUtdGaUxi3JZZHv0szUl/3ZECCz3ycDS4U8ncUjd
KanvnzX5yF4hINBkW7W9UL1kADmgeoVGkNR1l4FfK7jKzV7dcUj9WEP1KIE6DorC
zAnlQg/LNBTQDmW0iZnTHEB7ItZbaApZRMFb0UOwFn8aRI9lKcSHCx6AZGLBXXtk
ngCqx8RzJZJUMOUCi8ZRzWzG8uaIbPwkb+3W5DmKh6q90DH7ESWv1SiLOWTvW+q5
Q7j7QBo7YD4tdpk8z7nrbIoxFIgKM1OrvmW8/FHDR7nLQYJ5S32y10F0Vg1Bn6PM
Icvok4Jf4YEK0KkIIPnIGAqB2bLKey87mXtdSZ4z1Yr1tcMWd1ir3chqRTaXZGr3
l1kitnnXNes6X3KhkUHMhi8ADhuFDwkTTewyVJrsMF+ZjBvT65Bd2ssCQQ+/S0nF
2seOyTrgrKOZMIUmhdpi70O9LldsAaT0fI9IdSY/qMxD04bKx7eD6ABfh2rKe4jX
OsK5xHI14T/vTkvZJc3Dfi2urR6Jl68LqUD2heIx4YkUwJQvqNhnYAZT6oQkhwf0
7ZDOLe5oSuYctqQeN4HazmcBxCwknlajWdOlIUs9iHnp5I7SeJqfdZMx3KYgwdcp
Zz7tg1SQdG6T7EQhAivhGXTBVlSxG+BCmC4zL+cbpCVrN83A5ElDPOdyV+gr++fF
fIvdbp7lnPFp0aCsQvU++IBzU+qKoCrs4vZYTJrpMrildZf+I1pId7BjpGMRV4CZ
LrXXpNDpDgoNJEkpw06Uoq/bbHgJc0scHWyDq7b8AN2+36YGYeTWpqh/LMy5xmkd
WcVxjI9+gvtwwYpJR7ZQRD8lb+2hvi5ED20h60RVI8KiF8KAziougAkdcPqCmvnP
Ve8P6fWhJlbCql/9nCy5KukaiylZ2lZHxD5DCWpPVBOAOE6AbQjLXtdyaJvSmtSR
frzcepMQ3ZSar6/+EbueFnr3unEhUa8ZretVE9PvlsY/bV2iY9kAqJk1SMryyr8G
zY8nRfZS94+wf3acjyrwtQecrBZQwU+OT3a3GvlA6tYh85P81Kmkx7R1yM3rWiR1
OecRaKOXaK0x9mhW6YPSIKPC9ca1L66engcaFF+evdRUAPQdU2HQb40mqKJYJd3u
paYNDq+O1PV9cKOX6zoCguw2Kyock31QomP8LiEXCJBeiV15L80lQOQdG3K638xf
LuiYJDtTqwIH9hbrYfoenam2HlurHg6Ujj+kHTuSRvlf9k2WqguAUWlbU4E+SxEa
Sphw8BqYOHUxDw0g9O0CRKocfGqweXDGu7BGOYwF7kYWoyvhpACywYCdssi4GDVj
uktqZXXUbTJjic4FFAtMBru6aDGvWmogqz2s/92FxXZdvUSw9uMnd8VaCn70thJn
+Lwoq1QEoFKVYT+ESqKSXXXMYtQeg7+U0XuGpZ159dR5uVdgiRf6zFG+adlOQ586
ZGoP7GxvFoY1VvuQOjiajGsLh5WCDEL6UGasC2bznKmmFobWhbHtg8TMEbDe0rp5
T/ejxv5ZajXeSx6XtnB7oQJRoMTpFWS/ibWVxP9gn6zV65rvHjr1KtT3uPFz41BX
F5Hfxop4GbT4Da+JqcFu242L9018c5/cP1cRAvnmswqwKmaH67rZbsNkMSzjwaXV
Gl/fe456NiLs5eAnbx+imZ2LAdQ1zGPuVorBIu1+EfUm2UQPujCBTC4tOIWirePQ
n7AkkLzELqXgVRJHKBccIG1SQaCdd8T3KMSQAyXHxfpfCXm+jXfNjwZqXS0i/cyQ
jmaAh1HxaalDHVIYbILNWHWMo3vHBrIqS8Wur/yuwO3WjubmKUyzUK+Q/krGItu1
+Lfq4/76SizXXJNiYUAmSyQ5W9c6OGaebGvxtBVy4g7+zynUoLhkgmRO0ZDnniq1
HUb16fuxrJdzOz2d1BUezg==
`protect END_PROTECTED
