`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8N9cXqbClab+Vus1Q0iaAss0R4nP95hn8d+u9wGJnjmyBRDLguKOGYbgpLgW0EU
V0xyy6Y4dOTRoYgQZ2qtHVK+gMFJZw8PNW6j0RLfvUOzFQA60ms5PFvxxoxNIoRX
/jUZqQgzvMg/1RYgaxo6yVxRIFgbQcV0/jlPeKmnBG7TIkWf+JLqTnzsaXNM/pow
Zodlr8EZL8iWLQH+sVbG0+j3rXN5pLd+9uc5S9k6w/5W3cQ7ThjyAsqALVMCUk7/
oCCLe6UKw3Zx4L7i5XR5iPOw+yNCIIPp+BXrjTIrVRMEGtMAlN5pNuCfoElbGJqj
MIbVN54CTe7ExhQIzLhRpFeG+vPmwMuMoly8KHlpkx24ypnARWfybgCq87SYPEIC
mbZx4b6p86SAvkLX+h+HoS8R96nqrT8GApJFcNd+1vo=
`protect END_PROTECTED
