`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HvJrOUm7eJf2GRWD1uLgBmwWA0Y0ldOJX9U8YM9Iga+7n275jvU/bszXyoL1bgwt
HFUSBLDyXmrTk5UB425BMvMSMLf6OnzdA6DmDts9QinpluvTGVF92dzdpaTk8+7H
ReADArGbviMhyshWKVcbn2WQj9nJrdQSLNggIzK1ZJpawztQB+zReqz6vudmudxR
qMbCUcYDua9DRu0sj7R21mNnc5ViKdDbjP6yzwaFbsS9TE6nXjnNOr5ZlvVGx3Kn
JgBHX7somvg48AsWCxtkvZ+6CM6m+BSrGzmCZ6QgZX7EzxaatWJ7gwnJoPuLvhZo
0U9b9egLtG6AY4vcOZvjQS7siNQzZGnZlf1fK2zUZ3iMgJnqKTrBptnfwTb7z9yH
pidMRQ502XUfF+XCon1/MApebPh+t+tbk6BPuesVu45778KzQjra4vcvTqj3YK/k
tSOWzL64JMqCAp46mJAcEqygziZKJFOhuMQ5CUenZBqpIrAglbUvRLj3GRR7Xvho
5KrF2CqToRtt6Zs52dCcJwPD6bZnWmoqTTDb7A/8hhxpEEFZaoRCdCOUfgQVO4zf
Zw5FPZ8JkcahgZwP8PrJzdPIKw68Yp6NwnswSHfxe063maAsFiTVib0+vNJ41eQg
pK1r8rfWLG4BmbdPIwPkBKPQFw1D8Lz057nPrX3lDwKtKdrp2gTK0Cwkub0AV8Lq
L57Z5cko5Troc9eX/CyiRRJKmO49MWtRQ6NYIMtKPFoDXzJ1s3zBdmRswEs39sZZ
2ck8Sp0lEDFNWI7OCk2iB6pa1NsejuaLKSaeDoLi0we/W1o+V81jgmyjBT0zEcsf
muJeqfhzQvpRFquMCj+aNArhrpn8ZquOox/Th6uE77r3AlRZN0SEj6D/sdh/CXjI
gBIX0Kr0nb1vvfcxKII9YFoe+v1lXPFOUaIr/FWASbGyc5WxuIkam273Cvp2W/4v
Ggn7FQTPbJ2nSr01nGFAV8e3GDk8JYz5fUSTgywEXpkU3zlaF8qYU3HCIw/305o1
7Y+yuJecU24YbaEOY8awbeiK/VnQJroEqNbcFLD3ckOCYRhqjiXklZPxM3iCAFja
OkwRLsiP2M4/8QvU0bxPYHlcwU8iJwmM9ZMMfj/FncxIy2UGLnnNAhqR9XhqEj0d
0sXtU00p7Mi52C7euEwiVk0ybDMS7da0Ia1AYF3NfKuv9SFAzjufM0wSknIfklAj
`protect END_PROTECTED
