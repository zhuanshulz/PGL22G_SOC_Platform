`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WXkvdEvqM7ZMvUnIUjCQ8He7mEzA9CUrcJ6oA37XFl3wwTNH6gSbncq9KY9deFZJ
SPh8iw/9YlnqXxgYWVORg4tdZ/KKmo6BSGB4TLiCOHhJHVU890Pdw53DhMx9/EZr
wS2E58+o6sudtzzanQDInlcQBrbLOBdYVpGswNZfgWSQxqdFzhV2q8iMMmn3NImf
kpox6uHng+cb9Z6xF4Xqujra1H1jOalLfJFUVV1Fd9Jj0wmfT8FKXnH9NAJtE101
1/0YasUlQtqlDQuaGKIaFftuuAjvUK7pr5LQhInLFvwAYBxF5JDRFM28dhs9vrLD
nvRLcjW2yK3MMxEkhdSkl5ALmRV2AOt5dhRdk6YpNKuEXuShNZzEIcLN7S4zpWss
EUG9ycn7oeicwmqHLe8JJFSrzHV1JOSXeGXR6bNFvu3uGlQMfr/ko5kXX4KqFpaW
WZYAjHtjtpkKMKCtWw2Q06Fwl+cVcbi70yZoPISEtEAGZtQX6JGEdhrs13ZxHS99
NJ/EnnjJpWpl+ZlfLcvwp6fWXSePZ1q8u2tA3w+VZJlJqZSuWjHfqFE5EeV+dMuy
zvtoWr0430mYE1mZrXOxiCMFyoyvMECySUVjIMQWqLAAzE+JDNlessv5A4GuwIID
KDzXNXuDY15vaArCunqWBmrmI/QNBbhMptIT9obgGjChY2kaLtIUhAJa+m5IqhR/
Suf0qw3xsq+zXx1nxqah5Xerdt+0KgJXYwdmUDd7OTDbAthYz+d77as3Jc74eeXI
n40i6ePbzudoFrUab3B3C/RRmonjVj0YLv7u1yrZWXg8EMpSYQ2q0xYTPhh2ftyt
1Lpv8IUeMBk0PtcE9Ijo7pa1bz60hMIhvcLgbq+Kw4tQvmSgr2kksOhQa8DKXITs
P3nxPHtvCvhIyymvCO0ra/EZMF+6ltUT6T+tO8RTFSE9LRCl81VC6zAs0WqmQfdK
nlum9/XxXYQf39jRmqFcKMyPJ4ko6FMOvEZtUTPAHUUMVJ29rkwbegN9DfrONWBO
zk9SKym3/7jPTaqIaJKvBZy0US8rcgjBZBhgsYxCTYoHwiUjf6VewX5Gse2TELvZ
kAWTVDTXeYqGrTlsGG5zosqq2A8mZOIMiySWfTGRATZgihkOLvYOuQfsQCuymScz
2S1Aj1NZKGLVuQpYqveHOi9rxF5TbdOxfYufepB4bSTrxRcPUBctOfodKVQK33aa
C/y4ooP/H43h54ydAVWvK6KW0nFcgxLyfpGNZhEarRcwz+VKTEtGKrUZEVyHKs4H
4Eb0208Dr8QIeTctOmZF1K9AJmQUQN2kuoJ/d6OpSMxXQB4nAOG7Dwt/d7T87V8A
4aOOBCGWafrKt1fzauGKO8oqQutNav0uWChyfbq+ofuKnF4p15dKGvxhUmGpxrm0
KOzJnrdT4At8uMPMRa8rqT4hEUQrmS6PNjU+ZJoK8A6EEdL5R+/9LYVpIMMhxeJB
Qmv/3AefVaVtt/ANUNqVETKCuHAXhUPZ36lDWhTEuTzjyC4V/WxblAevnsU6gNaz
PGR+TXfrjsgY3e5Jhrk63m7MhI9UwWPT8V77TfuUQyazH2gW7DKqlOXKi0L2gYrZ
/5cWAl5sETtloBQI3P9G8t5DLw8wCrDTr2s3x1nk+G9JfuzLiZGmBcpLce7lyx82
KkeXKQOfKdStBq0jtukcslzOvoCtvbVVWSoCtkYA5CK8raC/p/0ew36yG/AWb2CR
HTT9Yl9cA5W0xG/cbpEX2+OEG4x6q+hjuzFwBw+rphSnD9T+fEipeT/MZdgUzTB3
LWX2hnzeKWTWa8d69QQVD/OS32NPDPpef8f4NnsN72A7WhkX/VYRRWCY4LXG9RqB
ccGANavWZITd7cNTVNKhFG05WOSkjmHESwskLgkjem7uB1mM1Tb9jwcvbDkpI95X
eDNwy7X5qPZjCai45ubQAyw9ilJCFd8PQzMqH3uoWXyaQBTzy7qlgLZ5xwEjncTx
QXLyvg76+ACZAjwe1Sub+tiU7cx3l7gpu5ky163CWqTjJXKhjgoVUW1F90qSa47o
tKJ7BknpYrCFNrGG5yKlhq2nsy3Mtxw3GYoVhP4nezWfGKWFx6l8fFsLJLlIFS8q
KNwsb7n6Lh4kbrLzZglIGoD/k6vhCmeX+yLHaFQ7HTphEDwZykaexzgTKASaTMe/
j7jGjENKfe3LGyA780eBV5NIfGYWzDJENwN1XNdD634rIA8OA0K/ioNk7UG2o9cL
2z9JJvAfYR2t75wrBAZOdc8pZ/1ksczG2J6R1HWTIKPgbv372lB08AQ3T4EkH1oZ
Eu0UiHlt+iUcTzCkzHdaZiEARQJwfuD6B9cLMmzHf6gEmGUbERVtwYekUx6U1oFA
Pq9rFYwbtUrDCjoNliQAFT38T0OmYaSfzCHtCQcJK+cw34Ql3BLDvgnqWIrva0Ed
1CeXUgt4m2GSLKDkR7SA7QEe5cCMhxm+sTWoIkgOq0xmnNxzllDxjiFJ4n9mdaHU
zgNlxOyxo7MITPA40VZR5MHSSM1PzZwBZmx5JRQmCL2fXBr1GRgNv+jiW6kAQ5yE
ZApsN4l3i4QRE7q5RERlVhZT3I3tuFxiftdBs8WklkOXKmNFharXjcXY05LwQ1Ja
M05oyCUk3yxcp/GyBtoXkoKj8yopfoBb0ALPIcJ//+5nqmDNFFBBADVXkf5po0pL
rcXiGV9fc7Xdmia2qFtV/a8yj/NNBZCcYCGqB7TkU1H5Ulgfa8W7zedklwNrEgsQ
b2OemfKFNKtrKq+IXThhGpgtNlJiIfvGZcu0oOQUv+euxl3JS8AN1Pntl4nuAicR
ESdN1u/zVE69Ke51lFmarvmHx+v0TNomemCjHsiA42E0GalyrsWmrgMMBtcdtMrF
tW7htPekmM/NcKYAfZLxGx0urPw3hO30tn3IOjlSzteZ0QmksZKBEYpwtP+q2q0O
EW8N1mic+E5aIMTWh6GCWP2Ci3Q0kH2I06yB16HRJw9F23sthojHRrx/dDBOie5i
dpvbTw007m5nRo/UHuEF5H3YnkPoDB8l46Kycj8TxuZrJXbG7gn32P7ZAx0qb5I8
j0wrjrEzJfu/OJbuyYBNe3V7g+clabcrj+VZ1OeeZH+GyPMeRhOvLtXxi4kt027j
npdEavbALLdVV1RFKz1jRihotgEBU4pTGg5+G3XAiitGK1DezC/mAPp3vfMYBt6b
7rUlYnCOiNkFeyJNXXCJJjJtPRV/QJIsqDtuKToaJQXuE0ZXPlZmV+51b5KxWEEt
WtXfLAYnzUnXA6/qPJAF7ysoWQuJxTY+qo+Q70GUk16Sit5KuJ0hufrKu1NpJ78V
AuPinT2JNdUQPfXEBnYeMYRc9UxoYc2Dl9z+UKVtxNFdMzMuDrDvDjjk/A3HMS9g
q0prYG1AWu/5nq1Z6VsMdvWfFLXlvfD2Seo235S0t3r5ZeFbnVJKngLQr8KMH2tQ
PkM+aUoWYw22NboKHS+v+yVuis+itT7uELxL8dl6bJUwnjyKspzW0Gc7h4SqwCbn
n+vG3MrshQzLWl7yODlxLbi1WvMXBIrRt4MPl0U5+LmLqb0J+iThmnVb0wTzKmpx
2rqScSfJKaRiRkTjZ3ZYdlqvQ/lBPuZtiBJh5F2g3TW2FRhN18UsONLjv83XLv7Z
v5rSPR4qvYWilEf/rCpr98Cbkx2rCxjhcKtTLrzdb8qbt7SWD0cTxi4t/FJBnecO
hdEMFpqn5nAgFouLe6ocYUVBmBM6zj5elKVAvIbUC/igzRtS9S5x9T1AXDhHSz6i
XPwp4GCoyPaDYTuvdNxC2C09hBs9XD7ara3fymHCRgb3KvHG+niiH+g9FBL3Mq8L
PjSvXojqUAajbmwO2kbSpRowa9e5tPwcGDy9MzSxtTuC2UZKea5TroihfbXy4ldK
HiXdtpWbHfk+5ZLDXSfKuzMV9fUppcy9Sf+NQ5+GQzg5/HWRfy5RbuhKiTwNGpNx
6RJQMUmIR8f/LNZqQzzDc7p0FKvXf/+M4Vx9d3iUwnsmlqKDC6pkQApU0LGiUSeb
7M72yppRQhW7WhQBqlelABn2hE7aNHXt4uSGTLMKrndT7dYI/IRMhQJDSCWl3RjW
PLPNMd0zAolMnfHQqMDuSe6RIOqF67RLldD4Dk81CkGMhQXKUnkdhM5VLzwgOmpk
bf/EQRabCWxRLels5NyNTDdtvSlcGMf1EgQQ3rzS4hlTAsPv8s5Uz+o68fr2wXU9
U9rNjFpJfBj5LJc0HrOrirvndosnu9nXsRCkAKK6pf6XCTYZs2VHjN1JHGL5CXG6
OzDr23kXiT/jnaIZMc3Aedb6Evncn6/XiqVjCldX/x5X2Qey1hhlHLjgLyYrr9rl
jzjITzw7rWpVybAYk4GPnalllyGFGt8t3n4dVzKixHE3GCFHbxk1CACNikJEOUCW
Q7tt5E/kRyoEUTU/rMEYp63jTHRk3iL+LuKhgQ9Xq5uQAyFVann7fV+33GKWFszW
48oOFq6AUGnl4M2je4SbChmzGcrMb7T9ccCunhmCDbuH1wTH9d2ZZzlhFwK4FZnD
z83SocC+/7rM7SnGs9H7gZr844tG19aQKH9T7Dh88FMnxqXKhqaSNev1KbVZdrlw
5Az1X+Z7Nc6MmrO8qrOJ9icIniBqLUCuDyGKS3zHI2qv2IaWdc359DUbl1tiENwA
qxXU1eeFVd89svhoTonrCzcvc/tYOBwJl7Aa0oPCanvCy7pKxkzfG5bgjg1txd8I
Xn53DaanWGyS+ZS7lDLu+uLnVTzdHhFrpZeKzvjATGe2pbqHS/mf4GP1jdafNQjn
7GFP8kCNPL4CwonJFzEhScL1QqIhA+X9F5LrG34CEj6DZFPCtR0FxR9jvc5IXoJD
Uq3e6/vAqu8qhax0WjSDVc1DJMlZIL/+EJSW4NF62AoJ8TA7JUJLj4tDDS/SRLx6
0ovdeRN+u33X8N3C589ixQ/H1d9DnJKUh4Ll3rM4Woc08h18SCrBUW8t3rBbuXvc
nCcmMa9Wnzevs9dVqL8RrxDOQJRPy5Wn3skBsp1TW3vfczu3Me2AgpbNHZaR4uID
IeE4w29VH3kA78uYaOz9vGGDQdzxaaqMn606OflHIbKUxrncmrIAYwWOmrLuVzgS
rMcDhPURL1vn9Xk9ZdMVW9fyGZW7HkoF/Yk8V/8W1u0M0OII+URbsnqL7J7eCqFO
I4BvydHShc7puv9/t7DetMAnZhIBP0RNQzx2SoQ//eveEWj1DzMbbRsieO++jVc3
Iokh6R0YpXWjt1R0w79WTwLHD4odu8smlnW8r8g8GApfIYVsSIF1MDRo9VUQwMLp
AbP2FkckNqz6rji7gtXD7zikFhGvSi4+Kn7D+kFmxCguDE8Vy4GgnEKr+vQKxO0g
+DfqahIqJ4e7ARgZ0O8oQKlSdMGPWgSCBr857xK4r/aZh8pgUBr14sBaym1zkqsx
iZ6nrQbVQc9K+q+XqO4GH2j1rKmbuUnPq6Add5pgv+M1QZoakHGGDn8UGrhTQXQA
K9n7OAkqH3ju/XMlbbhRn69eo0B5JsSW1lLhiCwMWGzLhU0paE09rR+wFWKbXlDC
+IZvBacnwXXSjl7KEEZX+OVXyb5P6iXJdB44qcLTv+Yp3htnFY+G29JCr/CjNFHG
ffN2+pL0pkDoHsB/js9801yCYqNZnHMzJ5oG9ZrW0qA10oVLSjVAWJC3nKYNdF3w
3VeTL4l/XrsQqLns0YUdaZjY//M4EeY2hSnJKPo8u+z43c7qZte4hMa+BYmj3Zf0
H21CNTlcZUvUVbJHOm9AkSd9PgB6A7u80pYXYaB65XLoq+zU4WmKYYNGx2QNqMTe
doyPbrA0hH1LkRWcq97Gk7ePuM11M4XRZNM5bfOX+XIcZgTLDreXPPINncZ21bea
5uPUU5IFK8LndQUgsVJ+IZtrcLwVB89z/+e7fGMr8rZrHpyVd8KnCmfwnWuh/pJ3
/LwTL3/ZChpRKXlWYCdLM+YnPw0KM/avI3bOq94IH3zkyVu345eyg5KK6Ln7+AOy
vVzQRiNFVtMjsA/cOCDJbrw2m8Oip/kL0eBhyKeqnpxFgLIni2jRseznQSA+Ebi2
TFR5lhMFlb6Zg7o13s1DcvKShveUxV/A+EQA9yxPAf5cgScOl7pUVTBSPSoCZ4St
QP6tQpOuICBl2bVnGxRwUyogEy0zi4TVwHJFvoGqsDa42/hqKCayGz8vpXkVytAu
c+THk6JcKlr3asdn4WF/00mOLX2u4nFSE7lyASxxglJU37wy2aZC5N8S+ePxuGCI
9DkZ9QhmQD+oBf+tt/Xa6yjgmCfLVOyWwcy1nrdA4iUvFnFuXXewOFIZB6+/S8sQ
Hn9fCqySepRpLvZIRtQCHSxa7jRN/9igVKUSN/AGNU662lAYwQ3VYJkbpKm74+FH
CkvvylgRlBB5USb44khv/L6LKEMl6lW8yySnD3ZJJEuGbO4Pr7gMPoUoWwSbKYnE
R31WPPhiaJeXRglvTQp/jMstAOz+UmeemqMncVjju2U2NQ8wItHZPH2fV1AzgINS
TAoVJdzDSYx08PakiYmdLxEwXTaPFWKgYAu1gz+RoaTTrrTKrdtjQvkudMwpc5zL
RWRiXGKcFJA6kkY3dXClG4eMVaztTfDnKuR7aCJhkXKd1MchjhBlZBdSoYlnLOHj
/8WdsoiP/YvMTxxasFvUXRuFZG8KFu6BrqkdfsVq7NPY3Ii/ZAt2Qkwdy4uR3ctZ
f25Aekn9qYhXLSkFAe5gOTbqUFE093LJGFoNqieqmTnytSAz6j8FotiEBKNGQCFj
7tL6PYtLiIamxpakGh0Rqr5GC6iNYgJsviW/Iea4tn5puguO2L5aTLH5nZxpO/rH
xfbDPWppbX+hubf9cnolCqZRxll0X+i7+pmgQJfYqCN5+c6pMrSM0dtUPbT0N0di
/5NqrVIZPnIZVv5DCaw9SPG8+aYx1T0EhBws9ZduKaWSAGjWJeEHoLgcmTKPA0e/
0WLokWZx0Mo79RsRhC3d0a7vVIqufirChELqbiQmldeGaCrAhcHNXIz6zYly/hH5
gqFWcZug/2hAzEqj1rAhlfsTZer2HDzMMTRNBYgyt1SnKkhmWCMN7YjCCmjCZhhX
0ZPx29sZVrpithr/E9BnJ02IDHqmsCL2LNorVw6oz2Vw0MMg57GL34A8D89bhn+Z
TP2Sk9CmqxZDSDI41ADNA0VCwbbku5DC06QTaH/IkMQCXaSdG2c+dw2565YZgTir
Kr4J31x1BRC7lXTBN36C1qSd/oSRyuahlKzjSWTcaFu5MKXY/XvVAK7kkvSCz5qb
8K+lBK7usg4r9kwQP4hMJ5s4S4rmOMRAb4LJcnsIJbO4ily3ilPR2449aWx7KL1S
PbGHh2ETEPe90vaADHjPhQLDFCE7t0bRYU6FOxv+iDwRx3McGW/XdOdh84rsTiAK
N+yAvUagzh5brh67nmtVXp/UEc7LSXG7qNsJBTDD5o71DMZwPNNQR+k6OtrrV+p6
N9XSnxFrTG8I2dgjsRdSHY4rkHZA9xL1/hnaOBdDQshoXI+oiQmygHoxQ6D1Pxc3
FZfaQeDPwK1/rl8KFlel5iQPlLh+7e6VBdegtanvpCmRnddCRPESt1/9cc2Wi8t8
4984CJLhLxb/6Kf2JJtYbh0kg7PmXuuRYbIvYotgosoZmt5uvNZU8f2fbEOI2BjY
/wmLYlOrTh0Pi2mf6M3iX3+PPHgHKFhxbMMiREyC9vf0bFuW47Uwdpq3AJ3Mq+W9
V/b9x8WMx3bKy3tPSpOpMx+5zrNG8NnXWNS9gs3C5rEsunnlYhQGIR0/P9qAaivw
0JYxCVteWJWv+EqCCVjlOwkjBJpHm5vGMcPt6yQy8wzqBSCmJJn/ZwBMUsAHULDM
qxHyqRf2CBxsV90hR0llcWEUndYRAE+z2Tf7IG43lAe8CAB0zRYLBJHNd4lalP1v
8DHOL4KO9e1udcw2Xru9aIhjjBbwqkuircRtDAbxg7n2sf82VlJvBNosdEmhhqkM
s/WEBgC1aZL6FYIoEqQvaeORvdpVDk2g0YB7zNC8ce9jOtYNK0ZdYRKfg9rw9XJk
UXl6NdR8GUWdcwfzXKcQBQS/ATW4NA+CnGLo1Dj8VTXwZ+C1C6KHCcKxrO5u/Mbu
X2GoOZ6Fij9kR6BQawVpV60RW/jvKFXaS4FUKjkqzqieGdNY9xjt+WWm1dF6u0nC
LMTzkBoDsjGANGee962fpcVORtOO5SqcaPmRu96EIvB52DKdaCMZqRGwB5nVCnQV
Na2neadVtIqvBqGpXgFP8yLPhERWrKhQ3hvNO+3yxldsi3NmgN/trVc8bgKrjNPw
zXx9Q1EaG+elR3nPkr9aUHxf9/K9f0BSfgiH/+8QBkV+IJ8W6aJbYlCJRdQ6xn5J
GerdK6R8EuMVWrpwb5pzFUE0kOyiXDjU6WXtyxumzHuVZaz6CQcZYbuej0MLGlAq
mGZYp4BLFs30uXktFKkxaMSaJntHS1eGGmtzz7gwsw55bZr8GTI10QTVWW/+7c3/
KHXS/2YJ6EJXdZfKW5EPYQh8gzZX6amPK7SSR48Fo5DwccToo9IP/6FxBdjPjzi2
cD+xot56Iw+qK45CdiFTUc2dHLVn8JUZzCAMJ7H6G2Zf8Bz0e+29L97odxPhHVbX
qE4fL05Kmdgzxifa9aILDbUitW16Appsn5i+LTRwJAXezqPzJ3ozOlbviaUGl3ZU
F3YfTx/rzYnebSrD+miKxfhs/uR7jpE5gzj7qq/CWBxenLUBFVzCrYskk8VWXDan
jFbM0mSaR3VIrD86eedQAmv0Ap7bisV3YUaSfJK57Kk3DW03aLUhDsKQO3ZgKvo2
jHfaukwfMNkxk8KmKLrD+huTKtLRKYKhs96XTbhUxi5Eks11oxVQlXcfIwn1rWfG
pCV5WpIbDok7IWlpY3K5wPNahlMskdfUkoVHxLoGWZgRqt9lwXG+hwr2nFeYWV6Z
9ZXJRhwxmoTCzpJ6Ylw9vLRBn1xNUw9fe/UBsinAs2WUwNXqmp+TUM5ZjMeqBEBg
eufPGIXZmG4rTV3sdP/HwdB91PNNw1MeNwVeTkJHb65emya1SK+Db+30PKNOM5qE
GIj1HcmXbMc89M1NY8Jt6ieFrqbkG7npWx3BGmyNQiYYxrKTIhwxI6IZ0g/kcvKu
jeijg6Qt0tfRC0P3j1O5Jwh3Qf9rLivYmxu0StLldR88IbEWHzIqzTlyGSchgeHq
p0UajJ4WsDWX3FCD67NZwIUuHTBY0IACOLmRGZKyDzEbvod3RSgX+Ywr+bKmgdup
1b01JwzkrUBBaoTxhymKu3LIWLVG03HpmYbex52p/W26DE3fpC0ORleUxLx3Rume
A+0Pxz8d7Q+cP/1ZNX+HVOxEP7Zv7qsYHVaIw0LZI+1dqnVcIF8Z6Jz/m10eWeqO
BgNSvBmHxFNJg606kHYqGMFPL6UN5J6+7TTpPQnXm4y68i12qA5NmCVDA7rMJ46h
TQxIsD7p2a5AM6Vn7zymwmEHDDXsAnMeVhDEHSe2BEiaFfr6INlpsrUAgU1sMRwc
UfYejLangyqvVBipLBk9LDYwc4N46jUqig7NaO1QOFG9kfoBDoaeEfgQfaauk4Sz
m2ZkzVksLGNmf3Jb1TwrxlpdI1voxaWnsbskC7Tts2CRCxaKucst+W4LmY0s1S/F
lrhT8kA1bdZVq5AGIgthfVJ/hZqdXW92K48ndjBlU7nzLytFWjthYwYUXq+nGXmz
IEKsNvl+Z9jVO5ZpfnKnraAu0zGz1Sj59RluSBLGJE5qtp4Lx9YXkq0k9LXIxP9a
eWsJyasZplN6F1vTa8eVaNIWEXlcc8qIYSQ81K+3xUVYLemeL/6NkWOzniYs2B4M
X2+zhTlA81hg7LuxL6zMa98GFCy0bSxClqJN3OYI1NGuyfMANzXuQWKyhFp8IzYn
uxf9aBlrpH2ATRuQSvM9rY6fkLUxJi5hIqT1YK6AZF6E/Lr9RS2A9Q8EvjS8FynP
ftZc2HNZVKZrgEEL+47f97es/oVbwjibpwp2ulJrGHllfSE9jAkCj4J2Y2t9DOR9
ARWWDswoU1F77mC5OgCSTi3fjCH77kEJJdIxkAEWuDTlchOkp1UWG1AhY/x799X6
aP802WUpEtiH1/SXjA8zeiydwedpbvU6mlHA86FJOm8rl93bDzSn1ngHwY3Y7ZS6
OB3MyEZMoYfolm1vgF3pkfG/fra1NrXdqtMdV5Y7YryA9Sz1GwCDfqWzihpVurr3
BG50BeAm//J9Y5e4vnB+Atitca7uqNPceFT6TB1GwzvRQ2XrJIrUpv2OdcO7U/9q
koO04S2jHtwiWjYcCrATXPbgbOg56LrXxn4hJvqlj/b63uSfMhjxIpHSmHgtl+yg
992+lKfBFd7HV9GmVosc/sa15CSCbfMkQ/tFkdaqYM8Ld1bZc/dFL3MwhjdfZaRA
NYkVvAh4tF2wHaoCZgScsqnrFycD4voNGEoGGMFNmH4vtjLF12Uo6rhiH59bRTDo
1dBgVATWbj1zqUNHRP+89fwKoU7/LiM7STuG6zrKujRYzsWP3HoB8vl2u32C7yZI
ska7Fapu8HsI3NVW/6zr8FzJONzppLlcelAxz5cvUV6TKOkY5gDvkmbB51XFcQY0
MBV7nD9YGfAQRidhgi81BpWrnKeXdb0kVPVqx97vDYPC6Bxd45zft3zjULjr0AdR
1vCSE/LMkVzWVBMCELb/qlGyhj5n3cA/7F+VmZJ/7xNssda+SJWT53JIKLO88jnE
5/OIAn2V0hCJAuOPNIX2bJegmFOmCvo4ON6qBtl4zkn3rQ/sKyW1mGq+HSDBLtJg
tC2J4hPlNTaWNiIr31dTC9CncmZ5RLLoTjkUA+z21P/ZFIIn8gozLHDHYRr+i0JF
2vwzkdwtFap12mlHsmPja7EbmXc+X/WeIW08ba217TatjCYPNpqz82BRzBQK/U1M
Y9Mrwrg4UqNSJy4YbiFWnyitc1NXBx99vYolFt2/s/rV+WU1uGGPjbc7e7DVpHxU
OtxzcHG4771gjP5oGblsUQvny/rduMc5bbYXKQfHAm+I/iyLUiFDe5QAquKSQ8sR
1Ay08uHQmUmXgSB65/JkSyx2xQgy5DkBVt2oV0tUELNqdSNGO9Zgwpxzzf+mGbL8
9d1C5ef33MVPVi7RtMogU3mjJg2eBF5oyMx+p4hcaMarVrR9ijFX4nnayk8MWJZK
/wfy1RleXPHh3rFAblMtgXUu/Y9IyU42/4+nCNCDY4YpKDmIb4xytfLOl8XmYVxZ
PrBGrhGMN0lpT1TeGeQCuj1l8n20PmLWp3bRza4S3/nUqHqY2NilONfqJuGGO6E9
ascnOUu/PK8YIeQlrI6Ndbg+gQDuYPWxhwJwx+Az6W0jY4VGviAhV+2BUXNlb2VS
jqvWrr8FyIHh1FM4YFZrzFqDyXJYaO9RrCFO9CbCF2T+Mck2oXTR0JZVkr9w3F3y
t8yL1ZZWRmAp10NotfwqhZPitc6QVy5oxaciUI5lypG57WFG/tgtwSAePsNjS1ds
uCFXsgiZBtUOhic4gZOSYlAbHMbiXDIvud7Ijmg5QAvcCsfUVyrdiRoW3GAO+TLl
x1v/nQ17AfqeEZQEkL4xV5GGRACRKiznIewGwt2xBxPrYdEEGhgJBzkOgo0p4gX7
EHq5Cy7dD5bzatojGBu96lXbnn+GpUQNZpn3i3fPm1zaMTlBX4c6TCn+RPUSJL2N
R/fAhwc9nuaaIAOOZ1egAYo/7Y2WIEtiRnSmWWgvzZsnmLTw83V95dcQVRECkCQc
sshbVzUIVhd5TZuw9hyjWpgeoAXoVDidFQ7Fb2EMaEDvxWNz2hdaT8hgEcL7g0/e
Aamj8sj8lUD6RkcDfXT0PjkA/0uCpwELgxYGmvYpswJHl9KkrxNUudXcgub5ZClO
t4zef7mQJ9o68OAegoqKZrxBk3yuV7urNtqn9/X8D0HapZKCWIu8cnzX1mBOrs8l
xLjr6ckJ+niI7knzgkc3U1nnc7eGbTC7Cv1ZZIhMGxoB5syEAed/GPRGMJxzBNRd
/g/tnECqcRm/lS64RjtkMr+LY6HcrrKSJ0xTDfvyg2HwZ7vGxTt/ndBLSHRK4fc9
aSLjJwQ5y5F0fyLzP8fty6jpA6h4ED+7IXwWc4d6Q7tyrx5+HNW+SEfK406R+cV/
3J0Kaxl0b+Z9RDI8T3nBlN0co6oz5hHyphrOhqvbC3+3G5lHcbJfG/7On4NsVeH8
BTYKm7DODsAqK6B7qei21l5mYEBsE0V9GWBRMIz2sRC6jymuvYDkOYP2KWCc+15b
xHW4nHwSsXGLfrCNN76jJDZ+1Bv0vEK2PtyrYtvnsckojZayyBXM2orhqdpnr2Si
GmKj0emu/phomBZIuVHi82BEnIVPRRRybnG3kv5Rx2UQULODVd6EVD0fgyxlAyLQ
0pR1QvJRd15YUfT75g2kSekC0lMtWATGVMtN3C4RQNQn6fAfLKkot4muadmOi8hm
RMFpOADk68pzkjJwK/dJ4d0zWNdYIBU9xM6bpexeL4AesCiwnpJbGF6m0CYQc+fc
9JY7W9+CyOO2ESFCvqW0/URI+PqjQeMK68sOwpqquW9Hvl+Jy6EtS4a1vk13+MJr
xzLJudATAcOMjMEft1Mfw5zcEUiN2soKpZEvQBT10LC+cuflnF0g3V8wbbiFiUw6
oIce2YMW4Rnf+/+0zIDFcpWxa49szKWFx5Ku03b6OlsTHdZushe2E1/xguV/7FPC
2AB3xhlDLIgh5YbsFeENkTcjjU7b8vAuAzI93uEv7xFMcTUo0T8AcFZAvWOLUsyD
B+/rqXkvGpCMppvW0CTqLi6NgnVoyQe5nwKFZvWiFDJ79QwUh/fD4nY/RM+uDxQW
bLzPTn+J0jtKhCNY3gPQJFP1BnRrGiwZt8qho6v8jVeHz3H+8S/2EUkBB39gEEzK
YKrXqPSFfCp6G4vGi78DbKc1fSuazeWVAxIT/ZwoZj3uJ3zpNlCAWX64rqn8WLbC
2mVqkba9+v/CtDxuxyxOxJ6x8Q1/C1iNtfpb+pPfADVtFV+F1MG0xOcsubZStIfM
iqRmWM2nDH1bscqBkJazLk0R5cfPuxuRvEWlAbVKTH9m3XjNKYGqEZp16KGomtbf
N4TEexiWzIUymlmkADyr87pEmXACH/dCpWPm1ct2Zyd2NUVvE9d7OcWRxEJK3EVh
zYNShahsKkb6REJXmeBpPrSsjeIw2kYnFhzA4e1ft15qY9tKbe0MBD743Pve8AiW
RVO0eYkh/yRX7+B5b7PGKf+ZPFbgzoKCj0lzG4k0lT/hVQ+WP6NMlMIuUIB9IVEp
tS4jOex0/yJB50Ngcvl6zvz4sIwtckxcFXOxxeu4OZvVaGEZUD2zeBP7aU2Rl5B4
v2Lqyb0P/NKxtMv6TZ9X2wqKI0WfAdCdoKY6lFNqTgyP8XRGHdVewMa0nEyRkEKu
HVG85t+Qv2n9zk+Ou0HWzDwmi6B3TA1nSo+Qf7jqNzr0LC3bJrX3PKGiF8QbzR93
zWJ8gZoRMmY5UX2+2bindnntHVOcItYf7KaAdkq4Ruc5SzRrQaCKRrwCLC67oiVT
cTt3Z76wmcFj+G4LE4ZVYL62T3WeEqw40B2+2lMpK8ZW/7fP0etz3Pritg7oZ/fQ
wtmld97aQ/3QGgHQblOpOkZ84nu7sBqdPhjTSLgaHF11SyIHZZpO8KC/WUhAiKKg
hOMCh2nusyNvsaRQKoV3bjejOvk2BxJysKgzJTLvIMRJQfsWcwwfNzOmMAbkqG83
0b+K3E1CRF+8syV5FioMYSHE38jjUyIR4vXEwZHIzOaHt4m+91CYbza4V4SfWzwM
nbGF7CBE8/tV6G0omAUJbpsL4FJaSAeP6zUbkj2kRV2jq/c4wLPcSpbbGboMMlPO
IghsT5tmZ/oVywhrUfFi7ou8AzYcShS5X7om6d5ZPt6teJOGE810UU9UWOdDvnz5
mVtIqrVJRPvqu9dJ9zQ+064oxGrGUrIyzWv/uk8pFladSJIZVPxC+M547AFfE6lt
L7WxgHZ0OxoGjhiI8uItv98VN04JTc4bT1o6L6XEoQR69JB3xpdnXWvpDJCHvVMM
D3P4h7qrMwC4gD/YrWzW98vOLIhwmvM/QHSq/wzIAGWp/s+Quz5bj9uJGenDXrpB
q2G3eLxUa2351yfEHMyqCrWmrz6oCEkWwJkEipl1+1SJYDa42olLafqIUDVNpcPt
WkPpaICVeVnmg6c8LOj1t7TYoToBdraBrhF0D0dV3FFsYSsq1OeYbBkv8RL1m0rn
m8w3J/ZSLSqh08TDzKWIybfNxU0+5ku1SfehC7xSa8+KHl6CkZnuanSeu6F1tg0b
X13y1ipJFAlf29NhrpvBZfwLl9JwVCv1acFJEO/NdacSqI04ekaUK1fdzFIUbC8B
KHIbkWi3KBbw+ecA9z7CnSU3x+Yrxg9/WT6fA1QNfJnAV7GkEZYKF2KfRPc4ZdF4
XXyKXf1Pv1WX4k5wD/g7QNcKTF5N993dRlBh3TkvlS0fuoe4B1aodhK9wxgIDuG0
gbwZMlx1fHvIKGJ/4JOH7YEX9fiOnTK2wN9fjsWIDRJZYZ5bfQqPcch03axi692o
09jUgzjMd0Dc1Lpdp5XFBNF0vq7ww8A8kpj95lrb22eyZm3CGy3xe3OlJ2B9EPE6
I23dsol0E1PiWqAoBG7HN3P/lFgH27KocnyIDHpQA2p54sfplSlyQuc8drzrIZWg
WB2Fk1qHjXe39PoUSEdjATp3vym/C36KSuGRECDqld9QTg/3NpcwXkiEI0ufopR6
wf2O9gRNwBmm3/0VpcgJ0v0e4YlZyt+JR/WbvPjPv/cldOPfw9KMxK9oMJnlTqf+
Xr8SEDnbu1Q2EJ/I5i/I3iTHeljynfqy2y1WDdWA20E3fwpzfN/Y317YbW4G5cag
RL4O/CUAtU+eZzS6CyTwc0VX14Rfvc6Zv4vDAOE+COhUDq3el/XHcTsGqRxHeuYJ
f5FcmJWXqRpbNXU8IXJaPvW3k41RB+DtH0+vdAuVLkGW6RPofoWGHD8xq0TtkRiQ
RI6lR7Pgef6HKY4xaH63vFoBvKj8DD5gUEmpuaH0yBcwM+gJVWs6wXWgDtXqsPlq
Gs6f3ifatqmVNK5Mt0Q4iWOYYIUMKkJPk7xzw0aWksoumf/7DkWokOmWWKpuvmLI
LF4ldCE9c2Ra1ovbwQPV5pdK+OcDpT3bgolIwrdoUaKQQYTDJbmpT0i+rlx1cSkx
02ZCZLySCqTUIsLfcBwJZMPwMh0QtfnFZE9f5Q/O4U2r6IFbK5On618Uy0XueXQl
AwYeKUsaoLywDbVpEyfBsGCeMt3tcE08/m3wfgGjbXCIumpE7Y2sCXvM+HZ7jbRm
5fOSe1zGHmjght4v4RSUacn1yoVCqEuALRNYEurDIgD/uwLAqkPDIm7B5oeqHUPB
8DObPdb7lCbhx/hQcz6IRhbZRtdklro5vwBxyW5vvdNAeEiifONkVQQqbR41hWMa
97/axSJAvolEGwC8/+SNeDNYS+MEDhskB+MGfhb76gjeqbndI2/9dQBJ2qy1Py2B
uBPUnP7hdpjc2IbdMf6YiwfeE/t8706dUulZsgU3dEBM84D3UppP6BAus/frG9BI
sqh8+OuSgYFRrQg6XGWJk0amoChvbMX3dWswNYxA+oDjJGo6oVK8VLvOZ4irxIIi
ZOAIi2aGqx4XWP8zbWrussIOdx9gdaHMXJbGUaPydj0MSdsW/wQIlGCRCeveYo3F
pBebpPsEWXC/GLWBGStydMmcYPhDCB7G6hq05PHfovJKQQUqCXyc2sCoWcSmUdR/
Q2F1t7rK0UZOY5+SOmUPDCHnSmbBfL5c+ldfG5CO9y0dkMd4Ca9l2cjD1w0gHAI8
2Wd0+wB64WG3vcqOYefcOBB6vN9psSN77xdImlvInU449LdbUWWHWRiaTDpgh2jy
3xleCuCRYFmE4JB6g27IF59ZuYC9KXQZuKebx5nkW4z1IwD2eAQlVjyxV1vdyLF1
COOOPvmQHaT2xFwxR0eXs2Ct4OKVk3XVn+/n1EA3GS/t7cmErDhnZDePB8eJXXi1
ZYhCOeowaAtU8zcSUgvKvOO2zkeHk0N8bHloR9Rzba0ziA4R6aokMjZGrTyAJOF9
NrJbQjOFpHn7h8r1xgWLoiiN2XS/uAQb1kgfMhjI9QMu/+ryY9GKzWxr85m5/+5B
J+KQ0W+7VNFg2ZOF7ZqSNwa9RGIZdRYwRFVyCz25BXDPKHc/TWxXHbkjmmlHfRc0
PmygnZKedH02rm9T+l3f1uemEzpvzr/8Yet/2Qd8biw6/43EdG/OYJqhNP6OK57u
1+KNEPbokpDpRWRit3C8pfoU5DNkLZSAy0jUh+bnFIzyWQ0wQVe4YMHgOglNNQxH
lgnJuyv8nR3d3QWj0zfeHq/2rXX2xQhU7KpcO3VnOomvqIXsiRF4NEIpJrC41g0o
NkTa9OZ8+m579IR6klbwKomTXl+4W5Pfkt35SKmuYnwWr9srxt1dAbuQP0SSehIv
JwDyNQ4wLDXHJyObKMcEheMUDMQg1PnGvfCSiKy3wJ94NtmTJvWVSftiFLcE+Sd9
JSO0SidBKFR1RF5RZuUtRQ5FgF3Iu4wSLBWHmB1WVmo1+Ov+p0qfR5VcRJybUaS4
G/uEw2I9fharWRxUGnBL9+pteO3BJZfi880Uz3vglorqRfSJt2FobTr7hjzobWZ/
Y0WhxAcCZeptokvtpuUNvinrQLZYKqRGlY+9FdGWqAnLqasWhY5Av8pa15zsSuau
rR/iJyatiZy7wPwnI3EBC40YMNvGnDfWCnu+42tfNYhexvRIDSSUBkCfm327C/za
1lw+R8F8fh3dlffkOxgy2LS1szuQfFKfDxMSbFODzkSzMCuc2ur3YtzdGRT+O1Zr
Y0JFp2kVu3bQ+QeVBmSd0sW9FAgTVaayBvVqYjLezJMcddlUOX3DEs4S5Mu+KwFl
0l9kjtpGdeDn/Z1y0sRzsCUdCxqC2JJty2iPS/XNIbji1En170tuHPrlTxxm/0z4
GhWGgLV28d5+3ZJzpn1TX3u8GpI207a/bpwZLhk+SXh94rwAOSluWkSC58iQgAfw
EQArJPKQcRlwPXI/FVGs3i5l/Ly8SfJFLb7fRxtCpcmrwePGp5FCtCECtKRM+qeL
KiTM5vczkRQvyZpMjJGArLRNOqJ5jFnGdJkVav2rHoFYMFCgtjTevLAfJ+Gh9dr/
5s8CLdNAb7zMi0Qqlcpnb9UDI0oy7gWVWOgpaGMCFO2fu3z6DBTJBXhP4mE6J5rh
cb3WnNzEiC0u9xAaBGEBW7zlj6Lw1gLfvP4XZ0NylNsPeS5UCeY7F30yUSvTcLYu
LJVPOeDUY3Fou1aF5EEsGFsVLAeq2nWk9IY1gANvuqiErgjXcuCVskUvbfgWjnce
nFW2W7rCyVM7BYG/HHFCRSyaK5CWgDy0/G9HZp0b4H7Aqd5842nlO6VuiWBPSkOy
VyVzUorK/13+m/8VgOvmB07/VkQeORQyyoKWN0yuCFOnrbRXRAlydZdJok9dwhpK
WFIQc1x8dG2dtWuc6ZA8tEcFLM9rKARM9sL/kMhqd401ryqr8D+RlDfWZ+HWLz7F
GXTg/g332ODcJEqFbvArewMXjtmtP12VUHMq46vDeYE+MiZoKcj8y6COHm3ZIXGG
/GQ7uRDVg422TlApPtBuQaweU3w/k1qkIUw/5bkmSwg1Umd3Ji1fQuM9NfXNovsj
ox7aRWalMDNdRsm1T5wzoB9s5sz/e9wwOILIR5+Qxj0Zcl6cr5oHyby1LFou+SCi
hTszT/1qgfp6al/q2y7LtP6TZjDYzSvy+fH5fTcVqA59fDF36rduHr2IpGAFeoOg
gIBJybour4HJ6IKMR2AF10klKkKYIUKJgA6+3IZbQl+74XvSqtSstCChAr+5grec
/Lc2cdYeygFzfsZNXUSxvmXeAGGurdNdHVgveAW6BPlC8UWp6/fN13USmRMcP0JE
XZt2/UnX6Ec4JpRjZZj433f5Gg4VD92SVuqaBPoTO8HdVSO6JuIL2eF+4moD0sVc
1VmRqvWdjvzYP8fo1TXwdZ1/6sRG0cyydL6ZnfoVbPaNNAupNQ5W6THD6SYnMxKv
M26l4+KJnUPkWl3y688Pm4T4Gg3VbjsGPm+K3YW04lEqqZNgipxfM97D5a/ZdHa6
zJjQSaDCJtvB5LHljR6Eyv9YFRL7Iz1bHIS5F0NH5tvhuICL62odvCH7eReHxRLX
Z81IlDmNwOFHERTa2D/H+ifV/nK9mL1Uqj+c63TPaoDD5m4CNfOGb7FkCXbK7cYl
5OxUlFyDGXc3wIPIPX7qCftMJrOxa4PZ8nPtaByQWDOCaaFQBMq2LMLu+dVayoVE
8ODGQ/lRtQyNrdMRqIw7Mi6L9xgr27lPufr9IOB4w4q0hNEjlEdCdb/M8LbVd9eU
Sgx3UujWC7bRbCOX4zKZ9o1x4QuoJ9gCmYi9EkZKSHmjzq5q6CnIcaz6+E5FucSg
Fe6atfSm8d93Azh/JTEtS6RhpCPpvGUvlsZ762kSGP7q+XB86foWkoDFBucURD6Y
D2MBk7tZMV6m4uusAD6CdS/kH4uQbnbia7WKJTJy5MnBibTQ3ZmI3mjEZhs7e3nq
LYgENsb6dqg/oikKZb3+SyRQN+VusmJBsleiCBxHzI62C219lDN11ETxvGusTnX7
apa2YYKgjF6FF5C3ft+Nbn/QXRpVKfAeCtWu6MJADnIG1N0MuZ764iyUawSHMeAk
aEfPYCNY8YdjMGkO5QhgKpehZbv/bYh2XUBPa2CYmVH5KvaWGMqxNO6MAxVnRxir
OigR11oPsxhhHy5mEI5A0gArUUPoLO1LTKmdXn/D/caOdfDHNqc/yo28dwHze2on
5JFgAN/ij+s7DSbTao7ekxaq2uYml07tRrNxe2XaH9C/L+M8LndPPv36jhTMkS/h
ijkt/1EbLSZMVGgcWxCosUYswPo2+8LNv9wYheRRFwoj0gjUyl054yNqOjK9TtED
SWfP4nvcoyCwoQxXsxC8tWjjDSTePd/23xLZXV4hjsTV1ON12wWDkJvBRHfnhHfc
fpbsRrdfGDoyp7khb7m2gd1czHyGrlmdRs+cax+Oak8SXwVckaB8n56cvVRS/c9t
x1AE8chl4yBFgEFpcR1EByAzJr0TlHsreVdX1GsJ0+7C09Jh/3UUfGwPWkE6IYww
MKk3mtZac+F6ySZsbimYZuXSXUOeWRofuaNPPJdjmbZpAla+0rP+zOU1o5KPQw2i
I2HOE995R8eTbUWQG/slJ+jD3CdRV+syNCOQvoUcpi8eybIQ4VCSf6B2cQLQSlE7
MkRZGZn0AjmDg40O3UcXjL0FBrPNDST99I1lmrc0/Owmz3eZs2uSgJfZ8rLCeOJe
UBjzar429wC6kfz/fVZPip01ygO24sd+5RDf6y5YxOw+I0v3yHTvyJnd9mew0vUJ
CClEgOTe1vD05OgQHiVB641FFpz77H04Yn/2fQgK5gpfjKc4BhokCIgQJYyhCzUE
KNkey5plCd9jUubijNF+sgR9L1sosXQV64AgWa8Unsp8edyJpRtAIO9v1C12RfuO
3S6YrDkWhXrj5p+kXAdcXJ8G+B4LwV3X1Gj6AvYcl4/CX4OiYx4DgyIJ3NcD+qsG
cQpSBN9SHHfND+gw0PAWZs5av+/Al8U2gSIJm2ROFfyRKL3QxkJxOHgp55Cx5Oku
EVSOyBwtlnMa07lySGCAGcXP5DVMh89m8rkSBmk2c3C0UBEUzNYhKaHBLe72hzN1
8RY0PZu1x3b2oop/pE1sFxKBunswId3Uwe/AHHDou467gPkviRJlf6u1HzjZ1rtX
HJwMlV7O6K99X5NRkpILBaS5DQIyS3PIsWKZgZ9U5cNuMAO/ev/nYU9o89z3nUF8
UsKPNt1/bx8WjOP1ZUSl9t6AsahkR9EONzgueVs7/9TZ9N0OjqbZysN5suHwnLvG
0/8VwS8tXGJ06GFUSnyO8/avp5a1Bpwp9ywkcKXUGeBrIbpQdK1Jbu20pnWeqhhM
qjs8IeF1P5u3/Cm+efF0ycijm++8PmYiOT1ve5l9F/bqx/pqxuQ2i5UTa5xF7DEE
XcvHc/jL79ymGRHKjY1gnwDBoB8XGjr5WCHKZiSYykSZ/85zTWnyzssDIeT7s0C9
lh0l1EhiuZ1UX5lFban6juLnUBQg1heHgVCOl9FyH67C8CheeRHvludOvcbNNeip
+xP4PtpWaDqr25LOFQt1GPMsKuP91JTdDGbkdkZCWwzs9vrra0BcI3tpmJ3+qlu5
uVmxPoF5xPs6WS3V1BYMB2MMQk2pngnS8IT3uZqH/7WHJoE4nyzczCRQLl5Vyjfq
2qPY/8JUFzzyVfMCIWA4xKMlvm9eUnuL4msGppb+nNeQStLz5pEKTtFLZPKxejfI
k3SASXnJRgPNgD+I+7OJi4dggTDO0sX4daiYKkQuC/1NouuWA+LztHF/7Pk/hld1
bhxCybU4vYG9VkY9eYA5wWCtEw4RVk+HJkK1FLWJvPzn1YaAHadmBTd1aexhyBXm
X6eQ3+4aO0vyPzHL4EDDZRMjl8pPQAgPJr+YGsUgPUHggodTpcF0drLXKQSYal7l
xVj02cRuYfaUfv8I/azj+Bt/6sqDOCs23WE02JcF81KzykGxhKs2NKgUDDB5PGsj
jc1eMkNpc0I14i9EI9FsODoUenqXTLGXq7B3O9omp94nnqD6KE7dixx5G4blQrrj
v0ozsdHdx4g4xHNm0V09Mrw6sTpLn4fsqUifXfzeCyOU8Mk3996QUYe5LqexZOxM
aRxK6G8/BOGSl3QVTCtpCaDjaDO/8eR1KRHphA9gDn+jpXLd6SLQf8r35EtM3cq8
Gakga3bo01wrDQe74ZLhRXFrN3zAgVq4xUUO6NX2+vLYp82QE54H/p5vrMJk7Elw
7/j+q+9TJ9zT37NhcRc98nQTrJQXKy/EXKA0fbUml7JQqhh0ya4ky9VahPa/8izC
WJ5RIbkvh3fKeZemV5YQWtBDyxEGZcaQV0j1hawiTcGmRjImZJgHsXegogr1rdMz
rr0ntKmoi4gCzVK7UG4e0OnbFckKZsu57tB4h3pAvOYrRJeIMOML4TX/yd2MbLHx
Bhk03LChLZc2CmI3nsluMPXK6ixB/xsElJAh2cv4J7dACIj/ATWZz3GJpr0C91+S
0O8Wzyliec1z6w9nNX4xLFJe810us/6P/NK6q5+c2ZKQW5Eq6PDQ2gPcO72NF0Wd
tzjRfUKxkFWpplhOTM8zPx8Xi2CTeF96cYD4wvTxeqfWbtF/xcLy8XQJWiWlmD6W
CcPQWteHMi9LGati58CDlSgoEPQG3U4dlyCj+0sBnZ4QuNqeJGmVJq7XCOCSBohM
hrIdbRdlW0Qz57cD6Jwh3VglTK9yLQuZoW+naSYC8Rfrj9aosKSd/ckC7fDwrMJd
J7VU1rfyM+Y2Of6sRLAhFdmsyeBmz0eHIBvH+K032+kZygGYJd/izws3EMpHUe8F
jzV5J7WVzERLDw8zB2c4IymFXGdxdWYhSYVVuR1CP7Uh/K+NEpXRtkiXUrjntE7A
vmBxoOQuI8DcJfmLbYOLQoe1fLtinDyt1Bo77p3Mw1lmitF3Vch+tTwNqoIna8ly
7QFZHOQxSEg+D+Mg4aM+YySgXIYMJdMfFt/FeYDedgst7vhIFqNNJFLwlmQz3aQx
eiGVkE12h/hJnQLWSy1tKtypzz/pBrMx9wp7yKL1ZHcUnw+vhiC5WqsqsnGAS/nl
oOknFUi3gJpD09mjGxCSrqUGw87ay3T92yqsbzRkpjtn/7xjaRtAGchyqzkku/gG
+gKQWsUHkvmwviZdtdJh6sSoFhxrrGELtH6GlrpEA/+C/xf0U6CDuphCFeievm4l
oRy1dyVFsOqfKlGgYZTRI2vIvGT5xUOiwG8KDhje6Y557XuqZ99XiB7CeG6uYWwo
oAKQ9DuBkMdo16Zknp6aPUVHyUBEBOSsRCCFwqS9badkMZCbe/y5aJl0Fvl5UDJT
me0iR32XQxkemQ6w3oyKp6Ik2cSaD8KQ5luxwg//9qvnsRnWwkUTfDMe5B7WoA3d
O0YdQPGFUcR9AIFtzBia5BWlD5ymk+NU/EJbzsaeN/V8QtiyAmDT80FxsZ1AX9V2
VA5YwAduZ7O0IcnGt7capDBCp9Lo30oBZoUO+XyxLs7Jyr7bLJLMYXKa3Y+nQhfx
Crx4nvVEt5JJyNfVgPVL/HHnk+Nzngf4EkgOq4DQmyCl30MlDHFEohl8Lzo/kyLp
dN7+GfwTaagpLzU+wBKYzxjSLG94Upjhr4zs7b1H2DgOzd9bJQX17WEOeHGQaT/u
oysTbuXnDBhTnpdDut1HAP4Bk4flG8IoFZ7S5g9adyZQw0RiWPZzW9Xm8+x6NWRj
jp+/TA2nmQ6gce+NB+H88jwTPBqeTeSEtU6fYenM04BSgUbjagfLIsLg5TfxzB4Q
sVa+p54foa5btlcJiFBSQY/rDzmU/DKSWEHmDpHU5kbd5sqP1XdRfvfkh1Ypx0Js
2AjE5UDU6WjvTfr9AMkxAA/QOosL5+YPWnlN1Ay3osxuVJYHSgJhdZpLLmgfEj39
KVTYY+JpKtb/HQVaMgOUXcR21vh2U0T4x6Z/RxhEfaFmAVVn1uEe0PBE1zNyWvTK
zrTwN0DDQmSsa/565E83wtTTegi9MP7th5eQ+3xJ5y2GQt4Cm4PsyF4R5FKtWNJD
rmdkS8gF9XpTx+Pu1zJZCmu5J3uvNU6qbqz5CwVb4KLUC9nRpkkDrC1w8jX2N482
gwZRhVqboFTyX67Pb5A9u2SxkO0Jz7D5GnjBExnuk/Tnlm0CPeWXeEoKL4ozTLDR
R6AHfZGFO2ix2WIOkISUCcBfNJfUVWV6+IjukTrp8K4UwmX2tK1INjQOHrey0CB5
IcvaKFaEE/ZP6Om8hK8tg8lWwvEsGoahNMF78im2ZzZzGxB1oLpq8s2wq8rOqiiR
vz0XdtmxsHO50ySDr8vEFZk7fpmK8zemhpQMwai7Qp5Y4aCctDTOQ9juY1QjnHMf
SbZHU2nPCNGlXhV0ZevbsDi69o5Y4wKL/P7Xpu+fyFPlHcG5xh/lC2Row3nO6t42
/pjtzEEl/qXX/u/q6+h/Em07PZJPJnY617ym+yQGuGsL9USpuXwMUWQ7QgOz7+gz
CSxsyWNiJnl29L3Y4W+zeTFU4TW3aFlPKYuumdPhEEfUYI+7f7tdPdg/nC2c7XTX
4K0IO0GVMaFs+RiikM03AGkzaTE/X4NNaDIDJLhPthgxlzgPRXnkl8aa6rWdiehK
tZLQ6wx46p0AgIG94jxxdlccLFAKjBcfzL8gAXVHB1s03VJ0QGIjEUszAKKN73ib
CNa0jRtALT4b94PZ89ZeMkzw4fFcbL0q1mnRqmJUQsGZeocqoXowRqnPAxPb1B6y
mnmKd+9fN5WElUQ51+OEWzln37SBe1BztrMsBtlX9OUkOVdWtb6LyE8nYam0qi4i
BxatlqYBIn/BhFdZD8EV8Ch9YlZxNOM+EBSfpltXQDrtySFsgpjnY/B+f1kY42uK
GKyFTqPOhTwccs/XqrXJPIyiA6FIY2A/AUXfr+SNBLeYRzAeEmlReedoZlzTPtAa
+pju8w7zla1bPE8J62kaKJluW9Jj9hC7LxkaQjXgAVgN5TscycEuanRLK8pjrsS1
xyY35tLv3NuRG0nbTKPLgN3MsFI01wwZcrFS+3s7eO+mbSbTZAeer2NEP0RAr2Eg
Kwo8dDzFyDUjXgu5VqBbmZf2PcDRcyq7BaSaiyEVP+uMQMhddCpDzoSPgbfQ74Af
E6sREb3j/M6ebr6YzKvtqShg4RhvNw6D0fButCkfCdnJWYFv4B2j77mhMBwQgcFK
q/KMFSTZTy9FO6etSn9E3FZ6U4YyRKEIuMs6Dg293F68AVbPwhF9GG0gTH6uFeFM
s4FW+/GLTlbaPhRAkLlXc7sOSWBAmDAdF8lKMDTqzjEXkhJG6IBXBHovsJRBMhCc
0R71HWkXxBzI5C5kjR1Jor6I5Ig8hLsa3tNiLxY3nDrkpO0FSxiODgriJ+SqNbKl
BdVN9RAc7v0TZacTV7DZ4MZHx5Qg2kaiJ5wcTDa1QnbzG011uZlX/Ifdgpb8snAZ
SccF2zA20nlN9JT1a1D3iPW3iUPk3Kef7kbVVFkcvvtcKN+DlXX7WPSqpu3t3J9w
bvDgPpFUALNxk+YH/2VmmAK4jkPJTS+tCdDO7/Bh4ceKk8r1Yws+IQpyVNQCU2X3
jfz2gICtia9sj0CdlrIDqy99lZAxalzC7TTOIe8sUmOh6Cgbg6KJAVUosnaAo9W6
Qx10Q5uwBPCETUcIMDzEQEfvcoh6RSv3SXrAYcPsh9tqcubNRUXRkYRW5wxS7X+W
k3U6TmzTynLuQD7qV7B3XV1423fbqJ/TnDH/GmhVz0ywJlIhKL8YA1P3gNh4Aaq0
r1oPcU44Ea/XMAEu3SXaaG3lJJgjALbktiK6o8esnNAtV2oaqHi+StqM92n0Kz2a
SVphjfIv9PW4qSM77/bik1ay8Ie6oqDjmSPbPuCDnhmSbGE2fdSTM183z791lH+S
cG3/QEqYVyi+8edLtGB+hj16NsxWFmaOQ4M6zKNRU5I39Wtdl0/hqM0PAW/vDCcA
kyQ1iPY2pV4Xv5mnKOHV5tqjz353j483gYCLOO7HNoVC4HdP/0RIo8xkV9mrOq21
V3DfNoCvMdaXHty4UPCRYyi5uD6cqV8bZMTnKgIytWOAjKJIxZ2RLIm/vuza7t/c
12smg2KQpkSPZykuCtnUez0USOIGbnAbVOzP9ir3CSAX4v0aIi4FRs68tfR87SDO
daCH427Al6WLUmJknDHEI294lAtZYf+9CmAZYtYA0DcDyfdk2rat8FiOBfokXghy
DK/F/g4CDXiiUDO9horxhZ77BZTT6a/BsHrMhtE7gN5xg3ST6BvFV76Ax29q3Wof
Q65Fcfb2etlOID7yT8RKT2Td8i+Om6i7QsL8DuCFUZQoNIRFZ6LhIfjR6fgMyxLA
V/XAg44uoaUpKNSwhWDWTDzZWXYKBjbTAv72NTquMU18hB3GyNGY4uQYJW7kypEc
QDr8Pab8+d5TlIwrI7cCKv0gf5yuLXOJKjQJWGduNEbaGycQoHVZMGZJICly0A2f
GJTS7U+JY34F9gvufouCc9R7HPbxCRP0KiWz1lYgmWhrt/pGho5LFbu+uP3830Yb
g57eJSTObNcd0fsfZrYdhnoXuVW7Ldtw4LozpkrRLS24Q8knbTJWqzScSgj99H86
mciK2ULgfhMqqTC+iX1Li9E4IWgJe2T/Pkhg6ZtA3bW6ToUVWqT/tEwmYosUJBsr
4diRc3NDcMDpDnUG7TBc2fEUvRq93LqrQQzGDrb/dfdPViFN2LcK+0t7MmfT8MYR
SH0K3O/kXPRBkI4o63p0TLp/nDTzCEhHWrMq6EKNzIhCwRSPuqzNEcjasEP3LUb0
eF6kIvKqQX1Uw8pbQx02EMj+uDRoXfpXsvrve8l9Tk/UdenXGLVNmG1HZuUaFZV2
ULRKKzuaBWARhQmxcbk4bp9crC+mz9mbIBGvmCoHCdhDmA7Ku51n8/QVB7JCMWSc
0wdC4GcPjSKYNfZPl3fpn06HB22V8qIxMvl8rgmxplQYX/Wle1ZorWE5tcxkXL35
GlW5lHvQ4Swv4WDqnTFXc2L3eVYufHl+n8VErjp3wlKdQZ4/0BF6reJHiLkEgDGY
EW0xBej/zvrFvdnFggeAl3YMwTDvTQ+zh5Ah5jA8QqBWkql0VAoqkbxH/cqU84wh
b/8crV+xdioIsWepCx2OhG0MYalge9Upb+43rPBym41qnkW65e6H+X3dLox6xpnQ
ghUk3kn1hc5F9GesCyb1iYD9yTqicxlrzZjtIYqDHwjx80F1ZmUQXA8MMUwg5MLT
sESIiPkbi6uAIqF3wcr83eZClzjUAE7E6d5KoWkymYoN7+lQASMyxXm+rWFnRFCx
5uZkk5pxxzyU0KDzPNTEh/fvBKzpA3A1Pj6jn7GGj9Joe+inVEZm0YBvTLa/J5Fb
QG/19Eh7A1wWX14HrirkFqrLKdHgsNzsURJVYq5Z35BN2SzPv2z8PAne8kNlrO4A
WzahbGgbKTSG1AYF0QtdqCFJXcZtBWAbYCgtKc5kTpyJxBgLlusU/35nx2a9c6Fw
NkdBIqtp04GHmT18Kwd1xaDE6IOCIl567PVPA/GPM0+xLRoQ85T3aTG3beN0CnrT
hxTz969CN3GBsEeegRU7ZYu06gF12z8yCzQQWXTEW5+RBLrb5R80Hhak7S1OhlZs
oOHYkPVVJo40A5Cm+l642dSI70MVDBd9+hmkO5S3KR8hF7h+8A3OZ5MSHG40IXBF
bWOd1wN6mdDsd/Z2jadHhBwnLCNBBfEJ0Iw8eKW3xha+ZiBwbqxVpqyPIYqg0IBz
+UhcGBvOkC2qGj1pKnimNE4fSvaY8C7paDSoxOU+hKJZk9YJe8ucF+WgNjEYCQ/L
DCKqEv4X0cpc9ZODEtEQ8UTUhxwQZcAZoPiqrIoccCLZBu2E4u3RvGYTF9OPIDVC
hFhtuzoKqJ1AQKjcjASBntPlpuR2JZOaV9QLADWGPSM5Izl/e8Z6ljPb2aK+wJUx
K1Vt/2yAeLC7v/cUHBYyKOvpxqs1H0h1Jbz7x95LBtbfF/UlabtWUx1/Ilg8vSa0
RwI0uGOm7+5Irb0wySY3uXEvqJBkI18stFLDsFOhtidepX4ed74LynqiEVcJI7Ra
O6FPPlEAXw1qKeC9NYTsQsdxALzqw8PITEyTeSqIsBSRvLrVgfA9OvHvQ5YwySOu
PyVB0XsxdIJqPAm4SAXOo+l9CXWMqbDI7qgbS4wHawWQf8rNlZJyKWpc9KlsDScE
1sxdqn2H0BLq2aadF8DmfxmTXZUf/hxRG372tXqcsIDAjMLohakVgnc0SYpElHeE
BOfz2mIw/mOYVrVe5UDzOBBtqtVvlfjLpslGIXtZVOjZebccEbVVb2B5fsyqQycd
CrtSt0VK27gkMCJYnJaNkr5cyR7vxZE2amTUvoQgyC6pB10kGUvTpX61LSPDZqBg
VhPaVLAdv77qxBAD/MWC0zMlaNm8ezVgZpRLGuW2QBtz9CxYXcuHSRLXZgGd+2YR
jvEXEajeLq5uMf6DkbadBak1qPDZ1e31LGVAVu4ukP/VCbZjEtmdiy8znnldedD+
bqiEqTls9OirnYF9UXYG5Z48GWXlOsSouki20c7HCqoXftbW2v+X69jK96SEeFWK
VZ9N0+qjm9lc/ZcL8DahOhv1ub0+30yS8fSfEVVxp7luPE9dhfqVyhk2ggxoXGcP
ICp5LaETaBO7GMmiIqDeQbCSEeA94tc8lfadjvZyWJo8XFal+g3cBq8QLa8X5zVy
ljUoyV7b2+VFvhPM3q9CQRkFKYNiiekUarHmG+elI2Ul9KiJBj1l3cimzFkVuL36
N40fmf5X2iDXQ7u/mCAjeGUD1JPzm4LBA/DFz7wE2PRsE8OAWB1Fh9hWvvXflq0y
q9Ztz4pjrU43VUexsJamnhCt7jJ4dAREW126EHMvE1+Bl4onrCs+fy7gXI8keu3f
Qe/nm5pjRnkiDwnBRq+Gk8Qj04abSasMEclNibMOBiDenqbcbV/PBJKctdbo2ubc
5U8xxDVDuk8Rf+9utvr1yOiD4xikIBYc4WEjf1/rRg5Gl03lG3OxaY7I0W3sdMSK
nmEyRxCkKsyQZ0DXmjW4QTn026CD0q6/DKQ9pqtjEQ9IInJNRPKjjqmFxtJbB3TG
4vglJ6yFQDRoUjUJ8WveQxtp/sk9QdwdpeWoD50QBlNR8wF3/GdlKw/uCn+9lelG
+sXmlvc9g0GC6Tu+26BRUv+VUQNkeSNRd0A8pO95XZbuszk6GPhMvZU/H1quL9kd
XqY8RMsHPPkv85dVFtbzdyo5fVIdsy5TkMK0PCIVf2htnVT0XLng6G7FdhHiTNFs
sRHTgR+ev7SC9IWc7fbv7yQarIzOBCM4BZPWQYq/6v+K0XTgu93IQ39cZRY83eia
v7JpgZxRgK8BeAxTgb6+IBJC//EKL7R9c0m4Dizkseoytb1CJt/9Di5y4rKXHRwd
ASvsIcTB9UKJu55XcT9zWEjmQa8W3zaJizFQ1WB6dMEcWhGVdrC7GdFiyU9eKNAj
z5Vsp2etH3OC/jAbgM4Pja5yCERokBgDKAe5lxuIgrgBgmRCaf262ZaMLRy0eBaz
ndCmZMxiRJ/+cJhnjlWXoweQUBAhROR0M5Bh1txrHy+svKqvuVMyqrED6gNXWBVr
CSyY4j8RbV/cuRlaTFnl7r4OAupZ90ey9lS7BNFwXJ5vgY1rxL5B/6CX4EAL3THL
rIVdAEz8VRNv+r3jlyXxwtrd04fHHVgfx3WK4JmDJdx3m+arkVPpF/huKNTzY+hL
G21hHdrEb91sR5ITKod8F+c8E6NY6fiH05wHQ1KJu/E=
`protect END_PROTECTED
