`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tt/puDji5f9bfjHI9bMiJzkgdkln9ySrqlZIbR/xj/Pm2huJ6wtM9uD/HETD9I8e
gpVQluca6dDUvkmPtTlIM89n3hwHTygb1oTaSn/p8X+yIF4VY2YZV9NDc10n5yx8
oDP7Z1wZvpJhrJUQRP/qQQ5ICzowe7RhaSUMBYvO68/XJeYZw4CXrWzgZvi7NjbC
u5YnACyA6SMG6Hm/vlM7HD5f2CeWIQoRV1ea6ENk2wOZjLiJVlzycBkEODF2fhUQ
nNzG5Ur3/qtxQCEHT6BmtJuS/th1C/rSLNHm+rCQ/9glYD+5z85+rZL/FmIYmtTJ
+E4C/tbcHNC25L6LJd1h9hx5qBA4qEt63qJhu+zfyeehdWIryy8TeWPfQq0Mv4Jg
cQr9IvnxG+0owX2nLxdMGW6fd94Q8JC8n+KleUJ/g9KxvcDX3wBdkZO7AM1QpN9N
bLW+9l6IpYljGB7s5kep/JljS4sTRQd/LORJ4aC0tvkIsap2lvI1kxzMVZG/A5Fr
A9FQ/gqsdgIPHQxe7pK2bD5v+Af52E4DYCHzePzJRv+D/PmLI6b6oZxSRgZWJKrX
E3TT/MVzo2R9MuIlEJMcprNALnaU0ztHe/a1K9MGb3LsgYshuoenNI2lrisk422Q
pjil44Qu9zK3Dc4OAm9W2NfpIChrCPiBcj30JSQJkzOKF4fHV+Nmk5Ey0OanmBYy
CkSqapXAGhF+tgZSvpPl4BokT5hKEVn9bST9wW9IbEP4unxaaUhCNuYvJn4vtwN7
4cEcinBvLm85PyuhJ7b4VLjfVfjwElbvAqkZwiL7btV/qlnbB1a7DGkOJuy0lHoW
31ZABEEilYutUz0kSGPiKZ+p2+ctMcNHSitcPWAD6dp5tQglwQLjNK6sxHUvsqNW
Rgy2Dq2gEKX2ueIYD5a6ihZwyy07bTyCi2gm7d6RiFYSBvhpsDTzRS2z4GPCoWgU
1hqs6WxV3K3Y2/d9H53k8qX3B4ErGYPT+O58moemT7wX4Nlq+vVmuftbOTQ0lwty
iMP3ideU8hNpEBfFDhLE0zrDXVpAwDrZFBNAsRHPIOLJEeXgmf8e69+pDfMhtHQY
SAatw2sBpNj/syAUsAHJNBXcgJsFyonAi/Jy+EeqIZr1fpJ3Sy0eMp8AvHGK7LbG
femUGlDqFsyWcIbCEUX7LAx5QckO6T5s4gTp0o081Sl+AC0nan490u6+3m8lgjgU
MZXFZAlug1aXPSUxoKEUvK6nEWd74bnRUNaxI8W9bxle+TjLNw09MNzxHXvATIs1
psto3miCO499xStqEEyKpuSBMq2VL44XmRDimMAuPCXaDMC1m4icajkqAt+cGEA6
hBrJ6SfSGl+c9fet1vIU7DgLCq3J2TMvOj6oRHgCXPjgA/6FAgvYd1Ef4lxZVeQZ
HPyw03FrDRwDYGHO8c3FDE2gWC99dYOIYNssG6DRFnCp7Ee9w3iejbA+ceebpWbD
qAAf5cGHQ+gc48WQX+La8CTR6JOISDcim+jzlruOfoNf0PbDdlbIBr+PhC+nDTol
fUjQuptWdHaeBA9jpxpYFPTNVd4gWzMYx4tNZDGfn6xJJ6kYAF8MUPMKdaF+WO1G
ukMeYZAseyhp095zqLRypoIR+rl9DN0sBXZIxnEmIZBzVrWkqJFENRlSm3lFG1io
Er8WyAoSX+aJQ6ZwcDO8FMLSS9I3hMm4qeBYYg7sMTcZLyA3iSLFvmJiRavg8K15
70TolRJBblnONPzlSJDbII23ny3nnOf290KYjikEM2Sr5gyMTpI4gwnZFaOl7SZ5
GZrAnz3IPfjgqAPEzf47D5Y/1IOpnWST2wIrhwqgtfR61gK/TlO7S9l9u4bS6psF
v5Wb06IXwmob5f9XUWP2N33yRsnnc+xIgH6lSShltajU6blbyidR7WKQSaavnRxo
Xm9wHnuXNpSDG8GkTO9BlKwdrUX/xYF7ZzD+QBtuIX7pCrsoNhArGc5j34MBbrnj
wDfJPlPgB6J0foSsR+r1xR2poUGAb0vChEIEiANdFZb8AE1FGukNm0ukAf03aQwh
qhCZAOcb0y7rkbBJCi540i/r6S9SEkB8p+jcAyUJJWj9uMId48UnZHgX3g0S2nV6
`protect END_PROTECTED
