`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hs95FASFr2qEvhY/PXXPk4Lr5T+iHLBriRZ5ggnLVoUiCiW6rRTRvArB4vnyxUyy
DjlwbewMzqy3IzsdDp6fTAqsWCuwNwBbaE0XK5w5/xSNLk1d+7WqAwT3A7DTm+8H
cRTXhuVSUjIv6juZ+nJgpc7RV5mQrra3nZFMcKCK5d8H/BAkVQ5f7Lv4REpI57oL
hv8touYgSWsCsLcrSYieyL+IaqzXiuM5++T4ZcfjICtjm7v+mJEhFFJjlGTfcQDG
eI+04vpVfnfc+zIPemzgvYRLW08VXcT88hq0s6uCmrm72Ac93j/1AjptZGGe/uwH
fw/WMein35xnd6GR2o4iU/dZuudsxMbmady7J5j09OMz/n0UzssIsFvNN2fBM6UG
ag2WTp4yL2BJwT4iTYUNCCqjmCRyhD442ajyhmKKem1PwzfP8BYmKPBodMHr1PNF
jPqHc0L/G+x4BHrxT71rUMvfIgl3/aNw0KnA1JC6lg+pHzVpxL7qReTSSq+wtyjO
`protect END_PROTECTED
