`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3Onc45uDPtgfE5ROhdHKKi3wpnYwcYkhrS0SbbZnkTrkmtQ7Ou6VuoC+y7dBiU2
Du4DEuPGIE8grsMjxnLPpIYrF0kBGJe8KO+a7DfNxPLkkRngrq0sQiYSeDJ381aM
/GpnhMmpCPe/EprHyXCEYGD4oAvhPab31S383DweSnHGOcoIz8D+p4laxXiU8M36
LdP1YKGAWZU+SQ+lDOURfnA670j3oZTGpeCG/B2+/RYhW1puvwe4+rR8GCBG886Q
V5/y39EjvhR8RrfPprxuPUqAJQWOwvGxLTtHcHL9Wuqk7/lS4/FysdIzUVJYqwRJ
Fgp1FP1xXohkYqr91H8zDng/km8MYaGeZ8B3xOAKZVVtrRARQVm5ZG4GBAyF5ji2
7/6AyhXw5RtvMr+clFNV6PrRCTBAPImwUA+36gbrmLEnaaUp5gA0phZxQhFKh7HY
lxo/gtnzqhidtStjWxI4msIOKPYb97yAbiNdWPGafQthGR6k8o7mLM4XNTX/JXeF
MBXkVY0ypW1npBV0SAYAlNfMm/tGCYN/hBmKcBgbRaSuCl8LSKdbrV629NyY5x7X
aYiUXOcz+MaFa/ijUxWAIhfMr0IqiiwGfk/s7po/wEXxRSpINcoxAtkBZeSxrfve
etEpoTaq9RermtSWY6JClEn3hPw6SUT7VMAYdEVgz34E3XG82+M4OfBYhLUlAGjz
Cm/z4cSymyxQ0/hNRDK2rp31k41fAF8fmg2Y7Piwm4cy9g5NEl/3WxzI2b/1Rbdb
vlm3gLkVpHKGQqT/BXXjNRpMxjiVHp8sWflP6PUjGyGjb/4EuvS1rki0eB5tqx2z
vtmOu9OvVhcOl+1PFaIaAkjEw9KTAeTK938fyNyCEjC6z+NiLOHJKVe0VVdml89A
SiondVwzNH53GSBa6xUNt2APYC9qGXgBxZVVPd3Uw/cIt2NAxwXQRdM8VHeLasO2
RkVOCpiKK6EB721mtHoDwAaXUJ2PTAL19xYyYQaZ/Uis5lPok7MrLa6361m1SW2M
ZnAwNTcKhPhy/O90ZkCW1/JVe/mVg9py7AyeNKHkiCf+KSJDOs77P7eK4N3fmLX4
rH56z4j0miirjMqN9QLN1b3bAk1JzuzwgRkTfjK63L6na81+hIcPqZ9R5GcyCEis
PZq/fPB3y7cySTIfcyvfS6vpexJLKzgN9EcZoCzKFTOqam0q/4Cyn3OfQUJe4sT/
g9DR7vztzumVU/7FhY/jweAVX0wJckNrhQoKQWtitbSIr3ZFX0wAM2o2mYmbpxur
xNJ8Hjd8ForQ5tl/Eoynn8M8iu/Lt4xrqeDZvdNDbjUN1kBiLMAzwWq0r1JtUIud
OgUO58jlDuzt1/kB5UsPvYarsVDf+225g7E9Kqgkw/4/r+k5vQGp8I8InBC8VM4h
EWbeOUXAhBid80F2I3P/Zv0Hy09NRdq9J9OuH6F1fD8Ourh1HjZ7QIqQPU8/CObZ
wlHUqAMwuFepm7sNypFt29PLGBBjyiRwPK3+eBce29ydaaDE+z05dgDYKNpkwMqy
74cFkg6mgNJjQ69IXdyJRS9D+fumsDQqah4bbYStR+37oEbggEz0A/zs3qWRlJTj
kkV1bhmMy2EQZ9josPGDxxDUob2joFAAMfxxxsda8bcse/t6cVsdVFha1F/ZBXXg
YYMPif3OaeQ8jlelfO+5FBeTrixIK6NuBd07hmIncaTtGrp1dax8Nem9ROq3TgAN
2tqigCfyG0mI9GX2a7Nh5/YbErmmWaK5+mhlj7doSnZpHqISxNv4hX32xttPQNgV
uHurH2qD6TtPPcjsehS0Qq1Gh0fNh/mq14nXYEB/+6ruThNhb4JZpC+nAbrz2lyS
afGIfOiTPIoST13WABsAREXT34/6InYFTTNjVkppHIvHNlzAD3tliLvtv76kXwIP
sYFlHuHGnt4rMynx1QCGDiMqj+byP+61CfNJlaQzUdubxeyiSX2PyN38Gsyr4xMo
v0RuqgIHFB+NEBuHnrwW+ZYXAdyIbpPZ2F635rQBd4mBEKF3q9l0uY6fQzK8qhOZ
T6BsfgZUwySR+ZE7a4spchPnwNjJHEtS7/ppOcdckSF8lyDUpaKDXIpswdiUn1iw
47MvXvkusAYOsBj4CCpgKsMFVOYo3sqR8A70JHUNaTXy/m03Pm8EDtsK8BHQ7L9p
5ELNzZIj4/MvoRg7UZfHQCvExnb0wO8Cce4kUPuNKRk=
`protect END_PROTECTED
