`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gr+6AFPNuqTEW0ZCFCGLsdzFGpNOaqmCMwat8GrFYrik5OIv9vjCE1QlCtRR1rwt
EZEAgNCpyXiYJDGBikNcydYu2OG88m4S0XcNfkfex/420rFSzGgR5lj9NNjRRHaO
mlaNca72307EvMLh7qtbK4i2b2wYG+2Yfb0XCPUG0GBnkQUZ8/y6+mNjGHYUe1go
wU9VbYDm2EMN/v2Uz0Wx+XkZurKBJWfNOjtHgnBhoSe9j9i05bGERxzyE86X93Ko
2XG4i9NLbzf68AAnPEODa7vPF9tFlgFpRubAyMYuPGiZnmWvtJ3l3RYnteCaKha5
Cr+QqdUHemfgFiZYjTvaV4GragDnyJLTrPenmmtpq+z3JBYvtXlJLGa1IPcnB+sG
xFCvul3DC24KFLAStKLNi5mq6x7Yw3348654PqRxMq+br1ywFjywuZ28X+sujwp2
qZVFxc1zRybO9zRE1lcfMCsNU+haxT+BKHCboYJLKrpXsFcX/tmFShWtSZOMGTqy
bkQU864h9sLY4WQYe6U5dhBJqzI27dJdb2YSE9RN1qfU2o/MXOlrvd3J/xt/dNVL
C8ExZgsaBXVb8phAu3WLgLxqgGr3ttGPqCGUoMToLwA3GW/9+CrA2bXWJ2Pd6xID
EIDUuzTIZrg3lZ8KL+l3bA==
`protect END_PROTECTED
