`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9gyAkwHGrqxj11BoFGJ1G3BlRj5yCWXL5K8LTTJrf7TxZQj6fQLUnwg+ovfoGmx
Xv0q6PNO/m9hBzbVpQ/1kSOaDVXhSC1tzm35umZrfuHKuR3jrkXTLyfkGtjUkO/G
tVzs2Hir7q2gKwZaS7bZbPGoz5Lauw866zlpgWT3fBDp0UFeJa3lk/THt/51qJ1U
63RsHR90iSGDJYTRdz6qmW/gc+2GMw/VtcaHl53mCNlJqomHFH10pPCe48Ir9AxE
XAa56PsyvenFsp5l9Mne3i+bVOrH2CfNWUBCDYI8UWvAWqIuFN4uJCAyunCMSWuz
q9Vlx/3gvR2LmKz9uWzV3kjqZn2rramYt2019jyWiXYP+e0CtsTsOizDVBYk7FKN
BHViYHakLqcRWr8wPWyCfL74nDzFi8Fvui0Hwvj1dMfpK6dh6dKJ1aigM+0utpS9
+R8Nlfn7+4z9IWfNd9sE0w==
`protect END_PROTECTED
