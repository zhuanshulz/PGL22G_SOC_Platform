`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pr6OhOsuyfAHGg/XkeHergjl3bN+KAMr+QAekN94osZraxWOrnWUZ371GE3uePjr
XeKSnI0lfHtVxRRJg2wyBrPbVvNQQKNEaujSOBVintwQR23aLd4gv6p/EBjzOb7J
kGjHAjC8+uUKKJuE6rJ95twz9ZH2c9X42YEtfGRewo3c6AI2aVnthUq3mZ++h55U
Pu6xst68rEvYYTW8k8mh4GWcoxzOMc4tfwVTDVWHmKkElVQ36zOt0Sx0ATHwR6xJ
ao8vkKovoqXMeCs+1zm/8A==
`protect END_PROTECTED
