`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFuEHCEYDNkRwHYIyKYG/8iBrL60K21BYA+EIFTol+DSrujQvg2HovxKq5rqU1Wv
JHu19Ysc8EwDfoJ8eSZ2f8/XJ/rslzKFvhC8NK91siQOjmaAZf0AWklGThsDdat4
a43ls2bIXvDGCdjQ3HN5m8Wv1lwvxBOCafLjFMX5BnBl3sgp0HJYOaGqB/BlO0xJ
/ffVDQwynYSqtWD3e7fAkvF/AwA4F7RJk3r5/hq3M6eyvjigpJ0370GnmWWMPH1T
wlJVSONdmuZbdpv8c7AxtaJqtzCwpx95fjK7THUQzhdbToJO7JwLGkUS0VsNn0YM
2hHEig5syyd89GZ/fjlqI2NVOUR61aedKr8BgIj1LY1bi7A3Rx6fOzSvtVkufGfV
nCcrw9zm3WL5AgRBXpxk7m+nagbhRtulrkdySjI3/s+c45ERd6ezYpAFtSqoztaM
WKLopvyBvloHwx4OD4HSZnOcjtUkOE8UECivf8on9vKmIetobTnDvOinsRgZSz93
lWBnGBgLw7dHcvrK4BzqJa/X/Rx5tlLH/e4WO2XyEW3ylfev1j+Zei4jk5an/uEp
O/QOcqjjhVrQPzEbcwfIg2Fd2Ik9HfvCvMM1Pc7h7EUZHdOWbUrar8tqRIbfmAgi
xuDbvW+kJxkB1S51xPrfaAGqq5TxfJdkWtetvwfv8MNroA+Wj+aHwHaUQccqQvjM
hxJW40ruhIdu5OQClxi6v+su3oFPPIxR49GlMTjcL5RBd8rz00Bh2FPNI1mN2HpR
hCK07CAN0cOKCpbZ4w19EmnUMwONqcc3cMRGnxiVyU5dvDfQfaTP7ZUuUZ6PPnbM
78mSgAtL5SkV6jACUC+Grl19eu8/lDE9OWKbspq9jRcD6/JFVxHhzxcFdZtq2UMk
/YSfxh0yzXCRVl6NLN2LCUnI5JdvHHqN4W4pPh/fj9mQ/+OuG/jAF4Oe6oIrLx5T
//l3J+1FhhrnWcBdNK6t8CWxG8MrYmkyxItDb5jyzWbFxFgPJP6sEfBauRbbWvM8
w5kbBKGbJwrQzSDPeMBpsPOdlLAuzG6YczXcoPK7vhdZgSAZDqCYbFx5j3jbSaRZ
+fry27jgpo40cpxjzrMVKm2BWa3HhCl20HcoWXDO6i38l8NzaCrcE/0fwzG2ZhK+
7nD5o7qQ9uYW6g9kWVpidcqZsNltSyze1NL+K27iXDJGHytnuP4yCHJiFaJoRogQ
DsfMikazdzm9iWn4DoA+CliUByHFAbILOQo3XACs4p0ebV7YUmorlZDFzD0JASY8
oOJVnCW1E54khh59ActiedITKMwy20bvy5UD943WHXV/oig7bshXK+qjAWJ4fRkm
XOfkHUvhGrqpLb/45zjiDUAte+UgVaJDprZoTtWH0FhTvnGHUSzbZUz71ox/5uQU
YdPLfAhOzRQMoEiiwl1SXpf0BKD92On061gM4No5Xyk0SMEuRXdKXBh4Y9kd7HUP
sb9xvZMBq75spuNnfgcr43lbKCkBjXspnQ2wFh37v95OteEZXX8yD0zCpiq0sxy6
oKz/p2Q38LQqan3SmM+hA0EVg3eENSfxxlyP37gmTitXtycnYuzR8Ib2Mngjc03N
6TlOzoKNkg/eDcO1mLW+gaG9rNo/G2BLBqYsA9oUXYPHwPoo5G1JJ0aAHqkYVPsu
eF8zv7JVd+1cqaaaHy4KT+quYJ0+nPQXV908DmS9gb6pw5I5qL6uQ5f8VvRXCVRL
eo5wGkYodQQElLJiw6LjDmhIE+6hfKpl0VmOPs9jZMTFqv6E99yzxU93poVPkRbl
X+sfwetgXyO5ijnJqE97Go+bXUl19ohA+ScG8E5MI8WvqzEnKAHGvqssrkCg+JhZ
xQUXQPz1Yjj0Jty+04t+5GEELm9grU4PtvWQoV+gf26OtyG+9+A2GypGRsigT2tq
ne5NTOUPCzD1MLMiMg7NEccHsTUzSEe/kS55mnxEiKwtt0ko1vRzWHvm9S+LeWn5
jW+xo02bd4ECckGzJXWUCT85B9sdFrXn43N4mZyyFZ2/mAFaaPOCMASInw9VyrXb
9I3ypkuZSx6Vejxfa/pISFqpl0w5Mgk66c08rIfilavb6h68cfpux+/IcoyFYu5X
uR7iMYGNwR/JBJcMkOTWfCpY9rYsro/1pVBtdKPXUBE/V+E6iE4o7bW6pMpCsX51
RjSJq6DiJL8YsvnsaWz8wtR05K0zFfkE3BK7YnAFoIDTdscouFa2n6oluw+CMl0H
15EjwxvA1LdJRU1eu7VPuf7TOgAVmOwddO8vOCc/R723HFSU+2hb42kLaN9a1sa6
bKRLDfib1jth4fho8etjOgmCZLxhHzDPIG78IOEH1hQJZIt5hti9qGILuNsT9E5u
g/tPLc/zqMG52qBtTRvrZYzOmOcSosM5dmIlOLzeVjUX1TYZWYznNRw7S2TmnAVr
+0SY1KrjrJmqaMRVvSZz205qOsB/QqpRhJ7dFepvyRQflU1ZkZExnyd8Jes9VRx1
ZTXXYCfiXvUzGCkjVdH1TMXZBKoEZQCWK2X43thO1KC/fG1Vp8PlTjtUuCY/V/J3
Z8++4XWTKdh5dmly+AmnTxcaMQyqL1ETKPbIRjzohxN9K1ARds2MGdHMj1dQ9gdb
tNY7CcQChMHVCrfnKkg/FXPL480+nsH1WVsa1y8tqUhUynNatX8vNg87L4rZR/P1
CJbxrMFsOcKlogFLlnl3EP0RgDONcunNDMlUQzG/NQJbYAjey7wssbFTJk8go4hz
8P76ZaA4Ik7CfzNmN2Pwj8aO2Nu+4LAl4kwh5mSBYEKAKBjBsD5arjcTvG747r6r
oRz5puY9TShIPP/7t5vzOxiw+6MmwaD/8Q1EqNzUi+UDByCX1HPUOTNK6eBLUgCY
kyrIsq8n7Og/z0WVDksnlRiXiTAcYHorOurP97eqx741knU3713RFpUae/TyLjUU
45KNkDsvHClZ1p6te64wR3DzgnSfPglmGJkcexQ5vr0CB8IOaGdSBKwYjv8rS1nV
UhJWgKanhTa2uSH8xka5v8hXaHy2+NdNJjKUoylQRjSnOHPPdhZLw5udNRtXVAyg
tQHqFgrv+DB8GOLNELIByfdXxklv75SmgZwvRBWVyF7bAXQup5BCDkpvq20HaDq0
b4jdi4ESu60IFN0Nr9q6RQ2X3P7FVV+vbqflzqVLqXMKi4doIpmaBr08eKoB4AHw
9z8rWQ7ISwM9qjyD5BQxrNHqXU6DXucWjTHTwaHinGOvpl+YsdGIvOeTV8X6R751
Qe7TyfIa3aU2bpljDU4lPXbs9XO1wJGa+OEfCL3FboK2WeohXrY3xP6lvyaMKL9J
0Us+TUNy4K/pHxbuHVf+KgdpjKMoHJXIFBCGRxYmznt4SZQ++35DXDbAXZQn71ri
juAy5HgKZqy/s1L7f9AFSK4bOw7Gwa4LK+MTKpM4ld001HQjwAAuEc4tDUFocJt8
UpCjjcZdOcTWiuytaeLzbiHtuf3oULHNp4Vq0Duk2cO32klFFAQrFaWAHeM8JXmQ
vNna7NeeRYFtF5sYEOFdA7xpcqetwpHu6XEVBtQOHMyXRhVU4MxdOFFW8qu4S2cq
9p4fj8tadIlIgqPKwhEyQ1iutNTNs33ZMaj307JfZytUt/NP8fHUVzGFFrb2RXO1
fKVgb+jUo8bbXDdf9o+mYsuVRgwNQm/oer3ojBElYCYMRqiozzq7z4MbpuLPds8w
cRlrta9gksr/5W37wtgjsWUAgHNjJCuYDL9P6zqMfoxfaWabYW5AxZgG7Bg5Gm+b
yEa8Ne8UEJ6KoJuQgA5HiokhvpD+QRtJesqByRLfRFozxYSMfzdYrriUNvG3yJUp
ypuPZTryK+xzCtKrHD63fuwMlFen409Z6h8UxHCi734tpl6//1/XZ9VOGIth3nyN
lHo1URsW8z+hYCuirujXCZqJrFu92Oo/Ru0cbhxsS2swnq85ne+M1R+f3hrXXkBz
POkW1cn2LhAiTUuQ/fyUuYbvVEJE0YOAqAyzQTXYHy1NSfHALJlZ8O19Apt1HsCB
8BRzKVU/E7X1kTK1e59Wv8oVIzVMdhhADLea8mZf8eNNuRNt4qAQm7wQ76etLxtb
4PQDci+uUtd10rGiw9s4r5Qx6lhZkRATG00PdI3xihthcvDDb4+aBRWo5weezKhg
TIH5XBBr7PoAzYt8jTousvxo0NL+ZoOXX8RKvV8jEpQTlNmipOeH+XpPdWzEOKmu
3tEXLT6kSolTxjmIJAQkIQoKdnLDXM3d4rtc4QKjx7fvzJykDntXWnUt+Jdv6nth
DUaMBTDugI9UejJNR313R+LkjC9L05/MQZIaSO6sNYo+gDjRgh6J7sqBQVYZUP5g
0AoF7M4yfQI5CApw4ChWZ0TkR4RO4WoEIMLFWhX/KVv80oKABeRNyLA/ofU4/qSe
I/3jNruPNwdqJyudO9X20khGrufqVvg4QCE3R/AS901RmLlbc1vqKMH3AW64kXWt
Tqr8AU27AERN3d4UpQ/FbQSvKpHSCvfYK0i3m407jWKhbkJQZVWgVsExBaKyg/Li
pEctUM39Uo1JfVBILxeKH5yrgVlvzZYPEb1rV+mu0yTXDJRgQtTlbut44gIMLMQB
gEEFx0ADEUED/tNSB8V1v5jqrYSTt4P/ykPUV4fgyKmoE7zxVKQD+WA0zOF8pv7T
hES7MHc/dnI2eXLPcDF6p4xZMR9jhb4ZfByMD0NjEw1C4DaDdCa5ygy5eaZKtTL3
fyBzljsJeCxkFR8a8Rc1iw2hYcB1nXYhvzI8nFVGE4dURr6e3mPNnvToBenEsZRs
UFtAJ/E0wQzvRIaOBLV7feMUPYbwGqwDK4/fYejURRejz/SPeNdbdGn2ZEueTEbw
XG/LMZK/+Sr+/q/Wnc+Bj8tVCAFZOIVrZf93SbESCosjsL6xxLv0eu2Wg1fP00wG
vYzJ4wq37n02dh7+2WtKZBq9V6mdHuAZNrlPZuVQCkLpEDp8SLAo92ldlwIRLb0V
NDmOHEakJwwRHrEjs2yYIgb/CwA45sqoqjPVbMJw8MY8brjQ3/OP8watk+pjRLux
g6IJvM/2KbMYxuzOXsuVulX6BCeLDoe/jLfEvc5TXXcab2jui73ne2KNRUutIDxf
tA2/o/pyp4xRx6fTVLNTq7/NUr5f6uMRDt/CwY6ndkPzYNDeb6V7Lu1fn/8sFZit
Pdq1QZ+kg0Q9Qprrifm8HSMT/7ofxlJ8qLJqpm4ixfVsJDT3YO+NN9Vxk3YxpV6V
AS935M09yZHsqpcdD76HZfTMh+aweqPCUqHkkx7imufFh17VWfe2bR/XkFtEt+ap
59GlMSRGi/T+XukCA+v5Jpmsa8bOVHy0bjSagYs7AkCaLwP1rVNT3mDS18rVl32O
KPP+oRAzzvd5+rv10BUpxkR6NztLVcbT+yLzrATae2chLoExSMdHWN5L7ITOuVnw
2BPXrp48ZwXmh055m81lulYx4IhX+LDeYGb93ehu4JJvyVFmz+aIo8cUSHllw/ii
kE4iYjVHin+CQE9R+VeMAItDvkfB6VDgNUB3aMv31EQmo7kdoSRN5T+aTlG411s0
TeIundUQBcmT5EEa8+Ta1ufrk29zoi8mxnQuAxX9BZSVQ1+q8gZC3crk0BC1eZFk
nVj0we1tn2Mc9pLseJsonFKBPBwPNFziDFVzxFSE6wz5Fw+1MdeKJxbml9ZVBZnS
mk38oss88FRTEVoBpVm9Xa32BeahmRF5g/+WTJBTh5SVG+ARqedrZFP8OymeYO5V
f4zkinKr/ztLtZJspXCVFf8G4UdoaENkgu/W8WdDJyw6jmAiopLhTAxuL6kaXw2z
+Ij1p5ahLELfDRIY8Qgefr3KuC9AMZtz1Qeov4DdM0UN/kiUZMzXhZVP9WY1iV7d
70PMVpgYyGPjDGZOOnf5gIG0uKYbAAax54Ed6bA5uqPq3/aHqYnZf00HShKrSQcP
zAeDzt03OF2mNhDBuGmVNtXyA3FNAy5DbsJpylow9j1xaL4Lwl6uSVaRbkCcI4ch
RjB4q1Oxe0IGwkVe922c+K9Ivz3sH23nheqqYEFrBLnHhxMS7wwrR7EmdMOlUqVT
1bRb7x1P5vWZrEAtE1fxMRZXXANe6XjUqQNNQ8fuL9zrxpvX9xDaT/jUIXoXAzOI
yjzgcjFPNtHR9L2BMu+r/Opib0ADlIfrGiAxmvLWbl7N3qXlSvoYwDMTu0n6grDa
MspOXZL9SJZn1CeVBvfZ3SyAnYcdH/jte1Mdb9bpQ/Lw7aoUAS+y8PhiOC8a17OW
RKk6O9/0CS0cDYS2/fQ0MnLNrZk51h+w22QKN+fsIwbaosNnofOg45L0VBxWd98h
09i3jpFvAH2TrFNWGrdmUJAEwgM4/C2Oejg0uAuSayJ7w8wMRvg4cgIUR0FjP+Ti
KeKFnu2FUfkfAx6UR/XFLYsMgiUGYV6uENR5HIC666VrGBSbf9XMNJIYoYrQhVca
XtxENomxNspEJk7Ie0d0pKML90r/tNRrieB3JiGuOYwOZdhmg8l/awNapxDgl8eL
+vYyjr092DH/ye+Cwj9vCjIzLCPxvpIQ78vHgqW0FvjD98M9xZrwh0aKCP5h01qo
Dc8jFmSAJ26CieuWWG9G3n2xH1i8p0mm+We/BBiQQ9yXamAod7/Ps7BLF3wsVX49
AQlx91p7FPCzMDVkEg317WnJodX7owSKNUdcaEElHjDE6ji32IXqEpEeJqSLbuMu
eiJehDGs8vx6agqSlb3KlvTbDYzK0AoQM7f/RE8L5y9KtkTC68OOWzWH0nvzSYrc
gDd8WiIKuvtiSl5QVSDZ6Csvp1toYptzWyF5qKgiXToQk33UZK0tI0+t0yC9YNsl
KtHCmC8fulZAlc+wrcHqkZ/4J11Wd0g48r6xwo9BSV8lHBk/NYxH7zTrdX4WgYHJ
Sk6o1RjA7RuTw67hTx7eeiBzVH+IwBztmpTz7TYBDWEFnmAs7Smchbv5UBGtlgCk
h2SFevbYtzSdcUrgvB+vPnEDcg6jejjWeCKygQ9HJDKDorYz8HoGv7si5NTREx7K
ffrjhYR0zznDJEpIIxRrfvEc7tUErjDDMr7M0AqeSTYcFay+N8+PyGzP8eopHd1j
LAEB1qV9LSfXdwJqVpmGb5BUV6jpTrHAlKHO4cbGko3j26T1f3jXmefPNrnUQHkI
UL4PuNia1R/5uFA9FVzLAPgvRGKrnmKw0mk+uQegPVKrMF8qnMEWv3l755k39IYy
4r0AvB4TgrfI4lnGG4/f12y/bHCyJWKIYK8lSq8O2qXKxlcZo1Ggf6+gRCMC7/mF
CZgaR4jnESQB8y2uBXnnKC528JLZZv8FJ9ZbV6wznPZQcyyuzaOmdfb6jCkmQL9w
Qm5+yUPxQSHay0zvp+WKydPjz9bLcCJyt3KLrl4KQcLsR2Tez1wO468u4pCKVFKc
sdj8b01fX+CGTsMNp29tT+M0n3kp6O/Lg5cxqQz148TPwyDTxc3bleVDdLxTV9+p
4QdPsiVXxNF3GAaKSCrN4MbKJPNoXaag5aGsmACLarV2Pq1MymH9SKsWRvNkyc7d
3J0ytjsEGSdhYKkGaxETGnYoaF8em9ku+UeTMzgjJC7AgxuKD2EOy2i5eqxvZ+Z+
IhtI/DevKgmklKqwkVHXoWXZ/rjFkQ+SRQ/kduLL0Y3YUamMwEGM01nQc98ueh+J
noQR5wNCjHUYZAHmIT1Etywy7qhwgK3fW7h//RamfRF05PoXoYH0VoHji6BLDZ/7
r4W69eKaUqOvyfqKC5aF9RFpUON8GI+Dw/u/ZyLBojZ+cm60Cb6DvSYBEzrGuvZD
9ATugNsSRhEPqCnSKZjOO+VQhd/lXyqRpf9xOxcznhSE2+QYoyJZsG5wFZ8XhoR9
3VwDHkHO/D2SN39KUqABqMwnf8BwAnTFRSlhiSU9xeRnhrtmIC/L8Hq9xiMCmxfQ
eYwCB8+P99E8/zQ2IsXQbBsGwBugEk0USh9VhIMClrqo6+rkdZL+Ey6k3ssa3Psm
Gro4nIeWpHNMRtdN6LVF/QHo/Lnt8fl8PP7s+GrgMcXfqE4wcf8dgrpIMJZdBaKh
ME+oA4IpqZaZM2L+Sud5A6P4HaI1jyNTrMfeDKXwoPYIjavlUZTToOFPOyvmDWpY
xzoZaZN3sMxTAf2FxvyFanIccQDWmuVxbieoIYhKXDdY0Uqh7LYEJMGYv9VuPyZD
b+4n7bbSYtg/mq0oCqWRpxoyzE6nsbyLK/4cSdnL2AkdJtinhdeAjX9Slbzg8ULe
knk8j8mr87zF5PpUi9p7oRpkb/hmJwrBWMG23acLdBvuLmh/3sM0hErlMbW2N599
Q6DiFkhcGv+h3MbovJl+847/YxfYDSyRkWP1ePhry7nKopBusrtRLSKhJdOpxVcq
q05wUg7kt5XrWJLd3/H+EPyee/8tgeXcCzOh6v3r1Q9aoTO9SZtQ76heyq7UpWvZ
xmrVYqeun7233RdCF1BJ1h/XXvaNIU3FI5CUsNpa0ItA68W0gxFhe/sMWu2Zdysx
MMmpXHJ5o4FcCkpkKsvI0a1ft+s1T9vhh3/KvLTuJo4G4ouAt1UHZ8rW8u0Y3tC7
4eqsbr4Qoom0vpdHEbL+/WllA2fp/nB1PF9cNmFAx9tez+IP5S/SnJB34emW/lL3
bFZVrq8tQ0CVUdr5i31O7uBIEx2H0VG0hVjBsQqz9n7CirwQrMr2RjSVM7l561FR
D6siTc51wkG8rOH/7qlYXRRO2AqKmTMxiH8UIiSD9uQC1H2ZdUxNL5oGNFPU/+1m
m2KUZDyOhcXzxTfKeyaf308bzYD8ABntCvCe6issOPoD3BE6nQzRhpgaO4vgNM0V
CSBaxvzvVd5C5DwpRd2Mshdrg1E7pDk2b1F0caRsK4YduDGkvlejEiukCsjINv2I
JjvkDkynt/IGqI9qB+YlUx87kgms8G5NVtGNyjDUOiA7ivu2CM2OKq9ddbcuFINp
KKBBfHYvmN0HkbQ183osT4w1EMTeESA8iMtOFKfBudRWIDwRyGbzRK/9f5bPlv2X
fAaW5MtwGTjjtWLro3Asnxd+nGWgye4ztA2Fivbk7JMhnc4NZZB1fv5NhkZEohaE
TR0kWKghTlH2dtGjN9zg1aCVQsetOZnwD1gx5vhFXnJ0PF7ka1qA9Ha+/X9dvueQ
JtDYM+mAjeTGqk6zNEBnx5g9JU9cdGUtLuohO7Y79hMdL/a7jeGJ8mEuG1ruVvVC
rn73SQtULPFgRtKvZuDN8TndwAgKtvL7gM6yv8GyBJ1s5NJADx7KwATXJM7uHT0C
ZJACn7yLpx71XWVjj5Y1Qb5SC7Rc60HXhFJyospHxVStxY0a6x3tEsDlEZL9ncNV
dHftBWao/q6HGfYGobAa12jk3vM8Xc63gfx0aVrFXDvueOO0PAbowV4u09jNWKRc
en6VcoyQLtvx22yq/Y+dSwLxIIa51lpRwEkr3UhI7UK880vqpwOtJIQD4egXRmMb
Kl09ZcRWw8OUzIMTswB3P9/57QgLpB3xElGkvQJ52y7h5zqxca5z19VkUwiotfp7
t96t6RD1HNic9YB7BoCOax4CqMUZnqDh17tLt/E8JCcZZs9Xm/gMn0oQy9m/HwkL
aJla9hevZbcttHopV/WpijE6taHNUQ/6e6rYj6uY2l2vvtL4Y216Zhtg2IZ0l8d1
JAWi6x0yfcFHvftA1NkEM8XOwtLSqgj5p7a28ujYXU4rjJKiuTSy1rK77+vGo0Bh
/ieTwdLrKsttr/yCsC1SEpATvBlzV0F0ITvPxMMXxNGZmbRy5nPi7KQ8WyREYOcN
MQO4WzcSDFYUlUwnOt+GkGKdE+IjITd4pWP5SgrBHEdUyhWgaNkvPqQOFqsshTA1
94tZyKd+qBcVzN70IqWqkYBrLvYuT5VAsRA7Ny52YY75hzmZLAQy5Omz6rgB5H+v
7Q+Nan+QfkLfa0CZUlWIein4evODvWE+kZuNLIhOuEG6AtHIT62Uy5+a+SzcwWD+
bCB/32aXHg1VZy+iOTgk5QPT/Xd0CyCD7L9G7LCdkA9dAfeAjkBuFuUs+ndty33f
oq1EEYNByOrhuwUyulsRaqJ8Bru8oPJrZcD0qkTffzAxm6m23qCvRCSfU3QBhM1+
dQCZMoUDbDHGQoIiz+et457+G29Bd+Z+PCVROaX7Ry0Do1wDPsaeHu6m621jrWk/
4+C/ztZGchJArQgMLYNzeNBf/PL/NDLwMYsR0zx02K+0fY0w4h52aE8g+wNqiVb7
t3PtBsQVC5EJ2etSe2fn/Am+18XcsTuOEFHuhXqB/cv4PNfFSHMmtBMfDhIWgg0w
TwQVvZ1XoJCV8UC+Qe+gv48gavm4T/yxG3BZsQvRzoMkX2XVfks+IT6cDomIltoR
P8YxJLTYmNL/wpXpxDq18zQQ6jKx+s8kIkZh0pKPbUMmfIZkTkDSJE2ga/mjqjK4
ibLQPj0EqGKMvXn6HnapQk0x2cve613gKqvFJgBAggUVAbIdf1AhllAQt9Aj2GST
oFmMJuS5EK/eNqBkpfFgg+YLjEt3i8KtrP0Y8dHUEjDfAQBfouzjbtJMirmkalMW
lffurKoRuyBZnJrqKpgEGZ1jzWv60WMryNmh4u27cZPKu7dhuzoxh/NRXFgQQ9wZ
D/En4xdYYdNa3CLnxG3Z/572477NPz4LTbQky3ws2suHufgA2CqEUsBK3vTiZvjk
i7k6wQDxZ71UJ6XXwMkEDk8hFe0EJEq/+AJkVxM0bujWtxGNLY0SgkyVhXjCWDUd
UjnEjEgbWJflbciaE0b4tYZwt/nKjtiiflBzYo6YwiBQbTd0OeMVAhcnaR/2jdWL
WseI1Zb7KPGnqnKXnX/ag6HE4VW9hl7AAuiupWzF/Q3Q86HfO+3kPZMDiR90JHn0
lFGa0ZlO8L/2HYhq04OWWOikOkGPNfycaqOcH8+u9ni39ASllYD0y65QoT0AlTFS
mDxkXmNEE7M1zP+azacsypvm/u0243gwHnKDyCSCpHLFEtufaGy0TQ7FFjklcP2J
s2Qc3RNQji8axFRQJ+YxgbmkWcgOGLJt3hn8QXH0yJpZeQItRQXKP0SSPUp047G+
Ahdwh1gPICaF+/vn/bqAJ9pCyKMITU+6txpjNhHGFvySzc9eaTcC4SkhFUwD/LUZ
Inl5RoZca75Qhvzee1jp+YyyXPy+b5F6yqJqA5p17+nw8k64YAnE0M/iqntmqtam
tcN/9BcirBdZV/9+zRC+x7/4WMdixiENSw/2Dak6JQS/vt+kOR4HXX+IIci9fE9I
GAOG1niZyk8s4+lpkFY6dNiTrJRi2Ihdf2/f8cMP/QW7T6ekJegPv084CmiNvNWz
rBLoXvgkfOnKL2BkkIlY45xpOdtFEPNU9J/uO4vYvd8DjNHWeEk2uOnbXY0dSdHo
nCv9AN4VCTgu4edxJrKsfZeqwdijIqaFddA1dGyTjrIh2bbsvhQU3s9e6FL+q4MJ
AhzzH2vyQte4R2Hd0uD/P+DBRH+CMeN8lSYtIpFaG/1IJylkoJLej0LClik2A8gE
WTT7ChijHbqWi0nl/WBAPNKcuVVv3IpTxuDz9tAXF1D52Y0NljNRfQn5J9yadf7z
0bHt2I7VzNEKQ/wOFWA4LrHPuYg/RJpHzYcgTCWZTz5T+OrWF+o49WmVQx87bKfF
kpvgAZ0zULthJlfUSqa9BPA9oaF4qZTCELCTp7iKqshmClAB5tK7mtcUCLo8fehc
6QLbtilZhm4WGTRRRr5+su1YKkKi2TjbW6PNSC481Bb0OGckYtyts6IGpaFBEHKK
xkXAdr6Yt039FspAzrDrmekYyUPMpSnIS/tIe8fJmxJw6t+D1SRjC9t7ij+JQna6
xA0qveLsuY5qfDMHuIPIzUVkPfxUB2FoQ4krQy7WB4p0uDDSEuDHDk/qQCgn/K5+
UYuJk5bHOcL7xTV9aVXYlEuWnFEcM4JUVytHLN/bhPZl9C1EDLSSOC7pS3w7hdvv
Wz7g4co9zLoE1FwgaCxZfao1BMZa4wqbgdmmMGTRStSS5TEKWH3MET11tIzCRde7
SKwhy62oowmFYeRvhWjvnlXP87xPrntvZaNpEoa0IrOshC/cQO6OJcQ53IFThNAb
OCl9lyOzqV2hREU/HiKtqlgpfNSJtEhDukZQJPZKLFMp0x/MzDpeQdX0CCwgn8f0
wWhANDZ5Gcr1HQbZ41eA+pLNNcdW+jndEtHKQ9CpsbjECb7sy9obg28MsKP4xxjY
z4auOEewRHQ02pQ0ITUxrsT1l515NXIyd+rXGw70lPpT6ww+YkXLjGhvpyLVVnz9
kTcZS2WSCYhVvYi5J4vgLAMSjp19PZ0SqduZFF9oFf2TV+Os1U0BpLoKixkR39Fn
sNs5RiellOh7SkHxROYx359rrpZemY++kd9QMQ7+o6oihk0/pXYosk5ua7N5sIq6
q3P1AnmQXGye1csPBFLBeM/PlCBHUXvLj7b6qm129Q2wa2tE//PHj1Q+wrtT8t+G
HpaJfbFjmAeq6mQDSPDs0AQy2lGpKawo3YWnNyAsiNL2IxOAFXWBajent8wHvVn4
iba/n6tXgUckleyaCys2NPhrbu9LPVfydzfcyVQqUaujPvESWS2QvvZMCmmN4mSl
p7pjSZ/fLaxNBVOy2YMXOL1ac8U9tcCihjmLSi4YKWlUeSa5eVmB5KMddxbxqmBC
DXzfWjXaAevEctjvnTORp3xto/mmBJxk2y9U4MOM1R8fsRMU+Hcs3t1ENn2aWTIb
1sPvxwHJB2w3U5sjJPTfvKRpg4imp1EYUZHBFRHbvr3blRnnWqRQyg+ozU1T78t9
OiWC810efI+Mooxw0/Ygwy5Sb96lcYJbed6gwwXuUzRjNjW6OzlPNKqPemOzV9Jp
TNkKhp/W6CYB81yMez6FdofXWu7uuhOyfgAHuDG6d6Fg6I/251IypysO5dmX4+dq
MJaGM0NiGOInXXyJP7AjebsC4nqF+rw0Noh29PiBjQhX7V5F1ZJMmqYs427RE38m
Lxu1bG4sxI8WNT+blt6SL0krdRGo5pxODUlhNMPgxQk/SNYfHToVP9TCyRjJeUlZ
ZoD9akjJ1SxG1sDuNltAN3/QGGfMQFyhJRpd/FyAisvg0ws8GivDrsNaAIH8hpgn
l2c4+0eNGIK0vsW+iMkBMfiKQ07pzvLcpBTQ6OQ0nC/IKZPtpNq9fJQ0XE3UDj4q
QxvCYVBwZpM2sz3vf2SP1ii095WIm7w4Wqqqa2kT4555dSIMjiUXOZRuzuT8mDYm
5BBSDbszJTwJVI8UvMS1N9qIrmw/vC0BHbxLAqH4wLngMn9BrUk24t4t29jr8Nh6
hU3s1ZztQYkim3c/VyeaJep/84uWl5E288xsmxwdm7W3S9LW7ZkIz3s951SFxGw1
21XhR3sa8F/CevUHwLsz3HMrQDXx0BQnm5F3dTgGmaacoxuqLTRwU5BB3l8wD2hw
gcjn5dPCnOrfNdFWDdBP1SBBJoKS3t9IQQJDtsj848tmh6pJasAb46BTG+fwrE4X
YRTcEZG+zvghJse1NJOfec501XSdpAloK8UpR3ZU3wUI0XveWaZXLbr0WtoK1Bn/
M424r2dcFzpj2ZQL5bNliZ9Y7KkXOUQWIE1r70ZX4DZJoVUWxEn3GGdIhy004ia8
ZGDMWjHRIbUNTexS91ivW1M8FoYbXGh26azFUDP/WQCJNw7FN91mU9tyiEgFYy02
8mo/yOZvdvMUHyr7KCJZ7u/8GGPSBB/taiZ4J0f9YvICysSwfbhQKDnNGDg8j/fc
EHEAbbwLGJ2ebOGH4d8Qv/BK6y/5hG1mI7JhLrHG1terBgZ3ialphpLRwKt+NB7W
I1ykzJeAfGcyA1U8BJQMvZxBVPXWH18FwGJV9UTV1Zmohn57otBuaJZ/s2qCbVid
e9ekczkyrUXBmkYPkUBwKf7O2Lc7uGb/y8wDI4PgkAoFl66Q4vUzqcMxXGXrOYl2
fQfoWommjT23SP5CyPRo51gdUBtjuJQKAf6VkTKLrBHgpSbHz6oOszrl8MH9PGy6
gpaQiaoHSSW3d2fYjWUxTMMJF9PKdLYZPSd5RSGfoxxU1s1+fRkc2ao7JDXSrduY
FT3pnDcslsVSX0EuaCrUhp2BFcI4kD7514CISXbxXnxryu515hEolFcawHuvY8uh
G0xkPFrSMxU7qrpUgUJOonIr2QOd+/gjrngFF+SHJ3L47WDdqdwZNyeAzzp3z+c0
qWlP9M7+W3XUYSkk+F6zECydZ9vmgsSx2LIRhSi9B85VyRgYg++Fr70QYxXAkhC2
H6XtPunS5xHkXsgN2UDliPAO1Xw0CAB8xfOLovCEMWW57MqROmyPDtbcLCcsGKKW
OYd02oSpg324Bx1CXzK1h0q3u4+ALlykkm9D4SDUi2yFFuSk23WwlB/o8UbPzr3D
D+ELicVL+X9h9rqn0egE0zefd7Sy6oVejesZBGHUsssRTUEP11wZKHsjzUVdvLH5
ECeYlPrnFzS3lI8ORDs/yYiKWycqhP4avawna5DkhdL1lVgZD2JMiYwOmySrRm/T
mu74agPX0UHfh7182yx23QnAgVTnOriJbYjOzDaEQp6URPSayq5owRMIEj9eiWvg
dpX4HGes3ydBhzoy6/y2MtleUvzF8tTgpFQNCtRAUhA=
`protect END_PROTECTED
