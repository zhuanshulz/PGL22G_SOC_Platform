`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
um6G2ECKtK+3noYRJsMIHtjM5lDRD6+Dr4NaKwy6thl3W+w6ArGSMSWI+IZ0LHnr
AXAupzEWzupxLZouotxfpVgHYm805IvmED4nP2M2vz979IjB7DuRbm6eXxL4qev7
yKmUYElKbd109DB6I7I06fI/xgAl6LkvXNKnzkL+P3ktpz6D807vYiVlTJZ8UTdp
kMakzUwS9iUmokX2TwaHiYt2AsWfgpMLfK9t+BbzUh8vozuOKRnb6Jb2bz5xKi03
2/xVPalXcac/9xKtt/63C1dwzuVVS1IkUp1PIPZ9k3/o+hsp3QBDtFUeu2efrlNg
x0VcvygUJj1ZMje8D0BLp57co4gz83H1XfMx75wPhoQINBoL1dZPxi6b9lpiwxT/
1U/N+lRwjqY6b9X7TzmDApBwYSu//rvya8A7JpfpygrTkqB8Li9EYz8IFxGDgK15
dU4joaO0bXTFTr2cgMC/RLEnfdytOsdNbFvUGyOroj1WKgLL1H7iLf7jT5pHR8TS
fh8r8kVvfVtj1jwFFxHMeFf2RgkxrTZJTigh5a/rhEbpbokg8K7bXsF4u9xqfUMH
xHoY2fnB9lGHVoSGK3OxwB3MMFqj+XU/qygROmaPGtAy5WPlpTAPc/8wX4C6DyRv
jztiZ7GcpL0t4TiWlEevTfsW+iuBQ+Y5OEVd5OYDSKzgier0m8jv1bVIzkajtUGs
NsUgo+S0dcLJAE0EXNssu4Ij/T4Nc0No+X2hsjb9WvvtvmP2PdxbiPK3ezUaNGPG
E9dl5H7OPhMSYBepGiYgeBe6kHbSz3iFZG1HDNlHQE7q4DYwJY5OA/wVMoCDOlw2
8OsdTX4qmmPfEicHiYjeGB01lGuF3Ge05cHp6/FdMWSiCtrdBEIAy8W8yP2xJ4pN
R2W/8u+tcooV26UYzxwZSmM3seJq43Y9YiDw2Q/xQtpwDNbbFYC47mXeAj+W1Eap
dfWXfO9yZxUrAYOthMb3jYdKzivoOjtVBNQrWAqb6h1y3N+B8FFBex3JoXCqefHW
x+QtX9R4ScJZg1IpbAwMmtU9Q3hcBpk4oFhh3O77VIpb0FhxiWWfXaFNKYbG8bCo
8r5fVx6bCaVd0N5uQL19s5jzzU+5ECqJcSy10o4yBWSnDpBtKeqR9GsLJVQjwqKy
3XpS4aQ7UwJomk7ZH4WjTKLYCqnPK8dnOZ/MrfNvTgPVa34Y60dqmzLEVNC/nRLK
fb8Ji4bK2fW+Ow/EX4VNLb3HSREcEgyDgx31at46vYEZMESou3Au940NGUM9JH7X
gwKsszI1PhPyEjKQyHg+a5icNEfgktIz+7G+Dvt5gK6LYc7pUFw8DbcHyKlzGKtn
/LUshCjSCYwSKxBH10yi5C5g5VVtT524hwfpersmBQSkgFIOQOiaKr55Q7VRmtDX
u6YYKH5GNIVceh/rdGoTF09mQOlth08fmYoF7vlf1y9J8nq+3Ec8vc2jWIdM6nW/
q4OaDKZnVOzA5Z3alFN+eG3KrCHK3h82esR8RFSFrts2ogJgAOp3xfJC55CTcEAs
ZVDTY1rtyto4cNDcve61MMCLl91jspQ3pAyso6FCjyyr+rVl6cm3O3/ksHnOctzp
EpEDkuR5Id/G8FxJk/g6ft5OGU5uebvd0D1FFJlVZwMFbXN430X9G36Mo1HWfqIJ
v8jlfJUad5Cioavli7ZCHZXLzCE3jBttTvLW5rHUlsZVDCS4/a7zQgpiMYnLVXLF
ZyDXP2k9+pxYer3guW6kgl6vlY6U1nfTA3qG63AJCezyB1pkYl81jZRxMlI6Gr91
ZAongkSRWtpfOxCHkdbvb90sVAd8g3j1EsBxaWppLZlSZ4p7l2ywkkjYalz9AiMD
X1+leGMhCVnPBJa77K2m/5nvZG5b8SzvEPNcssRyuHFvFDiiINbcL7LorAvhkGaK
TKVK1nXVMKjvBR2wx8Hz2MDjd0yrsEBS57dzoVVBO9VZNjpDM1dMCUu6RPgSMgsh
9//KWx1wSwaM0QozJvlTbgk/REjwzmp7acsQS1OGNmW0IuUNAa3TMOvuvwc4gnIS
dQ9vY3B+30ZqAGiNnJHQtPdpP6tMBXq5KIAT6N+9DozZ3u/An6/idopY04VhjzmJ
YYrcVUgsmWANK+LaY4CzrKgrbjTeJoxwuMjm5G1Xj7dBFJkBQEDgj0OS0RYeKjCY
YghDa5Pt9+aFd9nsslL9tORoUU8Tqdpz7KuVWN2fMo4T9U+zQLOVZ4KeBqjPvxZW
SJsJM9FNsBk6n0FWYffdKkdhlKDiyOLfe6loQTGgdcwFwXDGkav6HK26G/CbyMJq
nQjq/u1F419ypiSX44PZpzbNj0aMQ8SrTxcznQlEsoJA1nr8ZJT6rfdobU7biFZg
Zr8x7OEgzr4EcXY2Wazr3lfEfQX00aPhslvfpDfGA/e6Usgf/RsRkKqW7Ld4Kt9d
WjT8eDGU2Ut5S21ZsKf0DUtU2kCUsoiTecMtJusD+l9XLMPYQ2DLdxFUnRqlQfAj
TquUWMSVk8agvP9aU7mP4zWQG79m96jV9yzHUb5N4XRdSVpKAK04Oyo33+3z6e4k
wxwPuki9Pc/tE2BryVpahIO/AY7a0DvyCRG2Ko+DAmEgW0rifRI6c/sbYXk1Pf2o
EbKbvdS630YqQ2432IbqmLNIfKvV6iWFQ8TDNfX/OmQ=
`protect END_PROTECTED
