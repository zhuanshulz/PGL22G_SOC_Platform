`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8dlk2uidqCFGbi9ipah7EoGo40he7aKNWh2Sf4RB1Cs/vgVpklsC73DDKyR+bMyL
16MPjMvENRK1ewM2a57SJN9fOfXF19hk3VeJ+yXkaAWWPy5DMOZ1dI3mCP26E1jS
qK+W5G6vmG59XJAwp0iVkF0lAYQawGLxj/mzkcOzNMJS9cdAK1kEO1dRFG5w/mW5
kWVMFFEb/Iu2BH58Ba0KzKIKMTOwhcFDYrCph7NLVLlKyBRioAikU2DaIzrd5Yw4
J73K5xKzUgAjUR5Q/7/FQNg44/B0kGUBwot6rPWBpD59k6wmJibMLaS8jkPPHOAT
XWxPQ0XENKpTZWsWXwT10mrk0pPgGRJll1vHoCySqGW65dhTmmAnvC27c5+wMoRU
WBo40Y47wFPnC1f+saRT2r/LBS49DspoR+NupVg/OrYLHhpS9EEo4Dz5sXgFAIKz
5+OoY9aIItKx6d1DqvQ6rmAEBqXJlPKlsqgXswXmFz5Jg/w2teAaRBsG0rThQxs2
pv5ZDuA5WA6tg1v7fMYxgXZlLCn94uvb3zjfgvyVBPETCaWaghxS4LnRjl4bbUiO
hpuMqodI6m5lmMu9f+0C3HRLnBlVEq1HjHeES0X7yOJd8yeHmqG9nFbxVtUtSWUu
odrNFfy5/SkIAztqsA2Yr6I9A0o8gKdf65rWYt5E+XQ0pQi+OIjUMxUot9EjV5Nt
gkSHQT5MxUyQxSaHF0vGRgqOLfdBD08ZA+XJ8fxOCMj/lyY4jBZwY7hSwjOSBBud
Bzlw+MukNFQ45nxrlzbbCith+YJS77/ryF6TPueXT0caadcIkxhsRtQALYgMzcJY
a1UA8lLQwkmaZg7qBnhQO+rmu4/a9DBOAb0UseENCrz4XuYJ6+nKIVkqBW+f25R1
1AFxHmAjBpADjNfuMtVH7bcDxSf4H4gjRywrY0CKaEPsdinGCQCrJV9vs2kZA0yn
kLZmlUNuv5Fyci3FnEPqJpISy3P0lue9121MymQ2RB1sM/9L5S6eanWRLbfvXLjg
umjF427UYDPwTbdWBD/ijA==
`protect END_PROTECTED
