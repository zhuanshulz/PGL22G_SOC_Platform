`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ie/D+I+tL9yPBfUDYXFU+stMdHbFw1kYIAdc7xZE8hRtaAqEIVPf9PqOdat1RKyo
zVqPRpv1C60SWJjzdvA5n2X/EwsXe80JhtiH4XaYGrSZIMOwtcGFkhPSJVgnzk0S
8R9Z5dICiglLIj50yAmesYnCCuAbToifElWTK7Psj9OnJlv1abvqMWYgd6jJHnRZ
YIUZLsuJMcZyVzAuPZ66EWIDWhSTQxxWEZBTg2MePKhFpNsnD+f62q0LJ4ezyWpw
Qnk2BnrnJLwdYrOp4yGf7BPqFtQn9q2ytaJvfcf3Ewj+bNGwS9mRWWydTHT3zVzC
tmCJk6hA/mYFkzC6IFlinkJRQNEJyyRv1cChGBq6l2XQbJsUIhuXaaQMsUNvJPZW
4/lt6cCvWgwDVUGvGiEsYoFK/u39xYwkwMQscOL0oD4OBzR388dHXH+oO9BsASSb
OT2/MH1h6CNIBYUPlZbS6vDlCj6bXsuTRzw6Nt66dkcTolezwszZVK6uGfATEHUG
/G9Wl3jZwIsuGQWMPJvUrpYcdwIAULFrLWo2GrAm8Wbsc01O4TycXRyOkGCviQES
jXziVh3PpWazpUFbgv1UUm2pmuNewuIpP/d4YMC/VS8cZSOo558qJmL9QsYT/rkk
bk0zYcgViQRUVf2pTsNKJndHt73siIKYZ1VaIcSJtiMmU4Fg8ozJ0jvsweYzSROO
FOJhneg93hCV/YSrt1sWu178wWZhbMXvlWWlKaWiWKE=
`protect END_PROTECTED
