`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MyjY7UZ8eRTbW7JBfnXODTT9FhMjgqxMn8QSuH8sD7C7/XF3DPurQEfcJXhvJ3H7
nmSzlQdcKu+gRHoUr1ke3MYKJyVk8QJVBvHVrCbPC1qYWGbOjk49TZ99q98Nj58L
PtOp/t0/mZEfa8kWX40rC3KOi9PNYuReiZSr//wKlz1i3cJsbxzBCP0PJhpfk6vc
jm7dsSUN6lQVYS4l/6/sMFnyJtcUiIbyN1zUvIe15Oaqjtp4yqWa2LG1w8ahHgg6
Jol17qlKQoiiMEQtLnHDNw5+rEwJHNmyr43bz0vdlkBy3b3s9Q/guu+YczcslWjC
zyeUQdLr9oI0Ahqyada/vmqnj0ei6ULktmDZGya4ZtE545kqPbxhK++rDXioJYuy
/bZI5BYSIwucHHh8GIo2Q40zIX9BTqzHHsa7UzwgMJaWLgMbPEnB0ghH4WDP2iyu
9/Qq7DKdmG73McYyN8nIZv/mRMECgWnG+rUNnaByN5lFBIrgpTTsu++N7zEvx6Gu
tk7bhOROfjlYbvsAnK7yOZ3YffXqjojD3KL5Tgk7JpequG1L4SLOmKDOaFxOFQFN
fKIIxlugyJfRl+sWGRm8KGRUzugI9iLRo+PvpkM6LZ1WBbEjsFTOsRWkYKpiN1gR
kThH+cj+CNIYSrIJKvyd5UHjzzahk0h54iQa35DxSr05Kvwiaml6SZjtHdcUxHUj
8Q3SETj/3MH8WyvXUWBnlXOWTEwwdJgrd0Duwei5V7yo0H4Jod0Iy6P3PVcCnx3C
Um3zPhCdq0duuLWHGLiBuFcDL7Bp3sA0fj/QK3s3njUGfgg+b3csiXOxaGJPFj70
p92WMoB0F9O6q5L8wckcpIuwxnGd5R/hWeSoyBRIKd3UkiXN/5uYzvTiJX7I6tSQ
Tq7nPo0YtC84o8ShlkiS197D1/zrCH6mvq1YR6Wg5oi/sO2ePGfJjCgMshpQlu2o
p4uY/ObKw63qCdN79eepaPRYIvnK4gzpNWc1hbcHdoBoxKA2FpSDtq1HqnLYGrUD
ED+k3EPrRgI+VfJTCVdVN//PejAH93UY7NybVfe7Nssx1UWUI/oh0wM92gWNbayL
na6k4mOHq7tJYPOU07Z+mEwqJ1WJEDxb6s4GDoA6n6SDuCOFdv4QzELGT+tzQb5I
Hq1us2AxxKes/ZjcrT1E96KAVaCaJI7+HAviu+vgBPgW9B0zNG0dmoMk8+XwefoI
97bv9USI7M74EB//y3DwAxSFyRAu9sAox+VtiWUPCx5VkWXX9eRNh2d8Xk9II59T
QnmgXOXxigNc1ZfHWWNVEJigQgkkefApH4htOmnEqu+qzwMpP2b2JMyz7bcE5A5P
aPjut+AIZt80T+J+JNh51JtpjIWf//a4ysBjckRLrEVFz+bcaohesGrMPFWKBmqk
zzeJ00kN8OVpGXLjj37a80z37k6EgxSKvqvEPziPsrEmcb5ZyYYXn9wti9m5TnMj
oQRnKZVURd9vHrniH6iU8aITxSlzAU+jSQSeYz2hiSEeFDnpYY5AQNU3fmZM/xiO
Rc/OonDoazPrzKN7kSgms9DhEIn2r4thA1PD21tgi4jRUbmOfFJ+ldcrjnVFpzBx
e3WX4BRUmC1TnSHlH3BBeNtiXpiwS7lDaf2MvuFmqMUtjW0LBu3g3+M1PZm3SyuU
DUyhQUCdha59KU2RJW/QORZHRP+EtrMf2vu76yZ11LwHsiLKs/n9fz4FBkG/QD1b
crV1LxOJPwf7vwWu9190sx/1TwTzHPUpOXs6YX/QPpH7xdGb6jggjNGHRhdXCjYF
dixo9DQfY1wmnVYWaYkWDCyaUHt94C6t3QZtv37HneMbXixPvmiROwyZCoUsmb5T
u/WC9MGPZJnqy+uk2GTnk0Oag56bm9cH7+jGVFimvcrebQtgoBoMMb5QDYh5E1GQ
GmivgYpCfpEXHVnPrsq6hm64LMsO9r3HLkhO378ZWUveQ4lCS/QyEClbG4ADfNEn
MlPF5FzIV8NT5Mwf/OkwcLPDDHkDsfhFpNqONJFS8JLBMqkX7+bcmAg7oDr5r3XP
H5oc+p991QTIu8t36jooL1nOYQLD0Efq3kgNoEtAHExW8stw1hgNUlVHq6mvO75x
VqmKrWWaaoRWEo1W35w3eXU1dxdqq0Vwgb5a2lIFsgP37FJ9u1OcIqPVpYh6J4um
ucKr5SwW/U7OIVr/ajaKHMAdAgqAxRyrSDfy7YfKZE6mPBwE59vgNhffsq+gdcN4
YPXIcazkinqo/cfwzVpYPt3dgVNJ1wdfrL9UrhlO4O1hS+OTa8D5GuHeZQ14utvl
nX0niNWajPdmnkTkUlJe4/eJHMbhdmiR11nwDWiPQ5zMdI26JHiuXRdP0Lx6uA18
4Tvfc8QCd7X6s4mTVN4QFf+5KLSgQJ2uftx8wtyrnbAJCPVLLt5H5xtLAijbziUd
nm7S23n82v+SdMryRiKf7uvj/3CEcuhd3LXlqS0n9vFAkByL+VKD8hKb657LhHra
Scy/N1sYS2rxH8GWWDyl5RK5IVfmgj7ioT5ZF9rYzRkqTNNJKZlc+xpuiuDiGNop
lC9ivKapg8oZqQhKxInNOG8Ir5O371EgGGBFfCDQn9x1gUtdO3Ou6En9rH2PcQiB
zucfsvdOMHnI7xINDkBG7Wgzh7PeWOZrNICFzmAkNg27z+dmCqz0upZ98BNJ5ktv
7drIvGfjlDWFkjTMYQl+FUan5WdDATt/3Jziczm8OnKnu8Y9SwetTmQLhrqdxqyj
z938PvRsctNSgpXaYxUNBg/C6biqnDTBsi332Jsjadgc+jUMNyFVsZbgSl7El9r1
jdnp4ALJB4QRPBT3oxdw0M1VEblBmhIK/yLOe+xYpFXF69DnukMmsdXowr9eokbA
WyPZA559vm3Y28P7mZdvPe2Ii1Zx4HPkAbwOVmAfZDnKeFLaABxKA5r7mNK37lF8
DagtYYcL73Sz+a2q8uE9BMeFoiLI0iBs0rEaVe4zkPF10nkgQ5UVzsH5iwQaje8u
UROagRTZWK3/QO4M9TsPgkIJvUKSb8OF6ydoF/sYtm1IfqelT79nRV9pY5sN4bMc
VmcAGlBlQX9sTStMzcV6XeqaQdh+gro7Libw9WH1Zd008gGrVFw3WFhbwObTDm+S
F+g0Z04FbCQ3kPBZGZ33UvUGvOmOVo5elXY1DXA7EjdeqXLfMWhHgfKSK+vFIN0h
Ey+NhRbyubv9HWPM0QFjOgw1huzNv0INhUdlXxX7Ct/T75z3W4KZPin9lSs22/0q
/kg6zgJTgFxUl7v2ffJC/bb3rFGQ3GTUtpzlLLcZYasg3IfbpM8KJhI6U1z024aQ
WoEdLiZ7U/6VFJEXww7gOf0CORFUWkX7hSoWQrx4QFryJDSJ/033p9py2sVwMGuM
rYMFyyczrIn/rk27HyVng1CTv7IW9yQ0OImZxZ191l+n2dQLkDxjmKG1WlFry8hU
zZmmOKfWkE2yXqP4juvWBqetlTyocxVBaGkMpvIRP53gL1ipXX4oxqxSrmkjmOg6
gJKjzz/y5+9981HYH5FotYjxgZpUl/QvAi0je8U6WhI9mfwaPb+F64y37Q3Gkc+C
v//T2KQWabXRk/FvRI5GjFtn4IOzBrs7mrgzGhBuAGBvuOYkivA+Ze+X5zsbXlJ3
wxNiqXErtaqV69lR5pV45OfiUCrJCnMFmX6De/iG3a0B39bzjBYVOtjOROwFAXv/
Tsve48BgR1frdOEw72bA/sykuKrdcLJiSL+HeC9GvSTExATgPB1UfMXkxwztJy3U
/ff9CFhR9uBY5dd5hqO04mGDL4iZjSGQMYLaL0biVnSOHmHjejX5fHDCGJR+T1j0
BvMfdUiDf8LCKMRYSDECRbbpIkKlllahmqBZpCcTDoQqh64EUbceyh4dIagZfrEO
f2uZfiqSUogPsriR4vtdRtZvnNrQZcNdsEjlzeIBEmD1JkKxQgX3fI6evMgxvlC9
ditC0oNclEdL47qjsvZHd2J2VN2z7HnRYTx8+7RMV7xlzsZAuQofShLXaytZqt49
4h1gguWV97KbPeI+oHxi24ksuWoL0Bd4+qWrmegLQgvbPgUfgINoQ5csRc1WVT7G
+a+cFmhUTWA9J/UdkSs5Bqjp3GULCbEoHbvIZvcyNLuo91wB0WFru+lKWgR4OTbR
a4komcQiLp+lUxDNAiNVsP6q+ImEQMzR6YYTT6hXqbLd/aGoqLlc9nw5tM/kw8xC
Iba/6fkubYJdnV7rVldIP/6V8OrqmZNWFJaKnsjAaDa6Sv438iVpCn07Y29t+2zH
zu/ju50Q9rADxV9HUpca4SEcIgtOqyNLDzzTOAY5CjSnRdyBtgnQvXSFdxOMseEA
fMQKdIF3xjwgArpwsNubhwRu0vkNdkIyZzpYRGNHmY68MSh4Z/nWJvWTXtw7ZwLf
ndarV7KeCvFuD3DaRv7PoyBUaPVsYiYYihl7uiurM1tiyuZV4yKYxeLDyqKtcNQP
BW4MD6uHIlGlAm/n5fw9BqCyxZbbAhGXMbcvAhKPAQzEoyio443vJnn/iiWSwnsH
K2F/WnFYh6OwDG5b1Ro18hhXwziCR2SxNSovZg/JT6Dm0OBw6PuWzRjX+W/1nMhb
abmpHkPTC2spECNc4NhhZdn3Qa9zifP3iTVSvY3AOSMgMccfxzhOd9LNbt2Fwj8y
leqqYwAQUdH1/NbmwEK28cWBbQkGNdaIlkXDb/RXXm/ZvR4lwXiFIws6Jx9GKhIe
GJ6Ermle880kciiB4jPSf576OERdPC7mjJU/ayRcFckczHmZPXchZI4jyBkZVGOk
WCU+0DikoiL3woQ8N3amLUlryoaBp6gC0OgVq0FsuN9rdUsO6ksHMM2BleXUsJn3
lQaT9g4Iqi3OMWG6anPaDCJRdcgjaw+VQkdHBl0wEflHBqqXAWK8pFTC9B1WgZTM
ao4wgJpoGJtWlF0Psbzt45EqY4FMrFMX3n6jx1B9w9So/ijAt/cc3lRGOChw3F0u
h/NhCpOF9r6fLCiUI3bDOsA2YNmYtNEMVppln8xKmLc3o4uFX9wdgMGx0hMBLpqM
v8aHztb+kUpxErWV78YV8ZvhBq/sBVZWAa1HscgtUkjpk9KZv97x6cZlpHMUNbH3
1wcwCdZ3832EFm0OBWQqteqopklgSlkxWF7i6xKREZrRDUDTRiUuxR34vTL2z4Qx
Yc0lCVZN76932VeCmUCo8FBPOxu4oJDbXkgr9pxRtF/FxoU/gctOLorlugPI2DbA
PK3Q60I+H1QuhlJzR7TyU2S2efe7SyBlfjvYM8tJ/ndSjCYQ1iQ9phe7svxFKu+K
ug4mYupsMNLXFGj/zCccvNle45NX8cxU/Ht82MJ2nJuf4FKT4XJj2jkbWQp54zA4
oGibMCrcAEb42MRm2WXUJvFSS9pI3qo05r/93Ln1ulrHv6comotZpHhqZyhA4HU9
/f2v4TBtuIrbK3UgOIE+fKAQ4D0pGAImjBCowmCz7mZgqwZgoH5yNceAnWuLTiyq
ktP0tsUzRPpkQnHk5I4PN+VoDHMzhI00Ia1LVJ/MUve0U3bZoOqCJ9Mk+VQlxrXg
GZuDWtrGg5bQXW8rKij7yy02hZuR/HR+Gg+LjY8TBqk3/g5X7UwWjW8jh9VBADSo
ENwqOHq6B5sIwDNCb2wN9Dx0FBWwMUQo+Sm+8x6XIJW/ZAJKd7o3cDXp8MjVx/GK
f32Dx+oXhwmdL3rtUfZDLSx4TSUef4XXX5BTE6Z0qrXHK+RfCJZ6Kf6t0ZZzIbob
FhG+LR7J7OrVBy/B8LsZycRCHhFKbEfxHT74R7a+3bokDCkA/N7an4qzW7TkWcd6
L8ti8LG5sm7N8hrsBMn2eZN+fR+TlcveJ+P1MI4MSUCIfsRvnZLWoJ3HmP/tepJC
aVnBQstQ9FbeAJEpbBmqrEh/p9G/gelPlhavgZCzw9C8r8q5Uit61BAfFX2Mk5Od
7uBRNPiLd03ZOhYlkabM4j10yhtnmWuB+F2C9RywrXHaXKSpolSmUFFsJWjCm2e1
0yzknKIXdVFhNvY4upMQb45PS7BIcggRUn+0XgVWLBgpJsp8fwuWEolGrScN5kNz
0EK8n3VgKQHhqdx47+hXl0Oh7PCN566BIB3oHi0bbzt3IwExlzWmho9sXhg8mTLx
w29R3i1yKHX5iJTlbLkGbZwVs0Jz90FeyvjE2Ye0ZwjTDoG7hWtbYroK4Ds7Kue/
EzGahDtY86rsA2AMgu2CL0eUVYW3gNe3Jrc9vb9OTCWHSnHLnFXREDpWNYKMYa7S
yRNi725xrkjKC81LlsDh9fV/7f3qNo0g4+SOqgxiNvsPTt3sDY0miuQRO+ybq+l5
ZV5pFFd4PyAttR/RiZHAo0lM9SE4K2mR0efD8/sjnmhLcoI6t4RRHVCHLWnEb4xt
YtHsdfgM749LGH++zoV/5MkthsjGbcrRF3xJV+oibYKPWyi1NjeMlprj/m4ey/X1
7cLC8Vz8dP8VlJV7TAamDwVP9WqjcAxcYtEmsFRPGynxgOykM2aSoQYjsqIiF+QT
zcBtjhuPZkEC8WUo3i0QY707DlZpyptoGYvYQRmoNvAp141LGoElthM/fmuLtSs0
icOPyEmtgauruZEzrm8ZGnq/jcQHN3gTeR8YNyoOCGjrBdkM+bAcEJys2oqKJBbb
DXg4Zlpp67bl80PRASmePlzu3CM4RPD9lqp8+nHcpQczlmLdxkSYTWU2dy5p8h7Q
dxtsdDFs6CKx3JT56L/ciF1ftyky1dg+4DPxzpmzmIKXs2crVxRTLvUw9pjnDIiv
jQZ3FEFGklelWSrC3p6LXTBnD5N8nAjq0kKSPOOTmovgtOYj/3EY2yYYiqSv2lgd
vlPJ4uKsYkohQ9MXR7QmYtCjTUo3La2jr0BPWBPANyeYTWUUX0IlRH2ljbkGup84
8suS4jesZ6PkqTTVD+/tL/iHOwmMqwu7LA/qGIdDCM1/TC0rlQZT9RrSuCJZCMrH
1EOkabIGn/UeZRXgzk+clwJNoN7aGccvh3T9B32ki006bLjytaU0fNbm1YmbRhTX
B/XSfFh/a1p/Lr4CJL2HhgYh6BetrxDqZE/CGNmbNDzlq/G8Cz3SvGayuJeqfcR5
x8oEPf7Y5aWdhaOWBfdVFVl6OkXW/83YgJzzCzp8BEDiqd3onPT2wjzOnUBJa3Xa
KYm+r6aWoKguGZn+wqJ8tpKlUiue5QhnkujCDw6iE21jRgnFHkmrOcNlX1T63F5O
QIbltoyXVJDnvXVhFMUd1IYlcpJCQkhqCIuoT0C3TyrTbeWb9HWZgRLCGViykq68
hipcYoibM2kXFpzSbhUEWz7e+27DR6Z5mORekMO7V8nhv/BZwHYowEQYP4iEXegm
w/zG6HkkKBg8rZcYtoNF9Na+G5BTPHG3fupCNnP6dB6uECfbfqkeR3GsID0zRPAR
X9jii3zAIrT9PDrrFomdGxIGs8Z3sRkAdB/ewZpb6y8yneEWvwGcH/DIhAUvdATZ
qss97viHIr4z7vL4AmWfo0p9+3me/APGYexcOOftP6tCla2HL8dq1aApkZQCdm2a
vZFqOv09TlF+KPJCjfIjEd5RhdTkXlIrQSrPKO6rBzXMc7pEOSkTH2HlFLXEk6W6
M4C+XN32zRe603NdDelSM4zO880bZTEz7/eZxk0NrVKDLphvW/K2ZF6FgjvsUh87
VeyH8viYhkxG4u09HnKHNKVG8cYY6XOwmK0DNKZpDBE6YdOQQeKjxDeeIt6o3UVl
2pV6SP0gzQwJH4mOz+JwPfY33kfIIw+lQW+aqHzVkLrPU8uSmZi/JoAOE2MCltE2
7EU2P5Lri+YeabX6wiBePyUV9vjGJIucKK6c41MIiHX9dCprQIj8XOZ4c7YJckRX
gVWbCMTfa+BXHR35iuxnASZHKG9uR+3ZOcYxr18gTbqKNlpSYDa7hG1omsBdMAPH
122miHthrgP/4sBoh2JgRUVDSQf+IjvcOz+Tu0K9LPyGaJCjDkrxAv76UsN3YSZj
efQypPKk+MFZzFVexUaosX0t7bnL0uRWECVNQBHYJZZXnSy0iD9BnSOsAOP7ZVql
qQrHGuUbvPEr4WfetgqWc+fTbYcw+7IMIUgaxeirjbJbJwW8tqQZni8ZtvPc4Ltc
jRgX/5mqDzeMqEd92DW1sShLrizI9qK+3+7fQnd4xv7Y7sZTU4A1xSwmy8sEZH8/
FcqaQgEkLqkcLB1JIPxllL90d5fhiF8T3qUAehq8iNn0FmAmdnSjcLJwwELYux3U
T4vgdLKj5fmAAhKxGkgUEJezxVyjZpejabEpwka/MwFRqOYd0BXLMLb8C1wbRn7X
GmFG6nC8261TizBF764zsT6x1uxWf5UriC3OFukYrjA9RvzpOypSKXaHJSGQ5nQg
FRT2z1tJPmeTQoRW1q6FsWBDcxddgAPI3Cmnup8G3MJzOhLHvMnUXc6oMpBe+ukw
BI9VZDmO41+DjxsJk4Uf/mBbDTTUnFGlrK593cqbVYppAMfuXTXy67JooEEVYxKr
`protect END_PROTECTED
