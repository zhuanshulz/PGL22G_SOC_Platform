`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1iqYSMIZqu2EgHJZqY1Qavc9MCklHZG9uyBE62rPmUmMUuKKf5wwY3iPReCt/sYZ
/iVGaXARfU/i0ZyABylz61gZwTXH9PbVJJr0JFR5Sa+CZ9kXNn6jJzqINz4LJfVE
S214ON5ZVFd4OQXpARWMVz3L1DlXWB8yRopC8qWjg3J9VXI/C53pbkyurfFkNDyh
lrRh6PJnZeA3kWRaUWmVZKtE3k5rtWKGYIGYyO0d/rMGQlZSUo1vMbptNXq+6EA/
/mZQjVDJgDAePr+e9r/EYNjLbXDsV06ih1kGW2ncFAhJXyvufZE9/c/Ygo35CHQ2
1GDPMpPr+6yjKSiDKMS6cM9fdX9awxs0nRXCRTsgrmAI7X7OTB7tRO2XTdM2M3W9
KVO4ejgOcIdMNDxdPF3AhEhjdVX2UTaX7xBOW+BWtstguruPTCn0rzEgslfCwhEe
tVvBr3ps/o4SXcKJVOQGH2Jf7AXIxEz5/QJ7MS3aG4oztZwyHe+XcgmKfvXnjDZF
6bnnIbLRh7djfNyUVUGlxn3a22cvxO7QPP0T4mhkz4WY5JsuYjeGvMwiTX3P+91v
0oQLzJO/fvX38nJomcAgjXEtp2qhnFh/HEF6QqXdNjElYGtxDcsqHObDUnLPkWKn
pl7vx97gUZozy/rEa7NlTgGpngv3gAIZwcSuEqR+OkWgPSu2DLd5YOSvXePibe0v
1pNUqhyktWl9TFpKwuyvKptaKbNRKrs7fzHKIvaWXuzSJvhLHVYoLnnnPPNjBO1t
8QusyFOAuogi17hLJVn9EWu3Ve/4Dyhsbr7/TuPQl5flgyKsr/UAzkd6pT/L56p5
eCvMAaTtfHyKIs9C9sjJftRDQCw6c+Yy5DNwrFZWPp1uGzzDitnB6DuXFtIsYQoC
14EkoMP4k2tcT60iXTat2imrJNoJd+eejScjAVqh/Kh2DK6iJOPOe5yGD9a+Ap7v
zkHJi/93sRARdPGiw4E1vNaWbGYs+eASP4CeW0K3WEb/2SPM4TBHqijoOKKBInAl
aOnWc1uWAetfM4f81rJxUp/kNuoXGUgcO9e/TBapLZbvda3InXv+zv5bzw5MiacP
HPYM0sPmKMCSlFhI6yiZvHbyZ0IisbCCUa74vzTuJD3jaE1CpWZSHYlttUfyzdQ8
Jr80zb+huq5ZdcGbcg2S5HSZIeSABTei8h9rO6PnNfPe3ZyxgiN/4lKoneun9+eo
UXivb/mHq+m1qlEY1LDArpqIk+DL7cay4TcJ7XK1eZ9VxdEpGODBK1hQZqWftfAL
kALFZN13TSWQkH3ikV5qPaqQGIZQvFi2A27ELpecJBkF+WQQjXRpTV4+4RenJIPP
PZ3yekQTGoGvTe2JkRvAskoe9l3mLp5ESs4JA0bByQPdyNx8cHtAKxPQ/vXgycY+
dxb5eRHIEw6bFEbReIXW0FA/FmumPWW9Vpj/xxVBMcnJkRMLHHsrFrJnv+GDC1ja
Ed/WBi+NsR9RBbGgTrwSE+wwfXa8411hhPNmflDbDlFta5jXdX85DBHyu5CIuOo/
UWtQ7dYg/A4KLOlUvJCQRNJ24h0G4yeGM0K8lmbHesiLPggFoIv0m4eK0X0eCcCJ
cbUGZvBkkDBno8k8E2Ab+3mSe9Slpl5vdjXsQQ3qDZ3OT2BxtY3C2SbL6GfLYA5Q
fGBPVGhCBuoc9Nx5W5Z4mne5W+MfS0JDME1SsPXdx9BfpVGJKGcV0D40WaG/JmBd
Sv+9ZgPE1eoVCwZoCTHwUAY28feh50lnSjdGbtahsnBTJw3+ZKdcwBbz4mXSqjYX
kfSFB8RE7l47S1TvqWWlfQMSwv/u8HZb6iOm2nMsOVqBqTB456OFwr4LiWRmXBJN
ai24vaPAYml8hgCF6mmsUCW1pVEVf5k0Gbn0A25Yadtc6PW6c1e/Cdtao4YxVJrO
CLElbSQ7PpT4V5lQAeICssCy3nUMNp4nzt7oHMEMiZwRdGW7+C60wBNo+KZNgqes
bh94HpgfpPTcrGvD32+YREmsCkAnBOPDY849jniEmZqgEyIOJiraru7GGLNjei+k
T3lhDdW24b+7yU7UawpYIZP5p3Xmce1g0fQ1/0h34VC2IYver3D+nnBZX0fxLRZP
ZFXetzt8xAeTkKZAfNOFFoaGx/eeN5VRIcNIG6zUOxt7kcyX4UOX0+lxJMbo+yZH
MIXE4JnkY/AaR4bt3+lLaqtP5Jc7I6RHiU9xuw6LhXKHCM5Mvs+t0yIfeTX3Os4Y
m6qPNA3wpIqXT01FnSMhjLAlQV+jR6wpj2VgskebRz6wo5WXc+f3of9asn57jiO4
TE4PNxLeYJ9zvtdNJZz1Wu7ZW1dZgzxwGlmOKs5KiTtRggH4KbLLgnGkJnJKBads
Et7mRqEoPmpQkX4xPl9ipQoJ6qE31RG8Y+cVm8aY8tTKG6ozCpYBPwhNXaDueX3a
9Uo5jVfhS28VzalfHhNTwhUMORL8lirx706V8vvGlEjuau0g4kawdir+CfsgkGlW
iPoo+nzR/8NRG3bgqQNOXQrR/794+iPtMkhk5ZIoMinQR6dl1W8A0OUyhTVCeRD2
b8R4lIjqrGqU8iRqVhVFBJxXTs3lZNZ40MjHeDX37i9wjGSFAUxER2y1iFOwoVuH
0zf9lrI37SuMhHI4+kr+pDcvlMV/g8i+Qm1tc2SLEr69w7vNw1DY5NPtDbTyGkfN
wqzi0Z6gx+ZDb8uvzinwz35CATjf0/IFkyEFxnI/OJm/4a0FugTkjb9XclWzE+Ai
SBrX8N+cuKwN1XpQ/T3N1LXwEMUoDF/j11H1bZPumcBQMvLwVhXZiA04fddgCoFg
MMjsiBDkhscJSmTv5vyODd71nHwqXzuFR/PSA+n+K9SGedWiR/KQDg2r9ipSyR79
xribUBwTieauTeXWj2f7X+SNE4D0QkO8lhUCbwPKeBZyJccXKVJDoe2IXWdDNxyw
DiscoXKmwobKx7jq+Wb8Yfxo/AuZSUaVBTbbkdNE06dSuGpWv6SFp7yPRPLxy8aK
zHzhG79pXC0H4A3ZrSMIMMXYFBq2AuU0q40MJ19cbqG+WXtC++k6DFfuZjfqzzuZ
4D+8REnRxhJimObOqTrIEUcwJdI8uRxbq61F/rA/fXwc6GgRM+wyI76MSV0vMxAu
qy3JS+AQz2OQlbFqIBTWKsFD0wFs0jlU5hGZIRWC4vcWAEH2HI+Ppkw984GrHTj/
Uw054HQ8hiQKcdOtt0Nr9m8Z21etf/F0Ue+ykLw1DRsXIvfIuFUGGCjNc6uEJ357
DKEOJe6HFAs9Q9CIEf+QO4xUwPOr/FPWBeB3jdE/9bTRq0tdG9yAix3IvF/ZK6rc
UOHpX4vV1yh7u5LHynfTqokHtBImSD0Tr5/5Gyng8yrfS2i0U6QMP21MSY2KrgJJ
ZQmB7Cl3zNCAPaJEIr9cqKGW62UQAJl88TdiXq5wzBHra9e6US+ioOVyKqz6+gzb
Tj54xy/nSuWiWAkje1Ps5adTC1MCileAQCMaGvTT3IC3owmrLfA2kktbpxLVfJMf
xVG0QoRzovsFL6dG4kkc2w==
`protect END_PROTECTED
