`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zJAWbpkilsSmb9uLM9fzpDLqAwGh8EMh1nBkUxJflVXOVrJ1q8V7QujiM95dpBdX
uILSQ3ZGUECzlb5/QVG5grk2qEP8+emx6hCHBprCAEzfTa4CVUW3OSZh3AfpnjEy
BtNZ2Ws04pf4Me/xxY1+zKcWo2GMi9QWodo+eE5sr56/FJPOpjmWBF+Ze7Ms4HiB
giSacvADA1fYuUSVQft089rRLnbs6mge93EzXoEQmNMlPDpEkX1A4/jFN75glmEn
EEPa9uzVYWQ2Llx0fazcmwDkUASPwa9x9gOkmHJMrnl9RIC7d1hG3F2XIPF175BK
1bSNG0sbDMatR+IbaImq1AovqqxCgKOZUDm9Z5gV1v2c17EOUcFqsSPlfDln0BSr
zfjaFWvg+Fk/5pBzrkaCzmcKwX+xdon2sAG9LgAAVij0X4swSB5Mww+0PkIHDtM4
YoP+TbvtXZ1FfHM/PjjGlFQgpXt/ipMJ32bCq4Nv/DsZmqFnC7GNCUdCrN6Qus6t
tSydLyAJlv6mS1T6NPeDFR66bA+dlRDHRIWTEysuK0vU9ZDrXx39z3YKyU7h2kfQ
AAha3/BwDFAeVS91amvVlBGlcM+LPiy1LpGKgm0yqEXkcrN5t60GEehhHcnJ017v
Esz/MO5R/seF7K7XePaf4IZLzCajnbJdjQkEPef7g9kwCbie+5vAmETh6ZaPBqid
LRXEx4ecakf9IMUAI4MzEpSgBCD+soLL0Ycme0CR9LCo6LoV6Ht3HsCUqT22YNNc
cVUjYBXRIhxUAguw/xP5In4KIb/4lBjKdOW14WPp5BvH7qHxpCUOvPtfibO1Dhlq
BKD8r61Fds2aPuAC5UaiHcUmH0nz+N8w9okqYcCmtMBaTizkQ0l2X/6vCeZyl9ny
LTpVm+46r4g6sWrE/UjKggQvSH4nvkaHzxwM+aHU5aTlUYuh0b70JXmM1YseA0VM
dABCpT19KOmC6WdvwixjaaLB+KBouGyhuo9CYYg82hmUo7c6NMftk3x64BMrf0th
cXFxprB9pnzIwjR23qMBCA==
`protect END_PROTECTED
