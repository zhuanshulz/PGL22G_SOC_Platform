`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pm1nWOmZ+q8XDaFxAPrsQR5bEY21ubtsosvMPVKiizNlXFjCwXnxpVye9jyD8Ax
sIOn6v1D3lxnBPpHq0zjYO/zhQjek1wGbm62bTsZI/9/nr9fXcC4OPBNHatZ2v+Q
I59inWJPejeS91HQ3k4M9URaRcKdvDPKq7tdDD4A94L2A/4nB/sYrF8PaYcYjtd9
rBvc9+IyXh9oubNTqoNhZCJ5kW9qpQHpRtzkynWPPWiovLTOY9eFxXHOd/1TJbna
is+ev6nkgfdyV5YyU+PabqbDk6hBIVwiCJylhkxkW0mY4BjI97Vv6f8MEe2MEgCK
lDdZCuqrJE/BjR6iz7Kiux7G8WF3yoyvOSxn8IxlO9Gv8ON6Tjmss7tASp8norXF
pTQ5XYo3i3vobuK5liy65zYpR586r7hSRX359JsI7p0ySJPogTJZUAHz97070m95
AZJHNngsW6bxzkGaJEaJNzfk8codHtWNT0rBXkFm6PPwM8qSrs2Oo1pnJU9MX1TU
dFgWifoKrgZmUMnLDTl+J/z9adIA2uzR/Mxs1H3Do9CirwnNol7OW5hqTgwNstLY
KuQojvrQyZhRcpRMU2g9VOv4thcJJf8CRpFppO/4F2BFSMkIY9ruyit1z+HOtKwq
t0nw+i1XxEJ46wbpVYYCNcEBney+pSo+E1al1P2O7mB4zDic6Uvj6cRMwoGgPox6
qnJ/RYVFhQumtbZ3Rs6nxJjzJfpkFU5NZayS/cXFI67ajI6nsyIx5qVUYjekvqJV
TDxt29lEdcQWM4THmlR198Kmz9+uk7Nnfj23v7nmxXThAesUmMINgaqm2gyMZN9Z
g63FPxYhLyN8ZcQEL77hqUAuoxoPEOAZeOeQQdJ2f3Nut5RMaMKIYeWA/HmOQMco
CBpU8RIyATb+1wdUI13WBYLwaBbOrB7CcjlR07wM+tJ5lfli+81SwDtW6v/Ncr9+
iRspdoasX4N8scjGEjTaThYWxSVQ84gLvexe3pZ4UczLXauOR6ctpkvLJM1ea9Le
Y9G0GZhiJ3oqwz0z1jq6EBfJ7riK4wB4FGL/J0vRZUZQS2OTqwkMWVwQF0WEShaz
GKA3ZRBWo70lVE/q++ND0Dz7tCzktHShIZ8stG4cUlJ8Pa9AYQqiGKQWcmVvNx3D
a4vJPhsMbsNbrXtKQ9IJR6Y9h12dlAwr9amSOiQZU2AqPM/p8QHjvs+zx2NJy5cr
`protect END_PROTECTED
