`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Et9f3cG3+yHyJa52nJWBSl4hXpaXer8/PUUJhacRBp0ZJiQKJcSEQlmovo3T8w9v
LndaVB9B4KPmPv0QDPJmHSq25sCPCcXtxONHSGGLI1s6t20enaieeMjxVIwleGUu
Ocjom+sZhQ3+Vk8bpzIGNmmrbIfDrHH6TTF8ImG399pKy7EJyjvQKb7kTPcSViDM
ir3y8hMe6JErttCz1LMDK9XLC6sbUevlfpNtKzLhRGgK+JgEfYCxnIZyRS95XZGx
fsxBEt/HkGFGY+lmCBEl3J3WXw9zddThDPwj0xxHcXgb8ekSbedfZP4XOWZprqUn
ALVBz6OZN7MF3CW1EzTqkbtyMmjFrSRlhXceycYt7pHZgn7ajVcmQ8UHuqBJv6zg
AbJl+oFIjLztSaSoATQhB5a6I/Ai2XHFlDqJmAbigTwjrT8f7T3pm1/N+kgBUUIG
2b5+R/necPJr9CKh4WDusUahvFoTKE4RxjW+1X71LrLAGchlvrcbytfI2axAueXX
y19LmcBbIS5mLvaxnWuazBmcRKRE/9trVk8M09QIunuQfisySH/pCbcQQk8c+ZjG
RpksgEGYPE9yPEUQWGtUy2d5FZB20wSF5i4qplAKKLNNCrQSnXdF1k5kTXRwoonM
`protect END_PROTECTED
