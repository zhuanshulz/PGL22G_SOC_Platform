`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bc0AnQhOvlGtW0XSn7qMTi6etngvBOlf8ggoWQduysW9Aq+6fz8WkKolbhzX4bDM
S+SOFijE+sLp3Yl9hrq9bvH4bwmUFWjlZ2IE9CN2VC3N66wuNoZo3qiKKN1Mvk7z
8tJaDYZEFN8E26j+51Zz1f0HO0J06tMVqaqAJN4+8dNqVIUSXepYD/gnfkF1A7V1
uzZpR/mL/0fUamFB374U6pSYO60rnx2G49I2536AWSntZiyV6XJKEkVhOJfcFTm7
`protect END_PROTECTED
