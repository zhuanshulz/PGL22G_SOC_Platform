`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X5a7ew/MAsr1M1hoM5YcwoUQshM83iBD2lHNL+G074sX3ztzykV9qtDLjiEfnX2F
ar+XUWEM6vBDzhL1oib17x0L7I7ZIP7jznq8cvaDtasaY/oPfeeS9fv1MfovXqi2
+lR+N3UWTB5vNZIxWYHj87rN7pWL03MCendvPj9/LwSTgor00syObuRzeiD50BWu
WvBch0WF1cV1oZjEeZMU1eaLFxrClyvI5pnb00dVNDpoMAPJeV9Oomgn6kjeWdO9
rP7c7VKH+6IzoMeSWIdaEQ==
`protect END_PROTECTED
