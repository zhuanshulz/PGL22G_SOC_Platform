`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Bj2nCQRDV53l9XKk8Hoyz43vHSHSxKkmcUu1gBVnEJDl/5FdYXCkqo+9x4yjILq
f++NrgfjjP1sJxH1DMLf+4HFXDc75rFQ97FA/ygjnc5eLmcLchPjCvFThJJ60wSL
kKLpNpGihpkyRw09wQKRjkRpAmAasU0FCmAk1i7c/SB/ifjEc0Do0VI6SFXDW+tA
1CNdpkv1Cit89SGncS9dGlAcgOQEMJfuv0w9OzNvoFz5QlXyeNsEvQWptkObELZT
t3UXIAXdZAjJUr8O+zS0LSAA+uDPfR08+/zm/2gcoMrnDVVqibyHiSM1JYGLAqJW
Jh7hEtBTJhS2rWsDZpk10yzI1tWzYNk7a4Ns/YBMFh/zWXLo0PFXMDkGbBST/bUp
5y+uiTIEHs5sN40kzqurM3CLA9wxBLPhS/wbqY7ma117mQc6vkuqSd1vrnrksB1l
BfuJ63u2NCnjVQyoPKBo0TFpPVINH8OOPgblx/fbAP/OkPnzXMjW1p+wO+RkAr0a
08guSQ0RM4Qdorfzzj/K2Dl4Un25zV2NtZNv2gvjbpYM9mJuZpYgiySEIiv7Kl/+
WQMwluWR00vfil0S62SU+3l7Op472Xe2cehs16M/Q5yuuxUmTngUSjpURw7iiV95
5s323b+YBtyvNXZyPHkQJJ+6DVeCYbRxO4vTvijSPFfS7Pqd6RLO8aSDImE4YtyR
70zRQ1F3TJ+g5KzPwVFY8fBfkFKJuJ2VQuCkKLWK6Wcmx0VKHPquG8ytAo6YkzF5
dike3IK1OUCjlyDawDkE1CG3Ad2TkAwz1B9GyClPPuGEugrV6EaiD4BLhPVI+v5x
IEDNe0SKNSPblfeLeiBONDmhDiEhDWx2K0NknwnxVdYhIxbczMKWcfaoqOAr0rDB
oakm5WMyuGaGzwNU5lRI67sXOZ/GHQip2ugODbO7NLRZ7ZTT/bxbNQooSbO0aOE9
ultUAie0haIGSp48z/bwee01BFvORwLOVNxcAkptWucMZd4WupsTVBBxSbHZB4GD
hSHAgiq/T0RzrklvApv4OpDmL1bJ02O8h7PGmUJxwdm0Kl7yJ64CKYUssIg8QJfN
W6m9P+hk010hxc/oyMUdcIb+fOLZ2Q/mUNbfGERiHqW+8NHxFkNmA9pQHohRwx+2
JR63qjPvfuVr1FXyu67Xa7L332eLTsXmzdY3GQnVEpXEN3rEx0UhAJ3dWjEBLhQ5
1ZkVsML9cWD7vQinxBMgkQ2TbbRVaO8RXUmQVzmCtXgVruLny5BW/C5F+IgqI0S3
DPeiV7WoiqKDaXNGsjUO+UuD0UzP3HxOjD25De5I2644l1gX6frEOhr0IwVCQqLb
lQk/FUYpFVye9/nEr9EODJ/i89RgmdnQHQ5OrEV4kAC8P7TTv6RjjDULHq6aqon+
CMz2KyaYPl93A7iIpxcDJSXUN3rrwM8jskD5xril/9H9NY93qsLlgzbgG9yByTSn
JQzVqoqHXQqm5uSMxb1wsuZWgXSZMauV2RVELe/Tsx2cKphOEnY4Psqq3m0dOrwU
t6aUY+gKLpsoGGnHUZz1I1yLs7oZZQwNY7dVFt1M4UE+K2JyKuDVOrMIxv90PZdo
VYeMBtiAav5IoiuNvgSBeD+c2+4f7irRcIRO5Xl6ksmIuMvddap5WpLAt7NKGYj7
CucW9XlvRYISXi2OKQSa+uzHj+itiU/UuK8UdIfnAYu0P0xc5b67/+fGWiq8lIAg
1X3UUuVGyWodT0cud2tcd9HlV5HS+34VoZyqV4GlQqv2xbSghc5d34rBfdOAS58h
wYNzk2c052MjBEMID2jo4dgUToqY1+zRilmA9/UxNqlD1o0ncNJuZsypYyjcxKEd
iPj+as/qTedcMOMl8oCtElYMSe1hFcf/GxrPkAZtPAj5XD1vJv6iLEynzC4P2PRu
4fXS7rAPfGHc9+QNX6KvN3j5JlekXT44fQlvocMNtBQE19/PcxVfrq9XBtcEwbtL
effov7Y7FbHzJNa+DbOqm3h6EhDQaCHpj2a0QHZR90dJMJLQn/hNGwk+vygnQiAn
ghtDRpPycTIGOnfZzgw22/BvA9fW9+0hdu6dWtM9KnGIgzxpqIgJ2TE88o0tZs80
M47k3sj2GdxKGVhZoYE1sbQN7phYA+/zhN9A7TTl1e3ZBSip6UTJuV6SRwBJ+Yig
6AFp11Qtc5fxpJkPt43G1Urf5cLJpQOHu6qZZ4BCzBCahKqxK64PBTbGCjIP5Znt
WKX3OLYLsz7hUEBI1WvtDp7RMTpBFy/RWnyewyEvtI6czwuxKaM6Xju0LutkYzf/
O5cQbcrLXuFbBTi/n4JzWGy8xXXZD/QXtoQuwWdB4z4O+w8pp5DemJDPAYcGenAD
`protect END_PROTECTED
