`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i3+wjKLvw+C824IPCqf8mmqcVCU8mBaXABC/sBGU4WU0Ba/5kGLWCXblqpI+NL2a
ar3dbmLHUalHBblNdiNi2XtH4r0Owc1Na8gfZ3SFSZ3S8EvRc/hAzh13CH/JsDVm
0ESg6UcN3pQ8zlRBklfh/Ibw/igK9VELLIMdt2ND/ALJXTqo5vUO6MHZGpE9n+jh
5ltDaZ9CrZPXltva/tsbn94Oq9ndT1hmxJjcKG3wsfH3X4BcXH8uEwxMtPEWDgfR
ESmuboktvcpqdnCOX9VCVZooeADfm9/9MuSi8L+BLDJ7L7yU3hsyCO/u+TBEi+6b
MGXXb+wyFE1sgixLOstTIbDhLleYyC2lp0fUVKq+CFhBNIXGT9Rl5l9N/FCQj8Km
6dDc4vsatrR+MlGeHj2p7eyHDs0oaYUVy95ypmWfyPVCcduypBBc+GXdgU1wtAUa
k/jRkChBS4tkWdo5y1BxFpCzthgew2nPqd+vYnQ4l6Z5Eb1nIeU9lAVYn6bJlkum
JWSs/y2SGFgliFY9cfxjVmAQ93hxPy/kfMT0JdmkcVrl1zcuRKtOoTL2OBPmehGh
LaREF3MkY92Sg9Jv2kgDtv6xNV3cqhnmULGL6nxeRZwe0n+QRI53/rAnarlP2Ioq
qbbMRgeken663PwIJdA2NuJ/I/fQzIFzMPNgbpPnUB3xfx0YNGjUZxGZnsRc4jAw
N7QbhphMx7hzPYut/5zptjmF/F8t6jcBbq3Z/1osFPFt/MUwwcinl+N7pF9/Wewx
2yVeZtEMusb9apuxnGlBlP5CSnnyRwbJGDapXLjwAIo3Xzx8KegSvMTSZHtQNMEV
ifuC+5OM4TlyKFVz6vpwmYL87RO0lcnIuc1At6hI8p4YI6Kxh32fuSoJi+7gpPzS
JLPP7luvVUmqPnlpHnbAhSIzhkcNK5QLucEl/PgWsI28XJ6kU/svuzwbTyJb1M0U
29j99TnFVBBrbiZY05dlwjf01W1Ay3Z+OF9sEY26jMwM9PsH8K9pdQxdga/qP0Xa
L060ND09ifhjVzVcIF02Zz0j0bHbWzuMTcvyvrMX1zEDQPysvF6ITm2n8Z5LygAW
50RuktuCCyWrNd+b97Ok13xkg0ZYkpQukFXrp9uBqu/g/8IRqez3PTt0JehxkMt5
MwZAq2mbskXqiEaB/lE5Yu8pKh5/J8+OjldISeWyE8QPY/FQTIjduluJBu1z0gwv
mp5Trkwg5m0DVPnKI4mQtjQ4NiVItJZWHPp7RouNzi3x4aZKM1i4gwSIz2pWDoBR
Zc/OnCwQpWbrHRbfxtsOkWB2HqeWhyrgigaLHSm0VRaFAMQm6A/oc8hNX+cNmpIP
6Py1RH5t8M3XKwfeiVrCAAy63hBVXY+22E2tv0fPPOcJja3pCW5ORsXPkSXdtY2F
A4z3vGVoPk3WlAl4NZLUk2AJM/6Y3vOdRlJqjfcdJxtGf1IQWU4uUpjDHtJSf6Pi
/tZIy8bdBNnDrXuHWrcrtNHQ5qDZcgEfCX8xbU3hMMesxjE3ANNHJjRH5YQhNry5
I0eHiWL/tvMtBLdhTiUS9idy/Mf3tQVeK+9VmiQcu0slDbucj24SElrgwxR5P83l
Wsrv53JPe5qN1sLS8xpS9rM4e4ERPxjD/uzOY73kPh0hRDJ0wa8nFWbDZxqbOXCz
jty84/hhdQ8lj4YgZmRtdsG3JKvGIqN4+ZKRfU9RD8DbaUOBmiEy1OlvWzbDV3+G
cmHOZHv/5NzbGs5qiwNiMttAkHVA/mxCjx5cPUCkhDSzXKmykuGKG35jHBEx09Q1
kiN3nqSpcO4y2ZqFkMXw15DozR+oZGbpE0aJJWUSjxpyngm0cPL8AnxATkMC+b+l
TlItkN1viZTONxjA6n2uL3HpAXvEWJ2CDZpnwyGnUwSYQJK9k79h1alqMZ66etkA
N47ns1i3KjKouVfRo7012w==
`protect END_PROTECTED
