`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEMU9PYSG6luYXUw29drqxGM2ipv+Fho1ve2eRFqBdYaY+DBeFURWmmKxkCEwBil
mFS3jyIvHvW3LTacKicpYQCkf2EwsbQr8JvsjNav2rZ4VaymN/RRsOF01FYFuywD
0XVUz4DI+8VnNpC/RrE/eTSf2z0HtedsYsP7H3CH7272y+P+Zd0hnGVpEQwzghga
eX6arUmB1Qagc8h7iqFfKErmxKpV47SGJcRwqYi6N2mLyPor8dx2JCPqJ8Fc1BIe
WF8zStJu2aotNpIMl3nRFc+zRT7tCTL4LUNvhydyInCaW/9wFNPpTwcB3D1OCM6Z
juR5/Hzvd+ioWVVIdFfowzbvKICG+K1beCVvRPg1ytnEhxShdwqxqZ4779eczTmw
bO6wx7HKu9D4HiES4TejYkwASU8z94PmYDfgtfOPd5k8Fj32fBT3v4a2YqvmfVQj
JPNBz3I5z8BDOpjfn0yksvFNGDU2ePllQQ+41l+y+hADmmFRMBr2ebRpmu+mXwmX
Uez/nqTklFlM81nVNmGA3sSJPwrkMa/Rghyz6snPV1qbuyqam2Ggulr774gutWfN
vSwZgvops3M8UyCsWQquWPXonSlKphdCj97/pqUBLdN7IzpxWMSizkeBcJLhKYwi
tnq+8D1xsFAlxZzXmtmh7Q==
`protect END_PROTECTED
