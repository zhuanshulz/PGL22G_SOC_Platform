`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
efqTzhJhCRYp1Tuz9fm+tlnqap0EpJ4X9ld2ooV6upVZKNZqmwr9Ouj7XrB68Ps0
hmD1w2ZGUCQO50eZZZEJXtNnujoL5bx/zHStzN1mVDtAbvWWM64t9Ukl/NKFNpGx
LgdwgPEOVzy/JiBnuGPTXMSnTpXCl0f2Fui7pL56GBrdv0miVRp3sctY2YE1phoX
BsW+1iklKR/9aJDjw+1PzV9MXBydhIujFBRsDYy5x9i5GK1lv6HiZTXMhfYao1MY
UdTf2MYvhJ4qrdqKpcJtc2c0fs8hVZjx8xiZqaCAh17NyPHpji+wtc3G8Cy4y6Nm
19NQnDtyWeeutuSr+iwtxdI1jlCuVpyO2WRVEvubvV9qjF1NIjZ+iQNo1PaCa0PN
hbSspo20D8eNhtzZaSWKHooWa2btYSdzT9Rf4gKz+cy41lgvcGI3YadKaAE+M2LM
jnVw4el8okVoIo3+7M1ne7otbrmPPHTrvBXvu4tsarN73QcKkF/GMWCK/o3Gr/DN
CEg4YOUAdteRuVT7MrOAd9wGK0nKhGi8qi+0Z+sFRfs9/UTMIgcdeVX04Wf7Uted
XIQ5I66Lqoa+CAcaS3Jzac/atlw6iY7zp8EqWGltAxa85vCLssmLTmXD/vBB8jbj
yUsAXuLhL+dfMSog/3Q4Hg==
`protect END_PROTECTED
