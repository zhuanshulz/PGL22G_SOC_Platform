`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BF9n0N+1DvWCQQUAXQAPB69AB0jcxD1cDSvH7DrOhc94WcSz8aMuEvY4ft1Q60F
giMvRffA+YslmmucjpZSp88JiqwF9+Ldo18ZZRq7sq1GjRsO6JsqJQg2uqp8OpTs
Bl6RJnWnSvlcj3oJE+8dkJGvCM/5LmQyYLR7Tcslk/Aet/3oWojJ8JQnXKhJm9b0
+8fMEoe15N/qJy2H+U7Gf2EpPEDflhD95C8vaQZXVOkP87vz7yB61NGHUO02sNo+
OTOGp6udpfzz0kUdcXGWN/vXc568U6AS1ZjyULA9J0Rh7GqIo4H5XKm+mspYjdb4
rWaqXEVPBcc9Ydi07kO3kDre84Kvd3XXzLSQRCho6K34JZVJvy40kkcOmh3yBtVY
p15QKjUVW3jNRnvX87SNdw+6UjFQm3bNx4f+x83Ou/K/sDu6kEL1hdtutjo2PO5C
3CL78CijjubY5Z22GXasZJPA8lSvUVw8Sl2QKFO/0i77MprxoduEubEoscaNyaxP
atdxmNCmLOejSLtdCBVg5w==
`protect END_PROTECTED
