`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtmkW8kKiLMqRT4ECNbh0MdlhvVon9LJUO2LU1eiJSN2A5WSjrj3W9beQ4ZCGhHE
VmPHwLQAwV2XTILioOE3R6gHhrtHHkEak6Jomjd+l2rY0fRfPJzpb/9umMSETArH
kA5nCVPzNitkcPBMKzttO+j6pn9Geo/xtCp0ZCYJCIhCXtywzikZcohXxf8zpgva
m+yMBkFBiH30CkWXeG2J2CAW7KbM/t6BpJipBmPB57kIogj1tvkfc8CB507XTI9k
BFa3iR99+NTLGytBN6Lhdbaxz7TB5VYrGw38xhYOSxfPHfUrc8Y6k8ny10euc3k8
JDpmeG719FvHINjOpOQlV+lwChgwidBpXXaa3NMDNlQlyznUTBcwz1odIvsMp3oc
fAoZIkl8a5k2exSbQh/9cFqR68HqMCvB4dqoh8ZsbIc=
`protect END_PROTECTED
