`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OcNEj16K8uf0YlJjScHO5DajGaAwsi8fdpuYh6rrHjpLzGmrSOPMM0gUcKlKiGD
l+ttVmgOyIE6PPUDbJsHz01fUEFQn7KXGqrU/C8sZJhzXw6n/sLOCD5dtGHxR58l
JPgE8AK+AbnHzUQVcVr+Rj3kyoYGeWo4pDskYs12sXxKuSTN61moIpjW9I4Eh3XM
u0WvGfC7HnNgjg4qwlkBLS51dCnW5h6AKNI6TtFuufaagtk0t4PyIJaQXtE/swsj
zGMpmHe1JE61HIN2XfSminerp+OG6AtS4A3bwwmU8fnKcGpxetfK+kICGwN/QBxh
v/R4EGcehV4jtX7l906CkMNma1Zb2UR+oOsLPn3jXcqAywA2+hZKkFzAQat7uL0C
NpYh/XrpG4NtNrvf0TbMrbf9Pe7nexlxZAxwxhiy9Ab2vsiU2/UU47HBwn0oTCUp
CeVQsjJIDA0QKTu3PWOeWRuiFDjghoQLJA7oFZXaSdQBEFNWu0wGHMUjU4ejsr+q
YUP092Wjk757LCfim6FiYNJuFFqN0DT3dz1MhC3VJ3tYKL7Q7p1Rxs+IglqIk07i
nRqwjMwCPdKYP0b/kSonazfXUZ57fIvzp3gDqVBkhJp5tIXrstLAJaQIrCQlCw8A
ObkXFrOPEcR3i9l86/sH9FbUUvEe2CzFGqUXByHZBGWrCy3Bqv2j4cwJDq+oo4TZ
SdRngU8eIgOd0yDPwTuh08CDMFAs52rqpGR9hcye8wQNLRArJ3Q5i+adpUfsxxm2
pM65IJOgOqsJVfulyUiecqKlJqppSWp1BeU3ULerfoYoz3U1CeZVEMlyM7knJtBr
Ju3hbHwtZFSU+hkFAcCJYwYHxJobuC85dnVfwLPTjX+b8oKlM6+UcxmOtj8f9oPb
nirlrA0vfjy9igRfcQdO7gtwf922rYOMeqeOFIr7TooCgYUtQk6NFLKU2hMyegt+
BJHN2DP1oNUjT82t8l9iSQg2u6ZeU6VLN+7Iohhm7ujxe85KMxxjwufggXOGORh8
A6oyJ1XrfJmnRXMf9ZI8x3MYW3H4FqFBdb03+QGFmY+G2BQ5EOJGLSacrpjKdube
nn2bD9+2JlmBlCE3GKIhwgia46uEf0fUOu7etKOyRf0sx+HkqldauWtiv0nPn1pN
Kccrud1OLNYw91+lYHWEDjw/fsmFE/uO/bszjafZPPFrpb42BmSK2E0Cm1ilPudB
0M63nudqsD9dVevkkLRYMnlZO7PbrGCSUctqucF5lcjod4LDun7Z/1raVO54Cqcr
sI8tVeZlvueiCUgz6UvZSYsSrT0vczRqSfmYiFUJkQ6BR2LxxJ3+po+iSewpTsor
ZcddIHOgFlER9LW7dasCcYiO77GNFe99fSLVNDkdulkiYXeiBWOii27/5tNvOu8Y
PhhhXPgYRLV+IAAFt05TJxBA6Zu0/IVNDsrMJczhmyA75Vu0/vi+CPq6UqfVvfhR
HREXHojT0pI/qr1AVSRv7vF45JC3pNO1rNvd/BBTxCVpoTk8ub1ka/vgQyzbl9Qv
BJXWY5QxaPtjGjIzDL0Wfdp1pwidEwvr65sqGZ8/28m8oPmtNbTOHGIiyhg6ydwd
rcGPvDYXSEhvzHUHzOXoAfFV+t6iN98GJqj66a8uVXx2DNWCkEFGtTDdljj7oGdX
`protect END_PROTECTED
