`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EsqTM8v7JQi3ykbKLQ4Nw8J8YH9ctdm3N0+k2UpNEqCjkF78b3eTFBM9JhR95gEB
DJ9A4hzKOC69dPLAJu7pOntC2c+42uwUo4RuyjsTn3ubDw04QSnfSOqLKNB+PJeT
THalGAZNR6jrIrpxmWWVtP6WOpDuZZfgPQdjgoHazO63SwXt5deMb4qPB3qfgmRK
AEBLRa9zKAH1OD/ARkcWWF2rK4VgdM4zB8O9WGsa19SGwLZ6sg6sPGuw9o8Y8uiq
+zB0XiheTIHffbqfYISe/uvZNp4bHe9eGS2x43/1UsOXsAbMlEcri8IRX4QkZ0Py
WsRRqxr3zvNYIIIpMX+nIMKaOAD5zii5HYAOzBI4DdWjuI+htWP13bJ3L2UcB8B+
Xv9/Esk+irEiXRRJeLthdm/RZpNuTdEmro/ipuzjZdujPmh39XBcOPiNd6UGWYym
eMbsFpzttcCQcvHcXgXVbKC5mIPtnrsyQ2CTpkCowoqdKpxlKi4kvywoOwGSljEv
caiyy1206IuECUWt1XTBvwn3PoxawDSFvO79L1u/bVD7uW7sS1457Lx6tGfV0fHe
/77B4D7M2CL+4Sg8oLkH3tgXTqqQVpa2BFIhRk76A4MBie/vRfk930aVdwnhFToB
U1b6GXQE5bezTXpebPbf1PEjc/5jJnKemKHGDuESjf0vo1bsKnfI9ueAQxt54b+h
FMWJTERNItZrZXYMLq0FoyM5YB13dtIOMnEdMm2Y1MgTJwyaMHHhtKNztj7oee8g
vSOZDKjPPAt7sxLTg0KKf4BBzXgZeGjubS4IHVBEfHCyVzM+QqZIVqLrj09K0E9s
AOOaaxfONUojO+tT4CeSnRBZ8KraQDGWcSj/QhFoRlNJlVCIlSiS3pJr0IMRQMy/
cRM32GaP1OkzNJt+7cSVNIfDw7wY2oh+t2IvopLZB7+NdZs/dgoyQj8i1wQvKmB5
051obB5Fs5wyS1RmgueBxUhV/xvShpAZwn+tpiHyRHylqDtgWVpqfDQ9W/o4egHi
CIPDd36P5mcUCUXV6S/L42D6ZXvSlc3Q8DJVBcIkmq8ddPbbrtBvA+DSMMjmC3/6
t7OvYANaF9r0ckXegolJiTsO0HnaeH2jqhbFuhH2JldXDTJFNC6Ccmfbva0FEfoc
+K41llmBV3DpyvyKOtF3fvVqD3Wk7bQYPqsOSR+wiTpy3r2O7xMjYyHhRW4v/2Ay
2onYvRAoRw0t66NOY96EHjcx43BEluS38IERKt/IWrdIJh5E7QTgtfAtmpUZQjVA
P2eZ8QX2iJzLCOpD6QKuNGKdzOJaS7oSU6K/DvImCps7yOn1FwA3d6UkQnIIeeer
YYClW/Sm96OBzPXiWBBe7ze1/VjMVt/TM4BvI5b5j7tT2I47EGGgwx3E6ub8XW4n
z/9gR/GCJI6qoFfa9r/+oJh3gqFu0sOSWy0V1zj0bteBIdXWZ+E+isegny3SFaC1
33z+fcIGAJizzxfgG3HdHdcp2HLrZdzBY+btU4dsSpYJ+gTx+xytO8odS0rr89YO
PgxpC7VHpwK/vCXryIMv0uTLt8Rty7efS932K+PDemDc6DnOiO8R2oZwKqxHfvWX
SLHTLXHFJ+j5aD1J3lV7hdequteJxi+5nFmpbFKyDfx9LQjxhCbiGpI7HdrQweBm
MBFGBnLpno/6o1EcvxB8FpPI49MPkbL3oM/OYjTYchM37sITtxux7YLYgWgSdoLM
C+y/bTnkWRhVR0vleKub/PBE/NMxf6tcF6HDGXPUgiSui+wul1EVzkWhwX74yhGp
dg3UsgrA3lxUejyS6slLMboF17pImS3uo3tXcdx4WrB1ki5A4K2n+si3aR5HWTFr
N1p2K1YMsili4J4gVy406898ZKy/qZ0XJiw13sSBjS20st8PZsuIQT1SgRf8eysK
8LRA4DlDr4PR1CFMTVA+DHj4oC6cra9XMyjtdy+hw20ZG6UHaiKCIGS0j3nf3kKb
G7JCZXE84nM3LOJxWW4+qTNqjpdQ5a+3VzaISza1fVcIuezgllox/nDR79V1dmZ0
7JX+akHBvHLkKDrCAz/bXbW+A98D/rI87pqGQYVDs+w1favCuUZmGp6QilOyPBqP
zww9UMNntE7mEFDvPGkrArySjJDKVFReXPypvrxidVP8wbdXf/qjARuSzCmYbGdq
L2rXlHpsyIISl1S5BTzIBvlHHxBf3CulxFzOa4z84kcvXthPYgAr54+NVaINjtWH
yCSQDqanKypX2gx2I0RJB0fdjvHw5zyL/8YQvGrkxtqoiQewkT2dq4UWHs7ksbkN
vNdKRlK73khlSuH9miIdp2RJsgWtB5GPxiCiVaew8gwaJkBSdKGBXLuZS58AxIKt
AagwSzsFiT19Z/xbNp7QSxasHVjgqGlHvkGm6QlezYG9HeE+TBZ+RoHZ6dqquUC2
hu4P26gDLh4QdOTxivWPLiSDYe/xcJiBQGKpXHLrERMt+JEQ5CJTiO3AEMin0lJb
cwkpTKHKDQ6Ihfqeesh7n79LktS+eLRQX1NF9YtmLuyi0hAb0jb6KTm2eBxqpP7A
T4eDT2Ol7nWqcRmdsqxggHsf578vWd2XM2kyQjJMCA1jKQcAbWiAEXB7tc4/9UdD
FHiDRs7AQXINMjhjtteABiHVsSrgp+E5lgW4N+uT0NLlY+XUcVxe/coK5Y+mj7Jp
EY7FDVvNzh/FaKpQIpgQydYuH5vQTmP49uV2jKyrGlFU4exHWxscyaxbkYKQ1Y2U
ibtwt84wjILfkIQZyaT0R+d7ZlrpKT4PSsN0xgm4/E1lzf2x2EbPZ+EpWK3QF6fU
JrAjh/LBZnyK9B5iPN3YFE95Hni4AybdcpUgM6JG2UVm7vPo82A9t69WgJug90HC
sw8kqeJjQsSV2HBjN5B0xF7UsOoZcKTTcbBRnJTrekLWvUqHa6f82nqCRQtWVZak
Nirlxxhs1SrdpSXNPQDbDiep9zSqWIdj+Pe+mN436PzzdFDBYvt8LHSlf0st42Kx
1i96qriIBdDBWt8xc0cZz0jK+E14+jbVLbtYnJ0T4HMxTRcY64dstu/jcemcVBO+
rs7L1cIUqAkPvcG7uyyB+fQ/EG7TTbV9TeNHPD4HVhEzjr6Q8RTFPALagZob3LHq
8onxkoHIwb1DI2DEX/wjsHSRzYsCPKXKpMW9yQA6KVn3PyEWZi1cRqehqaUwAevo
ONeXYo/DCEKnv+NbzwY2/OEMojgab9NHG44VFnhdHQvlgn1Thwh1NrKOhJYWw6ci
JTboBW/1cWOu58iLsQPLkXLuXaHCsr2sW6RzEOqsaxL5TTcej+ZCTDVjHzE9Fcaa
KKcgDAsQKbXRJxZin16nR84bYo+19kU/hgLC1xkj6n9tsuHpybMiKMIZcxQX9shc
VjUj0eFWFdjT5NcCJr+TMpVBZ0IZvj3sTP85b/6o9yxYgZ82QVBtLl50n51l4Esq
hZ9KuBiaeo/4IdlGy7xHXgi50VPeYAkGtWBkySc2CaxHCc+lGyAjpGA8/HgBTTOG
hFuH9Brkt5KnduJZCRr9wJPCIufC7xx7PIczkCdRLtB9gkX/4o8tlQ7b5wUvo1PG
tZVqwYmGrAC4wtz0zN5+lzZoJNv2bH4IRYnUGA8Hl7XpoGgZnQj7UtCZUie0wcwG
rMaaSNhPMegrB9crBp4tke+k/mk7Y86XIeEDLi9vaa5cProtXpojvc5D5LiiFW7m
4IEqHGtXN2aLiofKM7DPb/F98vOgBfiK1WXcTJp0a+j9VueNrYkOS1GIgYbCurSe
SRvcwcIzBM7nZneflGj1m8OTza4bvUp54bfkWPLto1PQaXByLqbb3dmpRQ2FBfHA
ZWEoBOyqkoPOyAIexmUoGdAVJ68+yPO2zmJkU5pNu3ZBcjPfHSg87Y+UbpEbCGIg
kh/0uSyG7kbR0nrekscUK1zagL8wqeOOZSmQn4KxQHKWjYqtR667kgIDkiClxCGZ
r+/yRycs/zGgsBs5ulf9G6qq/d9qVNhMkO3RjWLm4l9b3j23owvg+cv7QkUEomd7
1xaiodtiG4O66R0EOL/CWYwefzWm+FeAA7MSH6xJjtQFxymHfpElTd5QVm61x8zU
rtGobSgR+M1pFem9aP8pp6MwE7/P8nWvZpUGZroRo3dpM7T+pjMbM32v/ljnZNr+
UkM1Nk3rs6SxMBmekaNY7HggPWQ/AoRcemToTzRYk/vcFwXuPVzJYFseY9DFdv34
hTazLnEOG863Sup/BT71fIdBrovsDG23MrXKVC9s4CdCqZqsEPq4wXR9Fa5eC+za
36Y5hQKgTocUJWzCtUvrSuOYMpwW8hEq1+1FWHeZW0XDkxGqTdCTsteGLUAd1ipW
KfOOOZs88Sd2fv8Kh20SuaMZ55GH1of9n+Ovxo5JEnqf++ySD9F5MDzLjtanJ2Np
DEkXnnNugcvvgzKhAiyl9+NJKW/GqWl/oU4yd+AOqzV8lkXDX7ltUWBUViMxB/Ch
wDbcI4/loeRoHdiCZtIPuxZx6n8IzPQTBjH8KR6Ndxbuy0XMNavMHlo9w23nMGpN
WQ7+6RyClyt1YKUPOZnoo77lm46roi1m2RDaoH3kQFxWpRPa0u1BglnwZ64DolTC
AoP++fUEB6NTa6jl/ddJNByvsOIvVm2JVAJk4l421syvWZUJjjL7Tc0FI96PrwaF
gCFoCkI65rVfDaQj2MQs70xqmi04Qy+HFKje61q/vtrwSd2UK26EwkTOoUxrHY/G
3ldjmH+joxV7WSfd8oZgPHYfxJg9wPQBZT1Ob9kgsDi3pyv2IkgGRwxyw0xP4XVf
G2HMwtZGoA8CS8lxA4dAC1+cizIOxibuMT0nDL5Rlqe0sP73qa9G7Tnf8pLkJLGq
diwqdkcOd0IypYMAUg52YLdyVfC3eB7d1FbFMT/vJuAH1lJ4ZXjglBlbM43ao0SV
5AiwjbRwxeip/WmIn812DV4U4br0nIMZ6c/NUruQRQ25TgPeBDFpiUF+8ai0Jvh7
6LBrtQtovLAUjd069biPK7A7MCp5fxT7Am5zRZpXVTgPqDPY4qZBvczw2pnDy70M
+puKDl05TnSfgFE7EgbEJdIAFfl+PSElS+lPE7/GA3qIHXTEuVLmAQWPh1E5lb9I
4oKwQyrzhjByOMykwJXyxm0urHHiZ26C693vfE0Q7QXyGzQFXZtLPXvAA41lBLx/
yfSddkpjgQzPDUZf5dtaKMZtNckupDZbOgBzVb6L3lM5N+GONLfajBrj/pn0vEBc
LWS/Tex5QZChWKGvt9ja4KOEb3wvIucHmqrSc6aL5elYP4IlDqkU1I/85xZq5mNb
GiOvwptl4Jf2LCNc5ZormwjsWy6AW2DOXz12XBYPzfEvyswaKGzM5AXQ+d2G71Lf
3nTwVr1nh/XoGxKbbj3keeHxJeb62pRt+IPEv5m5tOJ39KTLgMj0l3W1QwSHtdq0
l1Eu5Z5DEkEuEb2zCOx0aGNI6aSGLECQIs/9S3Qeyexfuba6a3LJ9llzUJEm+8ba
SMtavBngRVNy6mNbOmH7ziZpoaX7YUVyDNwvebSA/CA1UiDKkW1jwIvcbX9dkfTg
MdGumBOpGZtRApdOAhBBeq0UVxujSR2/2GB+vhPw7ly0gtG8CHj3/kmz3CU3q9qs
wpnSk19phP/3j+DEhX6+g6oN+b43gsyR+6RTccU7mEG3YMrmM51oGMnkIxPiYy9/
oZ+wSxvVXBOfOxk9ZfP+ndZLOope5RUcgzbx8/Q0vMeVg3Z8aZpxM0e+jgmp3APD
qWfrSlUq4UtElqzSb1TgiB5YA9qabxAff+MFatu62Gle7kflZdFS4NpIZG0/Znci
+KQHBxV/8pJisDHSjk+8TsK2SlR4AuZ1pw6N+SfGdttlJF6ebOB+MCGfuXiqJgMN
8GML4FmYxXxmQ9cy6gJgHSIgMJTlMXqebgfLnnbJofKhFDM6L6odSWN4FCKBKd6/
AlCPvpOP1Oso7GYU5MyI4Gyx67k1e6HyYIeGCztL7cqTdsFpWYVYUVyB8jdN6Bgw
zdXcI2YhaEibDG4QLkYl/rGDRqsup1mIdGaLWzwgTpMuimn0l66bBMikCL2v9aFZ
Te1ks8086chJfANpz8XuuGy0aAGmP3ZINsILFG2KsytTmOPPRfgJOF5TiigJmhmx
FrQ2djydlTnkVQxzlD/Jm2YmKwC3127FA3d0XhwEabR5Z3B8KtBCg7QHxzEhR4Xu
hCl/zd/LEJnbNNudehHoeZ3PsFte/9wWeiEsUjEVmO4pDjnPuK5J/bFmMwkkQsqg
xZHG8XYfgXMWPCbHg8GnqkHzYSpVmdc8wE68qsYCgHuvGfbUaQZ5T3GX6XWYby5u
A/ILx8QkJBpz0/dC2yNah2nXO3VlV0tuIY9xe2+if+lfw2yOhlbFn8VPXdXjACdd
4ENW8cCVeXonDqghH/fPwBILxSAN4xSWQ4Ge/lawsKPEXzUfJeERRj7f1Djq7iep
v5K8AZxuOKc7BMDUBr6ZTVL8H6xKHoYWqllb/0qjR63xbRApfNfleGl2FwsLd8HO
50CnopvG75WF1OenBdhDSHD7u4Ypi+UYiQGJ0o/P8noo3YEExXUKKEhUbvqLj6AJ
I1qeOuixCgT1G9wiOaZT+VX3JyM76Ir2QYGR8rc4vH2lYanjp8DMBCLjl7NTR3oC
mc1ODxKbQ+xy46Ze9hojicJzahTL70WdKNED8JIQZCskdHG92pd0NlaLKVwIK8gI
/qGoKXg6j8lGm5ETrPCwQsBHVNLnzjd4LaaBWngbISivCTcJ0pqAVh4P6zSUSbjY
2KiUCyUJwfjrEX9CufWUMGbPwVCB9LqZQEUMdMJhPfB0dghxiFtCH2N5Sa12eTZo
dIIu5DGoeaW85k5f19HpTV9ReTr6K9M7Wcjr1zSHgJGJFW5vP4suMbepFYU2wYjN
gwRDt3iHkq0f/aMkGb1c1Suisp88y7xvcbP8TWoYHxy9HafL61TeFnCQsA7/k0Xe
e7JapeUbXXMn3jNYZSvNpnDQHxYhq7M3nRsmy9SryGG5DwGBNgf9GzxzlwjAQZrd
HpWDBQRcdfT1F1zCvlU0QF3JFBoib6zF8K7bq8q8idGVhr96Y5zeZucVBgTWPF+A
zcfVa+M8xdDU2PBqrlEXHu5acdUtrVP98rs4a9L6CCAuqECF/NG+Mezc8+cRG4Gq
+ngOFPHPnqMPkFnUPKmioiQfkq64fqz61SBdSKjzEgFHl7mHU1O+Zu10koaq3osO
9xJlGheKCaj8ObnnqknEAvKZ17CjgPM0V+G4U88qWwMgjsHEhgx/F6gd2uYc0RaV
aMxTQcjfaVreVd8VTsaSJY/djxjERpOFOBPKV/GMOXIIQ2hfpANGdoIzbjSV1iEk
k/j7jKSpRduisIgCHOJWTMNZuUOtgiB9jXtUas/1dmQ2gCyZPS3j8Mwd+ITF9G5y
7mL5HrM2PMJBYCj2uxZIBvhpQwDoOoiNg3stxSwHkvUbkgejIGYR3hBcmuGAVBPN
Lbefo1bOVEvCQtNZ1f6fiOdfXwxYGTPsK7B948RzZM1PDRi0pe8BGcsx3boJ1KR0
fGfHc04Gs759Aio9UOFNcvEAQyFCwLl/76dx6AdE1orBo2r+ObQPx/fPyUK6w3OM
gicP9/8BOhtwGAw+ATmJWt5jvWl/uoO0FxEIYEidrATMj/mfz7qa5B5p6wHm1tz9
MJCRRysjGARQV7LJoZ+DF72dweq6XF3yWwpB530GkZA1crtcPL1Ecf8lrdQ9g/DA
SlbuUTcnX50pbUqUXn/bFg9vMv+Q4pE1UR2Km6KksxDnn+Qa0hMAEBZcW4kqTVxF
lRRmKf/CX1eda3xd2sxIsyZ1w4boarFLN1f8yfQ3EnbEQR9MA9HAYCMBDyWBr3zF
Hq9DETQpoUeeDNw/M1FaNpEGgjBg3gZZ6YGezJ2Z2cNvVNMp5ywHeB2y0CFNX4ff
GcyxtDI/A3k8Ec/hRh9sL62sFm5Cno5gQb1WOeQs24d7ihqZ9wZSDegiTMikRnqN
OIjeAmKZzEWlxCH2e2o90EhxIoVf703DKoEY6l/UTVKDzxxRZtqfM405TDaE6fRK
qkSp9csrE8D786PtV97HUd17cV9eHBcmXP/DHczo51+0sW1RnRG9Y0XyAhsmqM2d
xh8SLd50G7ye6JB4r0cR8KEkB3d99WgSM+fY/hCBK83ak20Hdlvn4BNFyKqdgaES
9+uZ6hk9R/28aV0l4Xumf15vQproGq3is9svXF6NzCQBD6GjjgEWuAOKg6CvDNy8
hq5BrRjVTizP5qV8E8FZHcuopXlso9OHplk+0XY4yyCEHx737dlB4fXqSfgJeGJS
/IWOZhOL1nn72s/PzISKGZgUrIg/OOONSyc0g6UhLnaIsfKHRV5GgFZJPaa6TreQ
QtY5b9V0TntsBtqjds8Kt/HAegeGVd1wcmlgUWfbegjZKEfmcTufhifeFWdox2ue
FelHREYQwR4R0I4bvyrH8o4IaatsfK+xgNhZekMS/7/6jfsRssecdqui3EEg5X3I
eAN/VOj49T4+9ZNrAwG+YNuYlC8A7XOkUIHtyA3zBx6y/Y9TJHDxJEwxKGHvzKlB
Q1CO/g5Mq46aOuikSKk4+q9MF5s8nyL/ZEVPjfas8ibNJz/bRbd50MNmPkG3dRl8
OWNbSzcSCKFWeGT1nWRF1PSbiK4ljzn4hEvN5HdTs7u3lguB5x9zZUr/LN2+BO1o
o/0YskaQv13D4HUyIit8lPtEcWA0yBQ8HKE2IglNJQZx/PP2uTt8GeuVdsXk4onq
hmmSfynjLNG+ww/hBWg2PbMsEnvWf6/XhET7bp76pB5dmfExK+Xom98VPJStcYiT
kG3ZgeafdiCjn+UVFjyXDOq7BVMTPOWU9IulwOqIvyUpWyHwHVYn2ZPLpKrQct2k
urFRSL0Bih0MWe7Fnnd3+gqJwlbW1yzHs6UYyxOLRoE2xXZrTbrO9u4W8XcPdaTv
r3LJSGGPigdcJ1sm3UgR1qCzGneFLEY9Ng7x1hCFUoc6H/kSrt3D0Jw9ca0VbSpm
+HrmJP0oD3dXhcCwQj+r5wq/tWVyFcXKiYnen9vorWhHo00Gnm3YxNsB21+gJbaH
1t3UVfMlq1QI/nwlkOCGldHe8ZEbP3eTALhoSBgyn9WnWjxKq9lmGwWDo5f3S4ku
Jbhs+gYXlOHZiRIiGAM0akk6D/GEwCIRT2rV8X7d6UgX7P3WE16gtr5kIH86EyQ1
vs9vs+wqyoj5fKBl5y8WY25UhcPMH+Vsskn8FL8SLcbMEyg1vvSDon7F4+mPu2nz
z+lbpx9Wy96nh6mTMWXKtIHB83C0zInpXy78g6yzGx4XhP+E3slUC84YW+eIx6tu
6hiPRV45q2jIuEGEUDuvxxmGrRepK2rVXAavnQB06shoFRrSqHpRT/r42UmziqMl
rm8Wrn7BU45TaEeTJ1LDLz90H7Vw/2utP1Pb4L1G9vGvIzgKmEv8VFqvH9/fRJ13
4SfCmVq71pEi/84W2Lx3CkCoHTRUgh8vtZ+nCztNR+mVltPRcSjZkVSgk2Ye+Eke
fSZFU7uBWYpW0CmAXexcRx0p/jAJOGAkNH9CrZDS8L38sIvxansvpvf/bA2xHdht
MyDw2sk7WEz26YqqYPZ1azW6pnsJFwtDna932ubEQncJqEv3sbeNagxu4SCyAEVK
KyfPZ6BjM/Sz5BnF3rrF8tHhlF4oVNJk5PHxNgkSsbgAlUYfjFe2ssNVlVbGx2nC
yulKmcxNTln67bL5fjHd30l5fAuJNIfUPwl4QZXEDbXzu0EZrbOaRBSaK6S9uxZN
xcvQxhWohgYX4NASxVhh5/ep+c5GCMEze2XYBi5TS2rPQZ+fUCxLend5AuZgivdE
fm4zJSpksCV9UIO0qHw5vssHyCWOpUo1358Cl0bvfcAavm9YG2ZVEC4E0AVXmV5l
3zwg7l6Rbjn576oZC70ww3codrHhhxhWeB0OlESBk98Cax2Zp+4Ja0Kv9E1EHtwy
d43tGlJ/BTchXfeqMGf1nGSw0rGZDbWdo9kl8enLblo=
`protect END_PROTECTED
