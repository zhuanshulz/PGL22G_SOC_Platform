`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bJsQhGDhu2nCn1GA4w47s4SCKahLagFUUpClPsTogPJZ5HAYfwnCaK59qCY+1ZM
vWOOlrKO9WSfOuXu27qTd6/RZPf7KXWvnCw8psAMf7f2GYugdNUyGl91RcAckm0q
pgtTEZE7WB13psR5TrCuaQx8MpUibRlRQGTfH60guNs+xfnycDo+31J0xVZ0oVzq
7E9WRs7NrLO/GJ01p7RCawSJla6hzsHlxdj5fgFJlXOLP0OToyFuYiKscx6YdriK
l9+CItg0yEQk6F1N28Rv86/7Ud5OvywcLBZ7hVrNagf/aBHuvJ7c+jj9k8e94nLX
flFVXwDl+SiGtpveJic3CLW27Bx3PykCyBPOSH6WWFhBEBo8gijOaOHPAbuPdgaH
pujbHBmd405UMi35nV6sgymeb2n/eXcbNn9GWUbzofw83Xjy3HM6XV2th8jO5RDs
+b/IyUTX9RKDaA52LpVvKJin/yTC7GAbZLdTU9JuTeXcjIZ9o2C4o/dxTE3I+iRv
OWM6fomy7vb0+B779ARY00AJoSkrMZ5mMpjYmsoIiFjD3zL1DRJ2aZkKhFR+gvgm
k6rErgalr9YP3X868P1iNpx/F1P0HULktnL+qfgKqyvAn/89AJRzvGq8rvqm9DZm
HfAne+RhUrog9+/kL5hMZrqGXanYlyfrKAEYnED9G3+r+oIWclcSmHS1Dc4j4757
V3Y5bp2mqqSipnxtYHPyYw==
`protect END_PROTECTED
