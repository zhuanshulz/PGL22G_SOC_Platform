`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AysQsL3wFv0xfV5CJwpSYmrrydJlmFZgGTYCHucmtkUB/KqA9W/xwrhQfxx664jt
Tdnyy9P7dG7SVEtwSQi2hokNJVmOsaQ0JPhd8Gd0OwdgT20638RH6mHplfTemem2
6+Xxy5Z2kNJipfnXTYchWCrjhjlABn7U3/bH+tlayq44qGqJLYmDmA6YIa9pNhzQ
fmSYaoQuHEwD6pmneQ3UZm3BfoW29hRQuBVWc1By4yYZCWxa+Xlh10rqy9g5WbYy
TUgvTQzTjGJ96HnQgJ7L8ADgYoAJ/G/4+3dotP+ytl9nrLElWo2RG5ybgCleEAsY
nInFEInqsLqrRabQ1mirjiOoVVyB3G1l4ljN6867mumRN/MaElTBPPzbqdjGntTb
wQWkUmOHSPD4c89H6gcsZbH7uqvBpK0BfnjUTV+zaCRWbx/qW1NhGO4iDd4TJEt7
WyXlTsYmy2Vt2zOZxf+rGd30Zj2Gwm6wqNSox3hCp2uYUDszJ9DRebFnm3i/GkdX
bGNwYxWQp9eghVgax622ALLZb7mnJKQwdSGyVRKTMuFEa+GP80zFCHZA58edjb4/
VgFaUNb15hoZ0B3diPxal7EERbHm++0C+lr0fNrX9AUaSdbfjr+a7aSeOAKvbmzS
F7wQspOEslAAhR9Kts4ZSgK6VHuwzNl6FA1iweNw9ysjg1kYeeSVmGsNZz8PAoe8
cGgxCXrIvsDdiNDmXrShqT2+IeHnIkBZlayiKe+BzjvgDTWVtRc6DcM82cd0hp6j
Gx+s165z4VpeBDjQVTQIrrGVGYx3MxCHg/hf4zIO2TfD/UOn1G6OlIZlvcogwsY8
Kjgp3V7yhUIiOh0eaU7ooiZrSRQLVTp0lQ/fAuMn2APm8krASUIY26LV84PZ+AC1
JDioGn6/ccXVHV5NXebS1tOJgi1UJb9tH+JsAmOVLlFGruye78lqgEj1ImCm7GQ6
ghT8qUT4yKNBnnEfNxn/2tXJbPAlH7Q901JC6HL3yj/5Exy9XeswWkbVNyESijfQ
8Ynj/pf6suSdFbQn9uGwEkwMyv7A87hWL9cIVWue5anKRoxxCAGylJf8zGCqb3nv
vTMtMAzb+Y9nBHPIO9nDqxWjQOCJWg3AQzY++l1pn+mhxe5fYo1bGsGuBd1mlvtV
Jvqyhi40ly84dx0eptEDEaebm1Y+P+Eg6mxbkoqhsUkfHDehKbHIrG9amylukmXl
lDkIAK/gGaWmj+4LdBXj6JVPLVhhqMRGvaaHtGengiwM1tPj+IT7qQ7XvXvvBJmZ
jPy1Jwv5iYBIi7l4vp2Ff/WtggKNO6ZT4SrjljnMWIkZXjRvmVyzaTZeyruZDuyK
nfYC6day0BHf9zfukmDPiGylUkFNRZ7q9XVzNv9r/YDJcrT9QVht+puYLsEYzt5p
8urSN++DGthmXOarwLVIJWsFRrWZKwIm6L6zhHttUsKCccidLcWdrxeHFJqE9hlN
3VphEnjV8YZ8u/RfH02ZA+ba8WuGozpzVWI1jSVMU2TKphqampWj54jTy63WpOXu
g1dF/TF5cx+Pt7AYT2e3mQLKJob1HJu1skUyQiO2kwlgeu1M3SCNheMeDiA/whCy
LKfduSRyyAh3RVqpSLEabMp2XPhIr7PWUBVLRBb8kY/fxHCLefEWDzxFpjfLIauj
hmsCF7BLXGmJzp9nbKJU0265xyZc2WLyaSwTaeCi++VnX5LCx+DxmwdWOdcUkrhB
zWi4ElFT4bUMm++TWmEi9I3TPlYpehT4zZyDZlN0desp7DgEiwtRsDrztgXFGIcj
yJP+zpC+v1yUj5UeRZD3CTVt+/sxm60KSBT5j0XzOigPb2HpjVw8h8FfEutG7vKT
35gClFc5NOM5MCKG5Nwz+QlJlL3Njce7mAhOIdwohDH7MywSm0n8BV3eZxKdaVF+
kPkem51pmoZsJ2kokcoYjcLX+GadnKw06H4ksvWj2C6FawQQWKgCL3WvhQwQsVVH
Ddak1VDCC74rgXkNNV1zXpLcgDndxcLvPCPJaV5kNJIlZ5w3S0WB9woWCl5cPNE7
xk1ajehS7sU2APBhgdA8lYlibnJn9jT+I8HqDPpTqVRp6SjMi5BO8j5/jzNpt8ut
E4C8RkrUXk4kTbQ0DDqKeQKiZiK3+KZJ5H63pMIGX59MZ/OMkKBTWWqbYMXs+52D
k+xBIDv0Rk/eeLIao1VMkzYMkncKWklME7wshXiXQY4SYbOisgBxrUdXcR7ibIDN
lo8NSLE0S70Ckw9B6CFA2ZkID6N+lDEKhduiiu1XCd0Sx+j/5E7N3vJcIe8plU5m
1v6njr6R/pMBu4gFrU9sxWO3xJkZrjvcLL7XTKwMgJ4sBbBX6SyajzQ2kcDQnSZR
6as0+y5gqQgxgOZI7ocn71jsiBLyL82KWmIKvBkWxVoZVYUQ1Wbi2YEoNQt1ui3g
PKaVHyLxU9iwvrG25M7p9paOxl8OdDHRrUbJJaZ7gRBddmxb+rPz+qhDpR0/Gt6A
h63SZDuLVLxfYe8bXMpU1SGRMGEOUgaNrIS8fyx4iH19noCyJdcsD54tWycMNKeP
baAAa5FcGYWEqfuDptaNi2gCGtRytqxhkbeOBtqktipCybe0LqUrQTRtA8ey3Yn3
qd+mS4lNFuQ7RJq40lYA14SynZk5FdF3tTlgdL7EIGs+1ln8I3cmk+3LC0c4DFds
9vqJNyobzKahNJExk+CfqBD9+6gKzRyzAE6RxEilSL0UIqWJH6JwIJziXVtkvumy
wE/pBSyU8sdXzgzRAgatIo0GE/ABZjkm0TVPpmXI0xta1UKX7dORZnJ83va9ZqcE
WbYEQdoJnVWWHb+FJfQchM1Ci2WQLuKCf2xgorek4f9T3/tz6yBrVKjcoFYQfB27
wo45WbhU6XzVZS5VVvzMIXmEC5meJemQBZBOAivIX4v33KbwU5dxa1GxbkmZtZoj
5veMBLzTJhkNjCS9pQcOZv4O+qh0CexPMc6QYiCjzTE3pXYgVvPB3OlMsV1Fe4th
MN6VdSdQrh1fW9N2p25pNV9afqD4xdacs70Cg1Q8JGvPee6oPXb6o+cZPAttan46
Oa11iHhjF2c2VJok903jrb9jzNA9fRPNjDw7c4botTp72wfAV10ut/U4Nta+imIX
PYAZ5AYh9O9m4bj2ZQ1j03KIhYC6/bNy+Hjn8UoOuusC7LC+A/GJR74CTQS2iiGS
HjUJ9oVo3N3V+WSZ2BL8rFUtRJZBaI1vUqtOZf971ni0YvnboxBeh0k3mQt5ud5Z
Ym7iesAWigmZV301ZznXO69SjSDtAxr4PM73HgJ+L26oslzl+xN0FBC6ChjrvvLU
ocRIaV53tCzy5tkCNHcJe7bmxQLmy08JV+aD5SHCiX/QCUFtCMvCpduVY2b9Z7L0
IPEeQnFmWmUw+cHTnDonO5C0/6gnpGttXgtyfRdyrCv1U4MgmnGZIA03M6gcxOkA
l0cqT5Uy5rEhWB5RRjeuV6lT62lt++CaAp26T+JywL9M5oVsNDwZcdnMP3SoFHFf
fFnwiq3QlzaZNfvqaLtJtlJ4woXDyOhVHwEMQ1yM/K18U5uk4QBr97hwy6oSA848
1FIeesbpyQIzhizYsbDej9buoPsCnBoaQa7AWM/x5aK3a+VjNf3PN+EdOLONCqZT
uD1spnDO3AxcUGYZkaU5ky9QRt+EVekRdxlt2wBjhu3JrVLfp2ChY2ZqDp13OQEz
pIDCUTVfdYFQ6cnpLNL8EbwknhEVjL4mKlZDM13r28ulEfdz6yjg9oe50SO8qNOJ
oqddodwWABlLKCi07AyL6nSl3KtvCZkT1r527tOGxZXN1tUb7ta03KRYQ5M2smRw
ptVhuv5cUT9f80vmtFH6bRmNw6CM32/XAHoE4boE4cYIDimVukvl2q8pqdhWp6uj
//aiSRvBbejR3GAjIIFnjlHxEdxoWQfkZy7B6kn2JmVAy5IqKW1xq4/Ff/4eI3Gi
pwoOlV/1X9X4F08NMlerp7co0n6FQSU8AEq2W9jVqY+OWLeF1FoJ6Tkh+RhRvGNN
a+lneLcltO+wF5NiJAWN1hZu6sBF4L7hiplbwUNYJvkfk7T0gUMXy8aZhcoWOk7i
bFDDqJAFhaBaW9Jv4ViCuQXbBtMz2LKFVmv35DyndXOH4NiXyKu+AaZ+y5UA71/v
BSoG0emPMZ1E8LIy2zEGs0cikE+r2skYKUB1Km1ZjQeDEcxTr3zqyvEaNZYVQfIG
aYPSr1hkGkC29sYOrhCbyNtHXEe2NAe0das6yhPdHj69QyFzn//6IMGjehdPCW3b
k9pwv57VywecnGAiUuWaE8S4CYPD8fYI+i15y8tpWILr1wUYGiImqhpuWtA0KRjt
E4S06vMYgFPl1qQBJMVT7VVpE/JPK+y2BItNiMLpDwJQFb0zer1G3IkphziapO9u
b2QMwLQmKrxHB8TBDZbhXdwVPlTvzp0xbhbVs8FaY8HT2k9wmE0YRjBIn27Uu+ie
mXwjKIvUer+Sba32eu15OgNKZTvsXupgvNCk6aHyuyBi6SPYObREZK/ThW8y0mr0
OAJt8+tc66dwXAhNdXIv7KGkVl3G1z2xhcooZqmMZWgVzc8LqsM0VntrW3lqX8jy
qJgPalxle/W4kPknVG8mqBf9tOM+m2n94TazFigBpUPJbGjtAfRfIH7su2asnXiz
3tZD1r/9ySwYcyi6M0faDOkjpFoek6M2SrxXXZiwxjoCIPH0xsyjchI++O7iCP/y
AuBEC1FnTYI2U+/vNJp4jZ7dIwIxkZBcoUqiSK97odFGD+ZMwcObwLLhDLlcFuQV
1lKJ0aJ15Fy6a75HI9XXv/7Ak5f/UXaXY9YFdFjg50KwlTYNNJrJ7O5Uq8LbsjGt
gky4lMp+VKjFadLyMcegEljAiPxyE4UAuRa2v1E2K88opx2WdiSWslCiSXUdPZeZ
Mq29Efpf6kpEO5aJWnGFTca9PnltX61+DHEUPlRhED4arTRDnAfXIH33PLglQwpL
n/SQweproNfezLrC2JyMIfQOsBfpyAjvT62DUD2mFN94li1wRWkSj1READAbNAip
/0ZncKCMx6QmT8lOgIEnBp7IH3MionQV3SX1x7GBPNtwsSUcD2+kmoUFWL+IFBjn
sD9S86zU0JHjOj5wk+wt+yy7qJeagqiM/mJZ3i/20mxhpxkmu89PIAVr9hpBI/vO
AD/qIV6WsruIp7DA6YnAL5HF+tHKvXKVgVYSqdHfaP4+a+DGziZ0gC6f9/c37zIM
eR8B2ZN7LTpWn4ImhHz6NmYVlppU+3ihzw6uaTsQfnYyE0TzrXIAmz5umr8ei9Gl
An54t0uLkgTd6MfvTzi3M2GM4VJGELfMQIa8RwdO3b4t7FBZOXM+3IpWloGqNDPA
mu8h6szzkcXa+ha5DfYbVjpIqjVeEALaY/jvI3yOtl2eSGn6mCF5WXtlyvpZaXtC
u/XUxoMNWYi2lHiHvnkA+jKDBXRlJKTRyUSHzxhqiHvMY6t0u1ZWFhg4zO9ikw/h
fpyk256vE2yiW38/nr4f8UIS8YwHqns87RvwV4fchCZCaNCMrkwIA8lztMlUmqcp
TrLKDcAmfWdtaepIsWJZ5qrebWYMnre4ylpkbztNH7F8A094UkpNpsHDLYYRaTrv
+wga47SkPwSwqhCoDkKB1TKBOyKAnVuEWff1scGVrXQXxZmfmXCKZ6Lb07uceDuD
7Xas+NrfpuV2FqBB5aw5lF7Shf0LyzDX9PUkxTscx8bsR6zTWo3hV2QqGlYLou77
yQ6KTvKSnoazRIE5ef8nLTqtfmwA1k7gVX8wIrLTTKQ6iBAny53RV1bLFtWN3Ga9
kwDauzHfkgb1sxl0qSDZ/6r9arqrwDZKsyCsRIttpSA+xpnisKwaT6HGK2J6vihX
7cPnfZa5EKOOYYsWnsYbpqekoXQMixKqsRGY9YDGrDsKppQblG+AXgqAhReHxqZR
SSFvVwZ6Y0d2WWvwzjLJ8j2rqOYx9kQQYaWkQu1EiM6mfOQd0xQLdUy1NyJuAXfd
6ATzrkhnpZ9NT273czSWz46YwPDEx/OctJDYQm/M9JuUnyUrA5ea5A1qxjn76Li3
ZWy0hUmvveJ0i8JHOd8VtDlChzSuNDaJ63iWTWgY5cj8+Zq/UdScL8PQFuPetudi
nv0hDxwOY5drmIEtD/vhCM3bSrH7eql/8VMkDdraE4ix10kFL/RgM03X651eMvHj
1T9UJWWA/T+6iYbNRog1Bx3Y0r5/EjeDPzWh5QfHkX4mZCvou/c9U6UZOs/JT9Qt
mxL+UsD1NksPR3OYZwRvQniaI4f5cD86gRkZAs0wAf1eGSiyQC/1c6bYoiEwwiqj
HAJzPQuFYcW/AXdMfZiv3GklyaVDvyytaoLrXRUlQh3wccpu3TXqQKLYxSC5Ri8X
YAsRjsmq7Ev+mdd8Koe7InIH3roICTzJCV/qARXq7jupOjY5cTBXp8XPnXTFGltv
x1/wX/RiFE06E1rR+rwXU7cfwpRrryE8oVGyiVagrx9O4mbrVsxCt+rMlvMoOa0n
c5P91RF4rqx4t44DDB+jIrHxk8fDNFo9VPwNuOGJYTnh6uTSkjgVSBpLcu+EzX3i
5NOtXOkfmI2gewv8hwg/IqjW+cglWoB9LkdG8FRKhsCVgQaCejoOMF1pKW5Faxxk
cGIQkvpXvibbfDVX/QOcu2ZBoeWmYIYRARkTQ2fOIvKXxPHlg+63XM4+6XrEqqxD
x8LZ3sXgwytN3HyDmV+PdhCKxuYvf8g9cYXPkz9XTBg=
`protect END_PROTECTED
