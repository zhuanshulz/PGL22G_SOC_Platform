`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AMJimhnF7cCTQcJIFNpTNjQnFu2fjLoFRaXFcvj44PujNQIdiAILWtJYI3Ih9Cmb
8pEqxUDgxZGijCbH/bIjlcXwvxb4PxDPrrSoVvqiW2jZF/qu1rCjwlu1b8R37c1o
YcukMWeHm5TVGgz2bOwIbqnYItF435SdF8lGcywUkWZR+Y18QfvTtwtZPTG76LOw
hMTpN1xuTqqPp1nItelg2NWNroTtutEc0fDSIiCgTs78vc3F0soZi4iYY0lmNGp+
I3DBS2aZktdU7FVfSFxSXIkMNAS/UzpitTAbPR0IkiCEnlzH6wXfZOARluHi1ary
L6eKuCjGyzxKwziFTC8tioi5dXVqIHSubXbzTv0OjiE6JSzpuE/K38zL9CCGvSq5
WChXJgTSd94Z5HqvVgD8FlUH28fBJeo/klqgOo5qlJ4u/c34kqcMtxGIF3vdl6Bc
AvORSnaaAK4DWQdTtQOYgHV2QXefr+nvWXlq9szn8RQ8IKD4NrLr6F8qF+HCkFAT
hypUbV381WoGcOpfTRDjh0XD275vGza/j2K1Fffuq5+soJCjb0ACP0ftcpnprZgM
OTG1t2k4h3c0diPuhW+7Ohz0yVf+HCe60zrRVogAHlE=
`protect END_PROTECTED
