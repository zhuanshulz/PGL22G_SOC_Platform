`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3vrZ2wy7t88ZZqzxS1qtNSS2dSTnez2N6sra+JLDtcvnXJ3kx5lV6nsGQDj0Ve+
sigiTiTticryLtO7EHi39QSQ5vTnQk/YUpXm+rYViTS/Q9lMN+esP3lSa7f72Ntq
r6oiIEFvSRL0FjsPVXcoPHcuCeu1S+Bevy4+MwESpz3Hf+kPYwCjTaT/QMjRnHLq
4HSk29dZppqmMNN0HfW1yFO3ivrn7TcI0Lqf9b326TqFYplQBk2jQhI0bzT8rodZ
dC7s6bgUMWI16/AxUb6YUZayiSCbxUMTFl2HMyM90F6Y5ELHM/c2Rl9U2EJ1xQo/
xLU5cEfnqRXf1Qo9cKQMBju2kgFxVPDnPBxeeifObTEhpeT1WM4jTv4mFTETUXKV
cRGt0vgHxMR/JNuExr2CiNVH5G3s2naEHmbmbOUYgMBHJq85SUi+tk5UXxM9opjz
g/OYUp3Ej30Xj713OnXktIi5LQ2NggWatUn9gb+3MABs+MmupdArtejDZsvuG4MA
EmpSWDwgqmN6dFuX+hlKM+yV0Ajbf125y7Njlv+Hp2aJXBzu3P+bJf3fsNRHr9S9
r2Zy825Njlq+Z+1XTjYMF5vShw/oquJWLU1Xiz5vMK1WJUl+cg8GiGexRLlQyh+8
Z2hkVkt20xhXKXK3qYTlGJGRo+g4jn4u+eXo6ia8UAb8XjscRwXMZO2WnCXnylsG
JaT2L4RhHnifJ/seRXUM3stTUBOd6sBwxlnopPG4BdCbZuTOL9nZskkem9wmXBKE
eZ6LFlnFOQY/LFGfjG2x9Opwk3XCar7fug6d31p2eHEbltCZPIDLTTc9Tqe8g9Tf
2rRp72RVCW8++3sKtcTIjBUIdTsfgsenwHE5gZXTlmMsXBQjfHnghPRtawokvOtX
CzIPQEwx1d7GVfs3i2EKDGGhLDy8G/2vl6lqrSvZGvP7C5GVOSY7kXohJtyHomWH
npYCF1ILH7n4N5XoL8zw1fGRMI+51UAjH7qw3XZNicL8zQNwi3Xjmsg0gPXSS/JD
EEramF9LQfZ29e4O3MVmH+W2QtO6S3/WNAar9Q3cZV/O3juQfqhcEQ43CEoe4/zs
ahgPVDL/0LoiwVFSwKFkks2o696b8tz1l8csq3xLFSyqJQWc+w/IBm0Tn3XufJNk
m95CqEhzL9WmG6ccRpRmmoxHJeL+a14aZFtV5sFZ01yDzLdq+50X3K3SUwmxlm9m
ERbIDqdqCVYOyt01ilUI0HJ9rFySZNxh95C5MKODCZAQ3hfhAvY1a8cKzW5QETYg
p9BdmmhBX4RY54dS5gE82F+ZJdgD/qub2Ipz2AMTykPALZRUELC5m+k4wpXC7xoL
VbgkwBeQP7liDKxcPrQoSZGT4IPsNcF6MtTZ8qaPoc+fFfhK6ogVInz6rlidFp6H
ibbfaChaHqb3htR1zt6rFQNqo5CpzXwHw3ZFFKRMh23LvjcgmWFGgxpHBoNO12vq
Hdi2eo1Jk4z3KmzAKqhkU4l9a5jDeUuBYb15flmCGFjLCT98w/kgkjfgfv1MVhL5
hxylMyw0Zj7ZopQ2zLqOu4IZuWjkm7dJr8oh3n0fh7npPVBjZBb6RE0vvjL3NtAu
eJmAB7RJzzV2MlwfQ5m2UPSmSIooM4ZSVnPBIKi57yfpRt7h92pmre3ilOaGuhvR
WnXy8jdvHvdwVXSdeFHzMOtms4rnWuLJRDp7Cm81anyMTxUZNIxIcSg0PBZRRSDJ
xKLgev4aWQpv2k5JAK9K+ytEJZElJ2YHrMfeTANOsxLD4J+aULgy8N7FOBjeJ0Fo
N8ZIQLb4k3Aldo6hTR0eFGeNc1Lqz22E9YAIyV7Bv3fewmrHJ1AHJtXA1sZIRM0F
EfbaOjVems55J/S677zkvrCPupFHsh+jt9CMjS8BPpfDqyRCN3jCY7LcW6ydz+BP
j8yovQTBYkn4Pq/GbIDHWcyW1bdSJKWJKjJA1EvFB2NGEpEpY13NndJp0Bx3v7Sb
jXpuW239613NFBN24fC+MW3HP3cW5vLwfsCPRFa1ti9xRZdXERV74QiFBYJnFKN8
2WzCVA7GDZPaNaI7hUoHi5SvKzn1LULhHxdAy3uipJI8mYzH935o5Bfj9APTiECw
O4DnwWd4DyBTclxyE++fKLuXx/64CBO9ocvVNwxXGgEgRkXIQzAtRWKETCRc8eiQ
gOwGqQRq2XcRi11/OGNjnvs8LE0aW+agencKN06e2oerydCMdcrGC2CqeA6YEDBy
uFmLwl58pZcw7/jhA4z0/8hTvGacyu/Hv5HL7Tl+7EkhOC+mI1M54RTf4gCcAqRU
GNzjbihFiCG6BBbS0SQxDq11bAE5VyFsvqi8zVW5anIxD9XsaFUFxInSPs1tHjas
yb9gsB+2vj+ctRx1npwkIzK2LEaDQLrUHNxBShL2AXFWMzqMr8pCr1o7927mFF1R
YEk2TPNoDAQOJN4FtEfDo5S7/qpDxERiFTnUYQe2MWQZ6JnIbkHUZrkrWE92tCQs
5OzvVTM7/tOnfQc9Y87oLi0CtdJyOhO+84fKYeZbZNUSkcIoOWT+qPwxEEaOjIdR
SSiF7/JqJKYzEp8nVS1VmyaSXbeZov1Wvro5q883IOqMG5FJqwszCkxD5OYlHcTo
Li97mjPQLiKxRmkmL6M0tOVrazieNHwuFtuGxwaBy0l18vzBAeComipUtUGz5wf7
0D4P4oMhOOcfhtH/pT6Fvz5xgvJtvtabRBkXZxsCpvJ4ttGxhd1g4DGZ4/Wr/TdE
ZH6eEH4/876bbMynBVD6pg3b+NXG7NoYvQaUjIhmAPHUOHZR0qYIGeCxmKJ4eOuH
PG54y3Hi/nuLTlm7YouE3ROMilAWPD9Eew3uXnVK1UFGShTA8O0iXvBgr6timQxQ
+gLgOjmInQEXmcUzNSyaeIO8UN8AAz3FSIuD0caWcchq8sFYIia0cxXRCxGS24qf
OtwooZP6SWz8RZF1+/7GZL/rRQtp0WOTOw5YgobZqqtYekiSW1A8MIA1h/juoL4H
wb5l752uREtD6AxDJLBMmggjZafu5/SQEhcjHAE8CsnOImCQ31LYiz6F1jGWVbvr
EEqemeu6CoCdKT8ZDlQAeoHJjg65ZOQT0l/NRAo3Y4r/Q/NCmo/TdgcSSyAsZTm5
n6OQo6yYRm7pS95c81t8WIQ7ts5pSbxwG1ncvSnXZ7GGhGCNAz046tUe2eCV9eUf
5J48SrMocLyEECbV3XndBhuzPAC8QTuj7r9QMQF7UOsx5ZGqngicTj/F5+RkvI6e
UOUPVUOqnwq02lYMCqCk/vA4N/hH6bY99fW1lBCGsLMiQsEFK0oN3PaySdlMRxor
TmRJPb6LuXT4BCmwhUMZVxPnei7GrPMOPnsoi3VBhPd3Xa6iusIOIgtseTmNZygT
XNHXZbAWKQjHB+WlkEwqSuZU9K2PHqtnqNSPENHX62lmGy3VJ0oRaHjEomcJ8I+l
B5l7n+BXJX7qg/1jSQEA4r7iiW9L+qIWpRWdCCDzfsiBxcIWd7GRXYGCCucl+qom
Anm5IaaAb212C2wNHPilspGbmRaNAP/e9UgHEztRQeP654WGqf0LztyZotGlc6Es
V+iqEQ+EwIKGgQ1yRAJpDvEjyQKQ7Pj+JvU1jhMKRCK1oGUlU7EjxmlnNqBiF2e7
VNA0mndiQwWZIH4mHpMbGp43SmZjs70fcMUSBOhwsBhLQm9HQ8aMhxrvRBg+yPLB
A16h7dw5KxUjl2eWvBv3H8q6AoPqnH5TQvhKddyKwTXcJtV64wuZTdvOu+qGUyWK
/BRwYW8gSBGf3pDA+23cmTcK0cz6uDv+VpzCfbe1FfPCWUlSnDqmo4P2rV+uofle
tThY58HTbFvu45gKo/ARYnVvGNeVC99CzRdaUUiRVSBwxylxrd6wRG36zOTuyJrc
BFM7LhB9/vk9+ckhq4J/Hb4Jf7KE/CqlcUgloNp+DIOSQaL+Yjf0CY56yzhZhmnB
zr2UskVup2F+oHEowViWu+GAOhEkSjppAVKy5SgYW+swSrJFcob7AUvE6pHcB1oF
T5GeaAAGjrQl07fdwF0GJcYjV/qWJ8n+PbGP/JtvygEyA2DtOTe9G0vSooS/+G/H
PQpiICDGIm36C9/c8siO92N54f4S18JvyLYCK6Aa6X8Fgw/J1fn6C4jOWsfxrjWy
j+6rxA6pVzq5cPrvGdUk8Ml0nzISmMKZHNpbxCq/2Pjl75GEwE1OLvyAfBDbVj2+
`protect END_PROTECTED
