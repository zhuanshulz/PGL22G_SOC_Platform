`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4pSF2Tz/m50dh1mxepAVKsmCwadgb9nCsE6DwnPzGvwgqKm5oQUPZJyCJVfYXGw
k27yOg3ZxsEqwRQD+SHd9RVVsb009b4vzyBiL4p1IsbbUfM+cSNv41IFcIdCtJoE
AS2QJ3YIlJ0n0xpuUMqnj4dk99GT0avnp0hSg0Xhgog1zTDLj+v7IiRDSkIfpaJs
CQy56x3rmPuzUvGl+eJ+KDsts+GnttYxDJVcH0PKAWgfsJVOAVE2QZHoy0YsVO/9
eJg76nLrcxSXCYa9z7A8b0/yyxBwd9ZV2GIH1HVhah4rQvVKGUIMQkrVEUOr3Fhv
8nild0pVNGbOnNCWpKbpSSy66WOwWc99A+5ULDJrPdTR5LjV3MmFvFUy5doQaCbn
Zx346Pw+io/GgKUJHr7G5eHn2gRWn0gLNVSfAmwXBT+eimb5eQ/VraP1Z3AR0ZvO
uYyDcIAgrYSt730VhLgLM9tscZ/GRYfikNCe2oZaN8uaxHK1R5Q7yOgArBF6/zAW
VAMWh0LOqoaavRVwG3C6dMZJ/Nn700uzl8lYL2EIC0EGm8SgKp3EFQwx1QXkCzCm
9Da0sikUfuoxXWZJDjJ+S7H69Q6LEBXyny7OTUT7yUQ=
`protect END_PROTECTED
