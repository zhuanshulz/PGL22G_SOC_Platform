`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S9btPBvBSyXySf0Dlej/wAD7sqYDOcZM2cx7TIA/gudd4IWSfGAKojWXYVTPr3NQ
WoUbP0nGx3iU1MmNtRm2rzF1xkp0xDOHTjNpsVXxUmeIN8hQGlltQOQU4uqdx43w
hQyj57zViFW/zfdtqcOJ12hY8TmpQhBKnrPdwR24o6X05j+/dSbNzndb5WPJHLsX
NgE5gqcUjtJJhhKFCnByeaqVnfE7eVKuvv4309JLqfIvd0e9MVmaSZd5I1uzjMYH
+gwzRDm8gniJiNnflcXUk2fc1esPY3N87nzwuLXWjU3K74coNqE+kHhXgLs0VNlx
HSL/Hec2TabnQbgd8/NRDVdCNH4PU4uZEUNSPoOMmNjcdtr3I4e1EieY5WeafDEs
hL5GO2223HXTjYyqZUREgLe8mT+KlknsKj0cD4R65DKBCrMt0DKQjsl0xFbJTCHs
HSxZJoC9ENtyJ44ATDRp2imBGEcCtGMGz4bzzsrI+9uRO8tVDXVvCZT6AyU+a/k3
4mx+cLF7Xzdgm4ZVWSMkTcxlmo8Is0mUNinfnFv7BQCYV7lFKATkvvi/dLBc8T5S
O6x/Vad52oXgKEstqIIjiKbCJZRbIJqY8smr0kOKVDQ=
`protect END_PROTECTED
