`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WAQOSBCXr4ZEvJxWV0DTnthnXdKjvuT+UWexYKQ7bRLJhicdVpFd3z/5xcr/HcmT
SgW5pXq1zQQYYcvd3Fh9i7W6xBN1bOinYlq16zBzR3Wot9gTqXetugskhY5e1HPa
57Fn/yUh6RTaS5sGRAJB21z4A5PF2q2Me5Iy9ciBrf6L6FzZOPRLwMOc824cqsiZ
8sK5M+U04VJSGbnaBoG4AmegNhOTyjedb+OnkCqM1rtaQruLNSBEpNMMaYneOTIZ
Qnwy1cP78ssX7Pk2pjamEM3UvyYSYbwY560n9aCa31OTnTvG9nHBB/jaoCFUGl5t
M/qC53YHpA87VkL55x6nhSqF1O1raVcBgDJhSk3AtyXNu/yTC2WvuFRLt7RkB+IR
JklcONbkPCCLP0MXNlzpmjlGOCgIYF4ZFyoWBpgFsSOmatHrtOz/Z8vMDYUefH0O
1P/dG+PAn4b30m+K6uWjVCt/AUU9+srAWrtLKiJQiqinHqEWe5nan0ALho2nxZNk
/eQe+aViQF6IR5ef22J8aXIbSFYOJ5iOGJv3WiLKkTrrAOpqelEwfeyegD1lLZnX
oFxaKTqoo+wmlAlX8nd3YDQ84ZEHT2fdWf51X+6Ps/tUXX5CBOTpRBcN60AY2LPv
yD+7l3QkfnV+XtWyTfJU1Lsh4bJuBgz+PPbVBHT/PlE2+/arYbFpXF0FJukRQ/TK
iAafd3m/oYgEvbm4bTqJzaaZe0tf+M3/fEy+CZqFrcKSbxpA98ybvQZaq9D3e6o6
3JXgNPz4T5alL59SURCv5lV/RyjSRGNNjpYwlXa2sqOEk2EJgoSOqjq1dO5R4Zo3
XTDYH9vJBcyN0gwOx89KQes5QmqS5nLxRuXXM1WWZaekLIfnmvBXozyXH6fxIoUV
olr5KiMT6o91zH/K//OXVgn5pNJgnl4E9UG9uB6ZqUR80jxEEK/ncUAnY2vztJQl
ELMozBva0EVisTfJUjH4+hmB9oHAo1wleFRyvnmC3coGvJWnQ9HYjTPX57ry35OT
lqX5L1IdG9ju3CZq1Y+jJkIr4MM14mV1bU47y/9ZBDXSNusDvC5X5qL3XiutaHBk
Z0d8SWBqFte64idW4PLpMm5ViKYNjElapqVzg/Tt66sIqr2hIq/uChtAmAEI+P/S
qRPtiWBYwTCkYgZiaPEzi2rbxVwjP1YEE+p7jpWwAGeUpUZiC5/WmMRO7KN1wwIq
HVRx3+n2z0kSLP5uFTFJmPCVDQdJscL/TzXmNoYJRFpaIzRZz2+0uMsof+4hIdTp
mvV6GY1lTa2qzWIrq2mSqrGrm9ZM+Bblz+FE8p9gYXLof3iALZj1V1HPU2QlzfBE
e785ILNCbN7anaX3EQoNWpZ3qiXiWKq1KnmnOJ6viaJpP4Mk9uQg+L7dNLu9JWRy
dGY7gjfU2hXoEctem3jRRBC3vwXfO6ecqvaHV/IEjJn9MUHfaOx2dwolLkIwulO5
jAAL1iEr6t2DboKTvnmmsRs8CHY/rE1fE3UUj+3pTkUqW542qfZQYFAejUE0+m2d
sZD6VFU8a359O6Uy6qQH/Q8guQwm4oXZ5CzyZyfC5E4roGN+i93GXiwepXDOaUY+
D1e4n0uNKNiJC67sAPZ78P8g5p8QiGrAjE1kISfiG4esA3Z4+jJddfoZDcD++Yet
HKx/54UIO+HTqLb+XJD1wf90go7UiKuPZQIRlgiRGjsUojeM+DLGxdu1Rnvaoj/Q
4NDkomCBEtKFeYztLCajUgpRmLc0DRVX+sikCetxMNmPVTiqg6NnH5ooDwOlbsqx
/snNWBZD6zPH4htQiLyE0VUY1IJx81+eExx2yXWegBsjkVlcJ3Y0aLWVE6obCTO5
dPOPxTEbOsIEDMJkT0ZYFkqAbhhDpu8X6wFhK6aupF9w8zSAO6YDdi+VAVYoX0aB
bdgoOYQwwVrN7H/A3VS+aefTcYFIC6p8MR+NsskxsuGoRnMgpZ0PseJEgA5qAy4Q
/JKBmrwLNnboT2FIfbcVx3Sy7rbwgPFeILZdqReHE1wu9oDmOUgU1YTptXLEENJR
1CDS1F5G+GUvfYtjw1s41o5A821159poFwqDRQ3gDOyAu+NgbPlDmb4ogdKpOfJn
AFCZ7IQANElJtrzEh0uX7mbhGmaR+TjstwZ+MfAArJxxCNNiIPoGn9L2ZDoWgCjs
3EG7bVUnDPbw2sv0JAzQ+82LxktPciUts0FkpnnDB+5O4j89AKcicuDjOtXXj63t
/mBaeseGL7a5ih22cZe3ix++2iVBPfJQ1BhBVkRO8NRcqfdrb3kPx2B/g9DfL6bl
UmgSn5s8vOUAFVQao1Vs1rznT40wOfKEitLZUgfXGaW/9snrYiB1vvJicQ/4Au7j
iK1O7WkyCat0Fb57MUscRuKiCr2UnW68Uuapd6aFrEVhz5GiNj5rbMzaIfnQedkO
cFxiflSt1WFy1IqN+ghmmhvZn56TeNRCcdlpVf56bbhdPDFQUtPEgj4D/qygBypA
28w+fpbCYnsQvapDHc3a55EimIsdPZxGo+BDbM08CnJcAfAIrCT5ZYk3SeTtYOiQ
JBekfCMjPKQ2saHjRLEGoBQ4yOXxjl2HGW+GY9S/ULDi37VgrRr4TnPsLdXH+G+4
CBif9ljPUItiAtGw7TvZesU8bIE+iScKWBgJhnBbkun7KyoKtrJAc1pO88HkBUQy
c5lA0OeacN6jW5vKnKrX0uVDl5ximJstIlCpCul+oSbjDRqcMPid+I1ATX5/KNZ1
gsX+PB5tObVsMJOOrJs8IDOK+03tM5V8OjeikEUPutRRSR9WLrQLo7/MAV83Rtd2
JNLPPjkrRXNkkLMjmsW0MAWK+rlxH/q8MTRnnQukQiGWYwlXJLmggBvbhx6IGdRl
CGr5pIIV1FMv/Prsd8ehC3gq/jbCmcpcUkzZrRdzfeI4PhIMDX25CW9/ldYVWW4L
cC9lMdI0Scr3Ez/BST948mF2cYjSUzRUJNTg2XwZzZPhnK7GfwJHvrSGMwDvKpEw
lGr5yMZ5fDe9x8u6E3+StB2bR46t04QIf+taAk8TDnrstEx6o81hWyW+R7eNDWGy
joBcno971n3dXsfX68wbGH4nZKOSkLSnVH6+VT7YaPAiKqMM5XkKUvhU+DrJW/x6
VSpC5G0ATg50Wx5LCFmzHc8Wg2/fZgLW6ZhnkJM7CUmjGAgvNskq0khPka8VhgKc
c/egweqAMAR5eYebMq7NBWu2HA0EQd5ykNl1LDxVbIfjFuN3JQX8oszGVJRnFoDz
Nud7cjpQQk8oWvscp3tq1+kX1NFYbRIRaJOJgcDLm1erkHaAAIaKiggFkc0hnJHh
AE3G6n8rjc9K81ohM3QrtiAzNSdN0FYLP/FvSnxyU4pHh0O4JP1cTQqsdPNklL1f
`protect END_PROTECTED
