`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AOJ0QyXkg6rmeWmnEkDYTF2c1MlVp0YyfwjGz7QdFGwNZ4cT9CrnlbDBa5SjgNkr
sAlJBkuVIPOnw4P9hWDCu/WCfvKU2VhF7totcl4jhcZGkUTJLj787lAr9UXw+PjZ
OBIcSxRmY1zis1DeUwZnuUEhuXF7GbNGW6BMJXkTW4Cvqj3JFUP3RlpORh8q3yZc
1QyB3KG6yR/tKrLduE0Wxp5gvjQdORM6k3dyIgH5sZCvAldREVh6+QmuHdwq3tAO
zbMXtuLukX9MekQ0U1T0BJSz4MkjFJEk5CjQWudGxxHq/CluyVaJp4m6bi6DgfpM
b6I5R6e3E8vgOpWge5EgPsh+62zgXqRH1fQo45A0yq3O64vmoILjgSmmQD/7XwP4
mEzs7pq0f5XjN1MsCnMLh0+8yYVryNEcmyBWyaxVWkVMEO9SDpGig7COLOZHJM/M
JLRVBHQ+7ybY972TMdMiL+aA8r25wQMlR6VQ6jK9CjHpUO5DCit7COFgUksBZIpo
Yjc5NtqGeyXtxdu3aW2bTXO/FvDQPai6WFfopsOmYe+q7dCNHD64jN2IbVAMRTkg
U4ddaQ5qhJCpLx8+qw6m30Hl9qXQZiqB2/aFQ7iZ4XcEhHmkpcLWEHQOKDq3/Y4Q
4wk62A/xJtr6tYJydy2Trf9g1KtbwOqAysVAIGXuRaMlIqY0ckKVue73Xk540PUJ
v9/4Vef0LGClNkDBpjmPXw7Vt7bJLDa1+8LJiqqTvgmKH8FA1TowHj7sXgbI61J6
QhdvarD274iP82KrNJMGnwntpuzR0vj05Zhga/kuY5xIgKLC6KW+a9w/40YeU8ue
3M3eewx3bu3FFNory5qd7hu7rRj0M64e1qXOedWO7JPekn+RarRn1uQfaSiho/Gc
RX72yfzklzYusyDix4hKK7GBo1gLQwsD0IWLFHxQ1BmKl5OdsFU1GekVe4lbDRJl
xmoWoyDsAJeLyARV1IPbKYKS81quocHEVanfHw2hB4s=
`protect END_PROTECTED
