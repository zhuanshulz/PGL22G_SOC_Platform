`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tnY4VQKVb4P/1WRRlYdxGQLsqSKrc7LYM3OO3OQsQ7IJhGcROSuVbU/kh/CTinfS
Ks3wW9iNqc14XRp2QamZdt8oGWOm5OB1NMOHWAMuPvbW/rDy0QHjMvLkeMxLAdTj
IfbMQ92n1eP+DLqfTOw/Rdr3igmu2+LNTR4r7iYVl2O6wFrebGw7IEuZfATloNro
q7P2iG41gFZqiQFsd6zCK0et3ejG5IbLvp2ZfmADnWd5kmncaolpQgFmMga7KLfo
PVus75gm8HnO8j4c18dEr6MHknYm5i1RxiX1zs53bOcprx6GYfARe3yU6WtEjBcP
nYINvVgQ+8lxKxsVug7w7EvZqgdeIAQYMmThPWMAEMv3aGi3dGt4J5KmqCZECPSO
W3Khoyl7egH2KJ8lmVz8u9i/HgiY/IZINKrmAdDjFjwLG4OkqPl1LY0M8I1/ksSQ
hHLM52u6Vh4mtY/lEW4BHEcGRytusRTjBY1LzEwVv4hBiSKuH2mi7uzEyQiLwk80
t/LNFUNA8A+IUpEbO8fKPKmq3h2vea3fDePGI2XRdR6YtyXjrUVsvgUO3cASZKaW
/tRWkwXkJ3wJSQn0ZyQ1Jd1Mnj1il6UV59VKBlca2xmRX5MBdqEXWB97B0Lq7Q8r
o6S/+1zYvVps1J0IibQ/YoxA6UcW1UamEJ+D6ohVOEyr2afnem03NSlD41szyjaK
+eP658a6K1fU9lDdFs4zfcSmA7hRlV91YNi0tbMdqhcWXjUt5ac3xlYFM9d7lELF
EN6kQSJhrceLeUo85HB1xr9k/YehmP+A0gqJ3fzUQQQYNFqhBHfwoZ/BdHYY1NWI
YbbyccsgMtLeQtu67X2p9nTQRY1ZDBu3dB0WtsuYUFXGgKYLwRGTx4ovGeRHKcYi
IuwHviu6LPoCG3jxUAk4qgMRGhuqnu9g3+WPVGJIjmuVsM3uXcJYX+VnglCY0UIe
CIlmQzdQ/AiuSA5nV36RJIVpjnYDaPpn+nLQ4FNBskzRgLZPVxk8Cggt9YNr8xaJ
EmNE+yG+VBLvyjjX0GMqrR9yJ5T2K56BzDP9oFwvnOrTPH5JmKPZufZSmIb8AOzf
WjIqju792poTpUDZibuYUMs1KqhIe6cTAuDu5VfbfqW5YZUYYVX8g7huwU7PRGtW
RO1jeYNHCcLcVvSD7BkbDAbSS+xSYYH/mU2/JogTwVTodDp6Gb+WdGShcXErkdFt
EKwclXOAiZ+fh/kdwW/S5wB8locsIlJIGrHt6Zs9I5Jx5O1vM5AL/b6L7Wosb750
vQZuS9R1oOvQ0iU/EXAXDNQEw05i9cZ3bW6kNqItpP1tezz8BUXDnPLYYEHZtfg9
hBO4Z/7i63WpCECSE7yCYWB7djLgu+ZAkTYnvr8AI+ZmeO74tZVeJH7x3RQgx/l+
YV0sGEPqgW/YKlEnxt4Fl0V1lmg8CZM9tz2/be6mfidm7dEv4ilBnDDHEs+1dIvE
/APQJcBEocP7BV88YW4hdeb6CBhmNvwllYoZpzCVKvHNUqYNIfTt5QdJXXPAvWSd
n7dM7H6wS7BY0cFr2NgBrRg3P9Qz4bRkWZSNNaMKyCTDUaE3oERCcuCMzrDmc2+a
OzScZnPKP1anHb4X/2pWlt1D7KQ9WRdTXvCJdvlSBjGY0ZhX1jcnGVtMDPg5DCFZ
SSkeoR6dWB5Rc6JZtgRFWq0YdcyrSBuwqNckgaMvj1NK1xpdTlaIGDTsSEeR7xQG
bUbej5tM4cr78Go3cKQSCO/+wsX0WejOQUcaOIF/CmlAQ5IvIhvfsLwrfzBpGq0Z
zpDslGvYAAEZetlO/T8w+Flbj3U5hg3pbrBoZ6ennK4e52RvxD1vlWa3UHmng4Sj
ZsbC0z7l2JsBn2lXdxATtqh7FpHHs28ziD0dIF1G4COkyP8ZeQEDcDiLZtsAns8U
+QablNv4McJPkP818Aq/np3uklyB0evewPJldzg6WDGGdODSZr+CvAEI21L+lWn3
gZLhv2BXanfPhMPVQKbLff38yfSAuBpBTM/5jZA8amKU1v6Y7SPyawWx+T/z9uJZ
hDZWB2BLIRTWtwmcULxYyqSDr6pmVH3t3sPLm+ezjLVmaXIFzOFv5ocGbNN6Bxe0
q+nv8cK57UG2NpoIanseAa1RB504HQA3Qog8xtVCSsoH7vr+OgcKGamGZ1dCkKid
5ne3mDRf/bH0ZMik2lCjbzfQhizT8L1ZfCbR3NnfEaKepSBJVH0ikxoFIRgOEu9m
5Pm/PgErhpbAz/vf4Ex4PrBK+QugQxGxoCX0XQ/bxU5s7u7KtYw//CnUzXNz4Ler
YLc1PWgPxymTHlUNjciomXF1fOmxFdpwQBjDfTmfxzvrY6EsyMebGHcvEpe4Gv8d
UA/HiwVJHeVyhAzCbSE4Hov+vYGs5YZ4XMg51g2hij5Iro5f21A0jC+j6dnpqTky
nm4QPLpp9v8H94n3+9mCfCbTYrWSXCHO1JlZXJkEEL5WawSrq8FvAWMOv2kHZCFq
Zi1iULy9NmTIMYCKCVSzNykhby70p5iMc+a3DzxmutS9Nirt50CG9V/eMPmGGBRa
1vieR5DozmhIKhtWV8JYo7iW73v1BsOZVzhrHwdQwUnz13D1VtrOkpzEyrk1E9gO
rMG/38oQTIoR3IbfYXk/03yWZOkwnnro7nXYCupTD3fy5LMM2rrR/fEwxRs/KuAz
uyeUHR7fP+ETnqkJszBglS2MbvqGTDdWVek1lSrrXopB6peVzutYnatPhboJpG/v
/OOeRvNUHXmYoQIPCumWfc3dZr0A6rzAKfPCXRcyb3wA4aesv/lAHd1rr49aUIcV
xslp2El/S8SoSBJoN4zQJWY+OZB+QMY3cXjGh8lOMUIQBIDPtqpz9fHTxZh1GzBp
2qUSTgG8cAz8HwJ5uCkBf1WxyHXF8oAGPLcAmFp9dy8=
`protect END_PROTECTED
