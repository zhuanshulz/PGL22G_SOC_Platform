`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJEOLjbgNNf5YiGmJwrR0B4tYSkXTNp4OHmRHK3Tr0wR86kk9dnB5p+AEaIv+YIV
MD+dykjI4WvialiKq/DQM4Meb8SNhaUYz8x2IY8uO/IzLyfx438g5o78yPeDN0/I
+vWzOeqP+2Ls8ZK3EVQ0VXZp8ekTTOOQ16hDV7Gg/iUw6kGz3EpsmvOlnB73g58P
8kC8ud5kEh7s/PZiIKwkVF8ZlpqkMM8n6kkrbHjjs8BTQkMp8FuDmUz6zi8OoMbf
Bqha9nnQrevI1UgMncTkuTB3OR6BYIi9k7vIsfaWkDtUl611fGOe7xAhBy7GoSAd
42nttrLccCqM67GSw3xD+jWTeUmqBg2bfEwD24DF9JSxMzEmh9GXmXsP1FnByNfZ
yHitqyzwCNenKXLqf47SR1+NijwjMFjH5LkqkYiReuWY3EWQMbrj8uPW5AJQc8+w
hh8kqKKVG0LJILdm2EBeBus9GQiI1MGVXq7VhO+s8AHZIIdYVnUs16ta7lEWq/KO
dYlpctXRLTsNm9O13hKq3NGR5W7pYkxoLfHd3ju5XqpjBKxS//ZBIAzP7MxdFI80
GiPa4M6tkt1vSxSBQDG/cmHNSNJBe9eNp8vCWTyuegaeZ8YDpjOoHRnURjjrw1zv
OBpvRW+G9c4bLlAYZ8wgsU5w+7Ne1DvYq6QN/ji/LNBEezigUAvabu9ahb9ZNRfB
wamPlw7V/Ow/274tKkyFZ4qd9UGVNOjuMLdK+wd6PNL9AGHn99nDKZ1SYM0nmFem
LMsS9fXvguKYROAEngWgyqMrSJW0WLm0OtAsxjMeMpbLqSHgcWb18dvOiEtmk/4f
bUfyktuQ8DKXjKIAwzw4nSZkbO0ES9+0WojjM0iieSEoUeBV26a7Hb6Zy4EdTsXx
+M5U5huwydRa79y1mk6psTpwZti9VQce57NAQnkzV3v9PHhczai0YujZkDK+ItEo
l5qdzTHY1y2IjdTlC3kR03Hqzn9t1dP1Lop/uKarNoAu+C4OyYTvsgQElPHIc4PO
jiKS2VFI6M/yDfVDxiSHVKyOaBny3kpnoUNqoM96iB33J/7/zJ9M2Mlc5lsgL9Xv
pdY9Fe6f1JsaNtVhc9zzqechFu+EjVyREKq/tr61vakJZVhXz4EbR0ENpyfFyA1z
DaZIP2wqFUM2xeZAkB0OEOnvyDfkgFqwgw2uvaaWVMQSfsnyzNd2LYWIXQPnt13d
pndfdsA5WP493j5RrxE7x72LXKJPX0AvRYmalyPco/vrEyfzcZy/NwHQvOZTUBmA
K4yJNHDjcdZD4fn4RnA5SdAJU8mUS/d5qGeZ3TnjMEh0G7CFVqG42Ig1e8RTvLOm
/Xw9SZheR0rSoN+l/4cX8DVX2GX/LPXvAimvbskNbEstxfLic2TZ+aURVnvau677
CvdFTYK1xTBRUlO7iyQq+6p8zr1FbZowA0Mz9XAYPbY34A/HATMHFZAH19RHZdKu
S+J4PF5aeMOwi20xRtfDttCpIY1/drA16jqotAQAdDWSXah9/JIEES15AYo5NRMD
s+BkCifYrojlQTeUP40SuvH3kE6oT9RdEw2uOcI7YgdszXWmW3QHo8xt3zAvE/ey
DBn3H5zkL3fgyZHhYl2/jzj4jQb1PCU9FcpcpmRBicjVY4XwsFUg84IejNt3l4Zq
Bz7lO9fWx1XHxCZOK+y8+5PvzYy4AhYa8kd71vRILZEWjJ5z5Y45KENjrpHDKwzJ
smt3dNyhMZiYeF/A78KkP/B3pgJU1ATMx6FYz+N1rI+FGFa6UUqln23BhAUxe2EX
RZXA8AMVSlmbwNy7zY5opypZdyaP7NH5kVmcqfir1fUKn31+012bRFqPPr2bgts4
8+BH9m44O3UsfObUzFK6urWbKgWB+BkwOVPY4FlK0Qd4AmUjgUBEFBNwhVt3i0W9
9yga7dt4MexxH8uRVoBSigwQDL6i0nz9pRiZeI7l2Zh3HeWr4AWkFcSYVGdsxXky
2w1zBHsMqB0AGvcWm+bF3U4+gpIZ3MyqXD7606K5pJmvqLjl4RLIbZ1fFrgbgOxA
AHe8HLhXUkFSAcvKRckCVD7tAX6oKLQVQGdBcCbz4lP2rPe162T0BIHVzLowRdhx
5bCkpccyj4pyx9zIByKhG+c8ZqyjFmEiHD+Pbq9hqDNQvESy6vAKGLFDd2RGYjQI
rPqZBOnmD1VAbQuL87WR8UjEPWR3eSR/XKUoa6KEOxf3BGPgXGXPJWakrO/E6olg
73JGFkg73y5N90+hh+lJ5WAf+XiN49dUULWjQuk1F+4AWtL9s760AHkE7oQ834Ol
xyttXkkjxEhyPutOr7BO+I3nMroz+5oKCh+LVA3ARmEqR4osymX2pmPiktbayBrL
FofbyApcEtZqmPBr29t9+MaMSFv7p5Uze4z32G9vjqcCJS1oDZMakaT3ujndwZK+
6aDstCNv9TuNJJ1Vr/oEaT+tF9f/2hBjpzv0ZZETSLT5+XoJK59mrVURCFWWptxB
a+MUJ0iQ/QM3ERv/FcwBIS0p/fvsvZ5yZxx0ZYpG8vnX0ZZ4AfBMQbkm4gxVPdDp
nyup8CrCqUfhU01h6sFqa5IUMI5K97cK+W3ar5A4q1PjQ0oF6hOH4OLNmlWdlHvb
gAKyzTvtd/RDo8BEvOpl7POS18h54/8BWXtC890k7OUb1j3a6UgCeUS931p0m/nF
jSV3jPhAAE2I15AskTqqiaQGJV4OhXAgZyNthrRgbPBIeqR3biK6l8K+1LQ7c8BW
RdxTn1kX1hD0ztXRapBlQEUAVguH0gHotl+53Yx3OzruMwiWCLTlWNvPOdwuGtQC
ajI8CUgfu78P2kxP5REY1zW3Gy8gOq/yjb076A+MwM3XjW4WMtGFzx14cZDWDyBv
6TcpOfMO1Sg+V43kW9ig5g==
`protect END_PROTECTED
