`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4G3hztTWKJZU8HhQ5roFJsgqgjwjIudd2zzO8flnvVaOUIKgNPRJW8FxCwJGDjkh
crMFRiVeMfYN9kk8NZgSD0Z7rbT7BAcyzQqtGoAe86dfs6XlybmvlZG76SfKeNhK
VGGREQULXyYGFJOB54pHoBX0faPS0dNyE0MrsRMCjPGIZYbMCpoBsXCodSNminGg
IX44RfTJtu2zi7/TZdaX82hKs7tSpR4b0Ol8ob05Z1exmTnp/d6C2UNJOjxFFI0/
B3XSHsvicdsJzoiAzqqyd+GiQBPh/hUopBpg8oyM49VX2bN2EUwBUjWZYXnFyIXt
7P2pwt9bYY2m8lqHH8l9hArabTGMxLjeJps+55kRkTd9PU8nKtFqkBNcU8QqTvdl
ZInyIC4FjhoZS1CiBsdi6LOOH+/lYXKS9czUqEjnXAUS5bli7Zr4qCg+QrLDTMB7
86b4X6Pa7kqRgVoMA122736JWUM32P3n/SIj78EK5jka0VpR0xCGVBIPINIS5QHr
dZZqJ6Yz0eTpapHFozfsYuyIfsIY9DK2m7kGi5wNsL1Y8wVXRTF+swyJTN4dlR+y
1lnQM5Zy4stBd+8fO82n1YD4gCk/XDqHY+sc+r6g0oQPyc75wLuBSCpQcPrvosUy
Xb1eClUbunsdIwWufvxwqPOw2S4CXdAhix2itslo5H1P/8ZILJZRqIG1YgSzH849
8F6W72OuZEw2ty26Ds8TNUnrrhNagK9cymHFHRoPUBDhdCw4eOjO4TNcn25DvVaE
WMFr/4KgXqmoWaCHIgjy+blXt7PK10Fy73QMMCw2SXTRJ7k/0WqQ8owhkgvnlsaK
0I7thySWXuskysOBVerH/O8JAF0iP4rXzA74Sm298mufNC9ySOWNWYmKujG6de6s
S/4yJiN4rNUWsu9J9kQVhanAt2OxyEW8+In+VezE1Ng2JVzHSgkfS37raXI3eKOQ
beVm2+DLWcYB0SqyUaYXWymocrg4WmhjSBmqVVrZbdphQKedCMaj53Rg9nkK/lad
Njth6T5+CjHubPJsAI20md/fY5C+qh3r28I4y3BHejeKZu929SaczD0TGxZcbvji
BuhR3di7RMO6/QpBFXXThEHO9RCOFqUVSBc8aCnxwAyzhtmkHuibNyHttT9y9gAD
6h+Vpp2/K7g7TQWW+qHoXQyRsaO0n/8JerWK4VKkNmf/anHovMg7ZaanQBcABUoI
UI1Mlu8ySWkNvhBTC0FFL8+GeU0UVibYqXuElT3izckTZc092mNSos7tQ6JCmNwp
FKNSvk+5bs5WpVbT43edNwTWNRIKU27r37AAKplzO1ToI52+Y0C5DjztHDpx4KmS
Dgfp5ZLcxbFJOePQbmvAw5JNqrhEvuRdCOjtdAkRCiOB/+GkjC85Yfasor7nWGkb
KP4A51Nudf5CDE2onrjxKsGK+ILipoV0LoMyuTgu0cxd35QbGiPvdym28o9dshSl
0Ujtkp7r5LgF895n4OaD+xkEakI2q0ZAQ5K0JIecCf7idbZ1uNtHakoSEvSULxaX
tHO90nPmjQfhfuh8s8xXjgGkOk2PYpyjnGvSzbyLmyCMEPJfX1rxvmI3rrr5ybxV
OyMksrjDyLqicDjGOt34PVc9s9KnXdfLDNbkoFS0jcMmPPFQLT+dXNiYVio1nV64
plc3urB1wFqz/nmFpRALOsVEJsskdPR1RGw8aHH0tneMLTDhmucDZkQwtoBbqeA+
mApwpLKcoVtaOgYwPPfaK3GdZQZeQTsKbKNXXlmrBPvqk2wwZwrzhmFtYzhmveLq
xJ9S9sa0dqB5xlCAYu8aatmT0Lmr+dySe9aFCMPRLyA81CuTs2BjKSzboI2aaqSh
CLjhebnEwkDKQvc19UeOdmWpzYuh92nDloxlheow8KGTDNvO49gDk5zjbdKw0GoT
pdXGS66HaF2kACweZUJdAZZ8m7t59VCiaRbFZg+8Fp5tjew7vxtpbmCA8JD2/59D
aO0NpSkCFex3WsHqEk8JNCL9SxHrpPyY0ZHx04WVPyoUrQbpfYzDa8uBWSjTDAKD
r14B2LURLk6VEPYbMapVUZQi80Q4TaWFNMoFYLRZzm1/QyRcuIwYfS+WbEy3cQTr
wFw45+fMMk6FnikjMLosW+C+cgOMHk9NTAEdS68pLZ5evRu6GRYCRrXEzrAGbRgr
RYtZR4l1MVDsKnbvKkpZHO5v7aKSge2yz/YLnoYrc6+h4AHgaZwg+P5Y+MQAtiZS
cS/XidugePkEhXa3lNwgdKI0hEF0cbl19udi7YzQiML8rteckF7otOI/SPqK0G1C
taH7fK2MNJ7adRRMYgrGiVO61djZSbXL6Ww97+AcFPpz8RVbzlKRwxjMQCQQGy5N
Dbk9xjJqzldBUtYbKJy1qqUNNjUQXu3kvQE9DYGto8NTDfSjZZWa00AlW1lM4nmR
BAHuYYBxzLCycrXSSij53YlMsSM4D7F2/il4fovzYYa/I1CDSPr14VPssZe4P86g
fir7PPOWKDTUdqe3+qYyO5Ifg/W6ciiQ549eohZF8xR8HJYLOJ8NXdny3dAPRsDH
QmuV/qzY/9IioaUz+OFO8HeNUKWAhUP5HqzhWJK2G0ZDuRxjlx8/7YLOQbx/y7Rg
y0ZWSaH2hzolAPs7FlK4GyxuMH6Fyr3XygTrGWjjlEO7V3ka2V4bC9io9JTQRAJ4
LYIgUQlpipnt9QSJSak9x/jCEpq94SZ/VVAJw5vYju7YCa9dy7SL3bJs0iiorvmj
p00CJ2Aeu8HEAUWA5lyCmhSk31q0z8Ow8YjaRo7Nsqb4xJD5klc2doSvTYOGpqqm
AVGScTsidH0M/uedM98WJqn/eKE2IkEfSC5ACEYrFeUKoC3Vlk4KFnoQ4Mcihs8k
mflngkivynCgZf1CXWlhZWXN6mIloqK5/exUJfB11PwDEQmCnFH01M50xQhYex2q
IfDwhbjWzSXmemIdiBidXV7ijL0v1oxSABB0eGaWGHtoBDBinuTtZ94yewdjyRN5
C1p7r2exoy+aFCC0aUqOZUDrPUNHjQx1qNS9fl94C5OpPfseOjxoHT235/Y5k1k+
utQIc4IWfIOoWMHZn55aS1Dj3a9l/C1l0AEFceIzQxW6/BcWApdx5tQbeZ8L0tAB
EzL3C6zfQZMwfoS6eYR/CzsNgQMuMpiLgXwQ0tOrMvaaLuOuaMMS7AkN7eaSNd5O
R5kxWmFJPU83SWOKk8Z6SNZe0uwKO1dWNBa/BzxuYN3N8SlXJr2e0DhRSFVfBT1E
fVRUwDkf8TjltW5QaHAereNoib4TrVdt5D2QC5IqOxvAnK5mOhHcqMveAzZzbmb8
PvE9oNpehXvLqhlqshp/O56+lUQN+diYOwNWnW+/XZiW0JZPkqKvqW81MbAbWJQs
/X36Nf1KToxwxJ+miQmzZBOxoCteTMaKmrP8OdGwLBTevPyEBFuMil05Cr8JZNLs
9g/4hkaRIuxCmv0D42rrZX7N05gcmM4WgAsD3DXmFFwCFu+mC3jHe9YiUdjLZzy1
298rF2bb8nrajG22NGKrjMBNinQVV+V2naMXGzY+ldVpUv5SVFcfvBJ/+XjNLuZ5
`protect END_PROTECTED
