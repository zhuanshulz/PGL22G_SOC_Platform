`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ms+2Y/C1y/9b73Kvn1Adx4UbsWBHCV1cpBq3bJ+0k4YJDIUZ7PLA4xCHBe0KEjl2
88AFaWGO+y1QgbZu2KYN1lvn/o6PByWsXL7JAPvQrrAuk9TJm5LGIoSCZ5P3n9sY
pnfabZyfKb5dARzbuMY5gTdMZaVoWjby0Ts8mtOdM31CSkE4THJuwr2IvsLNUBqj
VMBWtJp0pg4JcXebgaITXGx8DxRf6/uRHf/W5nxjF+HaJakR8/Ia5jRAw/gOOnJD
I97UYoJ37cymWMNnJ5OX6XTYGWpCaC5VvknTd1YiVHpEYNL8JZUmTGmdUELyXdiQ
0SWrtHFsbQPDIgDOSCwJ/XckJ/TShMl7C+ttunOxV9LvIKJrKuPa/Bxg0g0fyPXO
lXlfRD3AcSrQ8wZPsH7WkgbHsB6XtMmHuEZYl37EWyCV5fq1/CHYch8VhlinGzuD
lqfuAM0SPlZJeDm7JsGvsrgE5/2NHIvt/l5UwVOyjykdXCktGdSo6GMLCWh32vye
wH6eez1GIwSnXIT93GNRH3NHZe0HRQsL/FzZAfNqAeY0qvJDRpgtlMMjgZYxeKan
/l6jnWcmGYOTyWmtGcFyUjbPsDlJc7eal5/F/q7EqSVAWbo3Mp7kcqIi5ZdXgrsw
0e63RR0tOnaEUVYOL8Wteqw9kjbZL+cjncXkSNw0yYR9pwJK7rIXMxmPJoj0Se8J
`protect END_PROTECTED
