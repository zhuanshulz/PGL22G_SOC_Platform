`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pz1SAMfdX2BocPPXdKh1Ju7a8L/IC6QgFOzskieFhZbVLKEh9KCtlZBe4Exy7D6y
6+U6ocVVj1NJdaA1nH5s8Z5Z58+iZPCtrxlu41T8XwrVpL1T5LB1E8jgO43Kj9vX
70y+Fa4AH4QmE5i6GJu5UdWZDcIG/JtCNNlvswyC2Q3vmrVzB+ZiNaS+MPufiBCN
z83m2npL/Ij4721VrfCinRSiJcjyn+jr1sarf+QLnsK+P7g3RBXCENWL7FaNPqE2
wnooEubTMJ4tmhROh3qLH1xAh5tNdN+s8aZgZEvDWT+DbupHRuKwzlhPvvx1gY83
vJoIrvanh0+fSA3tMcidBWkdCDbLV1mAXofxG9u7s+1AJlR+5z7wnXCq+7QF/C1m
7pt7OlpFrzUsfcBJeMSE9j82GZkZvffh/0Kf6c0nNtNqaSOH3KyYzeV9tC1oXQ8f
sCSv/wKlTwy245mAeiEBK2Kp2Z3dSstiWI6brVsUrMObxrRiNMVA9f8MfzO9GIUG
+2fWDUkXoV9ZKasbsYslQHofTFBzuTRLqPf0ah5L2z8ZWC3kE+qfbnTjhiktDar7
jqQUonVjPDxB7ju77fXnFUXY4rrcN8iHmyiCBzVXJyH/PdVdgWzcSLfJHZ3mDk+/
8nUnDRU5Sl6YWmB2pkH/msfZ08N7hb/v+tFkXGCxy0leBGz4/RGfmZlTKeKuhPQQ
S4jrh8nFTup6s+ekMok0SN+9A5RjPuG3psVmxxIfsbQdGSvyGoGGzN2+d0JE/2kK
fvhZ3yM+rKe0XL9X7c04xvImTHxJdKhikRjptJGG6HPLfL7pIALTAZIMYeuLO+oy
NliR7V3KwgD0+l6myEkATvichBt8vpRxiLX6iZe1S0agEpaUM2uU4BzRqo2yv/8D
b8UKDuVyPCr8T9rI8nGYTB4u6K6oQ4y8oAOb+6YzHNZy+HhWgVjjpGxVLMvjkA9z
zU2a3sgqoXkexz325Zz3aELCtuejPtXiz1Vo+eCwi66HRbwEnE0WaRBXhZtjLGt4
pp/VLtDO+kipuDmyfzv+ZS+4DlMeW76905JxTgLTgG/l+APt25Tp5m7nPpsAR4JS
bkPDMAlutM9z15o4tgFPKhrx50k9bzPt5WpXPfiVuqYn0ulF+bULgj8sOeRcbPqo
7wmXs5Y7OFP0IxERvtggFwOAqC76b2Dix9k5ZvM78FIbgJ88HXSfu1Eea/xx5PJD
eZ70Wuy/k0ZoePO6brKpmN904b5bIddtAu69gJQirhoinQ9npfpDHXNmwUfBL1Ew
Zv/laOThK0faGS8CAFLGAEU+PS3m8Ry6RVb1Plp7bOqthINV0rCAeHhGMQv8z+S1
HKotrylacBJedF2DmAQWSkDdHXM73nXBI6B1urA0MULUW+Ed9b1GgM0mObXjSs8a
6j3dKDezpEMX6XAkGhOhUrR2Tnk3MMvUY65sDL0LU3YsvQOIbweVd1tw8bkJNsDY
fRtso0EzxLNNwFZ6T+FvbzjAJbhMCalibWLiJRfvfhzZSOiotqEN+qTr+WYQvDIA
pZOd/EtfC5jlo7VMGSNiw2bSszB4OCaRvBiMmmbHqRWt2vhMT4bxZinpS+YOkeVg
CbIi+gN5dCmrAz0SEr9tvbYebF6YZthyFZT524QexVwpba8i+93C1NC5yUPVb/IP
gRavts/EbAC4RuriZXPtInetr63jvUNsZ8a7dR3C04MYiDk6MQZ8+8NWNDPpO6hj
XADzHKRxGhMZ48f6nWv7g6Ypky3DoJy4PKaELmJdDvMpyuIvhmpy1qVfoGTFhenR
SxRR7P5D73UqpZNGsVmkvdWLxcf7V6KanUnF+NGRF94G6aPO0RafkSEuSwp7yfuH
8LKjzptCLJ+uJvfqXezSVXX5dIUx6caabF9Qr/iy5Cc80zivorw1yZL+iIBYUBIZ
28APF8rrMC6lqEnUFi+ygJ4haZIL49gPHJxQtNESLJ00SlPZS1m904WTFl5UDJ7w
zLl6qaFsHvWlLWAyn7HYuxh6vCN7lkFh6jjkDs3xvTYDVjAGlCzopwAhnSCYnaEc
vZAXz1Hyt+xZUwLYHbGeZqGZ5FihdGOSvn6s/WhQ//UL0BXLbwXkV6VSJ6vdGy+b
W9jDatgzhBf+xgCPJh09NJi1gLBSO6+QVQOV7LVCB9L/Jp94rdTPz+O7VX8VW+6S
z+TiSSP8Rmhnw8TAZUQ4mzAlC3mWzm7C8EqbvtLoKv+1XPUpuqH4f8Mw+xLnt2t5
BQTXDRF5LdK041HwcJhNKg5oV/fpbLvczTzl2lK3p6elu/gFhSKgkNaZ4vGLebvN
WLj2sW2n1IIu4jbUEnOFQP4I2ggm1EsT7SUgiSXQ3MZ7cqHmOHEJF+8xp1ELdc1t
NlrWWo85/ealAvOCzF872hXIU8YRFxrrRFciAHamyhz+OZf1I2U1wcs5oXvEivWH
5ir9MXtd7KFKzVVtEFVv3WUYCkXa8iKn/3U2eaL5CE+mxp5vKETGDMNh9iaZ69qu
Em0FDpnTR3DvHfEfJrPD+9GntObS3sG9T6DmAf6rY67GXUCszHHMPOLm/hMq3qhD
`protect END_PROTECTED
