`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vxCwXYZSdMkNCFPjI/iMEUTojZETr2KvrDnqS11afDwnWbBD92Zdl8TIY2naDqh
b3YHvbDstcvKQyP0CvPNQNrmis+qoxdKMXi4p9hO2CLxCvCim3az7HP1ktot7iKb
DJj1PvCR7lK96CUAb6sQO5epdPEoWsss1Pg06bNjY2kSLanMD/N8byhlZ5XgAaSu
4wtVTXgZxMl3u2WAWjjWodU7MgTMxvAmblU1NVB2OFL9gJ8kyiDq0dVaysff0Fkq
Av0ODTZoxEeVl7V7B3NBRHFPbw3BPCEz3fy4JqQ0JxMCjt4ZzUPcFVvH99Awr6/N
UsO107G0r5NaiWaKO7/koLqp0ySXTHRWZpzZUJ3U0BZJchwEnhTHf1fuwMDmswND
OSWFD1f/QK+/b8rl7MoPFy6G0iU4C2SGJghnir+26BCeuIF6euQif3onebh6Xicy
4gC41Ff/deX0OocuWomGKCrpSHzyoKFeUrD1mQR/7TKOSjXPiYmbLZVSRZdL43+a
JBR5JKeNLUo/sMF06M0GwmxZtgY71yuSVpzTJWN1ez2u53TLxdS77kOVoFUQX/UD
aLjaTvjKrW/x4PWjVgdv+TtmPT5UsrjN7iZS6C+06whNw1RZC6PG5CTp7oXp5bVI
3kzM9dOJ6gL5ThQfNUggr/YN3Ay0cQ9SEtVbGcRlmD57Bort6/Qw4OeK6TdjBQa8
bDnxYQPYCeURWHDfMdS2MblCUaEUsjDN1r1cvJvvjHZta6QsiXUyOMp1IZMMpxB9
kyiLArALIu8wuHjg7IBaSVbESlbja9Y5dPfZ+NtGcNVd4UPv4a1DoKAFogxBawT2
wRLksmc41e0xjQQgNL15SDVazcMEVlw0wVgR9yUBqyMbW2X7Q5ggVRfqCDJCd0xQ
8I2hw5oDSdPQv4iIBB7IO7itHVtFoTBKRXXahGdwJisYOcNUJqrj8u/PA4WMl7Ht
1SIdYlEJjpDoFvL2NZ216in8bn7v5TL4/xW5Sgf4kuhfojDEa+U40BQhpmY+V5nB
QkuoFvHpZrF2+bnA0lu9SUXXH5MyAybyRBTFyLzFlS0ReovJK37bDisjHs+dp+wA
J495HocII5rWZZnvF5MhszhpCXK+FvZ8HrH38Fzxk4VEqLBdSgZpf5GWIFqbO7Wl
RNTWtHlA9bU/mqQ31eTApOlQaemPja7bZxRhz7pCatuqc42QGfrar4cln6s1aQD0
RmabjLkhX0iav80+oamngbJOyeEWKBelJcs7Ihj8gJjVtCiGodifdZoPgf5WyQAy
dW31bsT6YbO6pB44nOBGfKnVmTLswQlyFslocX4DJF5pnoYkpsifjXzQoEduQzIU
TscLXbGvCskgzyMFEipfhz2d/j6Fz3pgW/TIDhbSr9m4/WbaU/FgKD8b1ANLh3Fn
Fe6Nq0xt82MPdPD99NexGbc1lteEl6AQdvQqCeGAChW6ljyy6L9iuWgUZ+1gp06P
pSW2h/Q8d0rvk7lA+vaREnrRanewUXmYgX+2oqKGlOQN9VX/sR276dkCFIvrp9ZD
f+NdXMY1WTrLx8U7thJYByGE452HLLckmhL0y5o8WhCgcoDYG+FlSy5jMMfSqgdS
xnHlsBZ4nWAgTM3Z5BYp+/cdzsPayJe2E54AQjYPpfIdq3u86Is+TqyjB8WUSdH+
LYICJvVeU8g6OqodM4qiNaoP60hdOOuLkt7fnukHanfND4/6jpYxigY7FRg9EAzz
YsEKAvL/MQ1Ji3S4oJNxUo8T0hXDw+rlJryXYax7KpwMGGKXyfT397knhrPv0PX1
Ccazyn/0gRUgZmvJlucGUlBzeJcSTqmPsx7SJNVY+fjp3UkDPl2msal0Yvf1qF8v
Q9v185ETbNNq5RBX4vUsH1DuuQFSQVCNFadK9BIjtdply0Uh740npCvafvxyCmZJ
uTdiBxtYX0APERCSmarAxQa9Fz8J1ItibJlxposrNtAIU7l1oTuamQ4d5ij+u7mT
58RMwFJlylNOdUUWC4v8hQwY4de7oyF+K7/MUzdCmPtpIP8gfyM0wk8+ZRYfo9Fv
3VmrbZpC/Z9OgXvr+WPH6JDjPy1TSUzXWDluZ+DRvYKwez5umAN+opudf++HA5CC
S1Um6i/mmkH/1Ts1qe/4osya2nADxbojPwgElQDA8j0wP+o2ebAuWlFtCTLSa1w7
mTIviE92Mabc5zrPpt/tNaajtXQCd8I5dV8iNpEw+wIyzzOkiAlf8YEyWvH4X9Y4
/9guPzLd02KUmeZ/uQ/ZnVMfSAb+GIqAYjT4V1UrxF8eqjf4S6todZzWdZUQFhC6
QwAs4HHVG4xDuCJMpVIEtqVYTLPMaI52cTznuMYwAdxUyGV5d/kGf7eRH5+KzSeh
j/HQJhkSlls/ZOeFq4n/ZL32y57adDq4dVY/4kjgBOE0ZT0NOJzZ3Yuw9d2gBhR7
7ur/YSgx5aAT/2IqaiEU1JcyCsx0N4pwJruAkYNPHhMR9jabwEIHEqAdh5fos3es
ci8G6wQDGfNEeBzJJ0F/mSW+wn9Xnn55AC2C0XoxQkNKO7rppBixisW8Pmqz5bQI
Felh3mcYKjRXUIBbPgFekRVda0+vjWvISl6jxTr3JjuCaB7V6coGan8hoJDsnfHK
clROllUgwubNnK4JSDKu7FmnP8SjIAvT1YYqdnHuhkee5dhHk3oS3DA/v81nV4/r
t83MrXKXXXUEbGnX8cJJLnkPY9tqEu79sF47vGCDiXs3+Jpe+YOYglBibFFuKX8j
eZrxnW6yQj8VmUYChHDl7XdA269lFdXWSCLgA6pJcvdIlIE77cqC5Cnk4Zt2dGb4
iFkgcqAiF+rG+MCNy6bdtaFL1+rkpW6Ex0YTX2X8UiET0pq8AWMJSa3W0CDVMr7N
mcwkp1ZAsTA0kvJgvyONgzZpIaeVyUvqgCdXM/wmALa6tGLxnrGV2AtI33BvhccH
woCJ1PjubuTiotBYsNnFGYSrvRwy0DKaQLFCTrwEpExr63JyJF7qp/VmNaRZ8rYh
LUVuZKNRr2t/jsdjsyQ8r8rYFcDlWCKK5+i0TrpkCAWmHHv15XxW2xORv5dE79Iv
uCxJjmxppVbeuc1bpp7Tj+GSZid1lqC2FlDXGPHZjbD5VLxqgmE/rCRSwJlbfbZt
PjjhIxt6ElS3YJZ/ggzBXhWuhDHeGmG2rmUYXxa2QnCPPX3OY0g1XKAb646+H8Kk
GyY8qCpIwPxlJzIx9TAF2xkNZbiBXG+hM7mfO5unr8hWsprCXOpuzU2herVl2ni2
FXHUaSYLzBvAjNjxCRDSCbGBKo7Np8CMn5B1QHz2C1J1+oQVAai1I43PE/mERKKx
MM5HArNsR+jtifmQcIIxMHR7Txw638inYZVvqicjRCxNaiXg8NiOGzA1vpvOI2oj
pXi5r40pgBuBFJLoFsb/wyp2iOiLdYU4bof3RwQE/owkYyKW/LlvA+NJsa5tIXLR
iaCTDJkX5AE2RWnbQeoCxwEqMokeqjapw/IcFcfN9Lo8/JpTPiAJ+t/EsU5bxMaq
/05ykA62k7CpClIRDSnJnsRa+P1EQKMXnpm4hrStOp/cn1Bn+FCSLGWQ1GpG36Pq
Z/mi+HLEoEGOGs9BGz9ad72oqzo0X6LJ0oHFfSqyBU/6PDrfvS8Kl6NykMs/A/rK
XvRL0kf6RzFmVbD1wjdN8zYpQH7JC0KXmzduwh7H8mqwnHVqt6FtLZJBs4AmBqLH
EKOTElZPJb6z8TZzn98hVJvREXgex6gW5b9I/EZRN6cP+ezgfMA/lbQNd5k4fA8Y
jaeh6QysOb++jkUYSHGlAv9MPkg4JFNMSjY6au7wE0jZmz0AMsvNV8VUcfouas41
2jA5OH2V1Chd04ebc8t0G6fFI2KdIzVwwD6Yqsa/nrwv8N7JhNcjuESuhzWqnCsP
g+ymrmHWyDTrXSzUIrl3dWG8rditv32AbjJy3qRh+GiHLls1kY1hKsjCDRUGZy1D
/IeojtiruJ23Mq5Sl/1J3IruOgoo0yjGSGYHqou3hSN3un5e0sH6jKlFlmLq2E+E
sAynfX2FoCizvHLKk9zY4XIVR9pv2KuvN0rG9nWGBGTn3SmFYKbxO1/sCybwf6eq
y2a+v1UMQa54DU7bnixxaGeOUpbmA+Kpo3AdSZFUNqEmqG9ykFjMCNqfI4K7ClOx
Q5J+6srdF0oDIt/RFLq08Sn8J6eA7iQ647EnyJ96ClQKmoegiyWshnVHoQDumNAn
4BG9kLuELexNX2E4jS5836kT4BXcgYnijeAdt7YtfOgYXWPaPa6D4YTR0C6kIJGN
YSRAxOW//kdhtBRF12mm+Mo0NTmn81cUvcxJ47/OPtQmqpusVxb6tIOjhVnLUVJu
1+Fo3jdH9Pfud3JmGmFmgit4XEVXB8CSo2AJHwZeiYTa9Q0Uu3vaN0blH+PmLsAz
PXMvdkrEYNwLXyx2Tz0e6++0xHzuDdJxrjLIn23pArCAuRGA5t1e4QwGPp22VaD7
OE+RTpyMIXWgCpoiIwF/xDUfI6m1RhzwEMIezCFoDun/l6Nc0pB054yL9LOJrjAw
yxQfba0u/1CsEj6v2b9LyQMf0STFNaKaQF6tLlxbFvlXheRvGH7RarXzuqfyJ9CA
fLBPqFD0gLOzSMnbkimFx/pkzUYT8mR0K/VY68hjvSHyv56EYuEl2ohUokJMznMV
o7juUgT/auLqWSoLPMdzKO3ZZIW0yzAP2YOGqkoWF9FN9DDIdk0xW2hKg6N4wgBn
YXMBY+TaOxnCjdcOBN9VxBzPE1N0mYWnTnRm8siSSJHz4mGd3QgHB+2L4jrE7PxX
WkOLlBpS/aXsjDAgRaDS1tMf/K+pXi9XGebwVmvZNmQvemaMkb2hYQU+126hqwHU
Q5EZnVkojBrcndyGsqlmWMxY2T1NZeiMKUq5dS1QNwtTrSfvLdaK4GfCgxWdoHC1
1vgrAJQpXasKHzgxN97IZHBgvWD94mbPaMJ0RSQoub8092yMUK0DyqXK+5L+Rtsp
6yqZhFvLXm147WfCw+E9I5qkjK+H7AEx6ldr8I4rc6Y1e+9WTnbN6BM/r6G3LdTo
xoahUq3M4CqnchTadW7OjgD7zx6eeop7RKr6Mw9VZ3ZVHK3JmSOOKcCavpyAjhQ3
9n8fOzsCgqMlPZyyswItQ9OwVTdYF99hPtrcm4ZLyolRDU3GGvjqoDvrNMSTTYtt
UnGayPbVt4wm3EoSLXM46Y7P8OXOSVPjo/f+G2DDaAT0+/upCjl0+HOK1oRPMifi
IYkH9fLOZTPTNmzVtzCzcoqOZxEpbzoFFmOq2rxTEPMMGA6HyOH4RoFfG7uHt7Rm
9p46/dxDUI2B3TR5vgFSfNRtMV75jNPzfw8gFmHT9/8uoMyOvBfXn9aWZO8Rws+Q
Xv9yKPzrA+cFSQuGDBuhQQqk4u+/GbzANAfPy7qXemT0oqk9VnY7yIgdnkREkW5h
g8XXHcT/nrDzG5a0oC0lewb+OZcXpPjpDyJJ8IlfXffpp1DaZa0MSPfbbU9MuDmT
RCMjKicvwqW0BB2pHgXkhjucs9HdoA9Dlgw9om43qBNvk9OFOSdazFVIBt191kwO
b3TZ0kTvk1ukpz7gCLZ2Gvhp34y+2IGCSGbFS+B82fnUd4ykH3WjsKc3riQt2Ao2
ej8hf8POSP1Mc11NkyZE6BjiGc7wZLh9jTx/0xhamrgg83qj959hirXz3ldrD+Z+
c/oNvFX3wOa1nmh61AQ0GcG7SbYv86LVP22RRdh/N9RF7Hhsnu63JEoWD0AqccU+
KeFAqpfvhpmqsPYMieXNUIT05eUcFGPMYwKnfmxSzihFnf3CTHhOO/1G0NDJmj4T
gd0l9hg52jFynh9sFf4TbzdUXSDgfZUCHxumMVz8N6xR085sigBTa4DoDHSlt/T8
C5nKNVuAKABq9CMS9tutzlX2mdr0RxNZrBq8fisC7bsjmDZgtOSbevR/7adjywgR
rB2gWXdeYsLttmVV7q9Tv9wdUPwtsfftl8C4qbNYZlE454pZJKouxA+eCnrTiEZF
f/bjNYD6m7Iuyz24soH+DzKEPE7WaPh/X7ckSq2TqMswRP5iP43uG9xA2qGrlV3n
9a/EBfze6CWfquNQS3sp99gmUJQ5icDbH76RKPYcnkplw9T8YEpfRw9CAu5hB/8D
F3QYGU8K2cyEFdcsi3JlmZZ2210Hv0UEWC06/VaYfFRYMIeOKEsXtRW1BQdoEq78
lgVcSed5+wLP+08PWrWjJXMb/6c9eFfPxqhcdzusqGZ7wr55nGA8uIe92PQgJKgx
o6z5Fpy4YbrT7fCTJCIrlIZR6a5g8GV34atZNH4p9vL8Zw+PEWElGulFikhOoQRz
oVm8x3RnPusvzkPYIF5nvgKNZDUkMFLhREJzGPDZU2uR3a9PneA3pAsMDywVXcHY
339TMotQHV5sC0c5UlpTwNmIawLde0E8DPJqh7OV1qCMB5xt2xWHeAhplXjURLfI
jt2l3mLnvPHk3+/7ublrzoJ2Nc3FW75a+C6oZS+n42TtVAQczHcuk0IJ59xgHmaM
qHBd2Xf+y99ankNSBo/79kpcJU9ybEn08v2fs4C8CMMGX28C/u0VCzMrYYYrJGSM
YZVxaQ18rzvis3/R4q95+4ulH0c3QpP3WhhiKoC1BTCw2I2glQQW45vPYXR277cG
8fc1bzcQnd7RujWxKn4Gz8TJe5gRCo0af6cvLQuT9SbrxYUgmli4ugaA3LbqHmZG
noirDAemT23lMQDhDd3yTDbDHuHXdsX2SkhiEElT3QmF9tVIQrejIe8volFqfK6v
F00ahG8eSxEOzsbneILwJ6Bsu4qanTAzTff0cDJ/G9b2dL/4kMGoKyu2UqtYdo2H
0Su5DELMoT7oGBQXOIJKtwNHF/SpoNXEdRsaouUKyXVbSXvKIHmijaHGzuVww15g
l7Q/MKxjNg+jx7psmQc8s/rSbXvvcZ6W5f7fJ1owv0xTdPgJMEdkcF0zV7Zv7lMt
MwgXJeiBhOEhtvd7QeqFFobS8rzbX8+khbRlG8XOkCQakrKD5+pYKVnxxLux4JRW
Ro7wwNvsYpi86Gzo9cRfhAXOjSi671ixmSLw/yr7l/+mUIh9r0s+ySqoYYHo1Oro
UuJBPbAQhbKm3DoXEMcSwz1YKBCiqjjv9bX+PodrtDrVa0FoEXrBR+RI7zutPvTX
CStMpKJYPfoYHIwkq+p4DIdhKs8MjFvyAaRuLk4ONirTR16ZcwnNVOYBXLgYAhfK
KoayzScKgmQDbhFS5UAT33EftdpXeB03DuTVMA0z3r7OXVgMAdc933+N7SKphof+
FgN3vPr7VH1VVwPzYeUA2s66YSyCp5aBZLdWsISejsiVR6UydBEKFKoxLGCzTOCZ
lcvxfvaYBTCygmdj2pLpkPA5/iiuhN1v71G7H95029Tkcqc4Ox4MdeEKOs6C9PxW
sQ31na0lJezexNjRpzN5HFf+VckNyxrEOj9WYt8dkpfP6KHjh/Im1csOUlzPlFYm
++7AcmBhfDWFyPa99cGGe7KZ7Cg5WqEi1mKQuMANWfPI5y1f0w2vDeZCiouRVXQ8
aoocWvFo0B6VM9CPTePv4CdjogiOmovKDYsu8H9qVC7XmkcjkVny5gsKcjlm9e8n
96CteUdfQIAe+T4OwQsQM0LpcSTuPgedHhbApCnUBJW8vYNBbt+RO8FAgOx+cGLw
+6L31ykFI5HRSWhr2T1iFAzpi9LORgkkNA/8EVizAJ/hCYIAMIV0yD1xFVcXkYZu
7HmjgQiVtnzFGKqepNChbsUHjCNuGgmx31x6nFj9mFo404lSBhoke5NWOJDnPceR
9K15miSKPcHQzLmzt0PotJm8QzmZA+RkTFIfysAolgesDs171XGq2a4eXjI2gxhZ
HlhuvSjfp3RWX5G9DjLbIpx8xjYGj58g7b6PvadsJIoNVuau+588s1x07fX/GkOE
jhNMVgvO+9FM+HX8K3zAvWneeyTy/wVsG6KhO9icoIK/Og7IgGJ5foBRXTTnEM8Y
UPpu3HQkO254VI2SMBDpTscT+28jbAETMG+jiHemjbBYm0bqTgafM6Ttyr5DiBrT
Hq3QR/mkaA9jZjxr16XosH29RssbTrJDZu1cHb/6xcQhTmDK8uNKOqiAMYwXt6zb
8r9FTQpCWzVRFZnf4pfoW5sXcf6LeWbOnB7O9rx6KD8djG9fdORw/BKHMrDJGPqs
J8VvtcIl47lmsOQUMcn8eqhTK06a46mcvuP+eqEVPkggkp5YQROKFclPdGfl+96h
AMSf+sJODJnock7ivaVkAQqDs9N9r5jOa+nulCPTlR9KpV8jD0Y5aWRw058grVhz
8s6Iop2gTcgd9pFIr00lLny4Dk5QgOSfhAJYPu1ZBYH3mbZ01H6/m5wQeNPPgtKK
ZCHGtpyAJqcTEQbGYZWU4OM/qXi2AdiSdyXkSD42IG7+iHK2s9lZ6HbGKxm/ni+C
8MRvVcqmNFk1zhXjfFFet7vMSk1MaDmEBCYZA9WkMaecXKCZYyQ0ekeFpQXbUqhb
pLDbJ+d+nNZxxeY01Wkaor3h1vj8WBFC3bpEMPRY6EwxBPZPa9AUv6+InRnUJ8mP
iw07VutOt9EmF1c8ZukIqWIKur4d3plCRLdM9jJ4zPaNTH8jVbjUATo5yCwr4ttJ
JVk4zvckVDbDc555MOtQ5Px1W/6UumJqvHonBYDKdhqO3enq8qQY7zFSiStSN1JO
oVLfm2tOMtyiD/OYCVvN3NcR7LEbF3v5fYLWCO9dLIO2Xu/2n1rS4U+Hw7RzWXQ3
1zwqC9rZBpHoSrIGuul3v3U/CZY6Tf3z0i6nzBubLkTyYQIBoyzOu0E09i9fs/ig
d0D8zIZaT6Gp1jmpXG8CNqIsbBwky+nGGWOZ5sKgUOrPCiOuDh/42kRmHG3Rj4C4
kbLBTbl2QgG+jq1mg6mReZSiFQKAObDj08cXRrTawsT5Hx8Ap5YuTmU+X3+R/X9c
vIdMiWXjhw5HdH0IsFm+oxMUxaR2bx7n4oy1J1N6QTUFTUdefPOGqZfYAesa/Y3A
e1ISyttUnB7ZD5Iu+a5r7/MsfkmNNpKWsNahd2Lh/R1AGz4DnjhRfD5v0Pv35I9L
rdj4wZ38NjChwhIYE+knD9ABMMNQUxQrXoXpQjTpma1ShDD5JTAePCFek/uDWr+c
kM0iqvojFVPqx+7qeut1wF2Zcqgg5p8nSakbK7pUd7DXB+IIpoeCcoZLBic61QrM
G24ASJJ0xbMxsORMr1s5JVNKc7OisXaa5Dh1s52CzAFsLgm7s8StHciyKFqHjhkv
lgMNvNk/5sEfW90823V/haxyZ4pql0ZYHJDXrWhiuII7kItQt8lCi9AxBQ3c0ejP
YY7w5khjfYDyXKTCfwdnWFJJMgBsCiPwMfwO0OdKwcsc+54ecHc6aEDhEk5+BFt+
7SAKHJeBOv9H3X0lHBxBrgxzTdd8vEVppyJ7n4cmeO4mDnSY2o4cnhPAgTMwSaGO
A27pC442l5jwuudIl2KOHFgmDRCc5mZXKs92JujTPIaD4t/8qRFmBeNGQ+ujTYoT
i2sO71qoiVw+V8AomXkearcy5HnlmGhl+/pr+pqRNRJEQmRuiXPRBCpSjgTsz0SW
i8MxOx7vgPCYAblzJcEPXJwPnyNXCNbu4wcphElGBo16fDSbfSxyUbebPbYK1K4L
5V4dQFmB4PDXOS/Vtqvomkot3bbSYOKB8KM2zirrU8fyBPmLEUPa8k6ar3b87VzP
XpxdeVPYZt6whl5PdBfvndwhXfq0wyUW+1f5lgEpvprCGYi220wUnTXPR4BdB0bf
xlDv0HzCo+1kmk+UT4rfpa0zK5ZvozSvHJkKKx73wYKRQurK9PW6SZ7otC8qLzWu
j3JVvqkKdx4PjQqqzcHOBT3j5izkXGBdlDpl6DF6k6cRTn/otCCuDFmNo4x+MjYK
vIU0LFWgWfATUI53sk81q09A1kp3NRTZjp3wGEE5LZUS/q4uSZBd4qMUqqYyYk0O
eW4ujagf66Sz+bKalgro6w4dgfX+U9fcWj1yXQMOqIlgS70oamLGPTg08fPs3mSV
H1HyORj481/9oCakBMgPQWjYaG0gW2MlqIgfTYnwUSuOX1dtvQb2bjNmASnha3v8
ijCxjBIMtbADjcScnaAAyjlvktHuFnzQxXLYa6HskwhBkpHM89ptlImgKOzqZcRB
48VFl3h1m8+jXDEe9PLQ5DN3VxQxG+tSTWQFDj5X1dZamHiOZ8P6sUgCFf96wzP9
hN0IbDXN8EJUjFSocg/L0ndBbGcfqOhzFkqe+TApc/n690O9lupzs/Rhui8C1OQr
l3PFkhyqs28KLaESFd3Is2o/BVP7EiU39nLIN6OqFFB+ir2bc9JmYcFdcJuSLEh/
biEkMab3X5jre7qBYbChsZZiyOF7vdHucX0q4wAHQj/H6JVN32R+4Iw9pP78ke8G
5gOAItFxCIMxtWsZRDO49gJKkl5FknpMwEk9boMq/AEBF5lkvfUiiCPq1ErG0j+o
48VVS2gJavhO04sGWNIB6Ft0tTArGlAAfcNULZqgk2QB+N//lpBUr6WteAZOHr4K
P5Lry6b5CWckciaqV8qVZSyxEbEyRL91/5EOpRny8lSm0lHt+JPzvNJ+rSRaPdP5
uBvlX+GkvMN8gJZ2mNLF6pazzHi6P1I9g12wbHySmRLgLZsfy/RMRG1kCZKJXQPm
dV1XWPmo5DuqBF9ij2heb20rLHwy2HYKiU3bWz2NHpePziuonY9kSZZgN4X2jz8H
67abMp5IIiiX7obl2zRG5qkO2DFa3FxzwEjg4J0PAM3VZUGJNfv+TSh2EPItBOSM
OwtbSFKE0E3VOmkbxwESWSYctXM+v7HThubIbwiZdcGqNlTTiU6dWi/9NWCbdMGC
896dK8XDt/4kMLBn2o8lJZbS32xXjpGcLKbxjrecgkvNoeoh+g26DiYMsxxxetjY
ZyvZuQXPbgmqeuuwuMNofzpKz8cp5ePHIKCn15YbIZFHj9UkGGs1l2NLCeIb26S+
OsvLpCqW2gLlFaplLLvnnPEX+lFfkiShCg7DoCxodoADQRQxd/OHOO9m2OJf+IwM
MXABeJeUf/J5BOGfBJ3edsRIl74V54DCwBmjXnHS+3cAYUrvp2Mir+Uh2Hhtr5vw
T3HgnpWBCZJrr3NJoJfaDp+xX69AexuItXDHxbeaCUXNycEVny3isQxLTVFIkJ7n
niIQOXO6HBlbyQtQgtnJWkVjMlcKIz1NUCkzmsK0QXGYR+WU2CmU0KlxbVABmuJI
o4l4nZn/m84jnzIyvaG+f43j5SUnUQYi3Px4ZD3sKr0Jk3HmKQ9dooHGeYyp9ssp
Rqm9id1egLW0kShH4GSHWNq3uq0vWXpuPg3BdYwRSgEs55GmwWb6/et73rcob4oW
rOR9HkdEmu2Xoy14vZaU/38EidtyoNWM72Z8oJWBbN54lmSjFAje5uvb0Q8TReh2
ODv7okOliApZGiTLcINmWLEdoGj6TjZvah/8WLYSssWTMol8PqbrcnZ2wapEJ3B5
vA8G4EKhQwNENvBJYlcWw9w/GPimYVbdMdjKt0hV3Nkw2ZLF0sCdGnXbfYo7bNfF
X+N2+yAe5w8DMeWIdG+1yDINYin6+RDrsyxm061GyvYNM3N7DY3yh0V9B5dSkY8C
eTXSNAKQua6iDeQkTOTQ9OO3lsoP6F8Q4fx85t0PyW5RTzQLpM/crmwjwAeiOYOU
gHcVXO+W56y20xNo8b6+nRqkmwTgT5wOlu31rry0mcU+gMIuiRISPjpjEAl9yosD
VmAlL+x7ijWk2bpeXaWGix2TSCSpMYZqM6dq2TZ5+gePaYydRAFEU9cqmGCikV9H
fwEV4gSWWXrt9uU4tasWGw5oKf4/QvmdCfeOTZs/POMppNNXDFU5456sBiG2Hn2y
TfXu8qlcYZnWB3+Pd8zIGD9mQpCjwM45p8uzEfRghOnIXWptx79PDrRIvzIctnBM
n4f6mKmlJDYv5yW6APsyqToPQUZLcmNB3f6YfECp6VbtC+uQpHYremJ1K8CzUXZ/
hLhFQY6oek6+6xTSQNeV0IJfEMvNK+CHnhYFb3Mfduk8B5Hf34zjfsPpc9z156Sl
lrxGl27C9U0pC8l4lpzZPHf3UUTFRGbZsBlG/g6Cq1521yKoWG8XQMfFZASwmMJP
XILJjMwGL6fnxkpRC6EzW69M9nYQWaK5Mnl8mLzNvdLvgOTurmvb+R93dd1VUs61
yuWcalpVvSmhmdPyhs2WINshu91BbXbhwwUxPY6R78C3yF2cPioMsjRMBm3CHOKn
wwnFdKNE9Iy51dxxqNdwLvEkNFvaxrl7QJIq1CE1zXsBKz1DXkBYAcjnd3oFDHpx
eXOwdzRlNH72osDSKIrZFpxAkih5O1vBPlfxyMfQAGBfapnO8drBJ9aWE61ODrkz
YXBJ1U2Ohy2WLiEqzRwgSSxPbbVcV4LBd/RJM+hNSWEyxDeTycH5ogPKLwRwfewk
stPd5ideVqsiY6KmGzV3/54YShpEB48VnCybaAwp2C4FOM267QalZBxOxsuCPUh/
Z8n11saHwYBBY2vBYVHnWpDNRcX27KGL4dmoypsLWbQ5ZDrxdBzWnTmoMX8N6bf4
3rE5XxfEJfSDKmc4hdCMOV/ElSOZV5rCsXmZfQyeFisr0iaKLeNkMOe1kF/pJd2E
/KvYZNo4OhJXglCSpdAYhDTDeWYvkYPsyTSDJCOl+FObcSyxsM80dnTlFQIVsVC6
CGGmZUK0RrmoyBSfc0TDuED+FHFHZ4pnYbQQZ5BlWpKw8PdfczYumMlpnGbvJSpo
+5oqltC24K9s9B3LAZ10ugznXgcayOcguDLtpH+2k/Jp5MmmNCgxNdAFfjRBLtqd
e66qlB665XCyEhqDBjFu1CceHdQQz2x+i8N95A7INn1YFGQ3eN0sLn78k+FZXfR2
aeEDcr5mJNw9/3eJsQdpFMtMqR34iFqZbC9Rz8CIfUPgg370rYZM+PIT/DEEvd5p
u1IaNWt4NTpc9+HQCsJcDdILwxIuXa7pKBBb8JGSuuIf4Q9inzbkanmHznhcNNwc
k7Ba5dflgAdSIsr9TuNvPbGeAia0e7vA1zEMelqEuzdjSRRfNTl0NDwqI2eYbKTY
wLSQZkRFzemqO/tQDm0rHT/Whwut709v+cz4hCYxMHBHGZQwlkcA9RH5pQmWKKOZ
L4iaTB2Ov/QhUjf9G22WW/AfJTv2F7vTmHrt7ADZCP/J088XwReR8yMRvlj9YEnY
hHqqF7n0paPsZXPqY1S6Vp3kPb0boI2Z7tOupFQtuMCw7mlWM4bLI1lWMcFzNw+u
jYwJbzeWWH4PC8QOyfto206RH8HbfYkyuXM/grs84hwQrVTb0W6vce5JhTi2ArAu
QlQJTyHyMTuQOdZOODw1CsQ9yQMqZGCQjGSEi0EO+CUi0zLT1ZyzXZJSr50qcmFt
F+oK3cz+NhlCLMLPRaWZqfZanvp/h8RzlWSjd2fSfv7RUU0ibw9sBzVKUOercR9i
+YfrpNIiHFVFaTqTzKFULTxhbDSYgqBAiUscPzI0CFyu8k8QlIWtVB6kpAc30+p5
d9uOk50EOIMZwIxrqzROm0jddTE9YKvarmBZVhKtFz7pT26H4WZHt2Oyk0NpTSC7
7+lOh2AospTtmIlSh1ks/UYOH2lVfew8o+/CwK5sRY6OI3O1d592l4JBMO/5eJA8
UPzOaYoai8DGJRlLi8qvCBqyzg0HwBt2LZj6phcKJzp+fIa8Zlbp+LwiK3SDXTBj
9yCCebL/974EArbotg2u8rsGgJUii1LHZr1mZZ3/5nRc54oFjr24nZ4UXnLuE8ny
Bdm/eBN7o2icnTLjueP0aYExB2n+xhqr+Nd7Z+j6ytxeNFZ3ECIxgFzOz8QwjaJp
jA5+zJQ3FSEEn2WqYq/ZcXs1Q2un38D52UywivYmEfyOmSvysHTyTsu8d6kt4pba
qsKRBrSwAM0uxw7p/bGxH1ZK9H88akJbcOaRRMa3LL3v+2UPAlLzMUggz6ciSrTd
TJ+5UQeo5LHETi9dLB9Xhn+6h9c+Fp3ZGg1AMnI3eo1QINwCDDEe6tjTOiP/EBV/
sr+r3x1Ja+UOnnfagSl+VoJZ2IicRNw7UcHd5pXa5pAukAdueidJqYcXDxT85WJq
kQ1xnMXVIoBi4crfWqJtdPO7G1ZXS2XzNxkG6kpJ87drOefo08G4+yCA0NhCTTU3
uMzHSQkp2hwqEYbAZ9zhTxqzSsGRnu2wLCqbaDfNVXAmrw9VEx2PeeHfiaMWwZwb
xDXLXcuIPgLlawp0e8B78LoU9oxzAlpFLRP51UeDmtmgl6GBtGfOGw5sFgZySQH1
Xk4naeL1ELhcDlS4j5qOREHR+LGP5VF9iPV5aH3borkKRq+pWZdOoGrM3I1l1YMl
IF/51ziwyPPBZ9RMKpEn5+urEY6pvTioEHHZvISJuP683P5+AdLdePsHDcPXYib5
BLWak8Q3Vj/l1fQoeIzWnJ45KGg2iULxuu+OGsvhUZt3Fz02gG9gEsFuzyNCM2m+
HXJf2NlO8fKyUhX5DOfrNvqG54KdxLgmTGBXDBD2KziZ20V6DBcGiICu+RSpEglK
UcY+wdz5HSaG2hQhvt7qswRqi9fcTUkDKkBUH4iBsK/LCITfbBAQHDoI4MFLOXKP
za9G3xWILEDslI7UmdR6ABwgo+kMY7+F3Lt7ks0l0Ah0ubGALOy9o9Rjtbz49vEC
n3WMPtiiS6qVmc8urGIVqan/6yeNdoGIJF51bw2MUj01i623niDiblrwUrHfwwtA
ia6AhFZHE5ow+1xFY7AJ3NlIjYwThHnIFq0SsUl4UlIas2X42QjPdUZueYf25u3w
GYip1c8HYMhsP4RncILktBdpf7qLSSd8pLRpsFFu2UiLClxOZNyXFqRrzMflrvze
EvsGIb6aNkQqp0nWfB8RZ4fZoxw2CEm/sRbJMc/nyvLsMJY0o5fW9pBA45QJJe6o
b2WWKf2A8zZm6GzSPnvqwQSxi8nOfdd2U7uQQGVt92Mk3qMD0kHrA/wVwkN6dNu4
gvJMefDLLsh6mWoYfBtmREe4MiVOBA5BG4Z3ja8AT3g1CnFO0WysWb0+WPdFFrbb
/3ilbtV0QFv1ULXywzgQlkOO+Pxxzr+mazIWwMpn8qSWEpb3axqg2LB8DqXkQUTL
1ytXjR+cENLLua2L5EzNzUkrQyQfj2gzlU1GA9YPdf5Agw2/iudyKPEgCh7iPud9
ijaYEwPC+5x8M+dAclZlveY/NKSzdfoxwRDNosI/bfFAzBx0AkY3oaknqypNNikw
/HTI4O6LRuCzhr+DESbspE+3AuV0c5kLk+5W0FeWZJY5aZWOsGnRW0rDhHs/982N
eWs/L46lX7t/HKnr3GibAWciVzXIL+j2rg8/FibOuVV8R9Jlgtmpwj5B/adl2Yli
TAvVzXxRbtqF1825a1otGPouTUSFy2xzplsLTUZAjfS5AuzCQgLaaNixoFjv68ue
hrTJcrfvz3G9cYWUHLysZAVeUD1HbTDmax5HP+SGviLmvQ5hjKxwn9i202E1tgZX
wN9svpL24H3Kb8ZOjANvvZYhzi09LOPdYvKapWHKmfUaSVZ50dBFvmq2IA8AESTi
1q+a+g3IyjzhgkqrRixSji2rPo3CRvK7dXoYS1AK6M7IeIiYxnUL7E2PfeCs0mQ7
GjTax3ZS+FHiu2m/a+63jqEHRmQ3plh5VOp5Z0TSDS5gFhr+RPTcQJ19VNcZjxe2
XF1pEzzZfUsAxtwanD/aygAd5pv0yuLAvflayoOY4OhfbxAmT6Rd7FJCpImk/sqe
QcOHHXf+rSbNZFET/EVzQifotsjQ9Qjr3CM+PYI+UMGPPGBda8NgpGPkKwLNu4oA
8+6oDXX56pg6MB0sxej+CxscFeHmU//+duLIFezOkndmmxkSVw76ls9Cx2NQ+cl+
SaTYVu3fKaLq1uDUC/2HviawebfLJzfzeDfA0EnYizdZsYWmHBS2ouPsvCGmaQnk
543CwxAmhYhWrq2QyR/+IqW/WAgQotHnJ0JOuarejjZBdVnAyY8MhuP25PaDVVLw
hEZb4w83VgxuTTtq9q/qmCYr7O3Nfqllh3gceEROXy3LE+/pBkAK/tNv+86BoePm
eXl4CwZZzaDrGDETQlKn6z41cfJ4cJ3NYXkjF7/GL8T0W3le//2YjOaAlQ5WrZ/4
cLm83qpLsGvNS7d0fOwf1VK8zYg5Xivv8FkWt0/8z1kXsHPeOtu144S1W+uveBUq
FwWFbUiTCukBDyHnikAcjILnXswhor97NzJoTN1kUBE1x9Twz3/zhiHhkMbDAr/D
O+svewFDGcD8LI5iKJlfTA6Wv6TAu5Z0frYfD3B21wfcmk+mkNC82RlIzqsPAN0x
KkriNmVEAXfeqABQamm1lebx2HivuUM8GgTcDp8VF8qYY2rheSI3IZvFaDmDn2cJ
1KBlMeAD3itNVKEytNRqOhcvvoRf/kXtMKP2C96aF+GG1L2G3a2ilKxm9cUB2Qts
pNRElQUR9R0vOZ0kBe4ry9Gas2C3PhpM13SpvO3GzJ+RCon5yEBslp9fC1ZJdIs5
+TZ84oYqJOLEb8E5dXyBwRaYsWXzCta8nMDsCGnrtwCcrh+UPSmgapiBWuuDlC0A
A4TKQxesImhtLPG4Bpfvwl90u05VphZSJiVzffRDIzFweQ/7sv/3+le8uSRa7LUB
VyVULl5vbSAuZyjRlBqzqiE3FuRZ2MlPc8cxVt2gFWUC36afMJU/qPL290hsW33T
HACgDiVyiDrRLq1eYHzVxbFMPQcqhGaKQ19rvLJS6khVeWbi2VKvdUyfEt6vMNCW
5wFPOBonHYSnAesMTXmONBPwtsOvKT2o5bNBCxz5GmL8nZ70zKHoIUyEJT42eugA
EiUt02bCGYl5qZNj5GM99J/4Mddn4gxvt/cGK7akICSSRmeCFCYWElJDeuSd6pbQ
2MaYe0L/+n3wYhieXXNLfqfRRmPvro8C8rdGbVmqAvBVdvFcyMZmmH+whIfEWJcN
JKjIaLHDo0M5ZpmvlKdtfo1ZOTEM519iw+q2UJHUpZxEi+zLBOdc3iLRcmdTXTzy
ED8suol5jZbWXxGAcPfZvsUIBTVE4Ydai9hXvSVfb4wgs8HvlThuENNSSpYd95FA
7aycoZWqbJH3ruqIdQac48oKxBwXhMc3YDpSLhKT5h21Tu7yDq+ScN8AxU9eYUUn
CIrJTRI1zbxIGLqtU9p583+5d7BD9gMNUghDtOnJnuLX5Uo0jkHtKwOAvuksRlxm
hNiyc812QUhRF27kyLgVqRBtr/rCkBkAs4+TL7WoHC/cVSLYRVIEdEndRoBDCAe1
OBbKMP69dU9t5RRcsRaLv3kvg9MSO9MLjpbxacjXroglH3DJq3pwmp9nI7ZZbm8F
Pf1AUxTEwcRz/gbDjgoa1IZqAZPH75zOZCM6oRqZvMkLr+SvA/a+Z8I0JK9iqe/d
2kueIIJfU6VHKSNU+iQMJwWEvCqybXZbkKjWgytsVCyFsuZFfPBlcoGjq5Hz8SiO
BihXo+N8PNsbMOLMhOLEO0mwk77XfKZKzfZrIusyyVPgX6mEYeNDOqWYL4RwVj0r
u6YWsqztv69tgy6QMYMc3IHSZAO0GByYG0Ea5XlGd9aV4R2y7OGJnzOZ8T65DPTs
goBlvf1BJX/Q5SrqxdZ+W39MLT/2rBOJQg1SMGdp9HcDkGbl7H/IKbNH6Q9GPyL3
Bn8HPoy7XZV5lzZpkGBVJZXkHXww7VVxYhTWznA+p59gRtx4baMZYpjUbnmKMlxe
zcT20kXy2QHdQFUXV0ksyxQsRCemxh3gUg93r8GW9PP30vrybbqYpF1Zv4SoRbI4
G5QlYzd1USrYUp3BMew08YXNnwRvER5Ehw2F9ezlE5hXEGdo/bOBc14r7NbxwtrF
PmtEdIIMihXntHdH6aODtx8hQqhxUtOSwTU90ZEft9UoMmGda9Kn0IO2owQE/Ban
xw3I6qGfj28/9w1LnL2WMKkeXP/3oOXnxpam2ruKtTVw9t0s/AOWNYliskUqJQ4U
Mn2Xohm/SlG14VbGv7GIzcSZUzwbKhVLqodOLm56axesgzkg1i+26qF8Dfy3F9Ne
OcfIFt48f8BW+OL4IabypZZktR6HoEgKQhpPUf66wY+haIpIQ/QJpPYOlyGLCx9+
lfJuFTJ3psg0BC7SHbFlLh6k0I/Gz+y86unSGBdND7+FdWdiXv897/2xVZ9VD/sx
+Kz2ylh2G73JarGUtmhWWqFLwINWBEW7t6Fh3N3e/U5x1te2SR4LgwlG+BGDEcv5
vhw+J6xBqh7VPgp1airdcehZ3VI+PDJxy6m+cd9A+UVmg7ZGoBp9fE1mMsb3hBeU
Ion+iDtQtxgQpBsHgy91UnSBgeZLhPK0+LfeFKgxzgnHIneZ1GaRZp32GehrS8JK
WZVRXwHXCn95qG+IZnRPxYoQ843xqvApsbmprLPhtIIOLWKmPPEphJmXM1SqwS1q
jJR2LUwpxugX2aZftdyiF9SP4EtThADwsG/QJD5It/EDUcZh8Z5ypeek/o76a8zN
EvJxmoGjaHrwuMx0hMbO3oGuC5N60i1QISzPXC02Rhmp1trs3sDz9W8ATa3PNe0w
EyQ1sAc/6qwFXR0DDvCKSZ/ugFVHIqEEmOMHe5TahS6y9p1lrpeNXBwB2Zgqk1lQ
IUNCtH9nKAQ8SdUxg8wK2XQPJYLBn7cxdSJL1fpXHMXtMD3o17OB7n6sT79YdtDT
9e00N4baDyz9koLwhzJoAfjyMRk2Jh8Nyj/kUuCa1ekZy0MrUG2l0B5WMYGwGSP8
c1nrWJGrS9K53KiS+IYajT3JdzANWcgdYSmUPN8KM33njTG+nerYuZHt4IXebkio
T1kKONXPoycfkGE2fcEMMwgGmXbpiT2q47/IjdUjZPrNfOLYun4EL1LFTkfky6Lk
QGnJB2M3pgGOBVvkmibrNEgwCyfYgqTCGNSn1aoS0Iu4j0+wenpZdg2cR9kOiKjL
4oZQ12spL3OdAI/Vaq+JDurVVRVEeSgAW6FRHAkTUNPa14diwkJ8fD7Y0UF7LwNK
sriIoXqr8hs16UQok9zXxqV63ZzZ4858RoM2TCe1tT0mDG48VwklxeLywbtaKqJE
YPvaGzbREWB95zOJnN1A7ejs0ivI5p2XZiS13qLak5tinMlb4m/8cnlD1eW25lvx
apxm8oodc7t7zb1D/qeM6iNk46bzak8z16z9WFyvR3enDoyQnjlTB3iX//JkAFgo
u/nT8pudmK6KJFJ0H4URS9zKbUcwn861lH4sI0RiMoVMofYkc1tuRmeV9e8dWC4d
v012V5uxxdSwggb9ONOxKhoEGcZb/BF1O9oD9LRz74vo+SOjBe6JQ/kJ8Dvb1BVL
0q7fEX/PoARnq/+KIdy7kY/rY9r8Tw8AbPnHY5JhEJATFdDuouw9AqBAb7Yi8WXt
Sz8DRG5fpIFXpSX+mA2Z0juy9kat9c3DhCfEx5wiGw2/B7nXzWtU8Zt1GW7O3rU5
2CD10AC/uR7FQpeX6/JgkW6NujudO0sG8Noi3XAISq7Q3jVvLyYUTSR5WGBAs2LZ
DxLQ6JCXxe2dUUhjMZm4/1DO6UQepvTB/P9P1wjboGJnyPdBD1pe+iFID+oOsZaI
JXuifhYPVOVqGnMSHyNizFJuXNBR4RQt12fqptdKJDNNWtUBsRu3jtEf6RkyKCgz
CXOCn8zLBhqd37YkVXcrlaF0xa1HDy0W/ZH849XVt39R+3k76/DlKNW0ZR3liCAL
qMIUaeIahZH28NUhWRyuO1Uqhcaj9C3l2n8PyNzkgKYSjGe6xpW2qq7le5xGsMFm
+RObUpR9B9gpM3DT2mxTw80169Hz/X1UkaTXk4uhB/0AsyoPzXo4Qq5h5ftdenhX
k06CA4IWMqqIF58DQVqTzyyezfgMTAfXxWcqnMkLikWgAw8vXotswSDPDveaJbTM
rwjDkk+0fSoQFEf3xCofnTujfA4bcy5b2G96IUmCi0J8qXSHdXUbyi5Vu/pBG0pH
1ZladVpKUGbj+ZnB4eLHN7nRz7fj3Ykia0MUedkZjYgob/xZ/rFxBuvtmR4A+q7K
N1LwXbFCl2/goAxCVrppx+qG1I+Gn6uWd55AU7RCr/TK7IGmbPdclTCSyszK5qkl
Eft/tvmGWCC5lz46rwXMyA7pQlNUogrIHmUT/p8bb7wDoQVlLq+q3jS8gqdSHb/E
4Ba63HT4bqr3DU00HR9B7VX3eudFgUAS+06wXkNseaTEj/e6ac+ZyzcrStS8HFUT
z9yCJhY5vahu/3F5TJUVWosbzOW5K/oQj8m6qQ5PqYc7ZnqEV+z+ud0jUb/ZUxYj
+SiYyn+VRiy28R57MC0wbJM1n2o75R37bfSkBNacoKhXn61xpIIrpMC2WtNHEEtw
CHqSC0QFcN04KZ+zVSSYwv6ElbCzF5LNyUIXK1TfVLlFKiiwEMQXS13xDaEVlubX
fRGzxWtu9EYpBho01VI7tuTdWwgcLrVuTXiHM5tMHTeUBOhgu8XMElrQG5BlcGS7
CQbwt6j/eycazi3ohJpPcUFkELQJMDh4sza4Uc/Yudq2ot9YbttV0pOtXXCAaJ90
9TDhyvzJI6Bbr9e3xoqIjM5XawlfL6oGRlA+yyDO3i+lDXvaOONywu0dbFN0l+m/
yx4o7yIZmChj7rl6kibSNbBN/oD+eZXaiNIh/TfQdDBZSV2qtQxCqWCe2IEHUpSw
o6xGbiupLJDxJezjIpipu6aK5xUQLUBhVWAxV1L+5YTIKhIsnXUmJdTBQ0oRa4bY
p0D9HkBD2+wL+7EpXG6ykSoSiE5S0G5QF5ThdChS95t3NOqAJtZYpZDvAs5yBmSZ
1k5TxwAxJOJUQWWD6+fO+TBRSQSxeDmBJksMGyXwpXvvyWOYJQ+OHP/WziZcg5dx
nN2fJSV/rbW7KkhZam9erj+Gnp70dXOgV1cxxE/6iJt6wxvMPCg/Kbv5KCZ7k7ag
Ayk30zswMZO8Zp3uR+h/Au3ukhPTrtJoiJxAMbIgPhpISGOaD4ld0Rl9r17PIYie
6RDQ4vZnkayqklLHwQvCwkrbfDDgns9ELODOvz+chQ+P0kMUDIjcuNp4XUy7Ne9U
ak4ZY4nhtN/Ga7HV9KXRqZT+wRiSF35NEOfOaEsKQXLBuooIp1RNynTb4Xq17fXU
5N6ReJsXaJdmDJXC2IiVhPL+L7vT86qOH8K8Y0nSdWr0Og11xpS/MhB8nE/c1wjh
z8X4xzV9X7MYAF5wFRy2i4zGCJAcfZoNTNWrDSOdHU1vHVE4X2CJFh7d7xWCjh0w
vzzPfBdQdK4Urxx8E7SjtqZC+1Y8DRLmbBkzJmyXLZqeQKgFfICYkekZqnkEyLtg
iA6f1p7egPdvI32tloEV0k59fDTweR1j6KeRvvZsIO3+/vRjBM8/LuPSlAEm8OQO
S3d9kJfBHzhc9/Up2D2SKJDM7p5efmLJH2Es2nIKKyuBPVyLEo8SOMDL2c36wb8X
v/mB1WZAFfef6E91w7UaqpEHOynUAW+LRBGcLrPR7Jeiwg2zdo72dyFEwbmtaqYc
fNsl9AdEL9cyrSS/KgktBS5l3OoFh6SN8/4krK1uL9tQdr6eZYoB+oVYNa4sry5Z
slmMa8A675YzTjdvpDxwJd7JOjSsxyKOohZcH3hN00QExeiBQCv8zPFs4rDB9bZ8
jhjikYpSGCtsoEJgMgbBTWFPleeNKjhNA0ZK3VHVihIIq9b+HquiXo5R0fcTbP3k
oLqyXmN60UPXOaVbzC1bjb+O3wRKSNW+alRRF7YNJC2CanzXvEXkCtFaBVxv1OQ/
+Jy3GtZ1DcPM7WcRKmlqF/TV4I/TqVs/shd8Hoc8h3IHrJUG2IpdVLhYLRqr9Lbe
yUUBnnhOj5dMWbiJJlT9SsGlhbexcPuxyOELAO7wUmaKJmYYQ2bCSEv1DRpquUYU
SP+pnx9Klqgu6mArjsvCSgwTZ9cD94iguiHpGSqS6jZpjn1YFFOA6WBIxinaX9En
IHRE3ZhqFJ422ma9OUwcz9d42QBg0xMc53kjbHL6TEs0X2SWBy+2/SaL0bNQ/R3+
h+s4ceS/TwuVY4HXFi+/NqMitnCI2Re8B90zhwO2R/ScIAWMVSMLpHL9jliT78qv
4ui+9YRtQYvmzmx0d//a2zK8xpC0AUavLchRbOEAETSrqrzsMWlf6xOuLRnNFEUi
7yV4T/17+Y7q4ZZYON56gOuWwvBQ3yMeLaOULXhrwGznz5GW+96bF5M5f+93BpSi
oyzq/YGRfN3uYu9wK0qJT2sV3RR70YrYVhOcO59aVqDlH5QwvPUH2ileHWMc9LA7
OsDFjuLGnGvQjRpB3UCtwSWZkqA5kJOzARp/3umzNId7gfdI52kX0ZRrQMW8lc5X
ZS2Ailz7fSkqwLa/sez3VbtA5d28pbhRVkDdlP8253BwpMo+x2iweRfb6euSKw9y
xO0w8qQmpJMv937Sf13nUNrxs/hNRaczvW6Ptb9tbO1OlFGGzCCzOhO3GnDKSlrZ
ogUiI89shX99hCg5MHNVI7UOFx75j3CxrdDAB75mXNo9TwZRQ/pPVWorvvqhkS3b
zWC7POdMDQHaWIM7YDYQ9Es+QaU6Uy2HJnLNjrz0Lsoh8XC/jEyAdtl/ntlizCqN
emLDL1aNh7ASPJSYepgxsF6ur9jn76wHppM7gNLyqrvbrFaCsp/R13BBsuO1Etyd
TzY/7EVQYe3xcEnu/PcWzuF0OPjn1Hz0orib9h5hR4WZSb83zEqngIcpPM8WBjkb
8MYuZ9QpR7c6frWRUWEI75WOSCZ/Dc6TJgn1qAyPm7fcfmb5XTPkypM/3VnY+5BU
2Spi+3jDr7/Kp4IOtL5gpOvfSQ6J5NupU28lwo0NzvghgH/OOmTaQ4jnEU03zLeo
HLlBus5MQisqMifRJBS8/evUaLtqe/AipmDu311CBzkUlbQ9Eg+KJ9uh1xFr+HnX
76KgVFGIXcoKkuhj8+iixvvDLm3regsiuBOlqFxfY085Q1C/2zzoyuVFXSwOuyic
ZXWgQP9HrK4OYzzF962zRkv/F2vkf/bRwPCfXasyGQOfWph1DpPhU69l6lGFw0P8
No8AkcOWMl6w2g1F4En48jmuJpx25wg74wb9tVKvHDYCj9o0OeBmadNlO6XWVJ15
rxV1RbBRcGnyWp1bMQViLHK6aT9Rfm5o49JoTd5MN6s2fcTk05ftb7jXFndvgc/Z
xiaEdp5+qnz1lN5U1C9DhRnmceLo5ggHYhJDk1CsXv9tnaxbpAELSf6qhFd83C52
qoNB7dX40Lb5oMPh/2fraJ1DSulDeGwOXJZHwnm9ae22rJqnwuNApZzrfpArb4KL
8sdC1TJo519kauZuXH4LqXheOJ4X7r/iQMhFXBXpznBK4opZv5Vnk7dPZKwSo1Qv
L/5SYXDtT/fPuxizZe5sFN6rXHeMbf9/sumU8KUc/pJtkc7SZ+2WE86nz1n93nwy
YwRAIvjl+F2CBzAqs7eWR/D7LrQ7vFnO3fP26B5L1Uj8iWdDz3ItoPzrtcLDNsH9
zUQcYGeWayMCWhAiplUupomwUYAFU0kqn5tGdvxBbWgzs5NMSuoC2taPql1OKtMW
Wo7JkeNWTk80K5XRL8m8mZfXNFEVHogktKw9pGC67FGL2oxXtGx6jDXdbggHQz6+
yqUfbVUIgJIENtjIKdRfF0jBirsSuB9mN8EeVOZE+wj58aU1Q5+x9ITHL+0Kq/8O
kP3IoSOAGIBHWvHgRi4VjiYb+QQPlzEkkcqeKGoKQK+bs9QVyHCSNJIPnJqCoZw9
uz+eTg0jwQBahXuKwTLqGKAAk3juGCjGfClmLzb+7EIU3e11s9w73VAMfo/52Tdj
sp07bE7vPnFzg3uFhaCv10I21JPlntKwUMeqirvtKhzBm5lVa0pLTT/5vups9j2U
RICJAgLs1q7o5eXrpDhaiFh1BVbR6VN52cWSSsjKPl/eWTD38fsqmkOQeAS2m0iR
xn9/KZgQsreFpVLWyz7J8KLsNvRv8D2m9TYBm18xG9TR9DSGNqhEcTcTWvNeUdyS
ID+7aVN/FWC8CU/rL4KgUNTyuBlLwW5SQXZ35hAO3LHjB4k9+jzCSUYGtdry3dW/
UqFXKR+awHl0qvZbRKzkSsrnxjQtr9MGKqbolfCLLKvdaaw/BGvQ3lakZaygdZWY
2dbl/fGqUGURp1u7bwe0nLzYmbIz2cw0Xr2tXUvczlJnWmlPS2Bv29qO2nvLimu2
0iUD0Prxpz2cvYQ4EOuH1MoJ57WU13Uf6Jj+jwWCUsWu5IdG5oCuQrVUe2IDE8R8
S5Snk5FpzjtHEJhIjZisPmsnXEqCg7c/hHekn2aLUSWd9bm7qjR9J8ybuI/wMYx6
I+lVSpM9yZZesCcZFKuhI+wVLjpH4PQZDpsWcEioopHMn7Wo5Zw6NFNvVJpl/c/d
PkIiFK0ONLj90YO0cYHquvGsv7osH5ABlBot74KGscGgB6U/yCm8mMz2jPGl0SVt
xV1E5p+W3KQN5X0KLss7Z/eMqhdjyRg0h6nVLNja9tsi7zybqxVNfzpUdsvE/Mxw
vb4k/tTyCpTstVTg2zqCXxdlQtePC650lU11kLn6sv2Kj7WzIhiy1Wo2pC13fMWC
ENGVlEhj+hOD0iM31A8GUAXtE/x9GACPLdq9sXgKab/OOpEWBJkC5S59qXh+sRF4
2Yg3YVQYhCWElaJsg8LUkp2LoSViIaUEiT+PEoo8q6HDyoMFRiYl3RoqMUEsOeRo
DVyh99xwWp1lKO3UwaDwHVWbgBcXM5oYBiDuL4V9n8VoNiY+cubfzUIrBFlKNgeT
viAqvL1h5hWQ3iGiGbGMo6KDwDptGN4pLJ5cXsmp9cqC8on5LiDEDXiF7Yf/TSY5
9gOwyQyikacAiztlb9mLBndy9OhRTcl3nClFR0GJuWSSKvV0hpvZ/e2RBVcHtNbR
z/cf+qKyIZcx0tSOkif0mItDLw94nKPca0VLpFhsWaihjMGJWT3OyEcV2NBz5E5B
xFRs3krb6l2nVFu0roV2Ac1D5YL306ypAxIibcg1N1a8inetcnUPFbHQJLXJNvzT
Dl4CMebNUeiL1ShBNjIKFOY/P2ZpiLDEBkZh79kiuXlIcUor0x0pxGJOwsvkNgpz
CRm+duiCfPwSTGW4kXPdw/TkmaYGI2LRuHM6g6pmKtwV7LcGkcyxZC3/fJz6K6RT
WbNkzUnq+6crCRK4iTKrTOwj5570p5ufIJbFmP1isD0KeNUOq+iAe0syV6Ej1W0c
x+Hpmxyq131PvMdU9ZM/wy2XPZkacfqSbKLo6cCZDRmI1+28BomQYzVXBOBrRf4u
B58oP1ekfkOSDvNCcvG6HmvRGy68bmflA+Ez1LfsugsTVSaqVfOBqHii710bxBUc
C++X1UgnhYrThTqPQgPR5BCu5T/PoHZkrsYoK/DUQnWCjzs6i9BE1rKmYNoISLF+
ovET/cwVJpdumh6+1jYbEUpuOqMkzGHOAKpwavENYRZBepBbW/oj8Yk8Lcl6Pcwr
N+GIs91TmH4iz5Qan4Rowa33xbZSOp8WFd86B3KCkdDghUt22hLiv991vZUvEjbP
7QOfTtXqzbw2LRsaEd2QbU+2RDN91d9de65NfmrtXZMQi3fcYeIG7H62IRjf28NG
ZOdBam7Og29L+LxRKBKlbYfhOudTQ4chKWsWyE9XMqgzRJYmb0VvKb3WhBtyGo0r
836u2Vp2xntuoXx3MJZwGG6lA18qGtHkNwSTs8mOZfz5YKuWyrU+otf5VvicoYSW
zIBx5t84j2a2HFHZtU8H53rD3cOZG0oiF4FNX6gyATPGfqfeByb9LQQKnd0Kxg1y
9Gmkd3GfasUHoMKNTztYETwFp/b1DRKQrSsVDgOutOt0H/bLp5gvIvmyeEgsbOtc
BNUFR6B80dNBCLJd8A5TZZ+IyfKeu5FcvxboYs7y/AmAEq8MFLnTEAcwvHQ/0F3n
OajA6eFBSrf4LuyDUPWgSk77k5YAQ1b/6UdxCe2jt8RYWDtp+2kVT1EShmjHUhlo
ombvfkH5GJgudD8mJKTX74gF5guyO5ZxOT0kyemTyNODRV1nWNe3zzohCG44fydr
ChVWJ613CbIf/YOnxXfQxJ58LkqxwzNz9nY6CxyjEZsAdYKhNZafMYB78YIsg+LA
uuw5Vy1qJmXvAxTQgPDIOfOSr9pRX7wEZcLEHAFiDpKvn6de8z4FjMnRmVsDrry/
roGLzVx47ftTA/FdF/iByofkWBWYL/lsvsSsUil3baaAaSlDg3mmvIg7rHRkr1Ge
c8eiw2DXjikZfZyGbJlxibfBdbZw/88xe5GTNm+QjhlVUMujzNTJFs3L3NagWPKm
MWSOvOXPaXn3KXRSfHw51H5eIG/ZvnUX5ocj+vNxVj/VYSQPHhTbWctI/5aS7/bz
SMmb6/k3h8V/NomjMsC5GReTdGjCS2aRpcTYdoaG2KmaUm8MuV2/dfYp6tVyePp3
4BUR/1k75IloYiz5ca9HoRD+y82o2H8A6vqb/BLTqjXQFdbHGlLlrCBDdPaaf6D2
GuCjINbtMujH07BfU2Iq1XMi5Db8mgutzF3nGXCkPQ1dU2uvDVV+fhtpdsCcE0aV
Gmt2JzC2eAzLVZE/zi709TrHVCTjrjYEcK1GL2c+QksN/NLO8/JdS77uiMv8waZk
VRgfVa9ntiA8BtJF1S0Pu/B1ivzgqi7kPjcjAWXYEC6qOy5khoHhOJ35V2eDlQda
5pliifbgUuh71h00u1PURDMyA4yNl4QdLkvVO3w6QQPOlnjL3W0JTZu8oOFhefE8
efqfAQfP9Y0UIxxkYVY3k9YmAIJGyysZ4lh3GbQnQiEQD0qeYTIrgaFb71LJzytc
SGpBuu/NufVaLsyduIVgNo7WDHSVy1H08eUiwyaHI/KD0+3GwDLw2G/MG4z6nDZR
NBXiLtk9VmxQYEedWRnsJkPWIQr4czWjKMOiHVCwXwWOqNyl7CE+S+ij/7S/2srY
/pNvQGMDiN0fi2yw90IjLZVxjrira7UrO6H2kW+nJFbqklHTBdmjsr3g7+D4QWNS
xumev+SWzxrngDdUMjxtG35sLcB0KBAn17jknVE18V0cVDhwfK1XzMT89Fiu/Hth
sHFhxKgT9eEOr46lM3gGfS30/ESUejyo/GpqSdjflswBPx6hDN7oj95NR33yTXTm
meSzxYVi638CAjVI6NUqjx8svoK7BSH2m8aaBo94AdSS1kWvNS0n6wP5RIk5Ai7m
tGmfDCHimNzpxX7ECDXGW4BhXMolQxFlaU6otTtHyaexhEtlCjpqBxPYSWf7+i/M
wJ997cBVF/f4xxaBm/qfhSCuLg911SI4EbhkLNtTYX4MG4i0iLBGBUwmD1uaH/NG
MC0HaSZYHRKMKpISHHAHQznRvRd5W7QJbaApZXyZ8LSMh9wZu3PjKZF01eR8OrnY
7FPgEGeCN97bSnejJKykb72uvuGDtfYix5EaMi98EJ3ME6xPMiRxhTirPrglmI4r
/j22VsicRDwtvXlLb0Gr23RvmCdV9cvNcGC/HOF8ZAJT2wqHu3GR+raGviaEaiEY
jS81hlummEq1b8t2kG6mEckG2GJ0Xt6c+3tXO/9hDWUQquDLKDVXwyGV8acV+aZk
sz4ayju6SILslzBzQL3nT6BsCsh270N+KA7MjwGaPkrU2Q+vT1qTIRS9iJZ6cLA5
N8j5mrctWrVMUIT9CfakYZmKj/CnwCsZdq+6/14C/qa2RVCv/v7DAgdTOq94umSz
zhBAjVbG+fQ7Zadz3JLESiViWQtb4nqrmz2ojzxzn3Itphmh97kJUaEFum8dCM3C
FNZ1I8rPr4oxC07Z4rDCbI7xIy7CV4/BjRDKUUCx1Uw/eyYPpeFOZQeg6LGtf197
8FbRctJYZ7F13K0gwoniDO0sSVCmKSPc22TvP9HPW4Qq22Si8765X/90IrzSVv5J
5Gf3HF6XenudgY65ih3qpDI/ofXmwT/nHCMBYQGg4o8UmyxSTA/6qKvi2X3JetW8
RE+oHop+yFrRn8EDtpqhlh+onwdQ7WRhNtKH/B5FKey9hEc8hDYvom+/cpJmq7kJ
JFehzGU6gLrg7eJoCf5xjhK+1n0oGRXSc80ZZDcQGuqqrGCtGfL8SNooTGvVmCat
C+kLpaSaTFTGU6Jyck2yXGzg6dVtE1GdsdqESYWohBeSFfwEuxEEvDGvXLKPbwQY
YBup5PMpZD21+ycpdfjFos6IkZ2acrLIQB5QbybSPiJgf1mhL65KrGXnJwD4fpg0
RlKCZG7aaYFOZFJQunWZnhezuFIodKb9VddZbO7Y36fX1Gsp1Wm07cgP6NZzas3O
ILxsTBye3lvM0mMGtBdIO+9q/Ayjp8FioCctxZmjywYyVW7XEeIG98tldX/a12OE
gLhCJXzM2rs4qcP89CMEXE1oPep2npcoDiuP39e4rJObY63XfbVDRUZRi2XN5P+e
CDkQxKRC12v3qF9oqrDn9t6OfV9OCD4RLMDl3ZSMnGJ2Mx4TZbiksm/WarljtkF0
OLYc9rzcGo2JAIoEchkHOTl5qjUv5entoO+Eso/y9SzuAgM99MQwtJVeCK9cDsdD
uu/+XrQvM2khvEZo/ZgVQ39kLBk2ltSWW2EFhveCIER0ytQUsAy9PuuoITEY0yzN
uKzRFeWuM9h+kXdD3sihnnS+cvU+1XXs0k+dFqe841YPt6Ox6u+jzRvB+wEjsz1S
jlLrc5LsmDDzfhdbRja9p8Jj5Tw8h6UXakag1FMQWH+bfP5kcMHVauRkYbeAxqAB
14DudJX5dsaz1KpqEMywgLEYBXTgIyV7znO0dLE0PN14OIN9Dr2xAJ5qPVW5YiBr
v4MsV2qbg+mx1Vedk1GMkgafW2yyNa1SAfUkNGP48HnuiQO5UNFrVz7eDXOppjYz
LzNMES6s7pPidMRsrM8FyPOi3gtunLx7VKdCcIcbyzbpgZwjYfApZIMw5qmlmI4l
YPvCs0cWWR4xdkGvK9Yl2GGAm/OUj15ZY2No0xYmRXg3RG+7dSTWj1nmKMaNBJvD
8EOZkajnfhENBOwTX1T181fM1rMKUMG66GXGezk52u5pVcUBH94d2Z9drwD9082z
fHnkkk+pRQPLB+xYhLUbNBBufjvqGiP5jomEmB7KawpLThED48NFArL2Ss5XrBXD
0SAy+SrAb7j1ZLNRBMlvcM0k7KJ6kP/39y8l/Yyu+maYIVpUB9PL8N2IeNOKuFoc
kfWJW4JdPkOf4818AUbtARELL54DH5xv1A0aHobkRKr+ftF+gbvBgCLAVuJHtpsD
wz/g17FjI59ZXG4fsGm2ITqcos4bprA64PyBoLanpAL5c7SIB+VmxQHmqbn8zypM
Iww4fhqNc2Xp6J0OIWjU50xJr+12bc6HAr3iAnd2xVt0mi6RNwAg6qwsTZKNF0k4
bFopLwoH3zOpQCJjMILYpp1s5UlBn2qTOWfF7ZTylDiL+FzYvRYGoQECyV4BAEYy
xFUNyHVcaAktFaDU6BeIS4tkrwt2+JQpbnPsOxBnYCAkoSF8x5pS6jditX4/ZlnT
RN/9Ip7BSsv1YqKDPEExauFvpECJnEem/gPIc4lredIy0jRxTakNRlFuc36RtgOJ
9MbNT6SPP4iPc8FI8cm0+gcdpRq/wC/J2BXegLpiLiafScNWarzxZ21XNNf2u9Af
z2x+Uz/qUmJ2NNOnC5DC1/pZhg9YWF8G9RuUVyZA+bPav02wuPZWuTQ2hWSIRaFd
gHL3Ei698rQ9kmq/gg5InH1p6pfvOlO5bldbcP93f76G0Jxa7iHMseFGKCezYGwl
WIcfVlaBQTCxutzoeqk+niAPt4zVDSIwi5o/JXKxANNZefsonH3jiPb6CG8g65gS
sXiqPrYyZJOq3I1+2vLdSHLbYVbw1zJEuhx+D8JFTHQ28DLv5H/ammO54cRUFNt/
suGVrH7jEStTdRncl+HKVnJfperW3E7wm0ledVhQXxmDHxRdiCVElrpQf1tPGf43
i49HHIo9efc0Rf5u2JxcFBRbQQ+ifQeYqqtpC7vjfy72ap8cICeoFQGxmFTybP/6
vbY1VnysQEHQ8PPTqcEmlyOnIjHbnHq6UpaAvnzIQ++6FjU8y0yf7sj4uUb1oLLy
vqhYVe4OrqIepXxjFL65ADvx4fa4fUYYGXtKJBIJYznT8MIVqgMEdWSNb5ipUVJm
M6Z/8HM38J73Upx4T20gIFhBkOfEItz7P2SC+DmdOFnrl9Z2OV+4jSv5+KTz/i+V
71Ip31cR7TylXHYYhDUsg5ChjlRuHnGMoo4Ym7tvcssTbp38HVkQdqaSJ4lDUCDk
H8unWFsrHHgDuvzSsT5Eio2Popwn9QUs8HVzBkbmnxQ/yNQMPAgJNEy3Tgatdcg2
U+5OGtjhtCvnwHKd8Ca9P2Svu+WSjKvqbytm3/9L3g0w7mtdYw6m4DYnnl7AfqPJ
hhUjwUmCLSgzlEcqLPigMmzwhyacy/dY8XZG1fdWrwpVZj2BjGEerJrkhvNRfspL
OvMqKdLRb8USNcCaVERevzFne9HBISzLKZximeozw7eaIU1ZHpRmfdvTef9XhLt0
UnDg05DWjuyxN84bvqS8bhfwRam3OjNVDJ+v5ctC6JUh4tbJt3K/cfhZUJgOeJ3m
5N5lh9uxZL8618GXZwkW8xXNVB6ToVI6iRoj0Dn6NMcriXBK2fgcOBGw+sAuDjs0
Lt0J0c7ru5MXpBeSWNmfJL6TzT2ZxwghgxfbuSay8bwOraJl/7PTno7EjezlCvqI
K2sWg9HLRqJLQlgSa+FRYHjifXHKBjgXtuWAsk6xnG3AsEIlTkenrAC9pmBzmuce
qwA3vmQGhQetTCuTTB8FX3sSMMggVMJGC87XhqhV9IY6Ot8H7Qw6B0g0EBnhLBgy
ds4L+fFkSVi+INUcCZvV1DulxkjqJ6+zCROgzn2xAeD9KwQojl4k2Oigp9AIYnPV
3XOiPvuapACoG1j5OOAtXqxZpsYKZ3jh4EwfINIuPtm4ptB7xtklYD4qOnahanEa
obcAzGMW1Rez19lhDfGUP7I9nSA833VPRo7XG5jc/vQa8rrdPep/wIGpLWP4lHep
f9Lv9JG2FEbHzvX2JFuSuLLB+GD3yH4pEWrEzTkVDh0YCAIAag3bFVDmoMiG56HT
f6Jd8Vec0dxqF/S4ba9O2Jr6IAyOKehbADxGR00RAgk01zp7z8Zn+yeBSWjl+HH9
ijD0aVF+T4aHvGKVVHb2m8e7awC73FZCpCHS8n7mjQQQFm80JbNwGaJfdfoVb5MF
wvBKXU5cofWcpB29YF2qAoov4zJxPBrOxjHXGxLHke1EB/GAbkhN/eQkV5oqfVX/
zEPVu9cDOoJdtCZItzzpqpA3oNaQti7uieRmxJ82ygI/q2H6vRwCTHE7q6FxzQnM
fsCV8chLZq/WLttDU/Ccbz99ZZHJn9EtbiqrcvF7lXVlQ9+l/Zuu1LaG3GfllKb4
IOVNpcKe0IV+xin+CAI8SDI3mequqQdKBxADrTu/No3ckH/ny5mbCEJ51n+w82Pv
L9gwWEHzg0nz8PrwBERxNGK/ZBbzNcsR0AqYDyKO82pVdV2a+2q/fDNhrQE/Iv3S
4QOuXi2EVG0xeT+lrNWMptYEYnIe7SRgVEv6GRfLbkNkAlvqIimJKeWHdxtocxp+
pomJandZQqP5nWg4OA+2XxrnPyAK4dnSK2L+AiRK+AjgXG39FqvVcFOAWE885aNO
JFT8U/+BYVwiEpDJBZQn3Csv3B35VUjuZV9v6DRLQkOI+TYjTB9urWy0VAkRtyXI
drIinQnPQmNH8Yel8MPnRXMruzYN/vy/YkpDLA9ejFKJAggvW5biobN5ifCgOmSd
+lV4HmXqs4iSMBSkVg0wyj+CCkTYwR3NogW6U7jkF3M8GHCbzHUWvHENUfNgM4NY
mH35JB9ZrQQz9E6GkgI2GJsemCMjMUT/RgTtdSyXlRyF5U0paQNIInue+inO5siB
+61jL2HPSJiJPa2ZvX22b3Lj61KE4S3fM3gJSePmAiZycyFf2eF8Fq1y/fFT8z69
rGfqrwMA47pO5GliadVaZYDFiD/XtQDNZ6sidOPpUohV572wmjkLV5jXfYVEoxn8
cty5fKi25Myb9o0t+X4C/eipaK+FFo3GjomkzhbDh/Zb8bh+MaW13si5Xjy708Wx
MNhSKc6ByImsHwlZudWoz7I2cMj7HmU45gmieAzgqMOSs38td16f+hvq2yyFY1rM
nABkf/ClYUevBYtK6qgNU97vHluhPrio31ptK9DohnYWj+RNtwINlskf6HQTlYdv
VikkrJrtyzeHCh8IwNdruhmPc5gWDdKwzQTL7xVq8g8GQH19l4B13TCy210Q3WhC
vLLiiOBoQ3RLZraZGOjUb6gW6o60ZIZcnS+wQqCzrwYcc6ISNDJJp675OnMOAh6N
4x9BzHDuY/IJ+sgWu6V+53WEyLBvhImFHXFQNiiKrc1HKpjflPmVVA0msfMts+a4
u+I7Qmx2cHgsU9BaQ3Cb6gCMTRkY6nrPLxyOiFOCpQkTTFRb2qruWtHw/ep3n6DF
66Lu8c0/DHPygFq1m0P5ruAfXZ17RnHZnPWIElkNA8J8GgWIiv2pRDrcPiDQmosQ
1Cts/L7ayTT5q4MVt1ORDQSvA4hjttY4tt//UBnSCQTN8S5Do1U5xOLZNqABcE5M
HeEDczscij5nwqwL47eyuGJSdB1BosE8aglkTGio7gZ/1lSkWyZ2pFfRwyehpPYy
D4NdFSZji/vbrh5yIyCGZtp80XZV9ml+LOTcNN3Mdpee+KkWB0XQKHIZ84QqqmWf
OyLBe8x/YeJqaVvJX+KPQ9Ro/zEf+uJGnKWbJZPdai7Bcp2F7qUSqznePXv38Sve
W154IeaVycbYu4U5TThIncBU1Yf4xyE7vgluc97GlRQQKZFpWNsPZubXZe90MF6c
KB5ZIULQfhsO9efQBHzBFvb5LrIt6X/qFqydyS3xcLjJ7iQfW7QF74LOb+HrRL25
2x8VZ+FhbhwxI8UTpcB5kBgx7df8KCh+uuQ0CgPzGs8Z2CcK3XpHVC7rpwd54XnW
SCcwbULFkor48eUDnYVpq0wVTYEvSy2BcgNHn2WzukrXS3RDzSfVjiC9wIJRwbvW
8FKw4HuG1dGXAP7OrVg6+OXrptdhUXE6pmItSFw//9PphuPT9uK8vKimgEkJITpo
KkITPvU1awtV8Pp2BV+pN+qRy4PLWpjtFjMwbopXjlbMTq552AWXbGoOgkGcjahA
TxQ4yltcZ6i3bMCmac+XC4mWDzXtXNcQe0lWkJzrpgJT6r0TtZpRwoej5Oez2tNv
cG7OkVYlhfEEy/Ql6jbI/bZexxSH9fDlvyvPGsDHh78aMkzY16awBXXwb3ulR2S0
leNzFYtYpE3KQ4bBgC7sarNfPB17yMGiBwDS2Nld9FyiBBjU83AcXONWDS8mJsoi
9th/kDbz7uUUC2ZhXlhRHY5ELJ+VuDUeqyHdQcAIwmmTDJpxhWmzxhF0TEIjL6bv
wF+iZqQTCjpfYdaezThy5/zZ2+KvmBL1zmrqT9EIrOHwlovnlUrjck4B9Xf/QzWy
CMpSBgY6CXMJCr07wql+a+1lrG0MaRntKbBY/bHTFaYExwC/OLtIjXzOtKA9dPVi
Dunsz5X64VJDts4qjtfwbKU6rhA4CWyCs0y/l/jBn3tsrdhPZkqWRAicRZcV9KUo
dtKh9SrWkcDTdlZWAwI4Xl6VzP3YJKyJooZt1cuft8G+wqg9p2WzuERsKcUhaz/I
QTcwY7YwVIutc8rcQit7p4HCqjKhY7WUHmnvhN2QVFmowlwTecCR+zdt24XV6RXW
gCmVwN3zComRoh+pU1kEV7/JwAVx1HCA5/rFAvwzeoK0eyaNXSfTDS8Iz+IzyADL
tl5QwaI5P9LFVb2QgHAfm3saOdGB4NfzJ4JHz0jOXCFlBU19t1dsayTWybZBvDkD
nLEx5Tf9h2RnsIfMrjSckmIorfy9npgl4nDvG5AytrRraUtpnIq3qa1PfDZCUR/+
JO5FtP3nKygw4S00xAEpDgTTkdw3ugS/IgNq9/mu9Mm3PhX6Fr021GrA0ajLv+8P
uQy4pA5mdtBL2BGD1/HAF1eitOeamT7CH7c1EGmEJG29inSN63/MFMiRxSORXlRB
H6rwtsDTtU1irWym+vAcneAmZ1zgXuESCnsfFYu85aFe00wpztYDqxacar86tlDe
Jmm3fkC4zy4E2TEKwu0RtoqFQ155WTKS6WzOxtzZTcARKTso2wnDvqP+Xdi9oxtO
MP3adKJUfugE1XIDnUanEl/YIs4MN20vFEluGs1SNuGaByE4zsBTFM+PFHa18hDK
hdVD6+ylau0ZxbF1sWZokSfv0ovgnCOBLkcbDl9kdMf1WVQRxb6EmQNwLCpVeiIJ
pWRO4NYL29TwvVqKBMhzDin7MrLzd8TfNt3ONSo6nyR1t5k7YW4z9D0Dkn63hD7G
iwiSUNFtTjCuKJ9zmOOl8GA2tw34o9Yrp36RPck/LuEY6DuX5RdqsT6I721UDDvq
EYwmDzlvK9OY9GR/cRMBwqzmqYE7K/mgmaD/BZjWx2nRnaZinkkg3kGXEq4GDDkn
CoE/ZuBKV0Rh0p/jngF4FHxqhmY+G+Jj6i4IqFDxA0i6cEzTl1XQuuGB9kPbzIa4
gHwEQkfkwqcn85G02AQOCo9AuMexbNCVXR6HQKJRj86RbV5RblDnx3W9hkQ1F5Pm
kei9FAb15ikvoreZ+3EmYNxSd0sRWISksmRDHgc0zAR5OjWx+Kap3m4pUuOk0x4F
J1ZDbtHZbhWw3ugr96coAdAhq3VBlyRT5jqYj1ehk7QXMMzBcSUQnFI7zmC02uE+
CJK+it36kqJRGb+FIZ6ydP6cdMwpR/C6jiqpXijtchYCr2BMlZETR7zuza4PzJkz
YvwaNE9dPUmrrUjubcbLQ9zhsQFhWzdCDbcF96EQoOD01VISCC68xYcZFbBG6gUr
5dgFKoq6egaXBDTz+M+dywTv82yIfhKQsIkYUL/IpEoT+HYfPaj+aPxz8ctaXH+C
2UHQhfDkGpUxvob4Fxo1qgU483bxz3ceZ3sNIRP5xO2YUEtY/TWL3U+d2riMmwm3
RbV/W8W4XmroVtdbNMo2W72odZCEMp7v8aySbCA4UXBH8oAKKFngbSU37l0UFT4O
RUMknbNQ4ovoMO8VH9FIlygH5z3U06mDG9sA7HAke5XvUrauKMLwbE4jtVVCw00Q
DByB1vf+ucnGG7Qsl67jn1Ui4jMlBhGdKWlPnMwiA7nLl2oHoEcoGBmdEO43xKCx
UIc9gY1GAs3/slPI1ase0UnoMP4rMVSwqbwoH6YtX0DLmkozC2CiWe3E8aCZDndm
tCfPWiZtXLdkgr1WfYmVuuv/eVHANPZAUXabRQYE0UZiiBEpcqPfgZukZ13Y9IGR
MfoswHRFAwG/ZYkLHamolTEw0wZbFXhMeHvaKvBtTiVEF2aPembJQEimvNtBkWcN
yqo1DCVREdEhrEwewK7InezrtcxooaeuCz2IoxAYpTFunx3sWu7rWao7DrEj65f4
CWZKVp1gWbJZ3XKXWhT8vB0X5jVvBiD7/oUXMA2dz7/WxrKjyNU1MJNag/DByKqB
HtVMqXry/bUVY9cKQMXF27RDIJA4vHAgIqDqRZ6szidDdPkjK/f5Wgv8J4CGvFip
/HZKS9/tZQJxLlNUm2SPT5jHx9z9ssafHxHfwVOHcue49oLWPa210Ot7WtItE5tC
3hmBvdGJhrY3I4eph3c08/mlKP4ozukp3F5BvOh3kzOCQqxObvrjuq7JBI8/gslt
BzZA1mD89FJ9S4PL1WgibhskezLJGr6rcO9N89wXk18ZbA+SKyW3SM5RicKoeBw2
pqwCtzENTZxPdX1vgAWpSEna3//c8cSNQohqxFmTR2SZiOLYwLmKLxIUrdi5+PAQ
KLX3Z+iAVHngRDXqGlA9p0OiU6WT2mH+7VKcs1urQtfYEDfcXOnrc2P2X8zSfU14
Pte8/SX++KsnoZRnYJUoX+m35jM4sveMmCQjYRgOpmSmXmcfU/9s/7jEXKs35X1i
VzWPv9JaMlwVKj0oLScx7zvsxfvdO+l3COoEVqQLSAGaeVoXMrskwsa1ItsVdJXP
PZ+asetTYd/5j2tavpM+Erv/9kHZ6VoU/SV1R3zmIHHg+gJBVCqjIdE3SqVhQhzz
gUQtDDjQmOkh7TWtb7CmBHHAQVxn3uMyMZ8QJkPRvF76D1ebXo1B83NI7x0wuHvu
emGGDDKfAAJzgdmVAQ1X4VeLvDsyB7dek0ty44JyRO72KpcYqIgt/GGLi6UsDRqA
/eNPdtZPqqdDwi9gjpBVs0sStZFw7UeiaiB1mRP8V2fcZP1d81eNiUOmC45QxsO3
29oMVJpnl+z5ZXfGKMH747kPiR62A0hT/CvtPikXuHNucQwA2nVSdWibTufA/aaz
H8qxZX6NmmZWYsCkwIKP6BuFYTZsXky0/5YWmGquW+VQA6Pjv4mp6hclrqVxt67o
DLSe6zfxFT84GsrlAhPC8PLLLSSeATnfz4KbIlHQfylWsgRB3H0pe/qE5ytkqEuA
zr/XbT3Xkr+Z0SPS6Vk5bib2zD9blxkfphDgq5Hi5eKMskI/IkXaaAP5/uckZjyK
Pkhd6eSJspFj2RO5Tfn86y8+NuhR5xR9HEB1pm63dKQrdo0t1stmSkd5eeBHdo3z
LF3St67tajAiEcbwjMef7Sze0zv6PPJMd++9JBJlqARr/9xlBnqeBykyH46pDaLm
5Owto62ZMvCAHpKW2qXbErKe8nXizmOvVlFH/Irpmnbc9ELTqSB/fDBd3p4IGXJE
6sbzGkJXtw/f0sRAo6vboy+3gW4dZxsJuMZ8TZb/cTaYfa5TAlYnDSm+fb4XyUmc
fFDkB+zN39kIx/tFE0P2W65mfUGbiQC6w48BNxfsHTw=
`protect END_PROTECTED
