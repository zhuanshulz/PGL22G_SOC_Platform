`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tiIdiSro4LNjPlmpoLweyo8M8j2vAUboharcJQ7g13wc8VYnoh75zKWoss4+69WV
HuldBZ6DMgbYdLzD8Urw/e679Zd0awtUzZcyO8Bap2aLzvSdQ8GxEns1luSPCmd9
eVqm7uNoZDPr6nvKevrgcznLgpxrplUkow/az2G/e4fFDEsJIazCFqRxsJnyFUhW
YzoFVts0yfa3/ir5D73A0tf0AMY1Pavk6U493mxD+Tg2ZBCauIaPGKJdgU7aHi4u
9lajYhZlkEpgm7EY/e9OjROBSAQDguZ19W4brb9pTHI+OznIHc39FWXU5O7Z5e75
fjUPI/cO8njFX4OOavMkNgEKk8ngdjAvdfK5LrEfsDRw3SNvZPS2INjWvje34DiN
QNEI3lhrtR+MaHBsnw4l5afMyd7BrHBkZXd1PY5FMZD4A3iiF2fIRjp5hSChjMKw
BZ/Gz3JcFB5iBIyinOMkXMU5YbwSKYWsMFM8dF9KzvVNxBdtMBcIt+AbTVQNIw2/
PupcRlWAlffrEDtZH6auoU7MlkXJKI27UYD95Jk6C88YlfCLdZhblVkARFWg/lzi
EMMYxx4Dw/QR85XuP0Kpc1xVUJR2TxSXbxgthNzakKCxruspJ0qzKqgNZSUj8IIO
/3K1SVkJx2ChqM/bocrctD5ydpgl7HSGSA/2DxLCnuyHU98o/BZzpIvHYGe41pDe
tpiDyaVm5dXbmjdXumyCOwA2n83dNKsmUIYNsb0WLByoU8PA6ZXrhazg2RsT5jT6
g+koy3fbF2QB1V9dmra5Rn6vnHFQ0z1Y9arWSsX+3K/uop68fwsvdyy2L08w5G9Y
6T8f+4dNTXBULUnNFSu3cXIsam3IjRbxPxxZqTpVpDgQh6Bprvo8fwrHvaNrm1TI
hZMvZIc6h1yPxMF1DlaZHU6oOlLrN71aOPn7zKjYLJHkz8E3OZ7BNLlu3qKHBJny
8MIj8ndw6XKDKJbp20onZO9huh5IUqvSCz+ZIMTjn2pWDgBuWP7qoFsOxuFLbb/h
oaBx/r3TtRKCmiKE/1T4BJV33f1IyCTSrj3FrAWCdwEskdc/J4pYa4jJY3OO2TJY
NDbvCpjyqO9FFxsyvOL7YustsJlPbXXe65gLQXTZPR7trUkDMzpitOjxiISRgfez
oFDGBIlw/ifqA3Bwl1cbsa56XmswBnMj7dew2CTESQYzhcEClks4kgIy0QBu4Mfh
+LB5zyVkJiWC9NrD9z2y/20F/pcHRnPcGOsaQczZVHDGhyfRwt4nYs106jaO7R1p
mJT9AX5Xq5Jki3i2Kph6IyyFxq5bFk+Mwu08zCPV+ReeLymikYwKqfY2ILw8O8H3
2KHw/YdI/U+hi2D3xwL78jzKmqTnaB/6iMJSNr4Rtgc7ozVJeKJqXXXWa9xazwUB
jeCgXPL4JQ5h5H+M2ua6zojUxYk8LulGMEnveTlaFeJt0h8D2vRW3QaLaFhreyq1
RBG/Pht2u4TI69bXsjmgaiOYDrT0qCHPOPBdrL+oMs+DQC4eqaHGGcVgSVXAqsKU
WzOn5ZeVD5BFLnM3FT7d9ZFW97S7Qp+YGdqgoplj/v8cjMp3S3peMSh0Y2nRhKM/
wdGovidzdU045gY4UnT/XMP35SO4WDKw8G2MZL0grudTEZBcSF6RYQJDXME6sYk7
a3bsYXmI1WjRPZQW+2vKilpb1LkUNpGMlFm/Tu6SnQfPaLYXGWHBBJGFy9NgbYRx
uh+DdpXE/0n5TdPuywfHbj0Qn2FUeh8HzdCSTtONFqKvuu+ii1v2MdRJdsW3K36f
cMckIzF4RbMM+sbK++bV/N2QMtrkpuwD7rhnAiyZYn3pRS09EHzv4JxjiaUeP+4o
twYRRJITqrGaorMbNVcIf3DkWamTIia8HBrmePhNVZCZ5e9dtZFbwqZPn2ZfxCo4
LCorHqBJ7np7g3w0WgcPLGSE1V8ovWCZIJS9ipDw/PwIBK7HLihcnf/oEraYDwUb
CJTmi+9Eja8wODwitHNpokegyPJBmJBLM+E/LxigNMpqq+FHGc60BB1b8FeoUiK6
RCUfpJSR8gHtApB3tXg1HcscPLnv7kwmwy74KbRdluCnM83z6EXDrd/OxCSAz8P7
PeNpU6U5aThAcZYl8yFY61tiAwl95ESQ6SeykiJuS1DwGK/w+ZsfhKx/xENM+K/Z
y0jxWpLNWCJ3NYxY7r1EGwAt2IxYKbpGwoIVcPDm/KPfOzuDhhhU3X2dUPUTYwOs
6/FwVMbQM7g//4bMVX6Xs2tz4rtOk0dNe5BCEZwcplRY/QRCGg688MU4XhuS1MaS
yQmdqIks6ogV1/X8hETzrZhOjiuLowfLeNDoKIU2TSvgTrvRYdSDna92XBNAGxHd
4frz619yggo9o7PCKYv0mEpBbg+uhaEdaFyHeRyicZz9tKsB68BKv6JJrCdFqZRK
wLDVgzVbtjEl/xKs31dbjym07Nt5dp7v4E+g2Uc+U+3LPCBtURfp08Ke9w1SqFtE
rhGffj/GkXXaqs33SWXDQgKmZ8ktqg5GdrzhzMdhcRxLAnKXTAGXKGV+z6XPp8lq
OrcdTqFlWI2dGTKsA2a0wDEl1HVnOb7dMAc27NhZJm9JRTCBIvn8edCrFGYcp2cn
89PhLWZ/rcc9wRCbxTUDsTaNcB7hrbQKOkjbrR4JjbIZbf0XAeVsSe82e8/MjRfJ
P6XD6JCkl9r8zDsVGG76hHmIJyAJKi5CZXQdupR8EJX9NtY0hll47zwsaqxdrmwA
EBT/4gV5Lxug5OCP7uzcATBHZoWu88KT5c7zYeSDWKqvkhbeGT3KS7p6sXoZsrEu
6TjV2FAUUz7xpbE8iwXDYAlU0Z+Fer/vUJmFsmnrMHP49Jbsoq2Icmaelsqy8rOp
KxArJPRfbl1BGD0Qb1Y0UWqxG94DS24P9+wCA2fBc95YlmhFBts8Wbgnhynzbb5k
bY9BSQkaSIzi9ncV/408RmbM1stQtx42vo42E2krYaiuaOlHUw4KFOZr6sdNzPJw
MGtlXepDkDUhpNFBpQcWfEC5mWVag3mj57TtuqIv47M1N0knDIosayOhrrozkWLQ
YWvnHR6qh0M2rzjv/m3VY1kUfJWfiAz6wzqqUFkquRQ/lG8ziUsJ4tWyFJWEMQ3V
fIrl/SThw9qFvANAHt+TXa6YSuyDdrVY4tAjgNWIZR8CaOnRWAPSPJ6ohz12tJl3
x1qm6TeQV/zlkP5hVzId8jtKtjzxOUw0nsR/klr6F9vBnLibvrls29pNyh87ex69
Uc2h13inuGTGtn4OcKT3HhZJoLKV/m0ylIx+CrwxDNuHbXskFFKQpoSNUwKd5Tkh
H+jCUZFGZFHebj6tN02cUk9PCqxWB79lBoDvEHi/GTzeFqQCChkw/Zr6RXYW+5/X
1PRbX1NLFrzrNXUhfyw1PdcCuEGJNTLPRw59G0iEMHDHbrYI66qfMk2OfyRTGgyn
2iVyg3Rx4Y0rzRAiuadSxct7jIsgmEUgTwwmwiDF4nk70NQMAl4SHzpCo47EbZCY
QCGHMVj6tApiDEUbpvzkSLYScdRr5RqPciQnDE0Qtms=
`protect END_PROTECTED
