`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+tn+C6iHsFFnd6/rFfsKch+Siph8KpA1ZHpsB8g8LyombXQLpjNTH22fxSKz2yWh
5rsxHdGQPS3NswcQyq5H6wbFDZsLDaS5vcevHNBMLdm8DuLjGIr548uo6I/ijcl/
cYQaTt4WjnhsoQKDKrUaUIuLU2Wsz1s4ZYilLuIyBIzvvT3cb+bA6S1IzTLiktUF
xt5l38GzmUw6zvClm1yy+MV6MvJOgJTkm7Fphhw2apN/anTMMqcp55E1npP2T+z0
5/UZlOWNYoEDzcpFMwrSkA==
`protect END_PROTECTED
