`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rpQHlwy3WYXLhP8gaD35rjJ/TG6RiK5yLY++vznGrPRzIBMdbwYDu3TjphhdNMxk
rOsIXkFyFHiT3OaCQaEpBSq0McnsupD5w+wE9uCi+jNr4vCYHAWKwom7ZZ8b6ehL
stQjThI0W7Xe6OefqgH+3ha3tRQQc8mYIPXzVpRi+VuOylVv5AuY6GUPOCgSHMgo
TBiD8M5EhaFYvQNpY3EaTfE+BrjUpAN3J3uyYq9os0P7vFQOFn7GqWwRx2VP7v1l
`protect END_PROTECTED
