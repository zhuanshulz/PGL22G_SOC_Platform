`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I7I/N0nzaKj2Yt4J2jtXg2j2whDiQoFw5bDXOC5wsFWxjgg1D61YlD385lcuI/Me
vwwwWYsxIb//+DzyqVlAItW5TXkhfLa/4Dr32PLjl3ExOwJA2vzE6zISZ8jiVygz
krLZDmW369kvq8ViwgRW+tEz3SiMS4QVoorOGaCxkSdvhNtP6S2WGaaL4E25rmIO
dIzXZi+HlJscITyFtSEZIibnsk5geG/y/iRGPH9i32y+KdR/vxE7VUoeCD+xGSR3
c5BMDAwkOnUh53zcwmz8dPkxoVM+IxYH1b6ockjILDUkNQl0G9iWrsvJolSV4NH/
qqOYbu18xsooGOfa6kW/bnE8MCAxZxyWQEieHTO2Vh3GGXbvop7sNict8QiHnBlx
MXadVsomkVHdzBO52brj7C7leppy8ePEr8dNyGE0ESkDtHmnw30vmspT04MDsQQR
fmG6dyznyuyVWf9bNceZCUX1F+T/K1Vm0sf8TbowBRKjotd2/F7gDWzfEj2vuAvK
LkImSyJo+gNACwQ1DkNC6/IT0lcJNkEMS7+cooTSPTsYw1Q5FRzUc+6E5TEQk7Oe
I4kZFnILuJhzumNU9+tu+HAHD/3fuAyJa27fraR1jQhyhfA8ONxCMjEdpTKuB0FN
2FV3Jh96/xAzAuDAi57dDK0K04YLASRCGnXZs9lpU70=
`protect END_PROTECTED
