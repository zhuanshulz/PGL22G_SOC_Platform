`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yieX5mHMuENBSmnzWgu75nMkRppuMn+hIx6TqUIniXThUNu1+S5eAaes8jEYt7m
gdeQEgqrIiU5FRV5AR7j+5PdjidOHYiM/GZ206ynh+RwyTiJz2dkMlbJHqsEbYJ0
ze/NNKaCRIgDclLtOBC4oYbkxgC0jevPS+r6oH0xH+bDKyws0pVK6u1xRATh7wOj
su4bYD2xtf+cRfG6soqO99EiXYEL03RJrFTEXXcBfdA5Eu1iLJK8FzIgzNA96S/D
l0WsnK7oHao4g/Ym9/Z43RARaGBzhZmlaBV63hxn2kAUN4ZK50+VMDPbK5/gDC6v
q4OkeJ9Vpy1UH9dog/M9quX0HTgXxfK/Q8vNwWrT2y89KzATxrRc3CeB+SjIn5+r
KbTJHjqj1SZ6Rdx29G1WhLZtLPNM7wmz4i4AYAd6ZMkRrx9ON4DMRUmIsVW/JNAz
Op0jj+fq/m+JFDQJrlKYQ5VfPf7TjarG5nuCQp0r3r2Uf4gGS0D5Psgy3Jx6C/gD
vlExaaV8byXRz0vvhZVlwPDp+VOuoK4q6JMN0cH1PQdKGEAqHRIVPdgbrsFm2DAA
D6IcpWca39SER0aWz1H1Kff1kKBwp/6MRM8TgMWu05IMRxpVJtYE0OREZ8M1MPlF
7GEFvpzdfcqG2loyYq9xHf1q3gzHB/rQCUdfpwy2w4Bvs9v4q4tkXqVfM2eYaddP
4GXz0AcF4D3hPz1yB+NwTa8eaM9KmYw2sTSwQUZp2ZQ8acj59zAaYkJgNZPnBSWG
c3X4rvOSY+qBaZQRE9PrAlNNzLKhj1fv/TbnsR1FlTNnP4GO5N4eyze3yhLNoSJq
elemFLqsy1SiW4279NPmQ1vU96FNmUd2avYNrszhP2C1uNTDDoaS80Uu+dkvG4gX
AxwBWXUOGyc5IqEyhunNKMmakd77Xm6gcCSDeZefnhyI5hbEXyBoJX6w6g7SMQTl
WdjBIoiamapVwkPZWez7S7Jk8oblFRhhZbsUJO+9noxWYJKy8WSr9gqFONikAWxC
4AQ4YUijQH7T6MO05jRnSgEXaajg6Aw8NXuf1z7pm6XyUZGk7+MlUjIbiJb8+/GA
K/CM8AfYgW9lgw7VFg9PcOdFZJNF1xAJNF2CmdwZR+bwqirGmrSjruX2Vax577oW
bRymFMJbjhZc/Rdt5/HsnNh9fqpwst65zaBUZIy6D+wcdAR81QXwY0moDdtQeMDs
sQhgScKIeu0wH9p4YqULP/bL9q8Ryb5MQ6lGlZwZUnASTFfnv8WB+Ehm/1pfhojx
X32bSXw3z+pgd5LDx7zVl4jEGVsXNWtNtST+hXqWbJ3/ev8dJlnaWFVEgztG+Wr7
kRQicbNpQzO5aEnQmJm5FpygmmCXDpyfhLine7KuqpvKNEkN/f6xEM61DAZYsnAN
ScgGOWQFhG9JjPqAY4oqzxniu2fAto8siFb433zImCk1L5q+qafDDtGygQmbf1ya
tMBVEiaXze7gfJfnwAAKwuekXTOQz0rmo+st15dC98oxnT9l3jxvbYsy4LpZKO8S
Ln0WvwHKcdrRDkY9j3b8qk4i8mTRiuLzsw216h2NE7r/2+ZLx1DtUQfDL1Cf38KX
E4Nqmk/QIQDC/Fc+USjMtlVA4JX79cbMpWqMFfunpd7qbQwKdAJrAe7Rc48dieA9
s9iHphIRQyLSousNZ3AtlWZDOy7oTXTsqJBRbTld191aLCTc8F7NJJl9hHBkDJna
TQYjmKXWBb2vOw9LrEdZJ+wjXF2sPDU0yV1LLIhf3TCQ24US8tpLBRlyNgYU9t8G
x+rBxn4Qf984MbD+DArwDJ+/SqHDclzPQ6sIUARiqMMVQXjSVjoxjbm1Q1Xu6eVK
rhh50eq6WLB3PamIxUi95xHF58f39IWRXxVWvhJTXoowMm9zUQgZzvmhw4CMtzey
0Azo1n2bqiHOAIic9ubFh0nS2xV9fWOO9Jh1xFtimqflOKq195x/Hgv0sGfyBpOa
HhPVQ+1TaFpAtnOkLgWTPA2ST7VLP0l9wgH2Kt/Q8ZcPDVSBdapl1PIBVsNNALE7
x3l56XePhgg5AyQ9BzRwcvSQwPS+WxH6QJSCcoNaCZuvHbNz9l292WpNUbIVGCRi
i89sGvJLlLrFOJyGQP8RKmR10CWDnAUkaqK/2DegD6y547wmVr8pMSNYv7Xf7Uwy
HqsmzySppqSzSEI0TcD6xW6JEoQ/alvy8TkrUlMhhGd3c6bLom7UIf3qToYld0t0
TGGvz1LadtmvkAgb9whTb4GnoYvlUzzVcQQVHziNSg5xeh0PDTBCWDdKwUz5Kjvp
ov38kSqowqUDQnb8Rb7BV1RSzn+E8tiU3UOWmqMZwfx9iJSvpNCGzM3Ilms4veKJ
bRR8kP286paU1YZ23VMjIDwosK9mRzKfCjOtO4v9bLqQqrKpkU/uJ64E6+XGwguv
bKbX0dIv2eBlQzY1q3XQkCyV+x4LrEoZu8PlEt0oLUmWBxhDUF5dnSBDz9U38JNW
2fyVMZuGZ1UjcQqmhxTbIrrxC3wMA7FKIM8VXPtiAmup1WVhIxuKFg4A/NFCxjiE
wnErD81IHfrtos49EUbVrwJmQlgKTAWS7QKgjMjXkUBrmZpU0KtI+/ioZNl7VPI+
+1MyaQqwaToWxEy1Wn/quGtpFLLGw0/4wPLt4MRRqoIfAWypb4Xcb1r9D3ZcPQwY
y1/Qu3TtA9sJZyEvgoyoGjo2sD+J2at3kHUAkubWCI92hEzceauZzIT5fnCbq7tH
ZnbFantYLfqM8qBVyZlcH4pQ7Msfo3ARbv3ErJsQbeE=
`protect END_PROTECTED
