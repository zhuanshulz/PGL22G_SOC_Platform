`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvaS2Bw8KDqhEjeOt8R/yrv903YOJh4sxN+MdiSY3V7e61J7oWbZB60I1pxCW2Zp
2RLjRUqEXAvy/I67SNcdCQhPf4Frfh3QKKKk0UqlJwyZCCuGHP/jiLt8K0aDRrOv
USdzrTmcEa6s2CudLfT6e7C3B8gQpExMjYiQ5OZtiM5/mOI4+tMRQl5Kya48arRI
PBoBPqutTxIP2lPHmBEXS94e+9F/PSkC4VVX2zfoXBFlKzHbvkCfXeFNB19EyfEE
JJaQYal+MSZm+mxqlS55ol0Zxy+/3XveMKXoAQOzf/L1oO/H/F47IlN/4Se5KGXQ
Hw2VfsMWJMrdqJ0Gcy6UaVH083wFU1H5cfqKG5+hMcPK7w9KB8OuTjQRWrCdyNln
fSM7JcP1rTZeMsvcZEYYY6RPHXUXU5vilaJgPERLmqoEHK8cvGfzWrGj57X0wSNM
H2tODq5wk8qO3Npvl/bJywWNIVtyM7rsPMHPy6NJBW78fDD2DOlJaKy0rJNMmyJZ
DkIzXxhIGyYr0E84QheGYknOtt04/sF496bkkiYpO4AepkIp+9I4Ib6z9Meucv+c
q2yUsqaUaz7c90LqkBlXjSZkMh/5cS37nHBXb490KEc7AasFFVFqpb71S9469KS1
7/6aqAU9Iua89NMBVlx+OkmBoGH3QwCS3vki6oa4WgA9RJqUN1kjgKMuCx2a1tSS
y/mnH7jUkD/By72Aglpu0kJfS9kTQ18tJIk1kn2brcn8SW7am5iB+Gc//HHsontK
Lp2V7F+Q42JDxdR+lRSF4s6YDyEZMi++1qo9qpyT8XRADU9uGc1dZX/GkCr1ATt9
PUGeGYW+DDgZ6gkrl8Z4di+eFYuAiglHefN4IaaaOkGrsps5c2Kjfxiinh/1RG3X
H5AiqJHt77is2CAIkPqnAyEuGEAR0m1xPuapjY0BjgOD1dtIw738q3Q/d2aFhFdn
rDGwU7Qj5iDqpw2kJ5GA1BoR7FWY8VyJTpj+xFqTYTOZGO643LjOTMZDhdG97gEE
Sjuu6ZDpE8bWJcvFE5G2KZeKpqXhw3KHEKcysXzK4b8VKxPx96Bz67n/RPXXxSwn
wZTg1OpC2jYfVPoFlqITZFnc1zuV+LnTw/NHwtINpPMXdfZgwnCvtzd0kPMyjVH0
HXX49Vwri+fADCgGgP9SyZAtxI+likh6ja1KG6hlqJJ74Rm4cMAxnLl95oeKmFpJ
1aXdR000jw8wEHlPV0mxvoqIpu28YiZ/wIMZdge/Q0NJ+4iK/CJtjkjVujpyf5sd
DoAn1ZbPoC/qkoV186C7NpWO/j20robPhGgNTZcStOuWN9yiLbi7ANxVwSsi6yMa
Su9l51BFMZOTtbQ6z2yeVDds68jdyvLcXYXThheGh3nEWXeYNyzIoV1W0ZbtU35u
BSL22wfU2aEqnDylSi2I5Wccx6EbVuwuUumeGvsLWYOTTE7SkHMrwTP/NmZspwRp
588YKeVe8PV9vGPoKebICb6abVWn/HFQ9o0UiYtvw+CzimchnNLno16XiBmJhkg+
lsg00Qrpw706aedhTypnn9lk60dgsjtNu4CFWmAIeGtLj9knt0SvL3HUjM5Qq7IG
uAhLpwtVP7FX/olMbynm391vOdTlRGW4hQh+gEgOTgye3SmEoEs89v/zn2J7v0V2
IyHlAYQApe4KV9e1mk2Gio+UdskB2j1V+XFKiZ2Avz7AtzCTJzOZB9QKEomdfmk5
M5aJ9hhfKlBK5e+6Tx0i5ErzK683rInpiaaWSBBhFn2AjRLJg/OM0dJuSxcd4429
B+825W8ZwXh8mWOu1VRrrLWt/MnZiPwVRf7lbQrqMSC4rb10AQioPLPe5E8kNcul
adG3CsEw0LFbyEzYR1Oj1loyZP9YFA1K1ZxZIUw/vl0mLo3L6oGlUtN74GZ1eLmp
Ejhj/bei2CKTA9sAp0Ch/0C/X5zX9AdRmJuBB++Gje664C2TzGkarAdMrYZ17ez2
T/zmpsJfB+9wFL0Esh13KDXEvSVlqFqw81HPagIydpDTBbGwO9D7NWAuHt4Co8/V
M9+vLgotmBeeEwI9HCjtgLRroUyBYQ2LmkTr+vgj5AQJ5FmzQ8qGDcnfqfPIJTEx
o7DCLf7emYaGPkL4kCPtuQmOdPZiRgM9eV8j4eCRy5YGU1CrNqipdn4c0X8EfLhQ
nbwd3ePa4jepUCTeWeSpXSPXUPy3/nk+dlJdNEhH3BETuf0Odz3cLQjKT1ZFsKeN
FS07qJyY2jqYMWDi+CNu1yAJXH7KCmEResb5+Jz+Wd5orqBDjQrG6yw5x+/WUjiL
3G7VE8rdPy58TmKT1g4uH3fiYq7YUdfqB2Us9bWgYlztDhN9KCXyoJVzJZUuVnIA
lO9PG6GXhBxwi2io35/a8m6cWA+KDa9HjvcNjEKKtIFlgVDgTGUrKF76YA09OJwd
e/5MjWGxjr0IqoEvgz3rjkqWayNzRhYI1FLTsu40mnzOtEvkc3/OV0p4PbnS+V5x
uo/m0XQM4d73FZX1MVamknh6ywgnTctQ/+tPa3Tz373k3WW5G0/sDGNxT01yo7VJ
rd7n+bPSSAzJVWJQGhwZ3tb2Sv9Z3N9usVHZqbJ36uD7dEBRuDr+4VExd0ZrTaab
yURVAJmIwhBVXaBuKbLs2RzY/4gylxvUciYaXbnoJChP/4EV2QaBMB4NwDbk6XCx
kLy1IEe7DT7/Dw2l7AbYvFiohgbIWhPKXLwCg6TXPK8P6ukTxhZOaL0mvglMTioq
UP136GWU/rVOY/DGcDNtDQ==
`protect END_PROTECTED
