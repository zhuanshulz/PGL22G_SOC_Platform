`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcuCKLRBgy3+W/GfnrryGCe01oHM93nYfhKLJ8OAQUlkMhNLH9HFPsqJsoeW3iy0
w6i+GN4+ju9SHkmArdgB2qYF6cZDHNSV06WJyLeMyj1DHDDcu3KnheE25kcCfel5
ysLmOFHgiVDHGG0/PSqrer8Z7Fo7jWpMmrZf365FngCrO5hSYOnV3S0TdLZeP/CS
PoJe+4psSFAJAtW1B56GzP1Zyacjz7txERSRo2FyfIKNstFsESWbIrv0fbT9H7w6
JzUhZ3HGwR4TxgX0KVkdUp30vC3SVOwd0RqBq5Zeog66n4OqdP7tndqcX8R9mXJe
9CZS7Juu+oy+tVXUWmOC8SyDyM0tVNbHbGjd33fwQ6xmYxXlnPij2sLA/GePDezE
w7AjiKOL0FM2jBs58JNH00prQc7839l6JpwExd4wWe1kqkoU9SXrMFimt2fHzkA1
IILYDh7TTPDImHuDThq7WN1Pa3os7Pa1H9y8PC3cIyQq6N7HPcQ0sSMngyCa1Dyz
tEQYKy9pmzoDA4PZZRokMXeRDYL1nSIK03p2DIc/FsF3t0dreo4I2qfqenEK3CO1
G1zt5XcoxhdBFiwN9OONw/QNGM2/Keb9oSuoz/QTmdKveph1Ker9Ia/mdiBmgzsA
Q/HK9+nPy+l223NBdXLGdJEqRq6+JGc6dT9qlCMQvKE0vjhsl0cpaKP1l2z55wlt
v1sWKdJ/RMn4J0w4tDq9VuEUiUaG9ASpW7FzWL4IdSpUkiIbkMo+vaddangSG6B9
SQ+KJOmF5EHzbNqjnJzF6UDMHsHRB8wyGbgVL0rMUAgSG+1zqy/nsImFNlWO8o0p
xOAuAEbPm8l1crAmOckNp8bkcGlJwhonMY8AiQJFpa/eEl/PXXU/wjI/FJoWE33a
+stvfHaaNl5SJgiIE+cIQEUzcsFGbtYp/qe8V46mVVRUzziqtzK7R/Y4PiYZRNU3
nn3gBi8feNqYx9fOVwHVdSdaowUS/rCqO6z4Ng+lfdB5cDMGzwX3Bq6tzBKvP6Sp
AxvsLZv9sQkIh9kcm7a/jb84ATAqB5IeP+9XKn1uatRqdOVTiLs1CJSR05T+HLQ7
XLxNU25WtjohPh0zF0Rb+iDvX0ZJ4ZNq7jH0IGk1AfEyXmPGP0Uo3vjiOuufJiuS
croMsJ0H/akJKvBaNfOZAdoQci6kVftGrkpsbhnsb9xtZybYuaXJNR1ubD8lsTqD
ymc2rWtXE3n943OfULCM0S0kRlXfhTl1d60XjZdxjys8TV3kUgaJ7EDdhtsB7RUn
BF0DU0r7HOdlfBTHnh/Qp9LO60fTwTMSKmtApCyTWflT3zEdRF3S2UexBAvHuzS6
W1Ygc/fdKhmxocT2MLca109v64gqrry5UVA/gQRL9p2RcuzpFzUVQeLeavGsoSft
jSQB9No/0llmSsGY2hWOWz/TBBYWpW02yl/vOwStKHt0v6IyLbeFzmwWE64IJKDL
YwLlp0NsThNsQeYAE9j4b7fo/D4I9tHzGjM1nnYA1/Yxf4mPI5dh5jP5qP+8HpVz
jKG8gFYaN4y55o7YoEATwFRYeLkhRfnC0+eRzXlVSvps0bMiv/8Rg+5dYO0jFIgP
aMap7AUSGNcjbVQ6nSzrbIuQ8Xf6kE9pctRCNqGj3sImhELNp/el+8eG9mouOrp+
W1FHYNCcpBLykSysb4+T/x8JzMdCf0NPubizB3mv/OFz7L3yi0L0/gCDfna4orfv
zkXzv+vc8CeGfbJ7lFri4CqSYzLnVL5kEIR4onpp5qssMbQHM9SI/9G6uiDOqFTe
H2rLuiO+Lh160MGpyc+eyCSpkogQ03Ovfyd+eXL+qTaH7jHZfhoKFzH98O+03nnA
Z9yxOxJ/yS/vaePKpcOfu/9tHHdJa3cZ4RdE+6dl1ocgIw2IlCjrKorWFT95ZD1w
hkeMwjRd67l/Rqx5yjqfHLVyOc/QKvtXVoNUUZPGK6qmrAVYYFoPODV3x7Rh4uel
RzzqeomCu4AkJf9YFXCm+LgtmISoUD68L1cpaDa5dWdCKYLYpGAK4GjPodxdq1gL
coKmfdwxJrZKqXU4ni1vpmmvcv/oPBgzEM86T9X5kr8bLxlAWcOYSqxPj86ggBZE
yM/MejUjTAQuhTxV1oizOtUHDYCP2i0AWtcftf02OXpPvOmbm6cdav9s5JTOMIGR
7w7HmqHKI7SDrrWmzEambfypJDGEKzkt6y/dpD1qSBJvGiR4v2Tm0iqvtBoiBGOM
tinqFvCqPCs+x3ycrYqZooaVgt61PEBdqh0MNhj/azShZFwuHONNcyWL+St6QGz9
Y6VI00c93HXJSXiLJ5JnBauYi1RuEd4kLaLV/F2aC0Hvrdk/DONM+WIO9H5V9Htm
c5ylw79bHpmYZUm/CCcJOoG7FPTFnpPFOSBjqWB7nDGdPjZteabYk160inqul1Dv
QWMwadNfb2ehGzqa3Jb07/jYV98t9nnr+MvHCs/UilBzlfD2Y/nw9TJ/p+5UApBP
X1emWCn9Wqt0whPzNAw01/TWAWGA5DUcFOJNq6gqG0DWoMY9GRGj7RwQ4j41nlom
AbSUc9QYEHqaRDGUpftCykVMXmYnCI4bzMHuL05tyylb6PsE6VKO1yZ5TLAsnM4V
t8PyjkZb9yPQSnMN4NAz+2HT/M32Nb7zujbh9KEKLDWgmulsNbIe4FqTM8qva1u0
ZyXygKNPYiH8FArGXsnfKqbg06Rw5JS6DFdWRLMmoMgJy6OYTQkdhMWAmt2oIEGH
SiD2hxNvjA3mgI1nuKU9VdT1ni+I3f1Ow+V7Bam1zWRANolDXzmgS5Q9/KruCwvO
SFHDin91b2vq7zLi8XOch3sgx8upfylIqJtDU+vv7GRHckuRbrIQtxtkUF1EzHmH
MGKVGDggWFnqYWFVE6p6jajMkCi70IxScmTKYiUBt9GLk+dmFs35EDVtbQUz5xxY
+jcctTFsC3AUVqOmZ2kMKgyXjMnCNm8kcEYtq62c9PAWJpLE3bbjtLG5HIriY6lT
dRLP3Og6iU7UcdoLRj9byVJDMGb3uIu8DjZXNclWsbKK32zYBI/3WxFckqXlK7Bc
xwXKz4M+FNgLt/m5FBXYGGBsArkNjBQrZIffpUJQA9j3LI2fv0nF7HM+VrDn1MPp
91NXnRRQZ8Zs7AVNrZH6yazlnGt/+I0nU4Wf7GbuHPnf5CEeweEjLe4cPYCUEjeX
PcRqR7fD56CzT4XdaaKyhV2eTnKIub1UKB9O8y4dpJ6xtgNym5g7FmoeFtM9JVTU
hAOQUuFCImxLqUZQb6K7pOc61+iTAMDpoAYyxXaBSQtqY3xpa3/trrHoHhU9A2eu
x+FgwocchTWZTsb2pyCEhRHPmaupPnVeNhFmjHork4+YyHWosc3UjzEBqJe1fZbm
IRxhID9Fh/YcDP9B2sgt1OIDBiZAjhrWeMtLqLvWvuvqO51XSqdS+wnBBH5bdVDW
hmud/mmBEpbLOZUTwXMRPs4jMZIq5R5OcJSxRxWdWUodihMKTiG0Rt8aAesXddRl
rngCreOH5AwQwGbz7kbRvbVf3Gb/AwANDtScq4K+odO8lIiDsSQNLpixiG2l81VL
2Czbe6Wjk5UpLI1Ui5SKtTGiNDT08jtsxcGTKWcdoi9vCu+dnQq+NexZHg8jXgdw
etHIoiDfSuL797GtRhrCAHXnzoOe45Rg+wStUTwVcw0nMMRFw0MlvSobFqjVK9lm
jJM/jW8NfFhbpYKTDKtlhMlkuRAEeV11Splu7AaoCFo6Lwfdkr6dqT50MVmSPgxL
P/g6k2RQJIDu2zJMMAcp4ITh5VQ93zTPher/+8NcXw5X4MN0Sxc+dwwSj+1FBKLv
/QNdURH1s3RPaOADvjDLgGdeT4hzbOinUXCbcCrtygg6NvVzFx3ggl2gXHqDltzK
A1brNfFHcjNaom/wD9Fwr79+Rs9hIgr2RGdtYV9vXD4gHbekUBKxj0EMywmhX4JB
h99atHqcshZ1vI+2urRBPXDEyVcaFFgige9Sye8waamixEUz1r3rlEG9Jm79GGAH
0TM2P7Daups5SvDveJ0FEcVsyd/9UBRHrGLj07mO6hybupWtiOsep1XFSm3Kc/Ca
Hx4KOEDAxQi2OmiKmrPQ8lLWg/owwBhwl9HKaHi7ES8/UO4UKs7wfBpK+nql7fcK
ONLbiqb/WHya1mW7d7kS3efY6+5HBwBbiWxYk50+BPwTxFy5KNO8qXdlR9nY/bWY
IMhjPFcBfRuSX80ZdRqZB8Kkz2zAAIPlQ9Hjz4Avq0mfvRgLTUjR+/0XhmIBZ6CY
IMFAwPBcGru5RQmMnPpmjye0lI8POyQ9iwwWwJVeYC53l52NvAETx848beYbQXHO
0DSRC+9GP0tKDchdNNHA0D+TKo0MUxQ6GER5GXs8LRRzxirvBzBEO2rcnz4KjZAw
`protect END_PROTECTED
