`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M26lV+dw7GoiuzZGT43FAq1bhazzHywUXeZkgxQjse/IXx0ftKMtsDWvCN9S/s/s
i/k7koNgP31Q3NCgYV2thh+fvj1n/O3Ylh8STDKgI/h1wyJ83f1J+WnNl+S7EhCh
LpuG8VBdW0JPW3ojNM0F2bpeThEoJKQLcqGlgPQylPVQhX97vFQygpNlaMpkluVR
v4Yd3/Ez0e8s0jdxkSQhSECJcw97pAZpmke5I2VW/Wv+sddUhDVRRxAyNQmqbK3a
sPl4xhGVy5CsKwLQP5STzHXnyK6yTNLgruDNJQxl7aURuy70+kpC45C4xS9mPjb4
nvYT8Jr4xiRhx4t8xw6cVt2c8G2gp3h4I3P2rj/XS38rns1hXEYJnUDe7r7pgSNw
9gKjujP1saVygD7pkmGheiZZElGOx300VwnmMiVieeCvZ/A7ggXdCWf7FHieZMfc
2c4+CaR7oDcTvvS/p9xeWCxl/cx2bNGAgtNzvJ4DQrX8KYEg79bAsQ9Ag9mVsz1M
NixyosQSZc4p8XPYLLyyYOdHDoz5sqtB7J+Fd23e+EP3ucdEGuyKeb2PPo64eh+R
3T+1vcqUyqqRBEsUonSlPljlw5e/CJuyDwzmzemRDpewqY5XBqI8PG2CSONOQVYl
5QJhxcAmTyRoQcyXQCDlG3q7RaSjhC6ZlWQIrvBgo52OVbbdIo8kCiz3zQ92+jml
iRJyZ9Fcv8DYg/+7CPO5OUR2KgbWvf0+mT7iDaAFhZqOuo2smdgSNjsebsv6salM
LLyXclJgFDm8MQxJ6H/68x9lrEOJU9PTXuJKn1pFlcKMsRq2euIzvzzx1Aux6L0g
pOj4WU4YqJz4QSNwPts/NFoCBasn8IMPZg1Pifdc3SPJE0wU+dQKvmqtqw3qtXm/
B5z8hFdNyfrexnC2xmLBqlLgpcFBibiGLF0BiFMGyaS16HFOO70tcPdcF66UYjFz
HtJPBSuuJcGBuY2f3Uvp+61reQT0VPFEodvsZoBtANAHFDmKFd/dmkEhRaD8za7b
v6SLmCqrl2QXENp5jvvy0xH/sc9xCilo/5sCepO1ni5HGa4VlbLXHO11U/Ue6zrF
ENgqUyWt8kN55KoU9Li/LUiWkH41c4wCGgTuP7y/8wJ4QYh69eW3L/yP7P86kWz0
ks4Fl8JLuJnDY5lFVx4IAubRkcnF1YEjLCCTwogOEXfzfkPrcR9m/rZFakcwiEDY
cFldusxnPZMSEaOOQO6LN0I181cBccbE3idrBBQP2D0hxEADH3Zp7OvGrMu6pHxR
EajerobOpeHecbbnOT2qHcgiKrn4cb3wwK/7Syv0nmJgQJb+eceRRwo77RNQu3Uo
FcZTeF7X3UiVcvRm4hbKhnmHHuDD8aBCh+EKc0rNRC6yfYx10zqGoP2avNRJLTCv
r+TQEITobEQPHcnrFIZPQnKOsmvWZQC271gjTOZumnMKcEV+34+8NkbQaJXzr5/z
4Twv44Dn2Y0TzV2E03ZkYHOpFuADtBecb6MKzDYp/5AiVoKIOHQ8FzHiFRe9fyLH
TqA2a/aEfMTsSPKZPuNuuRg5Tte+1/8Mgz4lYvazXvwL2QZXOcRZhZaha/Oo5niz
DDf/OkrDo8aLfzqZpBi+J+u9WIBHdKzrYQKsOMXPkKkFtmwqMxGN69XJ2nVR7wHC
e++bywBwhmi0S47NdPQ4QA==
`protect END_PROTECTED
