`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HK7UXb/ZNgbNa+urlfEVCFRTl0aOM240t2Wq8qM04crKQr7j3ab7JZ6QF/Jp4Or4
26YtSBY3aJm68mP/BGz+j9j8XMOGAnWTED/q9UK5ycbA3j0QFzCNqsnQ1s2rfhA5
Zz+JVvvPTLgmQa6Nkwhof4Y1rc6XBzbB2P8JQPyEMFiGwEKYOs+VbfMvxJz3EF/1
RP3du8K4pFm9jooEeo58EtfKb8X6zEWdD30NaOyNviabVuEFQAcoZOKSuA5j/omN
jV2Hyp18BFNiKauFylVETSBEYALIHw5k5iIUf9Wvp8UOFvkPH70IQX/pyts039Do
sVdzfHpCX0IbMZkgpzGzoVAg9nbRLXrsR6c6TR/j0z1HiOUhlvzPUyv8iSfmks5x
bdqmPOk2lmBuihLLsI1oOtUBioRvuyUpNNshtyL33bxRtlPuB8Wruc2MMa7dyf/9
un+99nPh0w31DYoPCrxZlcujVl7IJ3slcU7LVG4XZT41VdOSfyfzaYG5oCQ90dc2
JeFfeDv811O1eHeqXcb7XtQ9cL0GzlSskYswweFSyJOyBXDiKN5sHtZ7tU2k1xr7
QWQyq6RRvlemYrb5+Mcotw==
`protect END_PROTECTED
