`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CdbHWzYJkrlGWzNmZHcrGwXDLfLOlbxCONlFkxD0YmFWjTZRUvIBS3OlR3vPAQQl
LgeC1a9TCcaJpvKpE94ed405j6RhYK28MVNdpiYB8FLrR41K+gRKvlWYWrmbe7PH
RLS/e7AzW2fCwjbwCiS+x2zXQ85Vr1+ZDajsQYJBfKP3i/R8D1aCI69mPi+EJumg
bAUcXj7cNrXSh/3ToX73SpukmJSZbfP1VK1lPI7oA/jy+LmH07opXO5DgTHptXhy
uYMfYXb4T0ZYYKgFiArwIaxhu2pO/iHT18MdN+ybdRo1qbI0sv10zPXKprdBHcmN
AEm6WJkqRSWBK9I4zD11YYOUGQM44LI2UDpfHObhswwF8WDvD7skJzeAegOktZCT
b9DAZfqIU6wz1fWIBgFRiN/jKIGpuyLFMsSBfliU8SLkQIlWRU4mio8yN6dAbKmn
+/0SsbjoopJ4Qawd/z+3zWF4ZqtS8LgmXMkbmt3RJH1VTInFEv2VR9RvNsmupxLM
9dHbQ4o/kcXOYKa8v6+zf6onTbl+Wv2XUQTibLO3/CcA8lHyd6efgzAg0FQ++jIf
IY+f6K2ph0lYWKAhmL1Ez2FVItAyThYsZhk1zn1SC0htSJstqPQOzA0lrZ5dofA1
u4NisH5J/9yjhNN2bMn6+A==
`protect END_PROTECTED
