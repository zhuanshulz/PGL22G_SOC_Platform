`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qsc7+NNXbHFO/FdD7tgj6V2Fl0gi0ji/HmCaQCJMIHe7djMh/5LXrXwoDcZwmPhJ
IU0Bvm/yyIOgJzR7e+BKEkpG2xiWS44B2YbDE9FOMzeqIBkm4YSDg/eDRZ7F9SND
oRh8NRVBmC6D14kWCGZUoXpJedhqZ8gm8eMsFWO0Q5RnEX1SVnGZt+0HNRcZRTp/
ilJ74HCUSlxY5Se6+rRe9yJoCt8KpqLGiL7QrqSfDEe0bgKSYnINfN5nXW2ETgXG
LDrECz8qIMfdu8LTDe564/n4x6YyD7bz66Ep790u/z5/HaH6EKQdmRDnlgI+l/HV
VpoT1oA/io2ocRdAydAecACiYlNG7uVEC3VF1EI4lQ7AUqulh+UG5PiE38npYYQE
kEWmsvg3V6jD7bsvkYcQE4oBzkcPAyRhPefztGy6fgofNyYT1ppDmu2/yJDYUhDD
BsLqJ+fk7MervwQy6OnQASZbVYJcR1XcEoV7pkL/RMe4n8sbBhxa1a0HABKBbu90
zyfhSmF19tsPp1KA1H0KEwltFxRf7lcyDY2HhJTbkbq4KZN4kRL7dgV7ifjbeRfm
umUZpv5BP3XftZ+3/8G+9FyWbamFlxXva9PZUfytnmuDueBOxuWs/OQwlQ+ecGMo
oNtw+OcjiZ5P1B+rHrsyBAJ0sc7HI0OPuOr2C9Kyvwjevqetq6DXEvHuPK8sK4pE
urYt1hmfnIHjwPmAbrKPa8wD8qlogbcQUlYgn+rWqt2a/LgOYwnrogO7IRVp1AeO
G0iuNh9hdtJ6KGUmWVnVIhjyHMa/EOZXYVMlvl+QSstPWHs2lmwsD1skOZGrY50e
iOojlCt4LN+E7pVJtXlOcSsYAmQ/+5LS7A6mhVQl14SPLTXGOn3I+Kuxqm5D73on
3dl0oCnJpU/s2f+dAUSo6ZiiC+iYWmJpltNMVtp3S508PsG/F11/glDrnsuG5TgS
PfQRfS1AVy+XsQFgn19gPRz6EnODqZ/YqvbGVKC/QB4Hp202Ljr9nsJ4iOmXz9Bq
xjO3kCxJhx+ghCKrSrZJaTMGJZW3NkjzCj0oTiuAzryvDF1LIp7zehBVNxaeWrQq
/cRFfsNDn+xpjX4uK7XaThlhC6wV66PIgc+jyU+QyyJARzQyOTS4tErTyL+ihzBu
kVRhfnpf6xBwPZdRRqbkztJ78wl4v1TakhKD5f7YSZbm8xW3XDb9m9upqgBBCJek
VQFAtl/xRZMosmO8vwqfpkFL45rMuigLqNn1GMletGHyuv0T8wotaCqVkKAcQcYV
V083xGlYpCbphgj7efppHxWmkc18uy6S8WcQrNVRXVv9cO4HEXzVqzXDtBYMfLjY
AbqZvFugry5NMJ/TwXsbyXygKmKM5u0etcP/lSOoyVJ+XWka+qgoX1+MZJ95WrNg
QG5WCAqOTpw/tMjvdpFcgJal59F3mBtckC5kH4ItX30NHPCC44rpFqbkuQPxRrbN
zMX49cZCLq63BU4caWefazF6QKF0dTO31rfvtLUdJW99EuUWFRPEWCuZhBVKPW/Q
xkZMFTibpVw/XD3FYqBiSesJ6u4SEUnEQK2+l/YLlwIqex2wC/o76ia8H0VNXk5r
R9Ur6QrbEnrBszduJK0wx9s1BaFU1sR44VE5wd60z0vDE2crx9N9ANP0F5f+pxtK
FOisb1X7eT9ZhxxttnVF0hBms/LX6zBObhMuLlD5cnCVJHduEzcDaey5OojgfQiR
CWqk5VEJeFxL8LwjUIFE3SVXgjtq/BwWYa065TiXE2XyXsun85KbS+JvbGbkuIFu
Ht+vsrfCSBwtW3pGq5BNL/NkvIDcQl4KLvq+73vrL+oLrhFCf8GARqPIN8Bet/ca
aiITAdKlXWDma5xgeWwuXtI7OVPdt0dHg89sSYIGjRI/6otWoxzLYMBC9oAfvr7h
h7lg1jHJDs8lSDORlTDmz72nUCWsP5UDlIkCFh4938/tFse0n6HOPUelfuaggk8D
t7OlukVsjy77UgIGkatIcN/Skg+aD/HixWzdumirgs0J4K0zdydDLwAfLuZqqh4q
L2KniP2n3YXTbylX5Xjay9PPg1TCwP8GVAAEe7awXAumK2L3q0/5L4ycZTVaVwA1
vQ1BBy6Jt9aSN3PWD/JXPZJ9/edzR7dcGLnGb1YAMDmxalfGH6XexIain2fPsA8K
Ly3OaGUV+CwKrwSdPyw3jehK5FyEXxFcktFTgOX667wup6zksIqQj4Rk3dzbEeVO
HAFxL9n+KSkvgoYo87qYTjzIFBiKh1jhp1N7/+x+NWdx8MqSJgmszl+dtjAMf0f/
w5w43aeTxehoxA5Y75NpLV305e9il2o2goXkufffcgCosAqJrNwxXuEp0DxG2XaR
oHoqpCbuaZDnqxTlsSvvLaG0QaRWq+f6iY1vy25lebELmJMgmsOX/5eKfgYmVqN5
CbLLlu/PyiOb4iHQATbrbJxmVbxiom2wrP/lNI1wteg7QNEJtaD5GQR8+ELJQnG+
4E6bhHAdKkxLIUoHh0Lc9uMMEtiE5JagypVY+1oLvU7VocXPNsft2Mr5v27DPDhn
0fv6qHeKXmpQdMVAiTbA+krhItH9aPFI+ewBKvgNlaq8ks55ezLg2lyM1wHjupm1
taKvQ+pqQCl0iE7x6oS78rp08vdPn/BQTBqBw5JQ5yMQ+YVJZyAUwRukeg9tgyUi
xVqMn5LNkAXaq8yAkudZYMktQQ8gJYRgXDxz6cHhbCV1aeJGxhv9r4/Vu7i4zT4C
rEXMXf8rj9PLkKvHjn7Jco9xZEt9vm2Qc2r8askigdcZIcVDmCqV2ShUFEdAbkSG
eXNssj/qeNiZP4iMvDX3t+zGs+txsu45mlsi6Va90jZ2BrzFSgGA6XokY/EOVbSQ
QWleHS5aTl8UGm7h4sGNO1idsfJ5zxOSyD62bqJYR8ZFaXzURWLgNICtvDOqP7Xc
q9QvikStxHWocvpstMHshAy7CVnLYA4Fdq1wSrJD/OfsxK04NcWn0ZA6xTrJD4LN
YMdsUuHdG4tZGd8QCYUZK4oq+alBbu5GR1qNloj8RABlxZaVc/vZH7M9PxrSGQ1q
jpCxuECqwPHJELl9BFfhiWzQuzF8kbB3PzKFPcYxVZG2rXrU+vf7ti2tjdnyNMUD
LzjvKchVrpoBs9g8JK7HuizJsibhafUkKUl7GaytaGvAVTbnMWIm7yZnOTXo8q8E
jLItiV6Cne5rjgnB1FBa++jdTFyMizLhmYW5LCUvNwDBT6ts5FSLT64xdJ5eLhZc
CZD+yo1mM158cBheTWxtCP4DtJNNH0v0U8X+KJLmKwXNyMX4jxKqxy7np1TE3DBz
pd9QLDwPnDtP67lwiVjiQBDXcYN0rfgblFabIv4DwgObdDa+Qez4XVbfHenvIuot
9O4C+NV97cM4sOeLO2dsgNiV1b88KEMfx5D4S6xdGM/uge1IKxUPZ9eC9eMsx0QX
l8w9VUX1vNm3Bi5Bx0Z2Gi7buAJlpyxK7MiJCZPpj+B8kyB/90x0pXSEMfBT9NPZ
W3PVzZuTdsomhTmDn00D+DH5P/1wHHpeo69VDQK7+6kEET9m834gubgM13jJIQzr
uTfz3jHNYUMoFT7+qZXyNammEukm5TIeWgvCidvryfkPbVXH/mXCBN11rOZMvMbk
SHto2MJY3rGFJ20BBLEmNVkYI/HxRkt3EebwZJx+f/rIO7RSHAMQq3cykpvU4e+I
kIVI3+I9q19VN4xcU77G0VvVmGkSQVlKD1LciEM0U4t+tvdHfO+0Ahi6rAGT72iY
aIWjdfVM7eacSdSmf0ow75LySyqLal5foCVNp9l4r/WkCGqXOEmYLDUco0E2tKMQ
nEryxtKfQeNr9WtJwwzI+0B/OBjQKXX0UXKFipBIHVM40OF+yTXRPRf7BL2eQy0D
QjZ4odV7Gk09qbx6RxjShwkklg8/3X/BCS3ewxYJuF6omWGGv1L9qpSvFTuWCheZ
g5EBHCFANwJBVxVF/L1zghTQ6lu3ZJ6B82TLoz8LpbVAM4OcXGnTPaJMWc0qFNIZ
JohwlqCgdEMhu5qTMOMaWX5RcjjZ48U7V1qKEP/C7vxh5ypbIWLa41sEGkpfJGgx
xRcncX7DJIhLVoxkFnOeQDz/IV9twFO9CyPYd/uWFwWyBLanJh7BWtZDyKnLciaH
bcf2oe1tqeLKhYqOaX6Q+RXuiCDUoNvpGDBSKDbnP5W3nhPR+QuO29JhROnE864N
7zODGEaKmsoD6/4JN5Wc7MmH/YCGxe14lgsgsWh91W+bhB/o3PWHESdsKmTfc/g4
+kd6PLf6g3h5XsdINjNOWqrfHUDVQPndQXO3wMXfK54goeLl9f4RscvSi0xwKcZa
fxqngfRe0M0VUOHryWOEoz/eQDzW7+b30gBoIWGupWhIhiWDOM2txQOfSgD3Babu
m36vPcKLGuzFlThGb7F4ZYf85/gtu8RULdS9UOwiviJWF7ISy5VLuVb1U2wqfOuB
hPrQXCRChVFPd0YZFUMhJH8EjWSzxeh/IftlTdPulD3P3AdbushISX7WZ38Xxoih
mJ0iY/m83lZkVPUhlkuwnK6+g+8KlO/sMtjMq5XIFVftFQStODHajWJ7J6OV0RYQ
65t+pSr88FDzRyz2bCBxzTwNgiy0y0zfmuxqbQDn9VoLFD5e9o9k4M07iUdjjnMz
1r5yYBAITUUNjVANOtb75LtX405Xp9x96Z/X6yg6/cQrXVVfYgXIPavWeHEWkweD
0HB1onumc8JgT4aao0Xg7mGNrWn4T7Pr6Tk+mpDGdUdBqdHpjqr5RSpsTyX02QDw
cB77TpkWv3dwFv+hkjSlLuQFC2nZE2cI1BSmJsdy2DZrTfZZrxF6WXmK+SnMsZFi
SSSjsMntApX0EFJFndCjfQcrpOuaNJ4wFWBQCF95iuYgqB/WayAaA+0nf7mwsD//
/xqmTZUECAkIcGqTyk0euUN4QRzv92P5Iz3Hv6bQhyvCuzf0GsccByXNPOz3w6oZ
sVda/QVFBFP80YPqMWqjB5Ax0ZVfqf5BYyGNd8JuzXab7+nUD1++1JY2BRPSAxZ8
MCROviJP/u+nKvlykV/P7/RVcadgeuyoyvYvxCAtybTV3/elNFnCBAx817juEeQz
ko9hpvgehfpV5RS1AyYoIbBFwJ85WOuhXtxlb3sq2si1BmKKadfLmFQYgwXZko+s
ZETDHA//1ncbsXEeNW0T1AWGXuDqovdLptW0azHud7fHNbYv9VMSMQRs5LUy4hO/
UtxdawQa7kuuDLesfzg8HhHd5tgnMMSD8VvVuo7NxZ3XqGZEbKKuWWqs4eAen6Ia
+NHgm4aeCemHsa7RG5mMqVUPvt4u4FAmCiU+Brsot2hgI7DecgWmDBBWJ/QgUHGY
mf1GA5bgWyddr5jQk4y/gIMoMQhCi8a+uqDKyw2ArTnL0LYYE0yTyJ/l81Q3H0Kp
ONp8/f+gjCJ+Rl4cumWsUV6Oh66VN7/POtn2+1x7Un0i9CqtC/ERNuwen2ChaEhA
5euDEueklCerRfMv3sQANeh8CA6LsZIBpi9riHDEEND/Rea/ni3xRlykGiV0d+8Z
RO5LfSUhIDYnky4LjxmER6JrVIO4hG89tkD8kzc6MYcQgisl3q/dauOUrgk8c5TN
A1wKu+V3uUzuyUwtcT8MG5AvjSbOHoqM/BFQyi9GqVgK8i+hMH8bRCE71gJOdKnq
Vln3fE9O9RyLxrsWLMo8PcOdqRb94cFAvWGWJy2/w2t4sJy4w8hZvSABXakBsQaK
h3DReXaEP0WwL8lTG0RW5qUACJ+6UknOv6Ovww0WJshbGzRaZreJbrtAVVLE7+7X
xT3NVWfIccQrfTBtOGMHecYghsAEUeaK6jTmtAXLGxW18QNJ7WWYckMjmtx2OEhX
QkDd3ulVkHP+9KyrE0qNSNDSf7uKFnBOzVuZz1EeLHBoX0K3EQCs5ZggTWfeYqiC
iUOZ6CO4ajYtgwtCai4uM/drc+AbbpENa3apQKoNujjNaIL0voKvOZpfzKEm7YpY
YCEUXyDSmE5EV9QIjWBDpxhi8ZXWhpu2AkkGUQYmVbEvYqWRwFr8clpvdTrro4gp
jnebsIPZOi1hVOT452Bok1Z9osk0W5eilsG9ZXfDfotHJPZSM/YTDzDNfuYUROuf
SMh4qFj7S/4kWez3TEaY+i/gGkSTFnEuD179som7pucuhouD581+hV7Fsq1SYRXg
+MrY2SLlV/Y1rA9gUScuFQnIcMRWftAkXcWrojhesa8crU4zzQYMOR6en4JbvNiy
elqIGIai3KM2S4vn9RKCu6fCkDI0FP5ZwCuoxQtYvaNs65Xvr6wcO6/ghFxcHKa2
J0Unqxc1cbJSNSCZ4E3OzzN2P+b5bzHNOtDSTst4dPJpmuxWHHsS1DkdjqB3SLiJ
eJddx8OWMzYhCKpbOeui5JwMtKyQVPdTsbx3ijnDV4WSJ0l9wUPvF6pkRSuw65eg
v4E8KhcvFljbCfMFA5+Vwi2rp5ZUnQX3vEIL0PXWzEkHyJk+hvO8lrwoKXatJIb+
Mt97IGjYVjUPdDVVreT/D0rQnKx58nHIUd1DCmfpUrUI+eiobbVMDmQieq1EPYmy
g6sThGdzFy9SYTDgnxNd2sRu6zbT8ffoHvp9iBoR4uZSHiVqrnIqwf6jd5BrxmYR
/AFIiJUICYX9gcRPFtRCrmX6/xHn6rIMcrQgV/ZFvd8mLaQcf1gHkADpq457xqIK
LyG8YjvJUQJS/RTiJIfQfsqVkycD/sXAFM42utALa/A4SWyKBU5xxgsmjyLt1HU8
Gw1SxZi/Qf/A/ur4NwAEqPpEl+kck2RVzI/cPphD6fC9P0WoO8PoLJ4do+eShIn8
NKLoOOOPpH4CEC0Gc4ljp52ZrITKjvnO0SpXWJI+kqk8FFTc9mEMy+Jn/CK1gNdK
Udgbh2YJ1D5Sjlzp3fMOf4j3kTr5NNnb18FyIf5wP3naYT/vx7e17w+jXxDzMcgY
CscWKDZmAumAXmf1nfktcPiLFpxi0E6SGNOZ+/EJd3gA9GSF9Q+NxyDDD5/kReki
LWi4bDu9EbeZakGWelUhaFjgMaNWP2S3yRcgAitNXC0A2iPl82RLAaPkwJ1sEdhU
uo+4HWa3WuDFXNclpdGwmU7RAbl3QDS+E+5SKr7apucMhOODO7m15tg6kjFsCQiG
POgXP9gXiY1KuV+DHiLWa46TPi6IqftpES9KCCCBvjs9ceW9EiNZr9Yj4uwPU1jX
NxlULfy4mubbUWSrGJRIEmHQkvJPQxIvnwPA3ale3JJ19Vp1RLW/A/No5m6SJh+r
GwrJA2EUO90wbhblpkVrlSJ0f7eIGy0f2ZQDm2zrWBW4/9xsTW5m9ouJ3jGCz8zn
VtJogp6pIxxfvKU50m5F5x3n/2sItUPbNp+Kyswm2iz5f9j5bXAYWTP3sVBhFmTl
EpQb8Y5nEYFQiQQJyvlfL7izFwPc0/PnbtAPTU5LuOo/oqeZiws3MG1Y0LdPR6c9
0mBV1WtkqS/qWS111FjNkuWiCLVBL5OqRoZ8HvkvCQZ0l72AI2MKh0TqXy3hC47/
n77BM46UE2yBfl6k0GIHerFZF2KqfPeQeucHpT5kI/C/2g17Cff5WRfYdb2yVd/R
Ez8Pkfk+1asgfpCzJOZJ3YDMEEvnHEgxL+2CDw7ybRmlqrDtwks7QEMK7YMR72Et
zQmYDl7fv7HSZ/vLXzRNFAZmNIcn9oJbxboGfybFd7+lfNSI+SyX2esrxFJNp2X3
c1ZfXdCrzax9u4YtF2EogspU1qj871Iv4LE5IYVS45HSR/1dAy+hlhLGgFxY/Rq0
3tEO9axYd2JJI4/Zrt5mmTcfwJwhBjxzQC35VcxdjGcyEYJ68uL0L2k2bgVT3YBw
ZrceArZLduw6tdjVz6nt54RBc4zFMmOml4KK23yqx9kCV2T2UbBZHSFhJLXt2/mm
VeehEpDtk3B/KIX+fGj/l9+u499NLthEVdGQWmF2/dgKcQyPcnwWXPCHWLJMY6qG
b1EqwaH8XpDsk2YeelsWDfWVI6PPKdShN3Vx2534aMwFo6Vy3+pUrbY0e/olj+ZB
uDXX/TcmHkSUzOUw8uTUSfq1agexCF7SWrGc21+1Edky/iTiQMU3zMKCykDalZ8l
m4/1018fGVVpzBPesuNJ6Xmq/XIXmkLexbBNflfBqMSNFyAf/pBl8BdZpSl4/ZIS
5uwEjnuCRB4LvQ2FQ8h673oxmQfJrIV8Y7DXE+rQkw/UBx/a5zq4cHz3v36SPXjR
HpqyepCA3De5OT/ogFOxLPhnPcoVhqveEVCGmFXlrZRIDDYNLjjD0c/xSJ2bvzg+
IaEy4sHQJUMsO+G9IHCVx9b2se/2YJiebA9HDc3vjw0F8nrDV3wtsPDZEyFePtsd
WAW39PGNHq9DqRuvNGYsuC86+7mU08UI97uYIDzuCC7dIoH9uHIO7jB84dECubKf
vwGN8lUup97vtT8U6ITBe5nc+5bvGtc0RaNhHRGycT5XoMjyrN+qD/TCQdir5Oq7
aCDxnKoImWQchl1XQZHUjpbCS7R4EqBiQ+mWLh1L75Egh2rlsDbhdIAFgObBKyNB
tnSuozEKYEyRDQl2OYFHncJK+aiJivi6s7WXUMqfcqGGloX1kIJOkkUQcGPErcHt
ZzUt0+pVLbTnjjldkYbV5XSBlvSDWqFpzdU7Q8fWcjKS778367yNmXPnRIgqYvki
du0tVblzVvXwHzS3BiwN4hxWYYD5Eaht3ch4KdMncCXqe1o+6pWCsuO7XcGzkW49
VpZ6CWMc0T385cKCrJse9AVhHdnpwOUy0DIKIEioJnTca/0fZee4wO5LIf3J55N/
/2JbhRKyGfk4o9ryZ0semYjUNv2YIsbHuXXv5MlZHOrxYohdG12uFBoA+Tk07AXT
FQ7rCQmgpj3MSEX4bpwhY3OFQS+a1FBRZcN2tUnjugOjzO+Y3yQLVmt85hsesmtA
R6hszUxDKDawT8kxbUrg83qmx7RD1r5MtP3SkYthwkDoXitLHL4k0XUlYuzOvvKg
khRQbAm1w+jFacnGroVS2rXd4KiR9gSujXsiCCrMC3fZm5PYz3mqkOjemiRofjhv
9ZfXUYkdkhSLSVKP38n3dS0J1r39y7qFszRk32fDQpEhob4D1dA5nYkWru1gSHup
3HSNgkEeAJG6k24dEXLdnKc/+CBtockRkgvjVQxY2zWXqV9U1ELQ9/LS4x8ejilw
GKIK5JpF5pNklATUXITPf0ZUI/bEDmErRRpMHLbLHioegohycPc/sLbsfPxNKMCM
wmAdnEZtFeL6hJXDOAGn3at2zqL2QtcUjreWan2BdEI8csOC7lCAr5aVKsWBfraV
+yzhs+SZsLKxtdBMgkBB+mSOJAKBMcw8kQOwQft/eYZ5Z8sWTqFd1ME0G9bLMsDb
sWGK9QFrgfs/x33ldY+jbrNZyL5oodEuDEZCaXWCJAt/mdjdLXw9DVmiJjKADQqN
5lWnZUmzPnIu476UyBphylNjT7tPLdSwQqpk1vRYxm6++i5mC4xezqCsL4ltK+9E
gIkQvXVnOTydzmY5RHppvjUGdHFPW891fbfWy/FbNN2LsjaMZNFRNIU7VzytB7Dw
MUgml/m54NYZmKK8w9ITXRjLroKX7E95rfR8PrBsIKw9qY8h3b/1Kx7jCWFkllth
fNp9Wh6hmUi8uzOQvNfkATsDd3hyiBA4Khr/uHYtBCNm2LgETRD9iX6cwNOiOM1H
seovk8xQHUNE/gtOII708cRXmTuLs4sGesMcu7v2AOEwaeZDFwM5L+P2aCy41PZo
GOK0gz/lknKcyW6bS/uJ7LBUZNArsPrW4sQ38mr/Sv+rCptG4I8r+BtDaBn3/aX/
UcDo15ytxjEoJSr9yY9J2UXVzbhKD/qYlDY+1CYIbEP0+brBBz8ooxba7LBiqNRF
sUUW2xQcqPKwOuJ4N97/CamGmOXmSRodkC/sbEZVV1G48sFyspam0hJ0FEfzboki
eALXq7FQ21ML8Tlw9P1iil663nctjFAnvtT1//X7yXGcwsACqISMur47glThYXjn
yw0l+toskSfkeGMoQFr8bkhRsVwy7cwr2zeER1wfBo9FalI1mObbC6tWB1ZK7Xws
3VRh22NN3Qhv0UVKRobpvffXmB0uJ8lIspqxAiHBDEbruhImOQHaAyOtvOvo8rIX
VMq5QJeiJeBBLrAxsVCqA+RVH/pS0WVW8wCbcFk6UbFM9IkBZK9YdolaqfTEvnw+
P1OVTAWu+dX37N7al6kLkWeWtpRTUMhWKYnLwjX+5Ctp05hQPOrBdH+0UwdVmZ4o
c/cUplwUJLxATI4tEz39sDfhgurmW1wajzsxxGDq6cRC4OU+7YEdPapMptyFbVhb
MQRImcJW/wAj9wdnPxnKIferN7wixJ4qJRjRx5bKuqS7WRh8RK7e1mtota6a1JoX
XeEIk6uC7an6I3Z9J6k2m00/oJ28Wc9GBFtNxA7dQbKxQSNjleNhHgMFCZ6exsIc
aMQrYn1JImNj8X/ula/gMssi4g9UbPvgkaIQcBj6CJLkwNBe6elToOAni8q1Hnrn
EXeaGmbFrprskWWcCyKkSeOIae0ApHINm+mebfH+WzKQ8yOubMH917B69OqbxW8F
r8BGMpycstOX5kTfnUeT5usNjGyoPkNSeqkX/p72vDp3cVmyrRGBmLv2eQ3Mznm7
zujmTK77TgxsR2hgGyhONql+hIILA2JCT5rXzPw3ZX899RDvD8L1ZsbOQl+btOOc
7vB11gNfwAxf8Fyu6kC9HuA1vTbqivbapyRcWs+wdnZ2SpcUpVMSyAqf+h3b5rY8
GtwQSZrhuwwM/Fr/MfsWJVG5mqUiBLM7KtDoQaMqqat1LyNOvbvjOyYROL5jf3jW
cCvSc8TcLYjnMWHD+vCveC6dFCJVdlqIh6UbIeVT9L3+0YLjY8qU/jHw6EUT56xg
sn/UDOQChgYt6crty0Ro5jNS9ydI/Iu9Ql4kjhBiCYu9tz8Hj8RzYjaHOHGHzcpE
cJmXxEPN+b9jWM6IPWlySl3TF/ZSP9i6xLnpsQTKkzh+YxP1WVJSiczV2xehoEE1
CzFSGi4s/2ofN9H5zoMiknPeGGbY6x7Y9PfeOMxx/zWSDvGRJZB9ec4Q4WaVksl8
qvOFt0447L4kyT2ct7rFw5xn0drxUiQgIBcFsWelsKuUKRGEpf4AJKoKlM6EMPtd
gfTIsfBVWUoS1api6W4F9hWjZh07NI5tXD4vJVU/Vjks5I2QP4DdLElx2HSuyISE
pWUy0OuBERlo6wlcIbrsSUlzsFZrRcWXcExI/12i9Ci+BZo9b+LkyGsfwDT9NRh1
zOxU4527Hz/yFiyyVjk7/GLz49NpWePZDrkBL+kcdqrg34Mr+J1mRVi4vduiv/6A
VJfwfx71/LBwixDIgl6C/YANr6skQfEiK5N/j/GrwHOg9K2EAejE0jKVBQ1krbXJ
eyjA/1AOInslMXMxuSKqAWd2b+pOQWSoqs5Zo5gfoUiHi1Rs2I2ULdzBxld7hL9E
A4X1911rr8GupTlv4ypoNBeN3uT/jzaNyRDmFJ7TofJ7Jery07MHlmY5NEgi4km/
UZNMceXGYMrJszCC+96u0c1600B5iS7p8Oo/b6OHmUdhwqOcjmlNVQSmKt3ew44q
8uKfzoBC8riG5tlp4Ipo/WlPRJXm5d6ae6pMdo1d6W7gVgjLDUKsmw3Pw1eXYpO+
9aAWF2AEjALLmCCB3rlsVdzqu1Tk+PrwbuW8IGVC22/FCDoslOGRoNE8hrZP9FQ9
wu0l42+q+6Aauigx5eiRYTWmyRCEY75YG3NmWaPffC+2diKkAx94yHSEF9a7hFoG
pKUICmBkZAFc5ihZt1JXzZ+ZsZWYuGHobCFYKOiPNQqOsa0sTo1wjSjShTw8i2Qo
pxd1K0q++sIR7DbzGu7C+koh5S+daiFsLK/DM3bTPJN4IjTnp358DmIRLcXmOId4
OFxhgq+bUK5MF4tUQaQCZ1BnmdaPNhjob3zD9kFCLLKUY0uaQqipj0Du4ZqheJCB
xWGOFzk0Nj2w6t23gYN+ARO8kjXn29d+KUhQe1GBR+PluslklmpnaIYK5GxZGDGe
0XtDUb7h2xl+zGJBAGk6uzVAwnJGzB8jfzSsXIH6c+BPrDLq27lZr2lfZK/E4IWS
IIfCedppXAx1nqPZ/qqA6ygxUoIOxEIuI0yGbJFojfIiweTv5xXEQeyvmJ2j5E1X
FxbfAg3ATO0hcmjmSrQPJf/8HpRsiKiyiM7sjJ9mVl3b+UgKiYIMEQWIUHjSFu26
TgpSvYDwUfQh+ZaXPCSvPIeNlUQsYDwqN7ao4PK1SkjYN3GR8SXCaZgMYhUsoJ5h
MvSpFRYvS6s+sFw8Vf9eXvzjfoIsAHFxRKc2yCvxh1OzwGGGMgy/QvSOLJusCoZ4
lXCN4u7IDsB3IQxisb/P2Ia0k3iA0d8C0T+CWnz/iJJP0OgYDIOCpN4chSjDbw3y
8yTaJ8NdeKeQzDtmBBQtXKDMSmDs1FWjF/QRp5tav57u1xwL+v7R+gAOdNY3zd59
aahaSp+/trjOu8tBLaFrAviEu0ekY+sexvsU345xzEBgZ+3AbF9TIZ1crz9a8gs1
Qe7dESa23nKjvFLbx6eWvqI0G/3tQ1HWY53Y2VP9u9H7w5fc4Hzr17G4IxZEFh+f
I+BlhejdGh14wJGTqM0Ssn2wF5+xmrP2ylwd5dzHwtZjFXdiGzFKO8W3FqOY5jem
xDBqcHWItJ8vzUb7ZP8F/glNOROTdLTGHzovLY1+5WYf/DnLEVtiUWDLq07sUJno
OrQo13+DlFvQyXEe5iurVmvWYGfv/dnmDH4dkM24Bv+y8Ql0FlpKixn3zW/gStMG
4/5CU3WrIZvOZIaP4u+i/ICdODNz0ih67on54ZNNgI+tRT7JDCycCCQhSAU6ayL3
NElgctiv4ZqyCY7vyQhYxDEgMt/MsS4LIGaxdWsFf2pPtaUebQC8k50ChnlxVbqB
2myzLK+yFsg0nplFVDlU5p41T66Bhrye+6nGPunmZi+L+8hbM8Qq0e+azs0jzicx
NLSNmKlj0SvAJYD1/Nxa64jPl0fFIOeJcJINM7vmU5yvLebwP45+K8CDKZzGAZgf
LYrWP8F8CSjEeFGzBrnn/hREhx+GhxdQkTWlpXrzqCLMBOlzplpfK1KQZCbVa1wo
molmqDY+ss+/FoOAE9qsW/IjauYpyZmewihfrd/WYswN/28hqTYMOaqcy92nTv/Y
ijAKeR6pBcB1i4zX6R4XGA76SGNnhiWXZrlE1yUYDaBs2y/K6enQR7S8peujaZKA
8xhq11J4ktR3QOc/nAHGj38QuuruHiUCXO9q5t5fAb6bQB4S0VHvdb5bhKuJwU5k
AIy0wxeAPk2+5jOwqW1ADCWQ5IGAoWgIlmpHZIlEXRvuVp1uO30wfrMdN8A0IpaY
cakUmKILiPfxqOdedjuQ1z87znNzJffLYkwzRJRH4Ql0VE5u68notkkE4c+vwoMX
JId51e63Lo7Mu+LkN+snvl7EJgyewYytymuzzgzXs6U2PoYh6CeWaMfLS+Xgix2g
SWtBJquXzQG6qUqQ8YcsxW6/sAq828PvmWMterQAQ7ru/DOiVm2e0yHd6DgxVk58
yrc+nhXx2RZxz6rFc1UBDNMKsLuM8ELJsqtKL4XYu/SGueXTp3b5Tm/ZNddopFO9
D3a8dZiW2V4sAYtrc7nw2Y6T2gaz5w7O2EMVDTeSGtk/Jx2wnaWANqABiuEETH1q
BvluWaIQq78lDj0s8ahsFrJQkr51OhLePueGqNHqNhLCsUClyxvL4sX6d3PDufSP
Cr/1TMV8Cz8ehvF2VGjbxW21pUbcmWmwVhSvJsWYVgBjYThZZGZXlZ5fS4SWI6xB
I+wAjQBHZJWVwBoMTBKFzbTQE3jAyBn2/XUFitZqwxgEOr3XsjLyMYC7K080dZbl
PhCksTcychhEUaM8mUD0PJaNyJhCIhhYXVkS/jIefDdRuef2dZITCMr+XBgn7OXH
a1fc/Plpeax2msQe/fKuRcqOi4rqXqdQHAMn4EHda/DF5aepajYWQeWZ2QeY9qg5
1OYt2m4eaHxsIcBuDSrrydL3GuKpKqTILTIZOc/hUiTzRNbA+LfWLETR8P786CTd
t21z+H4zyViC0IQUqNxmUNct3v3qMSTe+KEVTdpzkoKXzsMJwPSLqZtyZxcpEjqF
cXYm1Yl9X6FqnGLRMxngcHL6ID/+afrSzhhBJr15KoJaJx9p/YmhDmhloTSKNjmv
kxFDmrWLat9GKiNheuQM9oDjsHQse1/1QNLf0oqwtvsw6eCZF1ZlG5G2HYNKj/C9
aAPpcvmACvUCGJppL9y5JS8REggis0tOSTCg30GA97/uLqBun6YgeoOtBrRC5NDF
5PhCcw57ovVb1j9wx645Wb8Tg+nUi4OF50U6kI9Ehr1ZNJ0HZl1cIcbwOQoioQZq
0uAhlvJ9uEePSQBpIqCrLqe4MDAyhoIKXVNqEGY/LfQyaXW7yY8fKFSWV9s4g+Ca
1jQwFH5i/d0gFly4oJ82ZhqNJU9tnOXm7BpaDDLUbsgEKLmJIUWNFm7QH4pyQNDV
qcddjQZffGCnBG94koR6HK76l/uhiklRic1nzruUVtNjpLshp53BfIRF5I0eOSyI
F32+R8TlT5I54d6OeklVcK2jrZhvMxXEqxCtzQkzMYSxn86iiWYJdAol3tJbqB8f
0qcz5WgeHGkEkRdzLYCPolCO16i2+ahkEsgnByDlfErCbRD/MR6JVRDglExcGHH3
z6M9AOc43YNCWhu221ZxyJypBVWd1jtYt6zSlE9xe81ZeXu9RDA/h4FBNaigvWhq
b++uux4ZkWl9U54dM1SL/x5K2MYxxXXfqpZbdVQPdY6lJ4fmjIBgyz2TEpWSuHnB
i+2V6d8ZpWfDpcyHSj+H+LrIfFmCQLbPOo+tjoi+hnGoQQv5vDHGXkMdRqwV3FwR
8E5AerrX2QovNBXCEcpwvbLh5z1SnSJZ8dbPx9OEy9nwF76p8FWKDQOudUmHr/SI
+3kenltskeSPjRX10kWP0MrcIfM7mUPVQ2HYbphPd0bGFRwk/mD0OL4GAlpmP00l
KY3Mggihod/H0pIcKw/kHCAiZZSBd1p/TUP2sglP3neXgplMmU9QCLekRdA0GyoP
TQlF7ijlB1R9RbLovgbAAQPTk1ZFyNlOUzWLuJsRozKUumoepFssLTLIOSsvr6xg
TNTqCEEST1XV6zr8W2u6pMzaEOBRi5GIl80jV4TAz8lOT9mXTF5LdYOW1j3sHG4Q
UFnJYWhqW3S8iFWDv956xI0kBijGrFtVPbMkmAfakKK5tA0xzidGtlLtmuPLjqKF
2JS7PDUxMrY7jOIGZbCiN7vhvghDd9oq2neRW0UFjxPJrZPPxN+PCoBjsf/Y37Hs
4xUbD5AAjHW/TM1hWoF0KBq1hrBWB2Nc/tS82rA1RaM738WJd4O6/J1tIbGGfzZK
rwo1hZoVERFOBlhqc9J+Pj8nAhe6wx0F0LATp4W/Mp8ISegj2+HYi/JVHKv9FSeY
v+vyhewN+nY0dWlab9o14TrNHHcZLBrcrVkz/vXG2kmoNpwX89BfmR+has+SHPwI
MWzOnoLt3xiCW9DLPBPMLHSoVYTadgwJjVl8VwVylj5j9qfcSnE+X8TTU02EN8yJ
efc+FUIivqTb+/OhymvhxPD5xDYieVY04dOQHFNNVI2WcRlcLjOWkQBdRjMMBc/Q
LAiBHwORPOFCmlCJrqVgJMSqFNITwV8pme2uLNiXUxksktNcEFFJEvp7VfBDMcwP
SlkHIyMG+zHfTco96ow/Aw6N3SQroqRazZBWuZAzYaGOPSTx4gc69KTVHRgrIznR
JIPs+2B+Ox9U9z58Y0ilsnNFJsx25nIb8sTzZivKaiuJka9Qe0E1euBBSMLPI1Cb
xeiP44rl31ZOeCl41AbBmMyzrBKL9EnYRyRTsRi+FSFCRtkT9RT6hiV9GNV4p3hw
RWp7OE1Iimu2HHLwibTWGxixkgUIDdLrDsyWUyeZ/xeiv85Ns0UjLCiOBTHAyoTx
SVUV7KvBHqM1NH/hT5GpfUv/8uLsADXAOrbEq4ia5b6m0YwRPMjXykVmmpqJ1D5g
1EvRQb9HrB8PsljsdBfQv/jtpKqN6BGc7OrDfyo2QD5McaN53UygpchijEPGGXMK
SiUiLdyf7uizLFZdXsBSfJAZSldImZfQ+k8HCudiDlvPhnFkdHdEqM/rQ7HB90BB
tO12MrRdBshBqTmHRfVlBQ/FCLO9FT7/uOqwUYxurSkHeP1LXpvajrqvyAawhFyk
0QVKRJWXHhj6CDymZXAXvDSZU9Mb/fXUREQfeV5DZDaohp7iwptXcOHkZefXOOhP
yjWQnzyM6k82pViHJNE0sgHrxpSh02gTMySWjagmZFuxNkXp553Z6HOOoQ4xm5C3
Cy2BqUmrUodCP2NFb2K9MV0a6P01S6qRRpgShjWvAdA+hm/lk8F1OYuCFgYyEtXn
WsJ+Ox3xOnoabDIaX6DN+DFeaUbi7Axmy0tfsw8olw14PiECrl1ltWGyPIIY7LwL
lj5NJh/Y6CJC7nH5EcH1Bb+/JNsAaW+kyCszH6vHQWkRyuDxmVQ0XxuVtiYZfKYp
ZMLm9r/A6j6KVe0aryOGuVAOM0msjO8NTwZCEaBFoU3WnifCpfzNGLb2sZBZPHpC
/bPX4AQZrHTR/46LWphPv7ebwL+khvvsShbLm2GXddzOyOhavff4KBgbjKy4Uwgd
j1uG4z5EShwguRKzujscCwtqYy8UUPhzNBHwpGF9huzilUzdGK2vipZX+X/45Q4/
g+etnZWKb9leEYpHror5LPkRk9kQBUfDRcNr1H2mYnPDoeScshg7zcjdLkXbZ++Z
d80MvRGB18M7eD47N8n0YwqBLSFKHHy+/bZ1R8S/kK5szc1lVGF4jeOpJTx7UJr9
ZHOneVJHEeFl2J15qzfvPOlNmiiEHFyVzibuIyUOb7fQDDNuc53b5uW1SIvrYhNh
ff9WjDcn/NsvecK3BBMPK+WzDkzMfNWbZjAOFO648rAFx95hf6OzPv/y1QWrnXh8
ocLEWcAQ1kQab8pUzzP13xzZhveh7K/U/wW36YVPHTDJ6Rbep7+q3ChR0Nws9qys
X2CI7r582otFmkZUfqYbQcyLX9BERTDD80x+OzFln0Oo24SNvAj2/2SJKs/gOKMn
9FYm/PLN6B1P3VoIeARWgGIYTpmn32h0MxO987gyO7F+7kFYJffAJ80V9T/77+sS
i/k8SJbP+QxOiXKSMWE1uN0HiDxJCwC3cZKre9bRCflGpS76pB5L/o5tHdVycOia
b+cMT0zjaiB4Kko2RZdNSIWyiJMYBcf7p9IEFb7ycxe2T4oY4EXy0ANm9/k7lcay
FcI5ZwhAR9eq7nBpbbAjTTB7mT++5rmNzTVmtXmvi48HNFaRqdk7royqfso/2K7f
WehcyVux6NL8zDVoG8yOAD6Lm0Y3vMvZAZL0jypkQYdm+PE2qdkSC1vNXfn8WuTc
v2n1S6s4nmWuBzWjzb2LJ97Pp1D/hyKAopqZ9Z8ey2N0BLWarGXuOaYPVkbKbSYd
IAB1OrYeIbugA+go/199nofJdhU7HMfKY6lR6f3zlk3DNViFSDZsXthpBnyUCn4v
gtrKlN7pqGbC8DICGnLgdbgy+rCpEOvvvjy3IAObmY7Wcp4Pywk8JbrYAF9D1L/k
l22LDYBLFdCZqj92Zjo2pIumEGByStIoog90FRfN+4z0CLQ7YsJBLNmyi6qV2ZnU
erv8ziHafXyUg29sPSrMi2TR161Wmb/1MfXVdw7DF5RYTK0sO7eE8biGUBLDYWNb
v/truEnhL3Ohm2m9J40//Cg2NlXRvesssziYORg9LneUCy4yWz2ijFJ3ubq7XlQ8
6QsUJniktPMcaf+kyfyB89uyrEY9s8v7RHVPVcPD1eBD2FZ0dIhFJnj69gRUVdBd
EJiJH5je0xedG/zDZSrmDnYMz8PbdQS28gik0uevwO3SHy5jPrnb8Ius9stcK72F
EQFf/8gNyoShi1Q9aHj5+MU/qzoFCsMBYzhdkfzKBx3oB9Kb71Bd2MahO9lZvI5S
QCsghG8+uuhODTrG2P1R7CrDqPo+ThHnnjXWCow7+2D8UehyncxmfccYvckA/jsB
JJc+18EuSaD9nCt2J6S/6lK8r4CD6DCWjIqvJVqHL5Q9yTTBNJYE1Uxm0deSe9Qm
TR9mE6eVTihd3VxbM5bh+/deLbQ/urepATvekMPF57CvPniGAATmoqFEB2Bjrgzn
z/y/bKvtrWFCwEn0OWjoQGh8FqqXPdV6kvJXUta07GNy7xC/UUtvahbd+AW0KwAm
lPFpP7NQha2Ly7YMRU2xHNElWLVN4lWWHNXmBqxrCJ1s+EZvWYsrsDJo6TyuXDNI
n/FLL/vuPXk4Fc6QgEDEK/e5jp6SOmUHUxrvX/5z/4aorenfQnNAziGlQIjUwz7h
DC+F+YtqkfFuxVUyE55Q8PS1Y8jc0TYzF3PvXLjAanTjigOV5UJuC1L15dcazl63
VHcuC0LQtDF45gU5cziba6z0lr+TYJyUSUbGqBzV7QawTuPKNZSuzSH+07uBRP9a
GdOsrB6e4I6ADnnqSYzgDS0NecqcDqG2w6Y4GaRQPDNXHPq49RZCHMaC3lR/LP1K
nFMYaEQ5KisW5SnSZBqxH81txqq/ZTel/a0s9w2DX4YFGYXwQIrsr4tJq3IqbBEO
Intb+zsbkE5F9velmCZl4sS3D0mAjK3RW9SabWn6yXR0AcMj40KrJXVV16GJmsxp
M73jg6G6tjbbg9GZa472DePy3HzCfvypYrQens1OeKuFvDnYOPGeI5t8rbI9/lDO
S7AhyC44L+2+huuSDZuGKAoZzxPy/9uye8duS9/zLP2Wq4V6EgwGrs3a4VK6ZV1o
l1YSjr4vNOKFtsZp0oKsz+0MfyTgiKzlv5FqsEw7QICqqnYsyP9MgJm1YEwD+YUv
JvpsjSk6AMLX3rCZPTUHYacSgCL+7uTsmSQCETzaZfCN+OfMi2eat81R+oVzA5/X
cbCBs+Ico3Sk1T0Ng2U2pr9onT8vICpWYpcRH6VRlheOdrI/VzBLBmfKC5YDRbJA
gwZIUElaZwrAiUsdZeFJ59JSR4k6hqdoMRqFqliyq0sbz5FeaZezwqFajib5NUmH
uEZKPFLYysLK7PzV96m4LsilQV/S9kM18JgBiJcN99hUrEop2VS+uEAO3y0ShIUL
uSc9oTz7JAvFGuk0bggi1bK1XZokjYZNK+jpTpFsMXrkVZVhoVCildUiTm6f5YSs
MeY3pCmd6/8wIIZWf96y7wOJETwaTmBd6DV/ma3flNwKu3KmsWHAma5OZTfTot2l
BOWE0xal+enYGCGpokjKFYNnskjgyiiRzsRj6HoL0t+hgOEEvJVGMitG8TzOi1oN
XhQ5lWMrNJky7GkccnKTlQOnK67rq4KirprGHxTA6J8lleZaa/2T+UfdTnG+eg5W
UUl7qninEE70AQrFFDhFg3SoqUeXAywcYegSORA1ntvQHAcGMF1RZ5IKIULJMH0O
LiuUekUXPEEHCbWu6AYA527y+a4Cr5EUV5eeXVbuEiQlrP4loFLVGKW4nez6dC59
AWQ50L4YFT22hKDpoFXSa0pQInJYdk1H/OCpXKdNYpZcZkbRm9PDoALmaBVmw7ZJ
MCRrcJwnxgNmw0lmetgPBSDA1zwgT8PS9fN6y0T4e/PkefRQ8njO1uR3KrDKne3A
Z0Yjg6yhEQ1oqLV8E6pDbI/Kaz/sKiTsYEIJoBJBI6CP/POjvbwVMGubu0839kXw
8Um9K42cWhtgfaWzSEf8FKLH8Hhoi05y3blqMM5/z4WSOpl6ulmPhJmFHZtDptcn
Hu09w8iLDGi40By0tD4NfGSnFIzkCzadWPNwrOx0jAMLdYuPdOtz3Tp/3QeGHccY
QjZ0ulrl9dWcRmSXxp9xYk18fSJ2ZwavPc17V2ceKPoL0SgE15Dh53KMAKkffy/0
Eg/fLmBgl4RTADNW06BpfrQdfCvM+uvh02nBovXaItdJ5Tn2Sq6of7qg56Hz+9Z6
9xWmzVr/fqU1ySRXrwLK4tLdoZQIg4Uk5ixqUUTbjV4liDVjC/tnwaDDe5MdD8ul
yC776tb3npceSaQKNuIGyjvHKCpZrraiZLQNvDNjkBrafEXdOn2gXuHSxtq6fyqA
iFtgpiq07XkTTTyuqPwMVgFth0hynQZAh2WxHmWLtXYAUMJG6tNhGFBTfRA053L3
ZEwvegRK61kbDSDdP/EEFcyAVkTrhaAxBprIwKVlaIkPfSeLb5T6fwiE22lpk+s3
SuQd1+Mo7uHr+ADCMPGhdUv3MKAG6cgKWSfjMLLRXpi/WJX/G8CUe+AmXDooYEB0
QtRrw3REx5V0YBa05cvWJmmeO506ETw3zTRtjl8o+DRTxhFWJAheVKgHyEEddcHU
hNs+xA3S/mIh/4kHoRjxLW01G7uddoaYTNTQsaZylqn5kLQP11pedb9BIuAIelLW
makbV0xyANTM4dKzzv2qsHFqlgXZVsgF86O4GpZ+o97xfC0s40uLkyvdWiK0vlcw
nWL+Imxndvhjl9P9UVUlUG2uEyfFxUt3egQda+LzXUtlu9UDnPZMDqJEshwlTDPX
N/0FI0c4X9dw9gp2bteoYnq51rRwMeddTU1b7tz2oV/Smme9BhwisQF64GY2MwLd
JSZ36qFIrkYmBd04sun9A8PaBav8yPSOqPPQsW64z8qZX3G1X/xaXXHRq3GKPWJE
bBJZaQiPOQef6YfX33MUdwyWvWXAVOzjiW6NC60ywPY7obFBinxN8sOA/7KEOuRN
03T0Z/HnbZcQ0Xj9zMxhVU1dDRJCbz3AV3QprbwHdhKb+jvLrUl6odTQFQ9C1Kxk
RgEr5hs04buGqK+MB+aJNK3+GrWbjIrJJEnsM+SqoTkGtG3pxW8NkmUjFFPd/nCY
LP1QORpbeOvphWEhQP+SCWn71ZZPdeIqWXIWGC67CeTfL+FpZpHkTF7K/v/Jf554
oP07yX6XOh3QsPl05jBp/RnI9dec07tFzoOl8fcvF0d+17ga5t9GKANYfA3pp9Lu
B8Z9eIIRcXu+St0ijdZ1nEf86V5TjlG5qFIdChVfm/liY8BEzO19pNILHgAuCExH
k95DruVNhShxOIbqXazXC+YCbtfBKhpNti47tGkCiJ1U+mp2GSmKnngXrJgUVO4/
i1LsRoEEm6a9NYbsxLY9IHXrX5xbnipnLbihbdZ07pnjGsfpaGsvoVpazvu2NZE2
NxcuiA8IzFY8UGUS2IF0/G1dqS52IvvRSf2SJBMoqEfAMAvF3V7PAwEm3HubsG8S
247KlRTbLPCO1fwzKnoXll/d1BGtBKeVEYva4td3/GEBqW31NUq5IfNb2FyquToj
S7SYQ6p08f9hcIVck2dp4pPWU1N1JOnAsUuZf1H9GHbeesH5X819fsdxunZb66Ws
5IfKVo8IrID2TBDB+mskaNqCWXktPp73LcYNUIz3iP0QSk0O8LxtQm0S2sNrPRMw
3A7YjnJjiBo73pND3RF+KEFRaPIQenUJUhFSGyTB4HHHSc4aPvxiHjH62kz/M0af
iMvoduXvlGL1JoSX+94q82h/1rc9w0414Yv6AZTQHKiz91Mfxe4XQ4ohZ0tHgN8z
`protect END_PROTECTED
