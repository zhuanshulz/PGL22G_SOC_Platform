`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SwFtsXNuzgOCfDYFqRhDiiPczoZyymcVlHi9tUHxzAycnT5sSUQ6jPOzcBFhmZRf
n8+o5mJLXreYb+aFAjXpb4AqHfzvwcF4Ldre8uY3DaSvLQ00dJuIDvFoiqVErvw0
jG/qo0Awnnsptr7As3gm8lRA9mEZN5X1x3L8wiIcrqZ9EQzXyy0b7GOtPUGJWy75
MXt9VduiadnuxcmBvfZZ7JLIFsZ5cLRz4aYnPd2HhuEg5lDGC1u2vn3R96sVfDEF
Z5c5iFwg7ELyoLH5kRfElfzmFrWrBQKmkEhnI9SN7/erpm7z+N2pAFm4mq8ewe36
+EI/1kTxnU7XwF0YR6VI4zMvunbOUg4loraqLViqK+nCgaFhFUBSJMWh5D/NEVNc
2dCVL/0GQqjE6xCYaDGRS8rQcJwTH05ZMKsbR18GzpYCdFx9bEpbi3eDcJnCTWiw
c6abGdZZinmFj8wSseIBb5HIluQNobW/IjPrQsO9NF8xL8ie6Ghle4dRVm24tqBx
iroPPXDS4TNkOZ9BC4hYO5LQW3ikBGQ56CqXZSWZi4ScU8YqKe6RWHzWG+sgsmcQ
lkV4x9+DI677hI1SbRDwCcGgc27mCWiGV04RzAuf5eag/kzCbg/YrxTmdrol/pZQ
6KerJDduIO8LANUxgrCCrIqhJeL9E08/7mhnrX8y2ADcAtB5mr5vj5e/6ExvfRfJ
NLd8Q4N2SWs5XnivgSk3KcEFx3coQtNT4FwrSVar/TY=
`protect END_PROTECTED
