`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+p403eyu7m07ltGge5As25RzYHb3S3IUHq56D7zYJ4nwG+DnIKp9ZQdPeyVZVitH
lcTxrfKiAsdW7yCnprS+X0Lg0mNg6HhdHmeYfatq26FDXj+mC/auxNy59hCr1r0k
FXoWF0mdukpZuF1+KUfnfsP93v05YzCSo0xxl/OcEq0pzWHVa1G7W7OMYAAGB5J+
XuxQLqE2oGrxOsUlWLpamzX9xqRJUj6+MS8bBvQ7lxGIxouDL2BgtrwbcZ7HT7tG
JKV2ZzJDKjxqkt/FJ9E5MrinhGuz8jNojBUYgmU1FA6cukn0utJgNAgafxmaNAXW
Mf81u2AHs5m0AB82HOnaNGFoeqTtv8XKQwdq/jcQlENV2W1JygLIHQZWDKNVqxjZ
GLNevT4VeMDYhZS8abCtFea16YHrTF+K2hePKBrrbL9CskL7Tr/5CdG5HDOJPXPv
h1CPflfr65795qb8AOWcOLWjaIYyuPNKkQsXnd6PK5KUxqGSHQio5rWoWxniZsI1
qjyQjrssEoxE6xhAr3a3whSk7a5hRMqsQDfelE/mDMCurEOqnd2+jQjjLD7UspJg
AgQ+n7a7tYsYkzwESNblWc0Jl5cTlD0HRlNmxq08Gi7N/ETfSFPZ/kYcDxdtFr1H
I9O5LTWoiOkz3cIS07XMB1cQly3+RHZsiWsmchBCkuxBrYdaZyraSZUTKOrrvflS
Uzye4i61XmGLpxXh+kxHZ8+p/fyaf0AEU/UbeS2Sh3cSMEPg8WCr/6OQ1CulGLWL
68aPYBNHgrBwvwJodsKyTNvWP+LjAx6+Ia+oLXj7kW6W0brcJyU7dBlsMkLuNVOg
+IHWnCTeYX5r+gJeGKrCo+9Ld/wRJbfNan53Xlp54pa1ki9xzVDg0AQn0MshuLie
DDOA3BBV0q+Z74cnpr0nr9itPluo6qkZygyXaUgd9aD4DXlcFQTAAW0I12XzyqIl
6exeI/AAkqFdF0Dc26M+jO37YXlSG6wQPbIMzI6c7ZvzGFvEKNiFmhcBBIMgFoxS
28TM3JtVlHt4VEQKlO5cHxCB9ZsTOCEcDL+tgq4nIfbKZihIiCG1gFCsR9KIZOEO
lDcwQ6ICsvUHEI3sKVsvSqGGmRImVH3pLH7RTOkcHVFejA61Zy4K27BFSunntUAs
yKtwQ2fFpeD1Eyyo4zaWzrjUIUXMXePn64lIxkewfmej2ezV/V1yhlPkxk1PE3/v
n/gnmmt3Ip2yVEiU73mtpL8qrA9slfuKHpb9yNgSI/MTFcISHml4wdZYlkmew+Vm
oBCo9DsJHU73WihxpjSZOe51ogEFSLHLxmDCnFM2OH4IzkAoLfM5AuXs4xGRGK27
ueXg6GQ2q+9PCrVngZH/y8+90EQOS3xid1LAS2ID1Pn/h2ewy76QGrpkQBlSAoZ7
Q/AdUoQ069n8RaK4xIL6vJuNNSvQvzeN1dDU4pX3zsNVVDCeUYfzfOwWhFi46i4q
CXNNpzZ4icRjIRW0MJ8qnuIj7kqlW6YmRkEA+klhvb4=
`protect END_PROTECTED
