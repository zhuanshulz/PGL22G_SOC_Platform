`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fvWrU3pwYvlxPFC1WlnJ4BmHBTxqUOlZT6SB7Zj59ZkM8Uo67Bl3eM9paDtTUmI+
KpCKF8sjilBdKPo2xrAYuq8mJKg7aYJ9JHo3sxP9TBI9ygnZLxFun6mE2RjVIk4k
YplutovNLpmLjF2b9Zgt2bHXgmMpljKbSpmDamhBGj526pOzYVJ0w2MmRFawWUJJ
mSgPODAbRC+hy+bd9fiaCqqL7LxBYYRbMmyhJtX6n0dYi6Lc2JwzfeOGi1bUXXsv
NdnTX5i2xLR/xwfIzdcaqVNgNNU68Q+vAQLzZSgqZkEJft60BUfjx82H4kLxq1MI
4nvkmiTguyRh8nOnqDjHuspPrXa8n669gDvJqEQdL8VyyOI0t/XbtrX5KRyQz3t8
pfLrIwJPgX8KNLG5mHY/SsGSZezrz1EQbM/ng6X8RC3uiBb7e0XzoCF7HMe2Xc5/
ycUdgC3LjUMBoWbAvO0jOrsB9QluV/XGYQ4Wv7jar5WzlGbt09upmkZNZMbtqBJt
DCphkuGdKfkXyC1PaWsrBNfddN7bBwUsWgZMX7oGHW2pa9GJm6wNyvut5Mxm/Vda
TfGrcny1lu4YFNXg0xEiN5kCzvb1B+E4darl4/1wGg9a39j/yJ2M5FK0+bdl229/
gvgdo9CQDv0DYUy+WeGxCw==
`protect END_PROTECTED
