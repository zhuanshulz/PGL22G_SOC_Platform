`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8K5sDCaJ3OgYFDHB5DpJOVckn5HOEEkULPMuW3Hrf2CRDmnPf3qPkaxVPxGMVJnc
ZpZe7NU+Nx8350yM4E89NmnRF3hffNTN1giOylP0RfEg5Es6+kchtnGElbCnYOvo
bHyy3Yb2Vk99JkkNuVJ2E2+5jTTVljS6JLP2UF8xCpwEOfkgNa7t8ULj5RzKtpWQ
tu1hri6VL6DY7mvsfpIEvCYGtgc5mavGvzky2jw+n9PeDCnX4iIP0zd1cSHYh0uR
W+iP0qjp59b/f0Vrpz0gdUUCZU/n/g1xwjmqGzkzcN2c/OE2q0hDuY35bYNb/5ut
nOFYSmuD8AUCZQbqJdGH98yWqCh17EkSy/p1og3wiPerol6Xk1RbEfM1ecyUSJSF
aYCtQhpALetboEEj+e05f5hwBdi3crEJkooDv33axHeroJTYF+t0QUXc7Iyi2Bv+
4BY4RU0qjXfy3j408MTNVPJKH26VZXgyQs3iB222Pu7PS7G5/wttRBapMSmnBSzH
azcdbOogOdDCbMEZWeM9VkbiYs504oTNh07QA5zaule7fg4muFEE1j2Mt9K2VP3u
4OfhFMKRNURqttUlajc9bc8KJTU0DSJYJ9QYMF31LHGyZj/Ks4VgOSh4rJ8nA1Mj
hDoS8A34lx8dAHH1Uz6W+pXJbmjYFaioQXd/JI68xr87OdrchLs5p19QROl/f9Ml
6U0+Rvc6xOghEi8ddvaNCC9xstP7jEgcc+R4CEGEPs9w8WV9diFiIa+bMfrNsubX
azipqMIisr4DBag+VoIT4bzPU4W4FMIj7yyy/39+1ZibPKIXwa2PzI/5tNV95lNG
CMPJwUVDhvcTDLFOPHMVwM6JI18ftF3ahXJTlfFB+n6sHa9tmgR1lOEQeh5B2U3G
wzzewTSVtTydueT9BQCq56vmJ540kKOB4Azk2kpJOK3Mg1lu4lDBNP4OFCFaRyoc
aDCL3uKLoYyWQnI65OPUyT6QRpLbS2dpNXXnZyjsg+yffLHg077NSh21XWKSMGEF
GwMzlDRNqqoAjV1zN72Q74mFs2UWDfitKRhpQosdmJSTSKhC8cWulhp3aSLkUlgf
pSoaoNBkbI1GOZ+8ZAZx0oPXtmy9xAh6yBi2XsWvKTRh52ovrq/JoyzEz0KtpdGU
X1VVoVyCysf0zSjkjdkBTN7Cb6QrUXaIKc770WFQx3tdT7nMcGzODI0muVOQQ+Xn
YKGLfvn8gEkSlAfWEOKBk6f8HC0iuLlvarbOQXtioFelTVySsBuIoicaM4JfqYtN
5O9jgmpHbqk2J2A+2HUx9fcPahB58sQUdF77OxmYHXG99I7JNAVl5HRTycNgIMTH
qqC1PE39yIDvIc+WQE2AQa/VpL996u+TV7+9Xl4RQfrCV6YODXPtSF0K2BiwDsYs
lKXH1SbzKOqPtE6+VzrB7xxjILt3x0xg8QsYu/jLoIXN5y7KqMjsmwse8jO4Lilc
`protect END_PROTECTED
