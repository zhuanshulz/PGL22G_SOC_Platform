`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pL7mvuqzUq/t4aqzw3kdgGZtJSywXQ5FQrquTpvL6FOsu8KLoncdf6Cukqg4YV6b
TOF4uHJzAbwW1O2h2F18fE1ZQscJ8acf6DzfHFomMOGKgSSiil7wHhCW2MIPxOXq
jok+JcYf1bWCxuNp7EFdJQqgv2kb+CLdHXyYdLGK3Z6HO0VAxImuXUrqw2+DcN65
KZoXgMGHgo0asuR7HGEEqy20hE62smOBE216i95gKx4cPymDnIkOgoAJxJSHPLAf
F6VkGmM+gWLkZ+bhEU31jdN4XMkcd1TeUzOpocaKQCmkK2aMjfbf1L+PAkSOp5aB
NBzlwXpl0NwBeyX3HN2TFw3UzIGZ3rcTUhx7uLm3HCqcseIfM6e1iUKxfDRVj6tH
A7S16wemGWvCafZZIRYSDIWIScPKCzdtWZBTCY+vNxQBS36gh2us4IkAwn69B1B6
oL/OWSWb5NWwlF3RXarFMyslYT9E2QhdeRkQI53ekLm7l5hznpj6c3Z7/YPqBvD/
9/xecFa1sbNMCOcs1BDMaPjFDoRbsFgUAOb2/H5rL7+rhNxYJPGLoZrayF1FPAWD
aTgtZAg3xyaBsGsBRHaedy6U92/by9GlnqLPZWAQ9JR/w4wwcOp6RnAEyThk+Vj6
aMGts/aQIN9aaKIT6Sru8n4wR6DK08FnZ7YRgIUzvo98ZjtKx6O+sYO7/EDXAqs7
BYp6vcMlM7GP3k04XPCzIPa/uoS0AEFf8j/MhbFTC3andCAonbG3vylRsL1paO9W
XMFdVfMEpUrwOWmpi3KfyPiJf4Xz/RRFd5sY8ZvhwVCVYnj0G2Ei94hZZOtyJ1+K
7g0QgjoAQqAnkgBWBbgpDirXcnLjoBPxer3KFZvU9heiI3qQOYMXgyeLWONPsAlv
b3LEBQtsBN4+xjKdvb5rMs5Bf5N5IYT7rOvXC7zewJJ2S8JQWKnjmDNfPz2hiA4t
HzOOTd9a8iVki+mfUtRx8T4mtxZ3nZ9JRFeTAximXqdg9X3pg3d/jQP9eBvWB+2g
CsNzVlyIkAxD+bRfE6GfZYfA7HBfpuc88T6MGECX5ofRmpWoKFlWjigt1CJa6vjA
D10org/6nMtbF3t22ao+xxubAdsK21KQvgEWdfo7PMWtZcvQv/6lxEuM2BjaQdMf
LjKkplGkmr8o5NOvV4sKYNIHfJwjT9OEpvvGrYYzVnlAxGalyJjlZP4oG4IEdDtA
RKPVNatoCzfADoO7i/fvTjhfVYl2DgiezGMVBZ6GSK47LfjeBuHOwLVaETZ9GLbF
+SQWBZPcLsESjDWt95eVFvk6oxDK+rSaWXLnNxIkFb1CGcIKXKyNcIPfu9+va2Kw
AFq77HmitCS8fXU6UZTj3OUqFqJ5/BfiVAkLI14d26FW/aEiI7c4T5q4kSOVbCwR
/2AkVShQO3Btar7NSlwXLsdvRjyUdNhdmgx3dBIH1hANlvYpZovR2vZXW+UM+daW
o5MCtqd/CvSORtxeFOQMmWQihSCrpv1Q91SFHP88i7nWbZWvxU1I3nz573X1Ghtv
BPmGGJfacrw63jHuDVgmDEQgfaEDlbXAgllO2yImRiWcg+ZH8RvvOjldaepw/zcY
F3QBis4Z292aIdRATmVgMWckvSaDZsLu3m8a5WJ97SnmRgeUckCU0Lnk4N54bDAL
n7/hm1AwHfmoLrzNnQ2bLL7DbSeQcO+mk0j5MKgDfpHRawlpGMSJYi1ONdO7yqEk
ms5hSWtJQmS4s8BtE46LRI5MMmAnglv6faK3uQdhJDUnDORB3YxClBLJXJxlWRyl
yjyAqVDM0ogY8OKrofiYuiI7O+5Hx05ND8yDa6JjEoqO5+fb2d43wKC1dmD3aqmI
kGE29cK1Q1l/bJ9whYtC67nHIk7VUxKTALxGX+RK1cDtoWNH8730YtSqcWxiOzwu
BTBu/gCaIrIl+teXXvSNihH6tpbQDwZCz7ClC5bBNOdrovf25rQcom0+OG6sy/VE
jy3bTaF6glXSWpQPfmQMS/cDrW5mHoYjzgvhsbdgbbg/dz5KIVClcWebaV2FmDnI
AUXNxeeuk3MP5SFtFJ/NEQTL6qHIo6CNNLgylrjCh8PvoLBnXyJ7ix/YmXTIhGPV
gpxDgqPF6zjfzIS29PcgCM0X60PLfum0SsUW2tEJWcfH/Qp8gQ0dzsrWyxsUmKdp
1JVTssYhLloIkhSCRo5z/RGdVm2PnX675wS4vMJICxDiT7UItoSKrWmLylUs6D0j
36xAvbmj6ozKqWq/BW3CfwPbd6p1GRQepunoCocBdQhN1kI0GoDLxhjeCfLv1tgS
SS8qxO8TVJErnV7G/j+I78Vqpcd7hG4MMKl122nWDhM+Ach/VNxtJPXFyasH0G5R
GVpEz56s6HUudzo3f4Bkox69LTja2K5j4iCYJvNRGLc/qI1kBKjfoArEvpn5qDoz
UZLU/BMUwSWDI7JVHS+N8kdtiNM2Zy0x0kTqSPOFRlIsEDC53wT/j+/u6lnBmYA7
S24vl+Mu/5eM5lUwYT2Fy08LdIk3aYmXJHtQKcwZ6KPGK0d5SneedvMJ4Ro9uFBy
yzJ5kCjCjJczpvjbajdk+Ao4sjraeWeRVGg/17sBR+mLFv9iJhntiT91s5N1zyDh
Hyl3o/pS+ruF3QtW3ZwlHfs+iojts0AWlVxnlyXwmOEdYSYizHC722zyS3TAX7jR
2rhfW3hfKDoBGXb2sEsTrEUI31AqKjpo0kTpOL+7u5MvcPdAkmWQR8acXtS8JsnI
6Wgwyhoe4QLesmZdw/CSnTCahfK0MiyCDXi1X3+IT62VKbPqdk1IbJ3tOxws7L93
TlDB8bddt6QnbihgXXPeVqmC1oo0Hkf/1Y7ntPiPfOyN/MmcbZDGPnYsq4sm4Y/5
dhNofRC+E+rY5e2qK2oaBLpaZN6Lm+k9phn4u6+iYzcDsY7q4UScPbYAhesGm14b
GnJMA+0mLarOcT2h9w7FuXod97+DmhQ3T7QLC6qiQNDtEOgjiDcGxYOE7tT1Cr3m
CsgdhMsqL8JUApA3YGqb8LOfCTVNGkIC1EPjPliDuhhz7f9JY4bvJflhZJcgcl9J
KHrOcDE79+OJ73y6RsjHTbtiBxUmk+PUPU5s+/gBnLwcNXPwTz/hHGhBjqFnYbht
MN5vKXxqGHc+H0sN/qyL5vpMXBkGsmVjVFRWgnsO8XtndGtspn6vOD206VN25PLM
`protect END_PROTECTED
