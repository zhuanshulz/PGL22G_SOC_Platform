`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ZqaYah5Tgw8YmhGZ+lPqHlmtY7jZAii+GZ20NgOY1O6AfWNCkrug+Fi3CJIbeUt
XnwgrbdpJAj7MiQQ35JPFGfq9YtZPStaX1k5Ue+CeawNdheGiqJL9mUBiqEBdcsv
t+pszcuBZTvY8p9yvkLn+FOd5yKRaxsCPjhFnIYsK3iSnYR2dCJ92jAilCKa1IIL
xCV3iQDv5X6RuEFaYMkCSQJybLI34pJP13IyPNzkbz6kA+7wY9fdZSfsqKCvzkUT
zwD8wiItBRAWItiPFJTbI+8QujsCWWumeOBCR7LxkWSsXjzRJypib0NnGNp2S3IB
nrRSsfZCGhbVDWhjHzT4jd752mL7HsmEUN689QTnHm8CCS+4tGMMO1T9kIEFEquR
OqK5xDAdpHrRXxZKOE0K7/rZs7REmheeG0aw8L7J3Qlyj6pq1kLKUertCOhrJ0Q8
hC4K0UryTy6gph8jWbZDIPLeWwNMduSJ+JIc+J9FQPd/HuYBUtNDnVKkY1oeWSzs
JVb7FzMDt5DeM5qNKqMXGxyzjLY4HZMtUPkfmzfFfApr/HYbxW8Sfw3zjL5g+gDI
GA0SCfAAMQa01b1efRZsrVBmkUApWuQ5wEKF7CQCWAwDRfqfP7QJwXjBx7eihG14
hOhe+lyoOfjZfrrDuFXS3YMvoWFhi+RLVbuQp9WBdJUbSxq1jd0uRY+OvHoYV5yC
ANyJ1+vdyjSP8DeqMnLKYnDFq8TCMdFOF23ymWVGsq4=
`protect END_PROTECTED
