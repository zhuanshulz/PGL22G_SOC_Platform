`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/P6FfnbuNKGvMXDszVU/ytu9RpZAb4n8RqSU27nShEh3peXOdCJ84hDOzFk+MqOu
VFiaMVk7Bz+OfYPkK3YEKdfrTSKiEIIOJGaGom1MMUZyu8/rg9CbwDshXi9dbCl3
eJzA0mKO3A0zH4X56GwOTKlWbfwSinWjNZzdOYaSOBdA7Ux3zjgeLyX7eaayNlLs
TC8DVAAqfpmp0YarOoy4Q0NFOxHlFVtnnbQSo+u2ff8ZnU+IoOqBMfdOrP9paW62
kHF0El7HQNTLF6ztaEQ8h8U31xSUe247eocdMeHNahRat15Y5Enw6CoTta6q2P01
94iKw63ARgofRx/dFXB4rW5DVq3ModB58hoWIN/Ql1e1AIHr8YPEnD8vQM161vNd
fIv3u0tS1S6Ef+2WwcPeQidFbtp/Oggv2ej/10TqkEOPcXmindcE1YOcQMbOdWfS
OfXwRYsBDq1IAcgeLMapOf7Y4NsHQTezzkiLb3wTFafPeUuorgtI6k4bx2v+2Qex
Tp3JHgXFs9SmH3uZIWtxTAHFkWZVZyqpMXcLfCeZAMWQTDa+32TvNoO12anXn6s+
N7qFhJxqOTTPnuG9gTDiZ3L+qqRLoZYtoaTsFwq0miinP9TZ5W2MaRENv/FSqM2A
j9LN/w3EJiDOh7MDBW9r2iBSgbT7+lonty4LqqY50zWIBwZmrBhanYJsrJ4tHA0k
VRM5RYvYVYPxH+FWG52R0z1PydaQQNU6QoM8vRNpE/VX4X65pEY3v89tB16p1sMb
2ABdIrLEfqABMRzzv9PLIdJAsqnJvVryURoRDOaXE5+uh3/xToCBz9JW2pXCulOf
bV6IWkGwNdhbpkOrIpa3cSolgeIld4ZbHH1aItvJ+zXhxlQkCd9BBQCJYxX+b7DA
YqwAnKSfRvog+KCtzce53Dw97aYK8MKsPx2ALP3DqfymRS3iBBaGybkAI5627oUX
7+2Iy83P3HylqGiRY7Do6+eIx5hwRFk5Wh+BIFDV5SkNpEHoZlr8FQaGCStSdJP2
DNRUAvc+DPfKA3rOXwLydwUUSPqt25C7VY/Kjaalxvg7dD+/q91V+KrSQa2MBtMg
x9Z0pRSfT1BqXW8kbTApfI94SDoMg8ADow49nYzki282toq2+C6ECOIG5F3NonR4
Wr3mQqwgUUyFHuWehVKMnt93Z1LBeTz8x87Pl9ohfX1ZGpojIvmVlKevTeVc5cgX
0NP78DTHTrq8/7jdrsUys+kaFpv+3fFo8XaNOyAHMr8zJQrj63GGg5LOKmG5FA0d
diVxvhADEOdc8PokKDIrtkmd6p4mVya05ppbVMVne27ygCeQdPl2HJq+NUjW0fSq
WvTt2pSldEjvnJSbQL/O0zuuI65cedf7TSqP4eanL4ncQtYypwGOH4TOnl4CaFAk
tgXdcoKQBkwfVIhe+jqIiOId9q8Yyrodzrl/V23l9CJj5whX7nZcohnNkiNzDeUq
wqGv+ZwMhmmz6TGgAeL28Y5oTzd4EJBIDuk0V2HHOhiMhQSAN/69vvhyJMA41mCa
ckbvxLtFRLP/mxzw2IHU6T7G/7sykF4VUKufUETuzhNz/0VpxaZ8vGtJ6xPrhDYP
dSoiQOIw2iBLVnYbXkyuyk/xeG/oThg409O4IZ4CddULehHVe2FiSDyd5gP3SSQm
7mXdUVCnA2hxC7R2vgmBgXb7P7v0UhGYioB08bg2ogCOlDDUAM1BwYacxrVwZk0r
ABaomQ1k58Po3nBknFWaaLITXOh4vtrekaGVT0b4lua16lt2i4gGU87hRQb+JAWl
bTMTZUc2YR9Fcvl13c+Dld0IobbWtS5/slNHiWx3FtI25kKxphVXPrByXq8O2xB/
fEiDR9GTXuCSdRAePU4ZF3kUH0RM7ecB8LMuyAxQ48wdYkFSi6acPduUaqxTjn2b
XUGK6TuJodHfV7u6K0iCrKbO57e/l1RjgWFB+DLW9RsdGZLRVMfgm5/DXYOAQ0NK
L0430cn9XcrUgGdJheBDF+e9rvJhsXl6VVayJvC6aQHgaax9WnzAgUUGnl7mdg41
dpKzKM/1sz6jinROn/vgIfNHXRAEMoBTqyTmHQGgIeH4EQFR71SiEVFDzQuX7VI/
NYByzhdvFgYH7YuXiSRGG4AIPW5BanInUJ1y/6eYiywGPW6PCG7FBBo/hgnE5GW+
NhHGRxbhOU44flnyd4UgkvSsajkjXry8KtDHpzGsP7nfwJjyoPOdOoNWcW7+Jz2i
s3lG5Sb71s3D/y1f1LsLuyfdbgbKiqq+c1OK8R933nAUQGIPHA6mAoz+dhi+UYF0
bPLrUE3OoKLrOX4oeWImQLYRIFP9y0TdQzCW5RKYQT2OBVGGhQiH3utQBfM9WPEi
QUIf84S6mlrxT6B0n7TV+3hETkGqeZXziJFhFSj1MSVyfikIXPof6uGMkSBdT6P5
j/2IVdZ7ghW7J5WghVmzYMhZUKEZQxsKX+vQTjqlBn1fH42CrYk6brc4r9Zsxz1z
/sCOwDW32bTzEZTK9T1CmjgQg27dRbPl1Xko+hxb81PEzKzxNu5SnaG60jzdeH4l
Mr2Io3mTLcFkRtpUF9EBdaKugVHk7idEomjvr+HiXRWTkmLeoqN/+JtnBYhibLHY
Yj6xn6VmOblKW/VziVaDPC+GPt+1b/Sh9bU2xD7pWEJ6nMPUwVDZlmyCQOGefB/C
MeLi3z2Apo6C8puh1mT9HwzLdGcZisGho7Tg8QNvTXbfixmIdEx+okWm0krQAgVc
Rnbikf0+g2bn1B5hfueYRHr0Ny1qeKCUv6/ZLa+yhmsVWx5ezKRm54H4/Xd4awzw
Xd69NDvYn4gNPKfFHEp1XIFhp0KVBWbFUVRuUpFmVPa4fOeodH6Noae+5QsVYPN1
P8BFAGHUUpxsDzFcp9wmIzxhTty8Vcj3o7RBbpFzrm/72NGHkFBF5Lxwmwonczfl
q+WCJVb5H2z3tzq83hDzcpaoGbUQRnV8Ux1PUj70wdGLVjBk05YaSPnixKq3SENb
wqKcNINNQR71TOC+UiJbfqu0qOfDV/K6CTkDjw4Ri5KbobIfubfbhypjQnVo+iPj
HZQhwVVBPTXrYR1HpqB7OY8+N+jHOa6HLZEYn7gZf0MQVOkiRe/0BQkQkzAbsayO
r26RCM8ClseLpLCEc4HF3SGnymndjuDAiuhcYqUyCvdS3vqhCOGPNlQ7LmGp6tny
AEbwVS3Z7ff1mu2FgELhbuf5YFJWysqvdUObbcPfFP0nxtneXlCFiiSZcI9g2gZH
`protect END_PROTECTED
