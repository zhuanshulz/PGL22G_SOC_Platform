`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFNaUxnrV94AK1jH+Oefmm0/HzJaXaotE1DkB4VWNUcmHOxt6fDR2eK/SlgdGtqs
+0Q7SpBG69cGawhINlTKEBPDP5a8DlM8oR8BGHX9tXwHCugiuQTUmlDinXvzDLcx
qSQxugVFXvtb4f7XNES9tWa0wtv0oNtCE25QiyZjWK0YjcCpc4Tm+mVlazoDcY7Q
YVdznHBRhkzdeunHH6JfiLOmFmftOjqng7a0344f5MGG7Dpesmg4jXikQroY9hud
aWdqzoYKNQoNDZpC4B+bBb79iiW9W63FQFrVFGxUQYWJOZNRiy/RXYb57aYhZ/bn
P2BhgDcrnuhY6GmK0GQzOQNutBg0o3sb8tkqm9VUJHCyRwWFW8UEbiVDJ8UJZWF/
4v2xwaEJfvGt5AjxzVOuRdNbPmNlji8uYmERk2cTOU0Br4qZYIwpPzez6AHDK4n/
y4x+6bg8UGoedbLDrkhbOyJGaC0SA2H1tmNEgdbQfHWHEaYf4/5JvODWw49L+Q4V
hvEWeDAV/6Yu/o0nkPbQ3GMFeCTn4KQTCaXiSUJR3mW3YWE9UQQ306b7qFFN/j/W
OMDaoG3lrG7oytupjNms8n6L0d8EQdSA287y4b7e3/s1HFGf0LCnuRIy2866FuE8
VnzbceprcNusOvf4Be3hODfzs5HrXfT212Bc4hqDLkfUVWQ9Qo4cDDO4QYnxfR2X
7rkpfVWjswrkJAHivqyaZBFFRoQOj8z9GpaJV+HXEP1p+F/BFWnPuWGEied3cSt1
7qOJtAeop4g291duSor8uob8j7uqtfXDRo5mNLHXrM7LijlZUjSi5MwdCd7AG4CC
KIRHelAL5Fv677blpf/KY5QEktsHUCDf2uhhS9fZ3nzf/QZKmOBmOTe68Ea/21Wo
`protect END_PROTECTED
