`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PpJ5m11jXGxBVv1DJc0TNjK7l+HOMlefYNiJ2qPsBC99WiuyF2oizjuPpnXBxC2
pwCuHo/gga/qRGVCyuMCSJp6gP+eqhUyfbelnEVfoJKkohAVfXOvounwoD9D6Fne
U2OdQCsLXpbVoqlPX5PHq2KlOSrJCna9RAOYKsyPd8q/gk5aIrpC6I8xJ2+xAx+c
4nn2pdOEKPiXrGSSOfQnccoK2tiQccP8fmaN0S5dOlUItkQqieV5Yz6CV2GqtBZI
vz2GWHFlyn1NadiguTs0ewdTsh7Xg/5Hy7xShL9hbvq8eY/IV9j6xbfQD9r9CUPf
iLDv9xdTG0zioPXS9X25nfMZHrJs/6v4bCP2/miWC5fybNbAb0sd0Jq1TJvzuxLW
XA1LcNGajnkHwPnq+6TfmOCBETlriOX5Tb5Qwy4j2wTh2y5OmxhFreNURqFWvLih
8f06mMdUUEh8ekoDKEEpTVtcGVd91k4fd35u2VXpS/ctlhyiNr7NX1UU0J0twGQH
BxB4LBvR3I9rO1plSLE37OdksdKuyf7Pq/uFXsCmomqE7zwUASbtBZxDEyyRgM8P
LhoZPnB+YUXgBF3QdDDTMQX8H63FTyH0WDxHrm+5/kuIkhAq8dbgDYEwmje6JYsF
LecQxq7dBYz6M8i02k87DIkquVlYDnK51f6bv84LEoEXk/H9fj0hMja4oO9r/gk/
8TK9GZ9kT+e69jK2FgCHB4v6jfQ9TQ0nCnFAURX5YvGEc+gk7ILLybqWTK8s1wyP
Y/DChefE9QO86DIEBL3+FdseD/HsLO56AUwriyR8Q0QPsU4vVKaGa70PrGyf2zAd
oPZ3LZtKRvlsEL4GkY5OlZzNAa1BcqvmLFXwqMaU3iG0iYVXHfKlRIfhxH79kYG8
w4F3eZc7mT9icLlTl50movphQtcaFrtwSsjDITkncC/WZwGPdUUH9Q3CD3dYv+gL
bUDDuiayCoXXX/ujauPbMuuDq0ZIHYH6HMNoewgbQ5HKbreotZfh3P5zk/FI7mtD
g9U8BuS/r/0cHQTllJtBzQNcdPEe82sBEKED4WGYlvLoqriZvAu6XpC40GXmA2BF
/fc5oO4btW73eSqnEiiQ+HQ91gl9gjeERr4omyi5iZ2M2T+Ya0GMStor2n5PRYbS
wmkmnHyEOw5x3rElphYCnDG+AOGAeo/BINISNvwSFUX7nP+qddfMFHJv2E1MW+uH
HbKkTLlheOAQv6mRla5X17TB49hahJ92Pk/Nv9relakqhk4+A+SCS+zLGinGVECg
s9ivWKjekqWftLZ0b2JcuA3DjoWXiOIIMHhU1OAZAGpXbIGIU7VYmnV62/RC+iB4
DloJtrQ4ouDOLp9v+J7I6HINE04mECzzS9cgX3EKUuJ91OcROU4iLlBjFvL2gZA/
tlSGN6riItvc2Q6lNzLUEt2uXQkjTamyvWNKDZVt7P8oxgWO3Xz7PsfUJcoNLArO
05q4ixoTyGcjjJHaqDEIDmHF51hC1iDs75AlL+nLoUGJf4IvBnfYrQFasNcqq4LP
G6OwQn+m4slsWWXYZcv1BMhzMXHmA1x9pdWJ12oNQnWnpUzjKa9YdyD8YHGXMbpk
B8wjTT7k3wmN+r1r2ePHIQcXAE9eXUdcXXRwX+cbMc9d7vyj6MhSpPVQ9n/VurWv
o5WgPcVBqFUw/G8OHSttbR8UoVv8aqYNW9GUMLi4KL/OGvnM7TV3WHkaA5H0gtMV
6ozElvopokAyE0wEjCAuZZ6TisE6oLYtibAgkXTTc3G3Ogp0S2FUcN+tNSsgrA1x
709Wk8904UygFaIk9yRlW5qiO9eLdSHtfgCygc1pNBu2vuiUxLNUy00+f5Ak/Vc+
E4j2GBu8wsLfRX81lOMHuwprE9CRGHhmHzeU5ohU9mL9YQZyJ1ar15+6jhNBZR0m
m43Vlc7SJCSzHg4XR8zD2ekoEdMstJ2O6HV57DCw1gDAi4/WKg8h1H3W3HfFB3me
Hk6NUhAiX0PSW1uTnoZ91uVhnM9f5yXkNiAL/qk23ZxZgLI128YSaAjb4BJsnbsB
IjKNw41UWnHi5pPmEMPgfY4CGW2OW8PmbdwXm1TllOZuwg1NjRKmWdGihr6U5oDN
efakINX8bUdreULq3vgCludI7t5hIoRncIoeJZ9Z7JTCJPIIFZlLj/Bo7X59+JwC
AN2P/WY5f/J6muZgQyYzG8QUaruw87LvkgD3qKd3nkbdvT7WXrgtVL/1ToATwYpc
x56po2xK3d1wfAY8P2N1aLzzAwDfNy/AYB0+8OBXtI+iil/c29a0/Pb0qgIfsLlx
2k2bBefO/KncKzCb3oO0lcdJ4ttdvXsjdKVEur5Jexn6evSItnU1n78HO9CCE3b4
jS+O9DGYM+FokFfrcAfeBeIAT8zk1ux4UBWC3L8ACLvOlD53bfXzdaZzwASbYrfS
HcigXxzIphwX3agmKkiwzwn1RnWM29P2ImumnW5fCqk5mNXMfIcZxRMN2C2UG44R
hqtYj2/NU3msNdcmaBeHNNHQ5Y0E+rsf5hfR6Y0i3o6YOf1WwZDVvpeUxvVVbZuy
44DdrzVU1ika/wkLJKyGJztaOInEhScBpt0hQ1YA7OGA7WAQmRyjwznghP/yr5/P
Tt0Ej90RvS1Xv3wEuDQpRiqQbc07ZiIx7QtHF1/3OKMSAS6N0tfCJm9XhGYFLN2R
U4xQqPO8mfwaVRkutozX++yE4sT9I8P1rcH76afj/Cmx1WjD90b1K7VUJ31/pVsA
EgRjNNjOWf8yrakS55NvmwsgkrjcvRjNtwyPpY1AXlaRYwl7kdbd0HMxh0pGLJbS
IRJjlo8Yj/SM6hRMdGYvAbmW25nTfYSHubKjudx/3HfFyJYiAmnXz8y6iBiIuH/y
dF9Di1r/eI0IV2IGbmsOURGvrISl/3prXjOP/dYSOUHcIuy6CFP18/S8i7FBMZdt
Grk9FNIcCahsNdcNlUjWg4/RA7gMc044GHiYCpjqUEIRD9vTpIG9g2vqRKT32yeX
sjBzHHMxziP6sRKcyQa73oDRGRWXaU6Mk3FX33J83tMXzJdhoRjiWuNnR0F5WN0g
LL9JwfB6h7jM/heLiGZytGkV9R5L9SEmo1Pz2rPxYnKnU6j4HZw7By/pAQ0ECjFM
2G2ROfSN86WBRtTB+eosd4cC3MGNdk1MQ5bErWV7FpP5fGLqeGj1wjrXMRMqW/xu
RliqC/UedwuzM632K9pTjFGKOQQgw8h0zgj4+h8ErERz07Nx9rxetx68On2zljDo
FBRpqrk5hD8B4PcA99d/Aof7tRRc9BZdfATrs7WF13Q=
`protect END_PROTECTED
