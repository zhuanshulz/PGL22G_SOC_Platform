`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6pTfGdR3uwnDByZVJ767yonIW4BsflpnwTdAUFLgKLUnBvodIlusKiZk/6PdVRxA
UHE/kF9x+9JJ72hewQYdMGt2omZPsmvTaLV2+MCQcvyT0uN7p2v61gpR8GOZ8XcJ
sAZrj92KhPd9Qlv9M79UYtyJBWwe34sdIsMtukQ0I/yGQAMacSWFM3bAdpyDUN85
9IYuDGeyWxBjfhy961jVZQYJ4QgNN1TwKk/PkOquRWnrT5BAM+A0N/gqlHaKhJHU
Zof+190bwjFcwu6XIo5JkOVpW/AA6CpEeJgiDJRRPBM4DLQM2vl2/IDfXxLAIkCj
M6Ldfet7lRQtlYv2neLYXRNsMxCsYNxiybCcr2bTS0aE+h8IFv8hoPWrdjzoSJEO
rCk9KcM71KBH3+s9RXkauJlze1jloDiTmiUTnSQHpmugTpIZBY/AzWdwBelQpBh+
nfikRcUWoykQi3KI7KhDBZs3fKX7xKKzCuzH3yMj4cTg/Ya4cu/fSJcYT6E4/ekR
OYyTRS7cDO/z8d3K0A+hqvXt3h1m3l/i5L47vBfmmTYkrlNY9WQqrtXK6Sg773TY
x5nxCOTpBGeL+BJY1ySznmx7JUS7OwsyP6jDcCq3nsvZKgOmEIZQju/0widSBVoT
bZUinoR5WgVwjs53ac3H605gybzP0gR+/5h+xiNtWwfuEpNNkhXlspuAgdVBhNNp
tDC9cZCZNF1pHTj3NWWyETcnuzrkLaJKSErg8/oq2dx2nRxVZoXIkjMUlaNXitxC
SyKVCIkIQMSYH7MNUE6w+zg6yLgesXW4vG9O2baahRydY0NH7deL13VpO5l1df57
p69HbnImZ+5DVb0z8dwuviJmlVtYKdB0AwhMh9WvUtKAG2yqfJWVzLnC1cWPwqg8
/xvA3TKRLubIFhVy864m/5x1SeGL2rDWBy3MpUhAGeY5RWIZWHy4QV2/gwL5tv2y
VTS+mfxTBvUuL00Pi6DLaxV9uTT8GP2xRau9aTQQlvQpQOf01By8BjCNXT2w677S
e5L6knhpMrJ2wADeMUiP1ZsYvBmxjHQr6KB6Qc4xIyocXpfdLraEErDWqtjuu2+C
1AaY7lRGxXZrEHsfZRkvjC5G8SkRFH/m0mj7G+A9wwZ93lmFMHaS9xdbAEQmCjt8
zx32Qc3QbTOib9+OFmIDoO/t/vZ9ZPD7zCRC2Cm64JlFsFjb9KhijFgFHsbYmcsQ
1LGW3Fd3LhOhi2qIAhOFh/hlaBNvyZraNWfFrNOuIh9KMVBDF4p7THgIw5a7fOUq
4qfX0qmpPnVwkDgc0eobV3QYwPNEXZ9T4gGSOAweoFTTI1vngpQJHhXl3LUNdxDL
4I3bOqDxyvsutc3VtlwnKQ==
`protect END_PROTECTED
