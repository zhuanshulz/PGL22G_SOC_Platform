`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ly5apFL/PSHzNFviFph2o/MBOPnmbX4ml8JRCsAA3Xy6Mh5oFC+94hWNu10FQMnV
8deaiUBhfu5YfwS9T1sAJjRii5cvtA79M7k4pTxbYtRoqrIpQmnKCSig+2HXzRIp
QXBY7oAVeLT7RYG60c3BMkZtL/+kO5ysYpRz9AKY4L2L3B+3Wzt89JbZg69RMYcG
q6BvsOB39THSpKw7pqtvn+S7SRZlH6Z+duHY1Nu3OKIWfX52oOCEa6Jm7aWJAan6
h0OKjCoKFVSSi+NtLpbdkerjIkxcRzsreeHgzIqCZzvGhIQ0/U1EN3I/kjFbzkPy
dNAMrPaCJ+x4ykYW76P443xi/DywkvElfBn67VHto7d9NRcSuZRQVxKG//aJeuBc
nbW9nlb3mvP+Klc3YKeYB4uNhU0kYyJztuMHIu6Zk28G0omMZIXJTadm+fNiTLor
REFrYEdpd3AT04p5GQ8EeUuMnpDyDKD5dTZczsptiP6ZwAkdmF++r3RLMp+POpRc
/1XuYi+s2pQX7fr/QIS0VbwBs4Wr34MyYT9VyUTLGP3NBCZCrsYntff8j4R+Cu/n
npZXPkYaMShj4XwdI8RLOv2bCjeXVainUgKytAgF8ho6yNtiGskWW2uI30aGl2bZ
Hp5KWUMyGA0555InyIdDVMjw9P+0vLWP/pGLv5Yv/msGfhSZ6HS0k2Mf+h8OzzKQ
eUYCdD22Mr1T4x0XJ1fnks89Oi7zx5SLh1s+bVRWjbNeB70jsPUAkbzXn/SuILB2
Y2EvMNcMSsGxUgWrw+8i3ABr7uSEN/Fvlcc650bMkT7qW076mDgL5woKNibkPtw4
XPhjE4e/RECLISXYYzkt4oemiv8Te3Hl8qsE1D2D3AOKWenkuPRDq6TobMT0KeOb
TWXzwTv5MH5KR/WmJWMekW+e25zgidfZ5JZNakLoxSbs0PtLDFEEJCR9UzxDq923
jILaGst48Tsp0K0wJjUcZLRsNjmVWruxwoAHn1B0qNhQ9oVm2Kjc+tinEroFVP/M
axhfcKX83+gMOgs5ADzonEiMlrhfk0hv178y9O74BIEOEViz2Tcqy6tq6T8BnqIt
kBHl0fIr+5dNGEs5/00CdMHo+9kEmZtHhf0230MWG+71xHL3dqIh+H0hQsj4y3sJ
dNmXwLUlF8q1oEfquDOVu5K321QMZ4cNkvpgyDgfCUoJOuLpRZCeptzDMIRpubf6
GmIrnW49IFCYHNU3m1EgWI0+mJtEM7ICLTsLwkPDDZsHfAoL/F86qPcVaraIC6E1
yuVTMcKCUcp77+VxFi1MijU+utkalbUoLh5xpZUQQVQxDcipMZHFYvLT+KBgm0D2
PIO2TdYVV2B2USihSGRq+FfxWS1xCgnkeJsfPrq2nsWJozMOcjxSewzvxdc8BLcG
CEO+6Ox+6Jkl8Mp/1/nB8Kixz9zlzIJVa4kgFNsI+2HL8l2MC/T3rvUrYT0i8RaV
/uagYG+x6v275YEPXZ1y8pj+yAsS5hQBZshWlV4jDffU5jW0ioafKiokelsH2IGp
SHCk+6PzEOsp0msCG7YE8csJlb0soZXl8ra4mIeqb9o2uTg34oDzHWRIShRBceEp
SZIgnQniHznP3RhuPcBlbJdybiP5tUyhgLppuzyaQAfK1fDLs0NZWb8KV8kpMqr4
RejCI5z0AMPxSpxzZ3X+KmXOa3wFiQB8JvQSfSySdX5VRRWfrns21ymmwzcNVKyT
Tz3NNdXLMy0Ddlne3ZPUL8LnBdGjgeFc3Tv5QpG7CRMjyKaFDHo2cB9nrhO9GdY8
sbOVKN5Yng64LNWdAflB2VKAiYCgYh4Bf5CHGRoYYVaYWQwhRASeChmuatbxrapU
OSBjead7q6ue8M/qksi/uoLWZugeCBJhkTUyIC3S+ljW14ekzA9IffH76YHbiHH5
AGDoB31Gl3ZkKyr4cGPy4DrH7to5C9FrT2zOQH03fNh25mmWKT3AcVqASSbuCrK2
BaSKhzQt9W5XlWDTTuEw6eS89nFBKnpX2uXUkDg+MLCz1sR+XDVFbcP5y1sKkhcR
hLmShM5jLHUGO5+nViOvOPbfC2I8Qq0ki50WaRWr6pb2FN/KkFVjDMju2l8PmZBT
kGXPk9XOqHArxRIZro4BI8ctdfS7RW05ScmRXDtuwe79mY6UDpzSyuSiGxsY4iRt
CUuUzbXRdqs7gfeH6RxedpLZ/AIRPOuSjlb4iRidoPImt19AZLCumaraU99CASaQ
kPIfIXuSvrU4lU7/L0nPJaYkVxY3M5r71m8t4A1asfZdwX5jGjeDfD37zudFNmZv
4hIeeK9n0bfI8gll1bu/3SQK/gWizvi1yBA1vR68CCcbZiTBXN8Z031MCv9Ydb7/
tIfeoIY8b/U7hojd0upHbtRzujtriLiSXORfoclQciwjXwOYzrxBWCCLsQ2PnHub
uNPvkInBLGoL4f+JEe+uElUBgNXK/DX6ru5SZsPgL1p9nKQCCvEYKQr7ZjElJjlV
vTV110/0l6qxpz7pWO1zwcV72/uK0mj9U0I7W/QFjo8Sc46d8UthVXZh/C0zhv4F
Eqv0+Er0SoeZVZR0/+HYv2FfAmmYgss88iJMJMSRFYb9CdEOzkZ9KlaQ2joODyWP
PjdRQpjkoVNRXmqw3aPP2MQFgdq2OitLZ//3gc47Lyy3l17x6jWXkR+X5mnBijvv
fR4UAK+kVj9tcG5MUSpsELnbcQy/BaCDYinRKFfPL/5hssRfEc3YpXKLPtRXD4ny
uCXV1VC8mJuD+qiZLWPpRZ+QjUMKjQ0WemGsyBJP0M/dgagtsXtZvJMbGUBziLC/
IwUMYwLM7N7MZmQUBcamRh/6R+YY6vwRV/bpjexAEyV7ihMcur1oEosdQQiGbuTh
2J/mV8wzv83hTYyBROg/tAvZAmX/RI70PXUXIdCPvKJTTTGV8f5q8h+QrwC8jBTL
gdQ1RFSfX3Tkuue0iRRRlCfGnfZdykLA8wFG9DquYh5PD+8v5+ubAUXZPtswDF3W
foNsa5AiAvt7Q7ZSpuXdSAwJjcY5u4QuG3mZT/0DHDE41cEo5GHRJghxPY5Au9GZ
ahfnqV16mHKa1ZciBaQ0h/7zZtseHubgKy5hmmQXCB7GpMypYqJX6PtrKVJX19km
9xcx5up2pUCf7FjWf/1hKTksc7P1QAb1HHKcz46vnZ0u9ChyVXUYGuNE/YKySdO2
C5/FErFviE+Chh68wAcuJKfOXGGp1iWC3i8VAGMNxzzcJWRCaXBr2KZqJXlPJhYR
ZbCyhCdnBABj2VmbXwJD6c09xRBfZChkbvgKuG9exLA1omfWcqEr0Ju9KYhRivOS
qkoBzNHT6/TLuM2r8fqmpn14+tpNgxTtA21l2s9kjXWSYtaSASSU4dYTKfpqmFW0
souxpQ7ESWGcNFeJLtuEFVXk6wi2E0/F2xTXqPyeeEf0w3kHsydfCnc4Dhnrht5K
XtIC1F29PrKjBLIx7A64PefH8agSshTolJubc5nntDoMUjwxaO0+kgH7wfOTgCgE
CYp4c7y7A5d2nVrPVVZced+oEFO9IGkopTwA9j+W1+DEDFNPSpo7tzoGMksW/tAZ
RRtrTfJxnrhs5UouB3P+MM831m828xIybsyVgIOGbBESWxpMSHECV0dAIM0/iSW2
r3BN7BG9RlefPxYkPaU7Wn+kMWPGnD1FQp2gpLrcRRRWtKTvCfpExRwboYfEyI0h
sLqYAzHoiok9hMqAmdjHTV5Z634J6yf9Xtwidc/v/y5DZR3R+ht5vcpqtI9/maEI
gpJ4CY3s1fm1AYL4fWF39oVuAgEQxTYzUcz7NgnwX++FrhlRmQ9ga7ptMy+EgghI
5A9wruBt6WJFqEDHzGNx2Ze/UUUD62V+OFpDfExLd9WcheFUWasptrJCx/TLpINI
DNVVVu2IazAQ4nwbgzhJRWnCrkqTwcA1nTgIwT/b05mN7dL3vnYSJPtO4jVuEfOP
LeEmMJVcr94FjL4thPb+8KBx6r9SehyPrUB8GLIjyJ7MCXfOLdjVwnnJE1opF07C
pfGi/ZobK+fAYDa2kalNRpvn2Gvqmp2JsEspJCmrmaKYLxF1KSQVjPAMKuAfyCzn
ylkRcSG7RPSF7ITvWsCD0r1RIRgzkC8AiEnf5Cr7R1d9IEnZb302IIitvDi/Bhip
5mgOZT6tE1JDgrnMRpkTOYAUpz+uBUYmIIvMeobSODzJXb3hYH50VqjOFSgruoDD
8OGmrhsYVSVjYfw8reD6bVnJYR+wq5sgkMtEprek7hClmIMyhhULmgdPEzMZ5CEw
nkfN0Xx/8XlpJLYzwf1IwI5hiRzPsuTIL3kjMcBbZ4uiprFLUFkzpwDl38XQJAF5
753U8yv4OAucQSimwH81E1Uv9oRgY4ujBrDUj2G5mQbDb/mheBIOpyZh8qzD5rc5
4klBXR81RSXnqKG1sBCnc7KaoRtXQGaL6xEsaztKuK87HuQHuuBOx5H2464DSL+e
RaOE0jJ+qvPkq2JQfNBC2qV+WDbaAeeaa5cmgODFeiUx15wmiiDokh7osfce7+8h
x7rVQPBgbbJt+cESJ6mY9EwjqQ/ZSb6qdR87bUCdpE20aPfmZGIodPNo+wxUCBzJ
j5GFN5k9g7+7veXCSSsB0/QL0DdrljDCJhV5F/z3ezyYwaHUYz1ogMDY3HPNm86S
JPZju1aU5HIs9GsFONTh+o/0fL/OPbyGRP/tXTSYKkPuF3RewrB+uf+AbkAPJ8u4
TzK+dueFHevVZ4IsUa/I9SRO82l4WSdyYvIG223fFYXp4q8xS0eEK5aUGT2Yuj/p
qhLSMxOvJTo8Oh5z1Pp1fMzosdnHSe/u7Q6qTY/QbOjJllPAF3uxZsiTtUjRt2sd
Kv2PKbvXQmCI3bx+jjRUOa/M0gRabQ7h7QkzV5fnIibdlcvRSGIrNAmUo1p3UWSb
5/nN7vP0lh718uS6zTCFP5rbrjy9JJzbHWugGHi2KX+UBmc2trpQlcPMfbfsiLI8
20OuJwUoL2iu7EB5ooBIiSU2JcEqFCykOSxVv9eFLE15om3zYyD205lFje1/flDC
HYxAWJvPSO+VO3UGfl/ParergKomh4LnqQdLx2UHD/XBPqjSUQfiLI68RvdYoAv5
IhZdeOCYIxw50T2vmpfCSk0EFixlXWP6QZWGgnVpo9PS5Jy9NKUwdK7cZsjZVENp
S+5Vcro8Mg/qhCpvCG6RaL04Rv7SUrv67In1/nIL3IuDGBjN78dQR9khevDDs6Nz
GwwIVN+IywgdFr5YZrv3wjuptZPwTJrdn678NsyLgyZ0ruypD1D5nOaulN4Go7gS
ZsfNkUEaiDLPlLYzYfFqTerIQ8675l5PkTrOeJsaFCMT3cT8vh0chwopmaVIAdLI
Es4Fx0bRyZ6ChXeThbt8wLKxHlzCw6gli+tGXjOmOsBQu2Zkxm97WkbqdsSw73cY
5Ea6xkvZhZ8w8eXoEdfnANeaqeOpXQIMikVdEwZTw4S7rHJGss+gJzFSw1OHJFYR
sE2+PIGJgJuKIMK9h5X6WndpAWF9pglPmMZXkJaOPeSyj6DfCweVhZUriAOaXg9P
W+lNfSZrgHjDPtjqn3LYRr19PiNK0I8NXgzWZJyvtgTk6AZcn92f3siq4xRwROe9
+QpuUH3Mz2eTouMiida9WxW4dSCtMfrMk9LPTR4X67SbkImsGUZ+04mSUkGJzoWe
otiqgXyPQ1cCLH42QeDfiaOb8eC6cpzEwK9VvUq77HTHBHMHuWM61k2f9/Hp4grQ
WB9hvxP38PUpnxXwIUgitM22ortXnocIhSjNg/wgZc7Pw1sIvu7TGdsydEUS4E0T
7PbCaNGzmIJZWyLoGE2OREuAvRT2+gBjgx65am6jGbOMd6QEfRsliUi338+y7CEN
E+8GNGYgXT6fL2YOFOUZM+EzO+uRaHPEv4z69TdUmMHeJIM9sdu+dgIgOdaZupIf
qUAQsCmhh2lPzbHIBzD+byH+GBkf114pauozZwRQQZHxjBhqpD8ZDQH/NVJhPEuz
NA+q2hhyw7ZDGHvrldFg6DH4eiOXdXbdwHGNp5VCrbwvu8toJKK4i1y7N2xa7EDM
cvdSogaJHVvLR7Hp+YMZMMptIV7eOynsayIvet8B9v11L3NUOUx9DKA6/iQCZXny
diZldtv7zKxpC3fcIH1ecN+l2y1kChhs36ySE9eiNBd59ovzGCu9yh1o8b/q1mj+
QBqx87pSTb9VA31eaQGW6BeDt8NIHbxRtIWgRB49WgARwkZI+rle4vJbIzAH5eSq
6Gx/uzAfD/xZWHG/npyDoYKQwMIGqFeNn+Kfj9AsDqlZ3Z10J9G3Dec3av+z8Xy+
gbiic7eWXMr74MkV9Uvz7G7dS3AVcMPTJEi5ZbSVk1lo9dxQIHtzwRdL35gTHYAV
b8Yg7LR3XArN14xgNoTznzxIR/tyogBGZa7k8ghP6Rb8NBa8b2YzrVE8634qR6wa
/5zrD7IUgnss5/oiN4Li+esSIpqyk85Z203293g6c6ZtdBPXioQBYFjcLvZmEuDf
qtBPzdb4gRqJ4A1wFR82Sruw2KLzzqIxHxh+AFN/suY1qwNhliVlGfr20CrXkOw1
YgwyvHGhm974YTsaORvGsSsg+rQrfWjkHVmsCPhLW0dyZS+ir0fXhOiwO66GWIsw
Avy04RWwNUCPzLsTSi4FJVBoYaYA3+5S0nm2SNV1LfZJkEL3Sml8V6XrBIIDl75o
AilNFpXDn4cTfovxRwEdLBkbP4rO9r0Fg++TrbXQfZoYRl9g09x1z8dwXUeQgvJH
Xm+RlaGJS791GE/EJSdVPGw4IcWvugBqUMXhe6OkGWUiu1VutAbYxu1JQlX99f7x
R0P8n7T8rawdARFvBrSFNQhhufnkC+iXBiF5Cq9r9DoXUERFOXvygzHDEhtSDecb
pE+Bdb9h+84MR2aT4RmkRAVOaZyicK/tjdDkPl/XDe7JWmDXyDCp7T3EqE1MLd6a
TFdIxg7oMR3AxFRGac+7m1vJ14zl42lILi7wCpDahO6ELOoixeMs1ILj9hqaqU12
1dukaFxXGCgNd5tmJZyl9lCByYw7yNc9UYU77+mNvD79kHNSZ7oYIc4GWQ4ELFE5
ikq5Sr9aOTRa4vdTheeEyHcqImw+pm/qCIvVo38qARjj9qDn2p/iQQJ0bq+k6qED
LeLdbVkSshucqz6eqioTPg5u09iOeCq3ManjLxl2+XvvJx2I4MpSlNTwFKBs/HF8
PgtfNrg+DPryf5eM9XeFFicMx5EHvx2yYV5NkOvSAbqUnxdjqnDZQjVMDijnHG/1
AC+GuZVZ1auMt9Iz3gL5gyS3M/KbbRrFPlzOE+SAD8kdZHDlA9PsE1pAhcofZSYT
RoB/LidGASEOinn0qo9H0ehhroffSPsnX1Ap0fU1iqFbCpu5QQyk+FmcFJP32kLn
N8+ybWYR0SX0h8e0GWjqE10iwEEYNmP2xWcd4I81BpPxiAhtMaPezrxAO+DwiUna
dLrrvn7q1zeF+ZXMQ/5ntxt8zBLo1uwZ8iSlbZqopOtnL14fo042Bf2lLWpHIegd
uw4V9ZmrY/16ER4s1VVBzyzdMHVM+I8zemgQHYr+W8SsGlDfMUuDnKQYNOaTiZ5d
F9ANoqVLhQII8gUqxFwkE1e+pE9ebDllCob98WWThFgJcwJ5nl+TDRMDpsbLItIv
Z+NP4fwbt0pt6Hr1/OhGWDwalilhWLUabmSQyVeYLyJa3KeaERwwC60MNRqJ1GQ/
mYNWQd5Mc4tTcOjlpOCdGDfMNlGOR0+fXiuRJT58CWBydx6N0ZmY2g/e9jBnNxqY
smlqeKmoeYjxW7LxNTsP+/CRoBHRMikq7fSuFg2676jbRIxFyi0zOKR/HJMf+LJP
sbDMksleOMUPjrxXa7W7yb4uIMQ49JHhMJ4gm94li5+uoQ3TauyDaFBJ3kDdJvXj
AU31OxBzN8c6gvu+kmwd6CgIBTvscCmfD5bbmv6rKYzgIiFbay5Sf2BAB34GmPvI
3PEgrAqZ+r/VunI8shhUVOU/JdZvYM29yUeD01U6MvTT9CSg3W87bEjOzJdYopw7
uI15GVvFBGFFTtYOL6MbVX1tsa0EKO1/IgAtMe2f5rXTfA8i30/dv9lVyGVMqqKl
7Jc0trYdtiujrbCPS9BVjbqP5AGxLL2Fd7+qE06/Gk5IhXQfKMnFyEOJ2d5MgH6E
5q/oyzM1QN68LfuiZYJcs+xFKDgvFOVT8ZiB7rUqQow911DBj9SWakOcrnvU2DNr
BXR4e6T+eYvUHhXHJPs8k2x3GnhGQPGKPZyo/3r7D4GYkimMrpStET+fEYXw8gDt
S3D/6Dr2XADDO6pohZbAHbG4GvA+UtLhVREzRshiUPwrtnvHd/15zTeWflPpk754
epplpGBkFF50LyQVuFF6Sl9AaZz8k85Mb/Sg0t+0LCzse3mIlM1My1YsT4c56Lzh
elUAx86sTrqM1EtpEkuijWybGp8OV1XsphhnQ9UcXVAAUILkGQ0vKTuEqU/mz2Wq
RvAELbHkqvfWIIzyqdaxJPrlDH3OCVUNEzL2Lu4i/Q8SnV9gBvYW55jPFtsGQ3e1
BmRdzuAric5WNR9YeADvFEQbIa8EWwndkg5u1pdeeZfmI8Cg6UkuMgXKQKm2VRSs
BShAI/ubuvlNJ+clFRW6eqJcpB/KbcQWfBDidDTlNbqPK+4T/DkAsBTEdSgFMALI
WoDOP+rHbKsJM5AN1xkr4MsMny/uEBxtygkNRqjbktLJ3TTs58ZBHL/OJV3nexvk
6wKIdqXY2VaJM4FSlMLtmQxDdA/zSGquLakGItVo27pwq5koi1CXWmMXFg9dByjZ
x5mROYx59++/b9OdX3UZvduaybETWQ0oEmqw7LHE79TAiGGyiL+KGI/fmKfHgArp
khb2ZLKylLhyg9gb47OrqPTUjDL67TkrQnzFBwPgaKBMQJA+X6oztEsoNAOxiNke
vblp/G1Ny5vAl3S3DZrnZtAR5qpyeaTUJJjTO++SxFFGiAfE8iLg7qwoMn7lvf21
winHxBfO3CT0fXIatR23LYxuKqeBhGIXMP7lJ/Zru82HZAEOQCKgYCGc95KqjqB5
UHh6574Z19RGTce4IuUMc0ffzjkXwNLoIV1zP59Rswf3GgrWNgxcPHC+ykXiEatn
HjeUIfZoXDWfA1njmzt6R4k0divh10LyR2hXfODXyeMo1nVUhWsFlazgz2kXyN6g
OBEHEQsvnC1bz9p2xuXqoJ5QXcB1auOq5l324jotAicInfAop39DRKgdN0K6+fKM
ChXxIgFRXTQk/KzslDyfKJvbjAR9eEN1d8Q/AKtixJK8scXe/E00KlPg4HzgP75r
wK4M7R49dt0SV+ntCdj5XxjkqxjtXD2l4QfwnVgmDQkRZYQJ3brvkIj+sudOKYgi
xJVbr3aXaA1/WW8ck4pxPryZS3y/qsJNUrXE6P1Vb0Oedi7OwN4u+06+j3sTmyZI
p9Lp5ZFHvPZ86K17LcwtfF/nOI3iN25rEI7d72D7fSH/0ZVJFxbnjlbdNKUGFhZl
9tAJfKFXABzkJoiz0k+ijjWaT0JACT/uXbaDjt4G+CvruAtIhFrO/0Kz1A82fnDZ
y4CJ1L2p5o1dnseLY80bSJKZS473ZUioyeNrQgev6luz/yHB2Pe9kq9VJ+WMCccC
rnZuXVtxSqce9mVAA+y8lu+wPX9+2RFlcWTXcvcUMkI=
`protect END_PROTECTED
