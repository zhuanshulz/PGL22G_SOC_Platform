`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QdhfSKeHLHQyikvX6kMnj9030sNo9+13Ttd/eSBqxYtT2dVDWsLsDgwdF5BscJ2p
EsewvJtyVK+MVKuM28OZjh3iSV7xRvSKt37K2xj3EWA7l2OnHVv702mFPTUmGhXW
RClfxkukvTBOT2/oD066qrolAQUhru2htEsJ2gDcf4Jo65+rFgIye/2OGbmmAt08
ygfUaO7mGJS9jaoTCgCqhZlHgxMS4qZElOfbS6QoTl5piujYxXU5V4JUJco3cSdU
YyNqgaja58ezf22crBZG57agwlr7of65ESjfpXHlIolBKigJcZccfGam6BS+lpxX
MMUOtskIZQAtCwqU5IcmKEJVgisbh7lRV/gPr2DekOXbjLGBpIqS6QGna1chgtx9
IeYhTebEudJHcGKbPz95WiDsCJ5x4BQmhLTcbpmykuRoNnQB6yVn+Bc1oQM86ngy
PWHXdgbZF8hE5ZVxdn94V1mYGUBgGNza2Im7QgyA8cN+fOvMZd0mNuhCtPSbXQmo
JLBYWhX5rD96blkyxXLQKDDbViXY9ZEosv4v088dqss=
`protect END_PROTECTED
