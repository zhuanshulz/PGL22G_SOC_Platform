`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTr+1yUk1W1INfiP2f0zZF9Q/NjDXR738auGjZGSKeBoayLRKeX271HgtikIQSIG
AbHTdrC/Y06NhqLnFDYHf1GjC3nircHwad16+uO53JIM4kiW3poYXZyRCYy8p860
tZXLUAtZdi/IxmP1LYTvQRq6q5WEQcduND+kXn9tmsTK6lqw93Dm6bBgoqAoEhXz
mplx6di2sY/KDed7ZFFFdPdlPUXN58wzaM7OH5/rghRZcFhm6Y7Fg39EJtDwvzxo
2ZXSC1T+4uY/CnWlLrkU1Ts+FY58WW/L/tyg6OlIeuRwvS0DcC+99dTFbw/5NzSN
v7oNDpxQ3njHheBidEdximXSf+fHnN/5/1VcC05meQGYHo4J+dL7Fcu3Y3b/H7LX
1fLAofbbJrqha5aRqigigoW4YwQ6EeGEum5jgdDHMJKQRdZaTy8HGhipsq1mSwTf
VZtJsEg7xTOwaoJevnhzFsPcOWlcmuDL1LHrtgPtXh9slgkwo0OEj/WBVJ+4eYEQ
LsmXlImXor52Fto7cLv20Xv65kdUfw9PMFQD0dM7hesPLjlkVOC+PYKr/x891/6S
APSdaAE/uiQYRL5LSlickLrh+/nVKze46Nvd1mVckqi/1phGEc9TbLE1H/ojv1JM
`protect END_PROTECTED
