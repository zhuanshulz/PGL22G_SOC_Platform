library verilog;
use verilog.vl_types.all;
entity V_PCIEGEN2 is
    generic(
        GRS_EN          : string  := "TRUE";
        PIN_MUX_INT_FORCE_EN: string  := "FALSE";
        PIN_MUX_INT_DISABLE: string  := "FALSE";
        DIAG_CTRL_BUS_B2: string  := "NORMAL";
        DYN_DEBUG_SEL_EN: string  := "FALSE";
        DEBUG_INFO_SEL  : integer := 0;
        BAR_RESIZABLE   : integer := 21;
        NUM_OF_RBARS    : integer := 3;
        BAR_INDEX_0     : integer := 0;
        BAR_INDEX_1     : integer := 2;
        BAR_INDEX_2     : integer := 4;
        TPH_DISABLE     : string  := "FALSE";
        MSIX_CAP_DISABLE: string  := "FALSE";
        MSI_CAP_DISABLE : string  := "FALSE";
        MSI_PVM_DISABLE : string  := "FALSE";
        BAR_MASK_WRITABLE: integer := 32;
        APP_DEV_NUM     : integer := 0;
        APP_BUS_NUM     : integer := 0;
        RAM_MUX_EN      : string  := "FALSE";
        ATOMIC_DISABLE  : string  := "FALSE"
    );
    port(
        MEM_CLK         : in     vl_logic;
        PCLK            : in     vl_logic;
        PCLK_DIV2       : in     vl_logic;
        BUTTON_RST      : in     vl_logic;
        POWER_UP_RST    : in     vl_logic;
        PERST           : in     vl_logic;
        CORE_RST_N      : out    vl_logic;
        TRAINING_RST_N  : out    vl_logic;
        APP_INIT_RST    : in     vl_logic;
        PHY_RST_N       : out    vl_logic;
        DEVICE_TYPE     : in     vl_logic_vector(2 downto 0);
        RX_LANE_FLIP_EN : in     vl_logic;
        TX_LANE_FLIP_EN : in     vl_logic;
        APP_LTSSM_EN    : in     vl_logic;
        SMLH_LINK_UP    : out    vl_logic;
        RDLH_LINK_UP    : out    vl_logic;
        APP_REQ_RETRY_EN: in     vl_logic;
        SMLH_LTSSM_STATE: out    vl_logic_vector(4 downto 0);
        AXIS_MASTER_TVALID: out    vl_logic;
        AXIS_MASTER_TREADY: in     vl_logic;
        AXIS_MASTER_TDATA: out    vl_logic_vector(127 downto 0);
        AXIS_MASTER_TKEEP: out    vl_logic_vector(3 downto 0);
        AXIS_MASTER_TLAST: out    vl_logic;
        AXIS_MASTER_TUSER: out    vl_logic_vector(7 downto 0);
        TRGT1_RADM_PKT_HALT: in     vl_logic_vector(2 downto 0);
        RADM_GRANT_TLP_TYPE: out    vl_logic_vector(5 downto 0);
        AXIS_SLAVE0_TREADY: out    vl_logic;
        AXIS_SLAVE0_TVALID: in     vl_logic;
        AXIS_SLAVE0_TDATA: in     vl_logic_vector(127 downto 0);
        AXIS_SLAVE0_TLAST: in     vl_logic;
        AXIS_SLAVE0_TUSER: in     vl_logic;
        AXIS_SLAVE1_TREADY: out    vl_logic;
        AXIS_SLAVE1_TVALID: in     vl_logic;
        AXIS_SLAVE1_TDATA: in     vl_logic_vector(127 downto 0);
        AXIS_SLAVE1_TLAST: in     vl_logic;
        AXIS_SLAVE1_TUSER: in     vl_logic;
        AXIS_SLAVE2_TREADY: out    vl_logic;
        AXIS_SLAVE2_TVALID: in     vl_logic;
        AXIS_SLAVE2_TDATA: in     vl_logic_vector(127 downto 0);
        AXIS_SLAVE2_TLAST: in     vl_logic;
        AXIS_SLAVE2_TUSER: in     vl_logic;
        PM_XTLH_BLOCK_TLP: out    vl_logic;
        DBI_ADDR        : in     vl_logic_vector(31 downto 0);
        DBI_DIN         : in     vl_logic_vector(31 downto 0);
        DBI_CS          : in     vl_logic;
        DBI_CS2         : in     vl_logic;
        DBI_WR          : in     vl_logic_vector(3 downto 0);
        APP_DBI_RO_WR_DISABLE: in     vl_logic;
        LBC_DBI_ACK     : out    vl_logic;
        LBC_DBI_DOUT    : out    vl_logic_vector(31 downto 0);
        SEDO            : out    vl_logic;
        SEDO_EN         : out    vl_logic;
        SEDI            : in     vl_logic;
        SEDI_ACK        : in     vl_logic;
        CFG_INT_DISABLE : out    vl_logic;
        SYS_INT         : in     vl_logic;
        INTA_GRT_MUX    : out    vl_logic;
        INTB_GRT_MUX    : out    vl_logic;
        INTC_GRT_MUX    : out    vl_logic;
        INTD_GRT_MUX    : out    vl_logic;
        VEN_MSI_REQ     : in     vl_logic;
        VEN_MSI_TC      : in     vl_logic_vector(2 downto 0);
        VEN_MSI_VECTOR  : in     vl_logic_vector(4 downto 0);
        VEN_MSI_GRANT   : out    vl_logic;
        CFG_MSI_PENDING : in     vl_logic_vector(31 downto 0);
        CFG_MSI_EN      : out    vl_logic;
        MSIX_ADDR       : in     vl_logic_vector(63 downto 0);
        MSIX_DATA       : in     vl_logic_vector(31 downto 0);
        CFG_MSIX_EN     : out    vl_logic;
        CFG_MSIX_FUNC_MASK: out    vl_logic;
        RADM_PM_TURNOFF : out    vl_logic;
        RADM_MSG_UNLOCK : out    vl_logic;
        OUTBAND_PWRUP_CMD: in     vl_logic;
        PM_STATUS       : out    vl_logic;
        PM_DSTATE       : out    vl_logic_vector(2 downto 0);
        AUX_PM_EN       : out    vl_logic;
        PM_PME_EN       : out    vl_logic;
        PM_LINKST_IN_L0S: out    vl_logic;
        PM_LINKST_IN_L1 : out    vl_logic;
        PM_LINKST_IN_L2 : out    vl_logic;
        PM_LINKST_L2_EXIT: out    vl_logic;
        APP_REQ_ENTR_L1 : in     vl_logic;
        APP_READY_ENTR_L23: in     vl_logic;
        APP_REQ_EXIT_L1 : in     vl_logic;
        APP_XFER_PENDING: in     vl_logic;
        WAKE            : out    vl_logic;
        RADM_PM_PME     : out    vl_logic;
        RADM_PM_TO_ACK  : out    vl_logic;
        APPS_PM_XMT_TURNOFF: in     vl_logic;
        APP_UNLOCK_MSG  : in     vl_logic;
        APPS_PM_XMT_PME : in     vl_logic;
        APP_CLK_PM_EN   : in     vl_logic;
        PM_MASTER_STATE : out    vl_logic_vector(4 downto 0);
        PM_SLAVE_STATE  : out    vl_logic_vector(4 downto 0);
        SYS_AUX_PWR_DET : in     vl_logic;
        APP_HDR_VALID   : in     vl_logic;
        APP_HDR_LOG     : in     vl_logic_vector(127 downto 0);
        APP_ERR_BUS     : in     vl_logic_vector(12 downto 0);
        APP_ERR_ADVISORY: in     vl_logic;
        CFG_SEND_COR_ERR_MUX: out    vl_logic;
        CFG_SEND_NF_ERR_MUX: out    vl_logic;
        CFG_SEND_F_ERR_MUX: out    vl_logic;
        CFG_SYS_ERR_RC  : out    vl_logic;
        CFG_AER_RC_ERR_MUX: out    vl_logic;
        RADM_CPL_TIMEOUT: out    vl_logic;
        RADM_TIMEOUT_CPL_TC: out    vl_logic_vector(2 downto 0);
        RADM_TIMEOUT_CPL_TAG: out    vl_logic_vector(7 downto 0);
        RADM_TIMEOUT_CPL_ATTR: out    vl_logic_vector(1 downto 0);
        RADM_TIMEOUT_CPL_LEN: out    vl_logic_vector(10 downto 0);
        CFG_MAX_RD_REQ_SIZE: out    vl_logic_vector(2 downto 0);
        CFG_BUS_MASTER_EN: out    vl_logic;
        CFG_MAX_PAYLOAD_SIZE: out    vl_logic_vector(2 downto 0);
        CFG_RCB         : out    vl_logic;
        CFG_MEM_SPACE_EN: out    vl_logic;
        CFG_PM_NO_SOFT_RST: out    vl_logic;
        CFG_CRS_SW_VIS_EN: out    vl_logic;
        CFG_NO_SNOOP_EN : out    vl_logic;
        CFG_RELAX_ORDER_EN: out    vl_logic;
        CFG_TPH_REQ_EN  : out    vl_logic_vector(1 downto 0);
        CFG_PF_TPH_ST_MODE: out    vl_logic_vector(2 downto 0);
        CFG_PBUS_NUM    : out    vl_logic_vector(7 downto 0);
        CFG_PBUS_DEV_NUM: out    vl_logic_vector(4 downto 0);
        RBAR_CTRL_UPDATE: out    vl_logic;
        CFG_ATOMIC_REQ_EN: out    vl_logic;
        CFG_ATOMIC_EGRESS_BLOCK: out    vl_logic;
        CFG_EXT_TAG_EN  : out    vl_logic;
        RADM_IDLE       : out    vl_logic;
        RADM_Q_NOT_EMPTY: out    vl_logic;
        RADM_QOVERFLOW  : out    vl_logic;
        DIAG_CTRL_BUS   : in     vl_logic_vector(1 downto 0);
        DYN_DEBUG_INFO_SEL: in     vl_logic_vector(3 downto 0);
        CFG_LINK_AUTO_BW_MUX: out    vl_logic;
        CFG_BW_MGT_MUX  : out    vl_logic;
        CFG_PME_MUX     : out    vl_logic;
        DEBUG_INFO_MUX  : out    vl_logic_vector(132 downto 0);
        APP_RAS_DES_SD_HOLD_LTSSM: in     vl_logic;
        APP_RAS_DES_TBA_CTRL: in     vl_logic_vector(1 downto 0);
        CFG_IDO_REQ_EN  : out    vl_logic;
        CFG_IDO_CPL_EN  : out    vl_logic;
        XADM_PH_CDTS    : out    vl_logic_vector(7 downto 0);
        XADM_PD_CDTS    : out    vl_logic_vector(11 downto 0);
        XADM_NPH_CDTS   : out    vl_logic_vector(7 downto 0);
        XADM_NPD_CDTS   : out    vl_logic_vector(11 downto 0);
        XADM_CPLH_CDTS  : out    vl_logic_vector(7 downto 0);
        XADM_CPLD_CDTS  : out    vl_logic_vector(11 downto 0);
        MAC_PHY_POWERDOWN: out    vl_logic_vector(1 downto 0);
        PHY_MAC_RXELECIDLE: in     vl_logic_vector(3 downto 0);
        PHY_MAC_PHYSTATUS: in     vl_logic_vector(3 downto 0);
        PHY_MAC_RXDATA  : in     vl_logic_vector(127 downto 0);
        PHY_MAC_RXDATAK : in     vl_logic_vector(15 downto 0);
        PHY_MAC_RXVALID : in     vl_logic_vector(3 downto 0);
        PHY_MAC_RXSTATUS: in     vl_logic_vector(11 downto 0);
        MAC_PHY_TXDATA  : out    vl_logic_vector(127 downto 0);
        MAC_PHY_TXDATAK : out    vl_logic_vector(15 downto 0);
        MAC_PHY_TXDETECTRX_LOOPBACK: out    vl_logic_vector(3 downto 0);
        MAC_PHY_TXELECIDLE_L: out    vl_logic_vector(3 downto 0);
        MAC_PHY_TXELECIDLE_H: out    vl_logic_vector(3 downto 0);
        MAC_PHY_TXCOMPLIANCE: out    vl_logic_vector(3 downto 0);
        MAC_PHY_RXPOLARITY: out    vl_logic_vector(3 downto 0);
        MAC_PHY_RATE    : out    vl_logic;
        MAC_PHY_TXDEEMPH: out    vl_logic_vector(1 downto 0);
        MAC_PHY_TXMARGIN: out    vl_logic_vector(2 downto 0);
        MAC_PHY_TXSWING : out    vl_logic;
        CFG_HW_AUTO_SP_DIS: out    vl_logic;
        P_DATAQ_DATAOUT : in     vl_logic_vector(65 downto 0);
        P_DATAQ_ADDRA   : out    vl_logic_vector(9 downto 0);
        P_DATAQ_ADDRB   : out    vl_logic_vector(9 downto 0);
        P_DATAQ_DATAIN  : out    vl_logic_vector(65 downto 0);
        P_DATAQ_ENA     : out    vl_logic;
        P_DATAQ_ENB     : out    vl_logic;
        P_DATAQ_WEA     : out    vl_logic;
        XDLH_RETRYRAM_ADDR: out    vl_logic_vector(10 downto 0);
        XDLH_RETRYRAM_DATA: out    vl_logic_vector(67 downto 0);
        XDLH_RETRYRAM_WE: out    vl_logic;
        XDLH_RETRYRAM_EN: out    vl_logic;
        RETRYRAM_XDLH_DATA: in     vl_logic_vector(67 downto 0);
        P_HDRQ_ADDRA    : out    vl_logic_vector(8 downto 0);
        P_HDRQ_ADDRB    : out    vl_logic_vector(8 downto 0);
        P_HDRQ_DATAIN   : out    vl_logic_vector(137 downto 0);
        P_HDRQ_ENA      : out    vl_logic;
        P_HDRQ_ENB      : out    vl_logic;
        P_HDRQ_WEA      : out    vl_logic;
        P_HDRQ_DATAOUT  : in     vl_logic_vector(137 downto 0);
        RAM_TEST_EN     : in     vl_logic;
        RAM_TEST_ADDRH  : in     vl_logic;
        RETRY_TEST_DATA_EN: in     vl_logic;
        RAM_TEST_MODE_N : in     vl_logic;
        TEST_SE_N       : in     vl_logic;
        TEST_RST_N      : in     vl_logic;
        TEST_MODE_N     : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of PIN_MUX_INT_FORCE_EN : constant is 1;
    attribute mti_svvh_generic_type of PIN_MUX_INT_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of DIAG_CTRL_BUS_B2 : constant is 1;
    attribute mti_svvh_generic_type of DYN_DEBUG_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of DEBUG_INFO_SEL : constant is 2;
    attribute mti_svvh_generic_type of BAR_RESIZABLE : constant is 2;
    attribute mti_svvh_generic_type of NUM_OF_RBARS : constant is 2;
    attribute mti_svvh_generic_type of BAR_INDEX_0 : constant is 2;
    attribute mti_svvh_generic_type of BAR_INDEX_1 : constant is 2;
    attribute mti_svvh_generic_type of BAR_INDEX_2 : constant is 2;
    attribute mti_svvh_generic_type of TPH_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of MSI_PVM_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR_MASK_WRITABLE : constant is 2;
    attribute mti_svvh_generic_type of APP_DEV_NUM : constant is 2;
    attribute mti_svvh_generic_type of APP_BUS_NUM : constant is 2;
    attribute mti_svvh_generic_type of RAM_MUX_EN : constant is 1;
    attribute mti_svvh_generic_type of ATOMIC_DISABLE : constant is 1;
end V_PCIEGEN2;
