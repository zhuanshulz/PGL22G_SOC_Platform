`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNDL+6kdKF+WYzIL/3QKHE8+o1vQNpGAliC80KSyeQIPSf2akIz3EKmhh4dZewlY
Cdf35rlaW38cB20eNeLcW2NglfAJ04xEUwq7lTUbV/4mZ36QTSVohG0VN5cWjdpU
0k/cbcYQEjAr7jXP+agQIJhHniJCAFbeOdT/09j57e9YAKmfy0G/fxnSPZN57t8r
j8e2GE85+XMZh7yNT3VTjWh0YU/dfPYvKsEzKswzB4s5shpQgGr/Yyfax4IXj/89
HOLhjJQ1BbZ2NlygsbVLtepo06r+3qOvZ29jEdKFS4RZj1KiW/tJotZcPusYSmih
KepjWMDPBNv/o4RzPbL0cUAZvkRdccWk9vvlEz6dEoEjiIOgcvWgTyer+1zY5v9M
yDcIdZTtXjdTiHNL3AuehvhNR5F+yBnLQWXxDZx4PvKRpZ7T1VqSpTrwEVa/GIKQ
WPuYLUrsvGpGHYZQArRLP1xgYpUgpE7rMRgQ5X8mV6oc/59LWgGAwigWxLkCQfGj
cedPkbjhrcNZepXHk3AUEHvX9VImnVxyVcTIRnCRb9Rl472fbr7mgwXeApYaLayx
6hcqIy4uNMP7Y7EpkxQjYoy0oyZbxdV218xcuQg6aI2wqE9GotshQh/Q3IvsoIkw
qfMWTMM4tDsUqgK052udFwpDIwGKStQtYITsqpp7HOPjSYqUxtL7xzx1uTXT/X1W
no49YwG+qQEZvzMoKxwyIMLp0JosxXIIKDDvkrO+6SgrXMRJa4A4JzXiOpApAc4w
3GVauIHs2tZRHLwoqdw9vVHH+ssEU4/pTR7KKrjodx9Yu/b+eg3OqK0HNxuXTbiF
DA1fnSe5A1tckM7Hb9pYngZQvx/Xt5L4pUkbqBjo7K7JzCuMiwNQoC0rtC1eHgjc
IVFOQLieFPLwAUAGenehFSp/haGT9FoK2UurajNkqU4/JsXfyg1rjYIBVX/OpvES
WgSgmpVM60q28UXDuKlN3vNhy+r3cgT3sDSHWxFgl/yh/oxKoRFC8FiN3sCxj+5T
0YD82dqdfFiOOO9vcURvkEbXPzsDW/QTOpJcW8oePvM=
`protect END_PROTECTED
