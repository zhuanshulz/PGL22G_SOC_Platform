`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aGhi1C8z3Cj2KAV5ZhDpILmpdF0Kia3H8xN/++JEySajJrRrWg2ZVdu/HuA+twuV
MSc4Sj4JeB/VXg2w9qYlqYwzTF+dGkuX2SE+OxbrwopFiUPREkqTDHxMM6mR3Or5
tusA6HeJxFVYr88QhpwfizcVURsoK2XfTbuvUffdDHpez3SM21gst6SoSJlxmQNY
QoY1Wkm+bELiizkELAJStTIMgjdSfkuuVigiCrn6fQWfOS1ULJz2pq2Lv97i/Ph+
cQmpTZTBgIQBnjD6qs0ouoYKYlQDsHIthXk6v2Ze4cB1KEXjVpW/5MSirHkDVEbh
HQHyKYzCX7AduWHnz+uy/rtpqIKibUzAWTIYjvlfqjWUKLQ49MtvSzCWCTXulvNm
s7LP8185rUmXjnWWRljWZbOF3axbNMNH/48UplSFrqd79ca2wj4Y2tdxYVbH+tlU
CEbbptQtPf68kmFLDoyltS/uMfJoZt1Rt077Ir3QT2ue6QLBNfPULJMG0mxfX/PW
l3Ujt/o8Yonh5gJop4SKk2k+XVAlU7mT0DzFFslrTre5HEKur82HcRkNp5BmI0WF
DRIryWE+PyjFBy70hSqpntHLlfPGUPd6fYUz1efe1X3zTNCHfSG2kvTiEFiJEgvc
MPPMkAGEPwRUCGaCckGnNpuuKSSl11003Z+yNoGRsHyoNahWffnTAF7Fi5S6mfTh
2XWLQDR0258mUhQ145WVWMsdd20NBGX3i0vCTwCUOQWdMI2LtmOa60jfmFSlctCr
zv7ZKmZNsF2crRrTKfRYHky8uMkDAjX50z9dOymM2oqUchSI6vP9wSlbck/LhKh4
Qpo0mlE/lMooTV0WlcSdo+jpFP9b7uAVXfy2vWZj+59Adf+U20/1A7yiMJTyH9yk
BI28gqeCbT75XLd85paf8kSUiaDPZj2YBkSyerh4wYht6C5h5qm49TcZuHSmGHF7
tVZl5ApTzzMui57cT+mB8Y82TJwnbH8ds1Km2iHG0+URIJyFOxr+kdNar24Va7qq
RHethdao+uflwo1EoH7iwDjaUZ+qRjuGR5a3Jes0K+LZbrxyIQml4ZosPbAZFUJT
EcCOXw5f+5ukPeSDInD8rETbmdkc1fXkhWdS0qWXzwYF3Jc60LrcpRhAoRBC82SV
G++1oHc3Y8UepxB89QyXP8ZuQT+UGCm01p3Yo2XnqXeOeusE67hy2LVSjnInkzUq
cxCoL+OBXJ5B5hqOeeHekRKCCdRhvytVt1SfSINbz0p29m3mMqT5HjqdmASAVpJr
BhzsJEv0Y3kP4fVirOTP5B95WleRJ64EBe8IVOy6KMlhmVGQbOYOoWuDLAD81px2
IiWBtNNkBG6Xi7uGc/u1qv/GNc/Q+RX7oUx1gXXA+HS4mcpoTns9YYy4YGlve/ST
ehbkcZ3DZWj01umvDIPSSqYUd/fyVQOj5ZqVWFRgpoSi2/QLVEcNdBMUoNZaHjqs
sCFjF+0nYyjwyN7NVdiFFGcIDknd44gwxkRJWalVMyFsFFO+KAcvfpNoIlXOtWke
SQ2yRkWVUz4Xw8EMu1jvsASHilmBjYsYpW6RwlLIj79r4PusLYDSUISE6pQci225
vh6oAfA3zuUYUV+uRKwhfOVMVnkxbP4g09o8oyaYhi0Zy6++/nO3c6B7oGnAtUB6
ZSVLtoRq8IHrCGED29LjGpjbLPMKYWM0zWkSQBvw5mKqQBPNSourZ7PIp9CGzseD
+PI6iFqSAJwn3PRBeLqkg9y3ZhaYSSbm8tBXKH2+3ECJmtQ+o0CpbtfF1ja/4QgQ
4cYWWcP2I93cmEUnHx0nkt5sJ7M3OI+qUHoOZwmXb1vNd370l+wZI8RppTNwqOgb
IVjANmtmGdXxqa8yjVLL2jHpvqE3hwwTy31n+a0ZUbxnzwm02qisEAxrWIOqq6Mo
1jHK870Q4HlrhySJiVbfvtcYjWfg4XNlZlfk/YQ7qLPjJBqkTIyDT1I5wbbMcFXG
nE9Ydx88wC66K5Wcu4QX0l+m2czpUAsMO5jeb/qoZ1QPIVXnhinkmyFsrIy1s7pW
M90QgmqrCPdr6UrMjpvhwhFJLd00QF5fzi4NFpM9Lf0Wc7oQwsEw+2zrFU3Tu+ZS
td72ckVAMolXIOWrQ9Uw5y1jy5uAgJFYls6yJvEu10yZrNe5yi+ng7g8Xz8bnJWd
xXjJqV02gklHTVnIC4rimDV77RbulJk9R92CfVvaYl6UjSFW3yHEl0dT5TYTaJB4
qM6KgdyD83rgoEV4is9E13d1lWzLScwyYnMT9n1eCTNcV8HGHq4pAlot/xtikF+M
gUFFHVmsFL+IG3B57XX9Lobh/4QV8v2tUWSUay1C2cS6VQ1rThpO/+fz8pD3QjXV
5IacHaqVAdxJKBi0jqzyRKR+7PM09Ivd1JgxRrCBRi1QkIyqgxTeKlohuc4YxkSq
j9MgXSEP9QmYRqtBd3B4klfCFzIfdlzNx1M+GY0wji24PH2THqgIvTd6I/9WyEP6
Rk9kNTPSC27TZ7ZCO1SyjEnGyqcwBO5Juk4LeqNl+fD8r9svyRqVqR3eyrSWjQmy
qR2UbE4PKbArPCYJqIsgFzk/FqBF9/EzLpTqcdBq6/BAh5oRy/DtTN8qGIfgS71b
HV7IWnry1alofhhnIlWPzymn/qOoscjMAEMIA7gAyQtytNqHtD0R4aVBwZNgUKPT
5xdrv/Krr2hgiPgieERl9Ry9ETpe8tZ6veMbt9eSnjIZCJBbhlGC/YftZ/9Lfjpl
kG/uH8AaBIsZzD5E5FbJAlfBmCbJfbV2FkaksKuMWYO/erSZkTZcKyEOTifXQKlL
aPv5MYIwyP8/3ATNfB7QpU8DUdZvIFGrJo9uwc7Dozvaozmz9NiyWVNpu3dA7pNz
Jf5LLuAAYz9BnmoIMQD3Aq5nLm6ns6TkKqDseX4b4T/CryMG/K38QjqQVnMELJfr
U4nE+kXZj9R/JVYuuaFtC3q8HmHVn2t0RpNSx82lJMFXWNzmRDHB6VQPj0PtxLc1
9ewCnXRDXBnX9Nm1K/dku3HP5qhbjfK1NV8a/Av2tcu5UJ2mS3eXBeRiOTV1V58N
SF0yyHrnhjsFs4f/kyig9nH6WNKm8BOfYhThK+z/58KKldGYh7NwTvorTFWbsRlB
UXn8go2uDAZqqt30If/803pOP06OJY6L01cyGDqrE0rOska+hstKbOU4brnocqR1
l1Xdk9sWHNIyhMg2nixrcLNImlyyc6MNTX5W1mJtWpXATXgqIspsa9DaN2ZjAMhX
4WY7xOaabbOpHv3+LOlIhM0kReTXdio+nqX10TlCjN8mZialb0YY/YBWrE50OE0u
GQzsJGPSRZ1K/QM8Cm9m6bKeEqSby5FDsh0NgqiyvYrvne42SJArKTla79VFJyno
GB6UBgRsOj0szNkszt7Uh3hjNaFQfoCEEKASvpB5VaUknRwKDgQC39rOQblwdJjT
5fmtC8RHR2t3CaP1FXjYjO2RzEE5e+83VmZ1d0c189tZ8/fYbWtTRO9usd1y1Tu1
OXfWs8dCZwnutIUgipPSjW3NZRHHM/nGLt06v5eU1zLxKLvz+1CfGTvyB6EXp2+x
8qqYp2+qV+1uwHc3SycNyde4+8coU/zRUEtM7dOIoPT6CidM3N6sX0w1Oed/ReHd
ly1lIg9Hk2R0f2vl27a1Js7oDsM6eJZHYQRM1whwV6OTumaJJxdBWaYZV5pwg5yR
jPTe/Ru3ojkkFpeEZthjswyl2SzcDHcp2LBBsVTiKX+6hrZGX+bRvnEtXICWrSq4
ZEe7/f+P7AWNxUqgTvyCcDOLXY4HcU3WwfyhzWJlPWoxp3e7ZCDR3Y0ARKtheVSs
YNHdKkSvW7X/DGPxiMPIgyZhXKW2Bc0yaC2TDLKjG+i2dm7n7ACXSz9NuhxY86bR
DpcEXbbmQgFh49KabA8O90nTEUn6mI926k+NWZEGTvnEub9hyKl/b3XLr5LZmH36
RW51AOXshc1KvyaFnZyF8UAwIsEGmqpRPUXbCtapbUQUoGKIJYIx8rr1h6MS33XN
mQPriE2ZZ7ZWXPhImKFtpBmn4rfUT1xYIAuOa1f+jFGovevxztq7HiOuSsOgdNgF
uvQMPFqYlzVJlmiKfMPcfQc6dwM/dk+PXfI/hw/qOmJoZRsuqRHscqQ0KAcHhMUT
qfRpNkDVCQcqcEx+dFG3u5y5kZbQrxesX3CsmvUvul72f0U+pSNmID/pTTylAbwZ
jhXb6LZOW7KVD+Dke85K3j+hX0eup0ESg6WJSWsxTkqZ6pF+wGF4gJ5I4kWVoTse
DV4DiumboEPKOhbOCwq5U0HO+Z9n0jNRvFhlG8sXKfGMEsjEuyMnF2dNUxnPJIil
aaU3FIMli8Pxir1ObFtN5RHLXYsgxeC4cus92ysodLiVDTFktvNXTGqhtcsjkBoj
l/3HvFqudT7Fj59/12alXw1SuthuH14WiDRA7O9eWhnyqGYuBQjavtebjeyWrewW
ZQb0e6UHbMEv05rtZz5wW8mw03lOmKOi5gwj+H85T6+pP0YE/oC7S6jYR0e1fJ9Q
UpyGnV3rgMY0iXZyJKjXRF6JUNwzJqRAsL0pPMwUsVxag6HrjekCo7EuSk09XEvS
iWqAFLJxVqY9pb7Z7V70BNezQ5z3m7tMh8GK0k2JEaXNQ3Kb31MJZNFx87B3RPP/
Jk8JQp1DehWuAM6GwLfkdRPN+NwkFuzxq6hoZgogqIZJ4Dfe7aT+dFj02YPaFyh4
WQXSVpdOyPfy23XKUjiGbCRoels3c0eirofIAp7XesUuaxy4Syi7Z2+VuLJrqKft
KkwM2KHJca0QT5mtSGgrrwq/K140FsOrlblRPUancgtjnqrnj5Q2XpMtJPygZX8I
NNd7i69ijUUmsAudJp7BugCGrv6o92qn6UITBFRZ32vkchyT+IxF63pgQ1iXNSA/
`protect END_PROTECTED
