`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0mK13UM+GtF0Vieb1NR8jcujxnZEUOpd38klDNA4O9XKe7W46RbvHZ1RQEeq8+s
BAkjYpZxnsUtYp1L6pOeamCATIoPfhY/+T0UlRuCbwqhj/uREXbTM7gXTeFI0aPO
bVu6apgqLqAt9css7NzhRHvBxKGtVi+haUAgfZzrHTIxr2GpRETdFR0yGaWsQ4Ri
DHwXum/uqGLUhRP9DKeLHHiBuIgSD4Co06AJ/lb13C30UiI+h95D3C1xhP2OZVfw
Knwv7hTcQsb6uBKvb/nIX6l3WO3TFWb9Yg19X/4LY73shxC0wMOM7Ckd7P86dXI+
9vCriejuQ7wtOUrtLcpe8VuO63uMFQAIljyYX9WZ70Ohszku26QGf9P375i0fryH
qhfzp3csmtd6nZeLzoE6jAaEKm9UpjX0+JJ2rsW5+WHr6FqTxU2kzgwcxr53G/ad
zhgMPSH9zqhfAdNKINLbDLj1EMZAcC9f8sfrXyjaLEnuBgoplG4lmF4dXc2qB5mO
b+BGqJNDb390VPLVMiiJ2J5j4pM4J8uI62M0+LAa9r6tMUYPi3SjJ+XVqLd2KdCc
D89/YX7sV3SXhzgEDhAgAPlUpSiuunt+SAkmBd3bv/5I/ux3HLBbM7SLhIc0hDl3
VK2s9bvFzsodvwMiFnO2hYVE4MUQ1Qzj+LLkD6Vn9WzECgkgVjR1JO+VwuGv+TO1
dLvMAzy/Q+PaDQX6BRUwutTfwPRPIoDv22zO4SanYAwN+ypTa34TNMariWiL8yP8
C++ZRP/JZGzUZKqoM4LN/MeAW6ZgPrMyKGo3jTr0bONo+K36FbCaHuuKfzVZny/s
EE676r04rF+YV13E+PTEAU8myaI/1JKvM+nXH6YWEq3GvZHup2TRv38xFC9c+/1V
/Q3Q/dHmNrRWzOqrsbDy5WRBM6U5zB4c5Gb0Obi2Z7IK5LYW8Tz5dpeo1QeJhddo
ImplC/FdMMdvkBSYHY9PcfP+Ayd9kgXC5qB76wck6EXo6veka8hJega3CRyccQzk
KRTAoUUQ0M0Rd1G+MWdbFg/Nef9SIoI+4QahZ3JiGYXzP2CEVH8VRqm/bk9NIhyd
oJWK8Oo9q47q6vp95ecshyGW2w0hg+1eBFq/fAtH4kT2IK0WnCj/X3Cq1lVy5is2
Z1FlOnUUCROAkh/xIkq80gfsMAWQfoFHCb6QiRUkFTo8TegOQ6FUoG+YE8AZR7iy
UOuMQa8rH6kXt+FxjCB5hKGaitxwRZIvAZyV7JBPgQMdMH+D+5sUiZymQmRxlXUQ
kmKR8CiKDrVpEf41pLjjxRA32iShT/Nx8SYUiqWWbdF9icYVjTZeOGIC4h6zBNtS
JxDXNkJFH2VmGdqbhEmb+KQRg3Di2lzPUlhm6woD8759ULsxoTdoDYTE1IPHPBw5
M3WzEm9wuGj5DQg88l/3tVNLwdhXvNYGIeyJ4jyNHM0zJ7c9ieBdgOwcINOUYwDB
OBmcmhjvV8EcqIucSxFfvMhi0ZgVWHgsnb+i9UADzfkmm7uEpC3F6UXyQKmbLqX4
ZzW5YOLIr/VqUfI6/+FSmruICKe7Aqkeqb4kzcNp7OuVTyUVFx7r2lgF69euCgDC
diSQGTlb4nPZUesnyugFVY3KVSx+gEJNlqY8Owddl5pRfDSt5bbUjuxZR7koo/nq
rMWFmsRGuE5bsEHdDusngFpi+O3lyv3WQnVptYWQOwlw9yD98hvAKH7EGKWBu1sg
T1wRYPuzVbbpsvTVdGTM8IiZWaLswlyDMRL37rzV47oDPvfIcff5dimyYAcRXIt5
3a9D3YVFSbZU72Bs7rIXTCoVEryXZfO6S2B32EApU2N6KSiQkksMK3D8ovgZb/m5
Xbb3n5xtVpDW9MTIRMYB7pCy7cjgUQpD3KQCJCA92j2VOj/8ZGU6ivzf05fVzjIn
RvybFHHAldhL2RZtbs4C1nT4XBzFY6cKIsgxR5GqvKWNlW7uPWnkBIbrvE++70c1
5ytovgZb09Ps93kOS3hlog0LmJXohvxd9HQAGzbEab4ATQOGDSZLQAx4KrNnvsYe
zHDG5XHZF519JV5fzcok1Qbct+HzrC+OPRAKpJsJavls2Ju53Eg+wO45l3MQUim7
rTuSiqj3BhC7UFl20o3cAva1iBrhsnKpQCIvflD4A5IeMDLC1xYAUKSCLskyC3eS
/9D60Hc/YnOGCbUOYE9q58ODlA7J9rWgVIi2pfwEis8y4gFGVz9RB+FIK4UfusrJ
tSF+Yvsfk2x0qwMkZQ8KGdmjpOkNUmqKKT07EMRmPZMcHDgH3DhmE5lpwxJuoxeO
o6FPmC3wIH7Vg1UlZVodEC0L9/Gau9AoxWgBUdrtzSiaEP8hK/ZEjpC86XjTV9bT
UlDowlZsp71UXs0Vky3iEC+3xMEHiFHU7XGEIyRAxmwkbiFhvGB9IjXifhXpp/C8
zODO0uvSpO6joq530lHCzty8qt7c1C8jg4KYByLTgKl0Z0gQg9l4XeuIMFe6qZ1O
/t9fVwA0lvMUidb+A+LI7XkhqCfbl1aJcAWM72/5cPInqpqWwmE+CU7zdDUYYsT3
ux++3U+NCO51mxCrrBXU1OMrv5fyylUaI4ba22dHzpfpnQSvLHiwNjh3uVseWw04
qUvXaG/KhAsdcW1O07eaOKp1GAgupcn+gF0gVY61hSgefIafKSZZEchuSi28atvv
iWjmG0rIvfuK3WjD47oNrVxIP9aD2kjn73XM01PAPZtkvUM81jHg+D3wNd1dZaos
U/gioimOkqJlLYbZc96U8/b0llTUx2muCe4zGjRMhzYVqz/P/CQtjiw3nS3XjZJR
VIhdRvoPssznXOZtkop8GkKcQ0jeSu+oyzejZv8twlu4cnFlBka/EojJKs09ZXFW
tV0BRRYpsA5A2vFDzNMEDbNgv6y0MPlXLP58EIRpc0w13Wh8mWdbcgiy0NFCPJr8
x70/OLTlseIBtf/Yjsi07nAlDppDdIwv269HMix2H9PHcArz87vheuz53tsGXQWN
YTKb4AADF83RaTOoVDv3aWaN4qt8+xY6N5WwWd+hfH7GbTjdQqdTNm1eiRUZF2sQ
CB3Q1QhctE0Koa3mHiebtKXgomw5165T6rXxscOcpmTBX2ZJmsRo48KYXy/wygXC
+inpJ0GcU7rdutPWcO9IjZ9gg6htXGA8tX47WJUoRwjMGSSWntuB8CVPhkjwFT/W
Q7bYaUc+cF/PwEwJWaoOiyIhj46/YHGOyhF93FKt9MId91Z7vHCNXm0PxsXQ5uyZ
mPulDshpwOB0+EN9nOIoAELXecQP2Ot0qUVMeXuswKVuYHlQs9Agmd2fZOnn6gLp
40JYUaxzm8sf645VpJCMKPXdIpxvOyYx58tvweHjvqZ5uvBdWVcJbQmYW8Q40cW6
t7iV+IBTXwz5m816l2H0ATDHm1CyXSYRLXSo2sRS5HAk4Vp5+OCDDsITXQaCQgUp
LBXmUG6umDY0pV7yOyDELmzCzT5/gXKlBXxU6l3sYl37fPnuNkNXXQs+IFLhgZJ+
9VREfx8lPAOzFKWy/xH0TVXuj41Hnv+dC3vVrv4VTHCcCikm6TClL5Tx6Z2FFbPj
EuAdWICTfuknk53O9jLErFFhhhW3kNKKyUEluLuIQe0Rzv5zokkDomiobL03P6EA
kRlb+Ne0QfyeUb5wgxEHboL59M8lFOFO68T+c6B7kF7dMkvnNsMLk7RDHzVeqOvb
1SeDx9Dy3in9rSIr2WBUzbr73ajxbxZUSEBhPnXk6NV1qKbwNtWwzPq+Si62OYu/
RGXwepHQDj/1meci+01i+HhkkbbgHk67y4SkB3VENSs=
`protect END_PROTECTED
