`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKLJcFMV88Br41Vmj38T3/uRprwsUvMz96TcaVrK1uv/Mrldu6qsjxomK9DldVoT
7jS7JvAIkNGt6VjuLCK9rRiSqhihIye2bo0fjFou1T008XWQH3fVMh1NFA47EUMd
5KcvE46472JKfigT9Esn3TjoYlix8zBXOsgoKoxqHK/O88mXxHBhY/q47SxTl5+6
Om7RMd8CR9F6Ql9D+buGSeE5Ww1mvn7Keu42qLqobqZvoV3JYFaIH6gBlcag7xo7
YZFS6UxYTT77rrcYNnyRo4Edm21PHGibEy5awirJqSUaJz9Jr6jXyscnhAVvD0l0
2+vvpQm4E9Ee+Ov5i3Vm752Lg93XdUTw6VilzmqzNQqZ/X4HHQNk9dVRt8M23oRr
`protect END_PROTECTED
