`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFFXyHgXJNe4i9oMUahw4b7WEofalRuC7dAiXda6dC51vYVFc00RUXLx6mqOl8wo
QMt+B6q92pP7LRTRMlvqGOi2vr7ei+lkIy+B+yVhSN3INKaOmRsT4bqsLdmyLPfL
x3fqVpbL39rKdzGJvHTIMW0Sv3dhfqG/OCOtIZFprId3r7+NuEraTYxhcsvT2iwB
EkIxMyBK+sHctRRozfPouz8EJVQEbpzLE1s1SfRvTBF6kh7qsWN3yChbH0CzLXKQ
2cHRJTxNHHDltdXV/3tsTsEPKXRIXVTg5bCI1UX7xlbFZ+/0hMWGQy9rcfFe0qmd
sEvLRRxS8fq/dTy1Nwdbruh4RMIy06fHaNTJpH3ISMmKZnjFitktXKDXmD3CY+bG
CHP9Q1tMZe5ZTNuDB56gNEU+WtMCvIS4Rr2tBc1cxO1jo11jDbuWpD3bTflUBoW/
XX6DID5vkA5gG6lLhs0SMet/nJOwz5Cnx08qfFVw5LdGy3DnL/41NqX7LUp2ms+a
WcXRmwm//f9hTFRtult6tMrbh6XWODpvoTQSkF1Bgw3htIUDAGf6Ej+gccbvrDj4
n7ZeNByqMpof5Wdj/YxfMayc1cGHb7ROsXe8C2chVKiDaY3rDemqMj9ErzLmdV7S
JyBRWCeUft8QAnzj8jAHGG9K/cwVLnDGCiEFKf0PtZgprq4O0Dx5DHigspLGKqGd
vhMBq55jIqWbjEEWqeK4V25XLJqredzh0cwvLrvJHaAw3z+snaPvI5XeOe1cNLtB
`protect END_PROTECTED
