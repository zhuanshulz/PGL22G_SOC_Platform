`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjI2UiFfHbsDAeZViYeduLvqEfhWPyUwpiaR+f4XoVuhKoILi880iIwZ1/c4M2J9
RA0682/PgPpZb0k6BD5fn2b1iOaOBYBcuYasyIQqI/x6B49wCMBD/N1o77PLiwXt
SBJFBQIxBXUZQsAfprI0wXcYUL/UEZhga/2YY11mgUfJJ1JkbVjXNIYhcop88Bbq
1aOoIFvKa/hN0jRVXAb/fjVFaqsPMDg06eoxjNrsppxpHM3TIpANZ6pUhWFhH7nB
QIYhcHtXQJy6g2hWqUkFqs80DjePFIouU/Z6sazo48CkEorKrr7Pq8Ge1sF73W+5
aVSTM5ERbws/sujPQ8t27lP0yUI/UP5Sv4BIG4N+6rUN+XKWQrBskUbQY5cw4t95
bgc5t+p4McidiPFgggvnSXBu5ywj+G2FdCCHYeX9b+IvhArQZP4WMN99RT6mBSrA
WzBbSm69BGE5LL/+o+UdZub1sssexzx3yovVx02W7sdE9CUuPO+qpE65uiPxors1
/3d84IWZciafWa908tL0e41nc++xybmZuh1Tl8b0MogjOSOeTuM0QBSeKvpmmf6s
yHBHWCwWMMZVjj8/+u3TQUL4Lw6WRfxCjnTyvCcxsAAuaMTYGyDVxHYdeB+mxh41
qBwXgj/36MHGlKFjNzIcjYzBEAvAsBst2qDWWrtYkrqDZigv76XX7MLX3hzYDUEr
jw9Y5m3NU8wov4qLZbqockrGmTKhdWAe1Ay1Zz/dSMgNT5dRK5i8rcZhc3XqUqPr
6G+lbeoW28rJRFYV+0VNEHl7LtuF8QKVjEihI19qtmoHK5PFXqSs694nwgcv/zr0
k6e2w42HEoi0WJxacJ5SN7yT8wCCc/JIRNM/USzt1qO1zVLzEP3Clji4W5c90JEY
QDftmlkDM4qm44ROeb6zLu0MCoi3pUUYXyizFHb0/EljcITroxTuUQ/grSb/LFM5
6diKJaVeUtzrLTB9NsfQ1hBbJgOb8i1Lex7YXnSbZ8VeLZgaWzUzyRgLydPhDTQ+
yCb2NkYvhYMA/tx2kaz1nRh/vM8O+cAEt4GFNCSOUIgmQmugaouA8ajNDpLnR2wk
6bK+Qt+GZeixLtt8ph+3Mu6EGkhZaDx0Zc5sOCy/T1AnGNrC4cDW3hvbH/2tYKWo
LTCAMNuDQOv25zbVRPYxMYL/YtJyHQ4U1ke+R1zp9yOlLFHaUE7Jt8goa4fHMBWc
p9ZqFYFWt+mue+gJDMrbnzBzz++hZ8zTuwa/hMYsZtohT/Bi8vb9m3WiqzZMoBap
uizX87UQ2sKiaCsDSYR6WBi073C7hS1O8SGkJ6bgBHbtcQmkUbyQglTD8/Dt0Zsr
LCw+ziIwTv4oMZNxuxDYZ4B3GC8cQntO8JW3sWBfA/JSznWlBZJzTL8M26g8MUor
s7a3uMmCxv4F0noT5pubg/FkA5peoB/km2RezLieL8A+mmEpVSQ5GdB2g3my451C
ZhF0sHbQH8AzUQJG737M2xUW7hK1xQzqGAKeVJOCSIFKHuVpZna+dPyFyj1B3OId
HqhnbxFjhe0wajEgNFS6oZQv2Ezk5OExTC7+5G3EYRaJipGZWNPVxQN98UuYapon
QkB53Phb5+TjcfkqnDOiOQEkeobOTbvtypnlc4SdW/a+JamA4lLJxNBOs+B9ARUy
p5g6IVwdXws6W30GStNfk9xeRGS92hN+AVLdsgGmrAt5bQcDYN5vNSl04l+CBI41
z970GUw1rboPUNwxMkVDMhlyBS5Rzrgihux7pWxABUMZCFRHNSedkGg+2Kpcmhsm
u+a/kTo3RZIkNll5fASP2MF+ygt4qxjfJB59Mrikc2weeIQmJYu7grukhBcooM4I
Qq4MNl6xs2ZGvMAbSXf3r2SGbOdI1gP5bRYKns59SL2WEFlP8kh8bn14gaAv2g1e
DKIBoIImr3AVVAEgolgoyZjAiiKnEb95u5OVAD7jKz5n7bBvY+3D10fqelTbKAtx
`protect END_PROTECTED
