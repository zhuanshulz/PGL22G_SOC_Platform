`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0MGEHcLLlxsRyIflAZSnqqEnc1Qc58L7Uso/pw+SzaKEZTjU9Gcozwbhw5iAivS
Ze5I4aR8kPvPlhepb4YBecVDHkMTZJGJr0HZLyFN0S1ua8vtO67Qm12983IiQE7i
B35aVt91q8SaIU6IRdcmePnPQ9+y/jpmJDmxBIFz/AXrtKtkkx9BSDDyxz4pcRhG
YlE2AvcVK1CG21N/+c6yYLbEOnV+Ow/iXk7zEuYMYUVNP41OaIPNesJFFMjh6IKo
jKv3v7Q7z016AnJyy+h+ICv8W+no+QrCkaTqI5pfUThebZ97gvkHIcuF1poEVWJ3
keAm8EXNwdGBxvXTAOB9mbF9e5JBv9g4SKUrDO0CsJWuYkfKl8zUebnQjrj5RpQ+
QbWfHJvH41is5NT40KsDr/f+MGGeHS+2ruAwqgmkC073ncKoV9GHCUG32wqd6GnL
ScBVZS/aaj2/221jEyX+0iCYf/F7AI/UWOrDtlUqozTomtaDL9mSwCenm/fR0Kxl
dEsJwpBepu7yZdetfJx7IBAGjtDYjHNuV1sC20NnqUm+tjn6SCBVYNWJOrjP+e/h
S+QyyCuJhd0BxiGI133Czw==
`protect END_PROTECTED
