`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QXVCZluHIRKi9LDD21f6BpFXIrZGJ5mb7Zb4XB0P7HRmgHDahBE6488UtWHAE5qy
G6AfEGkJkEmsRQH/utL3iK93LRO2t8//IpyUzTafIDsmo56hZs0loZ+OXHsoNctk
meQfPHgnJDJ+nvNvz1EgsaRciSOUvZYcVBRrWYmrjEJslzX1mGQzLZl3JErTNQHj
ijFAIyOVC8QcRwyTF4DHpJdC6ttS3DpPZl/RQmtFUdyzoWImM5xFNOQUgbvRiovA
ymxj6bTsN+f3+M93OLVQZFS4YB+xXgOyMbEerWkzIRp4nE0brGCYk+ok3JyBc807
HynbCFKfGfJtsD6scqFq02S0mZEG7rni8Od/ljyyj3bKGNHbCC8Am1Y5OWfvPcEZ
dk/iNFaoaISiULkjCNXKAc2ix5wHbMzwSfBFMK0tC+soBL/3+fPAPvZaq0ddyj/B
By5DAztDYKePxB2Lgixd+xtkXM7FhkXAx0QJSk6Sjre6GuDiWQQX7aUyliHU+L7A
OK37gPadjnlyAVqqEsFEIPKQyHGP+wOyMpAIt0rFeclxtRMkDnoHlQPDz5FMlMGL
Ci5Q7rN1GFVefBp1HyyX98HoJvzeuy5NPPWlmBKPeCnRtHf5djmSxdxirI9Z/BEE
HJMkdYf3yS2n1q/30IguG0CGcs9f1n6Fjsch5xzUdoWaYdgPbtXqMXGWLDHUBxo/
BuALxC7SLQfn+0TCUZ2Gg6zGioFIANl+7Z7iBphppIug5YD/A8H3SVNF0/AMGy/G
DW9k4BM7cuyGtvAMiYEHVPjOQEf+FEhlo4nlIWeaVdJirOHiQIlR1iCWnx96spef
O2/P8vN82hV6FwlDrWiNFjSQILijKU89PyuvUBPuP9uYUHyoks+2pRqpdxime+V3
BvljH+zCvr5C7UctGsUf2JJwVW/iwYeYJRWXLuztOWz7mAwOYT/D61M/ggY8Lijz
nSVX+FCgz9VQFbyMmx0FLUx1gjtz7rXwFHP97QYx0laOEdTdOwYCEZIGVws+P0H4
m6lsiFPtowZjGTOa7M3LwIUmsDu/A3jg+BiaFyNHlIsTzvLb0mt+kLS5rD0B5Xar
mnwxV7+meQrQR7fdjcTIqDqCxrTd3onHp6YrNbdoxKbYeZEWlZ8y5EqViqDRF29S
9KTyyNPKSeSu5nvy3JV6Jk6Yv+if3d+whXdUJy0D0oduztsvuIhhX7ArPbgZtbRF
fICk7GXSq9YY8OQRQ66Aa6pXvRjSUBesA2onQpva4BR+FqZMeB++/ef/gVc8fwoO
7L39lAPquPFd24MzImEMbDIa28Gwc2txne1PIGHXEzZp7yJUH6TBgDHC5SXk93eD
N+RxcYJIzr6EXXZrD5qg+v0RLMuj9YQx06NQoREPRpKoG1yQNbo2wErQeUjekS9H
Hr4lxQFLqVvMR6KXAG5ln3EHqDkEMgKY5FCIrFJxIKJd6xtYsNGGNfmw1FMziX9L
gljChAB9VEEKlhN7aqqUu8RfS3JViWNZYeVumA853kQZW/SFbVBUtGJrFLB5D9xr
t14vabhrm855nTPgYw37fyges/XFV8UuW6U3+X4krXCksqgS3VRTz+qhxGd6sCUg
9IhT+vwXD18jcryQSpsczIVFbZrqUj/GrxiNOH9PkFLAtdHtFM9XS3B6shM7lcHT
qK1r46l+/p+pJE4FdT0Hx7pKnufktFYnVN72ivcJbGEiGvMtDCySQkvRptolsuoe
EqJ0oYYO3OKI35aJ5yb/HlG8vVodmshUykRbFH8zbooRc+Jb8SjZ9MXf2kYscyK7
Z3kFlC0vfJVJMnpgaxVQoVgfxjzcH/6YpFf7F52PwSUm9doeP6HusBkio2lXAPHC
9PbiEnWC24crEmVtFKfJObICl33Xm4J0edbNlivgY2dY8if3JLJxtz8aLeFMWrdU
qZ0vhv4wR9nRrfxFfruKwnfCCyWDFFQAkZ//D5lTMS8FF2sw0OEphdeb/LyEpa2v
hoWn0FwrXHi0MfuoR0QmF8U9c6fK1lVYv67v5ua2MeIUXAUIgABrtBm4ZWsTjH8P
ur7dEK1iSPfWDfyAPIRI/uOinrfb+/dUsFOi2BKlsfUxL3iGtb6BmPZG4R6pwor4
u+VymjJm2ktYIXjaiJl5thLqUcP954MmtTji9tFMnGYQwkOGZ72F0IODTHJEEsoj
ZPZsfGq1JHm4ABHJSn224Up+zIM9VOK0vzIvzjsFwWT1Wp86LyJXUVvz2fcYmFvO
h1EmcNSZGoTQ8EcUfUVCL+eZpiTzioXLPmv76fI+QSzIGRLzBjZcJ5+v/HXsLt5X
QoNtIqmUKPVjus5yO6ppckJuib6AbT5W6twvT8tCuyOnKGSc4BuvWn4sK+/u3qQK
9qLLxbFtfa8WLeXT1yQvRyhlWHNLbkRKAu1MUQzyJeVWN3jOyru0ZcBEM/rOcDw+
cZATbWWLSn3/wqXB4iPRLtRMTqgSRya32qlMKM7uBmy9GlKLr4QLotuQNef4sy6h
0gpeKgkgXTexWnoMgaBYbdNb01+OS6KuUSUevByA8fhqfd/ZDuxpVWklAvDrZfXQ
Wt+lb1Rup0UKm9rl1KIQhqXjUQw7OAHNNOMWIt4gGUhBLgqAdMcV6os0JtJNIkWd
i7SG4CJAdoDBMX+v8qq6xF49W/tgCD5ykjEcSbAOn2wCcQWz+gnIQErzVBncsS/y
Tp4nsH5Fsit843cojPl/OwGbZAK8zVOrvKIuw7SiYpnwnFTolYTeeHja6Zkm++vk
xHWBhXlrMEAIfKGXEaq5kTTWb2P4vC3ObuIR3EOsFXI0vRpeVh9zspQAa1MCjJ/q
+LYKAxhSUuhlFwytx3pzvI+5rgAVogQvRPDqE39hiPhg4J0YszND/qBGBzvEcExM
b17XAj4Xyrpm7qigSgbvvTC8k8WK+RHR/6ydXV9gv+EbffB5G1t+yj4CHu3zUBE1
QnwgV05fqHyQs2HAGBJcKzF6r75pUxxw2Qa+f1luAisplSWntGFPuLEEdt/Mih3q
dFjNWY/PK46O0XEe+Nyut87ovjUIdupTC8+9hXh4V45tlvPMkqYxukqOGvi61x5X
7cgSIip2PBrOYsXZ+yT140zGDSQmqdGsbwUopCcAD62La4iWZI/rSflC9FZvckco
XRYsG8JH2o26dmozWh6MZg1JgmJ9J2E0b2MLJUFwv3yEbi/nFOG4GX3URnzouLEw
B4xlPmd8zb8eQVfLn4WZJstK5QJcc2Ur+87OflOtSJusMr1G/iL7nMfC/L+QjpXD
eCebR9+UPc8ZHJCcfxWH91URxDDEo5aWIezFwTKbQSZYFN8aadOEWmYuJtOaxHhQ
zf/Lp+wPKoiuZ9WuphdzEftqd68YIUcKY3AP3UtP9Y129fx8dPmBciFxf9aiIJ/N
DYsQxtXfeAoiU+iDYQn+Pgex8ssgLXXahS0IBag9vJog7EEyTU/50tHccprASmin
meoi16RBz1RUb6w6bXl0pFNKD93GB+pAcTD9u8aPN6TO44+YHDKMoorHS/Qf+34v
M7I2jU8Joik9l40jcio/9o6o5Ve062x4gHhHDCg7LRqb+iE1f+yMdMpia7oYlePM
u2kv083F1LzkAdboqCDml9+JSBAYazKUVRSpxy+ifkShD4UnXiu+8ZrkWq+p+VkL
9cjBXZPabMedQRoOYdDJRp3DO7Kzg2uWBiR4KmAu8L+RiazIRlugrrhvYzBpERaX
pBcIRCNRjCobq3bgMAOiT4TVDl46Iynrlky3ljEHRlqMPVfREUYetCiLHyNPq2WX
e203Ea79A5nzAnZmL3qYDUlMJIoaKS89XTbvtSZtUOn1MeF1V3fb0kFuygXTs8jn
wwCAM/XeGwjJTvb1kdfHhJWHCCYK9vtCheCcz3qCKTDCeo/M2OjUIBChptKMLgza
kHlObDhzxbipaFmxmo+eSjCr45jNrStP7lY6i/44wQwy3jzHvZlFYeHHnIXjYj4d
/AsXgWme9csvKcEFywz4vLHZV6Q33LCr9+znMO6Ouh4j86JibkE7AHqbkg3OmBvi
C+mNnBFWkrNoirMBtZzr4/gijd3hXQa8KTjiLvYxLV1S5AlLw0jcyPG7pBOamFUG
fHLuHD2aOf1PdKWRkVBJkpdzXnHcH6V7cNUzqBhRM4J25lSGJeivk8eh5Lef2PJA
L3fEEaPiq0woynFGF3epb56fReKwccKPbjsIXzrxzzT8zuXweAg6y3Uplv/QBQQ2
odQjSzu4o/6A3jURAB1Y5PLHA9+2H8NCrLNxQ8DuoE9iVkA1WQE8tnUhNdEcfsEJ
johaqpABriDy4G33rZwjgsbE0b7BLpNMwu7QzBPMgwG3PFXr1f0xe/pZxx6DA4T4
dywPoXBOL14vo/xylZG+dxviiOSShaDuqkQrEle8RtuELoQiDDItmUTig+qusF9M
J1P/PN6tHI9it3sXcv+RgxuvFehPMeZy+y4O1HKm3cIrSSdESAtlkM24GXO2Hj9S
XIcR5Wv+RqMv4wWubnEwO4cQSkqhm3DaTgDw/y2tfRJskoovzZYUWw2lx4cFIrjq
FSDLMTh0QbbbZAnm2jmZ2zYzwDAr6DRAfDeYwN9YE83dfhpFc8Vg51gjFb0vUzJL
xlIud6pUHi5tXCSeHQsphg==
`protect END_PROTECTED
