`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGyvrQATegSosMMTwCeRy5A3PbA/eJ9sC6dBDbucSwI7c0Opx46KgA40dkYUgPmV
NiG8HPYQvID7GHp8eJ7vD4jFZIFCy3pqK1DT0+oUnL/yFoU1DNwrI5QpGuJyWzpg
RNXKJlB06PhKsvpzXQKyAi79zbCGtz9GvfQ14d28oXDMUxxCnz6EUsDbCMKwvvIB
YP75eNZBfyruqasyRZcoEZYujFvaHf0E5Xg+JbESpxU0E5M8mxs6leM+HIfAV+2b
q31nn1BPxXGQgFrSFD2on4K8ExNqM7wfvjTu2r2hlRaygjQX10CqlwJHuRSxrd3B
KJztghNiRtYq6PCf393irUQ+wS5PPQXfe7/UxMnyfrcNHVPxIUWDmIUYB5mNVFHn
WJ6CzjJRbulVNHYragLgaSkO12GJA5CyDd8p0LhNCe5ZhtC9LaG+dNzwpiRho/yn
FJArWBDKlr5sKuFXxq3tPd4ErTIT6wByVoZX6ZzwmFWMUxy4ahX8cHF4tmqmkY8b
oUVuboq96jUSZuF3N+lSu3/nEpLA1+MY2+1Tbvr64QPaC2k8jjy5jtT2HMJIgcRO
3SJmqt1Sd4hdau640aA7/w==
`protect END_PROTECTED
