`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ff5sKiHzWcLC9O0kVNrahUAN8RnIALYqTmZWnjqyoTgQQaz+HVKBcUv2/0/RP/KG
fjqe/pb1r/v/6R8BWfUfS7atSST2/SI/A4gvMm37JLq3jF8DQwfZtFLRk27CBqw9
OjGFv3QfmckQ4gO5ewbtUdNwa5tjPO76pJG5AqtDu5goC9hB5Jtfh603MEejXjOh
bdLtclSbc4QUfd/+T7Soc8ER3ipRpW54Vep7nZRqKhMQ13Fw29sVmHTf2C2TNkW6
3uFuYUIfPpPj2a9qV+KrYJvWShJl0owa+7QIkdypd8Y8ak9zsmr75d4x+zOXrNBF
NcAVXibgHoxMObyUSt/LMC80pr6Rc3y0qFtaUtqBm5w3zJV67ckhn7TMwe+8RRK+
sspjislO2p7zxfW6LxB7cg==
`protect END_PROTECTED
