`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vE86Jv/vbzYaCGQLO0YtZJFkFz87xWAXt+6Kz5D/7x95lwaI0rnEUR5orYaBJYk
DOuY8gjoA8KqKC+2FTQt26BCLYSknamwbntlj3BuR3n3JWLW9//dkmthI02ZY6nD
4Rc+pCXCJi0mPeuDIWDEj6AbXojHjEScmU5kiT9oFdhZMyqwC76uiWsWoZQgHdDj
A8iaq1+lUX7/CR7F1aC6hjQyxRi1y4tzMun0WfC/OrVVZ55B76p2XrAyQFXL540e
qUFJTbJie/oum4oMz/6GgRu/9QVWA1pKJiKEZBbecmjxFzFUrWWZpYwFCkxsGeX7
MhKfhFMY496UkzwmKEb0WRG6Szf/gTrG4H3dltggtZXv4JZCfcgCC/wDyg/rHWpS
YGIP+pSLEqkEyboPpKO1XBKWEbTjOtAVJNMIhuXbHhV9R3w78ff5NA21wwQeIHXq
iOJqvM0Lsz09h42XTR2AJlhitQubrnM6MExXPUXjSO+G/gYos0H/PYKhSXFNNVOX
f3AY4qhVNBG3mwXGE0GzuXlasIbRxf3qhMTOkE6nXIDpc9BJSXHqyRdQro6WAmwp
D41G4f9R6jQtngEX166kinjOtlN1FNobrbKZMVyRmYiI9psAuUFN7IgWxA94p3CE
HFPxfN1p0c1OoMd/DO6bacNrKeqk3DbnprszggSiybCmn/l7AIrKotvE3zPaDG/k
5vipIH4vXf3eUXEhHqpA+cLzqsfgb3axLgQyX2/gGFlQ8I5+zdgYP78HD/tef2Sc
CZH/2p9m1CgDGFxwGG9VlpJzgRo/scaFgg2HqnLqRw1lkNHLydUkeS0+q4vqtV8C
JMy3SsynL8Ugc7tC6eTG2f0RfOFoizc6EdYu1NdXARvkaYfZd8Qaz3VxqkF6rsyK
WupXfGFo/RWZZVNvfwMKjf5ZQpkbpmcx4R2OAOesVPRMSmB5IKZeuJMtI8Mfc+d5
cHDRVIsxklrUGrIyjiinRMJk/EqgN/jZw3NKcWmMdnrbXV31Ho2EBHyVh+2eSjY7
a4P0AS2PyPGybFCm3UmnVeXG6gR140vNYNydb27vgOgR87o99AZKjMIZuUucTKtO
t5DBFiDY/GnCNwVbCNzoIOrN7njjdi5f1r0VsKU9YMXCrTdQL5rQfE4M4TdSnRlh
GFwPF7ukDNEfSnZwraiN3tw5S8ZYgwBSPB1x7TllUp9+nsNoK12Ks7jPzg+Dk9PJ
erFIcw8XtJ9Rlh2OVVOnqp66tgf4v3ocnT+Je2WwfiM3a/Gzt9iCHochGoXNf/TS
PYSyAFGbffeigDewe5qTVuvyzC37Q/nsfkGrNU96yDDowYRp2wTNAWju6z1zUb1u
bVM/1Zr3015YWRKE2z0ES8DF+mkYdDKh9R/0a8khaTVWPRdzbXFIeLK8TjxsXGS5
HoT2MBf22ET88yNDOlJ4b+iZobZXH14OEunqhNTbmY3xK/9yHdmi6XcvUR/tyYTx
qxDqopqRsY9yhWE8s4VAxoSl2ivZiRfHMC78KgK6xFR1gTzafWRM3kipHnQo+5ht
hjSXb/rVwzpz5VpWz/tS394SNM7ac5dtbMOymVqmbMaNSU1GRRVc8kiojlsqxnlm
Vp798YynrlBn6hjo86ZENBG7Bo3faFgrm2e3aSByrPzrrUm+4auu0MwVRo0q/0lx
Be9Fo2CeUI7ohAjoiAHrlDiRBMK6zj3ovlt+wG1rG/pA3cb5RcCX0X+TimLpcj/W
ErIN6mA75DoPF3/LSvLrdjzTJfHUlwhx8Pv8jinl4E7gEIkzXazgw1Mo//zWip/M
DZXSmaDTuFLh+EyZY4CQ4rASFcl9m6+HUQs8rGJ239zzTtVEbwlr4UOsXH5Oz3eS
lkSz4uUN7l6pbUIpZKkKn33BTjmiz4IXu1om5JreyOD4oih1OqIDnVN7dJ/Hrztl
doyi0gUof5F6PXjB27YzzEShrqdGAOJ0G9zETt4RejqlGgtdydbuRFXLfmzoGGl6
ULREtgQZ4RBxRl4Pv2wEHCrUuHmNpvpREZ5j71yQa+DYTcs88eROp7Rf9z8gjrTh
h81XU1oJrgiCoAqbDiYGxftgHwEZ2G6zI018xgodhL+zPrH/nblGzEPP8sG37lf8
MjnxtImEH0hfZJVkBghSgi5/K01wZivxyMlXrSCb0lliNhNblNKofgRad0bJfi+1
cLqlytzNmABsu+B2u8NLn9UaP6buWdlf+tLDLg/iOT0OVm7C9+CRR/OGimzDnvgp
NHnd0pgQt8TJW1ATPrA4yOAJCDliwfqdpCOCYGQXdmvK5lkplMCZJzS1zfSYVM6o
`protect END_PROTECTED
