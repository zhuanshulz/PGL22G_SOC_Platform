`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+g3NC1nWj/6yOuaay/8XrONlryUxtgC6ljVb/wqukEEBYUrG2YHmZM4jHhHOne5T
Bv53hVXNnyU2MCupJRSjyjsuNcIT9uuf8oJ3+PJcm04t7dWXlctP/B1XRTzbl+O+
WPWEqQrmOSXL5ZC5YDEQPZMhPEIIiA5PPWlE1NPDErDz+goLUNf7875EvF/HuTku
K984yxw28klAEAEJGagnZ1gaPZ0JG5Fd2MzOLI0FPB4BXqEfTEv1OEkkZHWeHhbi
RFiZhY9X7jEt8yJmtM/jQPRaokE8bQ2fYIOk3aFNiMGj187hvcGfhOazgb4Fw9St
bzVci+GjAWEkcEgNsylEcFvOvJMmcUMfYKDBG9ufGYpSATLbHve6eeIGHKUmIUfW
1d9yOTj9y74SXUut4Z9wGaTGuP+yiHZ0F4G9yYe0G/tjN4lsfHU/0BMMr1kFBebC
7aAkuagNxrjf3AmfOEf5kyts7whZ/6d5F6s6ciYXdZcWS2HZWXaxS1ZOUoOQLLmZ
YlUCWcLQwYTHTljq2gqDOZyNySAWik4MLk57NG9UgXhi+YbS3fatW8Ofhn3dv8fK
OyqyQO3dee+pgFqPRuPvNA1z0MQZ8d0U53/uB7ES68uRz6JpDJsQrydHG1FhUerA
CjL63oUVO2yVj9IdzyQ57PedQXT41Qi4CgChrY0o8VqP/a8f4VvUvvd7siaSZB+y
bd7XEnSG6qUsLGkTWlp9BoAt67TWXYydI2uC0SPD4YgZXS1mygmI8xKvGO/JcuAx
BuJL63b5b74nqwUmFe12oXJKtiflZt4VQNLT/http0OvEBzlrfJTtp0hfC3EQ8F0
c/e1hNjcw6oROHcnYPbwdxx5OstRv5R1+Ijs+/HSfyBxzfdrsjLUlbGMS1HzvUIp
9qX5htePq87ld2FJme68xJkWKeFIryvV8iBlKCjyUYoVJBMTh10CyPFKmTZFUJNR
FYm9rpnkFmx5DmjTADVcMUoa/zrbyhZ9aVtfFJOUqt8eXOvMUEJTEx+r61p7JT/j
bzMZSrwJDPeCRP4McIPndx/55Mgq3GdsEhcn3pvOIzA0G/NticPENwXJ6RzuI5zi
5mQURiKLjxTkh0qqdXc6urwXfOKUFp9rmAWRaYc8Aur/XhjU0CLEO88dywF/WB/N
H2PKQSIXzN2WcoazyiYmDCpi3hXuBGDkabjcJ5sBvFAvaFUSPbN3bl++aZxh6ARj
GpplnFlYhYutE3aFXCdcGAvZaYFTICwcc0sTePQYjz0u42sGF5K0/4qCycJLyMvi
od11cUn9is7wwxMGFl8Oy1FeOwGHsIOa7fux0moMJZlwhX0K4EJ8aDFlQmKrqtPR
5IQU8BsEtMnNKDl2OuWcWJv0ZXafNROVPtQeY+Ale19ZSA3LFPxmZHv1/IxZiUyw
LWCDAPfFXdmI+LaM9u+Zf1pJ/I/IWktgcIcWmD7nnjfqvi/8lrQj4z/afmLCmpxC
yDZ8+jU8Ao2pZwJ5ORYrqeviO2sT2BDOFmolg2Rwhcbd9c0upCl8WDAHRryHmg2q
`protect END_PROTECTED
