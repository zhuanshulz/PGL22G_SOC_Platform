`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bEhkRxJjHgycQQxVnw89YIhfoGp6GtQwENUyUIGXMKA/mVpPehTWmD8SuVrcku2u
a2+QSZWXi82xDS3TpYvS2Wl2jrXQJA7Nhoz8kFrz5oQQSJRb7qOFtZFNMuZvNrOG
XlTGF/7jXeylaN6xtauoV8uezJKMWQLKPYmI7TVf5jti5GoQwFGvFeKRTaidy+w7
qWXje9YGabx9QvbT2RiPl21JftolZCzGHcgIDdXtEdrrE7HAVvpMo6CAXG8jM4YQ
dvbJMc33zRRCUNjCKyJ9WL9z+geTm5T0wcC3A8QWDM+bVGnwNqiclJmClTEpjufc
Gd2Q27092FkRjr5/7j6qHFS8rbsQpw08TmebhL/G1klDEdqZmbEpDZq1SDK+ihKy
WkX8DKpnUuMWqwK1eJ6Zy5VRBhDpMisiRmdQWGvvZmtV9laQGUh670g+Uw7yaDOq
IA9Z4jcmgYpWsaeFnlbfDET0FDWgxgo27k6rKYVIPPBpZoBHs3qWcUpKioiFvhae
pdWbtkqq+DN0OXJfXr5ud+JvBaZyiAzUvJT3u5MDWHtCagyiFfxTbHoz624qp5EC
4ggpNcA2lAiJJ3HUNQSuYEi18k4xa2FnxMeDnUUVnRYL5NNpHeiqxQE1ZuKXlluI
J8nWNfgJmuoiJKMkmJiD1Yzp/kMsnb6KCCF877mP7NWprkeGU89r/tGAqEeSysaV
xxcEN43xZlxRQrNlET7UtuKiqGcgdfwFiyAGrLGO/W8Em1YxlMRi9cSU2kgM+Y1T
wWxWF4YV9IAwD1Svf2KvDQOhsTkSyH98cF/EWmX1B4/SeCCmeXrOwZZXuplRXSJI
9pZRzgqPlQrUJsPDIF/jExmfI99VM9yVqWDousm0smzJFIECEWwBZu0mXktKkhIn
cGRl58u+ZDKlWwBgsPohD53QOjyary4WkxZECmpzFv32lmdpXHSrxP9GrDYVGj3X
/cBQn0e44ehoZ2OywNgg511ICnPwpBWUigt6HBFMM60QMRvMR4r3ZCopd4J9Dno8
bO9HZLhlUHQZck+n/eh8erhR0jrUGfA+V/lo7/hDMqUb7ppPI4f8UDTjgm+zb0cj
XSrKvCErBTHNmV+0GpZ3/ZRtNeKvA6hqSrFSXfMppavXaLnfnKazKAYq3XVsZoAE
J3Tc8kiFrMH6gFJDjoRz47jfFkh1umfJI0KDT72Wlqo=
`protect END_PROTECTED
