`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5dX4cASJuua6fBJG9EK+nyqTmpG9kQndLrQmkfx7dJ6WyqR670BcqSZRuzQeUkG
4PS3fQl6Wm6TNOLzappbiTZ7wzMz+Z4tkQxbbBMQGcNeUqeBZRCSdTR1K3/pynlg
mLyTZPwuTzhzP+CQvgozk0omXqDnqJfBNFGt+vPQz+TDvPLaARP7XUDoTOZuWAcB
I7iUZcQ9bS5LZK/a/2QRSUOKY8PSGHMNSmlOSW+Gw0MrcT4ZLmdy6KfOoLqTNMtk
2wX275lN3lQG+oQGFg0HYW/i5jVQxdzikkdMo0Kgmy+kwVySV9Mp/JLiYyZdQ1rY
GXkHutuWaezUre9//05WIIhNZRhxt/WWGMVmnsksidAGF16XgDz8cbYEaTajqEUV
8KOM88v/+i5W6bIaDGRVUxYrWQF1A+wZ2iD0NJ0gi8FOoUE+L8OQiyAQcS0DWUiB
hQQJJD2rIfCU2hk3Z0WZLzAfF7uy/1fKhjF3eAzjnt+i+zYfq044fwEXjKPtJ8jo
`protect END_PROTECTED
