`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UD9pXS5Mio4MkDvDCErRS19NGevJqsfc5t1Ano8t3UxVC8rqIhAJ+QV4kZc72hgb
biqPBGHdEtDqd1KmgxSk+vvw7vn3zrLzEHDx5XLsuNlowda67sEC11fnWzawxYNC
DsIGf6kCsVhMFHSEBmPQHFFbGAsZI4kZTnzoDnmat3H6rSP7QfWEOU7htatDXy5L
dXy/UP+NZE1hm0lyC2/WxYrzvUYTmRkT7+Xx9fAoduKvV9dJxkPP7LV++INjxkbv
Xim0b+BeOD/quPQLKzXsx7AAMkX8sviDw0BPS9KbLXiSvbqxsPczRhZU++XCVmvW
aj7LGPYDDS9c53YGz8c5CTJdeCAbjUMFgzDR6OOBRfZIm/aRsflxzkPoCyUIS30Y
HV6FfD0mZx3q4XCO1IW2EiONcEdMLPb7o8jQ7f3sUYKep2v0WZ6ru3w7V9JfO0CF
teDGeU/9luRPxHRcb2y7fdVuwFjUU1eb7zhWhUitxENLSQ75LBGV4EgfsPBlUcH1
ALnS/I3tuJgoBoHIZnR4DUXWV0Vmf+yOBw43e4gnnRBVsS6enOC86i1M68PBqxfd
XsEvl2gX0Xj/nxl+rfb43lfwR1SD89HPeXw3XW+2bV0gjwVG3fMav0Su7OrQVUu0
t3RjqiD2aNj2MExB7QmtnbA4OFFxkLZn5khBLbDR4UJKDWAX2lNOSI7iX4JJhMIc
dolXF+JNZrWb3LNLInOFb+/qwQdPql6Uq2cGxtqvFBbwAwdn2lPdqVRC0KDQ2YBq
mgyMNNWW6SU9CXUAKoNiC8zW093Btye26nuZuDgk9garut1O0GLMKLVuofrVZOpp
PMiwK2rKcLitPr+SRF3cM10BdLdZJ6eHzd3M3+7Fg7ci87/AregcNlnL8QnTTMxW
kFySRE3Hc5lh/ja/zbyG0XzzYmy7hGnzCNj1+5SX14bnFRjAQEseh5cf42GaVb1z
artw9NLDpF08ADJ3RcRunvrFrwk9PD4wwHBSAhwqfObZzngRop6hR16HbApHyV1K
4DwAevsTnpvMjQSCWVXkW7HWCvKyWTIU0gIhhl5HvWBuuAJCPeSXGuC5S2HaTRi9
Rb/WEEf3F6jnjO30bEumfGgGu1a0c5ALIny8g3oGS4/iiH3EiXf776J2JxRRauqr
pgqc6wHP3Ihsjdp1UmCbQyJorbqS8fAhhxeBYSTuz0LGKBny16LsIZv44pa3d7U5
bRunJFFjH47tuadE3/5h7sLo4fDuf6nhm49NGcAEadu/Ae8DPFJ5dT2fU7PntWuk
pYYNLcKp7A3xYBqyYnJb5g==
`protect END_PROTECTED
