`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5o55HZgMYBwNVSIsz76y2q4s3fAj+aOUoO9kMrjSMrI3lHA9ILEvcRS3kOJNbJMH
Wkt3C7/ZRryKUoGg7hgbManiSmjd/v2390bOPsJCEQhICZDvOSI6qPaXHq1GJ1r9
tZegzsjZAlUsQWKjJJSnTUGdyHxpqm93rwCrvLyRFW+zOsQkLsHyWWxRR4stV6qq
vzZoXdojiFArVMno2EKirF+NzKl1DYSQ7y1gbYcjjtcPCPIB+f+kN0Crs2KiPueP
UL41199SZx7+bHzFaxh6e1I0bTEhs6yNVISjw+0BkLL6te396jUtMIWsyCBgxr2N
6vROIRHKqMQsvUujARlmw0gZpymprQ2RAgTHmSTcSx0=
`protect END_PROTECTED
