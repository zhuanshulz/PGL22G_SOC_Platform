`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZ0IIDqMa8m6AMlNOnH04gppYx0bi8wZ3gwEA23Nxz2yDdRl/Pbvr8FiTgbXrAf+
53VY/9QrOrzuQOI33DIfZzv0UBqB5mMgEW2WtdLRZaD9/Jpsx1KSo3XbocBPOmVk
woSjr1vvoDfR3MTG3T4IJ7aTCeAOEKCuiaDUxy0bCBBsRWPS4Spk3976HQzLSJhn
WiVh2mUuDl2I6Mj3ztthd5IDDqDfusj9hJ5wEq2tvv2Qp+VttnhKXZmHUovOig8t
POwVfJ9lQwtFiVHfPUFY0/2H0FL45lJ5BfJM8JL7nfsNu1Vy0DDigyj7D1ZJXSuy
dodHUwlGrzhCyfza8a5Ubyba4rK/fLl4at5X703NkrRfvIo+9s7zQZ012MHe7FX6
sYfk3PoKEPS7TIuSQy68s9b4cuetAFvXVNkBLiFXDbiu56i/hYu43HmbKW6WmjHM
hYkEjsMUjU+wJVw15MEee/Bm8e3db+aR2YFY0fzlQNnts2s/tbRtY4tcKSUbA2YV
wvIFhtyuZIyNSfjpNj3d+H1kUaVq1VjcRdnyPwH7fLK8HhB/zjyxMNTzPbBx5fH3
9Eg+3qdqL3kVwCWRhVTtougpWR/U4EVttFxoVsuO31CQY27PHA3ZEK8XVOiJO1M8
GR3OCd8xIoo5praNfWRlTzfNB5d8Q3Tn4SysU70qZMB2CwPC8jXcQAMH6xAS0twi
r8aKJOqB+ypyNu8cuoN9Ql9IIVKYCUxeRhw+qGqzrD7EAUv5Q2HZxsxh8BNu6TMa
4ZkxkHAdupwabnjGzgAtrlGCNg7U3q93naoFEYTvq97d/HHwISIKNUu3AL1nCb4u
E5lkXjgvBLJIPOpQDe9F7Qrh6NS/QlM5g5uXxvkBYiuniDRMTFVY2CHAjsGWAHHS
w722qYQ6WrGKKrL9hJqG/yLLJGYmyNblzUKOGgmlRQZ4L9zZIQBs5jLW70j00+T7
hKKMg/V8g5LEOiSjgVJ7jUTcoLPgpU9kZgB+9uTZB/yAwlpkv/FtkhFPeVA1EGGT
k5Uyy33OJxbxfFPcd6MdMkNP4oDsvLw+F3a0OZWMuJqq6BpF6ELtL/6UA/jlH3SS
2CR8xJIYQQZ+Ljpk3BGyQ4iDoolAWFDvA3ANUWUoymoqm25yJkm7CFmaoaJXfFKG
ziqGibtAUBXK1FeWO7Imkf0KEcotByZW9gY0fsetzGB1dpXPP39olN4Zz7cqwtAo
akfTTVoYz7GM1e2QHK70P8faqMKTNiz1NSRpMo0kH2XsWC9xawoK/+pl8qBo3IT/
vf/1A7uuQvNjXr2Exxh+1f8mmZAM+RH348ubXm3VgEj+meuVTIdzEJon275cP+9H
/vWNRXWtGpsO4V7QtTWMzcH5rCf626J0uZYOjwzDoE8zBgPL0+L3OUSlRXrt1Wc0
OkLUTfAhK6I566Dm1iwP41A9lBXgNYjUxI69qPMs4VMcWs5Sh1fDgW3Ldp9fJx9M
ynIffPkOS8tfFvxPr701eKmbw85aVvGfMUI7VdDBUkdFgBE8vSOlNro3bqvliAbV
uQRkmbDhpR5nHa939bY4tAGu3FUX6Hzj7533MwkiZR/1gZ2uo/kpxNEPzq7vo9ay
eRK8hCo8Wlrm4HazdJ8QihZlpuEzgA55I+Lfx7GBSW/8iCSDOctFd8oY252nZthw
G7j0HW/T7jULyObSRhk/eaWLOlYj3QWx4qDlQy3QWmcNdfo0SYJBdAMe1VyREz6J
b42UBJo2vOA4S2+R5uY4TL7zPM27MUmlj8f9bh4qK1Krf4TZnwxUAWesvJVwGZ0z
ZJwCmuPg5d7VTYnmni2NKNsnLCH0AT3D//9mH1juXh4py3LNjHnf86qHR6D+OxO5
0CHWTviegVfkP5HiLvi04174ulKMEz2hT8eT2SF4UADozeXwA3vWAQ4YTA0QnEWc
abPFziW55DcwJxygWU31r9GCQSviwtKPutiS7RP6gNG4nwuq017hy5DTRZGYBvDl
mRfu+CWKAp7MUlk79Jx1WYKFQzRRI2Sg+etPBVINJNNt67hMgCw7PAy5x0n61UAf
/zWUIsedkZW+i1ajMcswaa040J/Pjmz9pucTO5k1GRGLxIfSedujRskNkygz6Nno
ZT5x1gOHIyfJTy86h7IO7CUHed2/1Ofkky6E8c++vNt3FXp+bH77Nd6krzKnWm9/
E697qkCQRBF6tJhWz78liHka2NKoWCARb3/qgemdfP3OzhaBJdXGU7MPfFRY+AhU
ihUNjkuAGyQyS3pSSEk+VPqhNqnUmLeUFeYbxkSlK8wfiRpnfxGTFBeCS5xHEgFG
h3Ohb+aEHH8lNayQakEEjDRPqKXbtewhrP6e1WzgtJQnpQmcqGGyXcwoGvz3XSaC
d1/pQlqVqGtsvhtPr+49Frn6qAaRnFsVxVFh7QM9dOMeWbUjWCW6UqrEmP/6kePV
vvz+kkRAm/cwo1B++EhisLmGKicME7fOMShNDS1uyHyk+9f/tazFc4El3LO8zd+W
DuizDdPWf45s6p3r6ETtsrfKVH61n3zXdYoh0ElRHhUbVUskI6DCYvy2T0O3I4LU
iJPPZM0QNDHF/vpDwK+vHiAjkyaZ07qQbpXA0kKt6li+YMW5tgUs8qsGHcJ1rqJJ
AiWkY1U3GV1uP1yfyaJdqQANX8Iq81wHtlp3CxdZz/cPB4Hz/zV9m02d+nWcctIJ
hRKMnKxb+o9+vaMx1MostvsUXZpxvRNz0Uy0a7JpkmH1X0HHR9cHIsXhbSJNXrEf
I+xewIohlacahcZf8bZIxwpSABn5osHqCvZLTKzjAnEDfZ8uDHMz1+gXF1BxkKLm
GNuNo9DWYjAfQBFT3jlVi+pFhFS1DAZGWiNYsD4ojqjCZIE/dZQQAWZYIm4RLAqp
l1EPROBuH6aRpTDVQXQLy395qqn4GQmFVGyY5+qAJd8cqMFoMv2A4bNWJMC2Bo0f
`protect END_PROTECTED
