`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29/1KcGIjui4QEjLN3cVIVKAUB6jX82TLdigNluhzEGRuNuF0Mfvo/MaQIaYbDMa
1bCtCNwCs5fawxv1sFu6owX/VvTcOsYsRLLdy8p1OTGrS0rK96K4T2yT0V4ftCx3
/fO0xe/xw+W9XGGS27zhJvkdH+Qde4ArNrcpTbV2P/WNwFVymjQEgpAP/gsucMSY
G9c2MK+qq1T1ee7bXK8eHzs6Pym4M2mR5yYoHWYv1fG8hu5TPKUmQqSujfVDAm95
cb4K3K8lvnlfqPfN9klAzt+imTme1aE/X+UcBcyGE9/8LOkAYoc7UpGsEn30aysa
ZmIbaMzXI6XXKSgvbd85FSyRONBz8KQJ6ycJ0ecOys6EV1eP4Bgg7jvkwNfhHh3W
9bIlWUfLPj7Nk7qJWdNDG4H0eltsO/rFxrcvr012BUYrcYVQNmmlV0H7sqtIgtet
oJXJc2HWQ7DgpOwExfaUG65qLZHG+swhzfFTD3IkFwh6O8TCOt6sspgzCdJMUZAa
SBkSoH5XSF1UGYo5SZ4/BO68UJRrX8C2dbspXLQEHZzNV9BtjZifsUAKqmK3Z6Dp
CjjQ6zKp9r4X6CyospOdO4A48EunpauS/pOyOZexMlmo9Ie3guC5pyRMh9+2SiGU
TWXiB7tAlNl4FfYZorjYLkmHr60IA//SIOnaOch7IabpeGJgiwUEbQwG/BPgQccE
LyMLaeg07YH4vqphpQSXkHdwcZtrAQu4F4N3iMDU7vV2miKRXGnxLtZyqIZ/5rp0
MEegR64CZQkHBhU7SjPDdJEqz9Y1idecccoFmluQyj4GFkUH3iomnrjfPH+dmHSC
EviwfVIO683R/DtXX/eef3Ej0f685y5t/YSGDQ2n9zfZTkFgKUCOtBWmkFhwD6CV
KDlJfT2cJoj1FCSVzDOExlAJL5DRl5WMpVRnF+9/OHLxT2fE1RpQWuxMbx4bnsTf
l1H+RJ710Xeo5GZndcujhM8VZCjBBEK9D5kyIrGCODmv9p+FOy8eaADsehHUtzqM
Z9PiHhuiY31w/yhhtYAC74/0KWYmJdH1tlQjrA03HRxh1GWvB1hUQHsPZxynOlDh
Az48EvDV1ky/tJlsNR3YcpR8D/42GO3sPbxx5Q+q+sQvjxjnwP+4LA3fnjVbFBfn
c9C8NYC01Ps7NTEE+NqeI8EGf4EL7TLGY/W6A3zq8jr1EvVPBhplmZvVFTTP+hCR
LnYy5NicW9Kyqlbi5dFgazrt6hoGvnn6frLSnfE/sUJAJMqu9QUj8eG8wv1qpGne
TuhCPeHkand7tOImz6JARiKwfI3Mb7/UkwrcHOyHl7dISfuxoTOY5diJClnEUblR
GNu+d/UcKtx8LjIVWZh2AqCsuYPCJBNlFwTMA5giUJg2dMiAfM0/RXK1cXG4Vz1o
TLtOjR7/3azwvkSEd4K02iGOp5CZHwmVz9I726EdacA2nI5UdQLn6TIhnlP6MONX
ZInYydDmXc2ASPtc9E4eMqVBY4ojswr90J/M8SFrVwbe2/gBfGnt1khIMQoF890D
x9B0TOhskkeXCNfaLYyR6rfATGMnyVmVuwkHU1ai/mdQZ66a7pD9oRIxOegHnaCk
2PIiXg9qAiExDBKK6rd0KreQK5r8cE1SM/VRBXidgGt5piNncTkiQ+hGTvd8zpxD
m+gKqKyud+wxaZBOYpcI9lgULsIvjaS4SVNgcnv5G744//V9b0xbZ2JXce5wAfLB
DqeGl/iY8eXUQHV0NYuvNPt9GjXjvjiXfcViM1gcRzz8HkzgaKIHpACM4br0HZas
s+uSDQ2bfZmbhM3C7IN9rMklxAGKB9WpEz1E7H/mIrerRQIpAg+WFh2mYzKg/OWl
2H5949iUEz6EHU4RxvKfZowJYCVPoQ4mqSGlTc3dw7VXL/REvYzj+0qS3xkdcPV2
ZDB3MAVM9YzsJr73DQVl1SKxMasJO7pAOF6QSHNdFViFLEL1K7E9pT7gr2q4gi0h
YVKKNSRHmAZs+Gynk+9TM+FLhPx6AIlWNm+N36ZXBvsqPfJTD2HwtHUe8tM/go1s
FUKWl/kA+9QHy9XIVGD0miRDtVNrnSAsSBlYX+hNSVS9pDyxMfQRwKLra6Eo0C0+
ZH5+/9gwOHyXh+hZ5W+5T3J1Hsj7OpyPlP1g4FxMfI9NdoyaUMXCZYiyCRP65QnB
SjPg7F9RwqCkErUZLpMRBobdEVFy1sA8w9y5778/SKZARvCzootzkKiqNKbzziIz
aI38jljk3R42mxP/QBSEr8aE/ba2FdyFZVksEgEWxIZ7SDrz8Yd9ALI888Qptg5O
XsgiFESUVPyvYsLUQ5Alfw1poxH3L15hFCvacFR76NOxg9x1ylp1t6E0rcAQWnjm
jeXKEuMvSBiVNPXnGx1RhMrdD3H36txmWnNCA33uXQtc8JQcZwOeTGIREdLrQTpe
TOdfpZyoZQVvzyRm7n2FrTbjKtDKzcMHiSsI4sTFaSpKV2lnNUfc2IMPPUUETZE1
K63qzfZdUAgpDkrxi0vDLPnUSCftg1HbWeDNOxY8nl0wme9RyYnJ0wIBSVCz9pXc
CwLTlOg39zwnx6HDMY5MY6d8oKbedIOBCI+mACe41ha/nGfI6fHo3XXrV8424x94
zHTeZo9INEMdE1divYFpJoXCE9II1LZRQkGCaradp0zpo65x5SLNLM6sHtpp5Ay1
WSj6WuUfGNjGLxisQhiYcD0LLFYXjQlCafG6mgeodQYa+MycKkB22rSMaPt+Nduc
GFIzURqRxkew8QPphBAKTUyz/qB3AgJmROjZ6cCPxwpeVdCu130A1Rfq9+k3EYhs
1Ii9hczQ90wJmbU8ACmdmImAOVkZ8Vvltqclj4lbGlNjnwVBWB5ZZNzIfTi2vXHg
zXQV9tRu2yrSNL2Tu4CNmhYQLfqJLYVacjumVQfDOYgr3lHL99vnt+0ZTnT1lCg6
GbiO3J+oTl7nexbnxIvtKSzRGOXLTJP7/faniTdJivfdWRdcqR9Cm+aA8cRL0gxY
C78D+86Xr0pgaA5xKgPh8RPfSniuyeOCFULDNV2kzea8NgwXw9x3FFkhxP72n+Av
Mv0+GSZZQYfu/u//sdIAVVmPqi8jraIPl5wgcQoSYjsbMT58NYi1lHQ/DldSJ5Ta
tIyt8CKo/4qNaxOqtQk3Edj7m1+TZUoVGOZl8U3ZSyCanUBELE1ixq2N0X77ZlSL
ysTKAggr2JltLMqGTxZV9YEQJe+++5xn4X/F9bxLovnoHLjXvU+DrJdnBhhrrPT4
R5VkF5GahVKrTMuadpp1/5fplnIBAi+7aQdLyC6G3tXZKsRkQEQ/eBIhA5vB5+Fo
M/X0ADX3ffy1BDxHPxsmFRFv3v8nQcMldcLQaLBkIb5Oqkr8LZEIh049bAxyRcFT
LiWijaIaqG0TiTwPLorZUFNpeUxsL/Mj03hXSnnwRX3mV8m9p9Oss3nl80ZrrFOd
HLe0NFJxja2+E32tycoHMh8tuKd1LiDmgOnz3I/vR88MZl7LaGyB9vARG6LaMr3x
CcpKV+sfwj8lME5Ob1nXn939w5x67Mss/yPYf7VD91FAu4kkTwtIju565E8duBiQ
NodNb/HLUzDhhJSqhjomzdbaYrOU6oMuuE2p67DZSImt0bpjfPko3g0ahXpJxtGd
PKGgGdcYD7Vyec2Nt6bkiaWgOS0+NdOQjXocw32jdlMlrPI/NnVrkq5ZOA3Jsk8c
4tXISQYLzoqXYuMF2DjtCfc0WjXLUG3VzaniUWoJ3So6fBSytIaORYsbAtApm/ZR
W0OxUNP8NHXEVoDAOATLKnkpHZr1tCwswvreReHqGMqWOdEIRGQaTZHarVuWnTWS
+07WjuQNlG23kooAU8VGrSBCptW76VUPwGh79mlw54Mv5xMGL/TkgaNnlHmSwGaZ
NJDhg3YHhZf8i5fNdJfg3rQgyRyLiW+WR5HgpX24LmA3OwV8gpzGBpMMd96axXRW
f9LepYcv76Ll9H5y5U/PGVsTOs1qYVhQZWCKPq11CP/g0hHTKnfc2Qk69a4ZZwhN
+9hG4H24DRAzUAJwY2xi+wkeelHhze4cXn2oxiWiioQKicYX5rUGYUdvB8a93Eef
5kkqLW8zqP2DTgLChRVDz81RqmPL0uhEkusxvbzMdEepiJNn3JuyOJAUSPjzbzXi
/fUt2fJnSw+v0gSUJPcssvvx7wJc0XC11CoHQ8NE25Et8F8nOg/beoarZ23OQg6E
qBddMbYvqEsKixH4f2atGSZWWmosfip1lIFicYwNC8ONGKg8CELYS5TeqpiiXlVt
TjzBVC0E3ZX2kR6FpzWRvv6imtABy/YK5kr2pH4TV1FAXBV4moiF+HbxgWgE8Lky
arTwP5ATjqcwLtMG5EsWH85nv99sRfv1cXZtkSviG138xnWBAM4ZxTcKca7zEF88
g9NDaTU1hWSvmrRlpvaYnNIUvVP3UhTjSGvFc1VNos59HhzMZ9JbVXJEd8TEHjTy
+Baf6G2y+v13IrGY6nS3yVwc8cJ0D9VSqiEUj7U5pRozJDtKE2RKWExHqTLEaWzT
6vb8pMa1IAkN4fSMhjl43tUkJ8kfWXVjjqypUkOx+BpTjn+18PFPVv+5aHvMCHUE
7bopkZpSIKeJ7icYgv/23yuQsvOFP19Fm9LWUIu1uDj8/zFll1d+GVZSOOpm9HEp
CJRCA9RdM2D57507Wlu/CG7Ie246T9QnmEmfN1zwSzKKsV8qmODR/watGbhnX6qS
V4Kr1UrDs7AUZMyjHMPyNkrlu7CmxjzD01g9uVNkWeZvb5K06NEthgCxyP4cs643
Zwd4EztiM7xi3sq3NfWK5msvTNlnVJw5hEyjs73JRVggw9GDHw9kpNiDT0BQ+UOJ
adRCYax2SJfHa+M+uadvEk9A5ab7joFzBEqY6ObRSPZxv9xAiHzLFEX0UL0XcsJ0
omKyBBOuGW9Ux7VFyhD04lehK4vhA30ET85ukhcRTs1Oj38fXIoKGSBQmYPLNeLs
H2BebFeWM6qZdDZDNsz174TI3b9LVDdOKlHFJxxob+yOMvzDzADJqRd5PfqZr4aN
s7F4ftvrsDfrn5RzHJlFUckZiqF7zmVcEfcFl41ZjTGFIsCr1m/prWrSwPhPAmmd
kXAN/YY6X7ncwlKEWWmbeoTaQuUlbb01v+XgzDwR7d09cpbG9SoWUkqiAgpjbTxd
Mq2f6l4WZ/i9VkAyIWyX/3SS1Nw9r2Mb7hyOsrJPiGViAlaxdUVpqjW9oNTV+Kcn
0clPsSqfyo5V0adhhfznYzgK5qMcC7XBhIztjcBpeyigykKJQ6FV0BbCabMBT6GY
6UoRnir8pDLRIlyoo2MyrMhbFdAQBDY3eHgiY57u/3tGxPEJRqpBEp1WKAvxkPVn
3epgLvgxax84PaJmkR7dTmFXi8yp+yv+Zrln9O7rh1NkR0Yt6Nz2rJXozuZIcYOW
+FBT8ixlqM4hP8UFL/+ZxSecNC1bp2/bWf5AHc8TkwZZ29z3YSpLLfKCJ4usFyg3
R/LKgO2cnoHUADq430pUk88dxi7vr5r0iN2LZEjnPvhwkNTePtLxnlAWj/5ZJU3l
juARH3/UObWUbVe7B69tFuQnUFpxYdnuvZq49ywUGVrUT5AEp5zUOY5hKUavQsf2
SW+WX0D9RmuafUIDHihRObO9SqHTe1Fn7rianj5bNOvjVhUOvxTSaKW9jVeaTMky
uOqkPfNyy9D0t/UlxAaKZJ4l09MakC9O3MJ1fsnK+t1OJoLyAWR9mOagCX6F2q8U
sLqQ4u8/pCNIF6dpmEDolXF+KYt9O46W4jIcYibIqGyM71orCDWKta/4fBJ8N5qL
/z1+XCVvu/CLccbmXaCvc6X5PCquKZ/KHKpRciima5s00rfO9/ur0v+Zlvl5VVo0
K+TcsfBgL4mLtlPLyBBbbKm9RcMpOqQUgrHlHA+MMBq+2MnY1yL11wLuyJXB5aso
Efbg2ikEXimyL2+E4U2UoOJ2yw/2yjG5gaF9/YB5piEtnqMrGfU3fim34YNKk9KZ
8htlTkM5eJniR1I2riYr8F3rORZ/jPFgzpoWIoqbH/On+FQVD2R6GM7wOplFg0X2
Z4uFEPgRkrbOVwlahVNaGSFnzaeGD5tSDEv6pQCs/VNtqTnchVvt2OTf3Qpc5E5d
xwGsbw/5f+uQcpGMPUpRUb+86hBSGoWeqVdFLS53PxorwTbVaO6CIPBBeJzP7CoR
OSMqC80BGXBFYBuoP2v/qRFDk134qNo6vIxPLA8eLYoRcVLqxq7kWtMjfhdbafOU
S596qTo3Xvbo6INAldeNBnRtuF8FK4oaClRfC25K8ThVGmcuE7Fxjk5X7S3y/Svw
y3ktgbjQY76UkFOoqJ4XTaTDbK3zWZaMZEZCrOdXQf5iRHRTMhAEBQXq6W5cIl8L
pjNGh7ZvRlADTeVmE1CrE6PLqTZXMaynC6u4KzFLynd5YyGhjj+DNtCogFtEnUA8
rWutUOkcXDmMry+QvWmyMwQxj89QYWlahs02IZa5ICBV3j3UOJ+zNUdHn5Gx5gMZ
UpKR52OVeuL7NMtm9/jjDsZ49KbK3YT1R6JMplyEFaXPBiTeyAxnE7HgfKwUBgQy
0l/M5pk8xjLG0WZt2feKIRR9ZQo1STcTNbqBj2+6n/tOaOJWn1sxmhVT937gQaj8
mQiREHuz23wuI/3cYagmahw5Qx05hCcwBVNx6kHhWaoguiPig71zh8KAjy7ezRS5
f29kwq8dBdLJFkmUqXgKsNi+i4gpCJfPeUVbvC/q26AqYuiwgDtcJE3W94VoHXwN
RToRv/DWwangha2BiW2XnPYyHjQ3dmGfNij1OKAg78StYH78guqGEYq+0p9FtBMa
Wnc4ThMjIvUMTY7yW8eZfDW1K+Hv5DPB9dOFARqZAg93iXiAE7+LvNvkfyDhBr8f
eFVWWyOf0UtwnFEcQ6f4ZoaHfNmG4grW9wVokXj4IAGOyxn40eO16SNaQ6rJXw29
CrvG2MR7eNLlgQTON+5RwYnRK33cKcjhsioLrwvBl/87VEg+HQ5OOPvyEiBW9UrJ
OVv3x3x1LzXAlX7Sm7Q6UI6a6UURDM/EE3+N1D+iU8WRG7GOaGtbC+CN8qLDTYbg
BU19t4yBeaA603zCnOmHk3B/WkftO59zJ5msBdQr3EquvoAHAoDXOpZQ4AlxMmDg
d+h2Vhn653lzk5pBZ/mgA04aDb6K3QFwPUUe20vmTGJuGRXJX01f2z9J7obxm8YK
euvJTm+b6JSGYsDO5ASReaMb+PBpSPOfBBxEjHXqniz4Sk152yZqQosRx4FTRbea
bugYuRMYH8LWkK0ZtHP11mib3P8+YxhuAVs/BhkstVpxTpbe3Gp30BjDHMPhZrXF
omhtA73kOv7ARXaT7pJr7eEm/8kJeAPbpNRSBsUHvUdrg2ILpN6vd2c8bXyAln1d
hfHqj37eC0jcKp8F0qIcK2BwoxtuMaOFj8/LiSbkM8mqb2sNoICpLNm958KtLo16
XbaMNfICwnJvN+YnSqyhwG1hdqrl/h44jylebNI/O6QAjlSdBE3CSWzimst9oFQ+
EzgEVMz2AOZI18mdXeBotAMweES4KoP+u+FDgY1Mk822cvLTjiBTgNnEYese+1CY
BxwGCqnk1zVGt6guaJ8g+5c8B/NSEWQHaKS0Gj+Ue0kVofmLMr7FuSC0yAaO9H+d
CNVzGM8kSMGNbkSnHK0Y1tczzj7IAA089vvOQpzaxrHfOlgg5R2xbJ6XmVw9Zb/X
GjqvvrK7aCzL1r6MMt3hVzzSWJDH2uTzD7PZykjfeqdCM1uTrUPoVyFEPysw5Xwi
UHhRPEqYqmE3cCUZWId2O69KU4gateiYkLV3eJ168QBCWenb+X4PG6i9lirn+wZj
+6cdOqcln6eV0vlrrm7ZXjtRp0XalQpJEmyN9+sciFVYN9vpxMoyV8Hj0zr738cq
gtZzmJLmP04GdOFmNTwik5gq/N/1QUTWhNmjNTWklK7Q1BCAm47I+Z/SsedtPYv1
+FcC0G4BkDOnk7e+RQRDaEquL7ACPOi0epW31aHXKJxi48kzi7UH7rJQc4m8oKw/
/46se53TVPZSr4bCGepQ2mlFD/Tk15+n6jTuvz2sfrjwolf0ozlriIRN0q+rrxDA
Wj5FIFyMHKf+3KiTpJwnoXtSfucWAVzzeiq0gOcd/zD5p+yTWjtJ7XLkurPjL2A6
nde8Y8obd0MaEgbo/si16rux/gAgODuTD2NZlsB9PTnLfZnIoJX59g/+2ogzWXYv
YTLZWyOqBO4LcjoGnqjhGdGcMr7SiBSAbjrnR/Pma4A4euwtIT/VIwdNg2CsYpNS
7fivuBHxxdWihkuK1hh7f0CVKuK7lz3VjCMwJ6dqlHr/VLp1l31rejYhc3XcaXzP
LpZMlNxXiA1nkcjJ3QloQYwEyF7zydd2pjvYgZEYnh3sg2CzfZR6ufhBpFdBGwto
pHDd9eooNmcjrbIu11ttJYt/mGv/rQc/LMOTt98aA1x9lEvqIid90+e/EjKQJ18e
1amoEddStVUaGH54BxThUxchnYkQlf5gAj2qbE/MbgfztUC6pX5WHhNwns1FYk1O
jyQO8s+8XkegyVAklyCr3WhvQVz0kzogeJU5qte2Hu4EG2x/4DPLPKUiSX8ziE6q
fYt6uuVkYiB2saaueaFAJgsG7lnwWi953I8RtG0B3vnk+Dr6wCQC0zUQ/pReElZw
dbWqubNcWkhZ29Q3/FcBisKZFaj4S+V/8fIsS0yrevCwmdJyPpH05w0YdkvSofS/
nF1LID1XLEVjBumxT6rU4FpXziz2SJQw/UxCfJYzkf49zEupDuQpe51J8/C8ydjq
OwHtej4H28686dByCr4Z5TNukRznREy8a+UrXLYcdHaMxTC5A0sh6TyT/VDZR1BB
zrIIHuK0pZsr+Qh9AgFm+cTF+ciENKydJMCoTXv75lFYysyHzCkIjhvPU0Q8OtU0
MsOfX71kFtkDTTU8DDhXMDBAFCskQ8BH5ZGcoxR3Sx7qfavql3Sbc800zbYqhI1O
j7HeOqtdGThrRQvUpML785vCLqkUf54I0V8jDAkC45uhckJEgV9x8oNK4TGS9Met
H8HMpsSXy9ZriwB6hkRuDRIg8YvGpyG7Kpfr/KHgwkb06dBAoX9cvL2kkjcdkuEj
tzCFdj5RhU2AmcXur6e7/SkmeVkel0zdvLTzOTRjwRLWRzQwAsxleiaWTSi1FCvh
m4uI912F5N0wYHrpqXJKN61wpYTv7tdwyCjE8o5qglI2pIdUiEz/hMWJUh8onxSO
78BbNtmxcD3qtP84VHt4xEzyNpGXUIVQzmCMGj+vPMX08QO8sA/oeNONN/hQ8tRU
4E7KeevVHFd0watS2gO05n2CkGEDi33oQHoGZQxvXzMfZ3pUydXtJ+cqTTZ82xnS
vygRzKz0NRuk6/1pcaeD4yoRHubLzF4q6EPQqgELsHi6X6hRH+xS4MHQpe2VTp0N
TL81sj99htsWXJ8uxa2VGFSjythlh+IGmcZeiLzw4s6dXsm1iQDXxK4dOzvZYBMg
WIe/KLXgO2/TXhf1Y5VS5OGHv/uGYccgwr0DoocH0NRS7rSJZsx6z3B3CFo5RhKp
S8KW+jtncvvP4l7qGi4GnoFgqbTwAJo3mGjJEsGmhGCZ15l5Pd5uU6GfX3CfIv9p
+yKhESI9ngLNjxym4lbiNspS+OPutyfSeWcCITnBpLsZe871q28/165qRfwZ+kdO
y7CtueOOR3EyWYRsj0V6+xzsyJrwgUerluiAhM5az7Iav4nqrVYte7izJwiH/u3q
kTKZfVhIDwlVAqSzVACMe9y2RoSAvCf6QX5XFt3YFBYWXM74iVhxkkE99IfWw1sP
V27LNhW8fyivlYYkgGxVnl2ZHS+2HhNDiet2huRhHt79pVtS1whoLOF8GIvL+Ktp
yjEMKuyUsoE3gGOBe1oh8KH7I4HIir9BP8URb6XUXfSGS9nuxp+lR6TqGOEKI0i4
AWwqKfglGD/89NiY9M5Fq/tXWPyI2w6fMi8O3uoF9dNigXLKll8874iRh5f8/DVc
VpUBgi0637CohfPVP3MaS4Fkifr5/IB9Wr3hHyiJmau0T3+/ZIXkzB1UZBQIWWD7
O9YWrz4PrI11/JvQhTU++Bmo0vgLW2MhVCn5VO0VI8axfw2tOccRzt/BJK8ISrRy
6ns4wBTJB0bSxJyL+5S22oVyctL6JeB1LzOKrbu+6CfaXn+P6nem2yAIwg25HzYz
v3/xFPlGqQqYixUDp45btGofRrHOpNfOgXGTcMptPzvyzWRC8izUwiQPygFxphjn
+gvKkVVu0YWhr4xDof1765yTGd9m5G8xceXzTkKLK38FnOXr+GK6Uh7zcB3Llp+2
U4HktkSC5ZDjgVA9y9pw/ZxZYWyNUrzNt1qYHoHMADKfDzAH6yPW5FfXNdXL6wRn
a3E4MBdMw5HI7qBvDlUZTL+J2mUcfmEqRMSNj//92howe1nP4xUy2trQ8f2foj4A
Aq7iGG6VnEaWms7oUNuitTRTwcfuJ9aFZ5sh2o7G68jixiKalS85zszGZ+gWzYxX
WeO0qUgv//JbdZdH/8sJpvRk/UcKvBWCr4abqE13OSYV9ApMn88OA0mMNOM0hh/r
OhuTEYIq7w1mug93FofQYnJ2uQ3KOSznwiJBl9C8O+OqUqnswFUTxTD5DtIpBFPU
AbJk6LZRySvoz3DjTijHQP+Zy2pX9ErgE5Y4/w2BQWWzmwOGGR99k6+HMIgmWZdx
ZWglvtM1erlkW+VB1LDsiCZj5ODzDMzWDf4RSE53cErr2FvbeXG9jnl1MtnGjeB3
hO0kjEEcYvjMCyjIGoMELmvXihUWU1I0ORQuQcOOLFK1L4zwP1oQzMAMvixuxabT
3zbO+Ur4BZHSouCKurpSVVWheJ3UNc7Ayq7cYYD7dK3zTIZ+V7M4MM9yZQ7y90c4
sE38d3ymme3oO0mKqKAdUmjGgDBoBJyDcgNPbTJNqOfI5wjBZU8AEeXOKLaNCR/p
xr8YWGmJ5pcU7Q91IIIxE1QXtf/SdYpm1CjWQGJBpP2WPmEjTjkNHbp2j1+XckjQ
BEbSMNyOfjDg4OaB7hulnVS10f5gN1yDoKp7BVok52uHi7EwD23atOcItreZ8Nfx
Hnhzd8RT2U+H7jGaRWyhGD1CsawF5ENQkFw4MRXs/Rj6chllIih+6SmrEpCM0AmH
4hx3za2C0D/GJ8jo4In46Xten1QBGiXPW4y6ZZdhXJ6arYFk49oW9wQ8uA8UYrCP
3ju2BKmnmavBkYiV1bw0ZBj+osUpsfYMNlab7h3I1J+fpnKemKmoh0VaJgzYP+EV
FUP0idee+11SKfnXXJcoydEimgFRCo+XhZd8h6fYamwA/uDffBi3V2YMHO5dpiEp
TAzW3prZKXysiu72Ab4qHIQVPomO5m3wP1DFsJ9mWRV+AWW7i5oOUdDp8XYeFCcW
wY5rFslucpPXYTqNBELjhu1sdAZUKCYNssvLpIa+gzxSMcdQae+UmOiwt/bvCHUB
k+mFImTAz7kWFwNGQB4P9foNta+08RrU8tSKds1YcEU69kFz5GgJL877FYvmRRM0
E6o3vcm4eWg2yfCoBCYiyygJrxRo1Weiuns7JJYLmnwsYrqA3FzXhVZvWTbGk3Wa
AyhUnFjdNoMNy3arfSpxCR2zwFp8tQONn7lIW+EOkohVlAp29s63VYAjMLDUzvhO
uvrjtfFtEoqie4Lu6z3vdB2CsKA5qgg55V5Vshkao3ybzsRLFxKdqrL3+JU1d/Xm
uXfCx4zJkf22GZq7+SQ7TNWDjUjvz5ea1ozVIbC/3Jw6PtyazCYedBBx5vNAh1mP
5xcha0WjP3DltW6NNTDIXzfCNfqvWVCDLVKMT43VwbrlC51RrI6eAald4lekddGA
ea7JoRZOa9h/PPJoJ9tCbCP+lzHmZcqA1/fgW3eqE0rV+jtxQXEPs1q5QOMP/HIh
sA7WoE1dGKLtp0BhdxHc3IrXao3yoEgBiO6VvpVFsO2TwVrkMR1Z4kcU4cf+9+oS
t6ysuTPTfmSOD8cfjvTD2xDW1ge8w4pvjDST5aIK+9csd0yrUT00Dx3Nai7rBtJ9
KVpJrI0WFGrMeOyyekVwWWID+WEiAdy9U76SC4eL9fXuPhq92cbUv6vUSQus/PaD
SfIyEoDt4QINclkFXZ/jiewf/d8RgpVu2JojuoHNXC5+Br9WLX+uFQlXAFLi1nI1
JL/eO/tehEovdn2DMcqsPkzb0Q5YvMVPR5bR9V87QPCXuKAUJiUL/Ye1xn0nH9mk
n3LL4qsU9T6My752eRf72bYXf7Bytp3KxYi0y4dBr0N6+vcSDlgH2fuReaAdTuQc
0FodwhPmgJVmevehr+fCqsF7czGHKtRNeDRpJTZYS61uX+zvuVMYp+oFLA4JVDB6
edT+z/7zXFC5B4IXKZpBb3HUduUU40qzTNaJzVkYc7cqRpvikr7+bxcNad0xsz8L
jGyR62pmBJl/bCtVducm9cXCDbrBoVQSEhEeHFDj0BLBBdUCkYvrlJG8jJTU0YgF
xBbuAtF2z66tqGlnv47+MJNl/6cAsHePQRjYqhMWc/Ci8Hndp+BDGTxhNIa+Nt07
mF6+362ScAgM/wm2+FO+28ZKTBscb9nYgkG5CjpkEMcOVQglzp2FM0iUtQYJKfkd
xnadYiw2sRsTSn8EJ3QzglrjezhLKra1WVs/UEOo6TLARvzWiHlaPkMZCmE2KDMo
/m5EaoHdEjbMIL15YqJD6rT7Kv9GfBQaikirrQpcOxSNFqW6NxVf3SHxiFBk9mZV
YtYtS2DwpJFWt/xOcecYQ7ptXkBUBPXmrHlcf4QK4wGadVRPeKMhywm1OQrBotwf
9dBIW1PbbfWBsWp5jIDTFbKjtkETwJRwt1LRnKqSMKkALjq141TWFw78bz0CY7LT
kvbiVe3MnGz2tKK+0+Pj15DuX7OiApAQe6UbFcjZ1wE5BRHTXZK10yidbgyjyK44
jt3C7ZR8tIWaPceWx610dP2mEW0CoSdTeQePN7lUFYknaAh0SM2G8ho9SbrPXGAK
2RtQJVD8F+3IRJLCBNWiMVRY5MWPL9AfI1PoK4RFYvrj/wsYHPyDohcyLgWykGj0
ehbdDoH+LdNqUwjbxAUP/KjxEzCcPiAaLIYUtvoL/gCb+OZX4d2OMPEySLNwmpsr
KYepH6SsbN5HcsUFDzat9Vr/lIv+6AHXrpBf+yOei35BKFdDxdWF4Js7Q968SBjq
rULMOOyUMMrNVbE5mI7Zh1iLc7iMEYnR9U8TISGPQyBirHT/KqtAib+EfcO2Pquk
cBZmP1wKpnGQL+0yNLHQ8ZbZNe6C3y+NGG/qCm9yLsET07XWFYpYYXTg+5tqFNpO
N3cY2K2S3rvnvN6YeTZ/NOKfQxrcxoKNr5Fy/FfOVogJtp0MflCKJwdxn0SWD0B4
5Z6ax+N6hPTSpxMH8tDOL8UwfIqRV5EkxsjFumjWkceDa20a4s0LnBu299cuk7PR
GaN4urt6U7+fiI3dblIyoXAMxPyylara5BN7OkoLpMMmKMEsKPbux1rnCPftGM3S
z+0KYkR+049epETIlnxp9BSzFbXjISKiQBfBPdpgLxerUSF3PCp4S9Ef8vUapJQZ
VHPsDnPXNuBjV/627HAIFamJqgwmppS1es8lb5j2VFjEX6952YNJmMS1gLNt0Gqh
0yEpoUr1YX38+FU0TnXcmVQJzRHp/Nye1emXGuMkxvxTxevgzeYQwOPr2A5W7IYq
F6p8e9GRQ0IUT87Bc3w73HqfdK8lTNzwqRS0JklTw+L929Dua+XPAk5+hl18jD1T
5Jn+aRt8LqOaUGTtaUcYBuZ0AFq+QB+0+z1OJpT13ORWbTRIAcWWAqIcqaeUeHsJ
T9hcXGcN5siF6uVcHLWr3RF98C9fbyKlsokBwC3OjpFv6L8Myl+a02pU7IeygBl+
4882PHdwCbGNbE9/eVaKZWiKmQsfyFDLY3A3Q710HwyMWXjEV+h2yEUJqQDDAgn8
0MA+JldmeamRtnqnOY9zm+G3Rll3uBXHUkG51y5IdhDQ4dh9X5QjqELtFK9gyrKc
vjPfZXdalaX5QH4S7ievSIIiE4J0ZTSAHIPgYw4xuRkClgAop58YlXi0Ivxg9NmS
h4QG/ZkwgmGYZegSYbzo/1Lx91wsUdwPU21KfTouW7BYrDS2hSREevIqPEap711p
Nx9UrKK0+aXaHU+3fRdrjAjJWwyGzkwem4ZhErWLOJuPcy5uRZYWVZqFOgIg5qmf
GaYFIN4Ko37FJ21s887gcEvJEjftZAgwgBxaFSX23rB3ZJCJeq4eRAEA8m3fox9e
NluqErIihWhej9fQobvLTyjIErUfqfJUOrl89tByDavtxvgSggOR+nkhIMPMrOOd
09XKu3qrIgt1cdk8Vuc8ly4goRYMTIKu4NIiJZQoXAWkeHY2HjJZ2n5/XnzmjRG0
qatPbSTnPhZ6Bbru0ewFU2dfMA5I6aHNTpLaMgQFQMJ/BChUH5Dl0hJLfnMQ9yQI
FNN/Kh+Lf0h/CsvXeG8kipLH3EpuQzGnCGmXG2bgEu1ipIW12sF6RLV45y3H0/k0
WdDK0vhwnlrqmSb8YWUw8PGNVT3ZRcNWG7StvAVjiKr/n6+pAlQIxqFJZFI+42Nk
lqAHGoZYBZI6gYILdV7Od2dQmKTwV3F615W/a2AYGSHo4M6ApM90BALSWSvfU8Qm
BFxCIAruYuoHQP6ypLcQsIPV8hb68CHD8L2n6qIU2mJ5eKtZ/Q1a4RaPSC+76J4z
3HyPsRC65qBwPBDFk+cExuZg7WyGCYo0I84KOqw7I2ORuOLxBbUVGEHIqxe8Yl1P
Bynx2VY22act0hfspAz4Uuqcvcp2fzW3t9zoMv5weaqPEWHJQfwbFH999IfEAkzT
TqCwX0qy8JLvPIRz3yTEpOFKuTM1YhV3cuesOmzHB8eCHdLUwU9E4/KyzyuqrIkT
d5j+N3cCaa+Xs3aUO9u3uFodmpP7vHuRai7YlsFCchJQUVj2KIA+9zS8hMkhwDtT
Xs9/+98NzhpI27AeRFROvDNcUHQgzE7l5rpBkXSWLnbucigXl6KFBOldO6//oo7m
nkw8U2AzmBHTUFhhbe0x1/DAtzVI8IKw+7XWfXP6+OHnA02P4hVGgKoegu6MkMlD
nL2R9bcw1+YcfNl5v+cgesweP5BSbF366TldOy2MoHWfUFQe0A8jTEw4ukgV+bBQ
3YupuXFY5mXqv9sPxvBC9nnWMisLr3yC0r+Inf5kvZ/OaAOM6NnWo9MuCMELlwnj
vt3cDHHHAaf3d98wyXRf5B+xfXZm8kYo24SW7osgAyC/X4Zi1Y37LPM8Fjen9HHZ
EnflVlZFo1vA6rXVymjVYoVdATBimM3OY8fd9HK206+QL93fTxNv3Sn9mCj8Zm5N
XhXCx9emJgWe4V+wDzUOwo7tOJeWA7N17LM9pVUAuNYc3iT7ID09AmPzsmDlaRN5
ncfjyuKZcHMoLnVmJsoq89zRQY6G7s9HIyNIz1ugiirLy/9ZeKtcwGxts+/6UJpM
682NYQKGmy7Ik9AwHsIfZO01Clc7NaN8gjk1+IMTvmxz8RMR71HDoLvREEVtXkN4
GKydSqzmcwD8jdPI2PxHYwUwJ8NuHa3TqXlOwi3s+a/SNbFEE5nIoxvsNiK9qYrJ
hiGxcgnKxfCIbVDLw/oWj9sKs1huQFlaxG1/JQFji+LEdNJNk9T5wSyuXAP4ayg5
MclyoiWgCbDccNjNckVrQOs3w+A1RCw9QUh9rez/VOuwamlhYEYplTKwDAIOJVL3
OHmFkwOG0V2CesOZDgGhb44EsGXW6H/UlxlR5sV8rhHsIejUdlWjCrXS9oRHwnmp
pd6ko00K+7Cq12M7DfX2UmNkstLWCseKRmMQs15BsN9FRqdjn29hCosX+lJcxGvo
uRfW3guCbI/YVmRLfPAwNKdk14zB0gArx6dfPRaK1LA8FUQgSOlzbiyfmE3YhTFh
uqkDjjIUnYo+AoPC8Z1x+PDi9sip29jDab4OPFta6f3Kd0fNvGcqiJ0r9MauW7W5
AsyLCObYFKn2p39JXmbCYXl1FNvhb+gRTgOWlJ63P4O5+8J7n5mdKpJYWHMkScas
KXyX7BERsSIiItRcv3WD20cGTUCYXT/QliE6I6xe/NzkuTYWkIfTxmM7Flt0gACF
LnQnDiRBWwC4nhBOIsUJ/We8zCvwf3OEmzfEExLLaJy0qVKSDAJBV1ZolvPhsial
BdBQWBNNlfg4GZBBkRk8x6nJxgSt0gBd0s3GeVBhRSY9pTpAkKGTWdySDAM8J1zi
dPeEqvE9IZTLFUAbmPuvlWrvSybVbV7XvTUMVhEWgg/Ysj2Cx7Ytkv5NCKg0oju8
eK9gjpiUWSaLFGWMVQ3KERy7A3328BSn5dvRLT7KYUvaCc/d1pX0+6UKL1MhRPB8
gVHJ/BzKyZyZq5NzlkW/NPmw47l/LAB8OLPLWtWlcs485b+9VUfUDGITl8/ygb82
ZV/FHo8FTHJg+IHoZ9WryM46/GvccfIrpw0rdfWA/iQFoETSrrPZHnNG+0tfswxS
vS/RH9ybYhlR70RmovK/rVsLZ19Y9fEd6bhn0nJnvXLmgR7KCBi5yJ0nnc3fDlnn
yGRf7zwLmPfzYNmj4hTA0kHKBL2BYLEgaakVHioX/TsbTIOD5KZwdrSdh3NC4shX
rV2smLhq70Z73pknF5s4erW3YjVObY2WyEwkLf4gKv6Ldan4iffTOVTMb3CCukpA
AME/zYxWxXcWPJ+DCuju4ygenu/caUbCalJdt9fmjJa2aiFjXy/5Mt3SIXZ8/iwA
dRTKWih44pm75isYsZn3QahjA3TD8+v1Gbsg8i6bkYiN6GevT2FmjIadNfAUN8TN
Q6iF5hrvgFO6yrepoxpbXP5ykVa61uxCGsoRAo/DPqejn0aV05v7hXAAGdyzaOR7
uA1Gm53iIZati4xTptWS9Jsd8F82Cuulk8qtwHlQO5szqdnJQ7UMX+W6BfiFO9yX
qixWaaDg12LU9jz6w9y6XtP53tTvPyHUkp6pluk6QcTAZPkE0Xoor2e/o3Beek22
fuaR20wFIg3NrEIIjyvvprzeZV9RtYVUuZfvrgBRAqiw6JlVyi1nVHxpt0ys5uLV
KkW7MOp+Z6ino3s/4BQGBXKMuY7NqmlMdA5bzfcMCBiOBwpuEoe5x9opIP0w/N+l
qyxCLGolEDUDr9j/ssXfNpJgy9FnHZWqmekj4s41WNxOhiZMU0F577RTicp1Hhup
fKXQbytFuPkDN9ezl7eN2vqprd97xLbMgLAGqX3tSsGcCGnlim/Vw1ln75Bf3MFR
5/GS9af6Vlk4Lkujz6I1Tqm5CGan2Ll+OxG08bCZGQzjaJNcXnSlYFjG9Uh1s1/f
P1wRlFqD0gV6zUOAPny4G6cWARl6PdEMWO7tzzhKr2cWZG7o+JALV6wxqPvUuwF6
5k6sV6aayqIKg0kJMQHesCbPTldJ97+HKQZvw9y9CCMvYg2LN3YE8cjSMFCFemqD
4OxksL1y2snXzKskS2IkQIoZRlSFYI29PQybXNPEbgEl9DHf78i2LMcC7sTQiKza
p0FzZ7wj83GGhk89PNwa+mTtnuHJmET42AphgjWBid9Cw/7gVt+BLr+HxfgQuxii
VmYqxbtrPUJWwpgJXbLmSeMt290sIf3zmcmsdZBrrGXU21PVurE4b6eFhHvJDguP
8XvOLh/UXcDrNgS/nFcQ7vggyaW+2fWREpG0m2tbS0ayQcV2HkinWTMXIi6p45JI
/emrrySDIgDBBFGGv0jR1/3/3OgdVZiu/tqSOcDpTSITb5NvCwUrNSylcgS2dvpr
SDYZmfmvXFVypMW/YKHHzOahLu6td1W46YvJTEm+bRnfknKYGcwSP24fFnevkbxC
Gx2UnkLH8fjPZZe77AiDNIFndYJ9/wjk+P4tok9UpPC8Metg5CdWGEXvI5lFFm7u
hTF8ZEmQAXPfCvZc21ZSqpsqJPb8Xh5V5B4EKFUZkolkHxaz7bQIR4/xh5nNfK8v
nHEGgZH09rlVWENDFNre4JYY3+FIWWgLGWda0PsOjs01vo/2jA2pN5iM3O/EmwmX
n5kclN6IBIhhdYOSHGiV13Q3cBFZIl+gbJgXXzh2ZglROp7k8Yv5FGETfZYyTD8x
fnNhmSuYFcecOT3J24YjQXHeoC0bcHClZC8gwdbXj1fljIy6Vhq1qS0ilKNbL/1G
bPJizTO+9eHegl+KemQds3nk6ZJ4JzwCkC1Uf8W50V59iZzmhOCkPI/+lxEjrusr
35xMPzw7P6/YDrnbwcfYtpAHHs+qo+olgTIjB7N2itO5i6+3cVUdydS2CdmtL1Lt
OJ98BJEj94O+4e+2hC++1L41+EmBdTLE1+R+FDO3z0MWggPQrJsWtf2hdSahwn/v
j45idjApBsIr36/gWBDPA7/mpbUx/SEYnJgzZ6OoI4ZmWprEKPSYnZ6fdIbwOsAr
hXa8/TXNWl/7JUy8Lqjh71MtCIlUe9rESuJ6trIIxaHHRcaTtRuR+YdyhdYDX4qu
QS7uKOeXkETjT16jYHiwLzWIxKlcDBVFOM2CFRTrUMJBKc77u2HvudB5oAhhg0Bf
WJesGmdw33T6gnBW+jgWXCFFZ0W/8aHH5cC3+un7IUWtB2zY8R9EzMbTYlyUKy2Z
IaAgvNxPBzksmGTO/CHFS81qs5FN1zJEeQ2WUo/bI+Qdq4shC0YVJFbsTdPBFTf7
JrZrTq9yrkNZWsG6G2ydVkcWbkBL/JZRDG0AF2St9yhLAOZXHh97bMuI88DCC06M
na42JaaZNlDfb+rb3YnUZY4TF9VccocvqJHFA8CB5szfpEJbF45QSUzoLHKyCLa8
R3suFOQp7J+7AjdHwoYblRyH0RKDMBs80jPr1vt9CSsWK9c3LZSsZTBXYFzdclG2
mv0rESg3YNl4BOIBOM8JK+zcF4fz82d83xvYe0X73N4Ks1fXscgXfFy+ndh+70pD
Pl+H5GYOF9v/WRKJHl7TgryYQerE1mkW5KsLuxncUOpSxRorAiYwpnmaPG861Wqr
CaBEWWumWnG8qzAcGlpFQr3+LrNmTSfA9NNTLFXq62gJhAZDLvLQ1BzTlHXO4/ek
nYGAPGi9mGkGbOMYY9CyazSPzRvG8LB2bTFs5an9Ch5ETMiot489MzYdjCxe7opZ
yuoV1ko/fh4mNH0oZe4EeBnA1jwtiPS/zywDrKWla6m3H4Vv2Jp461roR2ZtViQK
RXonY2q4uttJOpSr1NPXlvJhwQaKV9KBmekKDthZqBG8agQgiTRrAU/VUT9cRzCc
gIz7EIoo0L/7u2OT+/4+EC4Jh1faK7nqcYvScxnhqt1YAaCA2U9J+ZWcrbPpgwXU
pt6qDqMtrXVyt2cn1MU969dOkAG4mxhbu0/KLZtxuffPv92hWe9VH4sORZO0ZCwp
gBW8TOGYoVIdRLCcXMMNVgKv/d+100MJhXwTCuFqByjqDTyOperksPLko+iK6duL
wWHAdFxlyFrkz2d+Fg/LIcZN8eUSChV6Ji6XEP2ixmfWK4yWRN33EG/DinSoQvbS
aIFtJgRLTjRGwQLrK4IBTsvW4Hyy3xEI2TC9PaP64fXxdCn/fHyXZ7LHJBLWSQIk
nFcNPtV4OhcGM7AOF9R5VSCsn9DHmyPrnh18MWat/wDr1re2zo/cX2ZAHRUVdTAG
3SHIkUrlYWv1HXC8H1LD/smbxsOMjaojWfUa4ru5CrIkUaEMqyZFM8MUNaDLHSLn
5MsTRg2xPqAsuZGzQjae7d23PP28eM8mYb4cPpEablFCK5Tq4BFEzuhOrImlo4QL
oFQoUxOyaKab1bYClvOxOMI5pm2fXs9LDB7c3Tsa6sb60eC3gr9+FKwd+n3ksJYf
UfaVrC1E8PeYL/gS20A2YF3nLIBaj1c8TQQaEDOxtQX9uNoA7afYsABF1fc9/2xH
LVtI4fSowMA3gSCnXerSuvytX2g7Cg4zWoZjdhh1E/uDlfaZpfMigB7qKqJ2dHlp
habjcS7qh1CRri3wugc3fEEYvuIU4PL21N06Lfhuk7XiNM09ROhELFQznmw7MdcP
GRa+qJ28h3c34/8dy0p5z2kDtbJ/oTPqiy6hZgmmg6gXsy0X1YeEUNSmaNBzb7ms
Ny4+g8JSQHQvpq56lIZ509f5hhKSHKdtGtHNEpqXy9JF5Fe6bU89/rE2684k08X5
D5st3xcX52Cloa10+GVvoUdA60XylI2M5XebuLd0nArKFlBfGLtPCebqK375U+8i
06tzN0BT24tshxFqOAJFdefksnx1d1w8fQzqF2WKFz+b9MQnyv4S++c4yHcodceh
StU18HrbQfTiyfoLUCIIA6UIZRyce2Cm4iOVCXYx+Qamow9yWVMrrJ/6kRHEL7KX
Mje5DKX8QeaIXfCuWqI9ZPbZo7UcbsW1+HlAVoCcejcNkbaKcEJ61sXC7GlEZyox
QMWK06JpWmMucWuRuS8/yefvXGKt61y6KPNYuDAeC/DZPI8CpN/AQoslWGe6zwSE
OGtxc/4toBWwXanhEQ+F5Fi296h4I4dO+LMmsfX3xkzQjAAe0oPBE45xQNIWwTRP
UBRLDUx/qyQ5Ukc0aVxGSdTyUY21GVIF5Yu6BKthHRF+L+UpgrcuV9yRr+gaWsAU
Gcr73QDFZXmfommtL/U4fRO9YwPpAWwzf9zHg+cTEgRs4seLMrVID//IOAFaUV0q
uSoVN4MoEkQ+xessAdT+UsOzu2ocsesxPczA6ca5p6C/331CL+pOmpeQ668V3m9t
0RpNsGyr0Kwz5KkBK+4CvfjKQjc8QI/Z+uiJviBogjjdMB7dJ1Cz578F74zn5GcS
7k+KAlrz3yLUChf+B1p/+pzs1DVWGP6rihDkHhYaOu4XqH0weX2xLX7EbjReO3qF
cf1PGR0HWTrZDuj9TlpMeihN2lkdL593VCH0SmQdgWtF0Tig/ZOX2/SwPxLinDwB
5zR4y8oaNkHMBQLdK8PqdcQ/mfwp3oWAcpOqe5RDSwcK62rvEd3c4dsNNoFqo+F+
V4b/YheO5XV9YSgPAMHE+t0nLNDv1mnMmfxx8PAR9bWukyzD4qTsss0C8dzIA7Us
yoJkU8L/h+GmlJTiFBbG1yghw8PUYEwPn3k8ISXHspgsyRKE97ZncvZjZvUvi/Rp
Vmn0jPyAzUJ8RkD2cA5rjmUnzx04taALzjC3OnyKaLSu/6kRl09eRRjBZHMqzaxG
FdJpWBsoezgQ/tZJCNK87P+3qjWdlei2nKIUHG0y1UmO9kVX7vkonOa7mmiceqIr
CT4YvK+3uOWwtaFJp+dQLUJGRvamuHQPorCqH6qJ0yDmopI5+baz+GkXoASO18E+
pdoY2XNC17Imjn474+wPrYv8Fo1o9nPY5A9Jay/Nuv8eKhu6fosRciPDlQL7I6Qn
utG5brcv5Ha1ExXtyL8w21P7qANUt8+Kn/8iwgMQ73ZvT3l2kYNOc0nPZnMmuH/n
vy9zE7fARcH564xneOgeZBnnmu4FyQ9Md3aUhBqlawYMoVnEJw3B3HPnDft6deQA
KMsQtP+w3l9WOnUoi8HEv9rKeuy6bTW9MG8EcL0nw1ixnOZ13RBHgBqaS7FyKjp2
BkhpMPqEaNo+IFwudSEKp8iUz73ZCWk9yq7ryVwUfjaZuwN/0APsHownm/LXOV9A
T5wWkpfc5Pce6x9o1ip3o4oDPmuipHWCgqFyyWBpza1LU2LZn6XZvBNdfjLaTYWY
VfeTJp8winvtti6ybCDRDoabAG0PlF/s0GZeM8TIiT3gu4Q7dduIOeA3cz0tZ1G7
+j7jWZpu4b978Ugr2wPAm+ay/OhRgtB4yeqrOCrvNo//H2EiEp01Wplx5cyWcoe3
kGQACUh3RYWkWJtDwrEbPKGJj8bU/R5THiC3mJyDE52NIQshduGzS/lT3kdp2EXm
gPKZpIpPIMsrs1v97XIe/nL/O6n9HZO1/LGxJcmvXjsio/V8XYgX0GkmtolXPJqi
OHpaERBJm2I4mCF/wleeXpo1M1ezTaPuU7GpnWy7goiiG5QPWV3cZaV6JkrTNDK+
xTNjPO055xlFpis0Y6J5p4slEaDK21TKz/io8caly2bou1NTf6JYrObV8t3aS7OP
HxKQLAwJHwnYiL6OBail3ZVPpb184ESTNX+MBFXh0wPyaeaFijjo9MXnqfyr830j
e3hTP+4jwPTwYVGJoZxsoZO7h1KLuiTeWjRjKGRqRYk2JPdPB4pbBGrSad1IYnZ6
c7f4qvhZrQEj5ovMkcVGHVH0kVWggUxkBn+cBUviTYtYrYvSdJ+GmHGcxInfqz4E
ulK7UTRGalOnGcZ9Ys3jaNy1fRcIX8mkEXzGx4av+JPnvhJo7Kj0V3IyCf4XRB+E
O4FleY1g9zSDKPvTeP6U33zxiX4avSM5lOjVh5+43I/wzYXQDd/IpSbTvjjnaNdT
TRexxYKiHup7Ak+yYBLWcVeoywoKCzyb98JYAir4JA0=
`protect END_PROTECTED
