`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtyiC/vpr0o2KqnscOOYXR0IJE6diO4Gf1y1RvkP1T3jJd9iCEKitrNBmOm83bQF
Hy8UXFuPSIV2ftwaDPGDuZqxFw2qfb0YB8ww0BEzceIK+giH4oYCfFOAkZzRW7m2
1FhPo+G2NnR0i+yTEHj8AaROGAGRYwrwpo/7QjL/r/tstFLTB7ROgVcGyU3X/9tJ
7rKmz4KuN4sGU7FSnaBXND7tzTSHxXMbYu3SC1z+ae0N5e7uiRz9Yv0DBpHLhRJP
hXY23IvuXcP56IVXxeYcH+G8RBsB24ry1uY/X1V/DzadQZA03hisutt2EVb+gRHf
/sfor290TlSL/fwYJRUXV2+cIFB7Nyif0z8vCdmfp0SOMQwnq2hclAnWFBAvIfFw
w+/helwLXlbxoxV2+o8tNWChr8k0wB16HYg8tx1OUspoC3aOCPzkZ24IDOaCYe9d
5fCJksOZ0J66xGz2kr6ov9VDT8ksXKsUSNFx4O7B5npuUknPuM6SST4OkMqHCliQ
aDVjwhFmhjIoj2Um87U4DWpdlYOOPxlmEugdF41twFehxM1VsM9+wWC6rLuPvuDM
teu9JO0kIBpG20Usx5UV8QS21DBH9dv/LIckheyZR+/JVqXdeRilc+K290AMlUzB
4WVHEkfkugD/NvPil+XfddSe8Sw4iUYbfORtmw8ejOnn7qjhJ3fLS/4CbwYl89YN
rbsfw7fvQCF+N5Yt5ZqLh/jKZhcFW55PAz75CKMxmzy76m6wn7LNJ4wb+MDPW3S5
b5KYxrQ5kk2M2nlAbbTdEw0lFkxbcBA6/G5eKgNFw+CUGXbPbRnZekXWHtVlu6tP
040PgJFocKmaGeDiucwteRYXt1NzuVTHdf5i3jYoQ2I1yY8PAckuve6G5t4B64Oq
Y+cR4Dbe9albetYoccRomC+N8DJH6fqWRW16tkBwMEBRnq4MAhn12Uh/N06iHjuS
ldeq2ZLRypRAseesU9oRhR4gqNiyXcjnwPfzHS3tSd4G+a+FsVcxdb/Kuqzg0YQe
Xhehrw/GwMbOpZoYJZg/+yINC6EDrddZ7i5f2yUU5KrcDkUmdICH+hvkPmczuk99
xhebINRZLxcpg3MXgL56jfJVjRNS6aBLI0p9T8/j2OdqEU5R9iwyPgoIoMMhALWj
uDbfu5qYYOuJzidDc+GC+pQcdi+YNoqZUzLeks3J8okvC+b/5K550VpWbRQ8806F
GKQAxxWFJqH6r4U5KjdB03jO24c2JwV6zk2mW/lNfuyTInqWOaIZEz4ECnCNobY1
wFexcMW3sivqea3b0W9VGZTwPOejannW9+bseT+HqDYxIjT3F4QUmH/6qv7hKEmk
/piSpDO3QdAjl92mP4mqH8bTdx8C7y5OPlUyq5WyFTevliHMlxqG58ZPFVzXgxrY
W+RhN7hohb1wHjYtcnuJA0xL1xjcJpQi0Un6lSY4AqDsH5ATc4eaD9Oyry6ydnwn
NrDiYBT5B8DXoGHdyX/p4o4q7loAESZHIerOyjRGgR6CnciZAFkUHTf7K4E78WO0
ZxI2aEM3iOx0tYwLcC+2fnVJI74nTXhFx0PB5LAaRnS1NckaKEdODGSNGn4nUaCa
nV1vVXI43czanI7sRFmy8b68Q1pINSnmcD0rNcqxUzgTXTtBWfwCxMCvsw1Uyett
RnMtcRPuEWIvDdYT4f39ytI+rBO3kpnCz9RtoSdKLDuJp+1CjDBHqdPbvSYoV+5p
OzZxBkat8HTTadUyKl6iW7PjU2xtO/DC9fBJBQ1bxhjz09qJhisqgVI/GMYeyASx
cqg3ovYVSdKEzRSAh4YkIxyQDqfCpxk6hF3p2G5KNHwi1Po2RQFOQwD/nWTNcp5z
NW084EJesi2NVojpb/O5/+MB32Qmqeov6Q5ytQHF7JCSIAxKUova7VngiB2ReeE4
K7VR8/OvQl1u+o09HQ5c7o2dGckZBWC/8ZdlX9/QY6wO2g65C4We/2nYt3mTeRA6
p9TX/iKP/dBbkDt6yZO6+WzMr7kkgmUQ1UKQ5clT7K/8j4YeEqE/6oAy4/5wG2WW
d8F7oZNJ3bH+2L9GPBT+fKQYhfCnZmLx06ROWsVyuLKsWOutaAoxJZIyc3/UbjAJ
ZBgBVQBgyNTx5sq+QZmOIozt10dpdp6A3/8zn3MODiBCRpwADAkxofQd2oZkZ97R
aPqaRYNvkTW1JDgI6LtaCbauB/gCYNFsCvRhwsZBcYpsFc4ckxRM1f9yUEvJY5CM
l9rteuQ9EI8O9YGoQtgspJrmSatrAVRDdE1KfKEZXgw=
`protect END_PROTECTED
