`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtYYwowWr5qrY9v2wjc5xaXAUchyr3I9uxESoNt4ofWlYbmwNgAlhxjwtUkLPqPR
E39A7RuFY9Ur3/crlAPURxFAsa75fGvU4CSGL3+BLYjN3dOBqtkaLxJixkGwP5r4
FNB9t8qyzpgeUA+oH38FQifI+T+2uCTW31y8JvUtleI/TyacdAlQXn+csoBWT72Z
XODvoiBisxGQCqqV7/JCG9JqU0HjK5sX4RvbFCy0Xts798Vc3QWQaxfF1cuYx1Nz
1EHdQa8sqY+a26y+ZD1MVlFmNDPLuAUMvgFI8UjnTWZ6k/TPJXsdww0kjcH9rEFN
Uyj7JS5WQIMeEFwOG5s0KTrRH9wqF4eKOJ+ED17Y0qmM5vd5sKRGQu/BeSFTyuqc
SlFvzioD4eLCVPPprqASTUZXCqKFiA6VDA8l+oFNSr01cC3PKSrPSOIwWOCCsp/h
oAHDtuw33oWPqK3gKb9aLxS25jQZU1R+5Jwx4yQvPmsmMp2JX81koqFJDP1a/7jA
vNkQWr+1BSnzAiGHEp+dkA==
`protect END_PROTECTED
