`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXulGGqSFGwc2TQHDnnJt5ElF6UaVR2RBJhPBDLKZTW124LY3Kt8PVzICdQgSTVb
NsqXwuHmrDOnWzpjaZ8C4HUSv1+V9P+XUbC585jI/a8aX1aDdFGEOEG0ka1UG770
0yETYfx+NJEyiqq8rtIAZBKyjIh1com0GWkyxyhqs/wqmL71NIRRfDEgPce+JcDm
y6RquVVFzP88e9SiFdvr6StaKHhWmYh26NXocxPd+xyURjEvnnYCgQVYHrLjNCGH
XpsEJ11umwm7Rv3NsNrc8EIPPXJjtotmth+MVLA+yfSfNyVNboH6nLxhrEYdScYf
VDWxfDE22DhuyzJn6q5hkZ4Vp+WXyDjxMuaHkaBemEM5uwlgZmRQ78bpZFIeqZQ/
9ZvWzDzpbwNbl7Mwf1VWThNh5Yeq35nbpOWvFQ36dynJQd0ob3bwgvVTCBW84Aen
QhbQIifJWqck424MuxEwoCIQOtJCI1YGSPYbszeT7m7vxWwU0OCrWAJCpwOMNuOs
cjU5h08iBjLZtjcsu9zBx8bix+PPa/aSR+e5VZqL9rMPXgqsUBm8NncLoFEPt5Hy
P4VzGEVKmsibNwG+3k3h24OVZQS60h60E/jGxwVDKxIE6cte7y+x6aosx0l5eDCd
vZK5MoS5LbGO92S0Pbw2g7Et2V/0PvqfTes6B4ClqcW+ThIBVDhAacxS5Av+fueI
Sv++MCSd1/+wNQDksr+gkkKQLOJg5F/l5HUlF/s3IKH9kvBoLoEtgOhuDvtBBAS5
r/awb20bwUljZDaEgAYszcEC82q9QSFhcY01eCq7nPBegzeazYd7oamHhbjfXNKp
GtIrfkujNM1ok9ZeK9gQWRllJfMmLnDLOAoBRg3A5sMU41GJjrxrKj96UMf5faoU
IGhTjamlzUoo/g7u7M/wmPFrt2PyVxgdgIycWJ6jnktqBxnS7o3CjEe4cRD2LOIy
1g+b34vvKS2tDxzIGatxIWY4jLIP8vSL8oqLV/PvFj6vf0l6hffs2S082tcXtI+e
ubX5wTml4FteRBGIxc9SfZIq4AsgASMPCkyTDqE4XHl6OGgXXCBa6KBZOHS3wziD
qz3TYN7eL/eKe7nhJ8yVZYWroTgymfD3LNK9bp0fjuS04l4T6HTP2Goz9O4qdMgM
XMsg/Z/fZZrMVBOKZXd7WMaHsVswtg8FgEXnUWffkjoHH0CjZu5eTTAHz/+srB0v
OeyiY5Kn1wOXlGv6o9BaXxgXq69QEGepBHY6ToRfE3pC0kuQm4DEROvrWzbczudj
fKU3SMj7SaQyaKPapHt41U3OGAkRU15fmewws4KoAKe49K+soIlBYce6ZR3R9NU/
1/aRNwH+mLht7NF0guf97Pq+eiU/oSQFIClUCqpWUc+pLF92iMkQHlpJSrMSdpMt
UYa9M+flU9/iwIzJ6ZZZzpWq/4bLLdknyDrHdlCXjnIrLSxSGrYt8qRtoX0hg4MK
jguHh9TRWgiOIefNAv6q9Hiyq2/6OUG40tINqO5WmBTM2LiftPCdzi6ipVL/TitA
DOdyIDJx2Z1fAJ3EzufJyXKPeVVAxMwGQLyL6EUyrDC8Yck0OnPgz6DuoQdlbnGB
YBIm/zmGNRdRsTud3yPb1o1xeegLEckDBVomZwbO/NlV1AVF8JAYYU5pSxzgYNwI
e633oQC6OUoV1U7qZ6chHYTfJLmIZUyWyjOQKuycZF/D/2Q3+aGG/9GldKAa/vmb
1ZROq5BUqNPeE11tQgWGdLCbQDHjVQb3bbPHBr6o4+g=
`protect END_PROTECTED
