`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5E/X3tPaf+GrfsQj50EnaAXrylWJgm0wxEmDlDbqF5HnDkqXQAVYA7wMkIUb77FK
tAQ87/63OYvhLW3kg80X83o9N3I0tx7A0uWB6r8ikk8rCdQLgyMThnpxOBGvRZPL
80/iIgUrIgvR4KcahOq8WNVunqPDayqURGC5m4JPRIl9SlHt4gX+6w3s2uIP977g
OLl/hEVTgSpWrwO/Vs38ab1GI4kynvo4mx4x6EzgGr7uKUZAdpPbKZ+WHk5WoBiB
XSo6KGtEiX8PIqQEPn91u0fYhit5V62i8kMbXWGVr8HIvMt3TDR3MpHybKqTnqG0
0I3zBoUvdo1HltVp4dBYSKQrRddiahrmYoVkvbmAdFcp0YRsmRlcdRSU5bs0puqE
mKvO10k9PsWEUhJnQgehbYtGTuHGsKp8ik5Oh8DCEmQwffTrBToJ1TeyoYG4O4tw
lvOIQRRNrYNaDFtDkcSFmeA5Dwfu5Y4i3cK2zqnmBrDb04T1BZYV+bb9XDn7SfYq
hKN4+QWSQz5kP1PMvMd7DWAndcQW6A/sBd7t8EkZvjEvJG8UghWKOu5kZQnxR2xh
obWV/TwnA2FnrojDtL5jjhxFOS/gcBoblNM8iXlixT4mTVp0wwhpQ0qQ3xWo57F5
7S/mrf0tGzAH97ye9Znx0E6TfJgzmrGLqrctQOTmPI9dzNPbw85iznW+k5EZ0fAC
SAVnw3dqubJTygMBNCrHpNPlW75obsikfE8JqQJAMDfm9JkR1qeJ1dcJMiIq5CXv
42lUFS8psiKW+Mqj93fXJQ8/PrXfg6aArbMWDHTxGldwHveOPGmy0bePoLXgDesR
2HykZy1lFxKe7EvfFM9ewWbPej4cy3MB8hgt7W2cZJG6tnzVQUCtfRQJyj6wvnvf
uy9s8uH3/snPUtfhUfZ/JA==
`protect END_PROTECTED
