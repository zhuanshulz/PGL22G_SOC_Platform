`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aCHreuMIt3zyFNEW2E2sbRvt1GuvWNiAz2Qpmc50xS8nRgGJvtTTZ03Ob7JVUzhV
i8xiMdZXtuN43NovpRxJAx1LPGaknpHQoB5REsqgdm6DhqeqesBzA2wsS1DFD3t2
20++xUfXuQwLjiY58eT854DRn141zizTpFH/a8TLQEEe/y+W0zZEgzjcrprP9pB7
JwtsarbSRZ+Riwmeh7RYUCzexR4gBwPYdT0uA8lw/w+8XSXaGY/OUT+vkKMwd+SD
XExxBmlHHielifVpQXM8wycBG5kTJNe/nppN1syTYw7Q5RAe/MGBCZ67VR4e0yrD
1FJeQN47Rpy6nqJMpZpX+Npi4bRatT2UEPTIA8vWFTyQNIJfGYjgiJsRB2VMj9fi
oFg+9rgKr69xFdVkcr2Ar69a4P5DdDfy0vs5fC5DCfgpUL4+Y1qYyTaovf9N/b+Z
x3VRb7TeK0Od62WkIflrjeTcJUNTj93w3LW6np5AHjZxS0WlzurjkC3PA3KOYpvF
XkmNw9PIe+OqutM+P2vdOu9shyxMfF97XICDNonkRf/st9LdI4iTjNaA+TbvJiOB
F7ygnwZTMAmQoEIKfTcgA+S1+G2bWYCF1Rq5n8mtk0fBxX6whBDaLbbBClFoRVT7
RYsDRZQEGQtrkFswO9m/zfO4ZigfgP8C0Y23/druI8K5DOUDB4ychRSdX9rIOd3E
pVQDGMCX/YJniwklxPRsW2Pzt/32L/vFCiQZOKHtajeLtimt4hn4dJ4JUtWnOlzL
`protect END_PROTECTED
