`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onWE5W/pGaCrZdrJ/Lq+YH9tVXqoft/VShkYUIZXuJMgLDumPRWb1ETMrckqOftw
PJI0TcON//g4rsdnaxREDpvKJwTeB2ldYJjEZLuKXVsfmwaVCJfbLUtsks5JuPA0
N07IxdwoMJOjP4fy1MejEAwEjGLnqDjUzogaaORJUNpjeAZRPCaRKqa86w8FzYVt
Jazo4ONigtBLWWcnwim5AB7zYiw6Sn/cYmfnXj9HnqYh3J9yzLa8vRhYn4cAqt2P
anHBExge4XVdbf7dQYH8pA+SgDfqoRnSuAcgsJvozYSXV/JCTr2icjIDKuNdY8lv
+tJrFNSkuHCBIvE/WE6T9p6cJRX/adCuDCc+Bm7XLUGpJkDv1lgdojPQZTDAIaWm
lvmDq3TUeY5uyjJGgvjvBu2hPi0rFpHvooA3ZMGOAiBkxeRb4RqUSaDSZ161yE2I
oZpBLYR9e7/OY1kwymrNDa8hbGP+paDOSY/nx0sh+0Yym2e1JOY35xfXPzkK1KeC
`protect END_PROTECTED
