`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2oyeHtNArwpmgSq52AA8wlCzxGqcwYs/swYy7L6Taqv8UOL/lw2wh08v/lcF8QDS
oZCXks3zEipLYv9kuqYKNfmSLRzjlOpe3OJQoROCmkNk5/Q1MJKbvkaCiV7HT4/d
0ulPchnsiusfoLFrTMYpJwucGTfk3UsNtHMHADlXo6i5R5sdvFgKEVOhDJS9h7f/
wdaUPmoTSMk3muwZhiMrXrippWQOENd7VynJZcCyptzLiQ10NWAEx4//GtS8XDhr
zB7VaYRAxpVONhX9UL5vWjR15a7EKtROKGMmWCo6mWp6c4VWcrO3GVhFno7Roc16
RVJ8CvX6goKI38etJvxL+GMhS1m40g5RbdIoaTJc+q4G0aPvpG4xe7W8kc9+9q7M
qNK9Kyp5N6s83qS8wPWMBMcIB2fRkY2OjM1Eq0Wfj8ew0mgisUNoRelLDOJBKwr4
6lAv0srQe4Kkn4quWRbiGg/2Cj8cl/n1pCyAsulTU3bZMwGrr2nZp9jKNlBQlmps
64bjSGZG5zwX9cQmg+pSISYkCkpVrB5vIf5AwFaxFKPAGLR6fuezxlBrT4AhRXVl
58ZTHjf9d0Nfuph8NWzD8wcr08IrndhFBlrk+4LK1D+839r6S9gN2Z1sUkGmb17E
`protect END_PROTECTED
