`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSnTbHG8LKNNd9+AruecciovW+x6u17TqlO9Ta9hScQepgORNYcF1/ptbYXpgw2X
v3wzxO2wmduCcMjkWemugTI2UzWV73461gVgjEAqddnR4Vu9IvGUTmC1SABucrst
mhiSOfiHLtOjBG1NLywu+qtadhaYgymcatwOTlmKi+2BcVI7vUzq8vZzKtJ0x91m
u2QWpTeZmPkBeuQ+X6ZRoY2CkdyN2GN3QcHYSnyvP4paGm/ITL5ApyAHJPAzs2It
sto7V59O9u+SpinH/L1sBQ==
`protect END_PROTECTED
