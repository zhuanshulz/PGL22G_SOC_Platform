`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ohg5kNHPhtzmQQnql2LR1HiJuHqgPrPOS1d1oJzx8yLWwPJMoWdEhd+FmgMSpFR2
Mh3iqQr9WuYRpW82VaFUq2m+r8S+rSpYWBU4dLOOy9LxdBv/1z/L3sQjXwSagolP
BULvds4APceCKxSFv6H0FTlDWatfCTl/VGZUQFF6k/Shy2CwE676UBT1DWdpnOG/
Yd0BRlbcvqbFHKUEO4/4szV95iehLvlQdKBRS5pwJ3OedbvgNGbKBp+lrwadTBUh
0Nyu8Cp8xbE/7di+Uqe6iz1s4Ex2JcQfchHTRWpItSJu2hSod8lgXwsVpDGss2ZZ
yD+oKmSC7CfxZ7jAHkKivmeaV/T6EEFaF3AkixT1xKIlJT7akzrReKeV3hn0fzS+
qvXhLBtlLuWSBRZhOGfv7r92CQnf6GnvRKfJ2tICzJHGD/kDvnQU2sE/zwe73Xav
vsQPm5n57vn9/2hZGm+Yt1t0fFvmq+DVfEdhDA91NRUt76KRiFLVhZbIl+GOqDQV
PTxzv1NuSE69Yy2shS36zTOoJQFPid6mhPxLvlGMpCKabQHZH7sZByQxocyN1g4R
bG+oINYSkxCAUcnFLIVRTxxYHO7xz4sPaGDtI5AvolLjvbJFMYLoOEXfMvzLmBmM
OQX/fR7ocv2ngOyNXa95ej6reK1BJFcAsUAykfXF6JHu4IMewxVKJAsRZ76EG6KG
A9caPR2/fRiW72+3jeUOABuwEYrdT3W9EM3+E6P9y2GugMYOLY3FoBXIEYg/4SFF
mqb/MaOynU8t9xoOriXLWob06etZejUyD3pbo8qGcBZDlREtrCYrqmjHNrj97d2b
UdVg02RriJPY7jKs9i1xrWf7NNBlfWNzIfpa/qii3aRLbJnJ4T18XKKLjDIwWv95
5YwwF+eA0l5nDkgV/uLboQ==
`protect END_PROTECTED
