`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LK3zNDKk+5kNp/oN/MK42FQwj9FaEF6UjgMDobtJGDc+jcRLvGWQYIZiM1mK75wk
XoqqKHlKnGw4HYooaCvN5wIve0OgLS95XO6sVEM93h176B+Lk8nTSp+tocRWBn9q
fZFkcAdHulLZUvAdPy/O+dsKjzPAMmOMhdNHS3ixwLFrguzp8ompEExmeanJHGIG
j07u9BkuFtjAOplKsQ8oS1Rt4QW63w7vvkm6ePX6VU+1zzvzkGR2DNRPNtsL7FTM
4odL/Q51ouOWJP3rwnhTFbQGpaRY3Bx8YqOM3Ded3UmkigZqW6OD3FzAs0/UwNYY
qcmGP2MHYnQn1fWd+cCiAK3akZmbtaLv0pibe/D3BmdAyAVWGXQ2tMQ4/LZCeWt2
rOexJ2kDUPY8TrRF5KWoFsVGjB21UacnMpnSt8x5SRC1VFcmeg60BN76VNaBG+M/
RIuypx+Sy1a7sjIxjnp7dpMAR8wsnZbTDcEzx2kxgO7rKplFZ1ECa50nL3ytGAmC
J3DkqsQNoc38/mcX87+K1CRRKB4m/IP8E5uDAXJ/rWkbjv0ClF1qU+WG2OwmfMZf
QQIJSQef5xJ/t2EmKQdrzaovxr2Bp1tYQE3wej+z4twQQkRVk8Tz4NktPmgz52rl
3SS0rQ0YnSG3peFjE8xft3iTno5BGYs68sScwFC7Le5N+rkOJh2EnTBAf9HhCs75
+wHX5pmtFmIjZvHJggFLGHb0ARxcj618U6nXxtRQ9Vn/7O0ITXYpMvE9SuFXq+JB
sqCLNlbGbv5tRC+DzI8LpbKssEqOw8yk4co7faNFGkzpTi0BGlQHnsr+TAWJw84m
TclKWPyTZQIkXJ7whk5M+fHf+C2zOJEqUpvDOroGtxFK9SolWgvrKzJZL+5+YjnH
DmGLVimCtfQeqaau9XiiMQUGO2SnSvyHRKlvEb8fZDJ/wGh7eyH3dEAh1YZkBk56
6s224fgNU/O6SUpNJHh4M7xYZECuRDnzl55sgHeqzmCrSI3aMeufmuRTwISFC7qe
flTyc9XsmX9OP2dxAYLWx/u/RCNuv3kboFTryIHWZWoR2+KO5EEKpkWXbwWZAs2c
JbZ29Nrw/klX3yrw8XZk6Iu2GFR+8CUcNznHHDI74RLEWSA8iTJZz3XPHHImuD+7
S1tvb/AB8psGJSk9X0Mn9TNTDD5wuK1FnImt1LemcTunwF+X2BIzMhBniiLGPFWF
Ptj/y8vJwglnQfCMh3qFKi/MUMMzLsVqHcetLw/WEkbuzDnEsDoeP0Bg0FT5owKp
IdcJZqYtTSv7zG8100PKbBN5oWV14LM0COiJc75jktIvQ7Ft/uflPwWTz+1qaJvv
8wCJMDLk9hxl9AfJdxFSx5MxMZV3VNllgyBFypSXDEiDmWtxTUFsQXpjknADb+6L
ppVIGHN4ZmpWy0o/CFoRqgh+uhSYoTcWdMj/5XlpLaLRyIHXDYQwuwk+ZuSqAVmq
Csnymo9bqHTlDHE0D4fq2aizZzeRHzyC9jCuCf+c/LXyybGZRP3BllNyiIHJV0id
ScFYEcNoBtJ80wgvKBqeIqLWFtWKqQR06QYQKk2FBlsPULEttqbiTA/D5gAH7J4R
ZqgqtjnqvJIOQvbtE+3vubo8AUbFMyK4+YNQdp9k1pkxo+AbWRjtSumakFaYgaNf
IRbIVhzHQOVsHaExdNCiXVnvnZa8tmaOLz51x/1w3/j6y3SQ7eufqJ9cCbfgsPRI
TiuHE7KqpowXISJeOE1vCRv4VQJvwohruh9PUUGdlG7nvdvZrqHCt3wlHtlD11rO
IELqIb/ERuHDLwkmQpNUAapWLMdtVkDFTlGmZoraugpgvUS71NH8I06Qxv/+L4X2
y+7K1fdhIwIMPHD12T0HM+kvcKbCZ1dgvSupoD6X1Fz3vvVBE48VoljTf5WcyHPz
94r/Mzb0wCmOGCPvjYKAJ8nQ1hh9kQIwQOh9ulG9wqiNJFu+hTdSH9KtxsYHdiNA
WSAj77HXSISNj6oi7sUxNA3LNc1meqlFAwlc/Sls5nuRIpje3FniKBhH/ksPTUGN
v53Y0yjI5+ZD3HptgrrbZgv9lsy00CzwEfKrFOQKo1YUKRre+rYqjs/Wgc1V+e/X
Nq/1k8mCpZxPWP6BXitFqSzWbe61Q8ibB35dCHnYkFjlCNQjy7eIc+xS8+RhUoEA
1GwcliDYk50LjUqDnDuBE3P3BOGjVfw9gwGL5qwfQWMVGRzHB2MoDz2d/e5tuvGm
YVvTuoxQ3pdibASQzYudDBa4kko8/Xj5hQHRDseJ/kS1mDL1H+FYOqYsEpStKf3s
ARNoHH9HmWwfokLx5Na1VczJggapEO9axJfD1YOOWE4zqa8C8dPdWVx0/FbULYFy
+Bdm2a64R4YHalpAAKbDsad7V6l2gmXkPHp+ze3KiIA=
`protect END_PROTECTED
