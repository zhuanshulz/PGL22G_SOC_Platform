`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SKgm30OQrItOEoJ4qdpqlh5GPK6z68yMHwEI7NnnGovWuzaeWhb4WFL2mmYCU2dV
X19CVyRuJC2qJ88Pdc5iC1dH/aiY4YenH89Gqx+qKcrHdHSrMTYwOfqmlekc7hs+
tE0ydJagRfWFtf39EKIWJeTY1Ua+/HorOF0Em5bEjDuqlKLtlqAAmTWiADFr2vmh
sc/287BEPhHVrVF0xIAyvFLA0ea8WzoQZK88XbasPSeCcBXmNKyXekXh3fjAq1Za
Le+VywvaOPx9qCFQkuqOH+mwCDOjUQ14X7E7wtnoKtMRraB3FIUUG2edqXZvWwmg
Um4O2CmW3My2uxTjScvpl9MsgI+orW8/viRZVViScW7nWxn2zKicMQEr79jmF9Tw
IQz6mLZSy8Dy3VDP0uUGI3pcm3pP2/a5pDHJnpXpYm5hrDLovBTh5W+cf3959EPK
HWlm3fvtDX8AdaXRzFW0gqiQqSr5wXXlWXxMaTqCI5rLqAoxAXNer9wlmMHzezlZ
ZzEguAgMLcBgPlOFCeip84a3uem9dbqvo9EvUniCGvuK1VPzXquSy2mdb0aEbHFS
RdHDyXOaWxYfl5PtZaG2e7uZOGakIdmxi3W0SGcRK8/2MKAol4BzjmBwSK8igrRD
084lr4m5/z9QJwT8Ir6ACWti8Ks+CQ8N5Vo4tqyY+IPu10YXyhbdQ/WI/LO+c11O
gejANCun8Kgda0UUwFIquvJc8gC1xRB//cQAX8J9TMlIa9XDVFEk4GyPA2b7oAaD
6NBSm8rRgD1q25dRyCNVgQ==
`protect END_PROTECTED
