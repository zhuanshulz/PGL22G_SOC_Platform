`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpdKbc2nO6uUWXMRRRYbO4jsm5PzBAE03SGAVMbunr1PcZ4/nLyeS1ynMHm8Axpk
KQ23X4+tt0rIJpaPgocVvD1t43C0vnfufVYPU6EL1DSGD1JCm+Jv3ifsi+O/PA/P
DUxw9khW6pO5XKjFV3+YPO6hXqa3VNYDmdUYXKXm6z3NWTQvQOrxGHSSpZzGiTOn
kctd4OngsFPAt8bbImN/95eQnKmfCZSmsy7wF0nkLLMRDkGiyfBCrGqtNNa3tKAJ
E5348g21qOR2pOF2dNDT1wyXWJ1s7dSg0nqUSgUr8xNXxBwJK158hs4k2UJauujS
+65H+B/XBmP2YNzt60SgsgxB/iBEJQT9efK2PDq8wCEbTRjSwKY8SvrYSyOC5R5q
L/+NhQgRYW8/EKCwiOUpw8TlJfjaYe+Joun/V0TmeAqQ4bTNynmEkXnSOzRt1R2Z
DDMG1AyKQnmcbsfXnU2c8CYkkWhVhCPyTqSTT+7L3H9/kOmduytWEfH0xLkzJh3P
p9zFWFWQXCCkrCEj+7q8/2M3DJoMBy5gC/o7J2/kgFKrHoNkPnUX1LaCL/zCmHYy
0BjnSbWYIK75RcnuaD6G8Zny3qrT+fyAh5WpRuJdKNm6fLaaOKHA4rPyAI5KBdzN
obxpuIvhttZfqhr7TDDygZLvzSYxfCNPMW1nrHjqsRmwC8XvTQzQi3GoTuRTqbzc
9Db4PD0KY6Yz482BWwcJ0kwTJZ6U//ZraaImwAoh4sZFSRJ2+0OyvVmLbSt3flEf
1ThgF7R5Cm7n6Zld+AK9uDriCl7O5nxUnxAqWYUcoDjJ6HXNvMWx8rb/FyrCTRye
UTOfzvL5tlYqev+OpN6+NzC6czagFhmVyMHXlbK2ap99KdLGqdtO77REsmZa1v0S
WJrCI23w+Tlzydt0NPJD/2U1A2VSm7na7cyZKLg8tqteZTjvI5WUUojJ62Va6iXT
051y9noG+EQx/h1fu+lxo3NFMEKlP47vIK9e0YakYEhdOegD/9HPExpu9Xo990jN
zsp4pYrEJApTObjt43I+3MpLBAwXbEcKK/zETaKNnAnKgQEkdf7SpYeXGG6/bypq
miUleBZ2a8HfMyUyJ0NG0IKaVhCe23i8JATwEhU/HPQ7ZDVU+FWrq5eCLmgGG0VR
xkriRR0I9e2AVqcj0au/RvZrh091nXCfTRWIMMEx6pvidRDZswoAiY/NvABVLe09
xSJYjk28/oP5CUOhSH0e4kKAEJ9fN3EUv6P0aZHyHKhFAUEuunDYtOeXfDPm4D1D
l6j3YCLs+ngVhpL8A76x21Z/hqD/SzL2m4oXGSGYqdAZBNTtWArNdREB48BEKiZZ
YA5b3VgxF3PsYRvRKfl9Sug9/dmwUESCb6c9rFDuokPFZ2gPMZ8psCKNT22FL6GE
LmdbWQl3Cjipv/Ogs8/qTyK883nuthGqdgTw3pAPgzCrM2M03b20eF8rZa8SAvRR
o2aDF7X8xk9krH1J6diR3rApqkLh2U4hCRmUTugWZD/jZVvu35YC5JyufC5tJjlt
LT72pb+t4IXVvAFCVnHrxgKooVcHitk2RMY0CXM8Qbm6sT6fQcXsfcNeZZoY4iFY
YplNIP5X/6g/2dabiWaF5HJqWzdSxs+Pio6PBoTTGkvyu7QXecK+YMLsrwIvMJrN
t8fgFllg4HSayrnxNKepHd4+Ucuaoz1OhiPRJ96JVRz8AWKP5saEyDLrKpIusW5V
uTppYnjnhpcIGZ+sO57eBJvGs5pbKeyiDCs8MBmV7FpYnLbsKGQvznlxgd1Q/iXf
0Qu8qcqFVFUNNyhhmqHvH7qOYQdui8jmvXpPFq0ig61v6zTQheXna7P+2UpO4Mab
KXbO673vvioXCkgnfsemuKUuvMnGplosM0aD+i0X3X36YCAttv54NzZMHpunXALo
S3PrqvjZzMjhpad4qIruBr9oSvH9Nje4IPREoR738GNExdAMwop1lVdcnutYr63x
nXOYea2fTP8TbX95Zy6Q91AauF6pgnTmsKDTXD8Vo1nhzEcapzsLQIIY763Tc4PV
04YAXthhp39L6PPuQJyQesIZsWc8vnNlrq4Rmn1S0DgABg+oMoO1ta2W64PbQgdR
Qu8PA9IC1WaLDLGP7Gk+HrBLafVjStcxrd1n/hJVZX0M6BTVrgBKkPocJQLCnC95
YFq+CI51nN80+1KbLWyUg6/c3B6kgD65SMY64dkVwfiroDpyZOsXKhj2wC8kruq/
H833Z4XaDtNwp4IuWZg0xHuDogIAFiZmmJUMEtpfOn01DhzjhR0wtM3kJMbee8BA
8kmODiLQ62zh+cJ++ri7U0L8ijkdcleLjhuOMzIwHheBLPWTYsGGKT4mxuTxsbZo
c1AzfkeQwPW/FQHPml4LmnZiN7RYjkNgMUXMI4vDDqV4+8yItB4b/XcYE/5EasLS
mIbLfWwEJXvKvHZqR8KE8xlij69IO1RZUQF7FUeb5UIFN9xDmHvRKm5OQvE3jJMJ
pLfANAIHjKY1ktn5CvZXwGgYZPiChdqCHoauxa0W0vZrnFmRfppkEe7GfuPmO3f5
MzBNZCZmPL3x7zamkYcap1vyDw4y5L/VddYSlW8XEGrNkQFOtsMSD+oF9OgIcfVF
2cSNWBdYevCct5q46ttHppO0vbHmLBoDsEjfQKnj7txYj3JfBiWnqk+ALYMsRYkb
0iB35iBgjzgx8ROioh7levwg/7E7jmHJzZxL4p78CWolD2DUK5ZaNEEIA/edr8Zz
zo0l0/aSgkCxE0bHVLK+w6gQDTc24RGhROoZSIWJdlOC68rGLahuA5Sp55138ll9
7Jk+7OKr0aE7J9NFEsfDEylVmvJSF/ZROZBkDgoW1B0e8ZbT1fJno08q3nJ/RHW8
1NIQur/nndw//3ATZkJ25ilinRP3dmRkHUhqYNjOJCIkKFPjz5V2LLHX0aScfk1i
Q1OC782XKSKBSASZPWJZeFOMqqh3YWjtqprSUVVEOmepzWnubU+vyqBObwJn+bIW
Yo0J9Gs04YwX14f44Ho+O/0IKxr3xnPo3/sl/2ec1v8SR2z/gLXs6ECOle8t4Q68
Nw9vBGjoQbWCG6iUAmaqM3JbNNlvwNRH76AobXhbavLOTYmPjcV0oFkzu9Tauw0v
MPU/49CwmdoZCQXBfoF7jrmE5jxUsxehjcYUw2ojqI5QSgKoidkv/oz2tq+8qqOw
9RVu5FuBsQI9uNswEQNkffMHT5j78M0yrjCEbdy/lXkOW1FRVrTYHsOwbjw+Qaw6
NXoxAz+Z14Nu9y1mBbX5+suJ2HG2hIGrG2TspfqtAsXuefXAGmrI3uRzi5TZ9sFQ
k3wYUI/8zd/YYd8njiG0evsYk+GEmUju0Xb8XFx+k/t0yqga9ZNVDyHSnng6wrjB
Myqvp71JCdIntLi/Q8/qZujwiZygbBAQEGRNUjceVhpTc34Ot+jzgTE77O3qIAQe
znww/3dvR4poUUiA8vBbzhscx4IOlR2MyqpAfxKqEwvQim9u4ERW6AI94AJAAio2
0eLrLVg/FiO3YImAxlm/Jl/UchZx7vGsIBoEFNwSuGlG4sQLrb5Ei4ZHrTFz3Npl
vIlvMwbrAKTmW5uw+pZcikT5B3DWjNNw6sBnbzLBXDQxtSQpkDP0xt2M92rMW1Tz
83KLVHE0nkxWbUGOlocIx0XfwOaU5b9eOJbVrW51EIv6RBgQrMnsudjHGpxtOlp4
mWWeWqXHU+QhEEOElHseoHy7wqLqjH6ka7aQzO0fiIMHVriiDMaO5SEbgLo8XWPw
wqPw0JuTd8BRMvkWzW14vKROM83MEo/grpUHQPRb5IeFJJlBXWQjO0UEI0Tn/CPw
JUUwWZptCb0qab11Bm6wQ4yApK2OdYRzvMCNhvdrv5l3PtoDprCeW5jI5mviE+MB
Od2819lYB0sShcE39n4L1tMZkNft/z8D6rJsmtFnuWQLWAzpFu1BHCQJuIfSYnbI
SST1t/GRfCBATC7vl1LOX1wEf44a6VWYXeiXNOGoktnkXXv1mcyPbtXUK3r+002o
ph2i/j9LMK03ERSCq1cheVMXqcKATEeFskyNhpdoBVnJgLbKYC6sa1YJuVwqJZ8B
VxfwU6Y+GWidG5HnIL2FpjmNbL2qoSTEXCcEmrbub15EK82r95mhCwS04JI+8NAE
4eAeimKW8UQOup+vPRZs0b4cFFldLF6hsyDHwpmU4fmkjl3l4zJ07+qxKr9Mi5dj
6B7TulB8a65F/fK4MDDP26aePkxzYYURaaa0hyLewZJKWnXqzu6BNRRvjOAULcdP
OTNToL3QDQwnyQyqbBqsk7eoJo9lMNR8xm0VYNkxdDH4R4/Nur8q0YJsT2ko25oA
bCmZpw0368dQIzW4uUp6S1qsa9O7z62UWd6JoEDxvRMFPG1yJz/py5BvcCzsau2k
4UQ3tvLGb+Uc97B4RgkxgP2IfVDXQyxfsiQzd8B9J9PqI9/siayh10SrilyuWcJ5
gL12+LAX7KMFs5VNa1MxLuuKMwFhOVlorWCUvlsiOWRarV22Jcd1qNDhcEKwDhN4
MlhBuZqDNweGc5ArfgF5izb1/xpraaH2Hszy3QLSjZveCsUXAUJJ8G8oH1hepdSd
1pqaK/txQZDf4JL9sKhPSOpZlYRgQUoDFreXTn+58SS6czXhuRjsv4RrYPSPj+6k
4qhJaUDj+X7tDCTR8LtIpQ4ndL6O+5ED1R5ND6EKyWvrXHvHY/8gxqJdOFY7Cd7a
0BpJqooXBrq//4bzmgyRmV9qARv2CWfFw6PkeIGJzBQXygcdkIsc9vnn3oNpQEfJ
fHXzLvX7DefvDSDYjx/aAtQ2/00uMUu18mBNcr6rIb/CtxGlrBNl2KF/soxrQUX5
t8qt7PAB0Xxa7ECoyQIINJGiIgEWlXTqWGvOrQghf6zD2dbav0f4zhTPo6nvU1O9
YsABKbGR2pxY4ERpwBhIogXhngS4poeddFDfJKkb+l1cZL2FuP/JOcyIdDas+C+a
ulvo4uWy6L6Z4SYFWjjQIWaNbnJll99p7zHTIaqakyY4VaUdBGseXNB5bQngtdO4
cx8ZI3mS7jLS1INkqT4nGRopNz0Cs4aRXrhunRq6ZWrVdkN/fscfLVmpZWdg5bdX
gdOQcPJlkIn77dH1BfxYdfIz900Iwh7jPErkhX7aUSugKmDI9gHNIzmwV7wvwC+9
mEV7szlO8Dp5QkLaqC3uI5cfTzJMtX50ivRQH1EOKlL4oKw3xebZBY9cvBMS+vnc
zX0tF0XCxO4Fv0/+pYAhF+xY/wlepXNyWV46mczzhBPJUhlShQKKtC1pG6cirZ2+
UmK0UU0CVcpPBW6RIjhibOTwg8Mmkjw9q4KP46P2es6wcHovKTwzBv+e1Rfi1ApW
z7gMi+pulNFLzQmUJMCbsW79McfrMyYWANDylS9iir3FiBhHiZLtM0ScI8LUbQji
WQyhCnVFDvFsmJ8GGfpolcllFCFzNZim84JBz5peoQYdDCHut9kMHGuncm66iqSN
uJ6dOs3WgFtfM83EsdEA5Qbh+AsRzaLLtErEedd6jZVnlnwt2+jKm9Om4iE3H5ut
hl8dKkXYAVCxIu1I16xvcFAlIwaEjeO+G5rc86OMf4BSvMSyWSnTtVthQp3dl23G
rj8fBgLxB+Ixlm3DwVvco/zsXbbMqqbkxTEU9AhwS0EA+l9LH35Vt1+1Hmio63JC
o9MmXWQS1Zt/0em/cFgSnz5KrGdkchpGYegeNHINQaxe38b1gUgmGWDNLu5F/KJ4
NDOA/99KUhS/ix8ayt7WUm5HQ/LyC7tZbGSyybRuQtaPAyHuhUHENSBoMGs6zMmA
WOtIYip4MP96CjAp+zzyvI4Yu+f6gHBVrFhOaCs5rLn0/rDf5YZlwuKFrxlLWtIT
uCXNpA23p1DAz1zIRBTD5fg68/rO+21S4ZfN7F/qpqDKtaZys1d5sumtspBUmgxw
j/4VWYP72gFFNP+HhznWXZsKWZMbCi3Ecyii5ekqNJCtmw7o/FeBVkc2uVmvoIJw
8BcTJ09J6sPrgpMNwOpDOAHg5NVPIeZURVAljyiXoyPBfKzttdhIMkOQYxNmhE7W
HNDbib/MH1GM6sFwZLpfIRIRqLTciXgrVG8jSDnWyUmZGkL/Qj9J0+1QY2FcUXb1
IDVzG4fpn4GHZCO7L0c5Y8uqTtiFa0vAvqJyJSl+dHj9sFUn1S0Igyqimc8Pu+fG
CNKUN7/DP6Bsl9HmW7TWEhaFT+7MUtbNcCdL3hnJGmAm56vCEOJLVno63eqfPBv1
nFiLdSUhfp+oj8Z4+7P8avwKHKc8g3sN6kY87OkZ7BCZbF5idSX4vbIZFwiA82RW
kPVnK8FTgmEBC4ajLITfaXh2FJSf3OItz4QfyKjj4n5jYrOuhXh4SAfx0cJAiNU9
lNok/d1PQBwcYntmFl+uPGtQvCppxTpiJoI3wQskAml955/NHPhR6AqP8NE8dQ/W
bck/Oss2KVj/79IcRZftbWYFN/POSzKozlJdIpHzT+w/5Txb4CXLErELh3qNaVwV
pFyhj7dybg/rp0eVClhaOAIdJnbImgdPs38O/RIUyV4LnTr3wQdMjfHVtyB0yrZ9
0CKL28gwaJBNrk5eYCvmb7wLIJWK3tOLSg8cjZ0FtSSXzjelkyKnsN6rNo8NAWHm
v8qvMs4phzeZZTFMCXDFj3zzGLrE8k++k/Gmg5ex7dblY1rqwav/znX1B1zvEIV3
LLra2NXNHxNzW0yEsexiUJYSt0Jcgp60MLp7irh8vpHOz7KFZqkudWqzBBjZ4/Nx
rZkGlYTEhUamL/lUf/mS5dq0L+FUJKjKOc8YT438qsoywIxC669QmFNnpyYRAhSF
9nlew0v4fdO4AwQh+kgxjvG25G/eD+qUZt7cF6ptlQRodnCOX3UWaHOua+z3Z1ik
an3m4L12zZgCmrlaw57ZjI0mAm20+4kcWyXRCC+0NG/E2StCutUv/5D6cYWiA3+8
UueAAI3u40mPwgzS2p9w471/gulhEUfyS4XLbb4atRWDSpvqgC4j2qx5LutveQLj
VKBmjqEiFP13oddJhK/1aLwUl9R1TFjw4mrZWc7ZoEPR6kBMQZ7uoRdCCqliM9Jh
kuVNjpj7Mctr8N/+u9L3pUd7efMr2BbTC2AIPmNBgg2kmF1voP7F5ZxI46dyd71p
whIfOr/CEBUQVvBgufV/XJpHAp1lwnl+Q0+Krug9lZ43q0xP4gX+Lpv5RNrdc8Jh
W1NRPEN8ctQ9bwlzz83UOTrOjFxEilIlDkV15rvzeUqFRHnvuavwl41yBEyB0ysW
wHy3FkF88PTAXJ9tOnmwh1oi5I2F2C/fxN5Trf0SqcUpE6hPG7VL+mrqQsjexIQK
K977YnjKtijtOI+i2QlbchccHck19isdiuN18rWex2ZLo2WGUX/ycyqFH8wLRN+m
kx++//R2KoVcmgywXFk3X/pG3K1wfJmRup/h8kGZ7Mo6l2/OK3GAqf7+DQkMA+XV
8NxmcctRNsJ1XJfEpuvLqHSWgiNVkWlohu0HGd1QIjMEgvrjvQgIOon8EjrdBG1s
qmad+GaJ3E8ikk5U8Cjs+dMWcQrXYWWwCoEm2M/mlnFKeAvY+tqH3n+Kt2pGFHFN
InFdTG4X+RbkR/ykwcWdyB6hxsJknwHYZjUokxzWSR/rW1YMHyaeiWc9ltn6AK/a
bQ0QNgWP9ltdy36koqVgEAuMWky/rEEu2HnOKaA/b4SFTq7fBw4UTqTmp4Wiaw+K
QeNb0ZijnSGu/SzBtqUXqK7bp9kG2PF6SATndp9mMv1VO6rjfAaDpvqMIcUnQDop
XE021BIb5L7JctRlrlkaBO4Pp3zK/OHEZQWKr7Z4uRJAvVtJ/gDb/uNB0e2QrOwb
leF1fP2zhE5ihZXBiWhjAuDmglUIQbIc56vghwf7iq+xyRY2jaHhRJNERXG9dTzG
JR/pxOswE7cfTeIEUAnFIL4OC5eDzNtL+hw4t5HYpRr9AxhMS+gCdqmw/Xy5yhhj
7hqmWKjL8fxPrY9zGVQ5CYvtYDPg3PPg9UuFd51yfMEZSHMLXNpeEQ8gNQvLUqGV
4jc9hY8ebcrt4idH9MX2CCbbEqO2q+ImqxW8XYKS0CCUcNn6bK+ozB1cCvPS7/vF
xVp7V7eo8lsk8XCQsfkwHk84nqfk/VXMP+nXUFcKltrRlXsG5lECkDpyA6cJyUza
ALqi8U2VQhxJBG8H2sUTr4JJiiq5uihMqLCg1g2ks+SXHsQo3INKmCsEaDYAvEc3
NLrKXCOPgGDTZoroLhKjBbulCxQ7Vn75IPavXBFYuMq5P5jE7XBKk+E2zSTS9ZZx
hx/AEDQzHnKallbzANzSsga4wPt7NuhWaE0NRvXi98/roOSJ3RUGhPny5gaaIzz/
rf7g4TOHFQKsXE/X0I4SyCqG9jzeZ9CL/Adt1w9wQb62yVscM1Ub9A8IS0VZhDVg
ZLuYQqRujTCecGKtbsVgNJnoq70RyrqXtvMv05YHqpN0sXUX+yYYT2okhHVKs9X1
vlaxf3Sq+xaoJEKItVOVcTGkxgB47/2raQbO9wSXjaKVXgLojY2oBECIEgZ6Q1J6
BiCqLuZ/QeuBEkdRoWPfR5/rvJioVYPeKWdsb/EPuqOsd2Hxx055C145y+sLpDve
ECwJ8pai5nd6trot25Z/MNGsmY0XfB1JbKeZtCT68xlYqinLNCc2nNxBcTPjkj7E
Tq3WTpleuF+xRwgWf+jL9ssqUXcMdYMcXheZPbGWgE1g2rWdEytZJn/XXkSbbgFl
0kjjaUbw1VVj2M9XG7WCD/I5+a5Q/hC/3tvtIopZB2GzDIoOUI9LxRoyFASVf+o+
p+ZySsbUpwhLOuEhf3PydJOVnX5Vbk0p+R2za/ouooH7qo5ZIPM9oQFAJ7H2HGpI
D3CKGi5HIom0HBxSponBDvBlQ1WKFQA8A2Wio7DiHWZsTkXorNqHCYCBOFjzyHyd
N2y7WwuoQVPxfJMfelljkolpfBcF/1Z3Dvp3GZj+0OsHZ31PR/lU1F5s/YCIgdvo
oT7++k9E8V2oNkR4RMgpFLj3xTIKWua4auqMUgcvfcOjIcl2GrX4macPT+CnAFcN
BrejoJj212Vw0z1CWUEI1RaEW58eXbt9rbiK7e9oP7hkNm6ov36CmuV/Zzmt/OdG
IF+spzRsqamR0ZQb7APeNwgKm1we9rhCoYheyGdcgtyQWRd3g95ciMCoY/lQ70q7
J6dkLD06aN4BxGyJMDzDk6XdkiayhKergs8x4ZpsoC8rkuQU05jp9jc2cYUhT7JP
IEm+y6JLQItlrnhj/lyZrwR7UeHx+10NuwWgwakOcb11bK06vUV7Opx9R9nVlv/4
4xlXpicGBMw+61viwzIAovOltbF12WJFq7NAeCOi0yXGOHlWFlxcRsZ/Jiy3xqjk
`protect END_PROTECTED
