`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+w8XlUFUFvTkf/AfK+9XO6Guhy4geVcSTunyIUhba0jY9WSLG7PxUyZjq4ndK46i
jMMpcIPdrXT8o5Qyl1UPDOg+BlQpm5748G5oJl8RKkRGyl5GIVoBvJy9NJYccFjH
qfrjl2TuMHmQE3WMCLSF/Or83M5a62OEwrmIneP84TLe/OOsuCCm75VmZa57xj3Y
Q80FpFdF+rju0XF+amW/LZi1BCeI3YS4SKYeETszBiFCm5n9+Ntj0JVuqSQE9evz
nL2zXhE/ua9ubtju3zovmE5kApm9vHHPvUzu4fe7CmVTM0A1p6z+CcKqgRvLHYyA
EUmMsSdjv+67pNOjAoDk0Q==
`protect END_PROTECTED
