`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naQjZHuEemz0QMY7eowmvoUHTV+pSfyi0Mcn2T000rEDZIEB0uW06g15oQZrKbdF
LKU0UEQZ1AeogeRhtyk18DStiWvAyg0+3huH3UZ1hn3gcAGjXtuKUxTmmbVngZBJ
z+Di2BqkTIC+f1aGHne24HTmqBORjt7esdecLEeo2lqRJ/JJ96zu/vpzsWXUUk9b
o3d3ArSycS7eaQG/IBoY1GytSMfyqDuOPMmd42mMbo3w3wOyRQmfAuxhYc9cp5rZ
f8ctHjNGbak8nEJcOacUDZi6UOzmJEX9b4UCJPS0BL6DJJ44TrX9S7rgUzcmPdxc
Va5aLVaZVIGPFHbGDWy+gE0turxTk4PU8s013z4K83oHj4W/eu9ZhCKq3rJ5YflL
eMzW/2jYzHC0GuT9ooTB8YBJqi0YDrPIfn3Zvp6+ad+4nI1nI2Cbl+ZSggeJe7E4
UYNMfhgEYpKHGoLz78r2A4Mgyb/LGUqVVWjytXNTECmQenz/AJn2kASR8r/JYscf
880y182mDhAW0j6t1nCsuA==
`protect END_PROTECTED
