`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0AzBJ/vzKzUydwSVGIkUqZlB4KOaEv/tOfAGApdSgLuXuyhJfmb1P7cx9uRHLHv/
L8r7cVwz7StawgAZu4dwwRddkgO4Ls+f8uoyQZzqnagdc9buDz12f0JPADuncvvN
wbBUXI1KgHNPSWB9Y+Iu63wCkuaz7cPUHQ0yxMabvNQenWTCIyTnw615IW37LRKs
WEyUp/1IdwrG1DKmfO46a24J2hTartto5UpySN1SyPCzGp1pPrBO1d+kM/KqwVzJ
AF0cXOU5zLhLc8XE+5vfW1VgKSUxQ3JnhCNFVf3FyRdoX88mb4Wp71fZOe3kxKUw
n8Bsago8LI83tLwTNs0dm4TPNRoMEWOW0clVSPnzEj3rICG58u08+xZbf4BKtms9
7Bcve1dwQ5Ym1eLuvZj6EtDBGoZrjtVLUfZsNxv922YIcEhAjTYpImo/pIVUVMtc
NSZXVDG997HS3OwQ23O6eLmNby0M/QQ+TGn++mX86jQAy+lE8A0vMgpEUtQhTQNC
9jElFgIR/UUYQ1GzxMRMtw==
`protect END_PROTECTED
