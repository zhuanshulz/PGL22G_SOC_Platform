`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqlhaGq041FV5icQNJbFl1hTtb5oYqrLjc47sLjANLqHjiAB+ND/VtnHDNYldM1i
GjPPEpzpf+wj0z3B9PZLWt1QjmCCvemn2e0a1cBUiUD7JctFAZQHICFVZFo0pZgd
tRbGZ0MOe9o3TTcLe4GcSGJLAGjCrWgnyT8rp0Xtsn7QneW2oSC+YRqLoMMno7Zk
hejRB+0FNLeJk82YIqKktKtdBMBmzC8St1ek3hzUNMsLgZmQi9YlXZAaMHO0d/aH
ILelw2JWsX6S5uY0KO9NMntlmtfDwA6wg4AyH3f+avLs+zn/SnvowLthKSvvEZZd
mOt1gmDKBIAGL5jUlvvWVha5iB+Lks2Yjg2UTd0IHSJBiAiGnBZ7xfdcUGLBXhtb
sX5f1PFTWVlQN7RSSVfVYQ4zMqp8Xn4pJZrvYBvNq6qvAbPpJrjc3g9pqHhk2iwn
JU47QYgCcxoYl5L5F2wPQyAU8e/bq0Xy26Qb7nWzQd8p2X2+xBiu8MUNYdC6k3HT
nk2E/5WJkfbRuNFMy0ODLYOEjjy5N7t2TEx7tJU1lUwOh2tCYusGS9B+hBOxEjLD
9KhT2KvpZZnxniGR3CaCNJzgLgUMmGEWryFadFYn77TVDyWfBiuEZhT+fMtM5skt
f7s4CRG1xiO6LFY90ZoRtcRMI4xKdAZeVXF/8cC9ahxFy6dWDjQr8XdqsgansN+z
6hG5uyBXYxLMB61PDoXiY7Bc4wBUtekAvmekGaJNCyrfPdy2iiKDtjw9Dwy1526a
ZYpNOm2Z1JhtHb9hP6mM/oBEP+hK31mu9L9bKq+8cV+POk7Zrii/549Qnn59AV6n
rZXDXx6mif8z6xBy3kUiZQz+PMr4nE++Em6IUJNGtITmLI+LlqG14z9vfLFa/uK9
aMkIXyWmdpbWb6xdS1cyXu8EWFB/wFqrUjOG4+EOlF0eN+X5MPyH5DNQ/ZeEMvRM
rK4DLbVY4NJuHJu/kY3V2y2sGkgHNM/TpILLZ//gVYQ9IEJhIh0kgksnTdJPMaYC
rqk18tZ2OiB+toZevj2LSo29uah63VeP0cuUzmmoGMXl0XI+g1dyGX5rhaJ9y9/6
NL5JMmtj6qPQ9wyyEA2HlYJFAK4LrL7CNga7H16WJeCaEpSG6sIl7ZG/gwCjKO4A
6S8cYzGTXCWeLVt9b3DY9Os0oGoiRwwh3jn5baXIgt0gcnJIAg/KES41SSi5D8HA
aMv1/wv34qJEKCl1rX7kmMqf8cHMu1A6wlrwZQ+qWTtof+e2Pv5woJLOw1uTTyGG
pgBq5MwX9OljngBmFf9QUMq1HUmeygo0Vl7a9I11F2gZiEIwK7QJl/j7/o6FH0Gf
lk/JiKbbpy+k8MwIdeUbiCIKqMOJ+lGHkNGyar4eNHiW3oh0whB8njfV9qspWOSj
1Z68O0HTMMJD6LXg4g+se1xq3oaXxufsHvR1ldUNKcf5D+V8h9SFclQTEMnncado
8/FPaYZ6zbkQjkHQcZoXmpqccnMi060EZiS3B7/CuPx7AaKkZRvXO/4c1/hFnr2K
xdIBbZwzdfVDfb7E52TvtATJRh31D6lj1WCflbGFIS4myIrLwXCtfSFCkOjlsmtI
cVUYNRIbtdtF+xK23hO9ZUWzx7FMrrudJUo7v/5XunQb21+Q7e+xtHclgSsNDLPS
OilvF9Wn1pRSaZHLWaK5FIRfOPI2/P/av2Hciwr4V8D8OCjGMP4d/5ZyXA6oIJV8
SAakrmmYPUwJqkuZsg5GpIa1QkAh065fr6CGdNJ7aq3GQDXe8Ybu73HByzVu2EQg
uRj0R8GXXiW6FHlBRxbFq+N89lJ2HY1tUYO19S+YtFRL0AEPjWNKZQtdKz3/0K36
n2cJqY+AM29p98zNS83k+l0YjuvLQ5CCMihGfnnbW5BjHfQFMRFzQrBk/rHf8CdG
r1roXpx/5tFKEheo1Ok2iBBruhHEZ7Jd3GZL9J6QVhUItd4TTYKAcxqTYkPe3JVb
NqnCqoGa7BIeEHcTXxGO4PaBO7SPYgDGJzwuD0c1oFkHXLskwLGrW04JZ+7avdJQ
q9OW/RIdJGOEg1I4/nIEMwU4hfIuFpxsY4GbxSXO2/h84vR4h8/GjdvGf1NVhCzI
yQzz4l/cf6j+NDGKX6rQH/I7UOtWe4hgaibmvdh+hQ0I8BTEyd0iZA2+LVaicscq
X6rt/nqPpBuUlveHXcGV9AlPClGCB3xOc23GTv75cqkRd55NRamk060wnjrx/sDf
lWPb4lOfAvBAZiuPYowXwu0ZtBT7UtzSEmgHELyCtnIVj9cLbQ4EwuH4e23+04vl
XczLlbYnpxqxKv9g7BpOC/BJmC7/Hfc9kTXDkPDObvxmOGJ2Pad+uyl0yMHXyB75
gbMXSVwHxFjEHyWTO9ACytRRb/ZxAlTnYlhuxdrWsIvq1Z89vgNg6IbrA8+1e+Ln
hJX6iz5yuC3iZuJADbf91uQyPlsDKxM1fjNDxjviQu4DOvmANWIA32BGgjqySs/o
OtdjcfxlJ8eNyQaA2LUHAF/rylwIvrzak23dKy3kaekTwgAbyw55Hj6naPtfifdF
F15MDgJZD7LIk4bQD0n52YK0ftCJJ4FPs22qQ03QkmKEXHAfNwWn3V9dW9esGRih
kxTcFaa6avr0Rhs7+xkOWJElw4S1AInK42iQuAI03dFbtuCEDgD1yjDzzN3/Czwu
VwUTiYFNkYqia5zc6q95gVYlCCAQRQ+46e5wX/cC0D9RU+p6yWWx4eTGuWlOSxLW
+4aJX6JOmJ5P/UM7ZBw0vg==
`protect END_PROTECTED
