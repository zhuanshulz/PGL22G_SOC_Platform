`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+PZtGB63Ym9/oKrRmq3q/ulx1DXDw/yFKawcmhqKJaap6GSUfI8n8aktwwZ+HRul
pb067vIELlpwGZ1GuypfR0GjzrQNaqBRSk7yNJG5+aQZq3dZlDSxCFzh6A1p5cpk
zBqyBm2va3RxzHcOYmpK1fgUzGRvUDMQxY5TyWAiljcYGhmbPQqBwRTPdQ2OgzJC
EMhCr/0UvnTK9YbsfcjZcHpPQW3E+hKqIRn10WpNceIwXB6DXTq4t7vGCZlKpy6G
7N1PD9xo5hag0cId8wKdsZHzAb1/NCdtd5Kqd/AHa3VonsQmAjC39COXy1elkWKJ
dtoLG1I3/FrXF4PBN08rp0gUhhNkQECLyBSq6lfsvpOB86AqMMp8FNdjLGgRZ1if
FjYe9ac1SJwOauQwDcBQ5l4OJEwY+TxrHF30AtMI2EtdNLsMzA797RFy+Qd1o1q7
KP8PKKJrWZbrsxZxGMy/GDYUpQTEnRw78R/knwaMGYRBJzdeWyzx5wyy4pXjAhle
B7xMaieOEybTSWN5vgFuax9F2Zw9fb7iFcgnFDP9he5gOg6l+WMQbxCAocaR65iC
YGyeVHHcKJADnX1mrMflWXKhuiSFDS2OallQinL70HsMGlhuFljKNe/y4GZ2iUr+
rHQWK6C3TeeZ3uGYH4Vm7UE9NooikEKcNV5NJ+cZtJXSfpihI6eTUbioi8nerDnO
qqYJ2X4PdEJrtkNBCafV/8P1aDUXNFm7C1wzGdujaPrQqHkF+ZoH8yXDXmoH9m4h
HyjAyeSdMtRZ6KD7KUXvIYaXV+VtT1PLWhRRChWp5vN7Z3dvMHWJ6PVt1lZbEOVd
dTVl1r/cB7A14cX/2+DIF7OO6DHc9Z2a6+BXS0eKI7vfqLTrEnqeRN7d3zNaoj6t
px4rFTOCRGRqC7K1ZM6j6SNFCE+aOnNfrih3Cc2V9PQ0KOlu+bJTzgCZv2d9D0aH
HPyd/rlTLrW2lDDCs/ndFSRoQfl1qiCDI0UrI10bca5jjNY66UCezVE8/osHyYU7
QON+azX6K9ZB1/FQQ8+cBZPbhNfSDkZjJJJ0+qyULy5/tQaXCCRSN+bpfvMVKb9o
ASRhvGwUliO4wlnhQ1Y0Qaj6LJsl6max+Id78OY8SmU5Hp0/3uKB7bw8zFHEZAYm
4Vrp3An/CmetuvDx9tpqq5rzU9YJz2phdwB0LbHU8hjR8ZQwbM3pwHABOONmga2r
uz7AR2vKFXxxB94aButlZ1+WGRZr1i+xgCzYLjlqcMtfOPNAdF2/C7r21ETdzHxg
/6QbdfQZdyqTPz57Uv3CoRRoFG30c3A6ceCPQGMivl4BkCIDwnm1w22ItA3YMUPw
ErXW8H9Nl3uh9wlGfkrzjaw6aq6ypO0Q3FmlTGaNc2v7J+5pZVdVpYq7Q8sITDPV
uqX7BAtw2GG3/LKEjuiczUgQ5GxurgBsE4jtbtfsA0zdKJNZshk2xdGDmGaOEiSh
o0OK8GFekUgARsgYCE97ZBn2vRh8JpbmR7JkF7c67l5mRQWSLv8/NuJBVx8nnqoC
S9OyH62broc2/Wsrmc4ApTIZTedw05iOTkdWeZF+EF8QwNaLVZRzOZpiN+Of63yY
E/MsJljBOwjhKvCxEy0ZpY+lzfmzn0EPv0vFU8B+vkS87fmE5C/Uxk5G/ODGtRmc
zn+D5tzrWRi9Oz9kZ3r5gTt0mHJR63n0LDfQ6T+F7uVqWboeSQuucHieJWTkdr3H
z2/u2+oVuAu1hRLW/lNhc5EkRIjFXPC6jN2dSg6UfYOiWj210GzDYeS1unXhv2SK
op+4AKQCXzQUttD2Np/rEqUJkJ7VA19SOC05cu9bs1rbPgoq5k86D5r+bZEx0xoy
sSpoSoIiP1K5Z3Kgh7J/13tbFeNCaOOaw39/wjBtarah6ctaIjocA8J6/kJVxR5a
9s10tQBMSaWLHvNwGgldDZ6SfvhN9pIMxekb94V5FwjDM6eHD3dh4v2evFSnlnJ3
x61AmtE+t8/grgalmAp7jAIadIzceAUnmizPjxVQlOwrCTlZrOv67gqlFBYKop3L
Lnob7DqWZWtZaXw/+qKBCHivlzPgTLbsG2itiEfgKQt8GAMwG5bEoWA1tapFQ6Tn
cki0REqcjiWG3ufR9oLBYQ3BE3aa6MFMIXMeyJ/XbgRC8tTLDYA6ElLteDSE+3QW
b/bWW/0Hj47bfgADFV7SwkWmiGeDl211D9iFv3+nkHEiAVCToxsSk4kSmc9MCSa8
wpoMbhSDSbss7OOVUKNQyRAfWVE1O6b+rAHkt3iIHT7iXrWDO4bT8Hg30z2Ol8bu
gWdzjEAMjKkRbsV2awcCf+RU1bdvKvXD2xA41CyU2VG+UTjF25H9bAUmSmIjomau
K9lNnd2cJx8vINi1e/sK6+Fp4MrDaadKp6enTTJ+Ds5jn5VylYXa+i+yAz5AflTX
k7Vr0KI0gS987gdwloXOOGipwQqoh5Kg3LPrABxjkFsi4LPjXBmBooWvUvMGuN59
Ob3tU1cz61mX67Od+YCCifozB0Y3QiYZgP/Ilg5WkSt1wJVcRe6ZEYtJXLHptpFF
SBL2KAEyl9cp3kihM9eofA8bivWRsQcRsvP06P4vp5Se2sfSJDdJdpN0ML+W7Qf/
76EYX9fpz4AQpeiUeCGZ762IKO9Gor9RiIAuNRka+oIdUVwYTnsQ2xbtk22JHZxd
vwSSPHkz0ezYcE27mKHyuDLwQTW/0TvJtJT+MCKeRtwYHBpZstLHUAOO4aQcdnEL
aiYaZDqJ9zYHiw2lwlFYICYAfsAZdanJYPv/LOpVbEpjPQuY40HHI8LBhDdMF62b
iCeg7hEOhMX0zgN4vVaBMH+gj3uXv30F1by5WcuLwJ8Y/4o9o9MxQEmA6EmxCJWt
LtoaholA/qn2zmy+VKssBOzmfetclfTuo0r2BGw1cfv//qfNJrtJqOEI59VrLXFs
EjvW+hfZkBAlFQAWFcHq71Z7oicMFC6DQnNXB7fjE6BG6sY//kS5wZ+1H3YLoYto
adYN8hEN1MBcq6+tXpRkjgKhW/2hbqA1pV7Dp2+u5QaANL3KGlMEFAukrZIrcEPq
Kt2OfGXM9ky08wcxYT0G9kTV4jz6AynCAlrVd98s32OMVvzA+wiWlVObLONInlY0
yf2vw/kF8hhVsyXDj2EcHAYF30numhH7r866Za9mGP7/TliL0JgT3u/751DQzme1
zN/qp7KCJMBOhfILv0n5UxDMChxVcDfdn4yydKF0+t/5lL6ngm2MCX8BlutZ0ydt
PFahzzJbIpsOryfjpReSne9VXpiqYJyE5DKw6Ue5ktgfOi3X0mfkHjbKUxIbOTal
zAmsufdp/PMHJmaJQcZ1lGDcy4BQNzYoeLyiaMPKQeUbVXbVwyB/oCw7RB/ORo0r
yfexFzY+1ylAS77piCC+TKc/4ZtLJMpEf0hNwqthUN7DLGXzGbT6hlJxT46ARtIc
pvcymzJi1I1wPGnvOGlsyNzjUSlwUCoAtw8cdUwxDkOoyBK1wGFg4YcxB/H1pvSo
kB7NJgbulvE0QJZqCD/6IKLlrdeS7X2qQufpe/ygqkFRlO8A21Ax9bDNnG8/g6aJ
8gfhCBDCbCR/ih4pm0wfQXUCEu3JTG8SUR5jtjHgCHAeVLgytahLdWHdTs6cOF1S
bW0Vu436gZLibitpN6sKGQjMgMJ/kI9TYhagMNipqos9/2tFobfLCYVU6Vax0lte
9FYRP5fjCdyUMKtN5mTb4JGAjUow6iQG7bN2n0QNQE1svjy4TCRUlJhySfZu/4P+
5n0NFnDvxZtO33Blnr3QXnjlXghl/8fC5bubnlrS7TFumE55hSzLqeli0sxFnjvJ
DyTYYQejJr1+U/dK9ZD7RXelOg8EYpOa3bAkpPFZzyxpsP4YqhYwZDF+0StGNbee
SMYrq1ZGIKgmQG9BjjVJjJFPCF9xyPh08luPDPhXpYmC6alFswVFMj+3OCb4cy+v
dK1WzwrfP6o47P5cJZBPtxixrn4WBOpKkDK5ldT0IMGmUU1cZFkE1I/VRk3GOLzK
P35fYtYstUrEAbPrL47WItPGtPslDHabvD7MGF4mYyLIQNwh3Q1Og3qmzAM3huSB
Wjk6MxOXRMYcrtvKHOR7Z3R7XYBUdEnIrjG1QOPTy14w/p4ySZPDyCbMi/vxCogj
LnXxg1DUoIb9Df+ONGujHawMToAg7zreEEYrMKQVYW+RRsNQDxrUEi0RpB9G0et6
tna0j0Cs48fZYZsBw0FyQZfgLGcDiX3oGpz7N3/g31nZ+IX6UxZOaGgRARpsYccp
sHIPjOEVtLsQc4bWDfFiAEiQQtK0eKkGgldqkJthk76l0FR2R1whNSlRp7RXTntz
S3GbUMyDd9+/saNM0fE1aLvR+OMsKHfvBzE/CMxkzmmMiahzNADjpCMZX8iiT4sY
KMp7lVYhyzSrX/oHJBlpqhM8DIWC5OcTX1UlDR9g+ePd90FQ13qAY7H+AHqygGqp
dFHzkpSKH+ZuqFAh93oKhZX4gxIgcTt9t9Q6qDFU8TVaO8Gmh/HqaCeLDpKsCaUi
jBHFN94qqiHDU3uNktT+lfk2ABDbdRNp/mRVfEZie6fALY013Nd9Rszeui3dr4fY
GuLS7Apa/C1x4jdUcSs3W0jZmElXvEYF88d2t15Ys8MbgJO9C8oJJ6W6loJKl7BU
j9w/RH7bjA/s4vKAVZsOTHTl8qF0B11ci9kA0bRpyiG1sN1DpqHxbacls5STSZ0n
Ue4d1ng/TMl1nb4P9G3I51qm5xm1VX0Cgw5Kh6a1nlTLhdEe/ydJXw7h8B0r7qbO
j8RRX2Az3KxKqH2EETIl9l5g2pyMo5nU8e+usvKXpbuKeRSw/3iIMvWCGeeZFfG6
lRQtKzWhcJ1isdbm1Y5FVxiVFd7jc/Px2FAMHktrvOfPc56sZHcN8gIG+R8mWpkV
kx3/93KkNwxlUq43+SKiZwefV6Jtan4oSFvKPJL5vdceJ2Pj0abWbjBOXOOCJaP0
2nb9SSJtQoZcJQ/vb3N21o5/mI/JMaQ0W8f5ORFr4CHVWYWgiJescM+S1ffauT4R
lRhfcHEIsKUzyYY8Sb/U/+NJbTFf6hk39T/s199TMay4EwyURmILy0C28oQsa0Z1
DcyfXeY43cDG6ZkKNWwxaCC6ILZd4x5R63QvRPyo0e6N8xYd832Dj8xuXmV8l94+
9J+iyxoQuQg9ldtgcjm5zlCgUj02BntPr4M2wxbX3snswQeKjCbb4Jzq4NuGSyKW
BGl3PIFr0Nj0nbJJzhn7MgSwy89g9jjXAzJ1k4yixhDum9reLMtIGKNTOGF6e8Sf
T+ngZKj2jqpDKjagAOnTH3lmEPXUChLV99eL/jUAUUhEIPuR/K3wRqR1Has0mn7O
ekqX312873lYJ9OVYQjFCrXP+G/ehkHBXjoLXwR+6DyhD4EyDsSDynBnM5mbhOG7
Fpu1sBh9463jeP0udTnKg91IO4AK+oQFE8ynir351qV/cqMfy+yIEpZ/itoQnMKu
BRIbMCK953GQd/0Tj7RjubQynKLndwU7Bib9gXiA2LV1sN1TPuH5u8LiY4oNGUs3
eEd68NGIPHnvHMZlxC/hF3Kh+zvCYbukRL7tauoGfv1zT0UKt+E6hVtOm35n36yD
sZtwy2R1Gdv+bmmklu50/HgD3+6niDIN3SYZHqJIkEzD0zCYYCpWyYcqmnNvkDRC
MWzhdOVxCmopIsv2dQFX46SOdgNNsTlDmLRu37IixC5yqLuNSowzoNZIegyIkDUb
NW4mS2CO22/NO+VbmMEvJIt7MiGL/y8OAnzmvQF6b5V0lc2IGdrn7CVyr0A9smR3
iwSbuLa2iRgSbEweSijmNiwxudya5rT9v0l78tNjYtfFKa/7XXeZOhhQM2zCPIht
cTfqhoFPoVwenVtlMdEo2ZOmEMF5/SEHN2uNzTEO0Mxxzdo11v4pdqY00sKQ0gQK
/V5CrsNzTx8flq174NamW8cIcL/jyHHbdlrPwjpRf+ZLgeAeqlXuMGQU7cBQlP9c
voYTfnMQ4M4jJpR7E88u929LMisxlV5dc/o7W6NVPNLfBBllGBxoluRfvaOCxErc
E6pOp1CkP+PunLpMxGVrwL3DG1bhdb5D+5z7ogf5M0cIFnUx8LX6rzW+Gx2tybgh
YatKAizH08JpHWRGTv7iuZqEn/WcsVPtu2V39zzcYCOBuywegdz2hMYIWr8BIAVa
PhkTQ1dxKf+vF38tlCuKiyBybiAtZfT3sXYEOWQKcMIOGyL2LmBDBXNPj58tqjd2
mf17AmkEUEwZjgOb9fZwj10J3LPeiyj3QemXGcXFEFBIq+DBZW2/QRyelRpQCdFl
XCyoCsce7DYE14VPqcpVTp2BkOnmt0MqK5uBSz/APkkzAguIW6HJUTAk3puMGqI7
HArAtZy6BQvLtbYsX2P8pGy9Is8R2kTmdZLHvwZXXfkf5zvnIVMNhk62qCceq0R8
FWWuDHcoljiDzin118n0EllKp5jBflVZ3l/1BJ99Mbs9I0xWf16+dK/LctqWozMC
TW8lwua8CjS2qKuLIZ3dh1dRMl92lbilUi/LGTta071ZJRXXrnyv7Ob6+lI5Tkra
RcKyyzosOsPfdyi/WHbQmwPln228GHOpoxTyHg8oF5+RKc3eFDGJ3rv3yEy1AVs+
mNG9IeTq5U9dazL+8wDv/bMt+3W4PEpmDMy17Rzg/7fJ4l/SPjTViIM4/XrwKWjN
K1+7/bJE3xdOXtyVt8YLBlMzXcEDK4Jc99eNaspuwfUm5LBWPWboofhJYVY/dIT1
fBE9eY4gmNOJcUjoyx0xAREfI4gdCl7BC5WqEB+57BTVKoD6w14+wsTbaBpBKqpA
36jM2qaYNc3sJw/+2kF9VQ/AwsPNLV0tWwcKqXJyvrIC70OfuBnvo4Rkp7dDt0Sd
xRizT9Dru9i3IZHXViF8QB+ia+P+6QpwHSDQmKQ3pEXmf6CB0m0SRyGDdy1nAGUB
wEREWtfiO8xPcgkNOtZXjkNWAIXm4c8UEgarzwNLR1k+YXJkZ6nXpiqhaE2ZFGIB
Xl4fwQmNSSywlOmke0uHXLprPkXaf0N7CckFgXcruPD/sfAUPZxUICGspKqXyKUm
rrM0Z1rDEP9RIbvU0HaZ4JjykA3GQHNEGB2cPX15kmCta8tiuOWDdUagBbKcWE7t
GpSJpkKhPYpse7qAXX0XGcUn2J0DZrsN+9DOlHs0QMT8Tmx72p7dAvIWdjdm8xa8
sAnfnwrXfWWjrahZ6F1+oa6wOKjyHLgAnwyplbMkdzu8QqFfPVZrEold99H6ibg9
51ih3rEbSIlyiBeZu/mjqGrtaPcWE/+P5j1i5MYdrl27LX6sBpTu/ReSzOjBa0ap
6i0vvqtPHNrdl3Q6Q9gIM7lNkTFxrMrlYD+5WZvpqNqkt5PaPVp3Dwfw630xJUS0
SKN4FewotIxKr8NNUd5i/C7yNbEwEA7qIMRdOiockCWVm4BTZaAeQFIWEMvHMrNX
Lq7Tk7ZP8S3SOobgD96HUAUpmyLj+ZDoYI1HWpWPpj16nfPtHOp+OibvK9EFUJ9n
HwBd2IODHh9tLolY4mb8cTGp4EsMSuk8kQ1Yg3Uid5bIJ0iwALycgBHxHzLQD3D9
VtHmyyLuBTUGgbesr6zxYsN+oIuS5ZrexAkpodl+WLV/qwmHl4wVcwMjUAwYELCR
SRabr5FpgTDaGGWnKuePHeF1t79w6rrRz0IbB8J4Y+TaYxkA/LQ4vu/5gm/Ogl18
QuRMApHmStQFUDXPHnb/ImJLSwifHol0EFFoEpSSzfafPecjCnZg2ZUC+R5bCO4p
LJcklr8rWuvsE74nIFfjcJM4drceVO9cbP0cTfFrhz7Ijjj+2+MRwlHfwUd74Rmu
cHwVI9cAsCqbOO9Kd+mTyU9KZz/WeRTWq7fuuc3PdZgiGTfou9Q8JsyRTKIHo5K7
VO8IKWDrAtotPaFLcPbai6dEi2aFI7vSa9DOvnVlqRxbG5bLHcSA+7NnhPz3dVT1
YZzcPqQ/8kd0bMwLavJD8twfhYPN6+jDdDjG3of8W/IE1joSBIXYkNb8XVtg/1+z
iWyHl9Ct+arvAeSy82HlUmALrvnZmT8ThH4b13+h/0/0NR2l3fRyOniOq6evRVeu
AEPehO3TJjHSZGqSvAN35V34MsSzr6c3wR2sG7GW4k7deeNvT/kEMLrOjUWhjr5W
lJWzmtZluSwe9kb6tnV+R/8dl6vQSIx6Q9/bDlOLbgPV/FrkGwFgk9LOkBbH6tLZ
EBf9hRrbmtIdxPngIGRJTn0gz10LnZHgX0yGpQtLeLYZhiEYPVkv0XXsbtAPr/ua
2i4X29X5bhdH5LOQN0W52N/YvpJwrb/4IgTEVHdVNVaZ1dIIPIzP1G7ECaytZJX+
h99t+vHgtl83HGMsb9QdUPY+EEttqh7wYvVsDjC/I8ym5jL5L6Iihq1gyGwECPwR
581iZyKmejVtN79uKyEP8lNaoqHjIet5bp5AoueOoxJaZ+mbJ14Jt01lRmdquE7p
V5t6BkG3CrmPqJqYgboko4nhc8nIpz3gDemEwpINbI9P5wZH+9jGJemtNKe5yK5D
W6Ur0dSatk0x0laZxZp6OnOH+nfSoCTgELj9DseR05m3aOiLnj0IJVzthn5iULNw
b8N/anIgtUmVJLrwFQZ2cQ3CUULTudQKpOz3BEcCTDNVazrysPzxjSEpp2+sHVln
Phgainuo5MIAK7FY80blRMM2mz/HStLxpxR2p2+TD4B3VuMM/jwu9VwWMrP36g3C
W27XXi06/quoQCsLEh9S3kG+bBmTQrygzI0wpl7NOo8a0GokX0uPL3+UYH/mUrs+
kmdSdheJ3+hPgofnaTs/gNiX26CNZPVSj1X8lqsJsP4/f2XtyUiMUuVSRFufq8xP
XIcuWmMKRuU8rJC+qvu0iXe/902AQf26BEvLsM9aXaso2cFu1C/F6DaJEn8Wncxc
dqK3pzoJz4w8jDBZkvpgO3OWbrk6c3KcPqWeb7/KdrjvNRU1TNUxlYzcVUGhV2/v
cnZTzGAkKizVPyRPD5Yna6L2SLsIqRZ+rGgQdIpuCHbQuuUYqr0kJJ9G/QzWLuww
bUd3Co7wWlLQXAAq/K/NCk1NL/loblfzn47Pnf1tEKusFbnKBjvea76g+XHmgKFQ
G1RFaCFF1UMINMGm4KR+DNPIWeap4EDwZ246jbwfQn/BH4PiemXO7XcjZZNR6Hca
FmockpdNCOMhw6hZHzIR6hH6/pA/RzrsD64eORNuoan/eYBYfktvRyF2fTik5j42
GFj7q6tRa2qjuSf/gIhDP8mnCeMorD5LBKZiSbATOC0Dm9SmAdJlaGRHhC9FtwOR
Ph1ngVgahy6CZdsFAbtNwX2JDrT67Eybz4WlpRRgFfILPho0O7UAYq1zvPeS9+gR
c2MPQ2ThzmVy1C/4y9fYmTu9BU6x/9L1/YcdReD70U0n/bmLaEVqVTKQLeNQsq+H
wk9y0W36+petiY1ojmV16mMLD8pzo0XnjAbOc3f4gGQC+y8eXTECmq0YgW/TD22w
O3VZ+JYrt+nSRyp9lyXCO3nGw8b7GnOftP+nhBKY+0p/VNfumtTb8NjMv1OZbIoh
Tt/hFDNF9920oXB0muoH28Vd+ChYZlkmIHUCzGnG3hWoz/Tt4A9jAGlI57Se7tab
u24kfYkdhABItqIK0wvsSHOP4y1SK1xDm/FMeVBljcccuUEo98BZ1Mwsp65ZlR2e
40YU0dquAqHMxwf8xa8zv5n0RYivvsgaQA5BwzoeyMvokUgdvC+0QWmziaNAjpsZ
TxIy+IB2BfpCCtLtcDDnjsrR+3Wq45I9C4VfjOWiCIJUTc1bth3yJmT2Rrgj6tW2
0ZGp8KFYegw7rH28Bbwdzd33jUeg/cG2hwuqIYVDJF5ie14Msh9qfhdxVFjtzKXY
4LH65PeOA6EtP+pAIMOpliRnQ1VrNVFXIcFJGNk2ao4VnRs64LEqoByKtXjfopRT
3jT19TU1NvcGyHYs5tF79yBv/AVw98rCIhFd7JadqM7LUQUdaEB8W4o8xsCGZ2iA
ihdbQmjKz4kjyYQhVS76eB9bwEkFhxpjNOlvR9fKzKlB6u0plKvTfcADHwoEJpQN
KIGohTdJoR8Kh9fbWzufTB3AsxfIUZIws760f/SBquD392FDbrp37s2RdsLxawlj
BbEezKS5wBaAuIEwY304Z/n60+yxOB3HnHrzlHh81Tk6DM3luPFmvJzBeeQcvkVQ
Gv9mqsF84vtcit2fxP4vppAW0O6tQcFmuyR8+nOD1hYYkT1Wiw1m1eovpWpX4oUW
3n3Fj1pQipjhaI8e/J9xsBNYl/ed0mYls9BSyb5iwwyd9+1WdV5rKHo8sFKUT2U8
O4L1N5XPEZaXzczpQ4Gj0H160GiPjh+AtOHkbDecGJT0HN3/13vIl2IoXvvG2ocS
p/hw9FKSYpVR9SCMMUhFwR7HCUJaRgHiFYTK5AODUToLgH3tsG2Q6EjgQaM2vITm
lAhFV91DEnupBcg4nrnSDCIW3mlH8hlAz9tJ760rCyf37nBLjYkn93T9KzqKxM7J
ohx1VEmkV7nGJbrY+96fkZbiGRqhtB03m3WQDwn4xUlXCXgs25RW3t5gIUuiZIdD
uZ24W/gUnaQZ4+480rvoGbW4ieYlcFjDvd9GbJZ9zt7sv7I1bHKhRhCPEA2vor0d
29Fc4pRHwB9Hbr/YOjZq/Rg3Com6H1XnJWm+5NxvwrlQ5sVEGtcBiuT30g7yRsyW
UlFdnXq/L3LpNh7bYcL/RxBkxKFnPO8e96mP0283zgwfAzLCVpXyYOWFXGlPaT+m
zztM7Ovbu5oXVhtjJSnUSH1EYaMjd84t9R2hAx1Fwz0Z0MciUOmuksUgEVH7s8xP
DzAvGengGhJNFtkL+JklbCaun3QgL1q5f7BxzmsqKRvMCFvXG7ATXqlb7DGZVnys
z/Yx6rP+IsKaVgmkxR5WuegaUyRDR862iMlcps9aydeRKKBeoOvfzs06aaKgHgaR
rufYz2wmi06d2jJJqABkJSkQzNCdhXJYkvC/yvFrOQofcRSzi/19YosYHoqZHmhg
/XvgANpfLDMF+7rgXEU5PUhA7uFl0vDHdnvgX0h/WhyChA0S/1tE6SheLkyh0rex
Abu0SI6Bdob/GRCQdjj9UkU4VSIg9mVhAMHqAt+s1yzwPCd/wlr4tbPb4fhaqh5e
NLDyrD9SZB5BlJ+NBnMzg0SMcRwdjcY7tbXUKk+cX90yQUamsVYHfTaBLxxGwSPX
pDA46ll2XZLsDHUymfv3HpWEQMbnXPwcAcCeOmTMhmSOoD+qHmnjDWlPA9RPirez
CESZBphRsywxJuKdE5KmTdsbnCmEAQCEExR7p25zJcdK9UavKTCyGHfuvyY8jcF9
Qn9SMdwb6rFpS0vKEzpdqP0Tuw/0up+RB+dY3AXadKq7hT5IBlXIewUtmvkbdmS1
MF++SKa1XJMIPwLfNWcC5fUA91YEeW8EQ3ehfBZCfxw7t8QAo9lQlluW2BisXt7c
hicIcPytJCF5ZSHp8QnezcMALt40syIUMUa0h3Ipmb4insnQNxrJ81rAiuQTXFvV
8EXgEKaMfRwYFh6TdXJQROmXXLXjG3rC+pUOv5/HGin+IC61MrhI0y+gV8EUyHUP
ODMWbGyvHj7kk/wWWXGPfMdUdTANCTSJbt/N/A+1E61LVXIP6Gq3MQPmcsdUoNHl
HpGWs8owAa2eiyr4oWdwqMK03/ibnWI6doX87H2J22Xsjf4u9iwoxBQD9M7Lbz/H
NoEbJKs949BDVzAa2CeXJwVLKOVr9gp34ED024rvPa79fp23iPpw8n7snzYenqEe
jR5K5ws6a70Qo7N2y6MyvHKazHk9e39A9ipYHGV81qjIld1ECWvM9wKr2C3mC+nf
M3DZRxAamgLQ55BOPKH6bfy74jTEwt7QbNQlAIv3v68WjljvqwZnv3dv5jcq4sNy
sxFTylwXaiFRP8mBe72xcFDDnnFDxChWRWfDNGW6R4Ose2LSIYea5wZLLDU8R82b
sRStcyyH1sR4041JbB8ZWFZuaZQnav88a1SHwWAJwIHPKSrETgLxowZGqS9QLEow
QBcUCtke8jAPDLPDxHSjE1i9KQ0dbm4tFtB42x55FrFL7/HxAeKIqn3PsMI61Zku
UmEpuTG2YgQb4g+Eg8MiReZmlCB1WW5ageNhL6q54l7Xy6DiMBeCcpive692EAXM
dNvDSXbsJaZijKVuvTdXiqh332PP+OFdree5V82JXDX/ksHr6hRM9BwSgrutF0KH
6Xe8n297ltugkDTb/7WiLekv7NVlzOk5wEKIoVgU1uTmwEVUvtHy5UmxKSHg7TOH
8J5Vl1qBjjzuEKESEBcmgRUW4zRf//YundvRD0pAEua3cV1WvWKAdA/x1roO6sbx
rw1+udCuoQjyAa0EU647iXDG07XHuR2KTk/kbh2VAyhOLL7RDt2l2ybqLc3+8MU2
s2mpkqHpxbBF9mGA8QM9sbQWh3valvaTS8Qo+fbPcKcL8e38+khagO95/1vSp/UT
wBf2Bz2lyzGzw+VQGThInhKSXtXDZXHMAKgIcwYes6mzioPWhr2zQCKMBdKX2d8k
RY61AwQ5xvzNpoTA8rTemb+1Y88zewHVcP3LQA/FzpGx/czTyLkeMqt3q4gf9heB
Q8iuJOeAxK5uIr1JVJoT5SwF57uxteHqruGmQ/j77YuecIcS0iUlRWUizL6foirv
//rlN2wqnJgjubRl6rEj5Up9oGws/ZUhER33SEmE/wL3qajr4PTSuYEN4WNbQH/l
v/gAGU2l+45s/1Jlkf6S0o1jC7AYXMuGZfpE1sFH+XCPrV93cm0f5SHx9XXS0lxH
r4p3HWeLY35CyOLTBh3QtDXA8/oQjaFb/SaGP3YNZTCkPyu86B8tA4Gw3DpyRndx
x0Pp9m1eTZsmkH0HH/vUfMEB/BFiHe4uhbHMnNbr6j6VMBLH6eIpAKqvhF+hCI/2
ivTyXpC+lfwybYs0HAYe2FQadl/rz6LJo0UK25NkUnLJvatylGhrEHOs+InciZuX
Ollklt/g9uakyAX5bi13mVTHx4HLRevkdWhsYg1TpnAUFpKuy1oPSgxVSlhxWrMD
QMoWHr/CTqceA+gClpGZxGbDQjX2w0/MBKcseW8dGoM0SD6KbN7x8cjtoX5ovPrt
VgYz4WfUBSYe4m6bsbGdHM507HZYhfd6J9vlGgs+LAENqyuoo9bp6v5YZl6U3ayh
0EdrPbBcjPhK7nYHg5BT1VzD44jtQW5f/ytlmtORT95J5sWqQweANEI86QBTOjO/
5F3QT+WefRF75XzcyFNiCnfl5HrMdrc4bA3lbOJrzPhPMLePjsNbwFoFO+fBmnyL
AxC1F6Uvgrsbix7St67wmO3ozCSxpOHAFoZ7LvozzpDRBB0IvydMgWcWWXp3GbQn
tVddXHn1I0Mghq8nSH4+7/raIrsMwpdox6pJEW56P6DeILFF7C0xVKc/qFJ6K4CM
VrIr11GW/I9b8b+xq+Zpl6+kv2v5uudBBA8NMeNQO+S0TeI0uMoSpQ6D3i94hYRf
I5zP04jLoRYgOdmnR4Kn1wAW/kYDcF0UfKMQGXnPwjIj2V7hgIo+xA5VrHUrtEn7
TH8pIWR5U5zmcz32Va/TwpJIgpWilvhBkEIVwp3edwPJjJw/OdkNayUfjZJ/kCI5
saBeuYZjnJQiKxAyHT4pA4vAYnKAwTRKTt1d2MVETgNOONViW638xbGI8bvfHITK
FLDV1yVDtyu9bYiWpCzHreJPCiMrt5UYKxQg41nyWV3Q+cgcMPLbtxhFZQ2F4nw4
poJRXz8NuVw4cf3yU6ickOjwqaUvqiTDvaRdxb/aUHG2OlLpgbqMjUG8YBkRVRTG
vYp/AmkIwrr8hCz5Gd7AZGrLQ/qX1sfCLo1IYl4nG1qCXNxoOk80B0AqrjXRcliV
gv+7/y0PyZjPGm8xfGPM/hogdvOdxO2c8UmK3ZKUAp/rO2OWX7uJ2uVi1OjDAZwd
eoZFwPmD51yZrb00PcOs36ZAyVidk2kspFfhumfASVfO9B9JACpMaJC95hbJQlpV
qV3ImmM7jxyNHTZTLWdpASojXQOBuAUok64O5s751DAdtTLtUTIIZWCWEGPriI0Y
4w4zfSrXEiINKCaqQSjVRlSvgHdPhTxKAeJ48cUvXhVWiXM6NH+QvJeDQtRFOPwo
WzEftctytRZPCISixEoU4bReemT/h2WzsGQ6rS4mnsf0yrnCrYVRHuMMqu9skFZ5
caa6rEGv+NHcahcso1hYNCjzdWRI+n386Xtm28TUxpycNhqRYmYPbCZDH3z901Ve
5ikP8R9ko2NkPoaTc7WAtYmyVqi3SL/vnkIQrz8e5p03cLygfqEs5QdX/yoxyscc
fpgHxA7LVd7TDqSAm4+mMwnx9LDjZGnCYMQFCRszW7rK662a551fBMxr/Ankgwyy
CXdAIQbkK1k8fwrs0HlUFAFEaRh2UyDeWwQVxDgnxsWDnhThi7KIg95WnRz2MX5Q
/SshlvTBEOtFFoMXQiEHAM1iq0/IBGBVZsh9NBi6CVLkN4aNOE2pAkHXH7b2Us+t
7vWZKtvLOgglDZQ/XvI1H9L8SUoV7fBxQPuuwnDr73Yav4PuNkxBb/xLWRwSYEYi
IUONwmZ4Wk3FPInYUJtNNYtn032vC3ZlicONrpNVi3q9ec6wpVpH2Ow11AgcrQXy
E1mEpcA/TTc7gnf1Y62rhWB8GZe3fM5jE80scBku8vgxAPyM/QSaGwwVzOEiTQXu
UB1mlwdYn2yVSsyrMgc5NywQhQ3sm6F0uZpD78KUnXMdzxXB2WLrxxhViV9ncXuo
GUnkpv3s17Iif0KEa74T98PPE/hswgiUatLql/CJwfEHjMzUWyVLI+AcpPQIL2nP
d9D6QyrykUD4I/b0zaXiFL0qc4l327VZ93ln+MmLdSoxtizHHeackdgTFODtYvLp
R7ztd27BDrji5HWEHgmRPqQwK8cl2QwKYOBQRZ7HripaTj9hDNKH6O4te3bRhcYK
IMQROvYI2GEtqWeshGysex7SlcUECkMTYFk2IdxxFZS13Sa483yJN5LFcjI6Xj3U
0el1wgjpEqhDitpsNTUNM2TeUPCzTqdTYDx603PA/UJrkuc40RVvi1HHFQ3Wgi3x
O8wc2hChKaEefOcDLp/zclmsJnd6EH7F/mQyXrD84SDk8KYgxe5upNs112ABZWPG
ali2d/3wibxKtANDii2QgWI6M/6YK0wim4T/VUowJ21YRUmWkVF/5esMo7JgBksr
c/iGRL21y0gVq7no8EOc6Qvqudm0qNPyP2+zYSmLHOh1BLHkE/xUhmwUumEraUj3
UjtXWO0Hxd6USdj3GxLuL5IIj8YhutSGXOUVh0mfP/0N0T5LQnXjXMqsXGp3DMl9
ftjsftBRQEwFQ/x1vs31FSsX8GC+EoGN6qA6v8KEkfGSvrr+q10rAg8AFktlrCYx
CmAha3lFcAZhVLMN3D1tekun6NwhoZiuLu5X8Yu/wlu0jRjX0q+Ghx4BQSqWkKEl
OXXNVEPwArd5fAq1w3kxs3moSoz/qTZYsZi1qyH2r2g/S6immn1nTYLTj/LInz/m
hCV4gZ46ELHZrh9oOowW51qNDxndJRZniI8AgF6JkuIlLhwoF/bI54KrhffHVDq4
cAbTvsC0Gn+aSj1Nw5YzsVSzLNqlHpV0k/ygM3rWxJW9FeKIhFOCNlnc6ryV8y2Y
Wi11e5Oj6q5qSMT0mvQA8MlXRtiVYGGZUN47+mSI3y75plT4tY7IG3kwdCqqSqhx
AKjw0ih/UkAwC1MNAC4o8Kt3Y0TAjVVHX3MYkCSALr4T4dKTadw6sV0tRGQb5pzp
FHd5YeIk/2KlOJHC7JyjiqrT6VlOgjWdAPN334KAD1SScsMHwXbRlinYZQZBkxXm
DJy/nn4yS5/yV8iQsC2dvfcQ/dnQVmezYBDodOnCv0KJUCKHhIoDLMaZ5AYvDO4a
Hu+ZNdhmJUAb3TW9wYr37eQ6y2Y7HXgu6flhjh2LO5qlpvealXkEWW/1QHzYfl6J
ER6U+uNprSqyjVF9It/zeLnWQlGdC30wS9sCI8oPanm/gcRIGfQX6RvhktUOkwOF
Ib/oCp3MNwclRK23GdK0AgDXW22Dxf9tjavnh8zPJ/tZlMCjIwzs+/wNT54wEOon
yVmjGWyHp2OA1ZhCsVtiSMsGKYHVup4rYIL3by3pPS3ph7PGAnvI/L5cZJRxrnaX
LBMD3yZLF3CzeZnuw6/56CyVX9K1+XwyTeaSVfzKbH8vB4KULpt+H5dNMolt12Vh
rxssB4UteTxZTRT98PQYKMqxPaTnSewFJXLmZ0Aw4FeI15oSoHuQz3SEhXRC813O
F0p/gPP67I/rHLCnVYGBOr30BFrAzaGc2QdPL9972V4wD/eUzDcTcuAaDzORNEvm
s1/rCGKazYTGK1f0N8VKcvnRwTCU8a/a6sazZyqPywVWxtDmo4RmrSNBCK9YmrVg
ZhKAwieJ80aEAViT5eztCRbTi417X2pKY0ruDYSrz1zJN1mvlzdeIa9Qis+kE80J
Wjs+RJYe27INZ5otvawyp/aT6WZxlLQJTP4BijOkRrwd4nfdeL6q/rKAlphm+gZ+
1P7tcghVsftcy1VNNMoIWW5J2lz6omAz4d1YzGQYqpawS1DGdLcFQpe6CShRM0x0
ht6cl+2PMziwDOiuaBJJxNv6LIQUiDTZtkZHnGq/QDr8INPIB+Pq6wRVeLY7BhWg
BTW6nsXwd3TdCeHdhC6XVXO1RhuqTfiPfaxrxnS1yiYyTWhuCz3/xkRXm88Y5rAh
491+zK2L1mqa78HyhHpWsPf+y9LgiV3MFKZEtS3czhSH1MwXH+0BNup6R8F+Wki+
6uhENI4FQ+fk3x3nRY1ozA5KIghS5yVtG8BnIBe5bwDgoQlOE3bicPpIY4jjoh7I
FD5lIFSgd9OFI81rNagvHcmOqgmjU4xa2TA0FrFBkRj8JIl/criynmNSH6TWrxS6
jGNJhmD5N/f41NpA7HMOLsagXa4yXI2n6u3Ti2wsPiXv5PSwwLe1O5LFV7TA8T7d
Lbico8KbCPfD9rDgilxa+6jN/dhA7ieF1vYxcwlR3SL7JskscW0+cw6Zcs8FgEMH
riSWxLiDT2JyeYhMdRMJLcUzddZhrSRyZsd83bATbaLxzcmBpYa24M8G61mMxk++
X3QyfDKWSrbN1/d857LABCbC3E4gm9Kb4n5/llh2y9OqV8XnLXlvZR5P7uNfK8NI
KkewXHSk9VYYDmRQ48ISO0UWJ7xTAY6ZzPIIAVdnvQH07OAuNHz9UXvrQ0iHZf2h
1J8sXmviTQaEqeUKhXeAPzR9rCaOkxZ5pWLPDN3zUwpnNkTSuMDDIR+pILKd2Ruj
Nk/P6dBqexO/Gv+r0EpCZU+WdPBh350aEzFNYccn+Q1wcUGuq+lQ5TbkB/mblIFF
SEsHWpDboLoN5/D741OOMiz96hjRiuhtBNTbizavqGy2wfSVWaFGCC1mGZqvVVs5
eoeh2+AeBrZOcpoWK1fUvMkhGDK1UpPDSvdN9jwMfUQ3BEV8szQOv0RH4wwrQtWD
PDzHv+s1HlzkFcz+9Bh5ht+uxBvqjguDZ/oDM37EOPGhBMeVLe9DOB0VT3mRA1jy
wI+Yrwgwtdx0tKyPCvgELTsvlEgzr/xtwVLaMhZnE6AyEJWomGaS3KKXGPPhxXvp
bQREO6KatgpBRLq8Mu7ow9SeF2nQwXc6N6ro7tVsd7+MXtbi+AJh5JWR6PQu0a17
91KVOkk9mvDuTvCWeSWGVd43jXnNkwD7N4nx8IQdVQp30/tpCoZaR6hfsKBBBBc+
oW1PVOydQDkJZOrbv6URDDlCMYTISe61DDIywVVZPbEweeG7Oonw9NI490c20y6G
7mKemIEVXY96fyUhm3bEP+SvpS63etuWZw30ljIVKZqgA8xM3EyGcGnmoUGP1lmC
dzrbJeWRLNiBmOK/iLUJHHa/P3tR9Ihwgq8wql5AQKzxt8UmZc1dRGMhJ5myerRl
YmzGQPv9vt7N+YpWG3a4fBVaXKF4WgdB/opnXCc3Z0pDHink+JjSUtgDN9J+5Mjt
4vzVpXAYyrCDfZhkET2f5SfUVFoYDNmdajl73YpbdIQXE37p+X8EkfsHxTHA5Ycm
H9pa+IXB+Kr+jZKGZtbXkwniVyFU2OFAPZF/GBxVPPintjj/JEezpRJ/USiP3Jmj
5jDjasSn5KPKhveR8wbgr6MekxqfjLKa04gyWJRqguWCgtwkdBQm3qbUXWWNQ16C
/W/dTLWZUl7hcC4qoVGEWfojDIgqksvZNFEhYvaNzsFUan2W/5ttOKDxUE6wzq9Z
OsIFMtl84oXmXzGW5zsQ7R7g9LlARYXLamjH06Zzxpz0t9pBb14ZBtmpWRER48Vn
b+jdRWK+IMxnqJk3vRcNqRTMSJUfKqZ9BEpTPfllV+ZBBEkyzLIOgK/6aiHFwcVE
aQ5mvnRK8GOfzPZDj/SpZy5fQP0WyBjevcNjL1PD/D7m6+S8p+L1SqUiCj0EagfF
nnMEY5nFHabnyMK15mxBERssurZIAe9gkoKi1Z0JvaZipvTEQCQ9AfzP4VYI1E1r
yFKCRvnTZ0cCT4Dv4cMk779RrCuqMn++C9clHGkqlmvXXb1IFscqwI8IO72dFSD4
Z3QoeVHWGgPTD0aZ3EY21Z52c+zs+kuBGT/BIaM2AS3Fyt9qEOXDAN380sDiBbwv
YDZI4tPIwtjOMimDuv/Q98fx84TVvmy0zdTIb7LMWJIIou6BV0BUdaVQxwJw8T+F
skw/6UcQWBI1iWxdQO+h0oUsVGwQVjd3XWgEHJKN+O8b+wYae7ExPEPyRN4aZo6B
Jdc+OkX9GSL3Ad/yMjrLYepG2rUK0mZ+m9tQg3aepxPtbphISj8jA0J2dx9NRZ00
U+KJTdddv89B+yy5mgM7AVSXcLSdRwWBiaTazbY6FLDp3HQ5YnGY9GbqCivwm1Tq
UO7lMpHUoJKgN7HvcUuYHUmx2IPp2hRaNQjkX19oSMCPdNOP/q7c45Pk7N+xAehr
0jKy0XQxmDvXnOXmicy+K5bmPGfSPX6zWMT1gioQwZ8Om6PcYOn2iFI4nyq2iKAZ
9w/D0geH3naTiZ8tbZn3PHqbQNU7954YoMQ/c7jdzmDVFhdN48MnSwPhZ25AH5VL
gxbKjnli1NrBGqcnvpkc3LJvxbPGiqTqFbIs0q5CVXBdC/v1bcJe4d8wKRe6oJ9a
XprHiUlr67FEQuQ6UU7pe9ahltP/AVGNs6bn+rJlqMdLLMQofJm7kzZDnnpwjFxZ
9eo7oiPmIkec6DvsdEKl39CPXQrw5+ARP+8Vxan6ONSMps44BjWBbXMbjS4cW4lK
Mnq29gip1fjWw9qe7OZuoKZHaXZ+2C1p1q6qAvfCPmUzpRIOxAZLct3An4To6sw4
6RGZ2exZclU8liJXNTJAI1zfzw9Lo0IrTB8snF4HnNpG8oA9F85edSsFRZurPvZY
ZXZZobFz5V2ylvPx58E4S+kJLAR5Ktsg3A2YbwDH0KFn5ctW3FtIL0j5djLdvBPx
U5Q19gbLuP24JIgFn8eQVYbjgRApP6kWOwnd5+dgISP4Ths1+qf4UIJAmJ6fl95Y
o0VnYoH+Ou1WQlZesYVbOcunyuWKRKng6Sr/00/Kpn9iqwhLOdCJNqdElrWn3L1v
ioYp0T5/cq3Anjea35l4TD5zYRuoDokEFoZbIe6azCLniTvJItaG5lYE/dIur7RL
mh2zxQNVtmr70A1N1Pnk1BVP4BTMbbJA0mteCY/H7gvvYpNAOodoOL/7WBMlJ/5h
pYRpCiekQQ/QmyprpFkffVkT+syz3ibN+dCV+WA+CAI41nlWeEFGvXaCWHVHc0m8
108Qa3u3U96A2OHURne55PLA1HAqk91wyyM5lUa0vt5cKYJI2Jc9Asz+c0A7YPzS
CdHjgmv8D+YKfDELyS0wPdwQjM9PjQ1l7cmfn76Ncu4B6SKJp3unlxBfEVgqTUv9
kzYGtNQpm943khmuOrMK5hZEjvS/aAKfE1ZmoVb28RYi9hHQwkCh41M0IP7i/IVS
HMeChx7ATd+ZjR5JWKMhTuCASCZ4xp35fC83s6h6iEbKO0d8psT4z2iwHhtLfUVA
fAO7T9HJYCrEbPsyyOCL52A5j5Y6dRauh/7GG3ISG+kejDahmjXLpgoYXNexi+Zd
QhjxyWFf+AZE2bNGhgmjyhIfbFclyL/ytPSQ8BH8HFdMXRvzRQ7QMz+KA7WZzsl6
WxZhjoM84vUyPs0POHI8APZOWWgD7+n9DC2xvt17n3bXNAz02T47wpEktZvgkYc+
aAHktcpxFeGFPi1Y9LzTJeoxCy+1Iw/R2N5ZtrvbGrTqN5Ic69C29LCQ6ezIL7c7
CitDrpDy+BrmHHFyKuYYB6u3vYPT11hCs1S8bS7Q/hU+9VqcWxKvo/TACKWNxfuV
dBZ0KiWKf/jw9il0ZpZQIW8Uae8J1sGdTt9tLvlK8nzo7Sb/4wv7ffL0epx38GA4
2Qct+zlpR2uF0KV0fjUqHh6krS2Jgq9t1IxAQzF0ln7h9nVVRfKCqlDwgUWvZjN2
1YfvH7Bh5fWPczOQ5ftQj8cK5yC7VTdLR1AhMFS7KIGRUSOkR8vqaHyxvein0L89
2gjxiBLZA5ymcIwIuJ7XzsTIUODR+4u8dumKiyPy/iZQQ3M0XcEy4YblaRlg8grf
fexvpfdoTJ51CQst1rKmUkO+s8O5XGnpSxBpuC4YosTMiLn0ii7fydoGWAqQZ1Ob
SA82UhiinJtX4kIzFwmwgKJHPRP1o4M6BZ8ThyvkeO2G8Ri/CGsUMtym2GzRSnr+
SDKscS1VoXdIHGC85hABgaOB9p6uJuKZO5Grpicf/BcaEblHS9I5RVzKQv0mAYYS
hn/qQQhp6okTdf1V+LdB1tvAJbur93i9azoQtgxFERZY+7g/QfprAJIpV+z9UwvP
7SPaGn++CMbz4nAzFculJ0sYTMqicOO6JPSCBl5jTwajsUrJKpYRJyep0tnnvLRH
t0bWH1bNPQDaPdBDdWzTaE8raAGfE3pZo6yS+8U+KvSMXK4f68bJbcu+uAu+9Aht
PmFkPjyV9a3T6AEiS75eb01u2cp3hKmPjTByhpJEgHDL92Un4xKFtGBR0Rt16FX0
TYGWFGlMJ4o62LkqYDecY+XGYUA84dK7oEtGaGSsylYsARYjSMYoSKztsHhWPgsl
oLBs8dPIFdt7mVQoB6tsI+uct4+zURY54DD+E91VPzUyPG5mFJiRSi5HdBOVhe+k
XLeg/Pt+Uutjn/1tw+/fmhzEuuhubFOeDXl57BskaL5XCeiEUZZyAfvVSbLhTfiH
RcGx8ay/QFKMEjvTnj+ez2gcqj0ctEMYstdAQWE4XeC7MOw8CrNqyxN8mgGBbn6M
QdP4i/G/YXbhqBcEqi0xWwmznTjLtjfidMdGD2HTtu3hy439ANjSHc7LrQ1RU9Wb
hxT6LTRruDdsdwzy5P5DChfNQJyGL2e0Dk2gYewmb74J2S7Y3imLpP1vwuIlDyzs
qtA0AJAIEJXfiE7COn33MvmWuCJ/ur4MXT/NhA84n2WJIIKS9o4fIShEI4N2maNq
oKM6PqXVkQ+W+iRXs+FAVRv480J+rF8AS5eA9idlNA8dtnJB42v+tzHI/2H5QUI6
jz+pswMT/nOzghTrNBrWZgsuZSIVKiUDQ2usB1+rB8tg1BpB7ZNrkHtzaNuMxijI
PMBBiifcjc1pqrIj2bwuF01efSz6UrLQfIbQQbN/EVvoDSgDYt5QhaQG5E+kRrp7
3NQi9vVwf/OVS5l4Qi0AhPlVwCwsPdl+xnulKVnVPcuSZQJB/dOilOqTFgjUeXeM
wdDy/oD/COX8GgPPD62PIkWcoGjXCL0Adi0HsUYqgBz8QtXp1jW96c/Ihmy86hri
usjCTSfgkj404Kh1dToJkMVKJKxtvyuITs6RBQih2+kfAoptux+WSUhPl80N3/Ck
VmyQx57NzgRDHelF6OwyQeWuuZkjY30duFBwfSmsyUfLks4QRCWldiz3kbciOXsw
CtSB1f9IRsZF1l7hwaRG3DXcXtnYUcQ4C2GHJkspIG6Wwib3IrAHAekLnB8LosLl
ltfQm6cX9WSCNKQ5LtgeimglCY0r4FZnbdTUmuZKKYcZBpHEqDBjfmFC7PFgOH/R
H7ojqZ7jTlOz/rtCz+83ZYKGyvuFVYBaNqEUT4375rW0b83dYuKocakpJUU6exyA
Bp4trovLCllFCvgvmB4BRyf2TUQRTa9S0SZvClov83rMgQHkmIvG5VJ5cvhqdc6a
8HhU6lmAH+mtRgLz4DGYcWmK0IdQi2x9vCy9R7vKmM8yXjhafIJS9EfGK5CfbqCM
xKX017xgTp0iDHacTSwltJJ2vYQY479yS6ff1668KmvYBVapozeZf5egCKKKqGST
lsvCv7ucxJ3gVEjWdo70Mg==
`protect END_PROTECTED
