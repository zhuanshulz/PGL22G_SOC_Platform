`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvVp0eHnk0D6ijSpnX9CV5mICrkwrkkeDKni/+mUQPGzQl1W5n77pnawQ/pLwfqb
GZ8tP3OY8wtU+i4QP3g8+QFMkxXYGryU5TT+QfIjTfzLD59G3hfXC43DDZsjGbWV
FpyUMpdH7hDDOeCXxNYJPNTwncckYbWuVo17HOCD2QYz1YdcOYGiZwJ6VqcbJMh7
JYk7RqAZf8SOYIO/BM6fhWf+CsI68YjtqGsBnU0CFpJLp55iJnkTJctocam6DinO
t8MBY5nqBNajp0oU0pUoS3vi5L3KCWX5WL3XtCKZ/dofZ4qhBiDfuomg9oFmyUO1
erGT0UKPsGJAmhFWg/jilc7moSRQdu+j8X07zOqpNPCPn1PZSvct+kOQvo6RgSeO
UfsMDhs01g8vatxSq4lXso5ul5OK7jUfpOPT3sPICYYxUGW4Rmf+mtpQtKdSIWcv
2InuRcYl9EAZhqjKQ0RsLSgH+8ggHrusTXLSbGGPwFI+tCkea25i/0R4UlvpSGK3
yZD5P8HTSiKRnaNJ9TbPpyTE4pVO2fjusjU7As5kn9ZocV0uc742LAfnPdH5rVrr
NNpeTQimjNKyFi1IHIVR2pHJSutmmPthk2nkwIvIF4nvpxbF6MMdrAf1xH3U6wP0
X+WIsP1xBKKGGobwUQPzZNsDK57uP9ylrfNfQ7hglSBDEIdC+J9BqKfEeX8s7wQY
TyAqmu5olY5udnME0LK6hZCQu3smtDirsF2WLQ8GfNfPeYFhsQYzeDx5Tv0VMq9J
bUDe7CzJwoyQe61hM0VIMQYClHOiMzjhOivVF2css8wv5JSy4j3GdCj5JwCnAxWD
0Bskb4IIXhydnqbAUS1PeDm38Zq1hSBIHrW9g6VNbf6BEdzroK8J8l/CYNd1KHJ/
jSb2HYwwymXqsJX1w4aPSvmAyki8AUGXE8RGSdeSg7vUqVq0ovi0FP98HBmKfMEs
kif4/xD7lXfoV01VH4LqoS1SLIC92DLOUmza1X8z56yiqKVTKlmwz30P4BcH57zu
WK3Q4pfQ7GUrQrjOA5CbKzaoB2uAjSZx6B4onyD2t1VwQlVYNCF4PHzwlICuL/Z0
3/gPuubd5gYytdTMj1p2DZsKVU6GtPrcOstfoBm0d2QkS/ZcNAGKwbsaRYMTc4LI
AaLKcENsie1r3xLqGnuFg4w3y+tdXPeTyB2/EUgMKYe8HYXyOz6mFA390B/orEI4
o+viCfgm30QszcfoMhCEts/iRnkEjnUGKUJsMSPuo+3opyrXs0ferNsEo2j9ZxPW
1dapyo8dlz6rZpHEgLX/pJ9sIpplnOa8Sw7D3hDlOJ10Hpcte3AgytDX6Ro3jvHI
teiUPGnFZnz6qwgo79+v6YkiQDslvJXKjK/HHIHIrNi132/N2RraTwiHTPgtvfrc
5YabWFms/cAlGek3Mq/HDIVQ9dUuujHAWLfDeGP8MUfopwWTa+y5Z4SyLWPHBbNp
S+URrZCPny9kiv0gvyGtjDX/Zox66n6hfRDEfM/5AvwDfzrDh7WJ6C5pK+yaBTOm
Ruz/19nAxSgHJNSAoflQdL9x7kVziY3a5e1szPHaY9EEjqPG11sVUnaqCj9tyhyU
hb5d3gYnHjFzjJKqAoI0LpcVpJOca4Z8gj2y6cPZ4WkGgwm9iB/wkE5O6L9Pe93Z
IRB/paW4Mm5tGj2Ty8w5XehOBCdEv5O/rVt8vtCwcvDx+xiowxKkgnUpoAyZNduf
W8MfATRcviVp3YS3DMOpDittMpyyf7f3fA2J61zBdoCsVjje+nmYh5sm54b6oM+f
Dq6eGABiR6x+jHfp6A9FZ2BxDu2WlZdSe0Iz5QziJTxd+EcXrA3+Xhs9F10P30er
hhJfVTlQes7yvpfqGmA+ITLVizxakBoSieT5wzkQ1Yjcmh8JmcwapVw8QMFcTNx5
B2xN1/UbNLviGSMJHTtU9tk5zFeEjwg96pFjj5Dbl1D7lJHRwMGqfzoFpgnzuFzN
HOMmLdzDtGWkTkrQLfIEjOAziMrcYeYZ5LtyAl39iu2y5NgNxnZSsPWUBsEYAQ5B
k2IE3oQwGQL9OWBGUWLHVKRxoXMHj7TTGvQaYdKvzdFH28nE3xjHdpOQe7fzdguX
2p0P3UxJW+mFNW+sYLf7cvmWcnSBBQTCIC5BlfkSuo9fHHTYP5tc/l1jAEEisUNk
hXurRfEWFchENPYoST2dwplTcMDxUNp7Fr5fTclGwnQk0qiiQDin5K2p9Xqp/HMT
ZYamniK5jidHq+FK0quqWSTgP7HJ/AvzvWx3pGpU+KGzAvhjhhXcGU2js8lXs2l5
R/FrP7ED2WvhYK5zhfYx/ApUt1Eu2Haw4Wz2obslpo1a1NlUXOjGG08JCUQLUhgo
ylmkuJeoPB1ncqPzGvYfzFuTtDeDUkiUaHwzkx9rvasN4szucIZqntROTH4+scNS
NRv12N6wOKfeQOIlm02CXib68hA3PbmdY35h1fGWU0NN8KjvI1etr5/I8sJXIlJI
mkykNb0SUdT/UMJfK85uw4x86kPS9jxNSNkPxro3hJdKEETk2hPVEklcKYMt6Nia
WenVTLYLkWjCWCJDysGjXZMTE99qbtn04y3pYqEwnH5l6LlEHe+VV1rj5TTmxC3+
bItSYGxbtGfAQd/7aa9mKUs78aw9skIcOa64lbYTGwDs/HDWBnptlEZNeI4krdsQ
UY/sDHycOKO5864oQjczRG+Hfkfht9XsUFWAK1+pHwm61NhnmSCasn5nKzv41f7B
3PNEPtEEZAsB2lnEiP67ylireeC/xGImq+AF0lBLsndID+ViSa1xDpfGlND+g6WK
p5hpwbXQ2TNCyhYhkU/95U5dWLnN34NAGtzypiCfc1mXRjynyKgWvHQcPkKbwjm1
zS4ObQFhJshCy4VLlDHHey5TAPcoTNDVgaW/QoyJF5BjXEI2jxFhVbxCW3DsPuP8
cmR+GPpq1f+TMpiXqWaiwa7xTY49ctqxc4xSXKPLliqY0XKIuMSjPdo+luSEEMsR
aukWwQyLVW0VHuyR/Db3Z5m9j1XJmo724Z+weG78qQ5MnNLVSUrAklyraah+96mf
NJ5UGqPKAaup7OY/Ueh8te850PDgS1hlF7W1UIYrRAaKfoGoeuRL4ILWAZgFQM/C
EvPuHosE20GARFhoUndiVFzqdYjPSGdm0b/qPXLB6w/K6WnRoURZOTqEGyoJ8YBB
2KIH6iYe42ktD1cE9YRYP+k51VkSYxrHDBXh9+ZC5zuVLlAf8SZoc2gIM6eYAFXo
OulB4Rxj5UcDCg3z8SRq7SlnVQ+CyK8DoqiY3uyfuOOhQFfd72q/CsAQ6hTR9eaG
l0fM7B0q6IlAANcI2jOOD44x/7ZkzJA5qMisPWtKu4o/TulJl1yjwb54Wlj3qam6
tpZIgPJiXYxNMrcmYXmYcoA+RFlL847IdF/i2iZZ8qvhMzcBLxq7qoJToE1jx9As
4ygeBCzRd6eQY+1vNbmBzUwunVNVTlngnQ/JD2dFyrE9L5ns29EueZjZaHg74bx/
p4yCC9bPv9fBxYbdt+jVgBtoL7aJdWgECjY6/ywigEmT1/+AnL5fivJx+OOGrzTe
gV5CFnISx1laF59ETWl7Wmwv67e4QhsvH6OM5PMZ5aeVt756WPe1ZKhZikdTtusL
T0zPJPS5sw0vCXZYrP/DkFcN8tSNTwzstSJYAsr94hpWNVoVv2Bhyz9c9gw8L8bG
U69UOjwoj6auqy5FQdtUgTZ5VvImI9Dm4OhrxIXtcxS92flGzf2Ai826YVDkZ7nb
KM2P3EUYZ1mQeuoMxuwKYuiB+NGU1/kLnE7jcAiDn84hntX6WoKsMDAaVVnuf4Pk
gSOtWmGgN3GXCgZyTUE6a1AvQhmWhC+n7+A5kE+OhnJOOqzbj4E+cpZoj2SD6Tqg
Y6GWcTp/E6czDFMX4eeoS+FeRrTLccaOukA+u/gVCkUfT+gIY9IpE7UWyabtXfp4
2TI6kKLbwjJe8CNHKl9MzBC4q2/vTDIjfbv5/5tAeJdVaSnn8P+MSyD6touHEWti
vRCgLdoSAXyJdZHH4M0Y1TXCYA2hE+4+ygqf6mAU9uMqtGegplzms7GfgQVm1+Bj
9AhFmAhTgu4CrIgL0e3whivbD9iZROqZ03XuZ0hNspuocCNy7Ehew+z3DgQ7MSP/
JTSZtXR0Y6a/8AHh0NMcM7MnWuMsUlTsf3FhgiuUC1+ELOV4NtrfUeyxNiJ3zLCS
29BnLK9Y1ZPLsCDvm5eWlHD+Geb1LFzoZ+Hss2XG2RDy8P4HT3JrWfp7+XlifO47
FcwIA483+xVsB5tcz5YARe49rPccvugJNFNtHEi8LU7Yt0cJQ+UTmlb6UEIU4Ppv
NdaDO2/jekC3D+h6ta4jYmY4APglywodFH7oH1cJM/SPnA82Neuxq9GDMvIKLTyc
i3w75ztuz2DAnxd3jrH37TkuIDaP21T11VvZAHCqxCGr+ofLNSU6sVPOEmCZY1q2
RMh6JKY8CSPUHGIt44ECcDUoLOvKbbVmO+lZmqg5g9QFz8w6lKaUotSEmb16gVV5
fqLz9epClRZNkLIWer24Fv5VNItSj7L4ZvyKjv9vVtdMFmpbm757ppIPYGHwMovq
udXtXQEy8is3oPdzshM0/Lc0T+NxXn80a5G/gKAk8X9CvZG2dDHod7kGE646o/Ir
T9hnovrgVh6HYosp14SsGcb3e/qOp18MGwF/KjNOcxRHRDONRwnz1b1YVVG9S9zB
st5vURZpeRy5t+AbXSY9cfJp9rCFXU6gm0qxQYGOwSBn0hqnhHw/35PFRWCrwdaS
5qYkDADj0eXhrb09rQda2VK0adahOxYNkcQ+g/mgPxNALR9psAvI/lejRKke1Fqi
K9CevAoRpu6/Em9VZ+2tPHxGMYVK/c/EsYXCBv6zb+rhKIMKYosLWf72u0VAPfVV
VTQwqcFHie8vtIglXyUc94XZ3Pf+ndXm3pzL2D5u8uI1aAjS+MysgVSuHdePs4+v
q//XzrZd64pWUNV2gXyxuWsTUQsccLZ4YCVt1hfDZJAqX2iO0vuqW/4X+i9uPPgO
qYeOezd6JxQGVcYKyxWOA95A/p8ycRjbhBIHw2j04vCSKi4wAnztf7DCPptJuqhp
AObBUFLCTUCpU2xweGbrsXBqFd38QoxpeBBDm4WJ9UThkRlKAW1xACZU09sbS0l1
3lb9zpNNxpJ7qnWpOWuJAgcwdN6pYPfn6NmfAjZKrG3Bk+ODalcPNxrjXj16Ptvh
HDyvgp2jJz+9A4Rfx32P6n/m+gON9T2F/TETQcfojTx9g+ppyzW/uRBE+40WuC2e
tBPlBOx8X5d88zs+Cbxh7w==
`protect END_PROTECTED
