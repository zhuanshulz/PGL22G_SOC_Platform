`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8y0XQ2SSUSjvc8P3WA5/k31WlhYkWQeanhh83FqSLfoBF/1Q3l4lhddLhU7/nwAp
R4gZ44b858e3oToq02KdeyaXIicr8AiqQPjf7oYcrkD91j9uueBJgxl/t8c8qbIO
8Joz5C0tSpymgaIg8T6LxR7oSzdmKJrV2z9tvY+/hPsLwH+U7NzwKpnJQU65mBve
uVpOaQ+LkcdfE1YePw1hzPgWhdFjktCttsHwJ5zIqBbCxvFeLYa8RbgRHFMQQZUf
iQ3lV9ADf19cFuKwRCVsseSdXApi9aHoiMREXKhjHznkyy5/DBoBgvQb8wg+YKEH
wR2vNFojK1UX7znkIwqqe5KRqaHb/XD/caoSVJL5H7UVra+ybikStOo5+nUn3Flf
UJPH3ePIhJmOqM9kNSnHylRAVCaLhbfVkMkSakieAimg95VSVZbS85gpt04FQztw
VpKmF74haa3xmNiy7ZeS2Oc44SeclKDVOADimY3ymqrDlUolV7bwEQBtpnGvJHtX
h74mlnfj+3gTd1Hdi9EY5ZR3jj+Pr8aKvXFkocWS3srKuH+MyK+3bHKQSFZRYRFo
8NN1dViHkBJffZFGy/RDNraCjdmMEHjUGgwn6OBwKQ2gQNZPEUHXBS+6oIsOvZpY
D8D5e+4v9MHmMYO7UkA0PZA8kVrMkLI0H7FP6PIZMgwEL/8YI66cdULClFtvOYu0
cz1Z9VRg2dKpZ3mX3Vnf1LrY0dZa6uCMjR7F+DC2zr/7dL/rEhnLpQgZ7XXgaqTd
N63K+rZ9jVoWrfMlB7r9He83NX7PB8Fyld4i09q/nmo9cFpF1iFl2bhdyT+pFg7d
WOp+r9QAhaHCUZHLgNa3OsPeJdonA05Mm/PoO4LI/FY7T0BAaHhjBg2JW/ndt4R7
r11+vt9x8x9kv+bxX0NopZqqXuIABxFBNyEdvBpTDWOez4yTsLgr+L6xfpRgU0eg
ljyubP5wPfrX2zbVwLo4LaUoqARPy5N3zKUQb3blyQ5PBbNdaUASw2+LJdanld1L
3blkiVOdV8PGGtV+W0pL+yv64KUtUxkRmwkpqiUOfU+twFA4T0DZXZTudNU9qZqB
iqd0svuzb2v/VkAugq+VgKq7ef5LUZRbiUXR5HABo6K/uKLYYZI/tynfPUnc767A
Iiia15+luKtuq9UKauABd6HFaJ6n/YKe06CJbVhHJ0PSsgMXnM20BrI3WOptxfrV
PfgwLFhZzTD585AbMVFqO1h5UchH9RF1X9NJ1z/0b5Envo5+wQEE/SObseTlB4RO
vsWkBu3R1dbAYw6IzOdP/Jvynp+Xdd410sSv7k/QFIkjU96UoTIuavfik0QRHv3C
FFxke/ogD5DHO3TAr6nlyjZFBHGh+vLYHP03EOxARgmd3gMQxehc3He3QESyC62I
FHOfgIq4HuiAsrwC/8dWetxh06Xv8cZ2d0x+TcjnWMVBkdduME/FuwOcIB4zO2t7
Q4NPinMV/n/25RJPlfRIgf51xOWtVlFFjpa5UakFipTCKFXH0eLlYT/eEnuja0jM
4oCgcrMRAOZYbS/AiZurxg9fvdicsm33aNrbbCgBqX0pDg15zCJFmDx4Iqq5+HxD
sFOWwGnz6rXqdVgRArpNC4/QRQUGK4RSfP+9FoamARbiXqRBEK2p2yzDp3X6GWEr
Gl90m9UA3cHXS1pAgHXo8GCssylZwhil5hn/VA11Gf/IYQ/Yv7TNkS8ORO59avuO
MDtPlTEYqRuvR/yEhtvuYXGCFBXJ1q8z8L4MZxwnKYsxGFlu28CmjXPPgID4Urif
WqxcniAJR7Hx3OKPeyxTxemL1yGv6LFoi6NvGRhFWnMrNvrTk6kZcjYVgbuYadiS
z8CGrCKtREsZYhp2SHOgw/rH6kzAAH9Nl2N6OCCYz3VlloRSK1rQhsM6fFb4gRmZ
NvwNHt7Inb/zfaMZJ3xZ/nPWQindy1MKcBWYBG4ZSS2x0q9xOMyiY3XoeRwpxGq8
QhvQywV5HLWea086V7RFDJzDGZyRFHKDir3AgPrZ0Hq0U0ejIGSyEurkCv/fmxjM
eGM3l0MD6rcLiUl2DgjCNTKWEOu9ix9QQBccOL7dFmH3WyjZAzZdOU+PU8HNIxnU
+tfvdR0JyDKARaDE7k6e+SBtIth9cl6eScMZsuKBux7pWs+jw5eyrAghNhbs8yY4
ddz28Qqm9lC775a7+Vw87ashXQaEdnDMd9nP3Jmnn90tGjHigljWL8MKVu0w57wK
NWICf5NnQ2gJ8D+b97P6845zL+FeigJfH/FaQeWdE5rR3fmyoZgq+4KOuTM/RORL
h6oblUMLdju7a7WqxS1iz366RjDRNOcwwFL8k3YJPc1l/OPEQE7rdBKdJUdfrVrU
dwS5he7OXjlTyXviti2WCmwnoHl8YR6nLjFOSW2vz8Vqi01Qo0RATSIjwl0HSQES
rXLag1aCZ1m0dlCHDSxVPsRY2cECyvPhcWpOXuF/J9N14DEadtDqr8s91xkzvJ9u
ZbI4eYfDbAPnpTaTcCo9ZhkCiPg9f6zRUJ9eHQENHn8n8B0kvjxP0ZA6KE1eWEGE
EvjjdlM13o0sI7wT6rCp/jb2vDw7pTEr5U0+2PSFlvKjyWGfeFp9C7TASTXH+VZS
5DiAnt5yUmP/FFZPcoIXergPUw23Q1AVD+jEALNUOyxjidwT0vNZt4cWKD9OdS36
w+YF6lLapTbH1M20IqPrJddMVWwb+2yR4iAU/Af4/mnULF2bh+3S7HPuUrydUb76
SxXgm039E9/++kAzWF3qGTUmAk4sTgszzdPCdM8YAwr7VPpm7beUc83MLO81E6/H
76etYPJvslmgvDCxbgkGNu0SFzwG/ca0g1YNccHaCxoYPbceJs0HvpE0DwA3js+i
9MQm/Bv+Cj/1kiofW3Qhtrhocqkqy8uJcOEiKwfg8ZqdHX/PkF3zbbTj23F/G9Rc
f0m5n6x79vwlNa6laKKfuI608ueDy5aHVxLFpc7xSZUKV6QebpN6wqiTzOZavcKe
ts6Yaye6Fwhr4GeRe1gHKry1yq3LRj1Q1vREfJPuyIFfS6DipfesU6Sj/h+d/ReU
ZXyNy1f0Df8JPoWFL533cN+PwpXugq5W1aUPIXkW8WCPTVZIwJ2z4lA0DndIpmIA
qi8wq3wDj0UbGNlTYDL6XnYheCzLbRpS4wscFjnyOybpbdoe4491kSPPfInEyNZv
0QYG/yU1zCFElu7tD0WNysvtFoHlpuiC6BDPyVcwNM3WeTOQt3bJn8dLI7yE4F5l
tA4xcdH5Nm3AwRjg1js8EJXRjHzhkRHtwGGeM1UF/zCL1qcpPoa1MfSFfKxyoKYS
4V2eZr+HA+BHsVmQXcQy/vX9kLk+n08K8BIsRFbHQYAB2K3Sle+cHEHT2E70x2tT
LuDWS5Okb9eQaim9Qe2GVp9mCh0i6q3rkzHP9u4gkqlDlL5+lpChll0tHY3JfRMa
GOLdVix6RsFcxcjVmhQk4OmDuGo6SBNmkIgnRqFJuw08FsiCl/NfBNp4C4TJvmhm
Sud3A9xvVOn/SAgSSFB+h5xhuenFgmDj5bBf7yyyCqrz5UoQGA3PYhRydJHEZqWE
BYtYRWT9wfmp5PrdeirWw9SJdx+XcRjFWZECLdxyN8RCJd/M+NfMavDdYFofA2q3
xW3no5u1OWrmxpASIjidsomHb2OM9G/HEASGtN/cRuCFasiAvnEi05TvoGVZisGk
6IlZOAZnmrD+c6UNWdSzF7iPYPgVj5Vxcm4bPy0mAvC6ajpvjT1PRafrVA7UXhQw
sDAA7TAUtl/J7DdNSlG7suA0Ki5ZCc+1ROjLe3akjWtd4uzQOQiMCdBHjSSFRn+M
XRn/s+sy+c2qT1PIXbxYDVXTvM+MVte0/P01LkISQXG0aDxWRHqagLxwpKI7B9KG
AvfynBk4o0xXpaIa2zJBg9XSWk/IAhdsyysaxecxW/Rv8/5uFKklESVwDcd9gSPC
a0nNa82PZjcSlXesTeGSdn/i7Dvku4NBZqO7EfVDMYEjN5iEMhoXz11/PhNQxKJB
RpUa9VTF+1o0TKSwJuM39GTyfhgF2VSYrLu/yzWRoWJ0sMpp0QOH0qM0c5dzHZLu
a1RVhsdIttLbq/sHVkqy2aHtmHUCa87Yg4911DVZ+cLRaiYQMJcVUj2Cd3Jx6eKE
Aw23Fbi//m/PQqMp2VLwV0D5iqWVqIXSz05v83ONTv2IsIDjU6VLZYfVJAIFfzxk
1RO6gYZGiVswr6BrS8NXw/MR7fcBm5hEbKZIHz9jg5JRK6RRtkJKHBCSCLYHuixQ
fZLQ12bMKBTUMt7Oe+DYoZFvTgKKhEkdE/VFvNGbmGAIzKnoc0IzKICr/hzb1vCA
grWSiHt9vPYG8vDQV2PJ3PoWBR0KtIwEawPekdvSss1aVssgYiaAzjR5f7B20iK1
5rjMnIniDkoCsreR6x3lFEQeKc/tT7KPBdltYrNEYGwDi0gjQf/ujchohijFMNvK
GOTBsi7yGfOvMsx2SPaPZhGyYHcY32gkhCifYiXn8dx+RLQbjTf8hfswXgcngV5G
7m9Hc87XHwrDZtofSoTtvj9j7VtrvAEHhSLvMOTHlGENUF9hi0J4G0boeBlfIiEA
5jox9erbgtZ818T3Gr+mqRlp0D7n5qzwOz3Jcq0Jn+nZ2vdjO6daemlR8C4uBrWF
7TiXdD/HpKeNQsLRtfnbFaKFe5QVXZGrPPDOT75CUhgHUMu9QuNx7zy7eR8ybpgv
YrNL+Dt7Xxr6cbQ7UMwXQ3j0UWaSyBg49hteovsnR4A5cJRW3GFWjAN04FbCoBxj
hImNDwG2y9IjWFg0cGbuihFKxlRTbLJcjnGQvi+Ze/1vhbtoVY3aywlTgx4Ujk9o
YNAPMOnma3lwp1BHeBQAMKUqHzeMbmOe/Doie9trMeUBQiGGRGugWRksA2FcETSu
/xRqQYQIFMvnVOmY/kCcb41B8swm9JFIiEfYl09stWqzPbofectdYuSsfUdeNGKq
2rsGmAvJn2StYN9kLvZBNYQJSVJjk16AB0OKl9sy0UhhtpMmAaSdGMS39G2BnrQa
xH4HteuagDJbt4URA0JE6ClIJeFPPDqgsLvVFxH17uTfizgpmIBS0ys7dtRjXvCl
GWwkv9TNUPYrdRIKkNHpQ4GPUVRp7Tcy2mjin51Ri+5ZWSslbdH5voEVN27SAbzR
v9F0L+V7Wzp1gjLMjOjbcAhgJjD5mKhJDG8o5aYYNojuZIafhS986NrW9lUgQJJe
B9cLBhnN5bq2lUaqTbPE0msejClnWZiGFH6KL4gbxYMMHdQlH8GzgUwdFwetmcEz
67FfwY9dBs2qhNMOT9KwKQxiYtnIHU1h4DBGi6rhxiBbauUXy+pATMnaYFW6Xq2i
yg+diWwX65d/IM6jWZpNkCQ2mnKcsQRCy829VOQGovtfw77BLGxtp6E9T7rxwVYA
Zzvt1J1SgNGTNClYxWgBVVKJY8FhZW1PrQelDp4hEBfGCWruFptCFz5sjSOfsmXQ
eQ+RmIfue9weul757nM08bQF973idCgkCY4aV52XQyW6YI2tdAcP3I0A2KLEvVI7
VXlCIBiVgCWvXmWKJhwWubG8bJU+OS9FJqr8ELIP9XZbqQK9BJ5rZgVKyvzls+pJ
4mNZmuiBRbTzTcHcpWaAjeWVlTiEMsz7rMn8mZ+MQRERkz8vwMlBS+nekxGjpTC5
YXNQky3BdRocFxRCo05qMbG/n18Dlxiz9N1KsQqbwvtJxvfH2PcEQzmXHgSUUn6T
xwbTwHhTUVEu+tYvi/m4ikVEj8hg1nQoMs2JpFf6+GqxP6ZYREob/r1A4F1qyS6E
ywp+yQFUtHAzHnly064wMlzFK2diRQbaPLSZqrJYb6qGmIrVbhZCLZqm+C+qEmfr
xPd14KuAonCXRR5V7wgKaxZV469sYS4dXDIDcfI/xJ6S8eZFN/ktRlZ4QsCEnwNA
n2kji7SDfKdCRHa+Tn5DpHKmSfrW7QtHP3P9oFM0+jqVSCJ2VkwkqA5LNy6zRu2S
eUI2qTiII3C2WXavvrrRuhdk06uyFU3jKfZ6SSfC16oHX+9or99xJYj8w0/MeWj/
+bK30asNHzsv6C6y1HGkkGB4QQE7gLIYDRNwefKW1HVc9dQCxenGP2PwNIhteNAt
l6jn2GCb3Z0ZJ3NSB0/pXTPnoFnjx953r2+sCqgMY2yteg4a07qC6uJDl4d0OI2Z
N5kpU+4o+VHlLCKlUS0GzsTgY7aIaawllS6XVxGKkdWAwXmPsaS39ka9WkNIyZZa
ok/qy1oZPC3DVRqBpcG6+kCRpv+YGIabTpuZzwVJPcXdFaLi+bik6AA4VEvK6LhW
iAogbUHZ3q2LYkdAuVB7mUSoOhEURazz0WZqzziV89iWUtpTpuCcuGnGZVbG6bTU
5HtvUUlP1fYtdQyzOpN84DBfaVNstDs2rIQz6jlMGHhGvYtJwUvo+jw0SmXFAHCA
G3zvzua25ZFSC8xDI3Om4IhZTGJ7pxJtJvqeXIKfDyaMdNYRFjxvYBwrRaPfHFIQ
ETNIdfN/KYbG0xfsVClifDMggRqy9SbG2itJKTI8KW++tLPdBkRiGVqPfkk0+MnR
+bxgXTnYZe2MDMRz5Ie3JGShENgMR9N8Nm6pDyy6kb+UYx2xtw2dtYsDCTsb02QY
MSeTV0pxgunKEfE9+BNXLqXQZfO2JLzFGWnyCvNni1TelOxxH+Svf6pLfKACnbkl
xd6PerjVG1pnON55ABMSmEt6CiFAjbUt5pc4eZ8gDXvlYuHfRbg04FQKp2b3a8MO
B0gU6ZcbhNi4OP0uDRC/XqpT1sfj3xwLu9AcZ2r7dwoA4CCsTRZEM30SFjIVHLN8
gWH4Ro0hJ4MSlkQTBz2czufymQiA47IIFN52jWe4DqJxHK5pCWc9quLpYbuJbd3A
Jaig+hJV5n5slgrXs04nDwJZOFGl9+stWWz6awqZ3PgfS9uURs7hQgYVWqCrVsaF
MnQEYh3zFnzCfNEQIkInzKNiXfxQAcIkcg8QFpTfMdGOOJHGwY0gXXgZNcEpltb9
70abC7U6fpRqhYp2cTZJvwI4ntR/DR8C/RytAs2r++LT5qj8iEfks0kI+rPCobKu
6lXv2/iNm2Knr+galKWSvQPRqZlAAFnyoXPClExpTbD7n0C7HeT0ABUHJUKq01m2
kPC1YQ4+oj7GkbuXTpR4WcaC/1NexcjXlmBqSkh+341vifyQfKVjz0NKDZAI6N8W
G5wslqEiIY80HD1NfsNTb/wfwSdNJ+zW0SVR6p69nlA/fvdVKG8x4h2buLFeEs9G
IwLhbD3Ax0cXYhWEaSswaaF1Q7rNlfQ5dt70iY989iMRXG5Ht7dlv2Yj7Wdu6gm3
WGMSzZZV5BoTyO4131uSP0DayaYCXs45lE0Rj8K3DhuxtZgOrrOeapHePMkVEyEA
DLmnE9Rz5W6ow82fUomFgErfUWmVK62M/urnG9vOuaoEx2S4hqdy483LOnOceFeB
rNFB3uoM93KDAYKZz3bV1WdjBMuxzQO6iXV7YriZFAe1CMas+gijOZ2MF78ViJmq
YbRS/UnUe3+QDIt9cJ4rGSUb9cxBEqS0Wn84P+TAoU6gN2aJyY5D3uKr/LRgBqMb
bc3GtNtt0bdTiZcBdWkGvoziLqf+HCdi9PTX+3/0FhSIQx8124lHxpWTqKW5OqSH
Ui8I2utlzAOl0xud1POxP/plfmjiALgNvJgXW4dyah0eoP52G1qxQGz4fivM6YM4
DIuC7yDG42AHWEI4MkTNw9c8I0l7wHHv1I89iGKpvwMlVUXooO6Fr0r3q6XA7QZZ
h0iNgKNoBad/zHPPE3jO9RLht6neiyt/ZZumpEwJiBVATLhGSluB/xD/CWjtg4fZ
YsAwLBA3MPx2f52bURaj9+ZS5hX6Tz8eV1YCKv7+mLCiemujrVxSrwJhjgJaH9wl
6v+I90kfe/FcUd1QljzWk38VhtN1RqjWTG26KxFFd/NcVfswIWO61EyqWWcSodrx
IZTMfrER8cqqHchIFCSARhxdBy8MIfRfsLXOwxqvfHWjYgSPlIhpHoFyTcLWJ4gK
UHDcDbi618/lMbgkst3hreEkY7FUhApQYb46avSmLHulDnkyEailqqggqUPkyg0f
RP54jKU3r06+dl7+RrEpQDteABNi2vTXwLFcjNjsFBAjYV/TvZ9joXkZM3WmY4C3
dcCJkODg3bBmLDZkQIhdttMN3hpYjICDnKBYwX9jR3tyPnnZSBSavHaQL4DeKDXJ
tlV6CM97FMNNwIZEmDJayaiJtdhLSv7D2NIG5dxsxFoSp4oix43FIwq+T9CbokOD
QWK4ZOUkd0XHIncQFZVyRW2brRi023bFYDcCFSOw7zjbiGaPTO1OcIDNxQf0yDLQ
DvH7uQbDwq9bwkpWQ6XM+8EI0Q7M3fXaqtUYWWUDAi7mwHtfFcljN9Cef2M8fp30
3++LMunl6KVIk9BtQ1LyiV4azT1MGz/aUqLYZsd1trhGWocgJ4xPXlxoAL7vp67G
Livvp/vf3PGVAKRtJbv4o/x40SLOhN7k5gjG1IUzH53EFzqG3QjuL04cqT24Daa4
BbWqZ34zOQx5/mok+z7pK+EIh3kLH6kl0ILTpHWGfCHRS0KYdR0tp+tPfY1uz9j2
jm6v0fQIKnhGAXbqrXalbjQrkai2LmTBeGwEWqmBr6n2cyVXsorKwp0YR/6JvR4u
Ce0YA4CnN5P25IxYkoc+chb42NIF/tO8R8iJzCfE43PYb1mYhK8VI4Rngkm+FmjS
EXJzMWrLl5Y98KcRdRU1GleGblKldWwao5Z2ZEsozQ4kWlKuYWux4nkj2p/gcvzI
lmuE6d9rUxBRf8tBCSVlC7Nr52S283t1VJCrZK1S4kLBxRivPcajPQHBBboQKTBj
9V1S0L0PN7bD9wNHlNN8RDLHOKuB7WjNT2hPRd9zYrTE0txljrYD1hrooBeDD45X
fAWCZ4kNzoVCD455g6H0GfD3whD9A8s+wnpFYplDoUXKbKafh3a+ztbmsq3RQt1k
c1TrAMRLz8u1g2DyoFu+3Q9VequhOLyhQ16zWkQ3aXJJVMvswvuHFGzFkl2QRgxk
aJZyTDuaota2JInilsHl9wi+FjbrF1RYEkrV5sGpj8iiHyeUJx9KKhtiJrK47LCu
8iHFnjfUQpAHSWDXjaLalyE9iz5kQSVbZnHbQGzIuuBadHnHWkEQttTyXUT82CL6
Ms4qyXi193WRAsrpE5Phi3O2UBbFrZNhGvqd3IhYUBlhfvVCXqD/A98hAyba02ze
Ph7NNZHEKTlq41drA3Jwzuz2HAS5B3oRsjy3JY5lPAJmZfdXXDPAPYc7EGI4NVTv
SMMbuTa1Wc8MwEDWRYJLIcfHNb9hZFnngrN5RziD9bgONHIR5eql4ja44Ewvx1RC
AIumrv4Hotu96ySGMXiR0AukT77gk/zfiP4QHK5viiAPt3uQdKTf0EcyrR0f+xSf
2lc0Gvdhnv8nf4aHHn3l+Ekyb7wBPJ9flfp4eRhQC3i78/08hYC6VreIG7AXTzrz
v420/3cjF4+CR0cOSUc8lK0nogK3pI0tRS6K4Clz0qhyISZ1IPBlcxL0H1CE9Mho
JbRaTc7sBLmgpOr5QNEMN87/L+MMfvfuYjBILAv0w38Bf2Yx3AvaXZzkBX8kPAzU
uBKXJrdetBYxkKFjKEE/fimDLOA2tfqwkxM7BeDUI5usRIw4fBR1Im1YK2v2Ubi8
ZfmI+kUpyhNo00lFg0+OELCdczbem5vh3idDOPohBk7HbKeQSeYKuYERC2+2I96O
v6gBn1G1bs3BNQxiI0beOZXcF5eztCY0lsKE4QbxucwwRt3t5/EFPB59hF4LIm7B
XU5OOu/Dq3wf6JvpUapT9txjT4dqHKzb1M+Wp7dBVDwuTIybM7mrpXU8PQ7tpe9W
T3SpNUlE6JwGgBIZw5YdzM/fOW6zV0CMtL3iPcszGUTwAynnjssbZ5lgwn4sKlKH
I/7Pt0y8LtFxyp8Gssq09dG0LlOVMmI8jlVzt05GDeLUs7xr4rUgL7U7SwEgg2e/
/xcp+kE94i8OOyczPXy6wk3eNHvDt4Pt3qwPSC4waXV2ktV1h2TPf1zhO9SNBqYb
pYIkaetfKooKtR6zX8nmbDooAD3Cpxw+h8e3XR8f4pklxzg9fd+UngMaaWh7jxRe
HWKmCYZ/UUXvDq9iZhnJ/P28IvQru3hAnmuyWWFgPH38rabXIKpeAP3bDM0PCnvX
l4C0xpCrfpmpHCixszyW5e2csxs0ytfG//VI/DCakJ1Uh9Thvvk0Ptjqm7tC343Z
eSnUilCuTD4V4H7eo4/EsilmHZvcs2ZGE2SAdbjPqyMkOQcWcJUktFwtvnVzprar
WJOJTRO4yHX61YQFTV/uw16DKQg/8/5QatbcpagWvoZZDxZeuLrtwSw+mmr/1Qhw
WvtjvJaokbGakS4EOFfkjGvDceNUam5u+A6OPkQW3uQyklXiDDN5XRw8CPxFocZ6
0cXpyYmbxkYCeWtO9Rp+Lpz/fPiV8szDNr26kUU+ZVRMZI2EAR5X6r5GuNbXgo1X
4Hp3jpSb0b8U6LMpnY8xqQbDAHFiZqrZ9EnX4txZccib1OmXXittGpm5K5l8RN5c
46dvZYjfl9fy24Mdk5lcQPnzMDGZJ58cQ/jqiu8HlByg7uj5QBIJZKjKJS8LKiOP
2zBNPOQqE7/ozMSiM6wG0f9imcfsU+lC9r6MWXpcWNTOyNbiV33ZpeVZbBL4O2wH
b4X+syvPHJb5MguQsEmFUjpGWL2sw2OtFpI1h+yTROZ7If7cmM5GXsXr/tM+yKeA
JgQErRFcQeYuPoo8Ztse8yIUdZ/QXCSh2TTYKBdHTTWwZxXR04CCV53PxaBJXrqp
unb5zqwSnKFYqnA/oiI8dMUnsJI3RbaFW4vCnAH+0RJ2jXDKF/PiSYKL4cfVKl0a
sZpMUUWNSD0hC/c8C3j2+vHcI3TvcWbfPiJmXScm1p80yG9xyOsikjosyiqigc8R
4p0XW9EPIFZloyjrKLMXA0c5D2hs7XAO9Yg4HBReepznbeG6nuuNOqDe8ZcZnAb9
J5L0/Q3157oDeVAtyr60KAgTBpmzp53wHdoUfkOcKLGXWeyPey+gaHMygL6y52dP
iRmCJfXcrlldQgje1uvw0ALoYFpf+896cHx3IUnEubz+Bp0kAGVrkT+mvirwlR4h
rvLqm96vznb7XzmS99uv0CVBE2ibAupFPzDe+0vJjFZIoz4480S8FPyY8QV/iqZr
ax1mUpJ4+nP6Ylwm05uzQd2MebFdsBs9GDcsQI95A3XEkNuiGCfUayVmzMI1Jtun
57udJexpHLP9anFflBd1tgOUhpE+v9aE7fGsblfwfR7HrarAmHnwjq6+AulvG5nN
DFs+kImtAf0DqvJ7+jYVQfBp+ZA/MuBlFq26JQuGzw1zxr2wd0JBcnuGNpyc+T0L
xRA4YBXaPgdrrOxKjcCeiWVNmCS0FZjcqFG+77SVXu5ijxBikh9SJjFcXF+oTOkc
EmgjidpQyMb/WS3nMapKY9ynTX4y02bWgEqHf1MsvrfTUSa0G6CJfcS+YFmK+GOi
6eP87qW2cS6UKkWOzQmnCVcObTkFpWzClUJqP09ovqUUC+F3qonmLJAJwbWbWG7I
pRz+b/0XEOyxHOvelFaT6GN2+T8/dewYiULdgdXYlAVQZNYoy5rCJXP1vg85qjvR
6aKuQhAH+AEowDxZMyEzNCKEzxP5bC+oSqyGxhhgTN3+hCh2KaryCV8sUXkM80PO
Y1X9VUrWhJ3I14HeiTW85s8Yk8o4lAkp13xxz4nVHBEeFL/UK6jkiA8nH+tvUFMq
WLDzmku9pmm4PNMXQ5ebJbiSbtsRf9FqGOyFU8TpYWDiGyFT3gNje+H2Dg1M3gU6
JfILzqI+jPfAkZ9k5kKzsNadHMizgySCok7p/qG5RoQ8EXt27Pyo3TWBk+kGIf4/
uxa0u3zVL4Km8UDUDTQWN/TEMB0JwZpy6PfFHZgL17ecotInkCKoNto5SLHjQgEz
ZlkaTL6tO4uAtM0+V/86N5d5Rzu21Zj2PpSpUaTltCZMRKAkZVM8JfJx3e7CqYaC
sFw3R5ycIl5qQEO1kSPvX9FxuKyzTM7IZGTNGfEnS2kFA616cKu6JnHlO/LtARaY
ZugrwH3fIqNVPdAkD8lUpg1ee5IAfio/DEFtk4VSxgD8QIi7oK9QQU5nDPswwj8/
gzYARGB9PtcFhYadMci9dgPEL6+l5ryil5bdY0exQbLPPTG1e0JGoMmOHH4TwqJd
QprEVRnBZA/EognrUtRr9Tiv7m2jHAjcsCJkp57+mz0XRmyFNFTlxkL3dyR6YXAB
ZTPXiN4xBUTw+Q0ntjfp6WySOfZFzQj7/3san/0Sr8dP20lpvrC5KPa9eaoT3p1D
5wJRrLRQMaIDS6drbRm7448Ow6GEjau7aQfIjDyXfXABrDIb/rmxzaMf3XxGJpUW
OrwQ8TCI8agrk02G3krF1TTl0l8a57TV3SKCRx1TpLtGknJ+QRsLwSzXbL7lIzDt
q3iaQei+818ke+VzYAak46fINfJAZSuVY/8ivoO22/Qsu9E00kut0JsTOqBk/AzI
MIQQJnSo+Q0DLOiaMs+naNWEV5DjeMHXJ6xAXhvcHsQ7svdr+M1oIEM+bgI3YAo/
EK9iZccMBjpxcVyCDNVvn8I3ib65rlpMtrgwfMLi/EQXA9na2oeIoaInpWw9tLHt
GxQQ/UlHGkrN/fA/fGMQWEF8fv8sG8vdLMpcg2vCmk6YAtKT+litwjgP4cqPUvGB
yHG1I9HSxBnn0D+YSkf7HdM//0lKqdRfLagLgTciR6pHH0CvHFpCiwg7tEQc+HrW
mFYnIKDyVq0E2eOe5FolajLv+ZeaRjiOpgAbDkRYREPiqkeO8+6A2oejiVcQj1So
Xqr6Qfs2B4FENEEoTUUA7Hl+aA9n+J95KASbbCUmLL+QkIZpM3G5VXTYL2FTaYo6
QmNiu+8y5U9HYzQDzgDNsVkHp9DbIX7H8kKERXNk+NVJ/wjeDgs05sPXoL6tJrCa
/zp3XCus6aIjDW1hL9rFVVe6ruJyQ2LnQlySuL/lX2c/UPb8PwlowTWbTNzr1M+W
TYJ057UkscRJZ7qvINfASKku57nFb+dIJXGfPg6bmos2Vx//Ty67MvjP6E1dtqee
Bplh6CZ7DlDaKs0BLAE+GnIUz84U9vSX/sDzVn6PmJDDOh48Fq8+/VRvWTcH6dL4
ZqA+A3UYDi3UirGvw3t4l8JkC+2uKaCrQPdDjZjyb4rVLKcCvXYfOxWCglk65rkZ
F2puvvq105LlUMcO5SlthZZo0DW1obZxMJmHraSLPbiOubhYYOPyTjYLip2zZYyg
7luJWDvAgKQvcgLb+RX19XajBDg+lymPPBcwPdfXKh6lHPJoDFhbCvqQFtj3nLuP
pxpTF7m4pIjcOr1LCV76Tq8/tsPVxSpj0IBmT43MliaeLBqDtW/B6rEEn1QBgIe8
z26c2rWTG6V2GXUg9uPMnZzrqy1M/fYXI+RZrOr2tSGXPjUVdmDKOq9usaFGqe5E
H6d8UB5kK+B8mq2TcMhxtCFyn3P55gjAgQbSfQP7xLTVAIurj4f6PqCI5OiuBdT1
jdgt9vfORscJmnuJ93IyI7z6aRy47mTYo0RFHfHPZkdhJm69lvXwHjgpgz8UB8/7
KusPIhTpNmxDnebfHvoQwl2iDhttVqLApdkZmlg2A2PDwIoj6fY7mxdrvjIujgJi
Pv6bc3a204AoxNbQIOdDGAfxX6Pkd2bDpYRqtT38vmzLvO6CJAbzTe7CNj+imPTx
60OA8uHNywwJnqEa+hDYVhaAFqzWcSc4tu7H1F4VKzUObv/3aZheHg9T44ibY9Vf
0q6Bygy2/NqL4TsGVTveYLUmC6JK4yTPg3PYT6MFuenZF53u/5y7Xl//obNQ328V
OwKAOkt+u/4PtdDixyuUgX65lZUxqmCY4QAU5r5uHdb6mDJc+jrmEtWxHAKY1z3c
kSUACTftyNWyDk9hpr+yrERSHGKdLnySwflune34HWk=
`protect END_PROTECTED
