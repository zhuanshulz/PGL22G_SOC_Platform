`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZ2YgKxs6oaYTTDGGuM/EN22RXyxEnh9tUiGBaoFAzC9E+hYzo3QFZmwHgNte8K8
3IONMXLmYrQT18J8vXrZxApTbD15ehYhCT5r2ZYTI2rB8QAYRDojLecfKT/ksxxY
TMixnjy8l2B/4+2TekXJhsZshnZiRNq5ktrwDwNLMrJpoA67/qtg3bhDV495f4Ut
k2j6CphgU9A+L312A8Y06Gw03830LR1FiJWY+pl9Ld10VqP/5qScgu3rlc8wQtEy
2GMxTXFHMcRvJ5eiMACWz45ZJck1ygBPZFUfsTWf3HuxgTQpfM2W8FKqAAVQB1/e
jOzW+OcCrtHI7SZO0O95OPwXsPZ9vJxLc2fBCEYmTJPnszp7zICcAlDIRvgwSolq
zRdkA67eCd7Ko/1hKEb1FO8rdsbbpPaDTBymhYOJd3GhSVDLmGPGlE5nDQsaQDhV
tBVIj3UJ8D/U3TAjP1TB6w==
`protect END_PROTECTED
