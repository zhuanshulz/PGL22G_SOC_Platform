`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2EPZD9V2QLcFE7FdKfxBeVBC1WDoavEAW+mxfNIxR9ksTo9QDZCoJ8N7KxIlTVsF
dgUjpSH+CQkfnoypZ9y+UsP946THzQYUiRPfnFC24vlZtqmWCSkrz3fgNq64/kNm
uYnBLLcxojhZCH5PW5GuFW2Dbwo3+PB+2Rb6q4nVRUwQGVdCrVRWVOK08ryZJrf7
JCzP2Rb/wTp+G/MY38Zj/fYo7ykQSCcMarMLIA5lIAUohkTZcDBGz5DV5RzblhRM
uSlmhGI53CGfmVQPQfHloBMTWMX4w8tqf+zokB5d26eDiN2KM1Q0ugMxgnFzqg/l
4JznGfPC4ODvvuystQFRrZDf8G7Zlc45IZIBM6isH7Qn7ij7pNyAJtJ8DTH5KeRE
zjsQ0HRHNP5cAHExLpmHgiN+gzs3Jj8KV0kwsg68ZjbY3YzUOFY/vfRkVlLg763s
PVCrDG15J7U87h2noPAdsVtZhEo5aJwoK7K0n+ekfEolm2DAT5szx1lKyZ5uWmMP
tqMJHjHLuyu7AxHlZaJtIl3TOLwR4T1dTk91WLYxSHVj6HmuevCnniaj4dGE4RCf
04cAntPP70XzsYsBxwP2AhENOAUHzKD/Asb5Ed215t7noZA/aupzRDHBcYeoKtdi
H/98Im76VzkJShXTBlYrw7SDhzGNrCTC9DCtg/+cIvcUa2jWWe4oI4iRAnYQ3bbZ
FHMSDru/w5LZqYbfEuzPX0APgTp7vKy8DDUt08lWL83hQw5td4A82v4jxr7+mDsV
g52KwDjr1NR3Fhz92B9l6reGEluSzriEKoEhSSp94Mk/k2Qk80WivwnyxKPHFyjq
TRi5xpY2WCS8MTMepWP/fKU428m1sxCJuf/SqOTAzTCS49s0tx17TczrEnARD2dH
f+RhdXdaXzMURMz/OQk3FyrTf7u5Ws0NBK88DpHiU9Q85MWg6fHjp9QGZqefNlRA
sJYF5f5lp98aiL5J8P+dZDo7uHc92yTKb2FxARZWzI7mMlMjN5D0tHIfsoAArNok
uK/Ymr2oDyFir/G78nRMbOA8evr4xzMdfVbvHpSoXFwRe3WZS9ZFsp4VtHjbDA9m
NW0pnYGKPUeKZ0Xh1nE9svHmHKlw/qGTrP7oBJtUZ4RrFeYCdRR+emMOh8GO64i1
GfSZNKuHyFgZ3dbdmJQxiYtBImyau6pGrcuPxmfZAmKHYLR2qCBAQH4RCivBRmQM
2/olv+DMIT7e9IyVtlOuF3H+6XtnVuvm/x4tkwviaYx8eFigyBJSWmuryjad5A3X
x6NoSO/kcJ0HPRBbLN7v+Z6zOt961rIUyR3Fomsqg+eWu+fdqhUOcWS8mnRMppET
XMn39sRfaCY+x/P+4+1hwUUvhfyMZgaxXiMap55axRe5JIYiRNtU/TFZNl+waBlj
9Qi7D4p17Nb456JwemRIDgSC77axqdbII4VB5rKIutOfkqBgxmJnoX6A0YtbFQGY
NstxuEJ0YqCXG3wiFEEvIPrCue8u2fHOsFUfGFyjojBskjHnRLv9sqGVN6TdsavS
Aq9TZW1d8ZAvjg9oc7hqju+TTwXsUHombx291QSqQ3R6xtIadFWu0E6CKhAqTzfu
LyMZ94jWv39Qw3i/u/Mif4DoHSXgDxr4aU9o9+1bfgJjtRmVI/zEXGDpOB3hEzI0
8scFHwUuJCLvoSs1zQXvpfTdBEgWBd9M5RbPpEEjiHEDyU6hhZ1qVUKhpZpeUQG5
LnxI5f5NTOxueKcl+CFx22oM1pxult6d6SuKtMc5K3ewoi+RsZCQTCR1F4rI8Kd5
Bl/OAE+LSrlqORP2eWJEJ11e1saDiouv3fnV3QRUyW1gspqyOmDvDqMrRSQ73208
BEdZTAIm8XbvjR2YolyUrx0z+l83zdQ6zYOkHdrkYGidx6M3kK6hAIceL7bZTVMZ
jYoDAzroofBcJumhCg90m2vZcuPJQntIgG/q995Pn1TcSh3OBE1yDp4DsmbQZUP8
439SIoPAuMUeNGj0on75lKCAlFV9F7tBIzlbnfOV+ho/gfC+pCvYAeTRShNRjev+
a5k26TsE4qOqIFx5G6dhAHVEaVxd+md7oeM77cRlBPmtBxB3daZ2Gbcq0KMplvDd
HZyNE2a0vTIzmJyS+x4V+p6vqxSYwbgBCa15IvhfjNVf1raJ1yVos/32v5mOc8Sv
yWo+BuwqDpb4TBIsSXgH4BlUS14gv/C4dEXqAi1t0tNckBSRe0Q5h4ykTuqbXCTt
PtEmHz+3wVs8Ngqs0r+OjO751FqqSq8Kaux1oTA+CXemw1xNHc7lhSGR+VSuMI9X
2IBdfiXFcBGg7u5oUFV8q2aU0DJkttbVGpmUoToWIn2+2g8TQSf39niidlR5J6AC
5tl6uCiTlKDi8Vz5HnPuUbbSjnfJhLu/kd6ngPBcW2CQeSDSF3EDYGM82FZn2+Wa
OJgjG/56mOKe5WgNY5bTZjSwkex+stVqPENhXcA4CYYCCHOtAbTS/OzMZb5K14XT
`protect END_PROTECTED
