`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVxUGzL4LQAMO/g4refTmYB8MeUDHsyCvhSliXmvmH4flLt1GXoGofTPiu6SMCfC
dBPrLlFvQa3jMfo2Kx2H7SG9MvxpvWP5ELo2yw1AufAMs/LOurOtQW509Mky3+AN
hv1hz6zpwHtEwray7B3fvzZBSFAxnRNIevWsFaMaaMqcW7uWoirPmuo9rkwQptZP
mnc7PgMIiSpwv0cLIUKTzqssNqyxBId/LEt2hfr/j4AamUED44hKlfspSATXw3EF
w7ZhnQ5DGenEdX27YSVKqFWhbRO7n8CPSsm8UcHOWtkK6Ssb7hRnbRWnTcD3AlSv
gEs6QqH1hYwc92uVPmKT4tuxbZseS2eyEEy7H/WHSHHXYLqMXQjOiVeGD/ZmocYh
JBN0pnHLSipsR8NTr4/cyZk6jP5AAUZMW6k5GW6agEKHLKW+EMpLJLB36IAD40JY
kMarhSy4DGKTpgeJaUAl9yHUaMshf8pjw0rYLzqLM70JAarmjkvDd71py2D5lqli
Ex/18Ghiz+FfhskVZEu/UT/w5XLmYU3z9SMf9qQPXz4w8duKwvDds6eLTSoEFbMi
wKqrjX8NjHYj6SnUsEpAiPlV89vSNDWWF6MY9rtKjA1KFh9tP4c9zyL39VXXpiRA
MWwCH8FJnqLH0CWfH9oiZsOxHNnCbUKipdICS/n5VLInU74tEkxWOCxlyZtNuVg8
AsimR7yp4VY/UcQTnaJ8d3NeJmGUibGHw/8E8lEicst7xEewGnIWLeH2MOQyhz87
pmqSIOM1LPZeqENYMN/y+FU1gTG2nvBMTvWbsUdUrvMBMNvqacjviGS92fGn9Ey7
eedT4lE+mMMOjQHsngYAsI3i3ruFjPFiMXocl1Zcj9V+0K3Gchz8RaizdOwRzpMQ
S5YgIVN8NT3EB5soUc25t+vK2h0j0y0FvkXlS4OfKt4OHnO7pZLEpWGv/8VikEtn
XCi9PwUqtLqr6RVhDoUrgwwj4JLIW+Nt8WByTVfE+57FjH5BqwLIGSblEd8qKloh
NHWHDN9ITugXYlnxikNcbqOcQukhO88TtZATphwQzUPePzL0UzpTIFeAw/6UGFUg
fKNXwQJvDl/RUPObVVeOs2QIZyo6bShql8kzyDSaPAe4unrZ2syVuQY05e35w/Bw
UdEZe9gG7VGKIcivvbCg0ngE8/1LgUnXbWAk+8ybKJyw9fCtE7oYQ1l5rSD3FLSw
rSlXKcSqjYUJqp3scE9XeO0WlKecO05DPKOCqcxH58h/dDDSE8N5lokbj9jKaefM
62enavsQuZwJtDvPtVgNpEjBUroOCv9ueJ/ONUV0WTdgQfS0rxF0ZW/Y4WjDar0E
P7CFpcfoJKSW+Daj+en1BvN6j3bu0DAGWnEmO/CspH5cZfT+Z13ELf+Y69AhvLTE
WUmkjdBMmOxWJvRF5tpfpMnjuodIZN7DgW22sueX4leSIbmrTYlMmUarnbIjjl2B
lNV/HZiNfSvOCIJdbXmxpce09hlF8M47PIdez951+UJ4pT84XQlCs4LIIgNGgM4b
My4HgpZJhImgkkmCupG96l7qj9aPWX9wgAcJb9CXGlMBVsP59d0pewx+wT4DLVCM
PvZg6wT1CjyEN/vL/ZlH0/1zi0gDU1Fh6d+ScSchW7LWCXrBvGToEp3+VFGwZdPH
7m54T84vCT0kVSNwabf1srotXop2McUWHy+uI78zx08x3vfr30bkuBj7rROf55MW
MmmaJ3c0Kfc1atVkp1Y/kS6yVEuLeYNo/9P08H8dHvxrz/LlgitAfc3E7+mjYcU2
Gc1H8jBTVVKUjSXAFhCEwUF7sbtyYxzzdFIx/UvErwreNqbjhR6heh4cOjCd5lLw
Hsa64IKWq+2ukKO8F2c5eZ0b/EAJyAFB/C4osTYLxDg3XWDkoqqOO1+r0g/oplWz
Uth8Q2YVIPRZ1wFT3VHkeVPn33AejOVTk6mYZ/FA3QnkJsQPB5snY5KnDD9ZRMAc
HuloqXKFfDt0vnYGSQFOkXGfnvPJMmIR8dR4Bq8RanM3hSm2hYdB+sZfctYb6rX4
/pJjeAjWYqPx/x6gNazfzt3jiDVgKCTu0VyHS3JRME9eFnVROD9z6J306bbpv9Pr
v53HYg7LqgSOxG7T/WYPPQ373h42P1OC6j63tXXoeUrVCqJmWpmMGw4QLYtWOMGc
ZjVEvnP5CqqSUo+q0bNoXGiYB6G0T3s1iiTUpv1oK0yKE0qsZGbG+dkrIKuVWhvP
LrJQ31NUGgVzv7IsVApe8sQoK+awTr9aoIgMF2RKdLHvb2cnShyPaeH9RHzypZ9e
3Zv889SVrfhgrFsHOvRR4GNHpANIlhX74H7H3tydk6LvhAZx+Jrb106PoH/AfsWH
9jzyJF/HIb95DlJvZjMJWUnfRhcBtwex8NtKwkS5jev6f15bUafazqCeVQAEXWL3
R7+eNWiwHKfcJ247h48rJSiDJYxhaRy2lNA1mHEzEMW/dLwOq38Ay9IcxpKxY5Pt
CAK8FFduLZxMPUqKieXk+Bzwi499zcJm6Os+rgFqJN7pIeMUPHfboCjKwyxHPxj6
EHrzi7mYZuel4MxhFisJD5FEIOhITFcCTjmeI/Q0xlV3nNCQoMLVNgJNvJaaNNuz
bhfKGjVr0L6xh0ljOnV/km4foJMTp7/5uPwlV//4M58PMdZKGyJsmiQo1Lkgivz4
dxveyX6DBMH9gk9qPjo8UXyaYPDOaiFNS3PmZK+w6EC1cfPAkmDJULCXeOIPzshj
IuOfhFtzaWbE/fhnJ2OAy/2Jyt90WZDs+qrjCAGxoqJbyd1yClZcIybAsqMBpgyb
uAQQWlTv8ARqTBAacXAzaYmwJmzUPcfeSx9RxjsdrwaLj+2rLp1NzunxyzWqaGrT
LH4KgswgoSbh8+ECJDcO4bpp95n/rBPfJ8q6d3EEfkPH/Nc0V3GIsUm7YBscgSUK
ZWc5CHy+5GbNpwGNS8fzgI/FT7TWqtvx11U57u91t/fS6B5JXU3V5OYwkt5MhH/s
lqa3kEWEnXWVl9cncQ6BBO6cS9HRUjrsSZZdux1EnpthkzVUU+7tvuPSFyv15UCE
r79KJrWODwbrglde5OHVP2jkQ6j+KsNufja0qrr+qLhbZLb+c+6hq4dPX6kGmYRO
YHvU8LQB51h64piTlkAMK6uE4mxyMeud2KIqrozSy6x5ybArnTt3rwWMyEVNE53P
uyn2Shke0/pUnamoy3jJloK7T4l4icz8YxxC2e75+2i0j81xTo3IKecFIomB3Iiq
KRDpTtKiTZ/4LWJvsdWc+JYgn+AXKn1PflVf+dcNB63ShZytE7hytSTbOhP/sR/I
uPRDn44swZXSSb6S3NZBS0rR2OFOkN+kVV8+R7gsr2lC/dbmcatGm7ZDbQ2WcyPG
M93VhnSFxYkAG5dRMgW5TBlvlo87m5eOQ/6FLYYsmVU+thMOGlJLyiZleX9ReKsj
0odIkg1Txd+PGzCVO8pkHDkjQW48xM2PKVHyqos+ejO6kA4RyR6wm03SXLuKAWNz
8EfAT4vaRhkrPPVcMYgZSuSMxGgLa0tWetpQL98M3d57uZFH6qWnbA/HZEcxAU4s
P2nBviEGP46VXUvPu3GVoeIRgpW6UmeQxLdq4g9HOY/TnaI/9xODtJFdZNqWqut1
0k92OjDKSGBy3Udd4ZKX++RrO6uVOKOU/IzUQgKNBk+PA2h+7fvg9g7CDuPIJcQ/
BRY4luFAzFkDGRtbs/xzJ1W/SR370fTGxzuJs1rn03AlaWM4MG3ljsjc8IiGAObs
BqHn6a2C2BsgmQXXb+G9z1Hfwbl16zGRreKy1OMMIyJkG1MXPFLNfKQZsjzFteNm
X8zgJVq0YBmmDaRKQJ1z6HRyyJdX008h/EB/lLQL0UMPaw+SkQRVKjnZVjLUqfOF
gNJGa93IjPQDxfXUPMAVixJp+hBb4GtkZLL4fWPiL2AuOj+di763FoF+jl0GQGqr
bABtCJjzPKb3Mxux1mGBXc3pWbpg0iM+cpRTSsrt0FGAnDvjXs6zY7JZld9JrM+3
oAFuQPa4Ur3TvHHzgQx2VZqvRiGzUzSMJqfhjv0VQp8OAz+gTkm343tV5nAOr5E+
Fau4cXFo2ML3aH+b0RbEWVMjWBQaNB/9Eijs9TiVWY66H/tWrN4lnixy7jtdcU8W
1EuGnXrMSzXmCITtqsOwZF6fHczjPlZqYNBQg1NRN0WUr5JUN5VBKCavcbzO1Ytt
wn3bLM4loRx6hdSu/7m4EPZ9H7i83xBGklBDlCQg+pakYkCmNr5hEdWVt6oCZevI
cUkjPhYoYe8gIhjEoZHwhWsv9DnfpF5ksdrRe3DPtvkLY0FXSQtgP5PYRQhuWO2i
fodgaYiBJzQFu2ytIZM4VE0pZyzF8epaQfwHOuAhLCMTEqqBK//Pw3WDzXiANJO0
vnXLersoExKzWbxPdHxOj3tIFoNITDk+cw+QZjFMcibFP5C07IjwDl5eW/W2U3PI
gkDiqXmIGZ/YQxthR2DhP4vDX7WZe1uyS97xg7quIqhlOvam8xrgl5hu60f3WoTp
2JdlmL3xYVSXgBBHdTd+IxBtdskIVtXHfxmfXjAZgLPZBiQ4odKTlddodVkbaIuM
SEmlkMdI0XIPob60xa9iN3MiLykGXhRhGHFh63IHAxWp2/v6P4Q/IfBpa6N5ljdD
`protect END_PROTECTED
