`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NzgZ6l5gJJusJ8rWk/Amfkf7pFDPeCPd7vpJFxfqSMRq05LNAx3NYrq7Toviz55
U6m58TuQ8MbxzjwyHu7OCqG2x6PQnD3MATL64W3NT5dfwTwunP5oaoSp0uFwtSFB
kj/G/DwEHAkGpi5+HjLM8UxTzQD+WXs6ymcSr4y+VH3MRnSxxjAXj2XiPuN4Q34C
Vuo1as8VoWWdl+Tjxhyk7hqm4b3KhPdkjA4AlBzY4ehhszrbnFixccymFkw3esI0
I3/R3TtscPMMiygd4KjoXAQHKsyWRYj5ku4cYFLfSStmxj4o/x5EQo42Z86djrcN
k7/AsfbZuSd69pR6PsYgpOUDCbUiefonbiPx6tkc+ewsDAlGIGYaVRpTpBxybS0e
qJScoTImolCiq7CaVJEU0u7RsO1FGlsf0FAasV1RYC6n11O1lTo4mss1my0Go4xa
sJjghaC3za0lGsJ321MQuQCCvJ+8FezTxEuLKEe0LqFTJYdJSSsy2TEgxTww67Vr
IixZltnHVoPSy61swtV1TdXBJjorBGaJUXiQvkN4pbJHKVdU5GKoFxh2X90StITW
u3J5HqcYR7MH5xbDPGxcZYAoGYHYzpCLLUg6QUALKW71icGD7XPyclzgX9j9aF4a
pfE28so4zY7HC8mOjX8nuZRPJ2zy2wPeZ0C94A5PtXA=
`protect END_PROTECTED
