`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+JIjost6UGEh7457u0XdoVwlSVX1cGDISSzC0rfeeWTjry+eBu3z1/ZVEqFTsQH
2cYFssQWlO/ONJ2rwE0A8DTPUSwnR08N3T6QhMFud3qt1GnaMYmY9CFgTLlqMUX9
fSCxVMiSS6XCu4NsTAXgEqY4kczpqhHbYgx6YH6oKIukbMvn/QrQ+VNFLiCHVuni
neFbTCkbzAlqwujkNrBOp0F9QLneWtyfl6vB8wmoGcCMIU17yaUT2l0iJjAosnGM
d1Z30MLm5llmU0lRt2teNKT1ARsUDqXClwkFtOfKutMm1ZelvWp0EHCJarBNnbkg
LmTpF1I30PIpukSO7wt+LHgPEn678xNpggEOhnhnWGFc8wQOXixfOcKfUb2ROkvk
PJmvBoQYeulHGpJf8CDLNg7tdRzp4BW4u8EjaYREEbL2XP0kYVoXE42ph9/eAWVf
1nczCs8bk1hmezgekBMLOhXPvztBnH801Jq7aINM97yOE63WhvZqCvJvOz0Iwr79
mTq7mH3jMkZff5besIGTwA==
`protect END_PROTECTED
