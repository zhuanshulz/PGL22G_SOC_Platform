`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0giworlhn9Fj+9R61Sw0c6qkNpMGiXWpZ446Nd0m0Q8JwcLUbdnn8UfNQU2Cah4
BLJr0y1MFRh+OmRCQqyogp4dMZq+EoiTVH00A3HWoE082vzYSCJnXYc6ylo+d16Y
pOaIeByRvxdUKWkBKLVIOxOA4l7BY6PadKraEJfWVFMSjX2EEPZrjNvvWw/w3VJi
dga8XbiIC/iRH8tzVfg8zerP47OUhf4GLrmV4+aJD9vNo0Gs4Z8tBvc/acRNFaRo
y2O64IPlKieKfv2Q7QuXOMrnNMVY7H6zq2f0VeWPJlIRQYsWsHIxqJteu9VvXK1d
H+FXY3fgPi3W/1JA+0n86xGGwU7O/RfOsezvQGIfML3jC9P7HEZLdLstMNmuQwaT
X/+sOSNSY6lZ+OmtWKzXuQVTst56ZKM5Xo5NSKwLNZm687ifawY4aAirMndmBrE5
u+FXW+c8ikqB4w6afLSo7XZ4EmUqC9MkXmPZ8oXboNMb/Vd6lV7D+jAy2nBVFpBX
5u5bvu3CdCU26DOShVRaituZL675t1mdUH3w5iN+/6gDNXB3F8drAk+Fvf5c+lCp
+S71NdXGgheVkd0iAl+yHe9AB1dXTUov/L+b1kYBn60=
`protect END_PROTECTED
