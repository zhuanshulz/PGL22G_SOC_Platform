`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AZsM81UayHFDau5PUbd6aBbysJCmU5CLMR2BcZZkOjpswOFeU+BmYU78K3sZDEBT
HQb79ok3lKMX4vkCTcnJQAKC7QdnOUAj0iwgWVCiCCwMd5LcgR1M+mPUI4e8FUy9
ls47UzgtmmmjNlUkcUrIwxASPqi1PwwE7zdoGu2fqvd4sNAeNY65NpkvAykxfier
yXH7dDzcTldd7jzIpI3Vs6Lr7KWwO1vyyJyPPcphAuqyEGfbPb3026yuCwuGubip
Ob0gROWvTd95u1L78DqKbDNx3IR9RqNV7cLtSqxzsfsbDDhkXxQ6UQc/PxWnv534
LaVzQUoLS8R+z0Y7RnRny1nY/sfsiUwzS0zuNDmLeK3qjl34d8nOYONG3+UJm/ZQ
DTzY4dXjHNRzvopOZqom1nfCen1M80m3tGLw5zszSVwwi0kC/x4QTwA+yc+YtSnt
qb2jP7m26Gz9lgvRSwZtl6HyyDE8i34BVjBMM6if/L6GIzBhrGcE7TlFNxWjQ0gA
1jBQW1Hh4LbEH5bwIFOOSy72nuzwDBF0f40BvpRoCrLcQbGB9NO8NBUvNru7Zk7l
gOCP+/uARhT9En55BNTmoDxGm7eZDGS0UqKESjvyijH3OvVtIFrDlWcyIqSt7b4l
I84pjpm/JfFFNMvF3KiZUll1sercR/DmdcmqujHSG9M9VebPhBzxdly0da0mHZ3X
cLt8biNG8XgY/h7ZF1bBGh37VkpG8u3V7FPdv6ZNa4uZpUG6bo5D6rZNIr3kgREp
E6VEUhSrKUrpD0wkRfdF8WP9XXOKR0RQRjqzdlJuDc2xIpVqVNUFOP9bTkVZ57PA
hgNkncgsjC/Eia6xemGSspY1iopTLN4siYyBLEXwxEcaQYcC2neMbZeKqvglDAG6
gI8bMD9VlFdGbE7Qcs62d3yKZOPwlhkNCDYngzJKc3Szfmjdh82XMNFBSGpE/3Oc
ShULPC4C0e8RHZjFMvUPb8p/N6xSzdQCel8cTPXKqCmcS9abxXw2w3M/R8mPWNSn
QTaeaq3FZR66TSLlPpKFEQ3xMk4yiGQjPkfgcTsjBfkd5OTSvtyqwo/YA10oC1WT
WdjWcBAe+snkbIFR//oruIlw/GE6g45z8QxOcubiUzOz/R4BC6+T5YYXS0eiZNd4
6f6nut+2e7/zDSJse4BSQlKsc/N0OTC2gi04acI3/ZM+j8NjemMLa/MQuWUvju2W
nViXQjEzL4rv9a4xi8S0DAqOV8r4xYx7TFV9I0iFo1nUAJvyWjT1GB5T4Rbrstor
YfJ5QHgcRLPfoxJi85w+Ql+DBxpgvaWhfHMivfwPwZV4nREGqG9Nxw41MUsKfr0C
nzUTI6eZI4wwSJahgKEDxIJrbRUxjOuMojhm3d6vw4TF8wMe7mFNcWa5AD40zYG8
g+qTzawsCERyGh5o0OV3EBwvtuZMSj2+3M46p1fBTRsP94xkNPQuMGD1EOuIDwZ3
cwH5K2zJ+bVTqD/WGOmz1qYhhHU7S91S8EfK1Tj9FY3Rsd1XPrVCS1harsR7hdM7
NtXWQBBdjOb+ZmEONYvqPHCvmb1O06/uCyr9+bN9iuPmsUek7JGaIWc4ZD2u8+an
Du5x4YSHBK+/H4f116LVQ/DBy5bcl8ZNC2S0eOOoivFiEh6ItzI2F7mJbAxQCCvJ
ak6l+5gAxvudLkx2fmdYpjGwkCScyUR3brJgQZElKo8LOrzE+e8nsdljoin3eqR7
bOqg7LjPhAqdGjTjJDK2DFgKkGwX7nmp5ea3y5cWc4Ob+htTiNwQL9DjF5sXZtNu
tMBzXVVa1YuqnIHxVn+lOqIcwvXZiSomwfTNMbyYcRVByAvuECbq201QJHNBSkdB
AzEH2NhU9Av2yZSfS4KKeaoXrPivVbj3c72r5pxmhaqzc+cFTVInJt2Jf/qy3jt8
XZ3fVuyoQue8ltXdUtJB2u5Iof/RIJIzk3LP/cVSeEiyZ9Y05/6FO9/0pb63/+Zt
q8ZLblrCqbNyPtLM+xhAbua0q69hALLaWxtpbP9aTPn+wGbxV38Cp6R7ZRXcDk3u
YrG3i/s5QWeu5FK1UzDXGN7sELwjKIR34pg0Hw8v962oTAey99KyXxpOmZ2orbaQ
ay3zdbjMvGFexCu/Y+u1IOSZHACvQylqExsU6kYsV9Z+HU2rJHZfJtH+yu4pDHMp
FdKaZFlTdj30gemP9HCB26qtrPM2927Bq3i0xzS1/5KSP/XF+U1AVL+Hj8YagzFo
kpUkQvtFpcwhhGv4tsRslv+oiUzRy9UJ9GpEBDL6mh0BtHQwfXbHzC3916hCnQQ3
FnWQUW2mxQlOts+wevoyhoGzyT8HxHUIPEfiMhC/HlXGbhKgEQLWv3rbCuUfyepd
dpXVRAuJQ2AZBUJp5Hyma83FCNqMPPDB+7B6Y9lSaWlocIALXcdFsgrc5inKdg2F
8/pGJNeI7nrhGIfDFSQh3djCMrImtAEOyGx/4VN1oAdkwi8P5LEkXNQgUEERqypj
dJhwy65MgQI5AhtSnLx4fTLjOu3KjTuBTUApGH0tVUJo7028aXqP1LzK2xcca2ek
xdQo1fEzRMkzHZD23ZznP+4h5+6j24OGi84ahP/vXzNuc0otZmQlve9QP6nOXklX
w0I1gOMsE/WEeymH48GAQkDqijCuDG4ADh9/mYNg6jQnZyhl1tSHFblj3X9KxkNz
z0ACCEFUeYaf/E5N9tF67wUUhdvHbshNv7kGbmPcD49Deh98qK7TbUwhFv+Um4U1
HtbJgF+iM+Aj7rIOp1pB0mlCI/i7y3czvIDJoBJZi0RGV/zxIqW19zzjKOQc9N5n
NqPiU111kaKGps76NToBthdO9RrPIXIqTDljYLrei9/deOmDTbec1Ot+5alqhold
gg4UB0/2qE1Pk9X/hhR8Yytps8II4mkrfpRHtxWCQWuVDtZyHVpQuGyOQYE2yJYb
tMKsUQJoEnPQsXEQobPJ9BQYzP4y7i8NeofgToM6Wb54rczkZFv4G1YRE4jZI2Kt
HxrjYhfm1SW4gDy1rs1F0UArPkktOBktvRODK0dNGW6mtnd+ZtXKUGOb4Loj0zvv
7SurSiM0ElWiIkq/M8cDzsnyOll5iUo4vm6nYSCCyf0zwBsPtkB6+VORVDJzPLUL
WuXhJYc7DFMch9B9kEMnWkf3Ku4VWoFLGzwAir6k/kTuGZeBlbK6/FvvW1M7kXWp
enbDcKiRbWPAtKquP+fI7qJEp1CEHeAjI533LhjXVs6bQZv/MUkDjI+0rpQ/fjis
rOCZeshB3JAJNvzjAgqTqmNhVi+hor6CyHvea4hlcJ5DeGocwvYPFW/kgD0EfgmZ
rGsBa9GYXI9lq0dxb15v9d6ggn7X6xkq0agAyxxU5bQrHkpUZ2gPMV4Ppx6I1oIO
pGxwRVNJy1W5V1lbOigkAa/BzitO+H3PvQbT1yJdibP4SMI7TQRklR9/4vEZr7AL
DgI+TllISO1zhdzkrmeHbGzKZfFopun2nl/f3bchMcrN8dymkno4QmcutDzzN4+0
vGr+VD8dU7/Yz/+FqlqlHg7eY9CrYbh1Qxo1RddQKMU=
`protect END_PROTECTED
