`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esUYqW0bNIHYe+XZSsk0y4VmJWj+08YWd9bdkr/IvLyw+7a+4zzJuh4JnwDHbREX
iOvrh+wTRGm4nX/PCdpjQpRcG8pZvqtUwKE5mSEVcDCpaommG8YPNSFFNW56X5G2
U85ofj9tAOFgcQd8F44/ln7BSOoZPPXa8x7Fw0ixX8xa1E4MPR6Od1pZbbCmkwCW
SgbC7FxMNkiziw66SWYoVGs0wbPmKXNtVYGOgP+7NxE1cvLQzCgIF8ZQJIDCbl93
PUUPzwIode1ABg1n5mo2MKg5mRcfruDnQztO58yMc4PirGNHXo+njZJygRTX9WoY
hvu6mXi8CKRTwJ9c2RYsaLhT39DXUkD8fpLbUwmOJ1Xnorp271BT67Zla9wH5Z+j
6epTEoQcSuRp63x/VfgDGy4X5ETn8vXTp3kqUcdkwVdNQQ6wEssLTVobEw3s9Xlq
MozyxtOwGdPqqpjtbsATIqzRoE+RbI2j1wTCk1wXCi5yTEVOTWG0FZgGjGbZWSjw
W+cOv3i41BpgXmkATVqOdvzi9LE946DM4IftrsCZ8whyeJxGstALPuLMlRVDcQsv
cLRGE3MnkH6l4uLBq6Prk0fqPvs3RX7xVZZeR5PVl5IP62mNKOPBwMzEwOKYxpXP
SvwtfJkz5eJJ64yB7cRuhJkQPdYZEHXNNutMmRcVCKc=
`protect END_PROTECTED
