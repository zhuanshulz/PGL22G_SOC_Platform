`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUdyJBuJ+YIE4NqRLqvcml+Aw8Fux27J+YmLrkxbn651diO84u1f3nsvBvq577y4
mnGxws7VHeWlt4LIxI09HTjU8nStrMxscuT27pTc/Load8ODvnJ9+5NOd7D+fRJm
CqX589n3OV+lrxqdiRwYDGgzXQODVjI6K92bUKXUlk/jXVmyYwlvCRkIuwVrtU5f
HxPPlJSIG9/lNOHkL2VSZfvoM7u23ODD+65+jGXEjSYNf6plvpnF5DDawro23UNE
rM4ow9ncBh3a1vZqQTlH0YO8Z2BmbftQmwg79b4GDCUqfBF2uPq1mN5gFZidOSIg
I53gtwS1tZBE7+DwYTrIwMJdTqkfk8GMBhMTfVKG5WXt7oE1nCZfzwcBVfyyBnsi
ur1MsJFLNhnrVQ7AbIYD+g5dXnCDlJunZ4I8TMds7j27TWLl6ZKDmMjoyPwB2f5O
aYv9wsUO4Yv0G53khM04KO2vE7Y6Yrd57J+UO8vLO5z4X5Q3smPOrT5UbSneb4/S
zn5KEeWqOcUSZeb+/AG7KciYm7ueyVXxBA37UvoOECu65a11DAgK63fVk7xoru+k
8MkLr3UoJZCyTuJIE0BXwKwJZmk5Li0KIkzQHJBS/KswNMtSYUZXZNUILRtzKeid
ECKLd97mrF1b21RE0abb1d1Od8S7uMi3Ee/sSkMZZD3Ec8i3E4OsqsjVWPDvCbXs
KVVQ6YEiGxXeEmkmIK+vXWhG2IaXJn7OMIAZMt3K8Oq9aEDEnx75YeRLRzKIWVhf
NiJjo0wP5x6Uhj0GwgTgkmTTNpsWwIEEKUWHeA901bTS78DOYVGkq2konyrzK1tH
yU70HCNmku927+fGjObaGRA37V6Zg5tzsQHSjk7pqlDXIluf1r842/oy3Jc9oema
OVHClGFV2JPRGe+gpt7aenamYE+fLxZJ79o3yaEsJ608eh1m+RrVcFNOLhbLuc8K
fSa+6vkiwflpH8tHhBXMFIyurEPwVKWAovAFrdNRoLxU0oJTOIDolBQjtdlUxuoB
YpnoBGflY3u0JgDkZfsGsYqARn7DYASViuNMgkZS05/tczK/HqLYaFzGNc+1SiT1
8jbWiKOICWVnehxdtu5efK1bmOLfIE4CB70qqlbdtmitGfLRNfaRN/4jZ/FOb+Vp
3mysre/QkeIv8KTop4LOQPXPzkx43t4Gup40vYx/35yWXuQGS/WecR9YaOoygJkE
tP2NqG7MAmoCQ44m/fSr7LeSGW2ZtpjaEmpAY7EXAdX1QCwR7apGMfDY1Yl/z1fS
IqlrYpG6acQtMy4Bte7YON5NpKxpWHPf54g72C67wKCvDZBPpw2i+QPMYqOdYVy0
U9OHzzKx9stiF5GZNsGToUic9fOletG/GnADIAe2WuwZikTnuJ7wJejUONyYzAvC
cuuASb7GZsTXJBymGH0e57IooAkh3TU1jTVRxpxG2aH4XGuwcSove9TA3crk9pHx
2avbkMgxotY3hbHPWXol35egMvVmBPDXyeAjSbD7o2+E+7tlQGDIJdy6/ACWg4dI
UNALyEn0vkaeVxFFCQLMIrHX3gaUNtq3IShaAGntYBECpUeR/b7est9FUkbU1D7O
VuUrIm9S0JiG87oHWSXJBbooUea3/MuhX3fUgL/kwbm1PtdmO+U5Vi5SKv9abSAM
5cCb4+JtCVbtnTFmQ87cZsO3v7XKN4NeciFJZrHN/FIqsmmHdvQPiIQR65WPjkGa
o1y1S3mxZRX+ILrnCni8cOczpZW5Sf94o5D9LH1zd0adRrNm4DCZuGr4GikeqCiS
IskZtzbKHSzYomik/8Z6PbLts8So/gmCRu61a3MSfE2UwjV37RpRy+f/hXcIuOxE
lYz9jG8U7hb51WEBZxYpxvQjo7eIgywDnOwrQKm+VAMGkz2fP9PC1/La9ZAWr/RL
dbKA4ZpB//GxI49YcaWk1ibVQm6LqJO6G6/OYfY0BMIadl8rNGlv3dmXdMG3Nrou
jSV81wYH5c5hGyaX3lsMPsPG8ar5+XqUHs2CC7zzA6pAlGsd2sG6iWfS6mir6M6i
Dm8bHP939QGNwgeXyJZRQEa8z6T22ZG4plxH9tvx+0UwvJAerQqF+mC7Rm4axehp
RCslkMVeVo/aq6qGUHS0fb4lFE42HfM0hNqvNR+IL+wsWBin5BNimbV6hKNbd3Cn
S33cMgefvEwXPduHZ5VirCbkLv9Uoy/xQwg3JxiW+h6BtFtxIaRGF5jlE8vrUkc5
q+3GNnD5lRy1XC9nTFFpK3a//oSBVXEVIch25R7RiHrTAYtN3tNMPdA7MBKELApY
TSQsM8peoyRvuXpMa1OsYTIUuchJVXV1W40Pjt5trPpURrhpY60A0jbKoU/mHb4l
ZHiTy5GV22qYfn6rsCtsS+VKQe81a4iIhDS2fyeZJpyZapc53nTVhMI+n92UmX9a
ixPyelWbMR0njq7un0sNl7nPSGCK+CrC7SQVtdgC6+ksID9kId3grtDmYvRLSkhA
6cCqENQYjva2ki0NLj/8YSFEc1a3xu/ukK4ylBPSxWUAgqkbubGqcdNVdy6FswKn
inCtCQ37+JfSFnUlXxSgL5GOE2Rj/SOcOZ0KSuztG8t3KIGqGJSoz580yFJBSEzz
JPuv61+qpZIXbBXe0Hn5IK3Qat5bVbU8fvs9gpzHq+8pBCCdhfnybaWVJ9arNYo/
zuUu54y6UrVszIWa/6BptKQ/6QBlVx2hQ/Rc6alU/q6++vDYnDWFJAPgK62xXQUr
BhPCvyWVEajda8V1qvPf1MCJyDu4xeuTwD5ZdPimZLItn++uSaUHHGa44B022Z1h
IbILl/7FpROP9Kt/dSf5YD5TsLBMVPH8oldQTnXizLYNr6YKR3oAlFEiUBigUfbj
FLivbXWSdFUi5OSbYQsDexkc6puZz1QdE+i1/ckO6avakVvRU+TpsGBiI5HUWE3/
m6g9uXCWBVXjim8uXOK67t6ef37wVw1QwzaVMhogJQU7MVgloQCw2um9vJiUnPEb
9BZrgPsQuj1/ujxaSk0OODJLFfb1FoVsrfyOKjLGefBJcjBUMdmN9rK68WdBRs2l
Of75oAJYsE9l21MmI85+mLkzLL3EPrandsLkUGF8bx3Iq1hCoq3tfRqMeYrwr57I
9zkmfmUc8naJyN2tWaJILxFNNYbiKXvC7Pmj2aGlGguob3NwmShcRzfDReXBnN8V
pNJvo5Mn9yo1VQtXlhSwOREZkK6bninGpb+1wJgzdrYr7Zw9mdvkZyC9yYafxuxD
aMEhZb+jFBiqf7O5Pm7Vn0o0ZutnRXXj4owOSOKYzgaDYaQFu1ZQWrmKYasK3fcX
upSN8ntly1QjE7Iwvpv9AtXAjTqnbuHq/zqGIyadcUIj5OMNn/lJOm3EOmpROusG
AF1IA4W7nVO9QWeYotgeod1ssJGeu7Gd41b5G4kOaMWIAvvuI6+auZrtp18w4jg/
pClbI0pFwLC9+cp14zrER1UYsqUrqjG1W/pvsK3cHcm8Z7yq/D7N55Z3K49Kbcte
xTmT4r735fU0GsUK19gWYH/XsJvKKN7BwYwWdVQipPexslnlC1xZ0gL8X4bwdJpT
a6LY03aN27dib3Qn5tKy3+hkEwFPdt4Ko5HDzvwrCVTT4hw9cl93XlAr39M4Pzo4
AIsADTzbeiN+qmSm43nImddS9JE4JhKUmpKfCltyRqWxel+FtRV2cWs01jlG8IMm
0551BTOgB2DD7e3/gk7NOGuMMYxeyKjPdVdXdw94mbhMKAU3k45iBb4oTa8ZVBj6
I5EjkI1b7bFPv8f+JliOC37cdJ6jYAbfoi9Ffwfrqfdr4tTgchCKTJjRPK5p/F/Q
QqS6awzK2EtBOUlqGyBllewXmsj+JALlyk5SIdMKSOQXzBtNmlhg0Hduq1Vu3mmk
ZDmCcnkAvDKCeMHmWp/NYSYfWA8Zx5bN/2jid9g0f4TS23PU0EZzB0cYuI3QiVvl
AGl2aj8//UGXa2wkmE348my/Nt7MUwceGPBGKlTjOcd1nQ7pzyxMAKrtHu4ynsfG
xqloHCvGReNHkGlb9eTXi0SL51D2sYV3x5pi+HV2/26lGCbpOjWhzLB2T5NYavzu
CU5u8YxwLcZxNZ/YtM3SfNOXGYoKknySVZGp6FowdxxVymEEGyx40jv51EpcnuW2
Inmy+oebPWKCGXoJe04QLRU2zmh3oB9xMTnSGkW8IiiIU2TEM1nuRvv+UqgMjG+e
CtD/+ohxZxo1wLkyoImjwwsjgd5ehteqDfRVuKisAcEqRJdK3TgRVVEm1pKaH30k
7/YIa9irqhb1z/pXZHrdUbWZctIjgnkaamDS/cwG3Y6X4KBK7tVmrGxiuZCme9GT
Y1xRoMGE1hK/WNG+94U/BRDAvIU5ZAoEQUxfPIxwnAulzjnsUIH9DZfPZ3toACf3
urq3wZ6F+r5AF2RkFdqtOMmyDWNGQ8MCmYff09d9nJzzu8T8sLRoCBztFnuesMUi
mnPN2NMyIOXu2EL+67Evv0+BPAjitNIRAlLJIWlW3kgngqpTTWc25I87YErWm9NX
COAdqXUZyjztt1CNPzQSy1H7nqVy0CcU/zgepeU8AaOmWsikk4QvhhlAR00svGVU
ml6jnqQWc/cEi8CnZfkiecI2MPV9j2ak7RkXXYG6uacm2YzXXAvwmUq9/3uksM5b
reiVk8kSdnFGMULMlF2PE+BoPQfwiojkmCjIZw2EhyfsiiZapvu/BV2q0h3EdNga
DPHXFMH44H8/+m+Gei7X8XtibLKAKP69mq0oJG4oga5sJfeilKXg3ewQ0LyYH1rT
rSBJTlGQFdreDVaZneqdWXM1db0CVOYlEjF9T7FQW+yA2R7OC9FSUR3jdMuK65o8
jq4nbN20YLkzvAZoe9yC/LjEqahCICjXK3s+6s0/p9xNqQ5vFta0k5Oe9OlwPINF
veRTTfUasHMj4ooMsoIbMF/w344XQs0tz08GFkNI9RqimnBNac+5W/EpoZ8qwlmC
`protect END_PROTECTED
