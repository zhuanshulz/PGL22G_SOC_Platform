`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGVH+xn0w7XrU3polQ/HtImjMLH9O57mCD3JpOL70o3wJfHCROEfrWO/XdcjMk16
j2E970QPwm3DlTymnBDIHYG4PS7BDyKKYBJMc7zIsIffLF5O0eRY2pGPyAOSUZGB
+vv/VAi3a1gv1tPmzA2HJUEclxrKfqo9W1Z4QPTFnLYwd3jBdozmwDMsVgHtCOlM
vJ8TtcFL8FmAgIcReNKjzzah2YB6L7e027G12PMiRzq5D0M10FmQluc6zBKvPsXP
DUKllHANEZXWeXd2cmGkAXkjor33f5KavDHJbdhL0Efj2z+mOnmZq5oUWbyYVJh2
dy6VhQHPk78si3ftBcToPAHaVpmx6vVfLYo+M5mZaIwas8NbYaZACmHBNyFCiuIE
C2/ZmsTde05J7LwHpWWc2iKykoXjgdm/Qah0ZwWB7SslFQNGXOUogQlurigPhaAi
qVTpum02GSOMWgBYWZSQ7lGxbwJUmPkdthiJFkNEjvwVFCSdEADbUYXbmm4/QyxS
9UdHL0pDLXYkKjT636Y9Njmc/9/7hWDOp8JShpk9HM+Mx4PT7z9yqSst0lUbNlEl
q/JS/frkdWpAYZbWo0XQgynCSibtGG/7LiohTDzhkAvMVBmydtSNoMrZbKIIZJnp
E8lCE64U8YdMtX/kaUAT9+RQQDRw4+Xk5cavD+Qst/+eAmdhz2f6KpYSKoVctQMf
h/SAIPTCDfuISVDeHtOhuYY1vuDTl8tpSmGC1WwBcZWfV5mrsc55MsC0BBuLgWto
Wqlkxd+QzLO/+7nxI10G458yAstY1F2u9pZW+296D3VsWxMLxdkops2gEAh8PjsQ
twRiC3+1CWfMiULHvUXmzopI07S6CYaV91hAL716kyOpuROnfvr68Epmc3gLNrIl
k70uZV20xfjsD7dHrYpuH7/wptk/HHxaJx8IPOeUsGIXJPtic9S9teIFKJuZfoyj
`protect END_PROTECTED
