`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgE1+1vyJBl2vQpnvvnonkFkPR1TiQy/DlzHE61tTYiEx1n2drb1gMmE7gopiKrj
73o5Mzb7BUoXhvN6p59Sra4nVByBFBk6gGXXdRANSrduZ+jeCmjJahWCWRDPxq4l
m13bkBu0iyFta6UgIxf1uu2EEz2/D/a5w/xp0zy2fNbEG0LsFcLunQmN8V43wFt9
7Yk7V+/GVqWZfIgWF3x+gFhIXZ8yqIa8GGK8SC96ufs5nsDW4Jnubx82yLxaSSuN
M5dm0bJ9Dkmt+/B3PSTvuqaaHN0+igHHJhPqRM0Q3XYTVR2T9/z8JgQmnEEbBe/C
JdzcrhbMzDu05iFyqJDqDBHiCCxCZt9q210Z2GWcXjVOKBpHlP0EuEZVsv9dTGI4
ileI5qgXg6fCliNFWgRvyOrk5p1j1voGWYVhHQB7EzVwy4pIzpwyLXbPBLoo1I/O
R7LqDQ5elz7r8PilIp+GSjxQRe8KF9iP4zYOQ8U3zwHE+6PXTPydxVmFe/GZDQho
BTxw2GrM5JCC4Tlraz41+9WqDrll+GNTqN2VRLh0tgkP9anhXek/Uz6uhtq0bFtt
DL+iR9LIE2uT4jvDXDAS48vfWo3zbGjIY2lPMbuYA4Ugw+B50z19hmekUJ8YlYSO
mHXY8j91XMuT43h0M1oGLPLUGNEC/0rj1JhDkosWwXLPFc4BFkkanZbJmJeq2wHq
7aD89oDjo5AdcnzlB1z5TDfzuuO0ti+wf+zKwHygJRf5P/HyMdRgHGsYfoC2Uyst
pdAH5zQXtb/GrLv98vA9rOcha6Ri09VD4pCvdQlkC39ESf+ciVKDQ0+H60PxNuk2
PuKK+2Dr8zrIYnqHgL9sRFFFiqqzJk29Nw94X7u3zT+/mxxFeCugLhHy9ZcWXDNd
8k2pjexDEuhcb2xXo1izEKkkWRiXNODyVPLyPeWKi4MbieGPFf/WzfyBDBZOADmu
rzILwTvLPzun8EQ2P2q/PwtXdK84eO6LKZMqjIdFi3Wh9MjZDnapN8sS99FTGIRb
dWenqt9yL2NzHAWVIZEe/rpiIRk+rhCj9Ucn4kXovnKONxu/0mY8cQj9jyFcLz4F
XNIu3KwYKN23MjVe392gBxmlSfzBXm27KqSS/tzLCso8juU5VyaBamy1lFrAjzlT
eA3tO/oSqZ+50MvRRxvfFKit4uBOPEtQ6llsu31PFLIO2nj53tpjfLjiljorud4U
jrmw/i2KkdLDYECL9SqDRtjaacRxjYoe9YOPCztdZz+Wat3MBvO8XREbl4CFwyZ2
BS07Umf5fmEU9/wb2xPWmc7uqG76uaJRcg56M31SleMubHbA1YGBDVT4TNB1ykVk
hLyo9h8KpChLYuT2xs9cqbczV0Sn4XLksSwPmAcNTB3u8EF2YBYrTruixO4Wy5BT
sPl0oE9jKJNE7V8akEnLNPSdSBbL2UtDLYoMXXNGod+4MnQ/TwlmqWxnSvrPWzbL
U/WbS1PYwE8k3f2lJldD2eQD0fhFcVbDiXqPN0h+JDrPKb6QNfU0mYiSKOulOVJ8
HqQOywlG3dGbkyLgRzlo13Kn0U7NM4myaB655KkCeJosSiTN3hKetMHWjp9wOBug
51YKSMczpxdF/k79Pbw668C5ip8Fh13VGt41tXpBMUaQd8Q2kX6k4OekWn5GSWgJ
Cj+eiD4fAwW6quxEydKxS+OMdltVIt46y3NLu205T0m+u9PF7ugWUXaZmmd78yUA
rlEUC69Zwyhbap4s06MFKnptbBj2xbHdm+MbEOmZLQtLgoJqZHhRmSwdHEJZ6q8N
4kxX1t75E9jvgyPlcsE94eAm02DNa8ZV2p2yvVjRbrxMm4gSQDFCD+JiD4fwjD7l
c75efEa/hWUizLNMkZoq0w==
`protect END_PROTECTED
