`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s326utTHdlu1er4ROTY6Zxe9fi/GRXTfJWuGHet3DBniRSwrUs0WXap66Ytf9Zs1
GVfwvLh4eog1siKslDP2iTiBS595zy32jnafRt3+e8PKMq7ysWIQLLZX9VlXTrsJ
VUdAJU9kss4YFsRnSIHAbq+0Fq2n9i2AYL9JjYzcHnuQp2Xy54BsHUKQhdPVPbBP
X7Q6vipAi1Tk15C2NQAQSaH/2o2WVfFxS+I+2OXorWoaRMpRq9nACgmV6UPb45jW
i3zEGEh/f6zSfFvnC3ZSFP1ZI2aOT/Jiankg1jJ1nRuSO17BiHUsKJL5N8K3nbmb
RhQ9QyrNLTwx2bcMJ/Jw5DS2cjLHQTvatMgxlMn3sB531NUBUyCu+DlC0nAaRQPA
Nbh834dQx0gn0YeChUE36rqOggYNnASvzCPRYeKDVoIPfjAFuXGnbHQfsna2bv6u
qj943TYQlF2E8xJz4N1DUiibea+crMDR9yeD33So6WLBzF8WjstgTXYItIL9y6HT
nxEVhIMCp83ChBqo+Fua4uraDZcL9jO2GoHxt2GIZdkdS/3wq94/tK/ggHbb7Sog
QBcFlPnrR64ru3K4RtFXEe3/ATcXV1KezO7BeM0ZfBxAy3Qy4wto1VBOTCW/nrlj
OsShNL9L5plkkPTsRq1ArB5HynXqV4kkUrS/ZqkQWj1cZGFF9YDMM8GKwOyqhMcu
hLjGGEAkqGy/e4zFP0ieuDp8sWR+HPj0McJ6ashxwuhffRfkQDZvh1/P0jwJzUMJ
rzIdS3AFrzrLCVWE/0vCMw8KY0/yz+z7fsshKvXL8bw5NhXV4gJVZodtPvGODTWj
Pk/lOIK67RFZTkNsIjLpo/Xie3vj9xNpnTS+N4LR4NQHXiZjTe01zNPokQH04aG2
`protect END_PROTECTED
