`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1p96FAcYCbFiJXHEoclBwjj2Gun8PyYR/1sRxnVYPSE/hV5OFR23LPed4+1ukYrk
/SUWOot4XVPA60HACgTId90iaRZs94BA1Id8yeQ4J7lowaNYozXFye09hwbMbJGr
xlkpq4uSrcoSdn9io4WzaVruBbiDBYg8RLa1iXqeE0yY/u1gpoMyIJ5T748EAUQP
Hl97qT1UuyU02/pAcMc+upLGlXr4B7iz3HPi+anlr6Md3j/T92AzBOqaYbpxp6JX
nVwY5CD4i6301DwIDUEVJaTu8WA1wDoRbwNbdVt/QfAZhkEjn0CAl/O+izPK04ti
FB23N+ON2S69jC5PYJArJDzyAOCsbWhWfvdmZzmQV/49esforAN0ntA4kQ3xwzJP
59aGm9hvb8grMCzi0oUEz1NoW/7owuaEZ/jDk8FszqjkOuk4vV1qmEQ6XBsAMLjZ
hzOv5c/9vMUGrONdDAKniImUNaSNGAiBvFDm7tV+1cV0jm9/ZanG0hdzAlxMRQML
Q38Nmt4aNmrzjvrO0erkwe/ti42TymjwJ2Anj01YsJXctOOHWCEH5Szx8XPYISbP
5V8pBFAEe2W2mobn/x9E04jLvL9Lap4oc2Pe4YrRHYUzCaDd9KNMu0qJXF1KKSTx
Xu/fwA6HPcTHaGYWN9oAbm3PkWARtUePxswiDBVomvgIXWbloje6+tA54khIPQUA
VIAzRkuWWAiF0wwYUgJgbPliweSabdLbnKiEXmx0ZCgeCkCAiSK5wLvpD/GlnTZl
9DmngGfb1kcnObUzAV5DVZf1nt6/iNb0HNlrCPN/7h0N5Mo7PD+BAJ2x3dTbGbk5
nq/Igm9wi9+zBnGQEOdJ5l6HbNW2JssphT5beA7HV4gH+tr6/cNcArqpfXGf5qOi
Xocj54GXLLSsCoDgRV4CT2Th1YwRKATwW1pExS8J1jrGJ2QFUz1qfDvDumik7Spk
tZkVmBaBCIzCn4n5L0XcvKHkrrLHIbeyfPYwL5EKCpfhWjIXf2MwIf7PjJY2Rdhd
/AG+Io/4fqNUFiC1bIekfp2EPC+BL1GEjxkct1tqJEMUoeX/09TkcMAvqUfVYYQa
CtM++oPyXi13Ctsn7spWTwiRLCTN0UbH3wXUH10Ws1JwOyd8lpAdfyG44XJs/VMT
cc7YlCaYuGdVoaE17U9IAb3e3d53oOEqRz3Gv/zJlNgeorXruiQyahzkUBlhFLJx
kP75L7WS5PiNU+N2FZaKomq0ueM8ZMiLG6/oTBw1+Suayp1JQw1bcVrhzaFIpYL6
BiGWBOqqmbLcc2+Y2vJYZrXQWhNoByQPD7rKCHUQH1sJiXwjBNDYbId2I91aC3Yr
im9s7IeCqUCsQ2366rNQmQKDJ5LL3wRXFBD7XWhiNyo8B/BjcqVLF504HlvtxBqy
QzxF8SMYcrT4xuFvQhPuFKEejk13tS9jhCBa7IZo6Y4SJhLHXNHT6kvyw5AKRtPd
I8P5gw4l+ZOnb0pQa/SwXC90gfyvdpc57JNtpF+VaF8P2KG9JSskMnLpwy6YG4De
/WTOa56xIo64F59ppeGjbNpi/zbqcL7G3r9h7dvRsXzc7F2xSArR8JH9p+q3xY/M
HI9LRbXCQdYrocaz+OcWCjvVXqat9TiFF5luJRjDeLmN83HqOVA6rXFxpPbf6bOs
hahpCF8KJCJ6XfknhV3OQHfYJnmrN+VXApzz9Byllf0VCe0Jhylxndbpody9dvHC
D5m4Lvpuhp1JxGpJebSSRUKseFX2mLhia6aNXdRmLSiA2TGpJEhjVC0WmYl+CVyN
ecalaasSmfJw7/BOOHal8a1HK68YRIZnAAPvWs1lMubFb4Zz9UDCK1McVjkFTaVL
afvmjIySOZRP513qzlL7QLFM3H7fk+d9tJ+CesnGbBXdvbod+1HfACFYmPefe5UF
6+ga76hUG5pxaF84qiHOC7Pc86Jr9ehIUS6cr5i9CYTzM+wjX6UlAGDf2yiMFLvo
o6oJJO0MeFbntNz5Esa+llErnl+G61e6f16WpJ6uNQQarwqj8kXBiMxD7g95/KDf
b6naWg+7FQI85NiC3m3+AHuZmUs5iE4uFt4CFYyDjqEjZ6YVsSD7mw1eEJyC9fz3
uDlryVNzRnbSZqPMPDhaTI82YPW350o5N4Le33yBQYGUUeJIlM9IpdXoiScoTNZs
Y81yOSDk0yxppx2yCmBnpVj5w/MiFhKnVA5QQlGDB6NYguDmCv7nf0BcLJEAhU65
tfUbkfhfnOP/GrTq3Q+HbUHE6B0Zp8sOtqExymBwWw3MRYoM/TRCr5hT93m74+yv
8pADxRsFzh/xjkjDBkC/em5RDUyOtu1BNfWGamEhe4iDR/3/THzlDilWxq+mtOex
le5ALg8P4ZkYd9bqGK+hBfcp1Qba3BdwfGthE2WMhaJHFkgJGEcIhSFUCTU27SNX
1nU6qd78EtcfQ5MnUNJOeAhAxAm0homphGjUpuhQExCizU8EN54f9rLPMO6jqAPt
cVXltsxWuC3i3+gORxRqQRNMua6vQIaurtEyhTcPQCjlWAIwfsillaP8jd2A4RVx
IueOUeRUwgHjquewVAscC/f/j8r0ruspPGwSLL/DCwegE5z05LBtDkMSir8epkjJ
E1jYvOfQ+9jZHDwezxndjVUhgXev5XiUd5KTUt4LfvWg+BnKw4BRPOwP6Ed14sj/
lQnaSJEkh1x7C1+aOaLS6ud4h2IAxYTjkDASBvcddsaQvVd6LF0INC+YdreyWYG9
ibWw5F1G3tjBE/nNT6ERmzDMRqxs72666FHyDFvtYMZgLRd4F3j/+LUOOb1ev8Uo
v8ouIOAUaF+wyYY0MHwksrKu+rsnQIVkHnvKn55eru7WtaWSn5swfDY8hIasC7Wd
vWSks2bBknD/RJ4boz0CdY3mkVMp7R9IZu1s/PpxspWfLOl7x7sA5LoWVW5DkNl1
+g3b0YIR8t876KyOObxUy71GbcVpiY+qLPbnAqHR8rA4H0BIyc4AeNAdaFFnIvOX
+sUh4ERM73ZOOnbqYmNUqLM9P4pdZY98NJWIvV1rNrjp7BZQYQCAJEWH4OwRWYcw
DvSE6B7IBNn39q2yy0k5mW7nBp9xCRqgtOryww4v+MIqVDrJF1U4Y3mBuNwa68Q2
PDMs2f+et79O9liunCZXIBWFnY8FFwbVnbNUX/e1mQ7FA8B15VSX3w8WCgGKsKg5
I/PnUuqioWtcy8In9Nt/F4/EAhER0UiZFUA74fm/V3rISKYMkJ84QU+75oRpMSu4
o+3YUGaN17KqbJXRNc7FOu9GWsSx/E1yZbM7Gpq+jhyMHPbCuHhdfzTDOxgg3q5i
Jbp/mC1KKFQdknjveOStjAwdIj3d8EYAzDDrxF9BZGUjYz3ap8XrVVfc44dhJBxM
ePBiKXnegzcnxQgFQEc+epWVL9d+D/92VlXLWH8y17AU1yq7F9a+iNr3pBEh/zd8
8IQp092zd/mdgM51W8HAmkR1zeSt5fmHkuIyvBk5PS0wtekRfrUHUPf2P0sWUNtk
nh+3+43ldYbFAffJkSBwGBpe99sMEpF36Sr5/i/990UheuxIePCo1LM7krhZGd7C
C/YI2OIXXkpf6xyBJfEljbWansHfaCIe7S06iduEyjIcKt4qdSUQWCOh5WgsvzWk
BI+c9KrnEj/04/Mamv5FCWHneGWETLitPTngDGLFEh/jlUZUGSxSEw99D2bmbFSO
5PtEmfI/7TdqVQkqnB0cEUWYcRmrmurmRReVTiyjv76DH+Wuwzwj+OUcDuLHOMYl
QWEKLfUnecHjkhFVewYC69t0lSdbZ42DBxftImNvkit9tg/2xgzy/lPYZUh6Pg4j
oZVv6fb5JTfXl8LqbUE6gwu1xscsslxxiiOMLIKdLeN4Wp7bUOdq7dZS7sCBiRI6
2Uc9yHpQ9EMips4X0wsZdkn66d7JeAJqUqfJl/xYQ3auv4HvSbYnegxJbhGow3hV
8pzdt3KDcu6wm57+qhRGgD9124hgVDXsvx1sY7YlHgImDsMS2HqU7HFKF88edwjq
0qYLHeMiaDRwn4xG9oXsJN3UYTxThz4bFyVQ6nF0xiyJ7PeHeOps3ax2oz6Y5rVf
RqdS/+L4sfB/OHCQuaeVWOXgAtOOLRe9W3eRYB/KTFlbyo3NyELbL0YAUirrMVZt
W6NSMVim7befMmxFg9I2JMeJYm1i81s5ELfhUOy93HKq9pGK//z9EoXrqZxQucmB
OZXrWpMaIAnWMcT2HU986zxqX+tJmWV3vtuquykld9gVXKEbggAHZcr40s5sNci4
na50Pt7GQAJELPypXge/VD8w5e5qa8DpY8Bl8C6cul+k6k6+NIvfPVRuNkPMtltN
ACwlJ0uv5Vm1sIabkPZdZa3wSzsDFKPc13pWwnn3pQhc3SV2wqUQp+FEyXYc3SS0
jGambpr7zkpWmS3PlBDpXwEOA31kTAtqovzzJKaIM4Mb9DTlrTPKOMTA8/iU3SbI
8iljQWesK7fNpGqO3tyAUy0OKPu/8seoz8R3vfnEiTSw15dTk3fMVhEXuXTPgl/r
2+zhti4FEufpgn/J0PRBZ5Xksd/Ia7yLXne+/Ktbq1u9lg+Jn1x6xL5Zs7YiS+s/
23js10cuhPQfa0xAuBrRL3wP5B6j+0/hDQgjYKaWush75Nxbi7VA5h28rdqUOLbv
RZA67ESGObVYyQxmRDTq7yant+rGsCFEcKQlVWZJV3hIW+DHPoBxhljQ//voduE1
+efCIy5b95h9Zz2F2zKWWuLbauwzLQOsZc2a1TH7FjU2nT06mcLQq+rgRhpnsyv0
zm+QvJM8h6VDierIzN0wJ7uUsldxN7chHkvWgUHkLkzFa0ecjnS3wyWxwfVkCG7i
e73PqFMtFTNWguo6KNYLOhFIqJueV8KOpeeseVD8a2/vcOIPqqa1buOysIVwqUgx
S4/ROPnt6TCLSpirvEjFOzecocG99cEkk0w8SFwH0Ffc9Yj0vW9BBk83y+r5U6T/
gbXzSj56/q8xK/TFKJCw3RTBZpJ4F2ELPP51rXHLuhrDpbpfqGsE0nckBxlBkEOP
PlN8SDWbIR0ccvD1JMMP73cWC4G8X0BrkciJXBwf6EeeuMdgBpwLfLOkCb2g3Ao8
K0YWbpEBRynO9dlWurdiTR5KrCERcRwdk4eM3vGXK4un2ehhAuwxF1xaYmAYGveo
jSIT0Zfiel6uy8Dbf2xPu0P1H6R/q6hn0WduKF0y/Ags78QbalzdotccDEed2gf7
kpKGb91nYZ2EVSDG7xrJTA3BBjCvjYkNc3N7ZWbHJZhFvch8B4f8/7Ld9mbkiKMI
dMOhPzRnhx41v0+1JvwHnvfCD7zjfu3zKekweOmsYLYugTanwZ9Cy7hca4Ce0C93
QDcRXwEXSZnsUqa6Ju9XwfeHyWWWMfZME1THqJlbcSQXbhYQDH6x+c9/tPZ3SW7Z
9tSkeWG2RisVpKdYCCM9IMJ3b1am2a1TSFMz+DNR2GupxgcYXqyqVHUAryID1SP7
AggugE0a6nww4L7CqaN7e9qxyJ4qQORfWHAQxy+f5vbG8woRnTZdQfK/Rf32at2W
f8K7RwMHLU824b8yVK+R42PWq7ubZKy3W7Zb2PXZBDoDDMWL1xCf8GYR983BixMj
gCGTAmtiPEQlcmsgudFOt62j52AYziUb7t+iiZUgk6VmsKIwPc8yLQ44YWIDZGBT
xBneYrQWmSbdE+DTdANXqhAmfs7jDvLiw/z1BeiPpVkko2GqEg7Hu/pR/0tz/RMR
EEEbZc+2zZ4gHWvCJnRE8tBtTQ1FkkuRwGq59ly7Fe/yxrLTNhX+8kD0iej3Zbp5
1lj/OVeUzpHwpbOBIpHACmEnUgebgRs2cl51iiwjcODlVoVd2RXFAwqMZves75wn
f26SVvKKbtBZYBEeeKSjst5TkKUI8GwnohH1aFVk+oUqEkLGUOlx6X4rXyPiXoWy
OoD0jmDShquq7tb96xC6RqsmArVQ8N0KUIVO/Y6Ln7JvAct8yrW9YO9oEqqPvElE
FDoqnIdzPH7ZOeCirt2ydhV5LHN5VnnbT8iaA/LdqDKrd4elwOr/uEu0tGFrHz7B
oLfJ1k88qkFSn28P5u9r0eFQdwO1eRKzUdKXIVMrnQxj66oA+4wrV67O/OB5biAs
5Nd4kMrYBlyjmjXVwyU2myDlTMbMk3HKWTWLJcvoLvmvgC0IoI1qd0Noebu3Uh8M
GAiPLJPfhjuoJcJ2/Rxe9xZY8Ob+v2kKisNXKZ1JwF/cnv3oj1HVZ8ez4rM2yOq/
26xpiI8mJJIoI72719FxUNfsyR/eVTkEOxNvlYfTeTzJfK6yAMcYWWcRW7vyyFLA
JCNUOEzbHaBgDu4HE7m7F7DVypVnKBZLVQubLcoY2w3udIVr6JsiGu3wb/AJPi4I
mejbhuwbY4FIFS/RiNO9qA2hB5B7rvJcaKlkRsI82+QZM7y2UrFFF83h0+2svEWt
3KUmGmk4gONghG1AFaywgI3w3r4WVDFxI0Y8i5z5cHkUmUnBmOQRRuw/801T5iwF
NgUFHNjbi8vVqsrfIhiuI9g3ab+Fgx4WUJYvCx0cL8ivc8PEzGWBpwdgJGXRx8F/
HzHFQ5I+NOMVVdNjU4j9Yu7eY8Mjy+6Bb+s4C0wNcUyB8lvNn/OpGcoCvew56Ghw
XvoFqJbUp/C/V2lkQHEfjQQ20HrNBR+lVTpkzcWmZMMdMuRZsHHwb/jpkseeF0Fj
8ADkDpUSQ5en/upIRUJafVRGBD50o2nzxUAOKgGqiGrd+4/EqK49aUbmfRwKIRII
f02DNxfdGwytHnT2ExEyps4rQq3MTGbzyt4uoU2nt6YOIGCs6gwWCBZEr95IrixX
//t/xjFLUZzkGC8J6XplwEhjMtoKJKtolhsX3SzEyh8GLhOtDmhO+OlDVkyZ/zmx
4Gv7cEyuErr3MH5HrixMPeojMe9AO7Z3F9I0tPp0FJuDr00RHV7QipEqFx4mWw0A
m1e8czG9H1rmDclpuzxJy0gUMpX1t1LQ+c11C9LOjQb9uPwEEQ4g9B1vRwQi2S61
fJl6mjbWhKONYc1pW45maagfye4jOb2U/7kk2o4C3MGXpAxv1Sqdwsltsxtezbld
eMOHPoFmt+cTKHmec6Br1bqgOpPiGyNHIiGX0YJ1ioLa6FLLKoXVekARoYRCJE1l
kcGEQtX6iOCVYlS2D9PQL3a2YOAnnkq/HFFT7yAmeUlJznf42TkUAsEZbBOwPNy9
Dj81tV8w6PnCnb5ud8IMt+tHmX0hr+PqtYsOJ/jkVkmjWH4U/eZMqwiU/U8K7+G9
E7laeogSCCDKaFpIQcg0m0Q1gXCVYkYuh7J5c5rtqYZ13G6uDnYefGY9qXokeSuX
B8YGpjhrudCCbpWzBH9F4qC5tn5G8ApZzlcMXm9w7HhdguDqJJh0eSWEhE72a3ek
sM9bx1UeTczWx1LwlfYJC4ROzEdWOigU8Vd8Vz/XwnvIYTxNr3VMXuQ6YUYyzxRG
JMtn1/6+4kHbilkB/bPOrSrJg52kNCkgfxbBrtYwai5sqo9Isl10MzaiEuynmRYv
5ybO0mRlzDQ/Iy9tKG8BitaqpDhxBWbeg68oKPokTghtNNqbpI/EZgDrm8mQMznR
x1BBRxpoJ/ey7k5NvPyWKkzkj3+bc++9zvSXTrwG+29oplPeNtG3lmR0II20wlFQ
khrILfN0+FydszpS7cMjDWH7LV9Ql0K4lrtnFeqplDNT28jncR1519clQHRDeFL2
RZ71MckIUKu9GE2TaE72bJGo7deXD+hxiEnnnl+ei0DkeGopoEyUi4zUZkg1QIGe
EFrMyc2jDLA/D2/+MkJ1a0ulXLe46g2LCCAm59kJLLcuuLls0u9b8VMWaRB9waBD
o1SuBRiYLrAQ4dyJMw5qyQZz8tchp3THbEcilSPVditHtXiWrH+Cv0B7Y7SKvLDC
B1IhQpIJ7F6Gwe6Nccg2s3Ks17nqMk4n++IP6vyeT7xiSyNg3UTJGiY1bbLHYbk0
azs42c7KnTFBdtgdvthzzDScVBO8Gj3aXc4AguUYyRvyEMN/JFDDBaWNszW0XzzT
AhBJyu5fZNcK92EQGQ7nXooqnygU5TQ8tcZn6ScTiOoul34s6ELcKwhu5FGouaU2
Pj8p/OuhRlDFD94UiVkMzFGYLtKlH/phooZDWY+O9aSB8Y6cCvkEU2Q73P+g6Cjk
pifG6zvH0qQWbO/BNZpiam944YhgAc1j+23Pcd83WppW6r2Gdas+JBAHRHS27knB
vbJD4KhKhDYAkjM1sekcP37kMHJgwmLFKdqPBotMdl6dIGVsVgPcDXIuxBERp/vt
7cnFSZOtbBbxQahNOUw/1V7m6ROo0YDGVHpZE7wDyCGBps1owUS4zwf+T4hDmnSG
BfqPrl9IrixjfBATatWAphPBIU/XOfH8x13m+oENY2uCsgsUXeJL2bah0prjRvLC
576iX3XUr1xh5/TOEvGsuYQpke1kqZiOTvDxN6rBUJbREo8QwMfS8vwGlCaF1bj5
GyzYMXQBbJ8WIMwft4cR94qaq/b8CKtmtsaiotCFGrySfqHskxD1hlF1kGQpFuOM
bBo9vXC8TvHTOizDDsPyFkC6geMWmaj2qL/HzbqG5fISLlVvzFJBCMe+8Jqggrz3
/UiR7aKAcvYnd1yzyU/KH7z/GUfd4uiwDSRR1i29sdBdQZ9+5Yti+4ZQ19I+GE4H
yIa3JlcppR9LRG4gFJ7wprtABAbzob4ad10P+J60qo37Q7uI8noToMuZlx0AyRgo
ITHAGWVe1y2N0i6tYhOPkxpq/nFtPGt+Fw35iqy2SozIgoEmUUSWwHTZy1KshPE5
bFJa7mdXMNa0UEaM1oPRNb6PX04W1S2wPd5CfB1A5E3fsrEgtAq8pWf4E9v7aYMV
8yBgRmtXcIcsqFlzoy/QYxFdZGs7tGSCNqi3OnphvmnugtmGnVfCGd7sSbNGV5vG
zu4YA+ljHxoqP3O/D8nUbBVzEbu58VYh3qDzJsXssenI8a14mQp8OfyhmPF47Xis
znkxT95X6BiyE133QR/hUiaPNS8pJIaaLNlKCq/AVYBFXPLWpfVPFAx3KTMWI/52
CdV0B0qqqPKgaZv9tI9Khus65kZ0Psk/jPoTRoTKTi/6CY/uEi7y/k5BItPfM3L/
rBXpLws9LjDtxZ4kUoO29o7oOmKAoQ5uruSEUR+Mwe8hjJM5eMwCCURx+kwzYMuR
V90p2BECWpeL1Hn3AUtGYFalLKGXoCJvIZSyk5AS8dF73C1xa3OJljQf123acJlT
pRoh/lQ+V2FNzNZLSP68sVhE1vIop0yd8y3j1pmqHtmCsYLuU5+zkc6nV33DWBqT
tPyECogD/dKrGnw9yIrq6Wv5A/0ROUzS0+PnM8z+19h5HCz39E2rhnxL+qkGnEif
rG9wmbpd3CIj9ECiTvJwAxtJvHvwWKr8U/Uqxy3pLaqtk1Fezdubz5AbMeUoOlGL
b5inGJ+xN9aTvBecKY5THKvkAvuVcupACeaihBRfYK4teJm68sneeEej1XCUB8sM
EAjwPFTQ7Oic06HAzaqLA9QZUbymf7sr/baYa6hQA35858GjRXLw4+jl/d8lRBd9
5+rton6wsR1Mmg0voI0hOPjyvN4FC1x0rqOTDJ04/PfMg1tOLcq+eO+ZT0l+VHos
H99XHeXjvZ3gd39bTe3plQIUc/edGoEkHPTiK43ADhUt62miCB4KdR9jo6wB0s8s
GweZl7CR0a1EyhX9J6kmH813oaOtDCUlQxvLhkgeQ0hgL3EjNO/d16SL3aRP12PG
HZPkEGQMUrS9lfalySWZHJVfnk4Ug8X6sCy9/2djpLKFIpsk7DvP1GkiZwcpa26t
kFNM57K4PGLxrp1JLNFct/9Zz8ofLw0PQZnTl85bdHE3cyYBWDUR9MvdGgUAHFBO
1n/jws4dAQCodxhNIcFGtEynDEVXhB7GyF3s81kiKCcumc3BmL65AiuReMfE3krG
MjKCGjxGp+c2qyulpAufAPWoRuz2SAwFsmysCQV2F6NrjEGJuiuBkhXTbp6mscpW
vjBf6wWdSwsLfdKMacBGuYxcZqcMIJV/NxJvsvkCboEGGD+FRX603eVQ5aepBsTo
snE1TYT818N9+7WSSJLAhASx/rRI7qroP5KVw60Icx1aOGFM39VtLunZTfvJjfDG
D555MTaizfrEkk5wuPmLNXF1e7DD6czbsMAgTkGoPyagt3AjKOdl5dEovXpangag
VFb24AAGE4flYOm4TKBIPN5+tRnqITH/uQ++TJSFAM/MBQF7yOdJ2xXd+bab20pf
I6c4GdIgN8nUSYeP88N8OP7ZeU9jFtCP+CvY1BouNGs6QCIKz53P5w4dcHO6JYWY
jjsmULcOR1QGUNiwdswQljshp25VKo3OoBaZjX3L1mzp7uN52DO05rsub4ysuvhj
JeewY2Cu3XEvbgWHD+go2V8cf/VIp7aqHImLqm4ZGg4D0KI8nXSImfSIpkOWrDRy
vGG4E1Lq3JYEJ00AvIou3lcE/D7Sz9CAPpfW7jHsYp7uLNtTwU+1oz+hSvf8IMhI
6WJu0dGLIlE6T8djZwqFOicmouLd9PJjKza0tRzNd86j9rSHm+swYIVRj03wFyNX
MSDSWZ1yqSMViCrDLtH29kU2bkRCtzJO1XZ6AGObmVm8XyFnYdFgItp+6ecbZHhJ
8dRoUenpUN9XGdQA9v3NvuiCRNc6+aD8Y2y900f8Mnr3SRoDAPpq1VCU5abWwEMc
sjygEF/0TRTuh472e3sNY47C7f62qHkK4ErIJb6w0xOZ39ABPldvQFJYr9nT0Nsy
vLTvRD/gBH6mtb9MYcl4W7yiqjDKCN3+sN1IGLTzAqmS4w06VZNkEmCG83rQcfTW
qaSxQsPMv6Gv/DOVEmhfZ0tRA2DDahmQXnGSRhbr79ICH5x5qaXZjVe1Q3AW0N+V
2s5zmecotqHfqN1srYzs8x1iqcCk6pyHZdeZqIE8QFGFevlLGeYKA8qz2374ZvEo
r98ykgSOnA3CQDFHquM2SsyBHbglx1hbL55RL52y8JLIo8Yw4eXB1dU+VIgiCkjm
CyfEcV3nmJ9uqfLW7csdQOj/04wiFhEfnbigSr4SBJmm7IvKIfd5psO92hkFy6VG
jTfNXgObos33+Cz15PgkvT8hdKbKNXsKMfxk6F+bIoAI6+S5Y/GhL1lfq7XZ+Ozz
g0dB5Lq/tLPs1TDKdC4myzMm2zsS9UmXIVvOmHhVr/GNXmp0kK/J5ETyoEfH8HQo
RM7WpZ5tUOYrpWsB92WTn/qRyVqiONfjLUfM9Gn2S0VMoYCGaWI+DYSwPIDIwPOC
d+R/fOLDZ1XXpXDu3gS8Y9XpvAxb7o1beCyDlusXB58N8J9JKTAfvoDVc4MG+gPR
5cugKHsTDXfDo4/fD6AlmGrAU+5rqzhAcP5kMKr0QUZIiZKzC9XHdFeSTug84EVp
LWx5PS+uIjAsqpVdXXxQp0T1XQ61+NrTotkiSRMi+h/r5L4i5SpUuxUoQAYWQffp
5a5mwEB8TO7OafUcqrE15xyELvSmnwRROnEZjiqFFw6+CYnYc7oRZeOo4KVaVieD
aXFROissQHQBXRfIlDdPahOW5IMF02YlcsgaYdODqAw+tVTYQMJNGefDVW9mWET2
BAvifXj742u2eXW1hjFm72B/dwtI91e+NTjslIQLDXCBJrKbZwpPGv/NEhOYqUP+
uKBavYOuoRhTgd1beHGj3Ay47fwLAwL90qnw3bTCPjnUjoBDzIeb+5JzhNaeZ9Tv
sVeny1M0q7/Sgv0ROBH+9g==
`protect END_PROTECTED
