`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MkOMvYOXORu86vfxol6f63wAVOra60lfdUJNf6nOL8MF0ilXAxsiShW3ozjb/Tu6
zB6cnQvre/89o/nQ7ZCkHeWc0MMmhSHGQDniz6JfM2MmaaBAyGSiaXkIszZaeZFR
gZ+eGtZfrD3tQCqUwA+RWLQJiTA4AXadUmO5eEsHax5C6r/53BifiY/ZPs0TzFi6
pK+facccFvcMFFp/KtAEIEB5U7MnbMoJ5WahBMvhk55ed+GvmFTp5xA1Bw1x8j5+
jzetrTt12w+h9UdsNCAzi8wMq9INcWPS9bxoiyLxjhO+OxklroNqYLp1oKR/oLNt
XO3hkLmo0zkdcwu2DN2g70aQrUAr3fjEU59RZ6TIHTh3d96lzAK5i/91qw01gWh7
U3Qu15j8pH6pMkXiAtHTsCXzZyQGskDq5AsH3r2rWUNJZ0yx2t46LFEhZ25x3ASJ
Vj8SjRZeQOclvczww0CO4Y8G5gFQCAb7LcZwcSKbunddrmyf+Et7dlXgxysoiCot
EGYBMj3L6gON21CVdEVJAqxWmcLOrqpBEmMXN73mF9oCYc8h5vQfGkvqWS6oSnab
5G7BuuyErXMKH9beuUlfStb99ytL5XHcO3bktD6eo4VZU3hsbC0rHgR9dIFZUBJD
33TUNRS7CResceXyolo/SH3d12YlGFeaEiVKgQhF8xecRmWWRyBUeP+NpFoy1wBC
CBmdhm12TRGGgAHkxKchigDZjvB2czLY6j5SKiBbKhiEALh0SjNccrx044d7eQJ4
Tv94oE6hyjF4mjZZTQv5yAs80y84fOGJXIkRd6rjnBuLT2B1k9YgLR8uXcL86adH
e5IxaMcmKGgd51efK8y212Trws3+pFZ584+RTchNcirB20ThAF3l2Z2D0RWvSn+i
phvt0FdA30CPhopHffJgPIXxVWii4n43Y/kElumKLfCj1gXfXPt2INEaNsmWHWA7
jV3zK3OdPSdCFzaKEJxABgr6OeLoKGX+v/U+cWVQg1cPN4ryqRQZ0ipaRmMSnzkq
Ko4OduUjAuTJKGAzUOqxf9iYYyClLNkMwGZoyUtjCNQzJQ2po6USWIR+HcKQ8uoM
+dqlFnRtE7tfh9xAHhj5dFaxvWxHxvWqse+2+8Fcczdb0C+FNiG3aG/leWbn10aw
RzZzl9x2Ia6osQAgqK/qt3QiUfKL+uZeXRoGdaeoMUoYc8B6qFt+WavjTZ36pExT
rUno/Vixt7+345IQYCXEv2GNDdYFYuQhMNKD9PkgkhFeODQ0afuXrqmlLeLAKIvu
3O6Jmia5xsQfke4o/plYz9UuD4sa8+woPc8VwyLJBPSTa2EEhoplYqhoHcPtiQdj
axen8RsjrxkWiC2fDwz+VQXWsjDusE8Dlzba3KFpJnEqwyi+0NSvKTYlqgQTc/hv
fbVqQpTQNA7Xd7P/FWBJn8IOE1UKQ41icee6opO2MitOsuKivFPJzwsYBuO28k40
NOE3cAh/cHDev0RmLGnzbiumWbigl37CrV+nBw6f4rlEFS66wt/Xej8OfRWHWjLm
48KUhiPC1zcjTZbyFl15iHNj+P6htKQ7OZWOf3lFJwFFADpoiaRzL4rvTL+aC8xP
vN2m2WfEbd3xEsQShfIrhO/8QzF4Lp89stEUBm/U6vRMqZJlfdS3KkMsaJypTlRv
VcwmCdcdC7TuKvHyR2x/AhWYZvw+mxcBvqHpQd4YDg6qGFMryq/wsyBNxSRlBVkX
RtoyirwXGwdxNjdJeyBC/ZI9B8tZ+Xjmii6To4Sr0c6tyiLmAZ8YPs8Gg7MygRsR
HRoPqxadi/+8wVOH+/WlZmsxGedTtl/UvxISLf75zxOkUrr+SMjEGH2EU8Ypr5NV
clhgGTILvymTfJ7etGsSwAvToa3lAHF9K/OZ+Cd1mwo/2kSso+b9aK2cIrczGLPR
doMw1KtctQ4wh4uTHRrt+f8Q/wr2Wa/BcyTRBXaUr4hWY6OkbB3n8zIBeF5Y/Uv5
WwBGWEO6liZCkcmYVdkYSXMRawWM92EuCJ7klcMBfXbat0iJR7KZ7xqPuHGu5FZ6
Hs8MjK+sVfydeCj8xpGAU7L+CeJHrZzqcR61TkWxxzYeK6k7NMQENViCSie+o0f4
3tr8H9FnMT3fbDOujHyqOTmVfRiPN6SU5bSiLSkW0y5SPU9qRh2W2dy0p0+k2zvE
pw2PWqZXMQVwbCy4tFrXquxzO6nvTPEMprGY2aVUbsZ7ALWILWye6bD4wZi6UD0g
OhZvmjAphSsQg3mLhNCx2jQvNp2pRk/1avOwoHB38GU5C83elA2uREpiWIL89eNx
IiyH1W03KN9f1fqErerrnXc58L+B9GnkazEybRkfernHHnIE5WmLZD6YqVh2sPTS
9jTGLxS1GaHKaORqLFbbGTzTaeFpN54pdtLTK037u3w+DzzOlvl2TO80ftXIiOPj
ShiEPA9LMaJPcPnHsTPZsJI3oujts7G98o4FUdQGXAsLl42L6JCHrFIUSwiVmGtZ
`protect END_PROTECTED
