`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eaotTB6m7qH3NDC7uSSFZ+LtP98dpI1nvB5V67HpH40PMKltp5oQab92EjNL2eE1
TqCEDbOKTeD/bHjLpM+1NSjryzka6kGdjWdeBcCuFzsf7npNchbi3WK+LNfVtxzX
7+KMeJBLXb4ycVO5snx52aniGrhNOVYWXdaBkEFEPcl5vTOsX5IDgRyonEfQ4hif
5io6u8psUnjp5uQso3a4Yf3P5Mo3gn8hXYMxLtK12WFLOW4bRxRD3MymD2nxzbC+
d5TPJh8+QsRjvFQQVrbqS6Q0yugY4ImhIRi4wVNee7I0C6FdDhMjOt/Egf8y+zlQ
ZYsSznjZkf1X8cJ1ql1cUZjj+m92IYnHMCpY4C7k05O+P6BOmj3a5QzTJBqXelBb
5XEw+9elEvrba4U45cbRmc9MnbY3PAZeSFY8RrsgZbnLA8oN9FVRUVj7yV2N+NOr
HzLboPnrWzXEHNiEAkpCLvUkvCqvtUgW9sOyHDTjyP1BLj81HFJPpWOcLJtifEGt
Uox5nJgE4g/R6/QVgNbUE49aOwneMApqMFnk0PDUg1hQw7lX6Jpep+xK348UKK2f
id1vs8yorODZu5v3FM/xIiUR5oh5Ptx4Dv9oL/tm9VeqJnU/ZOH4uD1uIcUi8XSb
XbRZL6i9nHpSYC6DHIXC0FTmOvXIfOzpvvQm5HXbtd+Nvse4HahzcL0OCphQ9w93
jufvOmG95chnc7oW0RKX63EbV6KIDEDeeMdEWRj9ClHqspecrbG8M5d3SsSBdTkS
SBIcp3k40/awZ+OjAx0MhkPY+hExUXp86BLIU42sD3A3+DjSfWUUBmUh3uhEm4i2
QbSwux8mDvLXUvZeknpPqeEA/WukUu3a3mWSvoMiNw27Y4xZjwwGMT5fltSTqtbf
0h6ioetkYIRezYqlYtqTFYBKvf+Je9p6CqpozKiaMcz4GDHFVapaqYUFWdl+Q+Pi
2f5jO3GiXYifBJbuf6J5bnFdjTHNqb8dkzPg8oYibrhWY2+dmFr8DmsYyQQI4+HC
m5vf/yt+1OgZ5dp6ihEiV6dtCYH0q+ybG+HkHKvo9h3ntCr+R3uxYHfBkh1j4TT6
hjfkBCZiFNeNJwskH5XUCessyzYG6eDoIl1TduUn6jJu68iKRPU9drvZjjmZZjc1
M3NrpkT0ezq8AqB58+CI6HlvREpKpgdrThHqUbPEwCaxg6I9rlKtTBZ2iljvLlTD
59pIQx+s4ITXlBImqG8W0VSBobYFH0ZShfA3Vkgt58vgq0xzk6OQ6qmus52iOsgv
s6YfI3XFUKZPNteV7Cj2yeANVtaCT13WCr58biXZrftQSy1B2qGYo3GmQAOD48jD
H8o9ypYOSimJzPH0EKSDyflzKHZKkgbfKIwToFHcscTMUmfimtDPbN2uAqkSv+el
KDN2vtSCBW6esiKPqB6Rnqk7z+hABzYtqcw3i9BamboWn1ps9ZkBy46h6qDEMS3e
K8HkeK9mgNCJe2EnGqi9bhNnggo2Yqx/Noo9/RjArGwtDTAbMS0vUjp+WNkcikiJ
JWgeMz1CxhtUu8uU7dz0Eo+0HCdMS7zWGP54DlXLIo/355vmFeudbylnI37oll1i
EHS3nJCWRcRZ9tk6QWfkG97KMEg2/Ly67tBNVif96P0+rh2ZnnRAWX9jfRmaheMq
EUoPvvqjg2o9Fd4XeQqy2V5YAxqxadAmfAqH7tJCmn+Vx1WeOzlNOfS/OvZW0UKb
scFFakJweqEbCOPItcVX1Zi8a4XssjBKyoKjfsjOw145iBEwcAS0JsXxVMKZdf2+
owiveDI+W7j++IM9upq2IMXRuvMR1i3MsNvzerwvLC7Vj+Xa8yDUOcRyqbwocxhA
iluIvEbmyL1JdiNdrfPcQvh9LZUHvGgMqM84Wj75fVIMCFmFiLga49vl6sI3wj3I
iiYYodmFUkFbw1TQwF/dI9bVFq+DqZ1huR3dWZJ8FkSfEqJkMCcOGP0924yE+MZl
Fr+MrV8RR7FeWLcr6LWO38CKiejx2Gth0v5kPg8eXZZ/U1q7qLPYKKpR95t9rGbm
pBY6/JYraNefWT4afF2Ba6A8S4w7hLP4Xfu89mvZk1kizPBytV9O84Cp+9LULM0R
1Ri35iTsRPFWxD2GJls+X2GqimyMl9u5RQSJsUCujoA=
`protect END_PROTECTED
