`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6FTB1Mu9R6XQy1ObrXX8eCS2aTZq3k0NfanhuMCeiHnODJVm+XcVO9iZ+zDOkICw
bXp52ld+4udlBEYS1KewTpz9fv1ulQLUTCEYwkkL73h9sDpBlLm/nNyFK18aE+7I
wKpTawQdtwEkK0ENweo8lb8H+5mKmhhC9oxyrjDyDWEbweOE5NUZk6ZSNMUCKORF
L0DNdeZFRq0lbvqH0g4KWVKV4mQEr91x/edtrQer0JEKoKi8rEMETeHmE6JJDLxq
67Mxx5Nu5x8ZOUMKL/IF/3yk+nB4KOr1CFCeuRKCV1K+9mesM4+R79d2GZDomDWn
JoAe+SfQZALcKfZ87HegHxiVBPSfXrARkjfuKAIPVX8MfSnQDSM62Kil6QTM+U8u
mNLVlnRCArK3tkuSP49FQuFU/CIEJffQaI4JjsaJOlRfQLqTbBvqE/2e7tkL09E0
StUCDr5FmxByw9wBFoju3NK6WdImayRmtzYkXs/MKLJCw84nhupfiW9HyVm0b8cH
cS8FPUD37zBFYnJRjwu+Ryrd6PeLwD1ISXeUbRfG4fAKk+Hk9j2liFmM2HBWf7am
YJrHHTfKM5/9gzGve/1/tzlhzmgBZ/qJzBGpUeIfO69iE7kF4kUbWURY/vXK68IS
3qt5NJsyoaUpbbtuKqqyZS6ddOg6a61AtbgQouoyEi14cb3y1w/Y0cxfPEvYIv1K
dKIv5KjOsIvQgxhLpIVP8lGEWAO2WbgWueFAe6uEc7r0qIafmOLHLF0/w0EDT45H
FJoY5pBgi+3Ey6cP23OTMpJa8O45XOI3HP8NnySYRt5vv5Bhg6JbMJb6U011l34i
/E17oaB2w38z1l2Y54xMh6IVH8OUo/OOdbObxZueMsKLZ+xQeMZKDbPDBDWBsRtH
zpCS/DMU/lFHpg3ab7BIfZy72cc9mY3t9O/ygl/mP7lAHWvknCaSyOL93mnHxPRw
xVYSYHiYUAKy3KMhTmofE28hzM2eDTbTY2WPJtba65e1wss/UIkh4JX8Kq/EcZVC
LepO6gPJ1XQOh7pquP2+cGdgYxRZ7apgInTQvY+tz/1YpyOAqG5NwtzxNTYbyb02
wxY2MivfjFC+Fk9eQ59mxk6UEcw2JM5KJD0ERtCWYlj4vgbtVuPvy/Qwb1HFjUiT
ggZtItyIePN4MwxMRoAoZbvUP4Ls4xQxCjj3KB1xCTlYKHZFhYDRba0flKzLhQQO
uohmEyG3AC6tVjWnL3aXm8TXNASThWw2vOAwBTKkf4l2vcMAKtA2nX7Kl38+ff9a
W1ogQtUOvBWkDGYm+jDq11GtuFtIeKr7yzryfnCo1x4wVK2BdTHU9yLDOrNcn0mn
tKu1Guu7iGUW8XDTyH6LPjNrqhzC3Brbtv5vK+mjFdEaDgYKvjA5kfc3uwWNVQNc
fIc51EYwPsJ3kpg0vKfqArzqrRSj4H9BodGZcpcErkOhf9pqMxS9LLBQzhnLKwT/
`protect END_PROTECTED
