`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QaP+Z9bBjn3KoLE0nWBwGG5WMzsxPXyeMHMfKiX57bSpgdNyVnZPpq+NNfz5jPru
/J2oPaKSxF6uCjsRpnPPDg10DjmmumIQvUjIFMygJgt/EHQEh4S1glph0OQmRL7H
by8PXRozJmr9jO1JMREVtaP678u9n7ogbvE00x4tfGQi189uZQ+oTXXsHUYRXhTN
eVDEVHiz3tA9eF35h0CPJEiGqLvjBHjuJ9oSnpOdFw1K0bdR+sgc9YF6z5E6kL/0
LOZWUAoFeMvonClAbYpjGn73XzVw9jneuKUrs2PcnCsmjAeLIVmpbPXXoOt4L00D
68FB0wP46YQy9kadTq+WIPxHepvTTNigEEzZSl5sNyiJ1gKARcw6qRIUPuSKxUcB
`protect END_PROTECTED
