`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TcLFgRsS07RrXqC7QVN4RzXtJTSleCOZQTVSyFbYGCQnO79bjQIFdU3V5BuW1Vbb
922IK1IYehWF7T2gwSe/4W9Zc554OzPfxbIQP+aZ+NUvTOSaq8rebl1oi7qLa1yG
cx+eIXT+8wUJZLHwk1wEVP/LHbZutIdAuVwrXzDSaXBwqoG5gYrfebCAwYnOL0Fa
292EIzF5QOZ2ne9WCxSvIv9oEaxZgWkjBfMfKeiyy7Pl3R/dmy3HvREuqdx0L4on
A/HROi4/w/RKjhemVMiWAoJFrMbehsK0omeB1QAfgejRD6G67hmzsowUG9uM4tcG
5NI+47InKepak316yZiNZzBR/flY501nYABH4f0r6chYccNEArzbndZ0+OQpbCdt
oXgbjRahFEg4KCq3FYMW4WbIKA+uerVlzy80TfqBWEnByOugBtVC5p+gV8hsn1rG
eKdSUS/obYxhEVX7pbjcldUbHt7w6grovnb2LK9KoxdPquw2AMX7ANFNMfzsv8Mz
Oht4TjUZcmy4bcCFZbqNw7CChoWD/9iaElqzv4DWBw4oI3uHz4nXX7xPx5N425bw
TmDb3194WQUw6kY7r8VBTDVEAvADg8UnQgTstNMtnwYLZyWJclCwiC0KCSqQC2sR
UeTH2a2dko5sezHpN8u1muWYwunF4udOklHJ2Kj/4hrS0Oj9VDU0tOBTe9ghu7Ci
3BP8K2Q5dwMGBF7pjXXho5Fc9+z+jVAsZi7M59NEbPB6jUhpvE9hTTzlg+8ADCNV
9BMbhl5y1wihLQLIv49o6yuQnKcrLD0etERq5uQp2fUlOyV/Lb5pykNtkoPh2W6C
pXqzvlDc5B0ftRsY9OQDll7WRtB5D0qgRiMl3jARKxX2puUN77w7KLcscWLpJt2t
9enAK/V1Nj9WNwmg9fiNluK2QyLVUZqEzkzX305AFLsvrvjn/fGm9a6llH7Vs6oi
HloRaKP3WJQLQ+qMjQK1Gr4CM6FOcCBjbTKvy1KgB453zlzDBa4lCXjvx8xt+ptB
9Ix0WVqTvChefbdUyAC6VSsV8mHWxvUFsWuQszCi3EtWcyfQBcPcjsEgm+IRlDls
byg30PFqsop9Fdy4x7kBWVvBMS+N/IAlIaHgJDePQ87Lo4nPfvyCJkG+uuv6qw76
16k4jzNv6ri59qfj7rrv7W1sn44ZAuCLk+4mXleOJsTORGoTwjeBsC3V06Ypj+16
mbGlers4/DvXHbLSSGLx2JcAc1I4Fb0pVMqLXrhuTgjGLoHp7vIiEpXye3DvjRWV
4RRtZrX/EGC8bz8wvQEub1nnZ0vYVHT/b3LHAIKRfgdcOSfJkF+6f+/2pgblkbTf
XW5HN4R3dzFQY844Ho+csejuuXrbH4Ei9zSTfKyo2FdF7uhCLpNd70byRHo64jXS
YIlWzcKo4/wFJfS8XlnmRC0l7on6mT9xv3YqkKu2sjVnCyBNTIgq3BTeFiaHP2MW
`protect END_PROTECTED
