`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gz7GNrJdLaTXvYDp+NYzNpAZaP/UwQ3Ej4+MsaBZlZXHlbzucpyqxvQ8abNjUKS8
KVSNb9UnebBzmf8XSlmRbd0co5JnPBCSaydI0qAAtkrUWvNM82/K3ZBorP1AsBVP
68n4RHTcftHMTlyUw1x45hD2TQizml3sWTREvJBBWfC7cd1RuDOMirabudTz83fu
9nG7J2/kATrMGNE2sX6n5JOxO3Q3VGPOmC8w3hvN82hk3Z5LV18Qre2J4eyXuMGX
pjzsEQBpOda7tXp4v+ZtQZW6zKzcbBFs6LTAEA2yuf6RJFaLm4UZzuehg5j7hn/0
YAgxJnfELOwIamlC/wH1hiNE6qquaNsiimUsvv0TEYcb0NBlR/8Y3uOTrc0TwHys
rI/YCEIfTVCkeTVVn8UODxuBJ8vSpKI78Bm7aT7TAJDyiCqeF5ccIVBoKS1CXEX+
QTc4J1uHs25UPwqqVlUtADi7zV/YTwZ/ju8TBzeXMuSqoF9EFhSdiwElz7euIdjE
IToMuVL2pjyLG57ddvF72kotb3guzobGFJ4HSWAJfzRGv6YETy6BE9lMOWrYdOqQ
2QboZRVpF549d5UoHsF/CvMKnxZHUD//hvaditl7dLPKY6YjHcbOsisgekLzWFr3
1pjBqzk0YYnGT3/tPdDyaq/A1pRheQFRff8jp3hG0mLNvzEa8y3qqm6O+hugQP7T
NBHJY38xg9ctnpae1fPK4nQqvB71adjMCWUimeiaxyf/qVoJ43Ddaf57/3ariE4w
N7d6ISvwAMBda1kEcayW4eGLVnDBVbzy/mdkDyAA+J0hsl1r+4XCmSieUfVC1Uul
ChknSQ2FruCLwUOAVWHU0sP3LdNzNRUHvF+H+1smFQsYlpqpPbHqPJCPt+qbIaR9
6a3jU2BtMsVwM8/fdcbTYzMR3GmB6pqS6e9tI3v5BkGuuXwBw4TWPfEoedDq8Tb5
u6TwLbzDqmzJJ0lsqs2r/Y+mcPsmPiXkaluj6649gqYnhkM38+x38yjuw0b5shIR
i6BSIoFr4xoDoavTdkByP0u5TKu8qdG/SOwDQcCUiWexT97fwkcGqRvA00RKPuCw
XSUygf6IA0MarriMSLekXqzeOT3YyaHzJ5EcVPSyePd7AbkiqUHtlyBlYZHVn22+
ivZK6acas7lwqVoewlGgUex4GXsK4kodaM1Sh2U/eTKXbsACeSxvHditNA+ZzAuD
Lt7chQJC5vagZuMUdsxoslqw5ffs/gXV59XywJcPBhLTZNr6Jht5v1X91sD0wYQZ
bzdltukZ9kfB69opbljmWX6tJts16Hm0nrigEoU+LATg9LORP5diK8ikndEU7QMW
zWhafSh97ajec9ygOqEcgDXoVVGt+02viTy0LeYqBmilMOVXFoiFCxNbWFpTOfYA
aiPRq2xzlzpakzVV2EmL6pjACituqeY+GRsT8ly0htCRYDmWSc9pDaet39FY/uLO
4U+v2LhoSFHeJLwF89ibZy9brzDW9hJRyI5LS77MO2C2ZHiiMeko2mWU3OeEl1z+
MdeHCYwGbHaKQrU0UpozGON/wxStnLBA8b7zL7nNW3uQT1u1EOJ2rxOStLzyTl0K
fA/8PkkZTjF6TmlSWl1dXAJoiVE9Ztkwtno/NiuwCMNNvsu8l7c9SGA4StQVwlcs
/sjVw/uWhl6dxUVUd5HCrrRxzchsGoo+Xf6QPpqJCDsXTet7M6HkbxqRLR8ceWTb
L3yjTpLPGIbHfGTuA/Q5CuQHpt1yeYv78C2iQNtkqYfi/s+dNH/C1GDIkB9PGD+t
EJncTkvqcEIcQ47ZZdRqU4rIf/GV9uxvA8QausgQQGhSvbpHpz6kW9vZqUSz+hxi
OnkOQZO/HRM7t+KRIoy3kWBb7TB34WpbtUSTQVzW5KTszBbyKTNExV8+EvJHmgy6
BO6BfdsVR4fxVRpWKl/0D3/8PGa6We6ImK3ZZZiWgVW7M51/frrb/JBd+eeoGd0H
5DYjhiWtlzg4unVAnCvevz2hyZREcQAUMKHXkX+ZQtvBh3NIdX6SfTDBA3ybDgr3
B7hXe5UiOhZYeRSTV6ps5HtnL1NIAtmX467YUU8xiSxkowQ3f/xyVd29dCyvXzvi
YdxD5Xy8/bxMFI2yvGbgPyqTo/eAQa4mPkzqripLLrGdeFqhzRfpMJNVKbGsCZ6U
DviqH5ctEhj99HAcBfpaa85s00+4MeZDiVLS5dcmn/wA3OHibGtHmrL5DsrScIbr
kO3nGQFOW+UXmIIZKVQm4CJM3zu2FDomcqS23S6cZjCVphA0NoXDthrNUJn+Vfmo
AOfzytbAK6ORcRiHMwMxvTRPVKmbIhBzxWyn1F1T33MNNb1LZBB7jFVISXzbRzUk
TikZaMpDmKAQ4kxLCn9Ag8K7Fj3hqrMriJBW7hCksWaxPDrLg+bgEuA2MjQcIB8w
EEKp/ruJLbDhryEuB3iQVCrpm+vlXVkagoyPJAD0pMlyFHqNsx6JA7SnlgPF1R+s
7fY7cB11QVJqhXj9Z+SqY5XstkcCSCbESj5t45U4uMYhARpeWc1AI9V9z96rnVfp
t8+MRTs0UU9ATSF4fGrvASSjsqJPERxRYi5mKbDSg09RwBg4kZWG6beTG4dpTie4
YmD4sXJ19cdbBOK0Djxn1ETCI1i93Do+0eun9+JmE2/rqgZlrfowWo9J+QGDYz1B
nBmpTR270BiynFm+Y9dyGlNIOAEomiwbWzVJv3KvytRfMzuXuV9alfvC3Rn589AX
E2fdOY04xVRuBSk9La2p8d7GeZ80AmGMuH8iDVzRG3KlSFo5mmxjmjTzY+vjzg4H
UsTer9iv/ZXD1lP1ByrkzqLqMWF4bKs1wF/yXaUPDpuSo75uVnHylowrWRzW6Ewz
yqtBITkh8PCmSn9LlcV96i3pVSwpUES58CnHK4gCEA4twQRnX3ogjo2XIz5VtDlQ
MT7xnmoNk+p4qVchPeAPFUZEHItnJmdaVCf/YJkeOCl+XAK63a0jNOHT/hz7e3l5
hz+ML4/NTzskdlZpQWVoEk88ojZBEgxlQLnLptq0YdbZyov3jOZVq6Nc1mnRt5RX
lWLL/SXcAOIV1clnYhrdvWSj3osedL6l8jfXe2zVifA4WXC/Qf3UjsWtKUXwTPMo
IsICpVLcdommiBZ8w/KnBkVXi7fZipHH2y36QuLYq2/fcc+L7r8yimOb3P3GSdTx
velt6VT/hRkEVh2zcsW2wSvYiiMBsOL87nHso6DGnOyniA8gHoxcfKr2J/ncnTtZ
oZhQWZTXcEF34x2Eap2W8fLYDqNaaa1YSRlMcePYbU9fL1AWZqqNnkMzo90bggUU
8XJeZQESwEoLVQoCNFldt66SaYPzsDMAz8PO348pcPvWqmZpv+RpSYdHN0Fqd2kT
UlnSu+cXIP4K5SkJwKj5zQffD32v+i2ASZQ+PK83ZpvbnkuyL3MERodzzBu832pZ
L29RIy3To8YsxFnY3D3jD7EWiUOvQi0yMGzs8yr5pAlco1Ni7VV9uz9z4kjKb/4u
tb3lrEW5AaFLjeE5A2cvcZMQrvJNvNt7E6wtzBFTRqoeO+CrQn4Af2u2wwwMhSaq
IyA6+jUKC6J3kewj6pWeSuQN53Rn5FOcSCcaxYc16Oh6QkfSrQMr2hzt/QpC+QSw
CFb9V/m6tta/YxFG+CTtQu/2LxQxsxBWkgLToZWVhBU8THhDjjA6f9pZrlnjBzkI
8PyCOGTeB0epbVlrXat3AZ0q3FbCcXOVo2fmxpD8KilbZUa6YqSLgzAmgRfKquC9
BXxm98HyZSIXBE/Yn6F0pjDTF+c056Vocz1JgBq51WFD4pKhFpKNOFZDFbRA4Oig
v/YiPlSJkNTa0VdS0k0LN6+83viXLv4Tv++DiMq9fF0Nf2pysZZYe/6u52T6jIXg
PgyHJbSJqx5zGJh2ETKuGeIwzo/V4ZfF050zH9HfdZRNDrxvKAMQ/ZV50RHyV7LU
GY5m4Y3dDcAH0c/K6OqBXWlV4Nnozluivv5w2mk3Z89AYyHjn6bTCikmlxBQnJeJ
ZlQFr9yUXzBmC+QZ7Vf9H2wBiDTbavhhrkRTg3loPRuik2SCrhURrEHNjfT/iXCb
DYcVUIpqT3v01dGMRw3ByesXvyGHKXBYWrkmScgEjvqpgInBIi6LHc1wC7AgZSjc
/Obx6t08aouLBK58VRD0sp0A/iiIOhgoX4ohD8ENDKF8w+ghGo5HsYblIL0+ajyR
VZmPAS+43J/XP7svhP4pc2wa2ELqkwqWpyO95GRhnnamBAx4sVlX53ZnQS6rs5Lk
y20Djaz46rxR0RwNDNEZVGiPv0b7pTMr+bFnG4lg6B1FnMInnBPsOdqbSQTgGHyd
jkzRemoEPBMxlcdAExAJmKLvfkfYVyjUSfNJqdJf7ojgDM6BePeRmawHx8FFx/05
V6sdbPxYqd21zkoa8As35UOi/xnQwy1Lw870eiClpVr9RGpeNv2HkBBVXmiEI3im
V6TChmXuYENxnVoQqIW8Q2gnVvCg+4zjt6fPqFJgbnFuOFeMqsot+rJNB/4nktVG
rgLvaZHChNPnsuH8d4E31sX8Ri3oIf+7utU94Kiq5lXXxD9kO6w3/GWpZMb/Wtm/
gckSqymnDl2UseHs5Z3/vGxNGm9PEcnI9Bkggfbc/+wfbPCuQHHenmG3VRa1p/Fu
SR3KB/xCsB6kFD1+a4zeIsRXRueAaGb1wlG1NvHFCZ8crIw4lWhVyT7P4y5V6fR8
JqPYk/s+Jzada8z1AWuMJN+aenpXfiFdtokQpCu1MWFZ/XoQOvx9bC1HFjXJu/m9
95XcqgAx0a1JhIUY739gMzE7rg53HagzbbhVGSF33IJ3q7QJAFicSryZKqAPlEb9
1rIrR8r5bA4piTbAb6X6baT5QFxsFp3F8h1MxAMqJgY2UKPV0/QlP2kOYrTQUA4K
Ob6JCILWqwYft8aCxSrtrqO3efDrEHOAPnTmtjOJTAoGEqC/nJP8+QJAawzz4fyg
IlNFhSZUL7vjFgaFEdjSx5Y+pKXU+CrTMYl/hsvDr2witqSYuJhvFo8G5IxSIsAE
Y6THjcmlywt4ajMtKvOWed47gOopPXLDFFJXESwgD446NkiGGdVzAlxgrFdvMJ+M
KLUUlvRCyg1SpIjdJnI0PBvyWRQh5owEQhdg9tlAgYfrP8n0LZJVe9Cm+0K4rTzO
Al0SCPbuI9JUl/88WlOYrqOGPB21pNZqfBQSBPEzN08Q+o6KGEFi9sJCFzJeaJFZ
AoYYVlix+Xf+cb2EIGLzVhQc1WV/I5EYj8ivyGwSmaM3vrYgg6wiK5pYD4/b5AtJ
XxN3Uzu7tcvxpZikHWmPxEbeAcIk4eL11ZaDdLGQ+/VlRliiOW+T0j/WqeiGe8Us
GPVDyfnBqYbzpd1sgfvnF7udwobI2MMyJR5x5ibM9+PMdhL0SfLR+18ib7XyiJOG
eSP+e9deKM8J4VQt1jkgnkqhUEGKPuwjw/Wu1K8NVFnPHGzV22z7ObK0zhy42hPC
2XjgrOlvyNshZ3BzU3PAAQgIkvyprIjVfqYjYNpQOIP0IoMpDS56T0mMlSEx5BDg
D5bMn9LecXiTW/gB5WhC4nTH9vH7YAzRWyFTBAh4r44nHsL0fSYqOctgqmOmsHKE
RIlDA9q3taD0XrFU77c29zxN2eY4g5KCmkao8EmL2Suek2krtG5yeD0y1d1svWJ9
RXfGRmtCIiLCLYQ+Kbvfq98M5HLhp2AVsUSqhOPIKtPetBs6MEZjiSJg2W07GOcY
VKYK0qIh2wLF88IwMGdsPb6L22Qhm/qlVfodlRQmvsr4KWnSY0yXM0o5cNTYB5oL
VFNCxRwEyo0mFSm6nP5IPeXNOXCX0qe/lxYDzZXAyF8olwZCRYtFtcCVpNpnqWEb
jez9d08kmkwN8h5xpEDkhUMxjZVFZOqRjOpEX+/ut+H1ljvTYVeyz5+dWUoXJth3
U4FrGAPMpQ7+dfrJea3mMn+pSkvO+o8SZoZ8HPi9QFccGjnGNORokAlT6jAeH3xd
WQAxGb8X9esXayHjCjo/2bpPgopxIP9xbhinu87CdVc7ZJyTgCjsMEY/s99vXKzM
TRfhcrSjA6rl1C8Bul01I1yGoyg+7/mN3OOFtwVxdfbGuh8LDXjK4lQPzPvrDgKy
VXlRQDlGrhVprs1cI60HucAz89LXnkMYrj6Iv5VNzJ+mRyVPZsG3UsyDkxpx7YM8
JeL1kPzQ5B8SI2zx9Bm46XtHxLtgB8D32IQX7ZXNELgmWuZD9Tkq1bOp7nc6FhKR
gtl4uopXb+cgbAvvHi1Ou3IhWYDfZjkrrpcBEDVk+Gf9i0N/EpjTawzukenArGJN
DMP4pwHGolNfKImJzfgmiNzIxTZZFuGWKG6fWyzmpD1zRG8lpgn+FVQ+YEEfweSL
A99ehYGNYyabb/2srwgy+ha7Lkk3ijVaGHxzpWVrrdsY/iVYMvp/NizWaY1Hv0c1
YqEpL3qcSMtotUEd8iOUsK3a5eal5KgRnNnevmoHcBbTzfj7LTThQYR2gfvRCK2J
rjIvGkbCdE3hNhYwiIRrNHzIRcgqGFu4XidBXc0gU0a9sfZfSXoUd8WTRgX3XkkD
yYbukzJABcpOY3YfOJtLup5wbjq5byfMF9eFMzEAN1Grl2H+Hmli1+9/HnStaVAi
xBh4z0Bj3Ov8+rtob3eU7yP8ljgQSODC61sWqJKagrptiRVWJ/4z6S5TmSC+gu7B
jyPgOt7HZ9kOd8Ts8AwNXr8sAgZP8VcdQnx+CyQcGKE4Jv3wE8EshW8pO8N7BhYp
SsqZ8Fm9UqPC553dthf/GTEXeRfCly4JU7ERa+AtGVTrmW8DZUHabJ3k9uGQEeV0
Hir5x3o5MVB9l05yff42LQAKKclpQpqWIt8DFbbUaF/xZMCvOVJ3Ah6C4jmFV3Xf
7POnP/KRGoIzAU1Sbx844QgSRfAZUmjhSCH8BcL4N95m37oD1D/j99CtHXQ9VP6N
bNtsgrGKG/jcqW2tes9WxxxgVujpyjUczpOzD/ViGrURD0x3R/1beKzeh+XSMDUg
tQLy0s1psFlkm/wRe+OYII/Et3/Leiavtu4MrBLTVSuQWSIz6+bT613u3bgVJCx5
e7TXevJqdcBDenjb2zVOW4+6SVbTnpNTZikqKUNGf2iEwFjBulMAE6ClKzetUrzA
5ry1czoCvOedGbCV3ozbqbO76kTfmK9JsX0WP9zjD1SisRscAIVNR/kJUY+Eme3A
jYisV+nkYaf3H7YrfdNQIM3pN5ALaqE/jlT0TIWylZ3kG42jRfJvPZU+HId3h+he
6A+pKFaplEUxKyoh96PhaISFBjHESY1YIrt+fBust7xiMFWF6flIo5P8I5cB5sUr
xUM44vV+SDVd4FyhXch0Vm+J4b6//97JBtzgZx5Dxmb/NRSqyF/vza3EJb+m53v1
Le4N+f9/5x/5+wEAEg4Zb8/E7AZjxSK5ucDn1bfxGjyKIeLPtJXMz5UJ9p35gVO+
IrbuTyNA1u1dOFCrSiAhUrMEx4MARmZDoeK9pl8RSH1+2m1Pp0k9X++ARzyK0jFb
hQoMtf6ePsnLu1SVQaFoPAOFPufGtW5Q6v9pJukBKzhh67aotCcaGm+wtDMsEd3i
WtE8KD9UyFj0tcjze2PI9R9V3NSIeDv7BGQEoKHmdZtXK08CZuEjNHvvX0cVOEm1
BFnG7gmZa/cHVtbBfQXE8EHDS5ktX4NUPBBWxm0Ph1Pke6yZyGQbpJHtNebEbcgO
fMh8ZzCl1sTtfXjOdlB7t6ltsOC8mWfPVvhaUt9ZNEfHG5C3CzyKqQtJOVVcblX5
Z8SIP1YRSMMKJvpNZyAKdSpHpf6JE66IF2bRSse5+mlmmEwNMdn09pfZ3zy2z5Oc
T99h3sQ9skmtpCmY3L6Qqrm0AjHLVmokUd0MtqteGUs2PFBOj7DSzFvACroqY1IA
EW01XFgTGAs9N9LYM74LUKPe6A/Hl3OLYLei0DfkmB+zA/LfEflaPHNX9hgPh6fV
tWnXtXb2DXT1K0Zt7RlYtZmcEpRbOAG25fUFcdAeQvfZOr66dzqY40zpTtxyaPy5
gJxMSKYWm2gBbN7VnoFN4y4ed5F6vvbEavpaFQxIL9UBksnTAG7Ne3S8zRmsW5eX
LeTYs2v8pEG0mDKwYMfw8EBgihlzXwXfa8t2LqO7N+U1wpa60hpgEc1OtVZ/csTN
5tbrtZtPTUYBz+ae7rUgpp/wK06wvfJ88dtXNTEO/JIj1h7sKuHjJkCLhoCH/5qt
Daq5OiVFCD7Lm0otKy1l5x5mjOLGxf/Sq4/+1UANfI7+hpLQ8ZqOckTXd0ZYqfmg
MqgQzP29dRafSUbmV1UQwcJvK+uvBdmxKkJa1k8t7Hk/ocGsh+2zXWo7eCNjvlJT
ZUDJrmAbkCusTtkUMyehXEMm+Bz4pYtK9bxGuOaNJWpv82lLtA5E+5wXlUZ9YSrR
LRqCEJQjLnfd71icJOjXjpRe56oRpjAQF0NNkhN4v6E52wQZBzMqTbVBO92vZD2x
Rgb3um0fV2uL0KxNfZpr1FCYfTjGakjij3OqKM+Z4r/IVW8AqilMaS2SoUgKGnqW
p/AFAdpbVNOJ3kPOnaUVexwNFyXtvtFeGRwMKFdzNjsWXuXBz+z/C7t8k8y1RBS4
bNl/xKey0VYXJk4/00Sy6W6QkBkQsqzH0ASWTgZegYZI3i+MIXp5PXQcGi2oVeA1
nxILRxlEw4XyTkkNADvoAmCJxvy+wqsu0CKfiIHCOynHFxZ259Cn+r5mIDbmrWey
/2kvTjgRXUG+Ix/gy6lZGhgI70pOc0MJgS7qQ8vQEnbFXjrKzTfoHd4+DwyqsToZ
p2CCCqsVfr/iTD07TFDqgj/5PyttO58fIRUjqZ74JVJX+6lQctv9sZQjB3lGCVJu
dWnvTU7gV64mOafQ542kiz3ik1k1nIZKP0ircQOue+0xhmm757D2l850Mt3oTX2d
IgdcLLe93WYFu1el0kRQg83R2wF6wcCYdc3oa8S7JRZYA8CYEpLj/H+5bljBWdcz
ts9mr0Hb+4zrX7Hm0eKO2C5QkHoFxbWy9UvnwzabjId6cWF/+O8qLbBRf0/6ZIKA
vVu0pnOm7AyAWfQmRUMgRz21ySv0c8sHcX/LRwiFWnALzOBBQEWA+TfPI1BLHn+1
/xHFBd3jVaCgeRh+yNhp/VwxwGQhfy3YtgqoO18zOVoFmYnpiaYiWJm543DoJDp1
7KUCCAH553IZNrBC4gePyvyy4r2iTrCBGhFY4DT7fiRvIvaMr0JDTmXRKxX3gjCw
jEPR2BwGcoAL+IrQt5If7j71Pw/nqwfCh6hj8hVJEc3YIUiOvZv/3IWKlCCoKHTV
lPpxG22eQG2sIqTJH30jXUy/XQyw2scocLJY+i6xM3mzifTNu/3nmT65VwKsHW2z
jdCDZFbcRtD2s/89gK6mpEDqma9wB0JN34aCxAYuXvzNjVmqF3eNnFjsjeG2p5EL
MtI51s6pauEG+/F5eMrLbzV9Sl+k/ytAGWvk9yHQtuAV4RbvLLkBAcd1WVqtGqJE
4X7cHBX+Vb1J+CGzKx7KOh5TR5SFvZd/R1BfRikxfNQsY6nKffd1GevCRL2VEyPo
b9rJxee95fXMgOgbIS0GHqvXOWyTZT6c5krCJVSdd/1ShpluFlgEh5RZMJl7pOBJ
`protect END_PROTECTED
