`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Z/tihXBriE2m0nSCWthKWc+9WzSQ0TWAsxPDi0ZN1m2+cJ7MVrbF1VpWzb7Wyqc
Qx1KkKLXP1RO+8r3I3rKcp4OVz4GJ95XUt2U/nu2CvNk6bSTo+jNoPdNRuwwxzye
mamuZCqaz/VL1X186wBJWHNEWjUIJfxi0ECqA24U/U1vUppv/x1hl2npbuYSX06t
19dCVDVcL8wDSEZORrbPM7vFAIB2QWWlhyOfFEyX/aG0Rf8irjwvpTCoFq8YLuah
dUkOPFIcN7+d5Z+eqdrN1HqtKyVGY8L/nJx0Ufd0fiPTTZTgZXAlGbsAr90H4C8d
bLBXEnUWueXoIDxdterGi3KCvl7V0g4/0KI6L8vbCEYSHI9pRD8oxfXkM3qF0MwT
mqE0/SAYx7grExoc2A73ayPgEoJnNGWRSNXVxjZimw+X1SvmRgTZV+OqCVSNvVZR
zsvDCiHCkq9l8MS891+3eiP/2uhE+LGWpjX3TgVs+SMMPV73tilRGwA6lDTy04yP
vF7O9hQHthnUqadpE2/e6h0CxIuGwszOrhY5wb//3Hk4Sq0jjm0g5RXErD3uVIVk
dCYdVFtrAs6CRuG2ul3o6vxawztoRMRSZxoAk80YDvlAuZG8Ru70FigGCR73AHU3
96oGWeNzcgDHscFVPC8xmLttIPwBoAafShDKkOTL8Zd6Xb+cPLNrFtirD4kKmkhh
kPGxMPTWy7ofI4ZLwyIp/3NsRqdDb87IOuA2ekYkZ5fSnzpROdxXQmJxzbJRWKmV
SIyyIdf5WYiGPb7Vfu4A7/QFg9FHUIdJ3BWNVkRPARxo6BLuxzPPJ/nlWDlafl8i
4i4avpBA9NXHD6DCmM4Di1CamZZ2ECaGw0cFvDQN7XqFLsdgJhq3+YOPFOpfJhhH
9Eih8J9VcYuhwU8rwuFiGD6ccHRoLf6pmGI3NtYwagUnwemORFQeHkkMJbsNQ71K
uS5ZOaMYCMXj2LP3Pc8aGK81aQPNpSgQgN0gl+V4boqmED3NxHwfRCHc5GPSqeZR
xYZnJGpgWEjrePQIq0CyaCz6vJpW8ZiUPCReMpFuiqywMTBznCYf6jWcVol33qa2
7vSSrCmg9yp6SEPUQP71WKe7kFfCbzPU8Ng7QCi663mjNzcUadAaGhYYGmCxdJEW
CCkBrlkc+BPjE19e+BVc6rSCZmI3BUdt7+RlZlqqdOG7rh+TywZ7b8PTFNZzXRAO
dQnVQYHjpAHOSTT1V4aOlwjzdcWxW0UPCwKqY0bfW9wOL4UPOF9xE5MhZHUwtKpf
tChrYQ4n58f3C/T+sPguiGeCGzQ/fG9NdJvYI0J8bhM5Ila/P3EX3bteq1pzE2Zg
`protect END_PROTECTED
