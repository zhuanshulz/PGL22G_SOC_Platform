`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JoJhECz5nT2lx8Ir70ZMWijBtZBXDsmo9VsYZdl+Hdadh/dP5cGlw90c7DdVgj+J
XVDNAKnHHsYO8A6/+d2GgKc63TBSHAnTSWsyRsoigkZmrHPw0iWqSQa6E+exLq3c
ZmqzQ1I6TxWJRSNU3NBV4z5sfKBHLOAFAo8nRQD6zq3U3cHjFD0FYLosKw1P3n4M
ly1nGRmqWxeZJJpkY9Wcw3EGkd1NmoV3r8Qzj5u7YtBh3gIWF2TTTA00xCfsKMlR
aym+JjeXBKDy2aEWf355flCBkHgyKiR53Je/CxkGTZvAHfsBNQZ0+HT26ABXevfF
1uiH6VcVDyx5qL2Dyow6ySpHKuate5xk+TpV/YLL2GKul+SgzvpEzPsJhGTJl+eP
eyBDfaWZLVEXaR4jqKlKjuGe34bRZRTf8Yp5a2Dh5Q60QZ53sHSF9RZyiulRXb8f
cq8rpmZboLpXJzPANrtn2CkjjkwiYERITqrsv2rM8MVze+Q8Pa+tdq9oqrnU9eYa
itEkPc42eSS5ApF2LAj7m7wANxVhl3FbvZxwFuZ1QVkCcRcd9tPD3gQLvuwk6kvv
0d6PghXMYqT1TcleA8H57PuH1XOZrl1ntCZkTtZ4xRrsangUcQ4/2SX8fET+bFZJ
tvyDzdLGdmK20FL3iiG4lNcPAsyaGp6zDBr7wUAkBG+hm2m7cKiJeCTDbGvS6Vzc
gWJB2ZpgLQt/6X2V9c6FJQPhVW0tUQyMNxq7i+aKBHCd9Zyc41OYx3FY0+NrPHMT
8NggYktKDUCVUKhUagKeUvFG6H+AZaoPbNfSYllvk/S1j+v2Ay12ad2MLUm8gaGY
Wst+hehDPwSp7K/2Pt9LVQgdZSa1N1gGiCL3H12JpZVut/6XUu8DjezghugNCoxM
U3yIiPEynygab7Cldj6xYE3ociA/Gul6yQNKW/+BRSHEg4vH8EfCgeLoZu0N2tDV
7/apM+EIgj0HC+xBzOuD/e0od71/3siQ6RDs67aZE2f62PEMPLP5F3kZ7JgwUfsN
BLGb1c3P12AR9YQuJ8eQHSMWNOOcweRR/sZc7tT00SCD6O1wLq8+VEdsnjei/Bxa
3PuAU9BTtl5MCIMjv2koCvKnJo8SejC9hPl8bf+Qq0BHOQQbV6np4UwSntpSsqwJ
IsWtg1MP78zsOHYcxrCO4iSz4EvmIf9hPrLChehFCU8C6Z02hazLEMp7oJN9JYRT
RVL8tylk3NIqctDWUWVjJWyhpPjtoC66g79YZ0bUvkSSpqxn6DLkd3Dz90Hjs3wb
LUwH8xwQ+swODiI4XOGVgqAbVr+a2jzDgpdVlra0t5mnFe84nyMubFB7zWJbpqFI
hpBvM3GYXYfKyineyG24FHPtaqPaGn6wwXc/jXBDfbuEebAUxh0p2kdiUkKB95/2
eGOmbsabR5+IYgYsPZo9Vb/Jl6YMpHbQGy3LjX16CTiucWN1Zjkbn3Bs46Pjzq2J
R506KKEUD2GSRfZ4LhLXt9k/ZnPwhmLB0kzaFPJrSe7gTt9/pPc11yQnQu6IQSw8
Luj0rvmgR+I9QIi3fUYVB9SPpsTpY5G0tx6/flbfcQ6Bd7O4Eq3RW5IfdcIPqatO
hgiVYzvisHZQZQRTVVoiD8MpBBAm0uKz7qudmop7J1i2WnCmBdPB5cK0HQif0PAJ
9wpCNB+fSkOwxtcJFrcrUPE0r7ZWM0Z5pK4InwiA0Kp6t/bEl8upHd7C26JZR4en
fiSqfXIkpspYW8tr6Sb8mF0Tnq9kd/QepYZ/g8Uwj5NH/V7gtOQSGyJUSXhCbckf
Mn+Ry0TMF+0zvqxS9tBeDiNlXhTsOsed3jzSaBpeSoDoiTIL532KhBUC2bkOyrKU
3pi652iAc1SYBXhc7V7XSYeuXlPNB1aVaBG2wLjm5qgLwZRHeWCvLp6ZK7gfWSdx
LhT/JZwjwP8vbiKPjPhJJM9VBNMbgRtQ+bWeAVj3FyVrDCIrDWdnX1ILUbMQvgue
bPtVoEjrct5Ba8e4QwtZBMku/CweEZXva14pdOnnAGuptlSApA2fYCV41uPleg8Y
x01ovCsFYYk1lbyq8W9TmLZQjsbzZlCqM+OitymVrxvCp4CuTs3kKGnG82/6CxOS
bZRS4IiTx+w7edw663N73ECgWxqdgVjI98gAsye0K7/bY6sVn8R2KytlhfVSk2Tu
OISpTrWK6ZoAg1JW8r2Go64/zskQ/Rod+U0svR8kKw24WoOdhZQfycyQHQZ4FTXs
cndX0auOQOcxCUR+wY3iN+hwksoQTxTeTJh0ZPwV2v9F+YL//kIoG4ItcwXMfNBB
zdFQ6o14dtgTPmbGlZFFOTVmCx5cmQihmRKQn0ZJCENXtjgPtY6KCN0MNplpFdyf
TOJiulJg7JgQdRlYXy3y4NpGG1kdNsejnAmUmCfbqSYakAnO3lHk3hhoDFNnTOCV
t/aNMWI50ZGE5VQCePsXdU17kmWU6/JFxwzZRHdcMPy51nRip5WtWE2QGXRZ7OQn
8vsFbjY6SuXuRkAzV16WKJQklxFt6S50Dl1HPiyPkPWZdoEE59Vb31auGMsFjutV
PsGyA+8dp0EkVgoTVIjUF+aoisbYtU3hNgbMyi44nKLb/O2uF2BqZSwW09V2htxs
M5qcSX3fmx5Ruxi6LV27+anBGfcKQpWOV6V8qxu1S7QZSTl/hB+3yrP723UNAo0S
gd2PiolF03K88qBpmZobNwrnRgrj6mZpDiJE1T1ONPJlJpJAoONZMtSBVA/NlCXc
rJVodkNDCZ8TKv8tO7xKuTIErT46CvkbLCJJTOmnxnQRN+bioj333RiWy74TjYH3
8UlmcfQQi9wHuf3C0k7paIVJ2ec4WergBexl0EF3yiOetjkQ1Jrnq5LLhSlLW3I1
ShzLE4TU36m7MKr9xbOnxQ==
`protect END_PROTECTED
