`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chCLJ6g5+y1XtJwOED5v4Q5BzEP2JjViEQYzw+eDkM5eQTaqUhx4U5E9JujD+XCV
vMZClD9HeO9Pza6T7YeCGqB2o07L3RMqQoyZaNqR37kjgpFDbk8DY9BfGgfwRzpm
mNJEcA6oCBaGYKmP8lX/TZy7xIOJnujcdzcqAwi+hf1QgXGhFqpXU/aHH0pwEnwG
DP0JGRC74F4VtXmlA/Bca/0Rp0SnD87AWduoEtGAxiPCpesUWU95oMFV87Br/L/N
10Da8avjtgXmTrQB7RxVtiYiH574YILku5MA65jAj3urv2E2pthRABDcbvn19xt9
Q5CkTiICncBJg7OUtIoLdhG0Zglf6N6ChhaomzkadrfOE5hE2dwdW98uyCJVyf9x
igUL6/tEniAJBetqpx1rDcW0S2dzYhJ0zgRqtrlnSi1Ij971DQb2/CsFNQOwzXkZ
MkWL5M1E64FucleDykNlgIE8JdIp+TUFOKUGYRqFsqloCP3NoHdm1zMgX3mdPhfL
BYnKO9j3yG3Q3tYA3GCFZc9GafSqEJmvjKgWz5uR76fzPtzyvAyp8ObKqlv8btPl
0cpqf5dbUxz9mT7aowh11g==
`protect END_PROTECTED
