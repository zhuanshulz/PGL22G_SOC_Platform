`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
90G5WvvKsXDdWZV1WsQCbhOBZpHriz14bE6L1Mz4yN/ADUgndD6DvrcRA1ffVZbA
L093/nkcaxye53fh0r90BLQ/QntvLnK8HfrqeOn4RCql6VfUz15fYTLQkcjqMo/G
iQxDEtFS2+g/y5gLQ8Wl9ZLMYBuC7BkSjCdRSyBaUIb4SKlH7Pn9hr1HctiXriRh
U00oID1H/pyiBalHCqUZs3Dexxkr9Bdi+ush7sPxJuKxl5k2IFWJZu3m2a7zFvg2
TbkGL+OKBCbXaWFQe/qRBOtZeqD2PWp3lN8/iGVdAKL7QiucyPgGoIa6yPzkBtei
ZTiPi2CYj3oo6r3ol0RwEOt5cQQxsYGbYP1WwFpIxDT+wjbWZg3bUn3HQSkjPd4x
+AU2LFokSjMWkEJOnIjVKprVNBc09lwI6jV3sWnchsd+cI3WU9r457uWSN+YrTTB
ruzKvxClrg9yX7OUo2W9X+v06ruVB5F+C8F/iDJfdL+iz39EKbZ++LvS9ZGAr0/H
JKCVbElnOp0ZhrkT1UY034N1IZp8FzW4iFqC1pmSJDL4HN66BvgDvX4/hrR7UVAR
+LG4MoDECrwwE3QdN756exSjEhV27ommfs0Fu8+TP4IU4PHbNYO3IQrDyuFQ9bZF
5lzK8qxA17qOnU8YyeU/c4VY4ElkkzUa4C7b+VZ0J3Uiy1ivYXJnCeyPL1Fs8BNs
66NdI2eLkiDQU+MNiJonAPeMwD67HMGWlPNYPYSmD9z+7anPvjdlH91kURxkdfIv
ffFJgbfezDPojPoZ/tTXGC1eeSGeAkorKGvAQnTTcV2Im41kQOzDYI6zuYJGEuR0
ztYsoTU0+s0bp3b71awHTY04rAAwGxXR0yu2jLupc6Y=
`protect END_PROTECTED
