`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
McwauDj4IczdvfBcoBPDSAhqzQ6jmhSlT1kCSQIb63wNVwwOwL3pj84ngWfgZD4l
iSiGU+5i0LpFWh1VXZNgRYgcQ2ahCEEy/wtOHmQVmrUUyKs9NZnc+DapgwPH/AHw
Dx5uJoliJhF66oODWHuyq5MWOHt333kQaXak0eUBkwDpppFmS2QXyIYGiQ8n8GHJ
KTKc9dIrOE5PbexfRgcgrJQby/Hybd9ZK7In+MfZP3kzimh3VbiL5gOl0vF/Tt1X
9FqnsLHjWRAGliAPuodtjBTaz5iNu8zqfuvXtCILUV0lcAd22UF42Zjz3siTqbxg
S10091KmHbWCe2zcS6UdIibq9UYrETzgQf0Mo0U0chUynVsYCdfoxcqX2580u4Pk
51KvfMohfkzWM/3CH3mAoOhrEcqpsSTDxuNSmhgIf/eQkyEfpVcJkkxX9QGDFIOQ
dgnRsNx2U85Oa42V6CCzWIDlkVfKIxuqpC13nZno9PVtrh2sn350T6HZQGwvUwH0
NFIqFg6MNkob1o7Mm25coD8c3DW30qKUgYVzQx/OMfFbiCmcvsn0wHWgYo88vYfv
TpA51AHu7ZmYZ3NK2sym7A==
`protect END_PROTECTED
