`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
56yhG3HYw5Q/kGynEblGnz8sR3anZwv+lSYZ3r2MeQ1YcA8rp1tTZ6f0v9V7nEci
VS7dJJxi6P6yI7iZUUzpbGM22FUh2Goy6fu4m95faN8xtYNAqt3FWSaPkqPinNq0
QJdts/gwGp1yu+I1PJTidNBuE67l2hOPgNTB0FaUAUVLUYsxgZ8eMp2wC488Jj9a
XHsD4K6hPfYZrJDRHZZ8FNdP2RqoAnBjO+rDZU8BED6Wpo/ylLQo34WV2MtfoAZ+
Yab3gGZCsOeWB1LHlY5+1P/iR3Xsn80We7EOkhXLGzdKblYnvoxoIFka9DUoGu/2
WTuyKl6S7yMwjMHeiWmd4KHK70/MtPYZtvs/HPzH3oUxx1/o9Hi3amtbXYjEv/qh
dirD6S1FcrPK58gwmWDn3UNh0bv4vCGlt+PvF6zfGQLztOusA0dVBfeDd/ZQ7zOX
WTCmT4YKkU+ylIwOCFf4vXZaH7ARJEGS8YYgXAB+5puHMbEYkUndl8a4BNt1JSvZ
xcJKM2Cf5UK6cz5nAfjAl5cwAGXOZrMQNfhRqZ2LTr62J2ItFp0B0mhI7TzkPw5F
7pJ6OEp0j9EKFq2q4vfGggvzR3eIjjLz59BS3PvWbIdb1lbQUrxIjfyzKLEGe2L2
J4AwoBwIMPQsV3z6fKOa1n+dpFVZE1PrToatwuVxPLr2rJ1THcgueaCkEe2Yl4e+
shDmHvxymPeO8WdmTVA5TCydL4NhmYuhnnVPprdOdcqFWeOtTaQBl+46CRDJAo7K
l0jgQGNPpZeI1K3smdrfQeTpZJrgTAdfFxj/9cN4AS+0p2fP4y+9t2QyE+ghB5bG
VfsrUGV5+9x9OF2HC97YGdUOQwTJsB3Y9anwukMYoyE+vg81/Su2RYsjOQx3061o
8pwsWrYRTUuVkhv/4ZOftQMETUMrfPBmVBr4MvVW/gr1MsXrDoGdW+SvYbK9IKuQ
21tgZT1Xaf/PPjeyfEArB4W2g19haFgvDhNT23s2y7I9ABRh1rXTuvB/CLooYsUn
ouA3qZCzpnxEU1Wey1QtodSwxLHxSQp+0j4nFvkj58TG/3E8ZoQj/J+9Cw4drkVD
bsCA01e1L/2ULFTVEMCYmEIkbGQHp8XZxa3y9pfdjh7LmmHf0TsAM6ryyqgjJnfG
bUynGYR90k4mLIgtQzy1zDzb+0gV25LvdU/LARRbf7X8bkz/v8BT8IXx+NgoP2nu
LvChoabu7KCg05K1s5qEgvoP2gz6opIPNIK6hQFrPRYvUZlF/MUhWo7Dmgvj6t8x
LPIbK1vYdasxJXtrwYqKAACNZWchsBSoCOp1Qq/3jjHmsAW0sL4MCsmsx+8NYZ7E
f+qyeZCZbO7AhcIMOGPDgSeJbG3LdZrcdYHRS5czoPHHfnZA+IhIZZzxTDvgM340
lHwPUhZQpc5Z2mVBnLiH5exramGKnJX900JQ7ipaFGFhQWApA1oEw+uoMYX6f2nB
BqY7PAaZLcZGs7IuT5EpisrHBf4jXt/SAkGPI/pMY6zxxSJlQVJh52WaBLgkWaEs
3o1FK2OY6I2ViaeBWFziT4A96svHikysSH5+AamlftQv16dR286EMq7lk/oBplZk
wNcX9NXw9pCbgm9zfmkAJ/ZPNXmWLo1Ihc7Y3j7YrT3NYp2v08awMrB8LAf2phXt
mIQQQhEnwE+Xrlghm/Mht7aD/6GLLKT4OIREE9/Zqa6Ju0iyJE7XwxhR9vE2tXEH
O1Gm1CrL4ASLH4HYnmRLCHayEqZgC81vwmpfMCNKCKEsp+Lm9jm5e+5mAQMSCugO
Y4+pInqeEZfu/kgAvvHl8zPiHiI15hmsgQZQW5aNidk42IlJLa2i3ORISvL0hXfP
+RoIe5z8hkdHqlQV4ojFm/H8LyNz7M7lWvWlSlgp82FQXMBACwybnJbtVwmrXZGt
LYyXoyjceZMtIQcpsv71UYDwsw+l5VWf8K+xdL1GtlnBh7uEihUjfDXTPFdcQTgT
Rdr8dTOoIj3sb+189rUC3Q==
`protect END_PROTECTED
