`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0LaHRUBLWzgi+zLKfDTcJwst/S9HoodarOPfN0X544EIAsVTSm6Xg+u2IYuEsSe
K14Bkuu9WuRJLo5Z+RTUcXidXh0nZ/iEu6j8grw25IL+LIL0G8nNTAvnaMwUxVNd
l1fjCVYR7+4jYmtWeN2Nveju8N9RZ0HdWAz4CaUy4eVZ575B0LJ6ebCsea3Ae4wE
qbqSWlTVSULNtzd6RSD3sg7swkkYlE3vI30/ZggZUCQUnvMLTSeVrVsR7y+qYP5j
9+5Esb5fon/4bX+XaUc5r8GT2376iaT8bJO9jKhvCaifMX1KdJgrG5q61roPham6
rk8Bwn1EwVpTTBkoLdUT9zQhRJLy/NhpyFx1DD0NYsD7UpkH9BvBsZWeGmy9WlCP
Rm0lkuWH4muxuP1uhWvhXoBxLW8sQu7cRyQPFzIHuEJl9cS+/3mXe1PgHp/IKEy+
4krROXPb4QKS9rr57ZjWOvIvGv0YbIJUtMsMvwbDD35mWmK2Gc+TEiOszvXfP2Cv
beUVBWcqOBU6EpdLIk1eba7Sh8vyWTOAjTFhsQIshg3acnfcGyoB5DdMGUI+HYR4
qNPZswWzaYjbnWb2w63Vq7B09Nxem3mYiffiix7Hf1xcsiSKxliYl35aqd98qvil
MDU2hXb9L2vglQVgYXJWvclw75WMm6Hb7h4fPU8+shOlHLGjuZEZeXUTXBW0FQX3
PNr50J4nuuy/HlDAz5jITtfJY64ooy3OBoVSvcCHwgtNsgVzAvhGC4yhB7JGkaRo
NcshzIalYrqgxd/6W+uYZGxteqlhb1iOkZTWOhOTXsGMB24o5suoAvk7e91cHIdR
Yjr13h9E8dk/I7CcJIcaIHvUiuKCj96qBSVcl0PtdEyk3stABspU2S1rQppb/FbU
AvmDLL1OYDPmttb8Pruk2JIhvcyxodLHeFmTKQObh55eXGWZBz/sy/996kAqwb3K
UYVbjrHU32EoH1cVsVrna9IJpAIeBEhrgb0vk+FXKZfqoHhxM0jUIfe5V4LAyvbb
t1un9sx9eJTsmfn1XjAhv3Ef4J+npGCEx/Lz5jut14S2UGjAYM4q4G7vnwyO9NTx
iBbZCzQMbRpSz9F07UOJusNff6ckfV4slNNBwsFvibZ0o76c0ZYGg2hYX4EyF8Bc
2YW2SbNVfG/qA2sndPzqse1C4YFQt5CivpjasEZJwnu0Q1sCNjNs1JcMfs+KzHd7
lquOrH4Ua1R+41OkneGboaA47ZCoLUcz2iihmLdIBWMq/mFrroSgVD01w7pHXp2U
p/C+5gYxNUcSTSG4SQh94a8e6P4Z3fqapcvdRxJpu2qxSXtl3xu98iSE5tiB/oJb
uTXdwPsvyAGsdl4NgLityuQLXv695cJfPORNBKYsTOplUOu3CH55SvxqgnTbG7eZ
/H0pl7SGG/ahvgW/Y+3u7P37eo+WgFPic5E7fsN/r3ODV5djT1eH4fIqYIiDV5Dj
cdhFK3VL0xfXmPfHaUld6h8uhl1ND+sdldOHcI3XZM/UszvodBxYFwNEAF1O+BM+
tL9o6nwHAxv7TAv/i7GPFtwCwSsF9POwSz/8l6uC2S0AT5ePEOkUUS7lG5zOXDAB
1vaUkZSm4WqClyCXQCEArKF6yq8BhW3SwQCFTrtO9NKF4+/GZKOMEXZdqHVrRRfZ
uaqLIM2jBgwd/wKdCsdYGlucJ0mNnl8GO/vbkyGe16oR3PjC5E7i0aYX/ax2fGHN
NhZB9Avjo1dKA/CEbeXn9Bbq2ttZqviFLS0vW+eBUAIOuBVtcjN0vxdJBP3D4bsA
3+YGWMkpdeihvpelSlhKusu/lVCXAxIGDF0amIv+BsWy3/0C9aMWwZrr0eEXiJ85
DY6wpe6NVuRrXY5gtYqv1PHQC2tzRsRO9qUZp+Qk1E2CkhIHZWmfdsAEGLegsgQc
H8RpG3qh3T89jR6kw9mra8eBg3mOBKiITDtwwl86Ogv6UjHspg80jMTPmI3ryTIY
uVHzO8eMX1ikIVKbNqndcUAjru6XaOLSMlkivxqKAZ7RxmhKnpv5dVSLahCL5PP1
3va8YT0aOqgHnObCFLamAs3Oq0SdXxqACnjiRAUqrHofgc+/fu/21ElLRdMotUsh
zhN/abT/enYzBtNTByA7IdZKUXAZbEAWvt68RNaxPB4zT0HPMJz0W/URjT6VLcL1
cbfpS+w1ZuAXcgejmDOX7+3fqgJyx+NnQu5j/U4ODodUiTcG//ZtfyTHROJAQquY
u6uiFWn6WVF7RiDixyN5dwic+tNIPYDDoksGDfqukiSMQ0qpkAwkZGCy6IK4JG5Z
xZT1TFN4Vi+7NyzRbdcot4xja11aIKzNQVuP+j8NMvdWkJRIAV3c3yRbHZ/WlZ7q
hvDAvWlksC6iKJmhGrhJYqiu6mtEHWQotHIC86MIaH1UonSVfEyl9tWM4VuZuWww
rwIr/8WzI8Pm2W7V06ODJsx7NuhOiHSyRxRYVAU9TWoeL7U2h8hGHyYDLmpuQmJ8
FKPo62XtuRG+C1LdSsDFnhya/8+/mOvNY/ByzXwDr6136SXItsFoFuwqwXAykI0l
dD1mT2x3Vsn9lboXZA5JG4u+k12FlccvTVYjwAGtx5AzsYFEK7LFcxCUQKKZyX6o
rgw10msme5ZTU+nn6NZfn3p90JwRXqxsK6RI2NUk2cof9Kg9UI3fX5l3wsEwtDcz
iMVhspbSnuFJ2tfbp5XyhPlBRCik1SbEJgxLijCYKA7JE3J1LA719vTOV/4qlHQ7
7eq6fvM2DDqjxD8CuRUcxT9Dd7QuowiLFM0t8wzHb5x3CT6ezxC4/ATK44BiPaiR
SmxUH6BayQWJA2wZR2/YTbDyLzMfe+GdNXKiiqNUVCs9tvnaOYHpOTy+KGwZVgci
cN0BYcH0MBOPBga1QXKcerneqxAw3r3t+pSgt5mXZS9Ow3b+gHWxoo0gwDPHA4bf
Y8q4e2TScUyr2u0AJiQ4U9rmR4r0+yYp8cyc/pKuIqPxf/I/y7ajGC5fZMzZ3MVV
LeuTaWPa4X51FqiTtfEnfbY4dtBq3I9CStV1BLfo684ljTjSrOOvxH+JmJzWZeMq
tCkb2ohtYG38OtzdGqG5mXs+dWYD7OqvV+7J3KGAMd3x8c1NzBenje/2bz9GMW1v
EauTa4FyPAYFP5Fj7qwTTAOQEbLS1IcplB3UfVHcvrq0O+iiXf+tn9Zg9tkgPViP
cHGHobNMI91veE36FbfqmIsDfrOx+PcvVCP52Rs2lpo1ccnwSjoNcIcSEJ2uWoGZ
r7J3zhVPymDJ5rYGro8Kd4u/+33eNIhBkR4n/Jlj01UwBdzw9o7pri6oDcEuNOf2
gLCVBlvC3lrfyI+xYJtuKQ==
`protect END_PROTECTED
