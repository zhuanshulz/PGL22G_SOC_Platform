`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
42sfOh+1ysu9oU0FXcYqXn6v5HH3aaFDoB7Le9fgy6wc9npz2W5n8wM/4EJw+KtE
+Qr5Vj1dVZD7L0YFZJES6nsrqtZveDn/kSmc+56V5z/9yG/YBfBW+nFaUdG0USDI
zLREmqo44yg4UfzI3476mFjjUfvth+HtLA0f/DA790sB3Umd/s20iYOFVetqi6BC
p1w0QRnkUGLBYm8z+jiIGO/oNWJU5KA6/5UXcOOBNJ0hEq11i6gLSoqgSVmwbKys
qsSl6YYsHRACgONf4NGBGcusaZXCPqjUIzFUSJw+zu8NfYKJbWgz2z26qprnoCcG
UzJhEnuneQyE+zey/3sJCPPXz21CV/y7J0jpbXAzUy9VPsvzYy5raBNdFSN4BY9B
0AT85ri8zVKyKQltQgBMxbPw7LFBXbl+oJrQ4cHLYFGSSJVVhPujWrSXlyz7oQHw
BQkNhY5alR9Scphg3dxghmkpK15UP7KJe23Wtobc6JivpmrL4QZaTyeIqy8PTKT4
rBGWXZ20z6/sx6EhYAK/lFo86lIAwpxSHx3kPOKskeJVdCqqXOnnxjXZmyX4D5I6
9oLrT8Uo94CTTuPIEfDNCv5Q6KTtUupB3cOvXuDc8QODr80C1spJ1EB2Lf/DVG3l
VprtqYk6ewaJHtxRLJiq0i6+d4BgUlEXeVQqpit5aI/M5VsBFDoC/sTpa4K+5go7
FAL280os1Ye7fbCuoYb41qf43eFrDRNJWPG4/qHFKE31sSOVngmnNAPZbXC8ia+0
X6NgYRXuujf3GoG4oyZCAsXDOtPAsyv1n8DJL7IWOB7+XxGXjRAW7Tuer4RTqtro
gm+icmDZIVEXoJQkiRtHBI9w/lhlqIlqNJBe5hYmSMbNtpnEWG6ctNUycdIA44it
UwzyJfPvoQWR8DxwGU2O16o5HUPmS1GDJbR/Wv6hNPJKWyq/Q1YgntzYMjdnmXF1
RLRTWhcF+1/iscmc5MBtJe3xlwIiESUO+ZxabizYuKD/RsG7GWC/PpS9OkoG+0yo
fDw0JhUBHGr4D+3CwASLbS35U0VlXINsaWCNa20pcfFrLeUwzc0V0hmC39fDimWP
qtGm2lnkOFRwY3luXFPypbAWv+nxLkcABea/9DCrQHFWHnr5cRXWgQyt5NUTe3Li
Nu9VQnX/+ejya3L+9zFWHlbGzGnA0o+3EgtFIE7lrZk=
`protect END_PROTECTED
