`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wdzE67+jyKmdMATv7fzoyL5IXBl6pR3jCxQQKyEtbjWPJTP6WuSLSWSULCnUYe+Y
qkeXOaRpCY6OAIi3QXyrKN78FL33tDe5Rm5NZTsWL5/BeQ//7pTO+ZqQjBMpxIZ4
3cLXTSPfD9vM5r7IAp86CuUOMLbAi/OjAT+TjrDmeJZPEvenpLbjTQIHpr3KlzO8
10M/mDhsDK9rKiHNcEHg7kuyZI2GIYjr05mpUNyxYQukO0vfSY8LxJABfznsy9Fy
eePicfdDt6WjY//55O6wy0Hk3BQfcaTUqvIkUdBjy2/ungNTpI0hCItBr7avpqRe
vm+hLSlI3ss62fPpJPI6oIjagE5b7Yu0tdaEPFzu6OwLzrupgqt4izDnDXKzQEfz
qjXILkP/xkKEtkHBLZS0G/Z1wiziv4fZxt33748EGaueM54JrQ/qOuUYosdMEeZt
VFfz66RQpeIB5iCUAC5fdByzSdKZkO/EV02jE3s1WFuIju4hUILwwD65El81C9+6
3cSqaPtkQvC95LooHEHnbavFq/xyPT4UNyFLmoPZg6k=
`protect END_PROTECTED
