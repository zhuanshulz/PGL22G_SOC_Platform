`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4EzmTCCSEHLWlQZ8OOXDEy90FDkeIBoocxADz+Ox9skSB+x9FGRR9Y6bHC5WWBm
upBTSKarmarEF880hbCKDpJC8SCw50BdcUiQcc4sjjEkJXP9lwnlqc5/uQkGoFU6
DPSs7daR8NbudopOZ+6KVb/vVaehHk+MUdePJ5eucVt9Z365InaxaiAbJ7iVKTij
CDmyebF0oUe/SQ5IOqLeT8JM1TFoLTOEsIHV6Ucg0QFvwqblu2NzSNCl9x/oOxmZ
EPmra008uCgIcdUWgdew6qmhQaFVY96K0dnkQqPK6sCRisBRx4C9r3FBfMRiPB+Q
kDAnE4dRTC7d9ZnkcRh4XHbvBiK9hDKjkLl+XPbhlNOcUgL3S0MEqlWdBLMvje53
jn9sj+y8wAyf3bNerzU16XtRrpYNzcdPLmMD7qClaMOW/CZet4/9ptR0qYWsaX3E
d3N04F3Rhb1OMA0z5wujxK5YOifgSfwNXj1HRcPtpPnIJbEO+a8DwfDJSJkHEZSc
H2QMeWeC6sujf2Uzw1wTNDILi6N7X+BQ/GegFt1L+DsfnPFnOeui068XxlFDFA0n
3z7f43vYyrzb9tTK1xKsuBXMi3R+6osBrdzL2XkH6xjpzAb+hlrYzGKQICEBPWZ1
gu7HexuawkU48oVqasbkMFlTLA05mwzNOx10urg55DMnlMiRxvnTZXKLRqyx+mcX
BBt1GIq1SNm17SzLjqfshLyBA/j7oyHz1d+OyiiAH5fn5XBVUM9Rxe0rMfBbV7QU
ifDJ9GBclLl95Ewkqp9fljgHxdM3ExONMhBIpmhphWDNA/gPMnM1kHSQdtjBh6c6
Ioy25bPnv+Fkg4Iq+laGk8k32ErlkMLy2RDPGCwqsKOzowUVB94AMGapk5JUInk4
RtlBLhlfD95vQkCwJMdZuwZU6DYo9pW7a5HKHxrsx9AnwN5rYVzL87FoIVQvIkAa
dHydVdxuZBCS/tdHFOZBLj/DO0hvq9aLV8/ygoXrJelDl8YHZxE3HKfMDAFbjCHW
2ZJEKb7g1wr5HvNTzSU3vmeXhseVZp5aMCkvYglovhVkzXEsHjv5aBmaVLmRPMoD
enXP/I7NBCsy1CN05EPlxbI1IietoSH4vmcmIpD/28BnU8z27nnviuaDjJder+9Q
soBRb9SFsVciWjCidDB6t9Tg/N+EulUPWZadgSB05wglAstCEjgsfrV0hyAE22Qe
AkJAYyQdzuatofIiGcHrtfuhI9PEG3DZgu5EnSzxns4afu679nojg27w3kCDQ+UI
6ajkQH7ftLXQzVThw1PXD++t6H5LVVBdUkGzaKlhGOp3Yuu0DSgth4DdBfSDkPU3
8nEYKLlXoeRLcsLcOAMWqnPv40rASMgyFSyJPq5FFCG/IxQ7HT+fvga2SnG+wKxN
+hlmDseSJfX3928/KFGH6P72y5CWQfYNXeARggcrD8jqrR7TP6pFFHUXxMdp2Jg1
fQkZCcaKKEqE/6Qy7pd0MxAWnzjErPQzqNcnVkcX3SObNJn3Upgw/bPELjEWV1G1
lnDUdfZwJhPdSAkuVNMUAMMa/MgbLMOX1NXFl4mFqTaIG62nzuwnhvmElSo+jY9f
hfFc934qyShgaAXfFhZLjxIPKJ1GQUf5IcqcRt4emw7hTYUqrmw/B82O0TDUDdVC
t4XgPCe3YhE3pmIlFCCZ/T/WpJmsKaexv/PIqSpSvGyYTr81J9cuQjMv4/DIkJwa
6ZTmX78q1mCoPrecIYmPy0Jbx8JEo7NX7iehq4z8gstpgC1TV8xGOAQSevCGImXX
bfJegBvj/rdMMJQ38udL0wY1Ow4RdTeOpm7H1IzAP8dBKU0zs+uAVftXyxITku+9
u5YcmsSSouFg07U7QvCsZh48jKDEb++qzC24Jiy2mt3ycdf058znl4q4y6a2+EXU
XAoHA+eaxV02xAGRl/GbSZOAoracdj/K2LqwfQpXhKZA+yt7Nh2YAIVV1rKXobYL
vovmNyI7mSpvu2n9k0bnvPm9s3u38DUoQhkOHRidc5XTRggZUe7RJjMl2MUxI8oI
RBDytgCg8nkEvg/9QMVJTG3CTwcKsLsmZmrtjjnD+oLXsHGTj1LWBAXV3eDKsjDe
cpQoRGPY7WQVWO8C7WUq/wc5eZrjoieSsBQkt6mCfrLb2NCwxSvxohe0SgTgOW2v
nL8ju+3SBwtmSJ3Godov9tQaY+FH0vTPZxB5jEyi3IQgnaFN/JoOh4p6OQVw40U8
feGIsKQU/3x96n5raNCaOQbE8iHXNb2iTZjCubSyQwAhnv98exz/chablZBBSyuO
USn9Ue9XnNdWe4MNFfsRgcFzcYaner9NC/e11N+AcSCjgeOE6u+vLeQ4Nv21n6y0
U/CyKILMpCdpy02a0QRlz3acSnWNm+sgDcRo75loaqFo501rLg6xWLOsa+Od0X2v
1gxEgCD17Tbdk+EzUAWUAsDKP8v56w5VAOVG5BtPFcmTHWnnH/AO9r7Xb81Sqs+4
bxWzmiAucZnT2cyM5eBBuLE+oFkfrHDuOLGZFqzHHPuRdhO0DqCKTdfO6sw8Zsdo
z3CEe6C+RdLCaeKeR3bhafvOcyyeDgDXJn24NtJo/ZkT7FVFeRuCui4AzB0f2b6y
1xYKtGodhMnwR295UnzOzqGL/gGgJlgH4vAQIOQz2wx0H7eKOb9NBZmkf5oBn45r
h4FhDvMMBR/3i3b7AHMoyvhc/EwCN7+NNDky0SJ1z/5GPiLHO/dUwJINDsUFJGgn
37mZf9PCkhXTwEoV/a3bdCEPW3Ap6uspaLeCVmvEZi+xQk8iUMUwv8/JPu7GNNpy
/vvjfjEBTAukT1FaspHNphvezmNpyqj8CM7I4jalssyw0HgQx1GUnOFwyCNF7HyN
bkzMU5OSCrNJuYLVRjN8bMSiSx3jOu/NQVLIG6Q6QBzc3Aa4Sj8VGGnVeLgqEoNc
iu52GaI/3lvPFVQA3KhovwXv7hDuHZ5306Q7aNIeq5V/zx08tFp9d6fqGzgfvDOw
mP0oZTXdXdy5ruLn9rL28Ir5DReieHbNMxqUnaLBEuVLBS7K2lISQ08kFY0cP3bs
9aqBu1Nqw+yO+K3zmeaq44eI9lxLaz7IPjeFfEIfhhlBWb2kSBel3sDHZabnTnWb
DWo1WvyRNJIm2ADFsZJmhA8nPwNXtebrUAdN5Rcc3YbJ6VdqvCW004Vm7G96QSHR
kYNHm0SnUqohuIPDCpVSUKIU6eod8t2ulU4tcKgk0CB+UJgt/V/2Md+ldaV1bwxZ
au7n/bWjmfyc1FebFc+kHBsikyoVwz2YZoBRQJfgPBTEFyt8JZ6XvQJmZCp2MF5f
4biGGzb9iA6tvsWaHOv23UJwtjo1/NHNJT9ymvNLBDu6NQrEJy/UA6ERr+VUvUWy
k5jOPb1+oDuR+CDyD9k09FdJJMnI3eF3abiTdntCrXo7+sDN96gWpkmBly1mfz+C
wS1P/QISjafqkvSMGHwjbkhQKchfxCDknDEIEIga/jUlNUfhkFkKd4db4JxqQk/v
PLcK95IMSBPVqocy8+PW3/5qOv5qLlMclKE5pgct5sDuoIwpeExXCxmBs66ESVv8
iQ5j0NImCMQysFoLhBxv7nt4Yblw0mUvtABN3Z+KBwq8xhVy06NqKbsAYctxwFvn
4G+QXs/E46X6KgxS7I2+Am9qC7QGBvXMjHp6lDZtAlDh2cf+JlmnCaClnAq4WFEx
TTMIeGiSg0QuACLPB3NezDxVfP9FCo2W4GEy4JjCEzBCJfpIo43BZBNSy7Pz9CRc
v+i5SK8OQWqg4eYFR4g+7tPbYItXUvuPNJOUT9kXzV42KQ4y0EHYAK4iMdi6zz7y
b6V1JaDvUbwva0OwvLl27GtaygnkVHN/kb03OUHAvk/MhmhlrK9+InvrBBFi2QXo
Ex4/XnsiOvzKEr5ehxDPKMULau3mfNJCc5RfjkvKpLFXGrmaJpBnw5PMUVs/dPyV
yACD1GXjxOz449qNZOb0zc/FkP6eoSqPevACXalm2mgnDxoQTz+Iq3GrGIhDSzUj
tP0K3iOe/Ce51ttIAFCHrFXANpljvfGsmgl0u2tFCzvKQWsHg7XbXW6B4vQ4EjmP
jDKqh8pa4opD86jnPGDp5B12rT1V+C8E5QgWVSUA/3q4fvRNsJGpw6ZpEsCLe58x
WpH91w5e1aZgse/Q/RaWDdx5caDjwHdZkCZA/94tUCeKGKitw1g7jg5Li429edY/
CR7pC5nUAYZpnuI9TPIOerHuEe9oMBTnzFWU2k7ZVEh70MKZIVKrogeEWYqU78h8
AopMtakWqjOrs34MvD3B9hatnncs93qHHTTuSIN7GD7NaFa0NNeYN1mfpAXj/A7c
4sGeCLWdeiK1bKdXwS9x8d+QhvIHqacS7C8WWYz7TWbFf7FrpAm6VZ6HE/gmdNgU
rb9LFumun3Jf3lW2ZTW9kfwIKaikWm7AjVV7xApMqm8G6eOCnnHIHGLXx7ma9+YA
WSwwaWCDXFtrbqAo+XDQqN8ezoivWJdN8JT/bb7IMC0zowwnTPeBQVWNQ0OlLGgX
QEGE9bVQ94u7FaTqFyDlPlh/iQCxLcodY5GxLroq+rGAagFMAr5k4u6G9/sG9D7d
wXm7eECbaV0DgvMSXydEIw==
`protect END_PROTECTED
