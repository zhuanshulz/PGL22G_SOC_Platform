`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9tsixffIR6e9No723J2xrGy5Ehf+9DTi344tvacKLzIM+D6DCP7ILnQ5aSDN/pYo
5SxxAxkAdw5LL/WfSAYrwnIsm+mPojB9rN8nF5fOUFL+JNqP8celQJ67eY+IFrRR
ZAAQ0qCRSLdKQJp1aQPod+qz7DUJUiOyBJVJGyPPaJk79NboyAb0AZQXpuz76Li7
4kUgZtvaLUYBWeGRw8oYAqnWvU/X6Z6lynwfe5eh2pU00q6oSqggHGoaE1NS/7u/
kIYEBJ9YmhOCbuwqBJ+oURR8tLf9r/DYE/Z/itVDI2pDoyHQf3ed2O3sQ+syy7yQ
YRU+gS4OfElCpTKp1nlZ2a8VHrwerPAeR1QpwjMMAmfR6ktBDShmngkG3rg4PQgj
rUAdGcundCgVnfFKlzA3lGHRwVarVzlxfSNBusTx5Dcaht78TBnFaIetA0r7YldK
yuBMQE02yW8+WVgW0EpvwnmJ1B4XK72+QjO5sD3BwttFMs4cJ17Bhg46UGcmMo23
MU3EZInyOn26C77gB9UHZXRTp4Gq3/ni+F9HWfWe47WcpXJvCRnKVw+xLxNyCYnl
V5acN2CL6x7dBDw48R3hSu0Y9loJz7OpjXYXEut89YPiPfpRYwrx192IcqKFQL3z
tw6uT5/TAKLN4D9iJsah9/cBVwhoynAFWaF49bk6Pw68WA3d/UtU4o30TGhKyn46
8zvdEO/kbPjppNFw9TE2rkGpMbHvXNQb7WwuuG6vZyF/+Dh4QIPcP86vOeSgMoPq
IOGY2A0WheFXJ+ESVNtVGbAtZpvhnGZ4m/M+AZMb7D4SOhrGWu+tE32j0Z3lgC0g
HsCncSEFTTRhMWVdy4nJGBKnmQkJZTMHHDjx4um6HEWbNcpCYafLmOIi92g07bSe
PJARjhufTaE9h8oUKpAXK4OOpB6b/Ocel06usmg8vMWEjwvzXTtq67wjcJ3D35pb
Jk6jNFPaz7Vyb2hJx5cfEOBEi2bq63Gf30hBRzPC6wN1VMDVFspjvSBOsjzzKLky
rrE5ICdSQQvwhcsSTmfdNifKzD0xzQtpfzcYVkpnsVo4qVAM8VhWDVmV4Y0GZu1q
fwR/L3FtCzPOxW9cLMWv+EISGZe95tTZ5zJjSeGuz+lcBWYRAsTeoSVIT8WcZSg7
1Wt78SZzVNB32+qDVwDU9cGCSIrs6jSaG8ezvr08iwBonmTk6mI0jVdJ8G1uZTIa
5RLWIpwO/gzsAXe+2VZY7hgpZ8Mrd7UJzlagjp45xX4=
`protect END_PROTECTED
