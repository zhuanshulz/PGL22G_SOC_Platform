`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UbdB/ygweVFxL6jKHPHbkp8rv7820b9guYK73EdiVJr9pXiiEmgQHKt1nqpHpYqj
TJ1zvs8XcHDme43bOynQACYf8LxUFsWu7YvJ7KlDpv8gfYQv3Lkr9IBypRBKDQUv
B/ArckMZP2THvYX27GRJeSGlKWjjPxCtj+peyyNgrV15KY7ehhBjFahk8DMOC7k+
ZvnJDvOJ+x5Cn9BVVRTItNV74x8xW498U+X4h8aYU7rf6txbDxg2n1PwYztGTjcx
R4qCCQwjhlcgcTCpX2lkC/1wbULmJSHWMsv7dxuVWM2oby9YC7yxet0MMte2+aMe
qsZ84Dcwwb7c4NAuhkP/kEtkdnsWhGFZoZL6ARjHl62YqxhIIaj7tM219258k0eg
IziPs+VyyPXAefQUV0KvQGGAIF9bck1MogRNkSLs6LFd6O0dQVgi1ElIiiczSDNe
FugjbIQVxjLQRGXx6ZEDa3lmejApV46q5FKiCBnU4/R/eORTjvCCEDVFcpYq5jo/
JeUd6yFvO3Vo2HKqfGwDJYuzhsG3lkKF92vtd1VWwDr0WDYeD7iLVMzm1Kti0TQF
O/ADajOMBtsv4F47dv4KG/DmKDaRKJUK+UpWXaCbcsuNCJ4e6mUMaC/5//MNG5oS
hguJ0Q6AiPvzvnkwhQuHQdmcMnORkGtZsLgh+esfR3/FH6G1X3k6fFlVZrwiIpYs
+0Qd4NEfv+FL3DTfJOY4ogBphJnRQsScw5VSJW0HlvlSZAIuSki8vcud+0Qj1JUW
XX34yKqm6u8daQkree9EYwmUQpbEn2YykWH40cCDoNn800e4PCCMjI7tksaxwP2j
WHoELJSLgvzRvANJCFa6SKnEVPQg8ptzLUjwE1UW377hrQEM6exS3GRXgDW66Ukv
wFKSYOBbHm5h2TYEpnQevki4PLb9bvQUmPXC5eyAZWO5qM8wOMexdtfqYelsPWL9
FbVJ0SBIf1+DiExILO0epvFmRZX4ZIYlOhEPhZDjMVb/Do0nGSAeh0IOpyvzQsma
meDpEBsT1gHnBNk217/W9u+g9S6x0ng3G+dI+0gJHpEoxPVFEna/e/gpDnOndwn+
hbHhF730X9973d+s3zXefkRCCaitYkDhW/Na89DbwFZ0Hlwm3zaVr0xY6E3v+C9B
9P/m4rGMfcusNpDEGfhemwsdis+jYT/pyU14415JQRUfkJppTPPXekTMHJL7eDP4
PtDPhQbXgQVhVy9l5Limta73p3RKVIkOcWYvOqq0XaJ+c5BvuOZ8Iad9JFJ9I2zB
`protect END_PROTECTED
