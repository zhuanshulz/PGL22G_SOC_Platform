`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xjZ1TQ0PcC0y9RK1qx7aiL6t9GUS2MFQmgnu6RXgKc7o59SKwX7s5gKe3GLFs6A
wyE+c+ZFBos1LP6dkWKokjb0bzyhZwewzIz6P7i5DfRHPY8ufMUZ55NJ+z2VMVmB
KnNhcVX0JeDcK1AJ8jZqPMzzKfYiUHwn6VJKYaaKuCkfKSjaDBJkH9FA/ZsWpEd9
e9LciUvK51NEUTM+iuLDscCq4LQYUhS/TI/7rpl8f5aHA5dK4CVkSFLvyjhRtlMt
Q3nkb8y1uig+TrOjTXvz9f72poniHj0zO/V+a2By/SxhKlbFU50XmSsDEfkwIcOR
daweS+VYRFZzA4RCwETToVA6IM5sWBmRpZmMknji4SXT93zcWlGoDO6UyzK8Y1pN
Q7rdKEiZMw01uEZweX6xIQapr7WuubEmkeGGjxulDaf143Hg3Qp9jqhVCSeJRvL9
8FNfErMbOCc+UR0cGrAygec60dsvcfI2jE7O50s5CgIXGwt+CzVtM0BOYB++aXus
48JaSDsppiMtHmXEKFkv3agqM/vNp6xJHIFGs3E2n0Gxz0Y8t760M3J277r8J+0q
91HB78L+82Xpn7OvIqYfPg==
`protect END_PROTECTED
