`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pllRqFiXok8DUXchnXOGzHujgK1PRVss51OdWkWvcUZJl3EuFfhBfaa5PDfT7qHf
GKOBeD9zHdlUNGQLKNEHoVxfIYUJ9q8yysaCUleI1YXGw6mn4STuP8M74Z2YRxrq
7ukC4TVUZMg55c+Sf9+DZxSgTypIIg2e9t8D/QI1Q+gt82EAN47wm8CmljhVVNxd
7xlIVqnAUlcJwaavxH5lasUkF3EwM5l+GW3F9FkQBiE4AHgncA3DKlC9/+CkpPsm
fdAMLTiMU+aaz1MujoTwmWOBos0mn1bGAJgnrPQ1jQLg7YraKT+rKhEKIH2GeuWp
CiKleLINr8b1vGH5oPZdhuWnawTIdg5U//vDvXSKRbPB2CMie2SqhXP9bgMcspmt
sb1Cwnqqx5VUxoxxsvaG4iFE9O8nL2mknTIb4+o9bthfQjq7bzixX0uew7UHUWPi
Hv+3f50TZE97ZKRq9/lBn64/WOqjbYCX+w13w5YbQnCu8Uwvf/XX1hF2MpkN0p0a
UXW9dc9fWWLCsgpnW6q5EeN299IQo6TPQ5ec7B6vVMqNona5zmroeiItprsdgKj/
ajftqX2fWkuv5K8kXR7N6U5Zc3cmDYT2KA3soS+Dw4Snyk/YW0wHSbG4Juu4pFcz
zfLztAjRuFAvnMjHX2GgxMeaOAEq/nfNR5Fw56h4y9pvYmS/v+xfmxYmhldl/umM
j5pS8T5xl4G5eaebRonj2NLEyqI7jydxHkDGy9eearA1glx7CjAdjSnnvUzofrx+
wNeyARqamXixPvzB33Caw8I9AcejzdRAsWoOyCHXRxkq4ulDOhDUD3KvjXN3uIyw
+Bt4kfloV1grDPPxvqiPFpjEfcHBG6MUAsRYTrLHkww71FaJmY3FtCy3gcTzLSp6
Xub1rtQf8OMhFzpS5+ESsGo8KhYJGptxiPPVdmvxNXa51ykvvkqEPCVE3OsMMICa
jddPBM2W9g83XvgYhRgu+0vne8Wf9/gFQVxQsvqck27vQoy8zudxmf4kdEzkRAgx
8lmYQX+oiYgxrtnnZYrujFUJ+An2/QOjIkiL/j8cYLymprkXtr3HNudR5bZn86EQ
xMo4GeEFJ6nLR9+IIpW2NIy4hQpbxwVJ3gFOxcbGlOLLuSAo3hZh/LyMa2dYdkY/
uGdgPVgZCJQpV2jWxeG4nNMLAKJ1A2I2aYVn1WzL8yCMefdX1JSzFTCsdBL4nHF3
1E8u8bMhkwN+nwzCBgCYNVFpErgf+maRUk5t7rtMBEHARePsYHs3NjgupLP4ga+r
2KqVHJnwQCrhbTWW5qfWZ/UeNCc7Vj9VHyf0dNCFm8Ho697fquo5GuH8hSQdn5eJ
qESX2ZPP7E86arwgkDGCfDmG8DYrJSTC9Xj7HL3mDZAP0w7FXLdN92ngwNDcRL2L
4H7GVHu6vfv5UTrsIoWZhdZdnVki5+OCC9OOvBQ2fweTwMuuDOr9iPZEXME80YD1
yhbcuITJDUWbRzN86SrS/NQrAR8PZrZDhUSwA7gc7Rii3qvVo3uBCBQQxFOjBnR+
YzOdapw17um98DEkKNUVU1xV+eGa8Qj/SoAN/2k7USGETCNkmwBGoTCBmqj3Ya4R
f813KVatTSVPM4mig0ND8N4us9vPerKRjYMl0vR7XKSMW/Pmz91/R2Mw5tFhiOst
wOQNzE2SJway18DYp/8lUKQlVJcjpEoL64NLB3mN6jQ3lxjjN24ANHW6RCMY8Uie
mJXJj8PaqQTR+Y925ahdudgRn2VsBzVBThH7pj59b9oCTugNLLNWWGC8QwFBOYmm
pQTurq5PERS0JV9f5H/qQ3KIvpUrWv994PhQKv6yWY6A4nnRVlofu6YnGc3K0nXs
ouSGg/d0kJ6TM1VN0aR9ptAuIyHtOpcURFkQBWjLUPvYo71u7FlMt5y9oEdkZthT
lKGXYtalo4iGMm7XebiDsFrpg8J450SnNJ8yT06e4GzKtaUReDAdbhhay5zNbl+6
VL2+Ql+cry9OGL11zWTLahABx9k1RjNTJ7x3rJBPaLChAtXBDaKKrYM/o22LZKwq
mcd5vW7FfkUTgleQBnRzLv9HAtbwiNNwD//FefzIlDl94d5Cg7F2y50ajUdmQpwx
ytW7tipEd278Cg0KAUkkeSKNtW+6ciOAj7hyYR6M86/mUFwhNRwDe4omjuc8VB0O
CnSpv3zAddsetkgncTviZjIMnZoWgYgVxor2cHxKaAV8oDrMndYJsAadyR7wKSaA
Q60IZcmtjMLGjq5PkFDK+HF5pIzoPvKZRDnnZHz1KCfXXbm2jgW2R1j8+qY3AKFa
SKferjQLCsYAQBrcW4p9ilkzGi2SgYhBIa8BUaqeYpr2KsGIbnmFj3lmYGwbyQPm
sDbpkpJQ6IMt1eGRRle6h350EMbiTn3YVmVXDrdyleNH7DdLR3MA52ZjFz/aRP38
jU6R72MDGDm3VP5PuqyVUjf3fBX5mtkFuTJQVKfWZRfKmMoVG1HWmpH3Mwaq7k5q
yezOeZFFX0CH12W2r99Gy+1E4Z9Qz8T/AOh+lGuRe6Hsqw0pk55y7C4qxK/a+3sY
Oz69qFuzw+0FSQOAXNX3Ykg/3RBPEMX9WaKIXD1hmZDavigwo5bkC37LxDLzMiSF
Y1FQ+j6Wo408NJqsL9pApuNOcQiT67p3G4cbhOCQTu7C0YVZp/JtEmY01N89Hzru
XK58v4X1WRL8RNnEHvWqqbrI364jgWBTpPpUk/xlG7dj5o5kC75oqS3oSvYsD04T
RdEupSbdJQpXvTSRyIV5wbp3u+pJALIixKqIsXVg6Qiy0ZgN4XkS8iz70AZE7it0
GGPEmfo3S2P1ydVNoHwc9cBWrmf0tGdO0CWVe2XI+OrmOltpOx+wRnp3HVQsf59k
Wp9aSAhVxrL7pxbXtnHhVNu74ReQsz24vWrgQEYvz9nyARFPk7/KvYoOWS2kgPmw
t0RnaXc6ek5on33v+ibSrAbOcICTIuzOE3xn7YpNFTYt1imYEolrfqZyys9/Xkvq
3kB8uphYIvAXOnFX/L3PbHOJOGnecyrXBozuCvVxCOupq2M7oHvM2ZM7qKyak+k3
1F24246cOysl6Kt0u7IuI/33xxpqwNRCDCduE7UrfyTzDYn6MXM+pu2NHVNpYiM7
1pknqNKZQWjBdIQCbJLBPrCVFRnK9mnMpKWApUiUkLZ34zaRqaxI99OKJMeXaFu+
pZg1BDPozHLBPgYgXa4LA4snc2gdJbIhU8LnC3aZe9PRHDkkglGF2UkzPvtvQEif
YLZAwP+mo0wZeqaAM2QF9/g6EjG9MHiAFC7FKkEHDXnYZzKtdrP+aQcdxKIvR1d1
4xdUKUScSc4qy539sxDKq4P3moz3gyAR0NKgK26tHMuduRPmgEeyQntoH9IdJ0HX
COwiqL8DKUzcwLyLb8Da4hA5YV6ylyAHCDhPqAGjmwYq4UhgOJcC5eXjKVLv0ucY
AhkrLrZGg1tllkZ/r4F1TqbwtPN5iIL4l8ye8N9YTxW0GE3Y2zRc1mIAXua4F6Xo
Xgu4TeZTDjGOM6VjKRhzROFKY/QcX7xP9UyPdo8cYhWMGUFMLnKwcivtqS4RbsaG
Awb3ULb6n/bwcP9q71/8rtkgZMXP69bqqjiTrT+mION0cewNY5ctaJyPpZnvz0lW
AKHv5AwfyWcDm/iVMgAPCcykQTSyfSmsgCHR34lJqIrequpvNsv3NpMDsoKQbK7m
bveL1WdhNaTHdL4J3R0hQxeapk4LrnAlGobA0ARa21EPpGZJDEdBII+1GzdTzHph
+iOSxb0aSUtpH/08Zy+qRYoMj1ClEeSbBHJ1XLQgOSQULgIzxU3ClchxFZ24B2PX
XdkJt2A1MsoGgAnn7ceeIIfO6e+4DIKi/bbPtSzaqFaNTWUs9MAq/997NkoL9s7g
SU4ugWOwXfnyXUMbckcv11iWrgPZoUVu9pd/zX2RcVSZj4vwSXojFRLLC1kOFiut
AgHu+NQj7kya+xNc8Hsrq7A4V3xEdOGWp9OoiYS8etm9MFyCc9RX6kzkDumtCuMd
l/77XogWXpxW0ut/e7AQPsEkd8z2sg72lVsim5FTxcRH3I94xUubwNsvk2POIoTe
Yg1I5nrlEMvcxL2XUtSjKKXiDxOrv/4LEG0wFioowcrVKr2tzyYAPG43c1/nXUzg
HvpP7K2xHmEmNapaXl9YoWeuRuy6H2IhH3Z26UtUpNBlX9q9JI81pwUJ67uslYFE
RRYRJ26oEUjE8urnJ7+/M2V6DqqwWfTYoLog4iLCuuqION57jlQfXGHmn39hzKfX
10nD2foXNxzjLtIPvVofcQfZGEid/TL+osoKsQRCUjxJzb6+e1BuoWTNlRHHPMDI
4Zsy+uUgk9DWhfE8Ygb4i8EjlHz9oFLgZrL9kGRjTq1Kxc72147sKAvGK57K2INK
a+SUJkjS8ii84Sk1QpIrv6v9K7w4pyY3+HJt/rL9qsvxosak7hIIjR04G7g7wdk4
Hx92LzjRuZoFSKtnxF+YhADcVbR449sju3BTbc01c0ZA1OTTsXRNzyxMR60IT0P/
AQ6nUF0UBrfYIljKOft8mDfqjSz6JWY9uc1d4o6R9tZ9zecIVaKy+QWAVWKtsdPV
DpqfJkQDefX13ntSlMTThKZsym8Pq4mExnXhPffuJvr9mP1QYL718gdOhak2mype
QDMjmuOMtE+ZTdbxX/pUAJVAqjwPU6aNY2ckBnwPMZ8ETOIEE5w4nTJKZwAJ/TC8
YNqfMFtaG8CX8YpV3U6rY+j61npaSOsVPHsfer2NiY2EgPm0ouJvdD5+qH+snd8I
D5MB+GGDRRmSlyAO5+Y8/wcN0pU+lyw/buxHkYsXZvBObsVLarJHApVGaLoi/eXf
64cBAFkrMvVdFvhB7sguw2UwZCf1uRBofVCTfiftdCOh+bDFbfcPLVc9ZDCyYA8U
x8t9JxRyr+L5KFhXs7eOGmuQaRM/ZCcLDJJBwCBLeh0yQSRL9ufBcQyTzjoFDitM
aZJtueuEJdvu5ZlkYiAzL06fQ86+dQ6NzCTKBmVDjCPXJai4PzPKz1rWbWWzYblE
J6gjEO6L+DNnUf4wq7hiifFjdDhpqCfzjPZX79LsaDgK5vqqwUGvQTh6XqNFk5We
rsQwD6FchQuez+Pw1GckPCsKhXpHw5ZVHiS5QkID9V1/o6j4goEhQD/Z8caRrb83
UH8U5BQ+RcYwmIOdeEAZiWXMIzY+nJqSGntj8c36J3zIQqU/jkhf7ZDdrsMj2kKY
iNSFp0OClEBBPNdE+H/BsDmDzjB7BqJ9eGW5lowqMAWRc2g3dpR5I83ptWV8FtRS
21oenO16+cx9fs11bmQ8ojvIBDuaWdBUv+hLJ2yZWmVURbJGBtOfyhMfsazrbhTe
PSftyDPvf2ttNgryqYYhVQR6mab+qNWe7oZol++B35PRdEDJoRwqBExV4dkB1EGr
7OqwFW7MDhQSYPDeM+Z4p6L4WdKBcAN+lSn9A7thOgjnUZ2XeL53tpeUFlU9G/V3
cnnFBQ8BAcf4sQDAzvCy5x9F4cvXWhxUCOsPuPIdNQQ42wijoTyJfxnZdXZ0o/io
ImeocEjk6B1HtUNj7anlkolY1LG+e++cyDvITcovBdfsXMouKg5/B0rMSheKk6NP
eHCvZwKzABLzdEDBIcH2mPGgpeCctkgeDDYq7nEQJg2UdLR0h9SB3EutCF4hAV+U
66ICAZufVplLjEOX3vTdh2swop3jzPJMCd2DB/x1syMCF3SXlfeHlhLioeyGn4GT
WVQ4d8wMeW4gNmFFJS04MVmyCRsmRf7kKbSZnZyoSyK96w4h9fMX8M09hNrHTtNU
TKRRWvgU9haHuVzgx1fdzC7dcTG0SC5m8aIikXPHxd9TrzDgONZvYy8dDky2wjMu
nNZ78dQOSsj1HWDpaExeL1+un3fhm5+JxS0UwEFMhHIzPKuUR/y5cz2a9tBgYzOC
w9VxkeaWwGc3sRo/5qm9olPjWB/PI6bEzvX/e5bsm8nHyjjSIdg96SHnmXwMYIca
dqSvI3KDna3XJekVx7VsWw9yHiQsKJflpZXHKDrCraP7U0eug7nSUuarzCQaivTw
z5PMNVuMs60yVeIKP02t88VqC3VonFCrqlOvIC1FLwGe6Apn29LGMYwvWnfkMQOY
Htmes0WeTDgsecxiCZFSqdxkfDV7zB9Cuuh4kSBzSPS7KW8SV9oSqpNY1Gzp1jT0
GiY9p0ftjodnrslF/thxyPf2oYTCBSVcvhOynm7MKjk+EyaaYD3ME85hquoOmcHx
+1MrKtIkVHciovX6ALHgljlD1cbNMqHOPjMc2gn0KFIoYK+vhK4tmNuwCYT4I+kd
ZHIxIDRJPnv/n9skKaMUDTk3g31Qhs2KD3XRQlVZqKTsJho9SR/7kEREeF9ghrsD
77YK7bu53TyVE9Dbd1kbTqDNjvQYsr/HtssUDpcr4b1zP+osSdXMlB05R7FSAXfa
H4iJfFSA2j25KYQcKaWhbM1m9Zfybu4Yctcg7kGucH8O9ZMvC6xUvZ/VEHPfw9dG
SDUMCi6K5MqMAly+hjro2RbaeQVS1G5uY9zaPO60qPl6QhQVA1SpRRUk3i88afts
q/fycSUGouCHKUqFVvzdKX1vB+bAuj6zO4OqjpG8g1m6kIPZqfzQW3KJbWIFPthz
BlaIG94CjdItkMZi5YZ3Hm7q4Pz0tV0Yb1wfAyCWcNRsyTEGhyA69zUl28M52Rdd
OlIowg0LMHyQ6crxJCjrPysaNObi8t3PiFcBymFmkEx38PxwWSCkCrncNFCANhxH
IEjiqbrpkJQIWqzkaok7thTjCOQE9LSBTGpqLZ1A0A+uXe6WeghWE7mNeShFpAk5
XmOYvuobQLk8mBcFG7js+ZzL4bJgMnGvvUS4nrQR6JwEuW5c8cHESjsvcHovfi8L
r2OM0jPmdx0/D5dZ3XGRPcls2906BEorvv+dTz5Us+Nl2x28yU/OYnbYkMbK/31g
cX0WAOpPGf1aefPGfzPDf/qOrW9hDmMqAJxnFWGFE2ewZ5T44i+aozp7xZM9JOFF
Vohigq2ij0F7k+LEX148bJHsa+G4TuCiuYKhG+/uuTJTFauA130GayHeLawGA5dI
Eec5wt1KAKNgIRWKTRvGH6DxNsdE0fwBskhT4PYFxeiFL1Vmw/MBO6pJJFOU/8MT
OerJ1GM6WWsrBU8XqP9Bkc+PGSvb6g1DRj8SpRXt9VLyWz4x0HXvFEs1lXok9HxZ
pjsaaNT9fciPKhahEAIIakNmue0riFN3BTjjznDh/9Yoi1tAcr9ER1IKAcTbJtAs
Z/yGLcEnUZ2PSmUI7y7OZtrCAg4L/jQZGn9CxmiXhoe6H/jAR+R9eR5QIuu27zFj
kRwunfzGkWYSR6TvyDnu9pktueCk5yhrwdbKgNICc+fzTVC6OLk6tZW36DgivDjg
CmK29qoTfIE6I1CPkD6hRemF6P75BsHNWpKX8Z1B0UHI0HE1wvkbfbNhvaWW2B+y
5pPL+zCQQ6fe4G/Jg7WXo7PzqcUxNkzVu6WLjxw95SJTwvvsJ+dhFRba+3jAVHsj
GV1mAEpF/bklGv+PETsXspTrtTOMkFdZJGan3h7cp6YKV57yo4livLrRE7j8cuG3
I5sqzSs2Lm11Uot+rzU047En7gt3eTHVQkkJat7rPlhS0la1cbr41tnTR99n9iln
sIfgCE3rMdo8/ZXW8A095999wLjP8WsujSlNntDyAFGMB72qKwFMS6fVTBcTrs0B
JV27BwSg2f7WuOvRXceWTNuYjXfVdJehxSBJIgtwJRwiblkV9c7iB730gfSuClo4
RG1O3yHuTIVljyqWKj3CKZWGMHsz/9rt/bnsTit3jk7lsiGOaqC51IpOsKzbrZ5K
3pAQdW5MgSPRTGTH6Q0l0+gMxaDNjOw8K0O3wgK86b5oS7IXm79i3fbrib7UgTGh
4AnenHk+rBTSHKDj3koYICXXgvz0aWgFaiyhegMnzYrU5TcC6/IWQ6QLQd4HP8dA
uA6j+Goql1ehg17LGLOs77Oie8YjPbKOn/hiLCfc31v4HUU54+n8v39jfvEK4BPJ
0s3lapHkCA/JTgR6C3pTfaaPIdXqAlHn0jleYQwNGJn8rQbUwOweujLXA5RPmgOC
91vf5fCjl6vRjnJu8qvzeZpPzzAuPqnt0IGjb6XNwVZMsaWCaZQQ+/mwXAuyAX8d
573USG1KHcLgH9INyrXDxvlY9Ox8MbHicckED3S8/el62LsrGro2vTLe99cbaBGj
M+tTw4eFAIu8ykOGtvKt+4FpueeWIFmnBu9FWrmRCSHoVY2sQnnMM3nnRxYO+PL2
1B35MjJqQfBWU/Av/hFzhwTnvaA7VVSAuxKYO2X1lYaF9HCyiyEKGytUZTHYjHbc
yJwV4V5HD9z5rGXWmokLviFD8GQYuDY7EBEJOWfzW4RmSYfnB40vdyKCunfSW9dJ
RfqDPFuzg8g1CvaMK6ULNF1ezcGQ+DUsZOmj1QzyEHLrSqrrKBXiw71aAjpH+vAj
mi/kY0olcEQSO9aBrw/u3hBhM1mI4GGD3DhCLGfpVsOGOrPABE6qE338PC+1i+yA
gZBOsNTdIrw0l1WGunWsLBmcB6vZJ8xgLaIxgGVVaXlFVmgvlOLoQxniIBIKhUFy
j1BXsJ6K0srqPH3kZkxd0w6svq7C4FmQdJCwaXOQhP/0CcM6ic2JOQ6EHCvQKDM9
ptCoiILguPSP+KZQseDWaTlkprR7tVdMUMX3CjCSt+1qeNpxaE0v9qLe+b3hJ0K3
hZlG7QJ6F+msfHrIaSW4653Y6Pq3bx0GIo/pcF+EUVpkhOmEb633qgwRASa3k1uz
1jLLQoQkhemL5sHjmj2uOPGlAa/Op1zovPqNE/92kBM08XVEyIHJm/P9+kZ524Hi
WeLSE8u8DjizCSf8yjqRlG5ZZMteh19Y3nqRLMtRmYS5ZwVc0QaffjIwk2FP2b1D
FKkWbzuHBSPmgVul88tMMG/27veY+MkFBZdRVUxUOI4ozzNFAnney0b5NEhZkT6+
zTAqidxETIvLi9nO2Hub2W+hFhT/6IX9vnJh9/lwQiRud20xTAu+e97aATc0DPbe
zIqSigqQ9Nmhb1qftCxWj92wg09nCFwwegbtfKynFA/n+tEqCA+/eNUByIP4KWzr
cU3ozFyEqCQQRh7fpIe1v1MPOzGYX3rxFOtbCb3imeCG5uc36a7PoPDo3EgN8Vy8
XWW+YVBL3ICjiBOCKjnkpRiiIunLuYuw188Phx1Q3E2jdbAjSbVE/YQSEDaBF8RJ
4voaYJKtGtuaqZOERChIgu2c/SP0STu2dlQQOoliFonIUJUE3PDN9qJCefAV9Wxr
8jrx7YDdGwxtH7fyToiHmwNhNvaAWeO01IoKETzgsmPfIHCafG7JiWlrsD+5MLrd
H//tH30JqCcxkw/r1jLYU+S1BPJAkqdA/PZuSKjciQ+gyll6yel0YreQG6mmyP3r
0ynZwmzbm2qj9pX/9VIHojYkopIMQuqg7eDmDvbpEQ9WGRhNTz6U0ADfXBQwCcVf
Jlk+BOQeO7IwkE1brfSh+88+uqHPQO8I1XWn7KE/2To7bBaYenCZgOJEqR7zXzJq
eCtPyiNk1QSqTwI8GA/yQPi0YACjmkEDhB8bbyHIXF4G3z3AJ9v6iqblRyQfMCO+
2W7zUIcH7lVmVQy8R2Ghbx4wY9UgR2MPzuUsqP1JCYvPc0nLxgFCrkHJbQVhQYc/
MclQm+QnyeVmHyBxGyVBVxwKihU+1uCEYybrSysERxMUk9FQyG8VnzlPJnnwMMR/
kwpS1i5ovoHGjCL3qwKYFCO1+/LsVCVRtyEWYLT6oh/5OFvcGfNsOYZfgMW13Z94
ZPqF7thY5+WtsB+NXk1NQGZOzvao4tk6SqzAJty5pxL0G+/3xRgompiAA0ESPJEv
Y+CQO/bDAV3J241Ud+BCKX6VzC2XnOm79Q3iKETfimfXP9y9xOIw03/Rlzn/4d7J
WNgD1pgscujpHgv73D4p9yJGGYcFRoncEKoQ0AaCTmwCtpxBIy3VC3krD3t13+1p
BEcvvw6Jt77fmYj5fbh+7pNhjl4msfhyHvjF+hl4Yrh8RMJFvLHoGkjwYVQV/Dyu
enEb+I7KNcw76h8dp/5/OJ7ozU5LEviEpg6TduOW++vq8/51SDCJwNw/roUs8Vm8
otz3VpbYgkCnQCrBK6fQDkisVcKIsfxu9MJszqj2zh2uKcwHt6qfE4YU8V4edzOZ
h8Uqd80gJeHyo55NtGQd2ylkiAlImmZPTvsFNlPul1QXyIJOER5IXcEXY96Rr0Ky
JMoRVw9WDy1E1QjEoxGgigd6D35a6Sf4WUEArsxboQ7VxQdvlwIiwLei8lVs9qrx
b3mNOEeROpPknCyGBmNE0q6JYboL5jgYhj4Gg/p7sX6+e0en4h4ADbcnboJKNch9
10++R1m5Mcbf4tUb5fu/DxbEZCYUgl1tRT5HQYB8HSdwRyPwaqdr5r73J9wfWIMv
TTsRO3aMyAzkMRQilqoLtL3AlzVXvlSlxuPdAfk6lnBBayVRNedg9ENBCJtYtShA
GA8sLqaZSPUUX7oA8sXtSD1xThwLReSotG3yKN/GtpcRABPqqHhJm20dOCGRfJCF
AFwKDWgHy9AaveWwTM/d5YkQpgMcpY39QdUTjFM75jWUg1PsF2I9Nnl0quHFCkP4
Wh2BCC80T3ehPGUPb7XklTyLHjMwzHMyKGqVo0hlOoXVbZT6rEgLz7h6dwjKQhTg
6Pd6hSzHGM2NNrNDdbg5PgfDBgVJQ9lPHMvUWUzfmq3VekMSxs/B0WbJVg+BTuVx
MHQB8ERvNxWTsldtIDB2b0rc9+PLHgafb6505pUGMYotano3yECvnrgAS2NRKktJ
4x3+ENeLKCnzG9vLVGcxWGSb8T2sCl9PWCsnReV3pkmFUZEleZzsHcS8ICYvDCgQ
8iS5g2zuIN6DNEFmRl8m2QFpDqONylzseaRtiTwY7IDsLqJjgP3AxP0vt2GjXoJX
WBG1JGiRhXgV1FmzGMe8NzwkEqvG4YvOAir4fM68udCNDFiSNsTHHTIw1XOo4UEn
BStROb5C5bJOTSjSXlKaFlfSojnoVg+RoUEbb+CZaeTMAVRvrBaSWQwaC5XmdlCI
c/z6hYrDr4ghNZj+AE20xYZ7anniUTMbiTE0vFacStHmydZV0GNkKUb0p88txPk5
Lw5hmjmAFyq++9zxcmWTyruvYe+iFaZd6gMev5MPF8eZmAqJyiw2ZcEPWtI5a4MY
SQS+ICOgMlMwbS0zGDV1qpy7qtkcqB9WBwfJQDmCzNnHkQaGBbMNiPZqtqbVGpjv
UKjfdHc2fhmSAq+68V1GYeuntay/SOa5f/ULWwFYsdp6RJPZAAbOluzAh5EeKSze
/2jBAyjQLTbRNWW09F55qOuny7aCLBREmJVE9nXKX/ugwPodu9jtZffZFotRYMUU
E8StQLWQienIEFr9PFEc+2k/rtlaoJ2dVh8aE9pgsDX24sz0fgjJbT/+iMDPWBHu
QdOPkqb/LG4eTLefTs04u+yd5IW11DRdvbTDdomOn37GqqJWOTxvKI/XuZaylamf
DoRa8p9DeJx/s37APe1HDgyuuJ0XkEFFrsOTXKaxMwuZOLxfQVMyqP5GRDLPAtag
tFd38sA+q+NxF6XpaTIatsSfCfG919W4f3JuFLcX/NrRhqnlzd4P5HzDZgqFaI2C
BT/01oSK0dpKj9tfN7fowf4h9dfBrhpVfVid8VYMGBAneP4IG8D3YtOpgjDLBGS6
tgqilIoslD8pXL7Pe6DbaNQlfzx9rwNPuvH9gONd8m4L9rKY8mODkizicXq68jo2
qJGwvEl48vOPM8KrqVAycvH033r28lbumC76JvElYHMqbzsQwG64BLUQU78MJc28
0/ReFvGaeodPUVes50zWYkEC1tkInalvBPZKB92iEsv4YNFAwQvQOyg6F3smAObg
QsYTXkm17G89FD19I6nLn6adQPYOrD8vXpZ5fGn6OpO+xLVNJ8TyK0o1QmRhZWhU
Z0jeX2V1bzvN0Im+P2Eh4SO1xLjA8+VzkQqSVJb2vBYdlvXyBFLyrVs8AOqmF9Qb
nYgPlO7GJnHk0DvsLtiMFn9QVtekv3JLJ2ORZJVXkwHVkb8jqc5nnqgiBjruBbAy
1XW6qkQaD/26ijY1HP39giTi9Pc0rYy9SQlon3HMvVTAlqkJelG4VRf8SThgLu/3
jQpA8//O6+evMykEOUwxD630ijrrijdvlstY1Qb7o8u/pJSlUHQc3H+Zgbr5YIl9
SYuko4K+qUEeo2wnX38pnNcDGdyHIoN49ohq1wK7SG8LRxJ60+nVskndxraIVhOJ
6ntgXrxi+c5KKLieWGm+rKLHygnLZgPcvWgzUuoc+hlVvnqjSyUwVfTdW7lJygUM
dTjeQDHIuYIgXPztbxAjOenDlUBnFiiteTeRj5w9Sh+y8HPXTw3HN0E7MdEJ6hRo
BgdUG0KdXDCpqvFvIphr7/4ug9T3o/LiZA7y9+1C+KsCosnsII/2Zu+QWKRdI/6D
PGQXsPF2czrLNzWA47ABhhgo3WShCzqkROmrLJJtw5BHsyc852HwwBR3QY6RGtDO
2sqVEzzu8Y1h6OnNvRdbFPOKWwShD/4A3tO6C7EdEyD4EHlsOinHn2R7qQgd8W9h
eVhgL/9VthFWz9Cmul/VGLdY0i9Jhm3IiRs0Hhf8yXCRUEqrJW1Sj4+zy3TRf2f+
6zygLW2KZnOEoS0tBbJl9+MVTm0GMpQeAKMdvzUK75NSCyYotACSApK2WUytW2wa
AcMZT7YNgBxgpG4Wu8c88f1jZEFtIiVIlNtAhW8I2eFirXLNNesGnezy8iX23u8d
86zC5gSISFUSAvb8igYvQbNZPUTDyK4PtT2hu0mdVNuaopwb6bkl1qi6Y46PWYYU
6V6qgkrDE1TnNmrHEpqR+mL24l4Q1z6nEz3BJ85LfhKuF7AiGLjZMczjTxQH+E2a
YExmCn2t3Tx4b8nwyeRx21MIamNFKGIhat6fvRTuE2NHhP0nWFQI6LWV4YyXfwyD
PXrrI/gNtb19YexPR8IcGaZCPcEAoeXQ695lCzpVRCXp4lizUGLiuVW47NH8hGQ4
n2gOJOZWtiw0iafK1cxFjAhcyaY8URO9ytzFqSbFYca4TcraXTUlqi9nn8sYjPws
IKR/mgvcIzcWPs6tkLsb0AuoT504IkD4hk/yvqQt0X42MxwC8nwnzR1abz/1K3Rx
gfW0cDlvTR66bpCeFK9W7Y979AKIsZjSj0cr8uKRpRAIiMeEEmV94lNjnTOWmUua
Tsz3gFv01RO+EqgoqfavHPYJpwQx+kPNcsoA3yyCJoRRGfrxVbEI+C5KwIYNVriE
0HMvAoiLv0cdduJpt9IlpKHDZNThTQYYDGFAY5g6oGV47KCfn9tLrlOAPX6CvcCJ
UrD6SdPmPQT1xOQNClJ5O6TRyfjLOiZ3TtaCZ8OstHtzCJXVkZMost4waW02gvy9
iA7BGd8f8naFXffyV2BrxJ/IVXgJcDDLpPOULvklLbTylVYP+aSF0TIuzin/kts6
OD/fuiKj0UJJQATnKrUNCpL4VKs79efBIC1TDME0RXj5mZvEViODQscB0oV3gmeR
cUv2tKz7nuJc/aYt3Jv4sY9EFM4FA5fSqwYFyw5GaWlz3N8d/WBp68xW0PYMXTxJ
QjQbU/2U3NAVlPFFligg9EzuNe1uN5KtSdofHzJXHOPZW2BRObBcMCDy0AnS3hoO
Qd/N8g13tH40AYFvxNVuyr7QKg1LFM1w5e6MfdT5ATVscy9wLcArdtovkxWgdYdA
g13TTWLXmQU4Nn9/5OhnNqiCE+ErJ18+EEkVgvtcWvbPC1hJKDL6QfBlffFI1n6Z
7lye9fnF/1bn790MnzSszzh8VBYvQENurBT7qQQvUhqGuORKxJxoAeIwlrWIVHXl
sGAG329rS9OXI54r6bE0lR72w9lxl5LedMrQEggRPM/HWTcmyaA+y+CvqgTOV9x+
ULhoeTAQZHD7IG5TuEDSlYgT0lMs/iy2tSBZp5Ku4xTwHngrKHdn/dzAsG0k6IUT
6OnDDxQFWt1/IXLFZfLI4UHI6Al0i36L5hK6DphXT83zFalyyWjD3B6o0rZuetad
2kyTSrT74XXe3Pm/RnvUtXilW9ewCRaui7lCdioqvkNz7bCGylyBW7ESqdM73OQc
MNfzYD6iuK9b/PBtIY/CPKa3OS8AGoNhny7ZMqO6CKx2Orn6ZYcHMzvVtnZaluRt
x33U4ljGHVPPo3LAdYF0T5WHiLT0SQ6ZJRbr2AYKCgdcZR7W8oWS9rYCGisb+5Y6
YJejiloys01okSX7KBNQfHmXadUh69E1LT0ZmOkMM7hB9cEf0I/iP9+CaS7y0t8f
fEupkjrkLBvBDzwn++N2zzO5wcnol7JWGyqO+yBf98ciiF+olLK5qqshj3undFax
IcrUbzQKSGQ0E5VXCzDNCriUmVShtlW/jqFBGfbmfJObQu09ctDlso9WqSTWhMN9
UZ6ZYR+HRniKAFmk+bkF4gaDxS6VddPGUXWV25U9Y18XVEMs86s/sO+NqzIUQz8q
Yohx3lv/Grrb5VXwbsa7TNqBuC05XWgjOF29KgMnjk3C/0wH51MqRa6hwqgUqFHw
XOgtM2VwJaEP69lwhMZudIS9AqsuWGSC2QUh6jMKjrCYdqC92UOwvTThJ0xH6fbW
9eL2id7ZFwq8AsuFA7v32+zxyQ/VD7Wuqb+KzB/LzozY1xFim1Snkxh1h/64rNKv
YMQVwSRWGs24K2vi4ckL3NX+Y3fmWNqX199T5NZ5VPVBHyM8uPuxO69CRMDivQz5
uXHNQJlAYXlxoHdLdYfUkG6UBwoWe69MJXe09z0p297REOhHVMPGz0VI6wxJ5+No
fyOsuv/B2v+rza9qJ3PwsDcdmWIpH+7k2hgpOxOEi/qaltRt9NRtookShJtGbW0H
QuG9WDfh0fva7bxVYFjz6DZrC4igYGxm3YRLUEeGZN9UWORlFP/Gi3QKI+g9y+de
rvuBv1XM9dYnDDv6IeKOAziw78MMBniKtgSnV6ScrNkKj6XsjJ7Ygu/t/PcvxUxI
67UvrE5GBUQQbjup291knT8zl+XUMdfsI5o1kPeopHm0znfICu9XtoHgKv3oe9ff
KAkes3yFiAeHRODId9t58UPGJSTBNTEONDHd3g6he1uI8g+U/lod50yEB486JjyX
Y2L2g4RLYML2+ibyaUhyDf9EfjKpT9h82nRVqrIUu/RoS6O+xiHrHlDhZw7D/rgr
+sVpivEKIzB98xGH8qmauRW54X+nmiSXEifPds7G/CDfXgsRqTaiJ9T97+X/NjvW
xNXcsAXNteqjWPiHVFcVDfZ00ENleFdi8h7TRGzkAnoJfqSavuNiRtdPveT1ATIa
XdY7xAnsg1UeB6C4dFpOp9qgGFmJEs38H/vNRbuprPCRd/zSx23Nl4NJcK1QWupr
DCA3S6Y8SO/4F3mfZXLRIPY/mihKG2yz9oP4hH3MtAvMfu4SugPl+7a+5DIwFLcb
fRgr3Z2DRbvtpt0WI4+tOQg4gmjWSp2McYS8rFWi47rN2Jq1CSu7aEzFIOGNLN7i
7eojSGyWaWRbC+Gi+XP16Wv6uNt7YgNnDGtLioRX+k3UYBldV93snk2kd+9IaoI2
DDdGN3exLpXciFR1fGvMfQ1YiyAmuDXLEDt46c9uyrHQI9e4a+6IqWEn/bJlGRb0
lrjtibh2ucElO0KfETxYmtlNUxgB//DnLRZpxEHCmfjRRpOTEb42kN7FoSrRAnJ3
H1PbvS3BfL8U7aKsIksVFOxT7MyOoObdvRGRZTPmfHbSVh9bfrJ5MBIdGNcVxDY9
ofU88K2unRZ3aKP3Ff+1F4ZH2aqeKFxehEmzwrs07pYNgAmgSNzkdbIvtD7vL5Mi
VGCDt0W/iYy7+gkTusktCxM0MnMdUxDReoN+HgAbWcaoTny4hUkQBitbuctapFZF
jNbal3xedRxlyzYNSzZFItB7zhhuCVpN0BaNkF9CLDbQINDtZUj0ZU5RDy/9PK7m
gJvG+jGJw2HvqZIn3Ooiij5DY7kJufwoinUDdE6XQ081EpCxwqEdiiE5ALWxSQC3
ZWjxUH4hDhhR2dcqrjAu1MNMi50iIRl/+Gvynv3TjUZ+b3VphVGmgl/tIsQPdbW5
0NkwKweVL7HyOfd4aLE6IbaqbuS3oK4k0ontjRKlovNjglilSonqvx4OF4geDQH5
W3BioWZvi3APTNZ+L0CcxQK6pihb1lGZiGpcAPrLOktL6iZxqW5rUAUGLpyF/7IR
zecPMWL9fffYE0ZyWPoQD2fAFrYGETr+I8gptYvs2BXIjwkDwy1JbNoEj/ED2x9t
MkGAhmIpj/L3zzcr0zL2443ZlRIv8QuBiOBeL3q8qB+wD90qvzo93h9q54OqgGDQ
bkyxy1OU2+npxV3xFqrwA1KyBI2JrNwOSdmh8ekyTZnbukvwr2nH26jzRBQNvgt6
E3/AbTL4xlcZ12oOH1etH3JzT7VloHd/x+vNgIgCkNCxJgl+K3rekqrljx6rRmQp
y48Wbqa3zYjKWrmBMpd7re8GzY19RqMYWx+Tb889wUqp0s3FcEbXNwqaLLJotZwb
q/qsVTQLPYx3kELdcYtIDg52X0odz9KuMklPZREfXzCVC1GJNGXwY2pc9N5X2LK+
IvL0XWLqIAcDS7sikwaAIBnpAyp3AFa8+Ky0s3UML4DfQ1Zsp5zmbvvGxNQffcbg
xxyh565htDvdwAt11HEelYJpE0by9FI19x1+g1hC59/wWkb1NaWMPoPNyToPxoQs
0/OwfWAguRlByj5j8Q3EX7PuccDxaDrPAYG5KbrNGc+8+jS40/zy1EBNlJ6WAOMl
CoOugMuR+FuIZYOkn/FL2Q9kF6Ej0okZBqbJx3bsw/KK0gNCoV9dcLFRJnViGS+O
iT80ArOmPskxgo6isquMYtiH13gqx7P5btybx9JkAvmBoa6evL8meynliGN9V955
YrKw6AIo1Jr/06YXW8Zf78klNrbV5cQrnOmrYnqE+hLM9DOUWK8vOOIS+HrmuiW7
jEo8tmSoQZmk6ywhQcneHjaYDTuKux+ZLuByLviCxI6k7M0a9FQjqMunoXHQT9yC
VWEFY3UWERkmtUVjWU4W2v3aTiPu4i9t4zTKChiua1GDtpQ6C8TavGTCvU9AdS4U
bHcIdg5iPdpvUueIBVwVoOOXIEwD8eh7AXvQuEa5wB2XPAtBAMYdgFJb3+sU7RRc
XH2zV+ylRjRQiv95+thpsm3haYYdmFORVS5/0fLIvQqgMdfOEJeVQNmtvGEOhF9I
Jz13N/zFoD230O8ArPrUunp2+Q/ALd+57ZkVywDc7L8LcoFzQGGv8JPIzs0D4kYv
WHsrRkLIadEgCmxb6IFxg3ON88/EulAsOq3j2NwUQkH3cCt/7hAAorXLX/yHNHRB
9EhFxC+nlEtXAzP1pIlidrYtqyAQeGIr1i2/LK84IxIxkUavg4lSODNflw1dIG2J
98Hu2l73V7K/GjlkOD5TG/Vc55ilNsfqRC9tvb8NP4SGtqte/wn4XYCIttB6rJIM
IZ8DdKdn98kYzIbTcyb9uQ/fEU6SWxsIQV6DxK9MsGoG1AvfWp0n7mKn3o/B5FWz
77jlFGHRtQ7Ou5WkRDw0+nE3PeswMrFTY3Wx1gPaksLwB7TcJcsqCuuSKG+o8CFo
aI7K8g9ZVOO7nVidtYJ7Fdclv/qp5KoMYSqpy9EVPBjTbi3yZDJsbOcY04H3hA7Z
/MT5x5jusof+7tKzvGmzrHEMMLbZTwZNDQ8upB68G7wsSh6QUIhIJx3QQpC/MXkl
75pgHqewxoAWL9gV6MgxqmgrMxUPcxtfM9QKyJ2kWa+TTrLFK/P9EngP2o490+d8
0N7UAJxqymSH5QYVyiRhwHyT1hWRS9uCUJC1UZAyS13XFE/kMi9fKhMpD3brArQe
C7d6hj3i7YMksPzP2na0t1I2uFlMHig+GtF5EfG8qIeQ/J/bFS2Llr0j24yEG92a
LWBO+Za99P3NWlkjorWFWvpqvmgkEpEEvE6qNs+0vChNXxmoXgXrNSY6LtRHssF4
5L0QZ+dBqbeFxKbgljuORFvAX3FG0ezG/Wj46TV0d88/066I7/Bl2iQNqTQ9M5aM
IbsMVQn7+4ON27ulSlqsQ4ACU0PbO7LywYWfPDNl0UN+S4BkCpfih3ke7ekjnSCT
or7Qz913SebeUxe57eYJsnJBO2AsaT3md+fstuGldPnomGblKjRypIFgbsKmC0x4
7yNIc3DctU6lEKVCcSvcD/PXC7m9StYB3Rbw+VZJFRCqI2Aixs9NzN3ARmH9ucKU
XoPHLJ43GjGhbhoGCa0X4CJaMhJXvBtXwPcu5dxg1psN2b7zcxSomTLDQveQFLPg
d+JSxx99k7Gqb0vvvWUtIAy4xCeVRvzgysDoT8ac7Ylwa6vQruWoY5jEBxwDKs12
TEfKPQAJ+DLYDA+sRZ0tXOQ28RZ+Q7/056THlRvKuRYbktKeatPV1tjb6OD3GSa9
uwrojYMAOVzPqLaRmZG8HYpNYn9LChr4JHqSn0pgwPrpa1oM7OThTdQqEmEC70NW
q50sz4ZQtkEJl8HlPf3jQ4EDW2S61qFtOh5sfWvPSwnFnqRiRM+mK5K/9ngBGu5/
Orm7ZcRm9lpTGfa+d10x6eoyeBAqsd4YE+Aj+UPfpcKfgzQ/UxRN++5kUhxJmAR1
9gD7yUEeqSQtyB5ASkVGVElRoGaZFyCn1m1+lWTLHVSgPkklaAvtHHWykvCyLYfr
tOQMv2df2wZvKE0eHkt0ukupOZyvDZgVdiCK+OUzQfvV71wpJW5SuCbLjjFPOmYL
K/5vLNPMb7VuA7nD15rmXvYqrRv7NLgGSxCxIxcyz+f0pmGipnsLZzSS5D9Hejqm
r6Z/A24kXXkrWwPKvIH3gCHGXrsdRYUvIogVCwGqPiYcCOzAlQPjaKnegLROrh/+
XEbORUJRSBz2ffPCtE3A/uAEWHtAg5GYJ+PpSjf3R6OcfJD471PRfR7F8yJQfe1/
ITF8gTpdiDpwphQ3cHsgx4M0gM77FO5a3gb/DTnoulxKz7LJ1CpRtYEa/gVCcne8
P4vYkBFmXQxnpPyraaLol2IpJWbsUwrUuU0MHUTOnnCYE+rnwQcb41bPKmqkVuza
pfOG60wOCmHeVyCsIgfI8rDbF9PjdN/8Z9Wp+h9BMav17Jah3uzpXKWf9Xz0KpVV
wjzlIzjUifHz5/KCan+Z/c6lEG3rjVCItlQlcmxjgYtAdrZMOxq2Nxebz6TSyTd2
eaXP7Yna7J6hAaiZcbhQ6ZxUfm9cUIUtkEiPtM7fcHW4YlbBH34mkswPVu3StKj/
h7wTev5Ax1qF2LNlcPRPOH5hEItKmglfnif5Px7nKgLmlBvN8fHo5XSyk5gODecY
b0v5WzCA8RBhhMUrIYHE/DMvNYuI0fJco6ykRwFK0170BOWq08L74YIEQpeZjMxT
l23qU5P8n39UpFdWFW9rjiAyC30faMqpWWz/U+am8Io8rVmZx4WS8yeYLimQDyXK
wp896YbUZuOTtGB/jH3o+IVHrfcI+LXmeiZX7J2Pu1zmKKi3Lg5wr96xTQqaUBUk
A1TcRHW2avyrPkzgO0GHyXc/UlbMslGkp8r4rMPn/FHu9GwIkSsAgXFcSWFmXCGk
PVg+K+5OtRNtATfMzoMRHvzFmgsKPNhx3YSN1+Qu/bt5GNJs8ZPfIA+XABphAj/Y
TXJpumWa0hhOSK5ZWT2H64rLaeUK00e127qHor2d63k/lCVKKPxnj8DpMIvX4OO3
fU3lxducVdzsJ/rAV9ngK8SckL+aW3cm9Te0NnZSTxirwelIgyM/B4YqtwY2vBmx
yVxC3pNVM1ewOLtlg/u9utEgtWRwEqf7m6mZEHCfYZuLsuY+hyaWLmNH8U+8uZMm
6xeKUJsQjQqDeh1thF4YwldzyfhPxD8UR7tNNkmVX283+2peBiTX2R5GojZCYAmQ
uzLYak2S1q6OaCjiQgdK7Hz9V7q7AuI8C/kiZLNv6Wn/hSLakg5OT0ekMlGj7ull
58vqNgiPcra1Mi8tVyqDyVXyTOK4GSNEQufAQMhiHCuNKpERHUFV81AmbpNIPLDb
HcDuDsyHxOXvym9sn9/FJoAzyWAX/HdX8pJyg90+Lp12DUi700kyJ6GhdCXz0Wy4
nYxv5Fg9UX27Pd9XhpJSoCJKAORzXbmou0dYRnM8icf370T+5koEaddpFFzRp8aY
jXLGdSEYQVHBOFvSzp/Wrv7w4WWBxKbvG6VlFfAkha5228KtECL8L59OTaNtln3O
eSfpk+PBzcBBHCR2gUXQKzu2BIFJtZ8ybLXftt6oT0OCEqsF+P86ycsp2PINvd2y
SPdIVIrYl0WHoD/GU59djlXygbMoSkiJfcNutn4dItwVYGryHgTo//PRd1jyKl+7
cgC54JLBXDYcTvmOLBbG07iuFXTwX8JjlEyvfhTnzVoUyiE4k0mBoyIqdWLDCINe
pooIIOmm1jsiJoVdUhfVqYJ/2+uhS+NUIdX3iWDQ7JmaLjOlpni+MjK9mtIt0V4q
NE5Bf5WzUZ1kVrBgQVszifwnjFW9s8nIz5YnvWuIHKuFS1GGwsNi5eVsGkRGr+1X
rMvxYTH4YkzYOKMsRe0186/suAWyp69i3nkZfBx5CFsEkesMokWRKkH7QDN+K3oV
kl7At2r+eQXi3d1Tdvqz4hJS+i/MLGHnoDFG55fZzGEgHektSUlw8z2w4zHlVsMK
wo997e/vv9Z94hTQvvvgFN+Fy1grvPCaiqczQi9JMzMMpfMJ1vIok0lvJ/WfvqfR
NhWg5yFt4wi5Go56ZEeS9VlmDvA03FEVlPYV8Qdse4FRLWKm0Cc/RkBZh2vkahhz
ImT7GLTvciefg/IiEEbNL6U1a2PupJgTY0bLURhFOgVJpfG72qO6PP/yyE5+EjI0
yqf8sWYB0tWuMBjtE/IaDSb6gsDnjY7bRxC22TvjWOuI//m4SEZiM0W6QQwrQiPt
HP4YSsL3avks5s4ftvlrnX+mkMzpY8YYAwk82ZmixeRmK/g0FRl4pdq2GPjtEL7Z
Zkqa+uD5GQBabtuKeCdoR9LvX4cJGWTs7bh7CDqJK1h6l04hQO05kpXIWt+2+3NW
SFC1fY/nFsRfN7MVQwMFVxBHwgshHVD+HVAjgcazLUeUoS39BSZF/NxpCBYYSR3B
8VVZBCusLLk5PkpKlLHg/7ePp0v0a9gRbDe8nExz6kxmdwPNkyndqFZ2nZ0flZ5/
nt+U4za1hI6/FCq+bFEhoIYANXid3NqCOpXU3R2pscLZdhvMfpG4aWA2sgst6a8Q
K/a8x7j9eWvP+ionKZudh4Eha4ka+zpBukoq6bDIdxD3fuO2uAA7CFSUk7tu/qzD
PJstBrU++8mZfWEtYkpgLd+zMdosFISZn08Pq6daQSzjWdzfLmD+XGUdAWt+hQLl
ArZYa0O3Or1cl8hR/hrysNXVUqLpztmEY46rVlVbLl7LIf/3jAnjpzmVJ5FcECB/
cjiHnJNVZS2oeFoUeQrMtPw7Dz86guWdz8kCVWLmsFGPziXDR6qso/y/GnmCsPw9
duAgKT1LyVzinb/4lw95EY7NMkvSYeGeSzyUuJ8CPWQeI6es74AAblg1g4j5Kk8s
rmJAzC4xse9Tkc7MtTppNRQCA67+VTlzU95wkl7Dx9I95/8Kym8MCYIPZRQcnYbX
vzNVNcdPMe1MVhP01Z66n9prixn9eGPkExpG0rr5/zp1fslyjnwkhElh9xnYQoyf
nKbJJCIk2uLk3ui1gXpEoBcAu3Sit0fAPIbj70QUX9kHFpn96WROxRmTDuws430C
xGlW2dYIYO3TqTb6ubkizSQU2xJ+fo13erXBJ+M+bk/tRPW60vDfbTk5TRojH1sY
l9m0cVsRqqsOzvlCzMzofvpRpOUAXKRV/jXiP7uXkA0K1v7LKrFwa+gMQu2f13Jp
c4uQNd+XUINdi/wXbym6ahQXcBa5UF1+3TPEJ3k+j3OSQcz3UrQ2+2jo7jqhIGbR
kY789gKjAsZv+UsS2mfdFEgyfhgAY21+YuQdfXOgZKlHwwA8MTar3mqC1qkB7fUy
q/R08uSJQGBL5Xne/EELiSBLh8nsJJJpM1+40ADYBPnes4RGuoc7dZddPmneOeKf
8J7kVcxHBGyq68L/ZsB2nd94ywc6nolUZ9pooQ+WBG55RW58GWjbmr8NYi1h66Fc
FEhZvlgvRILM6pyROHeShdQSXYaeT3qZMwnYhdD502DZkFnsOY7r7Ck1xni64l9A
vT/41V/Q0CAtq97Hhpw0Dmc5QhDzpcxwHHkInYammLA9ZyBRGIS0wm9T4AlMXAv/
Kh0ShfpVp9Gys01XxQGt1wx07kYJz2gZ0k81QDR1VGepBoYEdyVWOjiW2yGNcBOn
mh30iDcBrDarUvK4v2d5zMNEPVh839z72pQlno36ed75szUQCPM4/aFR881Y4AFR
HG7qO39mrPxQkaVpGy2uMgt2aBFHlkKJ1tkesWFjSwqdWLhw8HjsEaR/LbbOe0pb
jcEPRk+JKrIlHuAEGLfdy94+drw7BZQgoPBRiQxvtekrSioDQnMMY7nO2+YGqIf7
HhEuf2bE1a0bQak7W0v/IBruITMCtdZRB3PsIwiL19xjBtZy2F8HFwwnzaTaUs8p
UEeWSdpSlMQB76uipQP7VO7ysMY8AE3BdP9uHtqM2nF5WBebaallJBuYpGFJmkl6
p3dgwuL8p4L3E3BT7Qa3G+1H8sHYH5gRvP41SACHbwA/GQH1ZmEFP/Y+O8Zt/keI
9nqiwQm4wMp36qcZixhQjc7V+NdAFTlPkYyKOtI7Z07jqxLNEketwJS476/+bJFE
BHHJqISwjmGzBpJVU9MnGN9QVT7hHKeH6W7iDFMyf92+kZ9VD67362i1dnPe5cy4
VuGLaEfzXUsY62D5lEYWQNvoYe8XeVQnSIuenG5P7kjjPdK4bnhpQ3mo8nFo1PTj
Gt3ZfMaFwNxBHshwImmR5aLqhziI2g5E1lbRVsi2X6bDTwL1SM1fHq70cf+//hH4
fzbAANt1wzTGoioPi3hxToffMY2ppkS9cyIBTgo5nbSKZTpctYdPYLW3eLRavlr4
l7tYKepmOqZjBfBRdXsZii/XlNgNDC4FzxVNm67YPfYz8wXItOkKty8U7By8osKM
g2CB2N/ykzGvAu6ZDK0lb9oGj//PoNd9tLXT3zG+2xJk5pL0wfs8xVRxfdafatCi
MBVrOWzg0o+FyjmZc8m9kBxoJNmAoJyVKgS6RxQ9ZP9GjX7kspSfj8opXSWLK99N
7nRTsYyu3MV4xenpwfttan4OJrHOqBqc1v6jSrfl60IW5COjxiyEL+C6VK7/BJmX
JPzrIJA3F363Gm1JABpZLLIZ/9IJXCJrgA+FdAZm3qkNklzDZ2OqDhZ7Xs1l4VBw
PN8h2Wn/3Vndx6xkR+ylP3F+garxe7/dYngrLdp7XQLvkUyn6+omAecYmbAeRAwT
2tk7d/96AMJwmE9ITwBZmZF9DNU+Ml9t8DUylqdTIkIRh2Mfrq2e5MiHIIt+4fog
oA8UzX4N1XxGZY7V1AFFhFsNDR+OxtYw8rEX2p3847LSUvyyN8lK7s6yiN+gqjXj
7sFUjKVdn4P/kqEIiAExL/kYNIVOppca/84BnT6V+AEGxPwkSGF1z4M0OAbyXyVF
76dVYoTN6h/hU94Z1CjMxdcJHbKBE8bNGFNpSlE3KBmNTrtLjvUVavwmb7hUKqqs
1GGtZuvoGC62wRg0s5viIUtLSxpNqgNREjDLDSUE695RmV2jaQ+anNX4PUEEluo3
NAXVCbhjlnVF4Y617P/pLQSm7lyVrxVHsId8KHS/6WhAjT7jZdfhwX7usTbP+hfZ
8mmcVcaj++6M0Gvh9UgJiIwtxd7PdT0c0TVpypphOP9Uf5KbPmRt8QTdUE5LGtgU
gYmkjwu/HLzbmhn/fZAUvQaEbJEleeQiYDip3Bad3JhWqfih6Jv2DtirnSppO+gL
ThScItWPbOVzvcdKnCBwCvyLBzUOIMlAP/PuKKsxH1TWRLfppak43s4GbwZd5b50
bomttAYi3BNAfWkwVLewSoQ2CyvdBHMAQ+cF6JLErW2IC7HLmZndQ1cI5XDZxAp5
YKAvhIHzofzvxRZVr2P7e11dAv4M0uvOv+m6ccYW7xMAfstCn7n6qJTRyGtJlWaN
YaZ4P6U0ZjPlaYvz290Ad2xXNsti5azz+gCBjHSLRKD6IPSfho6oy0mwHqlXC2ZB
EMkRAV9bZxxk3G9KKfsXi6KCgB4SE6uh+1/emcYsvmhUFPGwjNXNyxiJV5Q81VFQ
F3thYY9EhZ+9jO8mWIYqFvIGfmlWd55fcshfe47vWj+VXdeXk8jbKrn4sho6TEga
lZST3RC9+DGc584rnqSVBL+mojbv5DDXy5wi34y8I++pV/GRPrE+KM0rRozs28Vs
C7w93Rk5w+dHERrxvZQuJR+HiWPg/3NgKvsXRtGdsyT+siYt4kY3Zl0SEgMgc1aI
HA/e3smi+YpAF05ZwlrFFYZisy+TWX/kycx8llptxSL3I5htRRF66gJXeHwEf/Lh
f5fjmbcu3yD5owFQ6W0PRSPdbefbQKvxCsxn5BAh3p3fL6qjDCE+gY4ixaMmaKjT
9sXtRUKsQvYhkyEqTEsgtJPSwb0o7+lQrLfb4uzax3JIx6rgY5nrHYuf2No9Vp5x
0hOdteqxW8seFmflNlAXvvexBT3w4V8G7gGWXbyZCXiSzyLUl/IDBev20uXRp4/i
yW38qB/pbUdlh3cj/wNMSb8pBw9tYLeJOlxL4J1qkN+YD6T2jNRKXxriJ7+asTXq
V1f2yJChO1snBpWPgIDtL6U1rRDtmA68u6TvCgLhlhfayC09+vrhMdrKI8k8/9fz
xVABDzXhDbv0w+DjSWU2cEUiG4BRMvzqnTx3kLVHFzPMUN0rrHBvifBvh0oWgpMR
ZzU7V8fSpK0nNMjC/cKpzG2uv9Zad2mUKSUNzqJeCAD7xumJTJTnjUUYz+uSCFhF
9ECbn9CrQoIAxsoM29+ATsVeTYdqKH2djp3bpPEhkgc+LgBGAuNiGLeubwfU/gkb
6C/5/vGV5i43kauXup9iYxASdW/4f32cTQPLcqGa3slAvmLQP+mjaHiZTfvqGbp/
lmyyVIo3is6BdGJz4TCxPp0Oj2KH8R2cj6MvXfIkEKLakV2utWtC/tmg8pGAjAou
NrTHDMZNxmH5jmjj3+AaGc+rCLrQPMRDN98tQOG5wNRPF0YBQ6DYLuA8DlmUMj+z
e7sls5Kvy8tbKB1aH8v2Cc1FSsJPE1I/j0ZH0hVkMWf45Oy95ATxHbyjUlk6xwvx
hG77NXsDC3Uh0FhWWdPRtmmBb2TUBp04nA3Z5KkRnRtjuOE+nu5h+MrXre094S3c
e/OMfZWTjLYe64sQMBNpSanv/fiFJeKO1YYnsEYyFghLclOoWsTns1z/Lzha+8RM
DxzO550PMB54l5qhmmDcLxpb7f3FSX/h/VZeoQI/I5Zp2W8Hw24pJgZur5I9nCsc
uYzlvyJ6oS1mbnsSpoaskDE+Dm2nnG63kXg9b9u+XSXcecKlAE8V21+Hwzjrj6Hy
IPP9OcnDcbMpsNR5ywYJa/jOAE/4j4wg7lIUzfBa9vsC2sSkSFyFuqhgI2YJkrt6
OXb4zOUSWw9+bOEbZrpOlZvx2S9bzf9PFHH5AkeL4maJqNtV82rsACjo3ednxn/a
qLNzqt6kDSrQWHtJoYAD55PYnPJ8YAEs43AMgZsY5jfkBPYaXKs91rw5xGY4SH/7
Y/GvR6wRVu5rLY9+c2i52k2cknD/80XTALkytJt6x4gyEkUJAWrErX4Q3GbqMEV3
148M3yvHKhS8N8rtaiPodKHWfybbrWnBvVg/m8+NcnYYgKo5sKXU0U+VG/wzw3KI
A3XQmuK3Q8GUty208akfbqsz69oXufl4jzReZdI91Sft+Shem++7P00/9ab818ku
QVOXT+3qRflKQA0TznbazRO/9AG7FmYT/dkDkNIHOIw0TqtYnZ/X/qEm0Vpzd4cJ
j6ZIxniRWJchyXx1hp3WqU9rA7pmhMOWYNo/D3+0vrDUMl3u3AUdkPloO1FDoIc2
UufJnGrqhKLmZ9uedWw6P1pziV14YVVvtNOpfX2RfWlTiSu32IUbQmWWs0ng+x0+
N2EDqzFewn9/WtkgZ+/FIilqRXn6WvsLl9YYHL72CI3uG6RWdkAsFA8DnB9X2FfQ
ZC32C1tN1v8z2ZAiIh6C0emwMnR0TrZS/PP9+NK3SncD+jW/qp1kQCh0lnkdeJfo
Vav24qDCkDNc+QwqOuaJoBalLqHZtP49FVYFPeYddWXPVGEo3uzd9bzZGCBL5+qO
79RWBEMhPRJ5QERhIB52FFkxvxN18xCax3XPtTfnfCJcpZw4UylV8MuQrSwJ3Vf7
I/YhjS/a0OTuH6c3O6t7CCeI57pT/Ivj2QbbvuiBNZgFO2a6TdCSg4Q5gJPSistO
wQ4Gs0t9iezJF7L+4jnZsKHCfHb+UlVOE4c6+y5a73gL+K1QjUzQyMI8ijxvnqk8
K5r7s8O0X7JbcGoi6s1rm9qw7DfZ6M9XXulAkSAlyC4J1t/OqCgNLvKCKkqG9e96
f0aDqHXVpVnBzVVC75vSqbfutXCtxziEISOE6pkjQlBeLwA4PPM2P/LfNS8PY1ue
4eeLl4VevMBCIIAzkpcgB/Q5BxQygg6suTsacFFyAxuoBo1/RZPGQEagcRQjWXpi
vtGSV/Byli6QJrRsbfgBgzdiH4TSGZj/VKlN63ZIMayoQUcTEug5CZBHNDpZLX9A
sSiK2xVaDMqJ9dWGzsxvqAFz05KaVbN6E8LFGs562+OXSRkSqXGHsyT46TBHBxrm
UUTG2LwCDLgftKrsStK5H7xFqNr2V0RiVDmM4/syXOcm+HbiclzUAZZ89B1gLgG5
m2idJrY6tK/q71V2VR00k+KiZfFep5FOXrAG1OeCi94QVdcjmq4nwufzLkpJzpqA
6RSYWW6OCKrAT5qC9GerMUOhiC4tPyl9ipExkxp3rOdGphz8JCMJZI+/yF1fsY7F
EseBtJ4feZxtdZmz51M1wx4vc0a54GwMlQBKHnWnW/fB1Rv2fzY6W1ZNk/7NFzOB
PCfeZfgI1Dq7DgQihaiK8ni16xOxunHl8GsAD9ycUDKP+cIvwTeKa1Zm4suyuBfU
rMEyHyoV2U383prsnCkrvCdtpNYgN79NmkahOz/2QdkKec5PPvttCXLUHr9Dt4dT
fmJiUjhcPUFLG0nrySkax2FEkfjkRbzlQEoExaAhP5eB40qAdsA1Gu4O1MtF9U8n
5Wao6NzY8E19zH+Rhesqmxwq1VZ7WZkWuNcC362pNCR2UmBKHeLf4lOdDHqrcuN+
N/CewWY5MpgbmPyxjlxxTnkqap4tGWAgbfHdk0DZ20jiEyWJ6YGURHb9gr3qAoiC
6BTyJBRLt1jlOWOzM5E7F8HBIKu7eSUvFK123+6zCrcC0Ddl1O73EbfcMQ5IYbw7
X6DwJ+hI9O2UtpbUkvMfKqutfQZXkK/iO1PzBEZDMscvMf8jz86gMTlzFq3nsL7H
szdRtX5q0CJxhv8pv9JNO7mjyu/Db2NozJBLq8a4Hov7Qz30W1nlefWvL0jcEa56
KTMwjrfs+u1hrc1OG3EKXxxO0R1yOTr9H5dissjpHMsY52k1fTVrmy/0CjSGBs1e
HFsgozSlwDRawg6pSsc25gA0KeLshwJ3JQmOgDFAfmUZ7JEWEB8kEcLRD5SikqkV
38cKTJBWvuarxqF6/24u87nBnn1HG4suncHWnw4Opwgs8X/Hr9vrXvH83WAEq5vp
zkEWuFl/RWRGNYIFt9MXE4f0tWJ4EKj2Mqf5D40k9n+8F4KUfnG6fIxt+p7Jhjay
Zcr/1Rv1cKRk9S5wi10uMtF3aYNjhfRy+08F51BilxXpt7R6C4qZXUzfGEDP+ADg
FEea40W9rqOlO4/SUGZl+LkPXyxjlbuCX+QCASv3IdV6H17vQsXV3C9VWHVUylQB
8e/TBynJbySmRTDhrkuDTPIyN0CM/hRuQFJOFvRPNzmbHfyVTX9ldC7KTEVMEd/G
du/LfQCzW5Yvxx+Beq/zqiXMKvxTFrgTiZ+GgopIfxJSiA0geNW9NjM1N+DqNr5K
imXrvVtTUAIavedX5pd3FpDGB+QwZr1j0J7UPKu/qd4yTog6MVubD5FWibOFIvKM
EMQErs1bYvZBgEO216lcPmBDkuuEEqxt29Qi0D5oCvDm6irGNUR0bMU7g+zGZeX8
Ok8a3wGmYSKFc7O0KRd55fLNfiKBhKk3fMe52cq0ERKfcUZ/roxHKhHywhNC/oxF
54uhfoGDS2fjuZDo8NDTWa1oJ/+GhMjniFzbfVDOx7Ik29h/OgUOnk7ATKVjqaZ2
31OBo5NBXEscum/jgTuSZXzbUKPKf+2hONVx7BhlbMHTLa8HeOQF/rqHpB/exi2k
s0YZvkmbG0wQg8aojPsnYeqK6/3uCE0TPv+j1SGdEZdkMFKu8GE27Lu9rWuQja2y
0NCy2rmOJMo+Ndsks53UsAV5Z+RRZkscXrvO9lLWhWvmL1fad64XsJ0QuNFmGWMH
U6EvWombqkLfauShVs/IWI7ktGkMAOjG63TwSNsWH4Lep54omXhnVHAVr48em4SC
he4MEnq9tnRglLdBYyvgZMTEc4V8b1SS6qgmmSIbHTCrEHmJz/9t0V9ahsja9m1p
y1W/gpOUuQhhKvLgpIb1GWeRn1KZnXwZD85Pa6XmsLuMyUmf9vhFGmNf4ZddFqSm
qPU1nTsJsmCsjseV1DumHY5SSlB6Zc/lbKwhw/LLxpkiDBnOxi+G6m+/uHzppAiP
63NW0QNVD8LNEoqBRg4AMcPHzid+9PRURVUNbk/8WjDtWE71TGgYdAknLnnsCqug
ILiYFbHYzgLtF2OX6Vd0MSsN4AgnQkgzVL4bauH5QLcejzIyYpRHthD/UZiCSwld
7okOyOW5LQZaNCgzuEK0qNA01U7Xi/VAZNtzJFQ7VALEtZ8BtoDqjViUU8SgxeQc
aFNw5HLQef7K34ONcZq38E8bxq/lG+DRiWg1tpCqzQ+x4P+M0y6IVtG+K39M2brw
SghPNH85KqQxfAqkRNCdBO/nmGuQRo0gBAq27d6jPNZRHM4QSz7OqhygyYDnm+7+
63OpSdRaY/ce6s6LqwdYiKjSIxPUOvyzMDiNnQ2bQ/mIHdx1fYNdjB7P7WxC8Czc
uMRkpwQpJLW400AHYpSWte6yD3GUY76uSXu+ybhWfiAKpGIEaGkaayCd24u/gSn2
8KuCpB88rjlZokMfEx4BqE1mRikXLUY517n8ZlOwh4VTvPXQqOjj4u0dtksY2/+V
5OBxI5fg2vMigoJewb0vc+Py7GfwwLplKmBlmv9mmoMGccrkRVsIQnpjqjHNotv4
ZfeyguRA0F6gNl9dibnyUMzu0gyHb3sX51xs0oi4hBPw/h1RC72z5jaVsHL+AY4K
y5blj91ia1vhA1Te/u3oojNXhH59RaaiZgdcHDZx7aINdfVm+drjezq5f1/flZRg
xRgBFsNIw2dONY6zPJjT2AMaM0rJXSwa3ADIe4CVKOUOl4z0n+AnevYvxW1emNUx
ObyVkWvWBcZl4iIeuZZLTQh36Tm7+4RHqu7VjrjTNCWmvzCDhwzOXG2yzDhucHyi
qSj/DZvPpVF1f6uFXzk0yZQR/Eq9DoskzEeLOzdNIQg9kW+MkEp8ah/pjfwjTHaJ
4AYTuW5er9Mto+NVyUdTS+7KypBXBmVomhg0JYpL3H3fsCs8QWmG3QRdUyFfVKYy
TvlV06zqKoDEEsiW/2x/SmTMahXfDxbCW+rdWEf18rc9PCVpletz7gb4gBXJrKKH
qeNJPHV74C5JDG9Xc7z5hStpddhrkXJ3j5kV656MNUaNoG/ErhudrxndfUxnM6bm
OgiiwY+nrBRLMbOgHEVzcQd4VhffaUlWpZUfgmylGTh301mCxHKZ/ORLGeIkP/O+
Z0YCrILBhis863cWPuTL5uVXLg2wgJ/si6JVLZghRvea71+senlGdy8TQ8D8tao5
4Ssx27J0wlJ0y5l1kptcRb4GBpytJ0tCaPB7rzSHiU0cbnFzcnCUnqhlybtgqMKS
M1MZKeMPCNbkVkI0zFJOMtnQyQbBd272bXW4EXz7Log61uuAKXS1I7AUEzX2g3No
jrpqBmo4zut5xgtaorH8yO5L14rkaCSBYPFDEo6R+W+5iakIa6k8HUJavcHm2QKW
SDN68SNV1zaD7f58wK/fvaJ2UA3x0Y35Eh82j0DDjJ4p7OcYip8NxKoDXRcMzBWB
DAB1lQ+iammvSYMcWCZrbWi3fSNEYMpFmBGlo00odTuE7BNgWF2cG64b8A16bqP8
3JckzM0XaHwZdsMwLiFWYe0CmvJddGceJ/FZq64wX3/US+2VnK5hGMyqNTVpg+D9
G8n5piMpMBR4AR/awdhaNc9E8HtkCUrztSrvNvfKtTR0HDWpRQYmHTmobXUY+4s3
iqQUVNKQIq6OkkwIUt24qrfLXd/hzZIZ0UJ+gC+YNOpdxjCWjZuyP9gjkyysKEI9
QCsreukt/2AmSM7za2oFGfR5LWw+MkVTcBCFSqSgypzupRzPN94b8aEz6AoGAQOR
Jz5iAFRvrb7z9nUHN+tL3dVTnvK3QCjz2zr+9Et3fa43UoFwXDlxy/myJNEFhvSS
zXx+IvFpBQLQYlL55xtoe+gqlPd4EeGp5MqO5YVUuZPzCLwpVoILZB18isrecFnR
inLsEiYLQmoBjLADTvBbIUh94RaAq+7QtDX9YqOYGJDm2pj9Q1DT6QrcyBqRjO1f
oXF8EPruHI6eYq6lzN4H0ElkK7VEaB1JlvZ4MpsYzerEzZ1xO9kuqeDN43bwAWqw
8heV2IZHSwqKFwSPqGoyVRU3DfsM3eTdE41iyZNc1xlewrgPyyEG3to1UnVJwvaO
5lCLe5G9QpEYXjq9FoxIGadkAEFhbWF3jPkCu/PCJdlpNrMoJvII1IXm78Wwp4xw
FyAI0MFb3+k2udrV+LPblTUl/2SNOsHA1bckbMsB46kK0tgO6vEgKtYaqvBn+10h
I0czMBFUX3SnXV/M9goLKHMqBw2LV3PcTahg1eWh7CXxSM4dIOuiYXFhzxqDrRIt
ihCuhzHnHiFPkbBJHfpwJuqU1EwSvMPUK74IBJvdQhC5NUWiAZ4GWXmSqHiqdEx/
tjJh2WWodq+G937IQdgwYT8+leCGFeS8Jhy0bFL7XVKnoieIkT8h6A1JLNGXTtCI
cvwGQpjvdDhxQxDfb/yoJU3w/zFRl2/wx0xYbiUVkwgKtf2BlHWpl4NbwvcWzmP1
q8vTng3sIOiocYO6Hd7BTnP2MSXbUMqd/PUQIXWkMQLi1WHmmR3G8zSClH1OMedU
XXeJTGflYunCCaAdOe8U655f924oYT565AWy5hZtv11JxlETGHgqFGayYDUO3Xbk
5AVbl0HhfSI/+UgInwwIS/bdXxkoxMiHAPFTRxthDpavBa7NYvfIM0Y60q6IywWC
EpNyrS10EnZk3GG6o49U8JpqKV6Lukat64NzDt2nyb7+c27pMAZsARY+lv4MPI/9
mfOjeVbqCygYhVoZ1NZjatb09cohC4EL9nm1u/fqfEtZ7Q7Rv+J9gpTAIXLu7laS
YYeDeoJZzP4z2k+01OuX6GWnhbygTvWawAZQZyvlvMwzd3AFPFcGZ79dAHIjr984
dvV4q4x2YiDWjPX39Aexal3rVYaD7wtAc7akDD8SEu4plRspnNdzj01BlGpimtQv
ugns51YMeXEyA6FTZ9lq+5TF4O5zEoe/1wuZTw3Vwgcrw3nRA/j1hLDJoCRkK0If
HdaEQNpgdlznblvcGWwlFclqykzSKehSkSoHgVkjE4tZdSQiUC0t5RSeLZvxHDZU
myBOfxw6FEX8fVFYvwmlijK5FcweLsnncfTcrepQTj5T9zTUecpf67MTal2iNUOd
J3YDHzbRu0JeeliMdYFTkLRGRAGGSzKbsVRWt8l/gk+5/0z7gD6Z7t4uiGmYy3Bm
cFpOhSaPToNRdWEtl0s9vzC7ZKfINbAtxshwFN5MT28wGAKZ07Ot41cxQNK5/5VU
l2H39sF3OY89jdDCLBbRyxcOqy7GVWSNz4AQA7SRk/zigiX3cPANib4+ZKMWuigJ
cLCf4DLxA7Rd0kaLiqB/e7LrTP/6gOcvsjde6tJAUPAoigDnJyqHeEclOqu+Cdll
YQdk3XDr49StSPrNVgN3SB55WBOy84Faf01Ox6pzxF5wNTyd99LWgmlxseCG49Bo
0/FpA4ew+LtvffKksRPL1JbJ2PAyxaYTmirxQFm1MdWgmnyEnAWBFVT/3BRAz8Ov
4316NwJvEu6WFlT4v859+oOHXeIGoRhNpAKNfLRonmh/gfpYqjZehroiflAna2cM
cKN87rKNwFOdtEDgfDL15o360EEleKv/L+M9mARCPGqZEBZ8LV0T1lFQby64+xmr
eIhMJ/D5EUKBEot3AA/5UNMtnQ87SaXixChWxvron19aykONgbym9/1eBZ28iDIr
3Nuk6M5tuFVIM+EFJErwRTJbxViXFkXjPhC4o+nkhKUULDxR4REuL5SrYMZ8DFXZ
9ZKd3g+x8ob8c6oaHoGo0B+sfM4/QUPsdkF6wzBVUZMvbXa+IKbTpZdZQAa3czWM
huOUiasHpnj+PqNX3boxaL83AqnWFuSWtGBjcJgJEov7KDs2sboL8ZlX4GbwT2VJ
6UBxQVF1W6IW3YiODr7WQ4RGTJ7FFaXWFoil+CCQRRD+eiH3DIAK9xRq8FDTTSTj
j1bVO/pVPcWvASoASfm6EwA2SNBzO0Cbce03x4eysvVq92RdHRaxp/Yy0i5LhlEb
fCENnE6jRB50ngRh/i+2BRXLkKe1Nwq8sWVARUDQsRRfswGEaLTq9IIKJrzaRZ3b
FZvvHNFhKyuQ2/qyw/7bMp0PV0D/BcJGypzHFgC4JVRjzFdyVKHt4SNOwlavR+hg
rYcoD9XItwyOkNvGXxjG8+wfQH4xjSa0dKZQPhQmlxMm6i1Hw9VDX8+gpNj+UMLI
/CiXYIhqOrsj/W3aDdg6iepFX6vg7MEoYFDF4up7cnya4v0r7RhWjyHPFQwncUXI
eh1uB5iQwqY4+BfdZxTgRmFbWp3i+9BI0BUl3E3BMbZSXNrX7E3llcgOHdqhcPre
EMy3K3dIOLLTrB6oUCG50Wt/Bg6ggPRPYPT+KgGOZk47HQWVyestH5fXYVsqgKeO
FmoquGI2kt9r9ue5sqVQvjDfAiBw4+CpCYQKVptiWpFK4xUoZTcim4c4umSDkrLo
byVuJF6TEmnAdYdI8uOSW0pnV1jJOyax56XJuUXb9OyJRdPqYrQZU6Udhutw/3we
6SqivDRubNiJBPBeFDmzWqXY2EVvC4Hx1xAEQRehTMj6salR0NUiUL0QofQC8mH9
zkoZKVp6H7rTHJYFwwL6oRZT+Jm4w/xd+yhb2IGYgnob5xQPyOHFCS1baEJvPOxr
agP8YADb5yHPrTYG4B3HRsMK9psZgKL/Uyq8mmyDIgIq/N3TgDpkY4b5DK854lT1
jYn/3h8ZqwXANKzxXUAdsyv3uXHkPFMtp+rLIqqK63UaX3xlg/rYTzTaom2nTh6L
3RUxWY6IQ+VXNKh+2CJJFCdkdAnjUIl9+0pLGtSsaqORqnHz+RVpqZf/K0ef6hjw
IKWwcxdo/Uxq+8LgkRzIjqFStQWaYkaEOR3ZkxvYsQKHwcWAFNAW80SGfHJvdHSb
VCnZDy+79VbrqHjP3s7Y3jjOuauPvyzB1nScRBCo1lDfnUQcG6re9bQeh/MqcGR3
BPEDvLab3QsG0OpYCecXaSMD/eUtC0TwgSIiuUHnjRwoAGnIWeXAnazbpvGAFLWA
XNtLlhuM12j8fYuTlapvp2RZR0qxnJNfQNv49M83xY2j6ZjzcHBMd814UHsOi1St
cujpKKSXOtVJRKrqn6U0SWUO3WtsKTEGPgSmOpRLqoeC/e0oL628HuSd0ntgKECg
gdRTVdkfH+ta6ZCyXPursW2C0HcaNxrZLyo+P0vnSepBZ5Vap2xE1XJPVYjDBLDU
330RtllV2v6qYxWMVI1Uz1w089gwqLJQH5HS1+M7AQvcpNNTRk9UgCMlXAqj7YQd
dgrinUiEzL7QSlVMaWPgFK7p6f1W9qIdTHaKIhaUh6F+iN+T2yyyxgAn+7nHptdg
8vwaKy8Yx4qnhPREPdCs88r6urI8ai9Pk1tVEksv3IuE004vbPFUUxOaRnKRF5Ey
Yl7Khqvy7HYDxhs/vwePkJCNSbEGBJ4rsWmFBJudtCzDHvGa+Ps05P8z58qAKc3t
Llc2A75metlqf1cj8NuPqhkMGZVAA6Vx7pA/V11PIbZzBK/72jqKSQJVKyilyhLq
oQScSOYDN6GYANabkQDN0Daif2ex7k9G85a0vcCWYFwFI6l6q+0BpORSVA/pdEbH
ghcMbyMDgNMkSHtkmUApsEQb8r1s5MyIXcijyGjnHIg77/vdn2n2HQzTTFT3PBR3
fDQ+XkeD31fsEqzI7t7WGOkeiCzs1dl6a74GGxQ7NhLameN/7u0oI0mmylalnR8p
5nZzgeeqmDgM0jdgfYCggtm7iVPhtex3z4CYsq0J8s40+t5BIkfYIOGkJGQaRc/8
/ic4ceOxcYqEzn++tMc4EaGyCQChtsjhRB2w0O9Hphzck7pyerEO+LEt8DNI4ZU4
ulMvdbO04/Uh4AykWpuKqdsf3sbjKeTKNEqY3asl2tDK1CJsF3yZmNlnpGMN4R9c
maAxAM8D3MJQfPISkB3pCbbmYxgpijU1Ee44IYPV+ZRuoKSBROqMeMiWONuojSrm
ko7Zx9LgLsLqefFpOrAeEVEEESxrG/zR3LZ0Y603oGb1oAuwopdnwGSU/lyZhxAQ
kSv+Ss5hX06ivaBBOv2YFPlx4MNjCRtoGCxqIu4mLuSR+8kDO1ybC6QkICK1wqCq
qlQgEJCxJWD/g2TtuAB9Yc1W1ZS8FcbMq1hUs322rBTk2uBQUT4O/krfBos9QflH
I9/xfONirC7ex7rpJ9z2isRLuWMIzvC+urBlGnIK79U2RJwk/anObeqL8OTZ/fbt
bYXVMNZa5auvh4vgCGWsrWfea/KVeW1j9+deFrCpuqBziXK78B1h9JlsA6VxO/C8
EscXCAOXdtdYB4KQSK7he6mW0zmjknEByseFPtQa0PUJMC3C/Q5F3F24zQT1kINj
HdfOM2bvSqgA0z8IqbzLcczy60bCBmKcG9q26+DW+VObheGBpufOBMMUiP2P36m0
pE4Hldd740OAVCSx9FqD33lR4j+yqOCSXrI3glipNSEUWDhgjqGxWhd92wUcv/lu
oTB7AnlRbt0VVM7hN6A6JS0cm7j7nBhkpc1AQyOcEp54+GrTcZga3drS6/oW09pK
4bM5/Rc2Pusc3GPgRo325uUQaaf+8CxhSOkC6AjMvpUBfgNgxCfmD1VW9BLy2Ci+
4uDVLz2/ZJNS/+mRIIqczL9/Tqy0gIVJw1cmhIaH5+WtmgHq+QWcYmdBrGK38YvA
OfHnRDt68PS1w7/7k1t31Y8du1EEssjraooxt/YgEgJXD/wjqEQgIBmrLUG6MrpS
maJ3sJnqS67SP9+3lMzpOT2aPQMc3AYb2NsKRe/Ar4gz4KMXqFXwe+q038h3DL5D
fXvVux589CrArPBhbBVs9fnZCeF8TqSrgR76w7dwZ5iZTq0amKPJe/+LnwP5Ldcc
s5jsIlI0kYfGIUYAQ+QHNc1CFZbrHKbRS3tJ5MhS/D/hntwK5yvnQHJbKeObgzf6
BSWW3xsIN1kijmR+RtAOdl0VFD0j+Y28P8/d3i10KCTltxOkDU1C99EtRmfnNfij
yblGV+OQtmgtB+8TMS2tT47H23c88+Y4BKgfZS6JuN0TNir530B29kObtgSPJhPM
KIKwPY9asHVgrWyAudDDS+bFblwd1r5Ss0tFglojRZhb1DsCyTfoQfHxJFMxU4cs
VmvLXJLkhUngO+Cy2oCzZ14Yq/wlBCK5yE4vOoZIZKfDpGPaK/PVQDlfmpW4wKfz
O419JNUUU9azsLZun0DZ5k57YnE9iwvcZBxCA2mSiB0nHOipBYp9DhBOE7/+1azi
7FmQl7HkiF2lrHTTMH4JGNEgx538VhKvnpLF3qmFX9Ebqn6QM3+e/5lehfK/9Kzy
6OM4U+5NZIgoYVLcwHn3c0qdRKBOf7wVJZ/8FkgfOl4MMe7zSgGPXfDxxHPFXROD
ikIcoZmuvyclOrH33X+dKnRMqZKEWOBRkJEN+Rp9iK4GkMOO8hshqjJqXbMD7f+w
HQSWNnOF291RqRsFSh0j9t0KOKHZJVGIaSvhHUI9QsrW7S06KbT84sUyycwNI3x1
OgpQWsscTKB1owXN9FAbK4yjZiUNZ/LwyeK9biC5JBSOlTGEi1kZDvjdK3cT5LGR
bT1D2zNgMsNbhirN8TRS0yLRAd1W/cXy4xlReWWO3bgGr/9oC9skdK4QqN/KLSFn
c0Qb/z7NEHLFHNrKmvTAa9mIXP5Czh3la5+NEU+oZZAzEAP2lAaMgyE4nazsuQN3
+bavrpmPkzVd6X9ccHMpjyXvMlg47cIKa9vVg+60SmDCTuqohizJ7jG78Qm+f/xH
UJXduQVrpzG47dTzZdZQ9CtJxaif+hPJYvt+3JI49aMQ4/xbA0mbKIQsgo5lAR6F
8d8m63lnAeU6jApjILRSxrikDUWfEUIAXtmUv/KM5K4ZY+TzK4w/o6sG9cLrXRR0
vj6tuKDsK/7BbCGLlgDsrZfTlYcJw8hF1VqgQkDJpYYGmRb+3EjF1ofHKRcaAPA5
8Lmm7MlpTK8JyGHYXRhhdTFo0EafV5QzXDpDxDmwsANhMxbx6YAqPCr4Wtgfop4X
1NWeL6Wf2CdP8VezMspT6q6sXr0vcE/abAT+H7tjCAv96qFRU7w3MsGIxXt/ktkZ
RSGeBPoWIG5ydVMx40IGwLW2jayT62TWrbvS2NOrmOBRaPawtytGysCY3r34w+Pl
oqByTf+nzFEaF2WQRV2RGVm6Ab7bmntp3TfkjIn9UK9Swv/cNo6TWBFrd6eS2XAP
kg0dMvP4eFnTNo3ah+7czxEOMB/DzEi+tyNcy99f9Zq3gQiMQDj6ed0AIoPvAo5U
TudrOrocbuB7a1hvhy+q4JQaIVkOdU18BSBnkoK7DPdh//oVLlsmXDMtH5hQXWau
GT8KGv+BM5M9YWnsk50JW3fRS0Qx/bzaQb3LzsHeWIakKVtAfz417aK6P/KKa3Sx
bZgYzTDop/mySrdgScwMdBmKZ5lxZsWWCBUX+sMG47oLcn60kYH+gMNoB1KOJNUw
PZSmF49ty2UQm7+9kUTeqXnJciv2P4/VJ1tbt4EwAl+DG3f9bOrLGGbmqg4Lbf3A
/j+lUT4uDTT5kBO1RcnwBZhY1Vf40s5pTLdvxE2ly2QEjVojx4bFPidbEDHK465V
9a1/aHgWwLGuWfv/bOZRNfGRi3nWLwLI9sNlLmRAJW9n7QyMpBAWk+50rymtmzRd
pkxghOmnSpKgD/n3saH7a/ivVuxDSI8eiyrhU/qNhjpM+gt95RiFaFvOhfia4Bjy
UOofHXThKic+0YzP33gvRT/mwfxLF8sIyrgJsLh/Gc69mwGlAPPKymc87/6TcFpH
N3mH45+nGad/5juUCVDtNUYPdKYpGrz2Kg3BQbD8LXCMrih8GvIXDZiY9gcqeQvQ
M+1Z/+BDp2Mc3yhUkJ24pd3PX0gKPi/WIx16EyHw/lrBf5EOY81yEMC0IQg/2zuI
yr4R3axPy4ao9nZ2k1AYXZdbFfPhZSKWySNuFPm2pg/O42AL1g7lJPAShQgzPq5y
BjdD/bkK0BY510E8Qcvikwebxpl7pClGrObH20XPnV9Wn4JK0R0BKfNbrKkX9Cee
75Cz0kgUXEI3svm863buvp8tTCWY/l9pmP3/yKt47B+PnEsxIhPEdbnOagnDIW1g
fHl0gHrhprsbDbKQ1bgsZfnZ79l+SWsmh80/UzRdyTsul2ScIcE1229HwkdTz/VJ
y6hRF0at7o7OQhs//4rMrfLJ0wlfKHpqlsigmY7cUJmZjpm2H+1cA+GEbSZjc4Sd
E2FDTWsFU9GL+R0Kqpl1P3y8PZHeaxj+7eUC4xinjfERKpGp+/4Ir1xZsxpjNO6Z
5wUIZBayeb/HRgxGDkjV23FP1tffNwr4mdklwZlfUF9RRlaAYHRkFgTCJE1hT8ak
8UrwmVe3YZnPgYfueF4dq3HNMqhadtHoOy4CaQ859l/ZNTaznIAqTDSOrQI80a4n
kV60t812XgMxCK1UfNJ4j44Bij4jKGkAkza6m6n5ecsUb8aEWk7j28DYykuOoyN2
eYIEyyhCSgWy5PYQKHbfD/aZ/LfynEguwqnKu6oTBOrX9vGPZp5kZo2jP33GmdFO
VxQT/1R0xl0cpd1Y3BheKPOKwM4EU8Fyx5VP/UziLSO3Su1hIDJzhc03arfo7x7J
mN82K6iyjYMPjTvRmbpqFmCD9yad5WnlPu0DWSvxUai1F+ftBzJQWOdeSITWe0pU
1xjQjSjdr/vuHBlYSNdxI3rSdF9u2oQMSmBZ1pjwnZnJMknkwBrukEpEjTaTP/hW
FTU5KYM/irNJa9FhEqc08I0mqFThq1U2sfji5LY8HI/bJ23mJB9Wsz+WF1T6Su0E
L85iaUrxwiABldTcLn5vi+cedjYdy97p3xx07b/xZPI=
`protect END_PROTECTED
