`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYDGf/YtEjNUQq0jVVY3DZU2hf5eFi4s1HFnMqitS3UbAZ1rgzfJ1Jo30l0kAOHi
/xXka5MwOHr+wU2mC0YtVD89RbqU8gb6X08JGXoR+XunZx2BA7XHkiiztMAsQ5K+
MPE/nluVRFWkYY2kg3HOrsZkWinrZ03kghSOlc6wZnh5G9ziNGWWhQaZF+LNDZb2
ezMvnfIhMv6iu1259TJhc5kJ6x7v94YT7SARRuJth6Y8EovE27zIfLSqnSffXOkp
88Bl5+T9izwnHRI47NAKWy9H0XczMZng5XcamiqNIHoocaidx+fFfZH6uWHxEKWX
/xG24lB5sXXMzCgzXREHH2e1eM7tgzte0UMe7njTv+cKN09pM3yYLKSpj2qNQQtF
wjqciRdq4Ox/6K5yv0irBRAOHP72xE6xMsnG8mRqib1nl0Oqx1aNv4IigxrgfYiN
lIi+iWowDHlpu6ZDCttp/zVgPE1ifLNZmBtHoQR992kirxqP6hWghcoMCr9oFMX1
zxX4jhsUaL5+G3U7IJ/SiSUqvU+vX5MJzPkpWGgodUebDro8HJxt6AY5tuJcQC+n
yXgu8urXOLIJdnkY39rw4M5My1GnQdI+KX3bJlMxvrkbBlJ3Vrn0btXyp3BFBDxl
ep+/1Mpn6v7zm6PYSMuJWZkbfT/H01oEqzMeXHBx7mhDhX8mB0ACbwG0ylMEltKN
HmtBG9rjmHwNWoaUBqRvf5UvywLkKOKG5WdUCt3XxlT2rM/dU1ioZ5M+y+kTZGqR
YGvkyBT9w6dKlfdlQpizq3gdbOwZBd6MXjSSYWHrAEuH4q6ugpzlbf8gx+2IF9sz
RZ6i0S0LKSme1WD9GxPzWucAMw9tzXy+/F6+dOFGAgGFF+FKZbHRLXffCeZ79uC0
ab+TEfPuFfQfRHnN4oavdTjU2zQK1h7nwBdUr8zmjiysdDxqZ2FQXbh9nJBRs89+
60hciCVpqE8IPwH3pxr0xQlT1SOpcDQNnwN/6yg7KAklqSc3AlP1UrCfguPiVfn+
Lah1cb5kr9OFgf94Ak3RMMskkAzTLz3jDLLU1gD16APPUC173dBPSeOm83xu4M00
nLfTXXeUu5y8KYzq9ppaWhpGwFnwpJCYpTikkRWRAUAen/ubPpUO+tFEqfqGdNdI
HyC3fNw9lq5PA21yTgEhJy2ysxt5dFldrFLVSCH5iVSTxZ7YGTQlmMjQbLd9h1vI
FwNs0/wwcyutEzrw2nxba6ti0xU+f8fxsc8hsI/9GscxR89QYOvMwkEIn0AfTA5u
M+HwRpF6j7RUfSjte9fjBJ6AtoKiO6M4vi2YbX09ghbi49b3QAcUF8gI3wkfwIKz
kgIzcnmqMG8oI6HfbBKQ3bWrTlrN3o0p1/rFbV9r59yR8fmUCBXCGXE+p5O6nwvI
6V2/f7k1JkAY335cCCAWTE0t6ZW5lpRL+lhhX7NT0OVEyWvuxgLTCRrY3M2tQBPf
clNlr4MHvK6/7r4IL2RzhPCIDqJit3BJZ638kcqHGhVZadg5nBMN+Dg06ewGQGJW
k4dc6Q2jBSNUwoxwyt9J4W/SiFhlxv2L0OGfrt0MYYoqwvNWcCMwYAV9Ji9EQp7h
Y7HVU1poQM/Qt0QY6FPeIfvjgFc17uiK1OBM6Ujq6kCZ7cgOiPEDV6m8tEN2xo9X
s8U6Wk76q1Sc9AyPTP+pKqH7jITG2eLlzxtrFcqlwsdFGi+e5vRYa5TvTw89EnVE
SkAW+L7ssOtH5eYnbXOoNmr7uZceLggRrUbmVWMZGPknqFj6OmfIVicJGewIwA/9
Abi2aeM8l2ikwU+udBwr2H5wc08iXHV6ngmFTVX2uFDMTKByAgiwBxBVytQsJjV1
zvcmWPokHVfb25Bvc9Y1AhgPQ1+H9Djb+ztbvGjjK8TJAThL/ZiJ+Z4bGaNvkRed
EgUXYOr07jlaVpz4NwtV5VwNK2ixQkZmUMpD6PViZ1UrgDXeqn+L4rRqyItCrQVv
dzq5b5Y9NW6ECWR6Q8Y9xhAk2M76sNR4t9iYWxk2QqpA7BaiG1u0M6VlccEKSrHh
zqkmX/cz3JfakWwzz2NAyCkDbeBZ4+OlQYe/DxggP3YRWZURzDDGpK/P0F9vk/7Y
KnM1XNZidQ5YVR0mNXE1/fSEVOEV9A2hHw41tCdNU5L5/JRxYcutL75Cc8oAG+zS
32QBfdFYnpXYEVUN7iEvE++/24TBiVBT0cUGz59wVAFN23PsP6ExEzITCxGTxDPA
j6zJ1LHa2uuFa/qkci+z3Qs2wR3EF4PFHBeEq3FpT4ILHYw7h6DD+0sHIX1Gw7YA
ndF0el+WeOwi4yk5eXpgmotATqraY+JODwcRDnqyiJZZVAmYw5oQXvvjUCmLhkjr
mvpyuFWogSPQcZGGQIGoqyNjM+NgyBvfjprae0gJdBANF6nhSCiCLezhFdk20gND
kWxIrN8jo3mIGw0LuyFu7SOULfIqoma2rL+g9yO55al+soIQBQYLeASXbOnMJQZl
UEi6dxL5zy5p1XqaOpTTYpXAZFBVyqy+1PvIM2W6ewUFbfW9KKW5rFXjJeo7EJzK
GjVl0/6E4lQ+5UUrqsf+lmwDsrVOP4vei/289J+6Mlc=
`protect END_PROTECTED
