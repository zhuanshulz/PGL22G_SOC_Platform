`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8psuD+qP3uvPK0yLkBnnDJpf9jyVJ8iWjJ3wo9HdI5pSF4QpkD/BrhdaGhcH+H4
vZoaKt/yqUGEZd9snIVc6x8ibO+mPECNrzypUy3IXWi1xIfhIIOPvIR0CjXJS1bL
YZgJk0ZWpcgOnyCl6qbT/2ou7XkKQ5//esKf/OOqOFOt+h1ZZSgWFdG2oUxdMhPh
DCyFmbwwdEA86UtZqLn/d2Z5T1V2y+E0pkjdwBvD/zt6GK4rpbXSKGh4lpHBi2mi
AgrePK5J8UWy2eKihw9tG4c4DpI9Y1iigUdLidvtMgMcIa9xnWRHgP59wlNPAxkD
KkSGsjBfe7CsHcVK+Cabg6tIITIBaKk6t6WJzA4eehtoncJAbSU3D9o4h/z5OF5y
aYzqW3qWiCzGs614UFWSNJF1E+MwI1IvBLXUEbvCMZF9ro3tUPLmOMAczYueEQcY
kg+G/6bhI9moPMDUKn1HkiGMA+vChGUmOLxHSg6D/iITe5Hl8MLV2JW06Vlmiox1
mx9RWAr9qrqIvfWYwOv/q8CCiNgWKcyiKlpQzrQ2qkzlnPG9P/vf3bm77/cijD6h
UorfeJd/oNfB6HS9ge9gGcBzFkA5hU2VJwAobr7KALahbJ8qmpipO8pRAyqqvkg4
FFfjScHhhNdTaMkCLeKfE7/0FfnHzesdqtGeMoLPxH1q07NBBAt4GnJwYK8MLAJB
56dcrSHK1HOGibOxfTFz3ycPKlNFQa2x/0t1+/JFNuw=
`protect END_PROTECTED
