`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICvRdkyNr/q9pzNjPBscxNTSH9kqZR2vffAAGtijf7AXBrLvTdXJFh7UXVZ3J/JF
2NDV6qp5jJGR6HiHxJFDnXpci9BboljiYWLjvaygeDu5+erZLSq1E4GP3Hm+bS70
seL6AqX0yNk6jWRVxW4+r8y96drzfTKWzQewFfMFPqUZt2W1gcm4qWwldIGxHUMw
cJNh8tAXVI8CMs9v8IFGGaKT7ew92N27cQc5r+0BRaSTFJqlCnTa0tWdEs85dUkb
mDs3RxDDk6R4L2FbjgGed1V1JICn+UJ29XKP6eJSwYFjOfHQzC1BXXF7nUjMt66p
8UaDtBt20kbcOLi3SXxpfQ==
`protect END_PROTECTED
