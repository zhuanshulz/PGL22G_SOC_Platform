`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxw52eB1SxYlHuTYBUvEx7iTvoKuRp9GassK3HmO9pGW0McxdGzQ571oT3BGpwri
//ieSsKjP0CI4HiBTNg4tW/uSFrlnQIWKJnY8Di5Fx38vZnZvke9BamwWGI3+fST
cywUDZ1/eZvDqryj0+rwTTWdX7J6ggNmpJx+z5BbB8/m6rBTXJdfpO+r8pwPFyUA
TQBjQyC0Ph+zqo9/1ogaz2ClguHM9FTj3bkYI6Ljhbthr5OQM+lPtthsvLAkwAtg
MkE6Zg2WdmUUgh4BVnMZuGObdujB/EqGuf/s1JLbjE6YSGskvqFds2U3TCiItJPT
2rHHFPlVBC5G/t75Nc1uk89gNc3zhTbvxCtV3l2bVfHpccxpnZaHGV70S92xRghE
kU/C3LytDB4dzgVclJPl5WVEZfSFp7XxxwJo0HAEmYzdBA8+U2diyCPU0dgkCiuH
ypFFYMXFc+WSv1r/qi+6kGsw8Ctq4wxbOcyFngUXHCQrZ+rzJH652OX6fngykBW+
J8Idi736F+d/+9+k+YZ/4aQXwYmxxuKkotZ9Or6PO9+JVexcEStRcRhSTSD+k74Q
mL616me7Z5Dvui6tqiaoTzL8b4lQ4WwNCUEP8BiHkH0UcgUM3EGfb1sYDZr/Trrs
WORV/16iRJYsdTQwMQ+2qb6kZw21FoJvwEB3htW2wihmwYvgDZ8hKUn0F+R7zLC/
r5acNcl+DFuHwoFmj9+qTpEvgnrCZB4RPpKOCPOouspcie4Lw3Rzd4QVIvGAehxh
wJ2O0sDSVVi500Y50GLnDrwtiJ74xYbG43K570lcY1ZtCtXcyGzoK2f2Lbr85pZ6
2VoWEbVKJ5fT871aqScKrbphAaHxfzjHGJbExzGfscTsnEhhDSS5M9QsWf+V8oWh
1zKLAYI28fd3QXD5GV69LsUiSmE0J37yPH0M3X3mbIir/oDffvA6PNWpKzyi+Riy
x3T4JKSz3gfnW33mXLbajrviNKSXZ/8C/kKy59/Kc0PPhrbBX8B6TCFLgzNW+aAt
HPktWT3fXlqCowvtTVzI/BEe//vQwMPzsas7/kRt1UbE6ezgx4maTKtmX4bGOA7g
HdWpOc157j3M1XUnHPy6ahJGgLxwW/F78GmG8Qq/mzC9NsmN9kJ4jbFNpHUEAbJ1
hyCZQv6ff+X/AvgngMgmm/Zm38v5Lk07lVQBAuYhF66cv36jF98noo/Sxby4UAbz
cvyrXo0A43aHgv9aibCpgIDkRdi9ZOVElN3zADoZ77mVL8FxgTgE61htByUa0RTj
afKhLSD/70Ah1XjCaDGNc+NjNrxBFHQq4JuK3sOiy0U8J8Wz/Gr6yee46PoslSTm
lwDFcUsPtoJUrgOO2hWhlvvTXy7AzFWDCAoVqta7Ps+3h34ZxD+gIKlVaubkiL4x
f8GEc8tGi8H4KU8TcCTJUWA1/OBW7VCuu0zMAUtgbOMWsBHBftW9fQxp1cL/8Ikv
vZtD5a5tFPZFvSKbXnhWD6EbXhuRoVlzX2A7Eu5xyb+cwhpl0R0ZLhPIvct70eja
k7UFgnGt9zToPVS9JZk/nfGbT6ZbcADMwnAfczY0lDtHWNgMGBBsx5IYZjeXs0Sb
zC4KbINmCmBG1MJFnyx7pzHxzw2Bl2+KQJR/FcFCWyK6cohHvBf2A5i4OGP1hYwX
smRr6si9x5k/kbIIItWzaDSufM191Zepx1/OsAa1GhEv2lUJLB4p7gUffe+c1YPT
O81kD/vHzP7zUWjcjNJLs6buL4Kwj3T1H7Zl81GGYl4cwumL9U4SS01BpSmadswh
9QldlPwqRnK0hj6XJTC1t2TXn0thEXtstyMiMylHQNMrQD+V9IU/XdeAPQg0VtXA
qn48YmfrJQS49132qIWvtU4A+n1BNEx+GuIH5aHyv8PxOF0H7V/T95ahK0+HbaBk
gBkRu25np1tybKxfAESv/AYSkPqGk/drt+FRnr6pOXGWlXEgBoSfCEJDUR83FgCi
dir7Sx/wCDYy8Fu+xw5iJ1gw+t7r8pKS/pbKi8TS5RQFXO0ZJGaE/Du4NoiGFaLl
yAUg9N1oiK2g+t9buNuS4XOYnME8w1gsJQEPJubePgt8/7OvMpM+nZXPfnet3LyC
nHu+zgbaCefbtWktl6X3BcdRRk+O8p9VhCNTASBjRa7oujDaiOZ994WtVP09MH1H
sQaMKsjQNdI1YmT9pkpZTiGQM6hOS9KCUyQlnqJe0Cf0Xzh7Dp7PJ+v8ozGRX9Mi
z8FGpDzVwIHqgx97qBno/RBKf+yf2otPC5NNtzWaBfCxPFKShr23LOVHZoPWwfoy
y8crd2KhH1vWsEXwzjzjVxJqpdz/BmrsEUKOqZki0t+lcCDqTlWUuZWAEssUyLhx
megzGkyDDITAUMxHSqy+YafmO8jYulluM8LFNqY0yCw3Xu38H5ky1aRn6Fwprj06
OoGvH/Et3hxC+m3FPWfyD0VVHuHikKpFgUx27BJPdnL93AetiLtuiw+Cb8AsMHTG
BtjXUd+tb25md86m++HbxBFI1Uo5RtW/cXYelfJfi/ZoDMMxNWxpD9yOGx33XEMa
FpBPE923p5Vuw7loz4jHySIdQncdJ1rH3IhOTmrIx5O1tBQG2uBXeD8HLzyru2qO
FItX7LrrkZ8rgl4Y0v2WZ+9PSZH4Qd4uuuJqsq2QTqOUcT5h5Tk3fOgZQc+jkWqK
Z5ExyAVmoIkxoMLjmdKTsZaPnBtHPGGf5o5HtHiGnEecOIUl8eY+N3RfzCBzpMIw
UwY0QKDaBOjEokXPzX/OE4CzwzYkA4xpkEFeLIwRqP6sQ2+sYOT8SX9X5SrFyAvx
RyKwlRBPwodPq7Ybb8SKJKA32D2BXCJ//M6hneBoaGd/B1SuDoyie8a3IahZadAp
Pyir2KE/2lxSt4znAguM/uNn7ewG0f7QUcM6ff2DXbYzRRy7m+9hjXPDNWkt5WI9
UvmXaaa9yxuFoz3PjTCsXNBz7sokTosCQf6uGeQbcnsVEuapkiiNbps/tgtNg3Ra
aNnf24F0n4jbBGi2WkGQPv2SO9yuJSKz3+CHSmiwt5wRg0XBu/HiY2rk1oJFZdZr
A6DJVo6RvK4CLaztbkwg91o3zaY+HdcgSYrdfz1vF2yPKfRx3D9PRPAFBXkYOrmr
GKtaAHO3+C1oufCya2MWNZjXo33n4pNW9TdVszdsDo33QXWUeH+Z7SsKBVDPDQXx
t1ywugyRrYyl+GTzHZZ6U2OGzrXWGpDz9xStrNL0IGEBGVTRKSSuT9GMqA9NNo/y
VeZznXpwF9R7b1rp68h1OXHadrH0XWGnvR1qVP/7n9Z1f11e2fZkoCrQdYEntk9M
qIQVBlQFNLvRq3thxgFtpv1g4sMqRxlm2lhQelGmW6i4tJx014oP9fg1TaaADicq
GtUf+gK00Lki1bhGlREJaBIofzSsXIbQulRS16TTSZqtNhsMPtMtPSnp1PAB8wDA
H2dARJgeEDAgMmOYIaniBeqeJJ3Hm+72SOC5V+2gIceoOhAFbSi2qcy50UHb3n6S
qpcopnvP8tlZKoNRXE7jfez17rCWDgNe1YLXN8BB0tZWzU4DnlMMay2i+uOx34PZ
WwaQM2oCZjAlzRYOwvHo9j5Q7lgIaNbGwzqMnDRRvmdTtGUK/Rv7pDGwO0kSpd1I
KqXxVB1C3oaFaPl35Enr80k1cIiLsfcuPwGmh+6gS7j04aE4LUoPalFGiwqSuM4W
IGqr535OlIIpaSR+RZqyHcqGAuFE+diBrG/kUGDk4iIGdSWD6QhBIkRoJV3yi5/G
l0bDdKHJ2jcQvdSHCuYSnESzZwZaJauHCWHDdVUGQpIH58EZx1w+/rVp3dAHY9o3
fcnVrC9zQbI0pMv3QCAbraaQEa1MXOLG/oQx33kGYmlY4LZzIXfNY6tj7VspChMG
RLsYmp/wp3MakLpegMzRBVfYV/iG467klF2237gmdREWYokmyL4bi2aWrdU2AiyG
6R6gPpYvwJpdziXXJ2Wv5WLRlJ4OAnWGgBGbZsvsZhFlhV8pDTcSbvaTuAlX9XUf
BqsDdQ3lOJIuxbTZE3TG+Z//1FCVZeFSRLT/nl9Q0u0eUO0sDAFk/TemBc4V+Zm5
7uqQCQpgfcrfm9oAw/Iz3njIap0nHEouQYXyv/ZYU22j1UXQuL032nFcygnPAtQR
AFYitDjxVN9Zr/e58ukSJ0lpHoU9xXTs7Wgm0DdOI8W5TaQKtjBq6SWDiiZ6V6MW
IbcZ4Dvg1wp+94VNbCasjK714OdbXASfzfJ9mLi4avtQ6R5mnfGvR6oZ97SI3m8t
U/VmFrApxSterdRdPvuir4ce++SL5CYfxoLGKYESLGoFi/e3Kgs4pzUpRU9oE2OR
L71oXY5CxT/IK5C4pKBlUnwUdlYEuORcCVw2XUep6LRVVT5Wmjzhezhe7hnfSX+4
ZDpzMpWg6v16bLqt2yWPLi9ZRvoobxlItPvY4WEuVIXpdHFCWPQMMDdAXLh/zv6D
/3q4SvhIiTeraHVx+KI0ZKNYoNUrFZ4JbyRvYkMxm1bjLrPC80iMPaUFCbf6nIC9
bdaPoUCpwrnEOuWo724vfiL5Eb11VrmQaThxdxXYR7VO6KenDfrPU0uVQcsW33yw
F2QWqvCaAp6UlAXFBrcZThAYPYBBoPTe14PLGuCzpJNBAg6IcWKtfoxUzi0I2K3Q
0uJTav/WKW26tvQknJiEXCqn8KHFta9JAHj4VZ5HCZSSccNNWCtRcWW1lR0B/lKZ
YfX/527gETvZ3EkJsKIGVVeebOHRsxLd4cntQX2Z/e1K621U+9QQJM5q6aTtXUnP
g2hI7B3hcFU/p09eSnujk210b7yTUhITPwiWQ4LECZpkO0NdWSEBTSYUxZlj6LRV
fQRydVTxphAiCD31MSDYqnjOiyH746L820+9gBn9MDUwvPG5YIXdfuI6gr/WaYjl
xsTcjBqf0TiaoZVuRIMIMkcu8xwBiDBt/tJOETYWFPWhlAT5hGk2b3mMhpGH6T3U
x7OMOT2AyyE66evZbG41sw+77GMThA8yFS3vcOqkDc5dHbDJmJ8aML+lZmOkLgzg
A5SKN8HcjAblE4ijiY4UwNRH+Plao1dTp4RAtxR58vbM8sJN6MM0WWFW3vKRbd/4
oib/lL5TCTw7qoMV0extyoEPlnVuQ4bPOcdK4K3CJQcdUcTfs3vc0bknxqwUJQox
Cre822HONyBTZAUTGm6dKGTF/3HGjT1RzUciUTw6h9DhXd2WuE2zQONOC/vxBLDF
56LwIhIyWp4O75wS4LYm46VOhcbyxVOiuF4dmHhDE2yfPKZ/rSJKmaX4Etsms234
tqRGeut5XtAkTeNFvmWZKFHxrrT98LduZSt6Z8w6o1CVp9+73nRDnMVriLpSSvQm
H7qY+n0u73cYTv5dW0UYhGE9iSkuoK4FZ4NLQ4nmJzG9rkc3Ll/IxiMIlQsm/xwB
+zZIBufURt04pdrisbwMVHd6bqeTPSCvFP+QukJPU8kcLHhxAW6YYnpan5RnScx4
d31EKpo3quBQEX6gqO5460U9cVR6/MzS5VMigNOs25bIzAjf0QNPAuICsE+saz9T
Z+l6UzXur1K/SOdjOoD4sodeUnvXsxfGvePLL53S4qX4wfjy89yCs2XMqNNDV2Te
F+SSp7k+3SyeR6mfr1f9HkCsa1K7RkcsxxgeflixJLYXDHgSvc9K85wFF2qETgOS
mv2j/WnTTb1/MhmCWDsufYq5trSguz4VAceeLlWNwTw8cj+2Ri+kTIvJE3ZaszV5
ZBJRJolQwCNGK8QYyKAZP8weeUhinuM8uqNn7NCUz802vNE3GtzJDkKkt2tmS25g
RJpk8tZmHcAlL6+Nb4h4z1lAB0WqF2dft4IK4+rCUy5tORGYZkw1wbiv1k4lmqui
nM2ghH5zlx1feehTREkT0FnEAPqF3DsFhNSRM0KO18CFD8MDXL2DVAnXJDvGN6tP
DHYQIp7DEWNtR8Jjp8QTAFjVPl361I+4cRHnkMC5iPf80h6ZAMO2TB2+Vs9ptIn6
fJidMkIdzetkNMo0OE329E784A8J9kw3lxnmrt5UvVl+9z7yWxR8quTlOtlPGZfD
xfl7OUhp39UsX7FX2yDRIaur0SFwRLZ5/hLt5N3P4ygI2FH6xeNQLXH5RVScD0N2
R0E6LA7xfcfB0wCErAo1Cli6nDxzLcOK0Ugb05h7Tk8n2INTLtzKBHm5m63rwluq
jgUqlH/yh5cordWToUGPsESyr0b13ItDYGJLIcXBVdVEvsDZ178y1xBzU6sDbgpP
+yJLB+5DVHQY17075cv5xQhErwCvfMzkXycr+1fAQKRf/6k9Mwv2kg3sGR76Ujap
gDbR0j029EKIypynG8/xoBvMu+P09dJ760/t5c19O6tM/E1YIZ3ncYbEPBxd+Nmf
lhiwRAuPa2xxGWROJm4Z3TXHNJz4IDgpYwCIFklQym4AE+lMir2y/eZ8G/4byLPq
FiRBU8jZ9H10IDC4RQTB8IW9PeGbTX3feHMdsLAW4ZPWM28Z6ZOJWyX/6cSHyB4n
8LB03yzLzDNTt0MhTMKBqbOIhEhX8MIB9zBcSiZt6l4xmJifzMj/n4uddqOqwEY3
E95lWqb5xciYIy0zzvwinfMTthM4FXv9EfNavEjKeCVdWwX+ona5uVXfPMctZhFk
l7WqiNQ5+Cn8NPQprDJgnQV8CsmGA0/1fwZn36sKXgu3GiYFyyO4eyN/YFyoJ+rm
EDPJjRQy48X0BRbRLnS6OJklcL6HYhfzedOmp9seyOhcv7Dq7zNzCrzEyj2Adz0B
YgslpXu8Y4RBfHGL9I2zN1cvXrRACgIq21R7RRiEQcViZxoHAzJ13Bs9MBHJHy3I
hl6qAMGk6+ijSyq8Ole1PCUtj3xJcH1FiVbujEcpOeYy86lpb4Czwz4xWsFDOjCG
nvttWZ9+bAClv9QNTk6XdlIIzjJg/XgZDN5t2nsu3XFKxJxcC8XTvyAju3NHCbFX
S1Mb6xddcOE6+euIbbS0mamhIl7B7LiNpvbGj5bA6RkZw7R3DzqJrHEzAzqbblLp
9BNjuZXYeomgsUVzjE/w/ZJY9Jnw2Ka2Tj12zFOEG7V9o35tnLy4rr1dzc3VxzXC
fWLpbxmsFbgSJKFWzvve7Xx4tuJQ3msslvnm/jCMUQ8tBf8yksf1JFOPB38VzU0S
VXB5z1+EhGBPbjE1alxzP4R5TFyHJckpHyGsj/ib65XOmHFhcHgugjq4YT/iM82h
mFXb1UO+NORdvIjNbUOEHjDE/G3G9KBaUyxbeVboIqQcCqLrCYs7rVF3yUS7sqqo
5K/y7Bkg/uCazBaSbPb8HihUTHsEmixaso/VCn8E1aUeWIvXwHuEIrwNAI+zGcL7
mvstcOxPoSAIaIG5hNc02M+bI6Pzzi2tgmLyyloS8oTubmZm9fg2qvubjEHAZtEK
qqTi+cUupc7ZHJxzS2hhIRVQkWYHlCaMyF1ASkULnC++m2Soe7e7g0ZVa54z+nbt
MuWVWsjmxiba7mfo7NjeUtE7dbqUey20qbDoySN5hh2Eddh9/0Zmm5CJPh3j+7jp
IFqSqOa9Apt9fjIiRrXh0hZsidSPNobdnJW7enEsRO9rE4RYIj0YORoSxKBDdOhF
Gw4sub9CJweT0vw4UW/kCcdOcA0Mba1KJpq+jB/crZvm0rkKCBKjPwjxjFT3yfyj
LHNCPoMat/tMijxHrOtktTRyFj4TFvAgl7I0Fjeg/ErLOLJBmMhS86CKgxTAWcNg
30/hfWEl8tdqPr0E4OdJl8T+RkMidabpBqqNLPHW5NpZvC2vXExxp+b2eUznvFIT
DqycRqA/AkJEWM1GNkEzYGUj4dtw3I2kXZLRglVvWHpcmxyfp4w6h8zoVEe9u+4X
nJQfmtTvP3E7YutNSBCvv0roLAPBkojFFZOA0eeW92MYwV3rBUPpvZOaiKju3Uj2
5zvL4nv2byrKPJq2IZy5sGtuz8yZYMImdO7WpY5BF3fhG8r16bD09rsY8vpFKIYv
+0HC2Dsr2LdL6lWyxxmUyZz2UzCcVQ/oNDUw6ce4kik0VF4QwN+gemZnlSQKrXAI
XnaMnmI/BHG+yU/ArESj0BRf/CqIMh6j8L3s1YFLdW4PTDkO0HhCGXZ682yFwPSB
IORP1Gv1XWlzy+59hVkI7A4Z4XOqUbuQkFL7u6nTjx18gLZW7cqVlNZwuBekshvG
tMhkLyp77AI7enMrGNATgkHSpiCTT5ngnRmTD13GaLZSUzfXpSnAkRTRKc/NuywT
/jL1DnkxEE2s5O0JfP/z8mG+zlGmnUrlqH3M3dz6PMKwo8NlrZGuvdyMAcBggjDj
2EMQgFX8uR7QxDfyLRTKW15xkiUkiKZM5rcy9RJ5dXFjigL2NocsnVmB8HiA4LfX
ut61MVafuY4JXCyS5U+CSLTK3cvDhf2krxAsPQGFdFbiGXDTBhbZgotlwnvuhNFp
TMGkRzdR+XreXkSY16YQHwbetY4xJjFRHzpDFBJug5aYMPPlNlyM4Rti+14Qz1Ud
WA+vXedmjEUZs2ZduvHbUgg25prgePddCEFvn5W85NsVHUEEDjMWUrAskNKNb6af
ZyplCwQNWwGU2rgf5a6otAw7tnyDIx5leMlxMT/sbQ7kAZq5u4MZ9nwzwF4NEfh3
QT/00rgrj1kEuSc6aYBKUPL7Z4qTpf6AuZQkhy9BiSmGJC+CnOELnD8mQl8mLGhm
g4xXbfj/wGQTn99n4mMVFGW+N9+u+GDSy3EWDd1dx6hNuAgAfxYGFYepl+nY8Z4k
+vuGdhH7jF8SsFKPYkpbjc5XkiSh1QVXRec+c+C7N1zkMr0WTzRqJnL/Q2kMF3lI
PFWJc0oE7mprBQ3WWiVsydFe8coPnWSwylT8iWolE2/tpbUTfxNL8YS/lvtLkXqi
8YCbai16/jNTIz8ARvy7Smqe5pocSW/v5KBLzBncw4mFFgmFjNgbOzdcY+B8wilI
3br336ndwuDlNu8dkFbGSPcjBLQkUti4Ougi/sJ4hJ9qLDW+bSndVs/X1tHTWwcX
ydZhPrLBg7AfLhC0Qm95KUWtoOVmZkUvGVrqrSul073s71t26etQFmC/9JCjYt+f
AEZ9Oz08op5HjSeelvy1/4PGwMfmz0jEVvMbjnzGpbp8U/IFHWRydvdDQTAa/39J
7g11H2Xh+G5VmmQzMXmCvffMABx93jt2fKE1dPu0Tf4E6iGL1RPE8E8CCt/0H8jx
tQWxxCL9lSzBxmpdwh2ht09xzwbJrmGPL93WgJ207VjW0iFQOCl6e+UQBCBwoxnh
0UME2C/vxOc3/gh+D9fTjoaYAzaRJAz2D5cLThzxeXDPG+x6yKeLQuF4UHAAyqD5
kinNkZq5lpt6DV5PhILoNgzYGrlLu0aVdsoZhRaUWontswPI6fkP07BvEmka7jmm
XZTg+bpJh0VGatF4rblwsJmFZ0Wks1WK2ms6cTSIGvzlGVfbIvmLfbYF3GK9hVt2
mMXsb4LGTanjcTULRZ465akOZgqjp2p4nSiiAn3yUZ5AAvXZxO1s7MZ/M0S494zm
V7bZs+/4cBvMF+ZF2+uKmgoYx6bH0lVgABah+Gm/BHJulp6pfiY5GaFM9URhM/lt
aACAUW0syuB8FAWRdGj4gvCGWG9U4y1ovtBNksELNGEw7Zq9BW0UzKpMcUtkEHuW
G4eR5rxDWS5irtiX+1ZJMKzeeVj7B+BbqvhQZ/BOXRxCJOqmOO42CS3lcD/yGxM+
sI8ImYBiqouWLIp+ZeD8OKA/BPjb6ZmwLXIUusFGeE1HTkTSj1X70jK6FfVwefJh
uOCaNYHtLHLRV1hvivjvxhdBsG2z+f/+aw7AafmGoyMjOZhZvfBFkyfQDXs8QJxS
KkQbLeeBIpp5gaCtRyX8EWb6XF5JX+ypv31vKEGC56fouqigAmhaLaBF6OaUQJEd
DAq/Dk7JNMUuQWIb8m2J6zoWeOQTDkLhghHLX/2nIKrzvtelA4shyP7bZWLqkhrS
syLEg+XXj1AysBIETyhp/fu88wqr3M644BRa7lhjcHnigO/IuinwE5cvHC/2Eojs
GBbL/YnM1lVDA+QMSlPxMepRq1u+FoGmULqp1HZbWkQ7nGAo4wv7I+yNcD9Ua+JQ
nG8Dws3clnpzMBDkE88VnCwH8U0WxkDDy5kjO1wjPZY4UMPSDBKJbUHxFSATIvTD
v/gMSgvi1T0F+/0GHtCZEuZ2zYqo3i5YM9tb4DxybDM10m8baSDqNEYf1nn2dF5V
mfmA7wX2COzWPLbH0jIddLqzGBACL04j39cL68Igxe5I5MVh/1PUSg6TATUnEffw
`protect END_PROTECTED
