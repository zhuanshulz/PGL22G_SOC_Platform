`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SEZec/Gjdh/JGeOFGaCC3WrPF0i4ZTK5BxcJesjH/SGd3UMO0ERvuL+EnoS23LH8
OThvlt1lFnXx2hjCQFTOVRgOHcyd8yXpKrjRsyWrxUZD2dD/I02kwWZbawsDPtob
AucI7f/m47gmRlaJoRuiGHpk+KeXmA7dza1RKklzXac7ntvU9DwDOifvbfPk/byr
GxB1vNEIJu01+ZtnaKHrf9hldfgSghLVv6kB8RGCCJfTspy77YEwhyxByCdzeZ5v
g1gt3WAahsguea5lgdZvuRi+zd11oxmWIg/mqIzLJdXqNdJs+9z7mQxtVjFzy4G1
cVX+FX1jEU4CzuSkU0wP6B5BIXvZrH+6lpuovW605iesUaMPBoxfInnM+nXD6hDw
sNRCEeguGZEkBf5DR9MX+8xmGX/MFyqgMM6+Xj0c+gerD1/uy8yU9mGm97L6/Nc4
hJp9EQlGFrCfO17jr3MJTh3a6iLQQWR8ti3Bjt+dcsTV4sykJR1yAR1SmQy1Pyg3
g2plh76GuYHC8CBkf8QDnOxX8/d9xt8YLKZtX+XAhBFYj/if875XrY9zPmeXyQjr
leSQGaOj+OYEjz+FsP7R86i/wJ3tgH1vXtrvTT5OIVoGNWUqvADFhFhSSlVV9TzU
HaNrkrdqUt4dyuCLn/R+MIJ+YeNqpKyZhXMo7Xsd8abUTXNj8nDEFNi0/ZqrbBCm
OX7Cpu39/HSP7kzy883fZUPlBN4oaDSgpzQYP7z3HGbdzqu9SILWOYWsS2ft24OL
zaWshggjf7LAcPDmE49Abnac9Os83EN4hCUtz6ye4Ny5gs3qFFfc6l0DqE76EDOh
`protect END_PROTECTED
