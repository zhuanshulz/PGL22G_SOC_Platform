`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QvAvY1K+LWgwLQ76cpyl9y1VNL3USImHgUfwvvD5ctZS4ptsGvNfMfftKcz8Y674
enHevRXPpi2DwgI3OBSOe3j2sYw4Gr6nbOeqltbvQk70BiTdRPSvZt8ook8SkmmN
KgGmrjJZ2l+m9nSfqxYBc6eyJX5O7KjugZ4SxwSHXEhrCbhrPnSCu4FawQhYj/eT
U6UDvugYfoPA3IJH0AjWMcvvw8vgdefVqxBzgclFvMGTf4lTde+21zI3Wdv11j80
Q2dArnDqm17VqomAXW0eMnFNHrLRT562+WlydMCROK3Mr6N+VeeYBmRQ06dt8Fu0
rVa7r1dk6zj0497yV4uN1/AGl1OtGo6pfptxuXBTnY+Rnx1z/qCbo2mc3fXfhqyA
z6hc8ydkqHGnpjoCdC58oZt0of98lXHpczdz47q8yXrDo4pNTBFLlvVGkIV93dYt
x9uw6Hj8SSu/fBvXqjXanFJ1fAns876ne817+z176PW5xItNvic5g4Kj6dXEfAja
Z+anPZm0wkcGS5UNJDSS1C7n6aVIN2KwFFYyNNOKMf01lVC9Y9g2VsM+vxF16++T
6k0QA8RMOUjxHVrgRa4c4mJDxg8kSz+c0a1KZj0hTvEmF9ZDIZAd4peuv9eYMeIf
wL3UXlQq2PWmb/rPQX5WSGMk9IIuAN9H5Tbxc7fzamclZrSGIRSBnPnNegc2YDWn
qJHMS6ubG5+0/bY6XyqibZCTSsJ4J7rSIx9TDjWfkMI4skoIdZaHnwM5TXS1FKZs
JaYIva22Pm0v7wcWleQPNrfZnWsvi3qoHMD78KGcCfkd0kOjnVmXxH5b9npGwgsi
wYTsUl3vhsh6uFzmbaIIoNsnH75VL/IwBM6VOdMGWFlhKVbn7KvN10HEOM5xohOz
IVeqk9j1u7VTkV+WlAZBYNKrkUbEENlNXuR3P6IXaZvEI2FgnWKimOY/+wvP+YSX
BwRulYcnZAdj2AzL/nTZ1eBnmcTqwT4mEb98okp+JgJ5jFhl/ZraMN2qZcN28Crd
BDdyGZTcuIOFOYNwJ+kYmzTlnq8UTHoNDjSv9y9u1BogB4+EAg54OvD4fcFLWWT4
VD7J8ogXS5VVigbVmoWyiXaWxHkQ/ffyaYvLLtuBl8f3LCvzuEgvjIlJzwKF7n9D
qXCT98YsF+8SEwHRz+75cRIYqjagoEa61fCqEh5pa7XBMCDVCLkzN7gZMm//FA3q
PT2lPAPcCXBLCWT3YbRH0oLe9AzCf0U5w6epVzPj1D1AuStVnqdRddKz0GOuXvm8
Oie4+Msee07QZqaWseWEcP+it1mP/Y3P/f/ZzCT1wDc=
`protect END_PROTECTED
