`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5b56DqZKRyqyFAhvw0E+Afz53eaozFQufIiZe/f3/XF0911NvbAAiG88UWILymJG
QIexSCDyNCVgbA+8qzvP7FZi9G2HzFEscJnk3Hte0uQxuexS1fpn8TaZc1QR0IFX
GTXgBFnaLLKY4nHMKfqQCVKKvoN+dcg6je/VGXS5V6csGTul+Dy3yVQC6AGs2WAr
VpaC4b4zGF62zDI56Kf0HGT8ikskaNRwf5vUve1Br8WURivilFud0WEU24YXwZEI
NeFEKW7NI2MeC+g75wCC4tl83HJk9Fsu/dgICYC+mYRbD4NhmE01KCLeJDeKVb/K
pN209Qo9Km/Y7UYD9brEUH/BsWtluE3U0KhtuFzE50hgQ8o7ejC+PXHJiVLs/5jX
X1r8dzt5bxCae7r3PGnJ6sLfWR3Aat31uNpCObB0Vj0y1idTu8CBB+LAggIuNKSc
TvkVr+rBMgR3fuuE9YVZTp5yHsY2ZhXFUuHoZhZg4LCNAzg7yvAZGhlmPzbDeoAP
ovGdW18rY7vDOJAbr2e/nY4yJKtBwWltCrmV7nNhu9Ne1QQ4fPxbNKaCmb+JSyP1
jQp+A8ODI/M06ekILcb2uanTs0qkcTkLvkuHfa+uiEesGSNYg13XDXm7M2Y/VxE2
dU1mrNS5mWdRcaQAGirELKqPDgGcDmMnfvNMsYCloiMTh+S31OA7m+rzKioLkEHO
nLNmz0a/Twc1ll8AdH0rR1uDTqrtoBUdIH1odRWFbxt0kGzpuQCrl2lQ2PZztfJe
RGRhYJG/r+aUEnacF+ZMc7T1goe1Rh0yZ9+i/7rmPcDC1Eql4NjeCdDBlny6NqAg
ARQH3W53S+XwnsFbZSdJk4lEdhWHyqz7nSKIkh7vDNHGIqezuzu2oYXhbOkt1Qks
u4qb9uDTfz1XVf8Nvo4R1PP4c9oG9oGcqNyZs+zM73gbAi70SuwaViTz8VK042EI
yDpypTPAlW3kEPbNDQTIEUSE9HIq5zU/B4hZDiwf7hg08dEjaNsvlGk7Y+vtPKuu
acSrMwKg9sMu9IGJVmsJAoFKxfwfMK6JHDw0gZJIs6gBaE18qd1LKN38Bgia/VDR
mHtCALASGLLrlTLReZH+yGi7ltQmU+CRPw2P+ohJJh8kY7wt7vJvJGV0EjCPI9Fj
O8vgzIrgKU5CJh5Ptsic0YvJplzlIaiWV/su+NjtsTBIut2DjTYXxG6jzU0xa6ma
zJjo/Gglw7WEvaxT7LpKbpJrtE8RK1i+2ciyks1dAoDz6b4pb2YOQYqWvqVCDbgN
d0ej4VXLIHCSHAHwRlC6d1yDihPXBENiSHGaAqgRNDcA7KAVL9LBd8ot+OLVwbT/
sPZFiyXj7SNFIsxMTT4G+aNIXNm7U3W059itJzkmfSYpZEQPW3f2o/aT8ACeiQ52
6T7wDorOiOxwbnml+RDiN8G1li5yIPHQfEyDhvucq8SKQQG4CUhHFlpjGEcDTa3+
kbcoOKkMQeaaGOBq2l6a48u0mdvS9iEMAS2iao+idpMCucBbgCvsGFCytnESGGTi
qEgn2rJASgaE7efevWnw17vyeWppZpUpsXXerfYcv8nGlD/mUTyZfThVkYLzoj6f
SgDMVUlmjoKhtsALyWOi7A33Lro+adIYMRjGiLHyJinprcjURN+f3Fv2xN1mCDlB
Y5LXDdETx6CPmjFfIwnq07ohYt7rGPpfTi/pLvkZGiMNJ1exLO4tkcPdh1fkBgIw
+NVwMa4p4FPbZRi4GYxYPNmSU0M0vn1Z7cN5UsYpGFWmVnDM1opOw0aiWtk4tkYy
HA8/yenL12phnuyxnhwDdChZJfVB0zysQxgnQt3r85Hw9Y/rD2OpK9aW/1oRkjxX
Zyj07cpVh6pvEaWgHOl2NtyCwv3KLRdIxBXj7fokd0QDl1CO9rlRP/sSfaMtXGBO
hJ5/u4EGViMmNmeLV0SekQBE4RZM6xmpaOtuAPYUWShejjXHtlLvJU0CRgCrjxXN
rsq9lZVsfK1AU7JAESYskf18//vd3n+Wr0Ewxt2gahgGmbS4rtWNMWI3mYbzeft2
9hMxnGPgsTqHWrG8VXbLtji4EcgvJ+lLFRblZpzcDs9vCG8ZwOFimwmKaGoqzr/T
GUElDqNcm/+CqltMgKZ80BCUrplLqlOTP901kcYAnZzdyuL6xwkGbypUuVVzXoO3
J8EZScOvRhMUHMGR0R7ncLsV/kaVN4Vc9UmNhacTK6AWmjWZEUnY4NJ6yGsiQIib
hwAk1SNLiGcDA5KVhDrr2vJGoqDkYm9j40igDRDoxtwQZ85F5pNLrI2Gs/K4b63T
jAHNmThIWfMAooIebrIgXyR1hJPqeoqqCCVHAWyNOigoxdZaaDItEIkDXWECPPJT
RQe1ssNnDWdPTaV5KkKq97eKqdhZuZgLXGvVreYdRwm7FYcFXLXV8lvbb5Uen81n
gyqjlk/t2kNtDmlyrIsTmk6ATlVy8rr3LSxazZo2cvhiSN1EqZGnWVtBTsZlrH7m
k7xL6UCqs4hypJd4ASsrxpKqtO0NlWiy9CKUzbIYRIteFHb+l2/+BgSSXXClskjr
ZJL/0ffu6165lISLQooDEs8t5jHu0DaTkEjvBmehGvq7Nev03rLx5ZfI4xlwBO9b
w+5f4XJDJkFSloj8zMMol4pDJ5x5S8yDnxRA1rSyYxEHBWui1FeImb105+oPOjNJ
pqxvhMDqy13nWYZosZhegIYr05wUMvNnGEx/JyaDbaWepRFTXbh3TBqE4wDU3EWc
k9EKBaFwR6cK8ngb5HPwTR35at4iZRikoLzdRe2vHwGfP4KxWxIXo3OYV+6jxJFg
Jqn/0ul6Pc5L+k2Hc7yEmqUbpdkSXFe52S3LvzurjtJXkZf0bdaSGe3qz0VKJ6Lw
KbX4TL+iuuP8jUNn3slJLHwDY0fwJbWwiVtWi50G1baa+W9b6pgzAMWFrkXqvD5f
LbRgFbow4ehbr0KOfDDR8DXwWBP57WmGCskx33Gau0UP3xJPHjdQtmWVNmxLMoA0
m7D4QpMENTtxWXz9LWw5GYORAQzzCztDNjySzzetelJNkIriKHCKibYpHE8ErhIB
oiqQpfCquY08wc9KDtCiin7FGBjWbIEFfbFPGS9ESKLREiHcM06FmHStQjkR6SK0
sF/MO90n6G0CdeM8er/DBXFqQsK8DhuF5indhgTdHcrm0Lk7o5Zg1azKJRSZVeT3
lOVyxp6HUO0JLSLqYbBXY11Ip9Q0o1XxBYdoNRe1Z58oYuqxNYNfOzv7gzHXsJJ7
mk8wqJVefzezSOLHNsCTSP0hO2Y7YTiQH+2sgutChJk8aXOXrAJ/bPqyHvKta//k
YoVEHFRhYsjJwIcfzKOOySGFdd1UHGREPz22EFPV3lG/ZMflLmCir8F7OydgI4Qq
czKmY6/xcI3da2IJz5m/5Ay0Ebbd4xk6z/WB5EElDHGUTgN7BFZEa5Jf2hpl+n6u
qCcUKZUVaYLTWG4/FMvyN4gIhvA6LwYvIDyhlR/poxPYq6zFXebqI91uTz39P7Cf
5PFbGbWKqlnvm7njz0dNDO60tnqav6YaY4MygjgG5exOVFxxGgl5tZ4qxkkCPR4c
aflaG3EZAHdUAQyD9f87eTzNCUa69QP7yZR1dipXbbHF4dq2wvzIzAfMGaQ1CWJJ
BdbHMvRGv434aDGiP/AHNjTu/gbBJoMTeXCe81tJ24x9dOXzRz3jjmoQHET+FEj2
G5QmTKih9a67DC+BJ6aj5DqpNur3CtJGbnHHndqKyJkUXSLfg5nDOpIQP50M6wJ/
Ke+2UkV1IWjV6sFwTNUxZZp5AW7GgdslUFjDazmIqgqeplWeWjFHoQjSel/GsNUF
MuXXMEtVLlz8lLPKNf6oO/5K0UTmdrwcFEbj24u02BJ2lS1ev4OiQ8LTk+XFyQlN
taDr+2SerxQdLexLGFc7Yr+pG/cyaRBofwddI90chrigj8YThPX5UjcD7g9Ezqpj
UuHloOlePbbapDGWCH0qQXzPV9Y3EWrL/BF2MoSlD6O6cb6ObpPmMj5WPwtR7T4X
azce7XQ1ok313Ci6Jmu2Vkd2CL9pK+wL0f6YiZ47G/tagffrJRJtywDEICkmWO70
flTTYGEJ3h23AmP0W78rW2oHJefKd76J4Vz/0naOPwpnRUuDxNubvyO7JYYbX3vh
fwZW4H4ngNEOAr9NLKTOVbJV0KxRRYj9+c8PzB2dPoyx2yYNl0d2UraDPypPemr0
TNjnJjvoaLWTXaIa5O2rhrYOn8U5eEqorpD783bs56DkpIXOthl5aZRPsQuwMOYd
mpbslStqVjdqWnk+oSoUbOmaTlB1lMImo7Ny7ZoUb55wl+XpwnMgelXxuFlG7uni
eQgwwrroKSfHtBMUckOb4yJH+G3pBOTGlHvUkMwHLfdVvJwyxfNUuvVbVTvEG151
uzAJHeg90lR4WaAL5jyNHJB3W+M8dycOjB03F0IqBgYstiW9+jzkZId9yHPc4zZF
TGhaT8KHEBS6iF1tMm5uQI942Ek36O3PyhfOz/P50wqEyOL7GmNK+7OsgOPmE1a/
rf9Z4QIOnwJCGQUEJDWXK+1GhbhRzCj0PXbijVzFYHovSIO1ELP9PLui+p/LXIvt
b3iUOfz5nCpeEFqcQHXd3KBZpAPzOYXSbA+ZdQqXYqmcDVt3Qic3nLtw0fFxNCQ+
vrjcK4tm3Q1OXKly+L3UASk7j0shrYT9xFkqOx6XAH3AvuBm5r8QexI9rPbtnrqT
RF/Ifo/lTbRkRfixgOz4g9KRUXzFJcgiJMFklXlE4ML4VSHnxo6su/vQRi7dVovt
MwQpUxyvkELcVEOXw5AluRDOX3kFzFo+wULJl5LSXWKTR8JhkuxccF9TnmCOU0/2
JuC3Ulav+H9w0EvROYQ4OXrry0+wmCJKLzz4czJB54/wQl8EX6RZTaltgAg8LrJ3
uwNWLq8LC4n4+8VPM1/xpmowlj43y24YJ/RzElUcHW2lwHIMzsd1YtoN456vj+WL
ze8Z2pAeQ5HO6aOpb6LM5VjDl+psjETMRjwwZZToAcMXExheIH3PzZrulySPq/1w
qP4Ud1lIfdrDs5PLqyWEO1ROdOeyeCMQsQTR7o6cofb+1s556KdCNzZqrnOKgMEA
chd0UOpz+MAuIauRSBkjSI6gxqLjL9pz9f3sHUdvWP7ovcJhmPPajLxzUITsOlZT
sAXhIO7qWFJMpgs1xDqTKGZJZb/ybbPsTVgRGHTCmrMpQ6HbfYwGbmqOhXNQHEms
PvTQpaaqajMf3vFRMMW7RnRMMl6dfw2KvinmSWbfE+ExpFXjSqNiOX/MGyzss0Em
TyUXCGgIDWfj087JyoY44ZshN/radpUwIkg2bVTW40B0GKHVRJp+qjSSR2hdnsuG
DSkhqI+iobzmQGqgCO+tPs0ra1amRnPw0bSCBnVB9ItG0BvaolOYUBDlwP+vggfA
M/f5VHBIGEEIT9JTnlT6DfTqYh1F91Br7CRUWx7mYpZvdg2A7rZyWegTJHXYKxPB
j9yVzFiIbEs/UGTP1S9jfyevkl+wcWBZvA+4WlQD0igNaUiP+AWO8hyEHWCE1BA5
KzF0/lcgWr4YRK2Neo0SbKgBBa/wrQ8MVPTY5N4K2W0yuEYNPk1fJqJwT+pztc2B
Qni+QTtb8sOchQapcINz4n/JbaUzbar51S3uyNWCwyUuA2hzXkp2MlIQSwSv28n3
MQKX0DPiRiX7MZSTpeK+vCEh3MUKy3bPYRxUKFMpRptwho2pFHE7l/RAXJZoQOxX
kjpvN3SWMSFia9+PdbwQrSzxAH0HuGqoFqqbIfyXeE4Xh+uqHUELHLajkynKPjls
GXGqC/xdD1ErpLrt1K3xec11Eb+ZzdiL7FdfDnW8Ro31hAMgCQQy/FCCBficFEn1
qRnFkRHii6dTgBRa0CHW9WOoaDUO/X5YEcS8EWywfLTHZNiavsVDLdXrcos6QNQ8
H8YvAWu6IvBw5MfVdTTOneEzHwX3mV2bc/2FX/2g06PNJo6ps9cUc0QnIdkP6GeP
D65Tr1j+OHT4P8EMM9VKKQZEUuUVWoclgb4FJvvwWy8dOLTb/+0GnQjLxTKW7HJX
cdkFV8mDiiShcCjMuGopqQqk82QwdunlKREDsO8E7KCdr/ibtl8JYjk8RaObsGFb
FS3pGeEqHAk65WqkAGplBakPpEeHkuVfFDQOGc0r+T8TqFovnBNLW6Wd4peM/sxC
KO56CrmgwoXTwvZfoEe3WgBlVdPOT3chnTBW4UO8sVsdzlQmUtnfNqWf1WGQ1uLI
9R2LT5MPbdM9edlWGvZc0IXMTc8+bLHAiMIr+gqr2yyLkavjXaBfXId9SxUf8tMv
84UF5uvW5l7kWmuydPwDTMah4TLFtLL+2vnKa0UBbYppdDLy7lT9F9fkYiHxFAMZ
EpS/SpDScTQOb6FEtC5WC18P2qjWZ7EcE62QKdvZK7pSfDRf747FnUzAFUv+qYkj
93QaDcXb7SEDOAHTfocizsb6dLZRU6qwrgHS4UMJYX2VAZ4TtHCYZVnElxTRA4Hc
OFx+gXfSJduBwdlLDR4leqqktw9T0FWDaJ/uhk5v3gPKmb95292ljslxoGEkb/a/
DTCkRXcmwMNIqfSh3Z4+vhpyLIw5oi/lgwYJYxpi3yqBEU/i8pFEPKfUgQanWbn4
ymPr6aP7yLNQ/zGkjQqsJjJ2+fVK5yASRRKwwdhOYAYnGCB9/rVqqp40ZCGxTDGl
YnlPtr3WhlucwsdzLuR2cZw5d7nIU15AE7P5tCAthxlebM123NYKCbMLHOCJWJtQ
x0Y0dNjO+YlhyUTsYnjIct8INVBhXy46Mj5xwDlSr09o99zytKS5gubyDzPXkbL5
2AaXxpR4di/u3cAEtbo1i157RUltozddIU/Na2DI9NFectb8x5CJeG9gOGgiwAom
pz0D//P/nN+l+2AFPFHm7mIEq41jllkHH3eGt20hNDPiWpq8ODS+mTrhzDT48RFn
7cPd2l+MDFflAEu2VVNTvEYDAwJOGjLGfddO5nQGPvSWzAnuJpeJof+Hd+bK4XIJ
9RyJGuIQ8IXYyzCS7UcN8FwvFq/YyQTCMMlJxIbI6WV943JNz8VDA0buRfMAbwYn
ah8qrN7nu+UwzkED0Lc0RrNICbWkJph8CZZ+QLRJ9Ns6tx11OX1eJfIgfTy3+oH/
fskruuRt4B+r2lWjJfD/04QIQVbUWOkzQBHpzA71djWKlNMnk0PrwhVbijjXW5lB
3XB7F2WpnUmqbvlhxPjEOte1ZAU0xpTpmv4oU+xUD/Hfx6ydbLbwj8Vtcl9JOjVF
Ur39mdhGsPGyPOimNsSxTzXXh9c9dcltNIvdeQ0DO2V1LlODC6hyEccJr1HqEGKE
/5kBiuGUQfFV8sWaoX574P0aRzlORTE0TmUJjJggdClZTaKyCicAmmdBg/macQBP
79uWCLGGU2pkNYTqlAYa1FD36N4qdVfEKxgDX+lLqbAFYGmgRCgAt78VC2WnRXE3
a/IVVFl5U6Srbn3GnvZw3YcNxBdYZeuEbx8A2K+i9vGz4E4UzXXMutfxLTwXZsVf
Lgao/q4Hg67jyPncKMKQk54v2RP99Jasow/HQ8eDzNtRosLL5IdfaL6JcrQeBASD
+2adnIsJcP9gaHP9xLh4xZ6IDZ7oIrHI2onH49xbCsqs+I06Z3w613mlFgR/ZEau
u9xv/aEEoh7IKAQiEBEGFpanf5VymeOJX57KvD/lk17XrUNhn0PobVIcGz9tlFjR
S+Qj/vXMB9NV+JUgUkzBMoQ66R/JCpBIV5y1JP6+L86TTU3Hx2ZsDjxUUdkSqhu+
13ifHg7l2WBSYWOy80fPB54JqPt8LsI0CgOV9UM1yy3C1jFw/VfjUw59spYHQmEp
GU4F2JSDD2ynUYi4646XM0wjc0gAKcmpBfZohOfEZkcXqqCDlG1flD3w+nJPkMwx
IeCkvp8wCP1Ey3W4A5BcTiNPkQ1L/4nKqcwddWamrCvzgCyopmKoVD4STog8NVES
aFzITamMdo37qBdx8OXC+yc8WoRIJrSnuCpTrXkXYg5sNtoiC8QN0BDRD+FF189J
5T1syPWKVrA2t5IC35XZrIJEx71IphrtWO2vHlYyQyhj9Kv2IdvtSo0vmmek++nA
p2FuZ1bkbQNUScvU/IY7bN6OYscolwwsBT31sWqA19G0vxq8HqbyuUOYlRfHXpS7
Dm7qOVwg7DTesizOG/nfIeOvZCJsYqT4vZHOcgvoo1zmWbvqCu1yKdgwATjSfB2m
rvJ9ML1BIsBYEvN45BJALExCWTtPpIgYFurdOyO4uOyHbrLDf5vhE6oSoPMTOELx
wxoa5lvlhRoQIDkQPzyXe5rfze79OvIf+dVpL+ErUhDVslSBOrpuZQreEQvF3fmo
AKuJ9Hhb0d3LoGJP7UNY3O4x03GIUUkP98+6jvjLH+D5NYQFwvN6L8BZoMktScR7
ZeGcIUC1IURGYdfLi4n9JgYDOUePIwDSZpVoMs6kZ07bU7QSqojV5Vm+cpwGxQKc
5UBbWFaTJiYZ8giM1n/f3wCLcND/SgXm0ukuOqgOpPL8b3TU4OwEEkvrh1uPwy9e
2Rk9OCAhrZkwNToMY5E2ybzXMzLAnGkHqV2uJSN21xLixF69wNgC3I9112xfD6D5
bwHCdUs501edwcZNWYYNmg6N4sXLJ0pHrEnUR5kpzcmBL2nO2nbk62NeIJhZvrjq
y4XOSbxsZkihqBOWeRwZCjPeXh2QH11wWoCJZ1JZx4j7n1t+NSdBbg5HAW3KHtwG
0c8tZVEDiU3BnhYGFIEzg2bUHc/fg9NkEW2F+BScZfj763Xr+GtLQzK6XEPSXAKU
rGGRYMcwGlXDQjubUhIhpbeoqpA5Nj9ea8ayXvsOyVS+29BEE8IljdCgXV3USezG
HbtKsP+wWGMMV2LMaAo3SDpjHrjqG81omNoBJZq+xxteJuWHNn4cr2ZmAi50eh26
5x9RO4dWOZk/sXDONShyeUjMdVEPskNQjZIUVmR7YAOiZ93H3I7rkNOKg6VN4NBe
mtocbifO0Zytlp861ae7q3R00FchSQPl9J1V8uASp2e9cXsSLgXz6SR1cL0Nxums
gbraghqcBpQPliXGJwdqEBI/V+3rNIwU/XjKA+5Hixv08OErSujKxoVgfd4zxPEt
0ahWAvomHZ5t0d8bSoZomJo50iWuJ6o5/xIHJuaS8Gs8uhUfnkS9p89BDJ/F7LDV
VApAXWekdxXI1vmxjSWj3IyjJGiOI80y9m1pCfHpI9tRvP60sqkpA3LYWK/KX+MZ
txoqFMIHRC0VPvoD9UOOLsHbMidfyx4TEJ3wB8VBV8malyMztKOciHmEJr4Du5Ak
WrPgoEYXGayqPX7ShdkRm8Lr0QpK2d3P/kaUgS/i1LDeJQ5V9nILrc1I10dX62Po
6cQHI60852vvLEdjuPcDJln0ngZ2Ep1jEqCEzHvHzOa1xlMKwuFDut1O1LoN6thm
rhyXLQCV6zTmlc2plofXqPBo8I/IUaS7E3AdRCiWg/GA+GO+23TrAQjwDcJ83FVp
VjRiCVCIrreJoEe4moAeRVdv07mx7Yz70K9N0Dn2TmLl7Z9kYNY5XljVXOMk638Y
e44TJfpwzwmTWvkXhwkYV91iijT98pOjEb2BWsWpOlvaJUu/X07yg+GnTEz86UqP
xQz2b/DH+1QZcan5nE7nfiSzPPge2CluqRL21Vp6GhScN5fXP67+CF4F6ozUY/8x
0sEWDyXKvYQkstM22YUpqxgTQSs22WthflNfRn3hqtPPIJX9RMLCp0zCfx4Nogu5
ktpFTKxJyk1UKAtRae58uNWkeN3KLX+K36igfteh9C51VyYl8c5T40jPOn6YXpRG
t4/V31hh0KImESB4rq1uibBvZXeMEK2DVNe8dVJYb8EGmdGbRGZzVhz/7/wcC9gQ
4Pc8C4L1q+ftP4tpfzx99hbqnqoU7c8FxZ3LYAtNA1MRrtqQiB8a7UuBFQIn32Hj
BNLGd/qsJjYlE3mXSn2YOLfMFy+RIaO72vRtvSNZHfxkys9+ZmvXsl0qfkUh1kiP
Ph2j9cn/u/ZWbkQgxc0D2ttQCBXL6dt6g+EIudylSdnz7AAXPNkycqcwlJ4r5eLf
2TnxOHTMDC6QEsjnPaXvR6RHsxCnEszeebdHETE537gNsFpwJbWXb+UwwS/B4355
Mrn0ymvKkH0YlGV5U6+JiRd4yBQ4PED3TateIv2Fu0gEYJkVXcDYTbQF1SWJ0oow
NWo+f6qHZ2Y5HN1FwR0xOLLTjKGL5HvUnIYoJ0McSI8rE+E4JKgaPLONRGYFLU1E
FCSFB3KHhdUEOyvfJyot+bGfOzoOX+IeGO2/Udkt9WJVBSdawQqXzz/XFpu1NNaA
NtJ4rt+BS/Jo3x5FIf4+TGjkK4abtNGQLTUenSZuvpxRcRzOhO2plSINUh2qj9VU
8OKOrKSQ3gPXEuiod1DZyeOhuT++OISSvH5xq6OjKhtwmbhcn0KatKrBw8CNoGgy
82xFBJ9ViDZut1//o7BZSIqGPuXsU5Ipq1GUzUbSathxS32BT+NDey4+7hdAshTS
9D/QTab3+Ajb7UvsO4vYeEB05cK9hfwUm1en3qFJTovaJzDAH5yUUKe4hJ4hb88Z
A4PPdWQ2ZXbTR92qgAV4DigvR6YA5/9qvnnicny8A2ctzcVOTah9ZotlpAOffx+Z
anh0J1268iMSferAZas3smLquI6PLHBnxOCWqdHSdFO7I9yYwhlWb0QlSB27OeC7
X+UjdvZR3aOpakW7CkqpH0wWwHogAj+Vv1QLqn/AxJwJLFqfaa/6HquGvKUTssT7
9jXLr9nbUVHQSmWFNgpEoEzHqmQyXxiFVpjsLnrSBbsX3MG4QxQmkUE6RvpsuzxB
Xf3ymTzPKGMyi8NR+h782Uovx5ticqZlYkhAV3Ggtvkk9ZGses/4ICdsMtFB7VII
YQc1LAc8DdxuFSa+zdAVSWyOcnGYTUmZKXtu9W8XuDKz+WkoyNrpOjsR5N35dOAJ
Rf5KBZ67K2hoLk4KW59UjE7r8uU+uTSps8KXcFP87SP70a+rogVG6A2XQJpK3pju
/TN+6LMtTtfxg5IxYRb/KgEtjZFwoSdtP8adHvvd4J1ryihRMEqFljEK/hUyIMWv
POOFOU77sFcZQ/1iYs8sdz8yR/vUXHvivHWN49JE2soUCrVu+kKlYS6Ci1AEfHpc
NvkLABuyZeI31JXRjUw5aXL1vLHQiU/HarCzPgv1o2qmOW03VugLGdHxXqmb/7z+
TU+hnwXGFrpgR833CdtdujS+/uu4FRRKaUD06cPI3ImvVV27nJwqmgWoSN4jYkqm
hcNY3JL9mdEprL/CsNXqbnYLRiGjFEfZfq7Rso7121gOKRKizDWNT5+K22eEi6Px
ptpJ6VvSpLYQ+k2zeyxUi5NUchfXnPfmhiZgRHyCRMB7w8SBAxMzj2fdhy/wBEw2
GhCeOAlVHnTHgOwbhGGv22gDS5jezs7waGTrmlNFSwiDHKNJufv1UagdzcSdQ4aV
44TLdf2WI90FPDi/pEdygyNWi0fILRGGM66E+uewpnFIj8ZHbKjTXF9fXlylA9Hy
zc5HHvju1CSM5n6+c6K5BDN7AGzv+3fv5uMlH/aD5WDzkHQ1Yz1jtHc/f1/vhVV/
LoFaGXrOJFG2shmhVRycstQqyQU3u1UiTsuiFTfGmpC7G9aNmihcH2Kd0gvlKpXb
e3+PxIbiqZkFLNV3zfeygqpQW2SV2eT7RbLjr5CTeQ6cC/L01TiWjDh7V5t20oPi
uqJTCpJ6RAosrPgflQ4DE+hCOZrshxQLkSnRqEKL6Gx/mYtYi9zu0S2jEwU3CUHQ
+mEQCe9b2U/nMUS8GiPoiBJAu+94fuCZMJ6X2pw87ifrn6h3ibfMLuHff14Asfxy
0+wIcfEM8+14Y95pQBe8j9zc+SSsaLyF1hTvn2+pHrCdGdmKqYbHyY7+34S7EFqg
V/83+BXEHeNH0uB+6GC8GkZgdgVj6/e38PeQ9okxE/wDYqEdRkriz7bYfRJISTEY
cCsk5aqtS4fl9X1p76UJ7ualjVYfPdH7JmVmHSB+hDDTC1ad+L4f1Uxts/vRiSuq
IKltyZOsY6+o4Uiu2CqTGBpHvsPBSXbuKVmae8GtocTf+sdOjyvhT+TZRGuoIQzX
0H3KFhANnd/a8iHekJlDqQs++0n0BR00U49htYsCOQGu9wY/gCdmktH8LFBLkV1G
3MHyea0nBErbKKeiiBDgVQfA2sv47G3w561VlzbewPjjRY+3vVYYWdM0hQcBdZXz
in7lokY35mvP4KC/kTsI/zIsmcut7TkFf1aH7FKdRBJLw740UpMHYWjzRhd/MM4m
iybs4ib4tVUkjx6uHWs3qeHcgKLnKeD6x1bMHVXTB9nDksCN77ziuBKHlPqyYnBf
qaInFP5hUegkpKdbp1oylxIbU8YT7qrwnm4Ayzvg1yhqBEKLMgpWa8My0E2UZRqX
qSYF+d1GX7plXe+IA2h+21h6OLEwe07StMnWcVW8pvJ7q7c9hYv8Fu98xWPTe3t4
6E40nC2FfS16KvbOhF9WQBOgbCM9YRZXJShYc45Ljqb53a5lQ3XnzfVerUMgciY2
B1HGhVq3s9OU4zUXL0SGeJ0pZsQ+S+Z2TAAGQZ4QlQPR8CDD8XVweGoi6ysa7M09
LDr1e7YtJJ29AdS+X1o8hjFfb4+oLQxlCSp13oYUiakukvsqtmrCnz5jQh3CoG3q
2DuW4myrXWqaYsiJF6/TZpyKS1+vbeE6PSFq2kOCwWyT+RNlzwCZLvqhbv1fxUA0
HtkGBZYtLw8XEI7tlX9G/VIugkb/sOF4u4AML3G10R6+Jd4ywf7C7K4wc7h+vnQX
zi84+ftwaUjoqQ2FE3nCJHoPk4yghSe5wUraa5+CtUEIeGZ6DN9QJbg7ql6uOcop
unzjlCsxoB3Y145T8bA3UzsI5AEINneye7hpWNU33m+Wy68EwKhXGrNpT9Jc4qgZ
Hjevz+YGpVGP3J9MZetLLZlPr/q0D8hNrNnm4ap+tBlKhTh0j1xaLNNQRKfMBpWP
+6wV03BJTb1xh+fZaVqtsE4G7S7cTJlujy6mgr44O8vb0uso5k6FQqdutKB7i7wv
mel6gQig+rk4dvAgM37AkbnEmbC0QDRIUVmJN3H+71Gw48G6OvPnD5sXTc9oeQWa
J9OhpaBtQRcDd+ISFFrDeNZTJ7eOIX0bQ2lB9V+HvOvI6BCWyjwfGfPsbF7s5h41
fx+w11plfwJtDGh3FWp70/63ucedr8VQLGD09Bg23DMYhachMP7947b9JjbL45iC
j/B/MohYImh0OUfeQQy/EVtO2PdnNvvY04dmGaGKZ/a7tr3KO3CC9V/SwxUCFgxH
4xMEH/Ybrpiz6gBWFWtWxv61YIRhtlazkNP4tJgz6MYzMELsqTwTxqM9bqbthWUr
+YMFJTeTobWMv2BCvSPd3e5SE4cnlxpCrzYvN1t9UfFXWZaebsuuqp0qB+4MPVrd
i+LK+Z7KOCnSeT8tbjPAPHZmHHlv8ISPv1hydeYbub1Tq/y71w60v7/dtNiIlZ6m
QTZ9hXNDw4LzGCYGe8tvTayN54SCjWIkE09OTkdfJpnNoCM9IpdW8Ltg03cSyhlw
fll77tJ24kj1jsICL+wFkx6su4mlyu6w7IDfYZebRlYHCzCqS/O5S3hDIe7ecNfH
EVf0IHU82YDI+FfatT4uA6uuTOAbLtIftIWNGpoAH9URhV9BlFjak/sJGMKh9UVP
iOIBhCcRiCDzLrBDhDNt8i4BmLvGaPdc3Srb3hZ/Nfwvvvocxj//4pfj8xdeU63p
i+L1dElX5wUTcePMZHAaAVWOeI2UtJy5k+fc3bm/jGg97+i5uShQoUEj7rhTXsR0
bEw/dIrLer6sfSlibZP2EQHGAWKWKGt1rGvD4hdEfN/ZwSCFBvaBeb6/T/U5IXcE
Q8GPe2n9GnX3oa0NHooRm1dvAnYZ1FSnllBiEd7rTrT0l6cpETpucVJgAx5O3tTg
BAAv6rBke5PPaVSkv9K3jO108SJmLDmwqPwUX8Ipf1IfCxENt5Q+wQesyNeuORtq
nr8AN9Cd3t0TBy0p0kaqZ5rGiTUk3UcUPbcm9THI8L1pRIPJB60bpCn8cz1NmGBx
J9TuIJ0UdbxqGD20fUSEzVG300rJKDY7DLX2pn/O88QJK7A7i2FkFMZsunthF/t5
LLfYSS/mIJJiycuGsF1llH1NxRkfvj5LsZG6phPZIv5pSfzjo8p7CcY2WibcDk1d
kXdBujEYFJg0p6N2omGhIn51sywHHIhDOUsBBTPLv4WyjctOLsec0b+MVRtY3INK
vutfVExx53RVA8o6TMslV7DWlfFGFahPVwJ7QpXoRuGzzf5cFnoe3IgFGmmF+qH0
U4aEvl/3cv+TKirbjN8PpAMwMK81MlpWpkIRZFghFmFc43B4ZBv8TtIAw1FPMI3d
WCRFFqUs2d5bq8wWNSE2DdHEGXCJWb+XH+EfmeIJEyPH2og5b3apv7O/a6rprwa/
G17LoZOM0LxhX7zyGY+3iPVdkYZENLjeTTgcf9weBDwifQgvQpo3u6Sigqkvraol
ahDFeboRoYRqPEYqVqr8FVYjGWJJSsZByHC/n2FlwGWs0+71Icrt4q3Zsn1CpPJG
o8GO4yUbYWi6mVpyjrzGENEZAEwd/WAYk7bJiCA81tkRxQ3JubLWQdUQ1t83vGoO
ZvwIw0/5k3sqSIqkz36pJbc8mlR4KuWhCcsxXUtUzdegrBBYLWqu9fFt/srxIb97
4RgImpcuJPuj3fdDfcDEiCRgjRq9quYCQeTiLd5CRWlqgx/cfhi0nGvFmPz+ChpL
lugTuuZJHVe8kvYWMrqkZIyu42sergdG0k5bOt7sRHi74HeU5HZB8D83RYJfOrtC
bcU2vpi5mw56P5bPVA0LjDQhqkyi/GSVgKcpwrjkpXktTyR3Q6jOHP9d8+L2ktyH
vgd28o43w7rXL5Pzt7JBqrFpdQMXfwIurn7ZvHPnaIftMJCTuyj66QCOYC7ZsMBW
rJwMk1k4FdA40FdESGCQrfOO1A5H2v6813q8YNN1lhjAAI/M8cHguaAUYu1oj6xS
UWIWgrV/Rsc9szudmlASUUisvy9aqaSWva/a8CsHcnvwLghPOQCCD7is1rDXeF9N
6/TMgtlPrv9qgR2qHiRdHDfD9rMlBmmx4ufyx+3o6KbL0rQWA6eRiWuRkFOfy1LH
EOFvJk35uK9aUBnvUEsOEXWFveggEEqxZLr0NYgOHBYFzdKh/ee3MSDR1y8WXV85
OaANMLzFM/J35CvGFjhnd4AxHuyvwT/5PvvxHBbqQlLmMjiw+jOFO2t1d9T+yqVc
NmsuDHglkAdkynADjYt1x/oBLUBmgy8MmPNLqB1U1GDtlXizGjTSEM9LgHzatanM
KpWFhx1EXUpXSZVjaArT2pbl8ur6JBozSQiWsQFJABNNu3H59PP/ltyQagQm8Q0o
v9Wl4I3j0KiFg9cG+5ux4B39WImlEOHUpH4VkW5jWruK5GyKu6U+bgKyhvvQK7oG
lLwi78Nus1likWhSK9dSBENLTFpjY4LX0eNSkxlQmgFNW9ZSkCDP/3ryEJ093aVr
e0fVYZ6fIcITHPGYVGaw+y5nRzpgE61RGYQM99jxdWMuQvA+0NCiWPXE9Yz6wtAy
XGZ8CMm56b9slS6hb4o+AS6O6SA3c/D0qcJD8usNlEmtQnB6bRLuUda/pb5R/bWB
h6mJDv6p9tC+0wyxqzOqxIMfQWyPlQ9wjRr0G86vmQsEWI1NoG7FTARAbp2aNEoK
lIoFjV8b0vpLATRW+3y6guE1luU0AC6H7lwHow27W/8sHBlPGz0+0mSPNQhXHV0A
p8HLbnCX+y2HuFqxqihI3hC8o7PhduUJUFN1IA9R5s/5wuHgR0rDSdlxpzGoYQwc
JEzQ61CGOpcZWgkgN+bKaTRnho2WPcjW+5GbRnceeRvc5tPXggl8NDuxQn0bHX/n
N9YztlfblzXEqBCjY4zowzKjHr6Tfhb83TPt5vecBBCXcNnehmkz7Fdsio9gdCZ5
aHeAqQ3Pch7e1gu0ZcEM04FSYWbX5WiMXGtDKXAlKnRNZNZtTJTwoiA93QYKN9Q+
f20Jucbs+h+PN4YbEf/IPCo0CAY8ahsRA8BRLFrUNYi/o7F8wYr3pcIwBY0jr5iu
HFc4ilxRWkZvYsy+Zm23WMATG/fzKSTxlt6aCGpn6CHpaAEnymU35tvY15FlKwJ/
3OQ++InzTcj01o4PtlkItRTXQiiWypLYrGwJ92Iqv0o7NWkB4jnyOL5YUxi5BbdG
LCVlEKSF9tR0PZqmi0CtuyrMPbPi1tdpp2vG8jzDQnDft6/NmapA6vNRPlyZQ2Ss
G2cqjYRv8XvIAMf/yImCJKsr0Mu7tSnHr5WVZkX/j2gAsomETnLRD+KdKqECevN7
qwnNVQRg5ky+WzrAB6lCGCXpbhRVQzz5HvIHtNrukWtQ3hTivk26xUrc/yg/CuQt
urLkhUOqfq5XTAFGkpDOsc1M3BUpjVDC2befTYRJPnvGEA1n16FCK9d2Sa7qDOa9
8Hst22LXl66NH6yK1UHtH0yH5QvEgIyYVCgAhcNbf4aoEyVqYsn1qO7Lf3DBtLTT
9Yn+TQCTFGzq2HbOpM91i4e1NTcDj15MUfFcQtAPBLgyxxff7riV4jikwfX3wLpl
yKNuskQLtvvoC/3EJaTa79JzkthGncT7L7+nGCAqNrE0e0aKp+pTyjCopaIX2UN7
t1yk4d8ESm8ylMj96thhuW2cZmjh1DsCohdebp9VBUSMzcPSW3dy5t6vfyihcn1t
kH4sNaaRf77qffUxZbtcnPInh1mbmydO+YFboFC8xUFoKzZDIS5ogd8ptRtLWBfY
WCkupUT8kAtqSu8BPlGPZVlEuFJxoORzMKHplWoHmilS6L2VAOM79g4iS2ssSUqK
h0xGSBANemNceC+dyrFEYzmpStuY7NmFYx+BLqiGccqdEEMMZvftWKi2FCbSNgIi
uBZcZvZIGIFh/WZgrZqxr4aXSXm52AURfVuZPwWCbGG/yk9jG1owCzJ40/D5GGMl
b0vMQu5nfCkF/ZT2zzO7bBF0/1hlq1tZTJNhDtN1LnrSQcFzCiO0j0qys+1cNz3q
xORVhpdkMS7ZZCZxWhL1i04zZp1Q4l9UNvxQxykw++aEXSxqxoHR6DpIvu4NlpZR
biUOdUrRi8zvYeM4ZnRigmCovaPYNb9x3Z4rOmJ2da3SWMpoMc0Cvs6t4CO0lM+J
kao2e+iHLxSw3za31pHyI6hIBqFJxk9j9+aQxWu5FLf5KrD+7dFOyP5nMHX3NqJ7
8lwKIGbW6eTm/vll+r5vfDKPAHEAxW4rNJtQuSHs+a7I+s+DO8ukX3S0iU8KUrJZ
aXqzi5XLmPLXJYc6dLqALAve9CRh/oYzlRLAySw9vLylSbhwJPETcJg5g9EYbNVS
ocZUPZp92TM+2Vmt1gov8r2/mpPVPuFi3GTQ5eVsiJdosK8dxzuJ/MBXOEiFZTHB
RD1CfeomVZxloF0Cr6wKzJ0T53JVb/kFL0Wv7eEtPyT2YMggsHiB+j1AnxYEf2T0
bFgWHtkiFWOO7/VY+p7/upR1sOkthOBMeW67kICiq8EZ6ZNio/o7oboTqQF+KKjM
IImKhQopRe2BXmnAiJ/k+UVRJnlqH6b2a/9v7pniY2qEiAjFMf1T8FHtpl5FV8yZ
urSaGR7CUIzseebMCabZClONQFmj3+D1FPH84Ar9BvaH0AuXoMnG2+3g5OuJaQXO
eiaUnA34oMwsgtvfoiEzY0ausYsOK0akJWa5B18EISqxP+sBAvLV1VGynXQj++Hg
n91aAUHaOFYIbjgkU9QqGTi0nZvGEC/PP774UB++NojxJsWyT0B7VkbqetbOTjFB
k2yyF1j/DXWzDesQYobvuYLPDsOuBw9alrZJ50Nhtkefzg4YIuv55/bQ38FElvO7
NtmYyOsH66MmTALQL47KYv4b/YjEKdSKFZCN/hwOJaBhcvR0T7udpFf3KhY4tx9J
HbDPzlDgcCnmzAqGRA9oAz3HAPVLB0v5KHHa4x+9IN3yWZ9x4UGz/TR2fHee2jI0
2BMAbz3Upupx0TTO4LQ1pDZr8gbn3Vwfg4CHkuIyWVDzE3o2cqyGYebkdtg1DZbO
wp7ONECukpYDhNHgIojZMhnkgos48KotOiynJMIPX6TyYG0oP3YLW66h6ngNHiSN
ZkYvUWcDhsh+FU9Nbkq134LL9o9I9BzYUipVOZ2rahYiVN/6D5MvXVglNFG13nu4
KCEi+XUA2TBRVSz9UBtUFc85C0MLXd2fPujN0C0PzwFViZFDcrA2I2MmPgw0tUmv
R5qI4KBZS9ckv2Pn7MyrIGPlSZzLwfTZPsnJdPw9eZeRnqCDcIcYYfCpcMR40/Em
2EyJVyijkwdWnEd3oBP/qmm/4kgaAa+LaI5CSnj2jqPwpWzv4pDae6qXpeXsCvHQ
sN73jQddKckpVl9v5Wq5t6m+n/BIPznXH77GpRdDWbCoSEsMCYTwS2uAUGKzcV/+
5TgrJbX2gAzjQ9ieadR5wxihd9tkYx0nwilFNTHufr41G9yFjgF7ZDr1Ns1iDVrn
O6J8dyS9NzYMvQy5lB3RnTGDLebTInDfHxZW8qASyK8FBkLR/FZaCt3oQG4On8/E
ciEhKx5B3lgQaK66YlWrY35R9W35NUASt1wKcbS+kdCxLRryLiNJ2whGtnwIJfbk
qK45HzqQ+Gv0DjFKKJ0ONbvSw0qWC8nUEfF2NjGL3HHhwgK6bZZsafL3+aDehbW5
N9EPCjSpkAGMHnvXoxE1mBN8rVF0ySQlnKZOYPS0opYlFBJr12WfACcnae7LURCu
Qjv+hW18Ha9/JOycxbsH5Dpn3uQJrW7Bi2uD5EZe1+SAKs++HWxtPlHD++/R2Pa3
KimMGYUU2TWNLWnVRR/Ckm3KQd0QCMCFkgDWUwJaDRW+L3Hq05BzcoWpXBDHw42q
VKa4LzLzCg+1LIx90T5ubEfy/Hzb5X/rhTTMr9M1N2k9V4UwmAKin6Wa8p65B4Qo
SDPKa2yMpZk3Cp+ta4fahv+nfsUt6T0kBF0thvu7HS0e8GSckvxfRdKyX9NfwAe4
cGcL3NgiCgZKJzW+6HMa/wNrASs/gcDTfxWd5qRrqRnhtXbJ3DAN8mmRVO9l40AQ
wgtOu1dGOlPsDObs53M54pOumgH19NgsI2TOFIW/9BGc+oR0/T4ktzXp0pispHNa
3EVgOliRny7xZwia9SSv5SLp9Z9vUfjKB2RVRQ5zktEqXGzGnn9myMydTdpYWoCD
JTuF31ztOVB5uU0FzbkP7BAH6CLS/v7VALwDbdAObGBmRLPw37m3l4THqIYCaSzZ
pdBJ/sgEB4/bHdxsOofpCLMAU189srVyi+EYsp0JPJ/6/hlUPp2RN0PdvPLBCw3G
clESQxkx3RIjW+0CySxednI/ZbX30RTqQZFiDUxlItldUKTUgRG9JrcKiwhPNbbz
5ntPV/XPgObABC3d8Zp0y/esU0B5UuuSZS60VlEF+y+zCVUXpfv4AaeUajI6Bp/M
3hd9tsvhEjDfsQY2HsxxZfwMbVtLuJz+mv9DVAH6uMxFpQrFMdga5wHyh4NtJt0/
8O2VuRd8gMR9jDLV3Hf9BrHDjChiXSGvlj/cImDE4JpRUPQEvShjsFFiCEuLY9Fg
wGkGVEZZTiWkHMxvyQmzGTJDVPboORyqlMZOTYLRL59i7ADsBW6wkMDlC361bSSJ
gAYyXZ1o/1JlTP17bQtgzc4yE8z8RD3DLd7/eS73RFt939PNBPmLUNLHjathYzXb
/UBnd7m6C1WRRJO1sSrcl7nPxUGmYh4XnGgUZm5QR1E+fLFEXz7Na2J/m4mYldpB
f/2VLiJStaN7BuC/rlx09ilcQtzA5EGJ3EENMj6SpMt8odSzD5+LktN4xp2TWhAI
lMddq7GwUJbImRxR3hWC2rWI3E8p0Iec5RT9z7JIXUghV5krhnpZ5z+ebVGhq/Wf
uCaTjRXIAgHcI7siDWub1Bc531P2+hzkE9FLOJz8tPRB/Gvgz1+EwRbKG/Nl2/vh
EOQHV/wV10++DgYHJz/0jotNE68cfoZZU/P1uPlWs5V8EQidf+3YJZn1VRR/h4LK
mSrH6qElWDgJE4lm1Cec5pzqgnxVHwLNIlJbZnJfnivp1fjpxZXz4eH0hHa7XkZe
iSj0QK7iK1usDXrkqM8OLER4/D0MNkUn3vmqSJrQlzvgbGelo46O3O6UUKMBezUg
og8VE1tcnNUtUpBXtfEuosT/IXYB7aE7nSLtEIrCzrjTjkaJNLpJ75wDwL6Fw75R
yUkaQSBYRV8o+xPFrgoqM3X5uU6OotvYFT5X3B4S9EG4hiyirReRnsLpgPzmdmJa
mxYvUzexWddLRT0Y/+CJT+RN2z8lKdncNGjDd7wjOPZAxzGVScW8UYw/XZ4vUgKK
Nug/qQl/xMPz8+u1/aBCZUrgSz3nW91Qlfm2Ok8hcm3Ygo9oqvrk17URW1rMdSjI
SAOk+a6FLWKHzCO98tydatS0kuXTuk/b6SFli47qWNfaAErlkvjr/SlTqrVAKRP0
AmPGMPQiz1mq9NkAOcXZlJsPlCSWlWb6ps7Btmm18VK7nIUyWKqzUMQlJr1krucs
1M+MnVdpfmIV3PmjrsSOHqrvwNATd8/iIvu0o3FweaWvGu2CXQ573GI0xG8daohe
PTNcTOUgIAvMk86HK+jPgBIJBvFuIOaGbEoVkkdLmpGgwyUh9iNjSRahbAQQX+G+
7zQgHSPJReFoeil0+hUAKaoXcQPT4Xg6Tr2gHXz4OthKR7Vcmx9j9Kp76DtxjPMf
yKC80+zipCUX905Lpt7lfrjeq8qU5y8+Uh6RHOPTUu+efFsmfPRgLxYaJCmlVibZ
wVEh6bckJHsFo2DmRdJ8m951SehFtNVv8lslEF923UOTmSQQ7TBr4bdB8YZjhapP
K6QlD9418abMLDmve7SFj3agPmWlWaNfmxlKPvMm5KpJokEH+XmKa4gpEE4W/xIP
8uIWx9XsD8JiiqUXLWjiP8+6+VcGF1fMqfIcE/HHUY4/Xy4Gd3blTm034RUiC7L1
+X8ZnQOM1zcY6HjIGaJwGsUjpz0buW+dAVwAj+s0z44Icea+Hc2gZz+nlECKjSNl
OkFzPIMrIQZKmCB0VepLtMMnXG2utftCFo+ZsDRdhpTWUtW7Lf9A3BzcBkn15n+U
J8qegLxD8Byl+mvPV+nAzHnUzZMlzZLrktZ5isWjl/2McBg9EZn7SfSDMT8qE9Qu
pWYujQXVO56EIW2DJrLR/o+KouPeTklTuCtPZjKIEq1EdftQSyUGGfFlv4OUZ+ix
LkBAgcZyr+vYCydW+H6VcvdNDCiXGWVtikXJDh755jqbrO/PlZX0K8AjWW9e4oeQ
B8jziIi/eEsEf6HZQFnCoB6tVzFPlMvlU78vhirRcYllHELDl4GeXyR+Gx2XAuDs
gRzHQjqJI/g71CZFG+e/Y+8+Xk4i1p7/3oOGK8LNx0aXMLARHlSAe01+cvzG8VNS
vUbBQ0WkO+rHVHUgxLqg+r7OfYnu1uhDqKi3vsqOXczGyUbO9IqubOdxHafjtGQ2
GWCgUJWXh+qkdR1mHn81i5SZ4xtufIXeYyh7cvIZDAXP+zhVWB4DafOqBa3L8VWk
/LCxo0iCPtW/MhYq4hYbjIREgmdubhzWmbYgtlBsWF+m3HKJUZ7a+FvRTSjIvAqA
RjYLECS9Ahveh9izcOFjrUfW9HXGEIcdBCr3Ylh6EHC4EWaZ1I6J9aVsHR/0K/OG
0bOFRF+YL7FmJfTcfNFr61BqGMBuUzv+L6Bxn4fupWkjgrKCA8IyF78Y6fKQlF+H
wjw4ZwdgE9lB3BPr3bL6S7HoOxOW8yO+nf5/b7DeIf/sftT+YFEQ3EMMI75PfkmF
CIBfVvJ449tV9EoE7OuUmjaoGi0bdRzC6vrP6/qStZFyp7FJSGu9QFf9+nU65wqq
ECVD/wdwbAvEZixDV5Zx0wE4H4SDuk6Yul9vYn8e7I5OnRyReFMpjMGsB95rk55n
523OfHf2FwplvbDnEcgTMQ66Ax1Bu5/6unJNIW7YMKAxFsATXxZiXNoQLvkOn+Z9
YR+YiVekSl4pQQrGgIA5mfqUi9ZJQKq2qOnQlFZ9aczPTq0WKtjIooMITzbhWjH2
0aBKbB/sXHg+/IRk8csV1VZuKInku+kKaeDIMpSn/R+8lS8Qt8Zc7FOiWUUTMWOP
HMitgMQj7A1/8kXcbBMtPk6KYM1dEMxt3F9It59WIt1ai4LPZe8bBJahRuRBxnKl
JC3ogFUIFhSNeSIR3KKoPURTz+9XZyBkMQZYadzY6BTFsvF7dXqVnPpof8VbtXzc
b0U3LcinTQu5GytFqK5NCCdRWmiPXYJZgxJOG9y8UrUWvjtDxziJMXqCMBiuH9MC
30RQ+XNmSnn3AnxP3Zdww+2R3mGF2AsefDXxZB99MYmLi7Nj854hz2rA5O3cSrh0
hP51vzxqWxaOziDQPcnDbN+Pq6x2fIKILPFZP4XTOIdC5b8sO8Org8owu9vBEdPg
qoH0LAVsxAIj9v3Q00UhDBMA13+C/vt19Ym1zZN6bek6GqVuCpRzC4YjyJ5MMr3+
8B/WLnGY6zFqsko1y+3BucYIkfLSTjUBxaYROdjtgoB2Cx1ex3/+JtoiLo/dOyQT
g2gOoyFVJQtq6gCr2lWFXnGZRtiz58xhULRa/s7vmMWCxqpss2kwm7bpR+OVQXUC
QRQ0/eLd3RGPWiN94iAbMiZz/6MY8By6GRcVpw2pYr4dMF16SPM1SRybL2EikvZQ
CRU+6E4PEaXLrVceoH1l7t1i5HDw37AFMcoNwjmlpxMRykIoauOccOEf8N3mqaQR
aBiRY6L+1MeF9Iw4UtR9iJzNLf5LrOqPcI84bItNEdim468gv7AtKgcjHWJh2iuj
RuySlzMNV9eD4LFBXKthNf+z4sLhtMFKhx+WpH+uqtmAhdP3vbr50SAG4In0izcT
7lD7sWDHOKqUrXe8Beq+DiuV/YQd3u4NAsC7oEqMBEvNqfP/PadsIsZugWFdNx+B
EA/P00Cp8KyHdGkYTsZxGx162ZreTNLc8LEXuXlC4d2Sv60afYFhmrD+Z0/6BJu2
0RybmN51l8xD8XaN5XReBttNPvwDhSKEyY36VzdX0oE0X6qRx1vXgvgwNW5nEFfG
c9AmU0WwGCrLJQrAjLCeudS+TWmmI3nqAAm+AAFqyCdtoK361eXVgLgfyuXZWUfJ
Zr6yY0JxHLEWDIX+GsI29298oxvfnPcoXigXVyzMfppnLQVydmMrV3QKIotPMJ1A
WU7d6+7AS7qN43GdDA2F65HyVuV/m5pezqC0aHBrLEHE+tWq3BBZcFxXLVM0nhib
tSZf1MhR+T+0dT3VKKwX2pgDU9wv/jxn/O2c0inefDHXJ3yNGo1N0BdeYZu3mAFg
TyvqmkyfEtGYv2TOHPIAZP8bMaUyrwD96XGY4G2GKFPYJco2KFRjR9anDjdAjPaI
dk4lgfV6qVqP9neotK4/+acAEWIq1eDAnOjPzifc0HNe30Pms6WYO011nNYVOPpT
1ic2U2Qg2M+OXFJa3qlARmEWrn9IyKmenDodBKrsPgokA+RRg0xk+nc6xk/U/C7B
OuMjuT/ekLNdubODYlik4A0+bt3iI9glD+pzTmXWVC18Sd7eUW+Z8PaPdkfbFWhW
Hp0wC3wPQtQfGRbPiflDp9GaeyUfC6dNvya8NFdWnM0eu2BvMTcHvKGoOFZDVR8O
KQK8ka+i94qAL5tlje6WxZjzFSwyYPoGQfg4uyu4SZms0hIpGYOyHRRxOCbdrGYY
TQ7rybJC3QWqJyvNhvM59aWXsxREZgAoRcGiekl9PtfRtSj6oo12bA0PlHpuIFPv
NgPyY1XNRsZQbCYcdCz1/quA1m25iJKzJh1Pi6yj3yKPcJ9sXNkzS46LMTI2qOx/
NhWXvUwzVvtwgzP+5lxd3K6LuVa7Eh0SiPj0G7ACFIbAmRyzLQIxc2JJVb+X3lkT
ld19uCRWE2PJy61cENWWdHNOPRGEWto0DCKR0I1wmxbKEj/djaYTJZjRhcWzweQu
RZv5tN/SXr72rEpkmmt1oHRAB85Ax+gg8hVAql/RIGB5Urb72kRoclwtUS9UcQsW
XWsa61rApVfjrS8oGBgiqOTpbvOd4UHO0xm7wMgZZP1vvA3VvUTjmZWThYSHBC/7
8MagahOvDLFbaCOMNB1KoRph4IonGdBR8+xXsF/+dpZqRd9Q+KRyYiePWvqIwsrv
EXD6aM/4m5F0u2FTNaqcJxMGvdXese28WvlSTqvm68UHbFDJFRTv+xVDcHq0JNfn
F+uDjTBB8REzynS6R48oXDhy7xzNn3m052P3GPeQYZguAsu6pCjVsWa0zNsnyFpv
zdmOiP5Njz0dnPGDW9ftXewKZmxFNkSgbDGSwkwERrIoDon6MImGSJ3yYwsPlx/+
VWmpExAlACcm645Aj51Hh6GNZRoCbFlCnKD4948+FxFLOPCMlHx9nWAsvzixzYuk
Tqqg9G8+APoUZefaXnXqsQCf+5r7pQ2WDgaR7VFVKfxWbQd2T58hetAG79Ola92I
XrqnAwQN5FOMTry+DUljmcgQ5yh/wm8ii8hYU4i1uI0fXhAz2Uab91ZY6t+02/OE
xgn9RhPVrteXsvPeQL+Q1UakLrDmZhHsO4x0IW9dkfRrOvJr6V3DebVYQBQj1Srf
SQ2LU0aSrWoVqOrC1oPWhHlmbyDopNCoTM/2a3OA71npMN5zvbTDtvcO6LXgpp7r
MQWGkl/q+LF2rGalt2DrCrIlcB8meNhpyHLx69Dkz5vaMDaFdOwbYza2f0E7G4M+
cnKSw5s3+2BRVbGelrha5UgoXabgeYPJ5Xmr9RIM3wsYaPcxyEvQs6woCJfXDmRg
SExTyqa8PbKXy0TrnEuMSQ4sRGyVCJQT3NoytGugPSaL9VZ6YeVBIUEknrhMxxR1
Emq3HxhM9vqIuKglJybY0AwxhO9xoIjOxXhcHvIMwGIPa9MOjtSJSNIIKE96P53n
hVKYdfeM924gDbJDE8PWXBZDW/Ht9KMst2z/1P3oMkJ4K1BU2BuuGxhKG1pX/iP1
W4NVdx1NF5rbb2kyP/SP/dTHF6b9yqj7Fw7yJhJ5YqA=
`protect END_PROTECTED
