`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HubiLOHVnhKj8VAKa272XwoE3UyeUPx+ltRvhKQXRWFtem0wenc5JSPw9J3dQpti
6caFZ1xHraXyOsHQS9jY5ccvrTC2g/bTIUNDZl34LGX/lFXkJWPFSN0Ku6WAgp3o
OPhzLnC2n5t54rNDzeNPJo+EC+Yp1i8cizokY7mnnBuKSRDC4rDvnbS26PO/tGpn
tvP1b6XDB5tDcXGt8NZNrX5c8/2DNs0CXbT3ah2jMbu8YQ7VorX6dKwxGCe5hsQP
VYrM5uxz+HPzHjsX3zQmEhr0jx4UlDAFdDgkgbBuNKZXIQO9hIoJgILPFKhgodZm
2DCDab4VjDVA5ZljLg3gJjMelBeLTqc2ZhxXSqq5A4S0a+XS8S1eZccLcLsxgv0k
tMEGIDeREmALDS5WKnvRxdqpig5JeoITeifSLhEX0Ap6jETiEg0ttq/bFFy3FcGW
2fVHQ0lVOxwWSGLUOxfy17mFidn9W+UqL3F9LTwL/1KidKSU/hfTjjTt/0ziTlzr
o1mR01IVeFruGEFmHu08kDj10mP3No7GcNGAJ3nW/+ZROp9Noo+oIL99DxMGakbQ
RB4krsST+EeWKKBzyuUDXIpkYgQjSSOL0GSMjVyWG9QhLKsLQ9JeEvBPwSL3eZVY
BNluej2T5xmmEuokdUK03qyk8qZc3v17+pLCUqCKNUusjgQ3Pq6IQsUetzMoWNUO
GjQzqa4kFD3mdjTGQmKjc2epgmo1TX9xPKc5WYnxddztEFCoDVXTXBAzdyscUFyJ
9bexla3aBpd6tkF03GpD2t8O94XffD6A57RFSQgoF6o=
`protect END_PROTECTED
