`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXBfC1xp092Ox+FiiwJAztC2HI4tnZ64b/SkOjl/HBQHoN7UcMtlw8yXtlDyPuBD
ptCWHhZUkTNRigrlYKgmOTudrAk4P3mAYdY3ebYYP6uMYR2R4416jmFbMWRwGmkG
kDFC9Qnz+keQDy6n0jgELSf56uSniDAaYC14bXiYC4/0+de7FPCssv7o4bMYgckV
yIe43cqqrUnvljK1YLUFnWBRnq+vRSefAU/asR4c/1RAwvawgh7qtlgqPcCiroiQ
D5u2nod2sEqZPpozb6Nm5LKZhz50n7UlsPlNKwiGyHi57HHarWiipjdx8VGUjVJG
B1Y7JsOX1PRt+819g4Bg8pVdfg3cuSPMyfwAaQKvkYHJhTBu2EhtlsgEJ0z5un0o
6FYn+E62aP+cTCzxprYaCcL8w2RTcUgciFsZ/xQcnlyhVwn3SpiKE3Q3z340IbKt
OJ5Re31VWWrwgxwag2mKqyorqzJtniFvh8XjCZKCGBf+GU9UcNIviEapXcu5wQHP
HxRCAyr9Nd0NhSgZYV/eNGxbkJHfHhH8RAKdtQPG9+qIrAuCO3vr40zSm1L/qyEO
DyKucH8rXqIbzcUzL77J9DS624JX3DsyoW0XYXJXrj7aYz0hCxR2YMp/bHlc3ZTB
KnI2Ikr4d65pbd/giFs6oEG4lGnckFwipsE1SNj/2V0yhaYBwH4XH7VRxtbJ/n7L
wLT4aJ9FFPLQDzUjarIIW6lq6Q/yCn+dWxANQd5D6T1gWTwEMgpxMc51k7mWW5+F
XnvNpnmBK9ZkflfhGb/PYes3X7+SXfw8WfKqEY+z7e5ZS7vH0uZaM1w0eaj5zlRs
tGwjCc8ITwee9DIYM0jP5ajfKGMdBA9Vpzuxz9D4jARrCid0sdcOXUA+/3ZCncCv
rD0BFN2i956Fp24HP1ctfZo7pRykwnsPzl7By+N8uUIdbeuVU7J4T33SMj7zHF6F
sk281grN+CZpTuYgS9/iJ0C37kpRo85s8mEvFmxlLvl9NA0jFYfuDP0hLMLED3Yx
wMSsIT3tdjjDdept2nNSvFMfjjsG8pAQcyV89c/34MNM2PldDEr18ZX33rA3HCcm
wAPT3nfpSc7wEsb2KIhgu+ybEE5cvBzzQHNTtNyMTDS7qdt0plH71Ve/OEqKzJCY
6O+bUzGEFPAa1Dpe8+chxCkwNpaZhhPvrN2istQoyvWzOd5fHfpSkMcHqoNg7028
WkYAroRXT+6fdZ+NNLGtbsX7qX/iMzzYpcAYAyjPaP8QDdDE/Zsj2ASNkCuIoZq7
FDPrQ6W8vo6CbaHQ5Fb9ES2EaTqe9NdEcrgHlqJorhcZL+QzqIZ3udtyR+Qvgq4r
SFCPS+JK9WEezLmkpfdkHDecmCujZBP6ipFF3Sj1gqTb0tMChkgxZtr51XzPFLmN
GB9sManPpPcA75I9Eka+SlLIPjDkuW+j0HsYPno3sq+mLgb9uGNfJDTGOoTR8Nkn
nHVuKPmdIZRsJ0LtOqMBWH0+AWD3tae3O5pDMmAl1m/XvWSQ31ISpBYaXX9edFuA
y1+4kidn/0H4VB57ZM6Uu2wTJ6cjocgmKgQ6KdCu77GjjiUK/m2SkBV1XkXZ6JEd
VhaKNdsjXSqdBaOxYAVIgA==
`protect END_PROTECTED
