library verilog;
use verilog.vl_types.all;
entity GTP_HSST_E1 is
    generic(
        PCS_CH0_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH0_BYPASS_DENC: string  := "FALSE";
        PCS_CH0_BYPASS_BONDING: string  := "FALSE";
        PCS_CH0_BYPASS_CTC: string  := "FALSE";
        PCS_CH0_BYPASS_GEAR: string  := "FALSE";
        PCS_CH0_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH0_DATA_MODE: string  := "X8";
        PCS_CH0_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH0_ALIGN_MODE: string  := "1GB";
        PCS_CH0_SAMP_16B: string  := "X16";
        PCS_CH0_COMMA_REG0: integer := 0;
        PCS_CH0_COMMA_MASK: integer := 0;
        PCS_CH0_CEB_MODE: string  := "10GB";
        PCS_CH0_CTC_MODE: string  := "1SKIP";
        PCS_CH0_A_REG   : integer := 0;
        PCS_CH0_GE_AUTO_EN: string  := "FALSE";
        PCS_CH0_SKIP_REG0: integer := 0;
        PCS_CH0_SKIP_REG1: integer := 0;
        PCS_CH0_SKIP_REG2: integer := 0;
        PCS_CH0_SKIP_REG3: integer := 0;
        PCS_CH0_DEC_DUAL: string  := "FALSE";
        PCS_CH0_SPLIT   : string  := "FALSE";
        PCS_CH0_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH0_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH0_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH0_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH0_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH0_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_RCLK_POLINV: string  := "RCLK";
        PCS_CH0_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH0_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH0_CB_RCLK_EN: string  := "FALSE";
        PCS_CH0_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH0_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH0_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH0_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH0_SLAVE   : string  := "MASTER";
        PCS_CH0_PCIE_SLAVE: string  := "MASTER";
        PCS_CH0_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH0_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH0_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH0_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH0_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH0_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH0_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH0_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH0_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH0_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH0_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH0_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH0_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH0_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH0_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH0_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH0_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH0_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH0_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH0_TX_SLAVE: string  := "SLAVE";
        PCS_CH0_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH0_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH0_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH0_TX_OUTZZ: string  := "FALSE";
        PCS_CH0_ENC_DUAL: string  := "FALSE";
        PCS_CH0_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH0_COMMA_REG1: integer := 0;
        PCS_CH0_RAPID_IMAX: integer := 0;
        PCS_CH0_RAPID_VMIN_1: integer := 0;
        PCS_CH0_RAPID_VMIN_2: integer := 0;
        PCS_CH0_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH0_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH0_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH0_TX_INSERT_ER: string  := "FALSE";
        PCS_CH0_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH0_ERR_CNT : integer := 0;
        PCS_CH0_DEFAULT_RADDR: integer := 0;
        PCS_CH0_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH0_DELAY_SET: integer := 0;
        PCS_CH0_SEACH_OFFSET: string  := "20BIT";
        PCS_CH0_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH0_CTC_AFULL: integer := 0;
        PCS_CH0_CTC_AEMPTY: integer := 0;
        PCS_CH0_CTC_CONTI_SKP_SET: integer := 0;
        PCS_CH0_FAR_LOOP: string  := "FALSE";
        PCS_CH0_NEAR_LOOP: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH0_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH0_INT_RX_CLR_7: string  := "FALSE";
        PCS_CH0_CA_RX   : integer := 0;
        PCS_CH1_CA_RX   : integer := 0;
        PCS_CH2_CA_RX   : integer := 0;
        PCS_CH3_CA_RX   : integer := 0;
        PCS_CH0_CA_TX   : integer := 0;
        PCS_CH1_CA_TX   : integer := 0;
        PCS_CH2_CA_TX   : integer := 0;
        PCS_CH3_CA_TX   : integer := 0;
        PCS_CH0_CA_DYN_DLY_EN_RX: string  := "FALSE";
        PCS_CH1_CA_DYN_DLY_EN_RX: string  := "FALSE";
        PCS_CH2_CA_DYN_DLY_EN_RX: string  := "FALSE";
        PCS_CH3_CA_DYN_DLY_EN_RX: string  := "FALSE";
        PCS_CH0_CA_DYN_DLY_EN_TX: string  := "FALSE";
        PCS_CH1_CA_DYN_DLY_EN_TX: string  := "FALSE";
        PCS_CH2_CA_DYN_DLY_EN_TX: string  := "FALSE";
        PCS_CH3_CA_DYN_DLY_EN_TX: string  := "FALSE";
        PCS_CH0_CA_DYN_DLY_SEL_RX: string  := "FALSE";
        PCS_CH1_CA_DYN_DLY_SEL_RX: string  := "FALSE";
        PCS_CH2_CA_DYN_DLY_SEL_RX: string  := "FALSE";
        PCS_CH3_CA_DYN_DLY_SEL_RX: string  := "FALSE";
        PCS_CH0_CA_DYN_DLY_SEL_TX: string  := "FALSE";
        PCS_CH1_CA_DYN_DLY_SEL_TX: string  := "FALSE";
        PCS_CH2_CA_DYN_DLY_SEL_TX: string  := "FALSE";
        PCS_CH3_CA_DYN_DLY_SEL_TX: string  := "FALSE";
        PCS_CH0_CA_RSTN_RX: string  := "FALSE";
        PCS_CH1_CA_RSTN_RX: string  := "FALSE";
        PCS_CH2_CA_RSTN_RX: string  := "FALSE";
        PCS_CH3_CA_RSTN_RX: string  := "FALSE";
        PCS_CH0_CA_RSTN_TX: string  := "FALSE";
        PCS_CH1_CA_RSTN_TX: string  := "FALSE";
        PCS_CH2_CA_RSTN_TX: string  := "FALSE";
        PCS_CH3_CA_RSTN_TX: string  := "FALSE";
        PCS_CH1_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH1_BYPASS_DENC: string  := "FALSE";
        PCS_CH1_BYPASS_BONDING: string  := "FALSE";
        PCS_CH1_BYPASS_CTC: string  := "FALSE";
        PCS_CH1_BYPASS_GEAR: string  := "FALSE";
        PCS_CH1_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH1_DATA_MODE: string  := "X8";
        PCS_CH1_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH1_ALIGN_MODE: string  := "1GB";
        PCS_CH1_SAMP_16B: string  := "X16";
        PCS_CH1_COMMA_REG0: integer := 0;
        PCS_CH1_COMMA_MASK: integer := 0;
        PCS_CH1_CEB_MODE: string  := "10GB";
        PCS_CH1_CTC_MODE: string  := "1SKIP";
        PCS_CH1_A_REG   : integer := 0;
        PCS_CH1_GE_AUTO_EN: string  := "FALSE";
        PCS_CH1_SKIP_REG0: integer := 0;
        PCS_CH1_SKIP_REG1: integer := 0;
        PCS_CH1_SKIP_REG2: integer := 0;
        PCS_CH1_SKIP_REG3: integer := 0;
        PCS_CH1_DEC_DUAL: string  := "FALSE";
        PCS_CH1_SPLIT   : string  := "FALSE";
        PCS_CH1_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH1_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH1_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH1_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH1_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH1_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_RCLK_POLINV: string  := "RCLK";
        PCS_CH1_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH1_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH1_CB_RCLK_EN: string  := "FALSE";
        PCS_CH1_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH1_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH1_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH1_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH1_SLAVE   : string  := "MASTER";
        PCS_CH1_PCIE_SLAVE: string  := "MASTER";
        PCS_CH1_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH1_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH1_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH1_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH1_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH1_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH1_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH1_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH1_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH1_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH1_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH1_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH1_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH1_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH1_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH1_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH1_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH1_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH1_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH1_TX_SLAVE: string  := "SLAVE";
        PCS_CH1_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH1_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH1_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH1_TX_OUTZZ: string  := "FALSE";
        PCS_CH1_ENC_DUAL: string  := "FALSE";
        PCS_CH1_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH1_COMMA_REG1: integer := 0;
        PCS_CH1_RAPID_IMAX: integer := 0;
        PCS_CH1_RAPID_VMIN_1: integer := 0;
        PCS_CH1_RAPID_VMIN_2: integer := 0;
        PCS_CH1_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH1_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH1_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH1_TX_INSERT_ER: string  := "FALSE";
        PCS_CH1_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH1_ERR_CNT : integer := 0;
        PCS_CH1_DEFAULT_RADDR: integer := 0;
        PCS_CH1_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH1_DELAY_SET: integer := 0;
        PCS_CH1_SEACH_OFFSET: string  := "20BIT";
        PCS_CH1_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH1_CTC_AFULL: integer := 0;
        PCS_CH1_CTC_AEMPTY: integer := 0;
        PCS_CH1_CTC_CONTI_SKP_SET: integer := 0;
        PCS_CH1_FAR_LOOP: string  := "FALSE";
        PCS_CH1_NEAR_LOOP: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH1_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH1_INT_RX_CLR_7: string  := "FALSE";
        PCS_CH2_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH2_BYPASS_DENC: string  := "FALSE";
        PCS_CH2_BYPASS_BONDING: string  := "FALSE";
        PCS_CH2_BYPASS_CTC: string  := "FALSE";
        PCS_CH2_BYPASS_GEAR: string  := "FALSE";
        PCS_CH2_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH2_DATA_MODE: string  := "X8";
        PCS_CH2_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH2_ALIGN_MODE: string  := "1GB";
        PCS_CH2_SAMP_16B: string  := "X16";
        PCS_CH2_COMMA_REG0: integer := 0;
        PCS_CH2_COMMA_MASK: integer := 0;
        PCS_CH2_CEB_MODE: string  := "10GB";
        PCS_CH2_CTC_MODE: string  := "1SKIP";
        PCS_CH2_A_REG   : integer := 0;
        PCS_CH2_GE_AUTO_EN: string  := "FALSE";
        PCS_CH2_SKIP_REG0: integer := 0;
        PCS_CH2_SKIP_REG1: integer := 0;
        PCS_CH2_SKIP_REG2: integer := 0;
        PCS_CH2_SKIP_REG3: integer := 0;
        PCS_CH2_DEC_DUAL: string  := "FALSE";
        PCS_CH2_SPLIT   : string  := "FALSE";
        PCS_CH2_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH2_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH2_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH2_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH2_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH2_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_RCLK_POLINV: string  := "RCLK";
        PCS_CH2_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH2_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH2_CB_RCLK_EN: string  := "FALSE";
        PCS_CH2_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH2_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH2_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH2_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH2_SLAVE   : string  := "MASTER";
        PCS_CH2_PCIE_SLAVE: string  := "MASTER";
        PCS_CH2_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH2_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH2_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH2_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH2_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH2_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH2_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH2_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH2_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH2_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH2_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH2_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH2_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH2_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH2_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH2_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH2_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH2_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH2_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH2_TX_SLAVE: string  := "SLAVE";
        PCS_CH2_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH2_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH2_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH2_TX_OUTZZ: string  := "FALSE";
        PCS_CH2_ENC_DUAL: string  := "FALSE";
        PCS_CH2_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH2_COMMA_REG1: integer := 0;
        PCS_CH2_RAPID_IMAX: integer := 0;
        PCS_CH2_RAPID_VMIN_1: integer := 0;
        PCS_CH2_RAPID_VMIN_2: integer := 0;
        PCS_CH2_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH2_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH2_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH2_TX_INSERT_ER: string  := "FALSE";
        PCS_CH2_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH2_ERR_CNT : integer := 0;
        PCS_CH2_DEFAULT_RADDR: integer := 0;
        PCS_CH2_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH2_DELAY_SET: integer := 0;
        PCS_CH2_SEACH_OFFSET: string  := "20BIT";
        PCS_CH2_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH2_CTC_AFULL: integer := 0;
        PCS_CH2_CTC_AEMPTY: integer := 0;
        PCS_CH2_CTC_CONTI_SKP_SET: integer := 0;
        PCS_CH2_FAR_LOOP: string  := "FALSE";
        PCS_CH2_NEAR_LOOP: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH2_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH2_INT_RX_CLR_7: string  := "FALSE";
        PCS_CH3_BYPASS_WORD_ALIGN: string  := "FALSE";
        PCS_CH3_BYPASS_DENC: string  := "FALSE";
        PCS_CH3_BYPASS_BONDING: string  := "FALSE";
        PCS_CH3_BYPASS_CTC: string  := "FALSE";
        PCS_CH3_BYPASS_GEAR: string  := "FALSE";
        PCS_CH3_BYPASS_BRIDGE: string  := "FALSE";
        PCS_CH3_DATA_MODE: string  := "X8";
        PCS_CH3_RX_POLARITY_INV: string  := "DELAY";
        PCS_CH3_ALIGN_MODE: string  := "1GB";
        PCS_CH3_SAMP_16B: string  := "X16";
        PCS_CH3_COMMA_REG0: integer := 0;
        PCS_CH3_COMMA_MASK: integer := 0;
        PCS_CH3_CEB_MODE: string  := "10GB";
        PCS_CH3_CTC_MODE: string  := "1SKIP";
        PCS_CH3_A_REG   : integer := 0;
        PCS_CH3_GE_AUTO_EN: string  := "FALSE";
        PCS_CH3_SKIP_REG0: integer := 0;
        PCS_CH3_SKIP_REG1: integer := 0;
        PCS_CH3_SKIP_REG2: integer := 0;
        PCS_CH3_SKIP_REG3: integer := 0;
        PCS_CH3_DEC_DUAL: string  := "FALSE";
        PCS_CH3_SPLIT   : string  := "FALSE";
        PCS_CH3_FIFOFLAG_CTC: string  := "FALSE";
        PCS_CH3_COMMA_DET_MODE: string  := "COMMA_PATTERN";
        PCS_CH3_ERRDETECT_SILENCE: string  := "FALSE";
        PCS_CH3_PMA_RCLK_POLINV: string  := "PMA_RCLK";
        PCS_CH3_PCS_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_MCB_RCLK_POLINV: string  := "MCB_RCLK";
        PCS_CH3_CB_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_AFTER_CTC_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_RCLK_POLINV: string  := "RCLK";
        PCS_CH3_BRIDGE_RCLK_SEL: string  := "PMA_RCLK";
        PCS_CH3_PCS_RCLK_EN: string  := "FALSE";
        PCS_CH3_CB_RCLK_EN: string  := "FALSE";
        PCS_CH3_AFTER_CTC_RCLK_EN: string  := "FALSE";
        PCS_CH3_AFTER_CTC_RCLK_EN_GB: string  := "FALSE";
        PCS_CH3_BRIDGE_RCLK_EN: string  := "FALSE";
        PCS_CH3_PCS_RX_RSTN: string  := "FALSE";
        PCS_CH3_SLAVE   : string  := "MASTER";
        PCS_CH3_PCIE_SLAVE: string  := "MASTER";
        PCS_CH3_PCS_CB_RSTN: string  := "FALSE";
        PCS_CH3_TX_BYPASS_BRIDGE_UINT: string  := "FALSE";
        PCS_CH3_TX_BYPASS_GEAR: string  := "FALSE";
        PCS_CH3_TX_BYPASS_ENC: string  := "FALSE";
        PCS_CH3_TX_BYPASS_BIT_SLIP: string  := "FALSE";
        PCS_CH3_TX_GEAR_SPLIT: string  := "FALSE";
        PCS_CH3_TX_DRIVE_REG_MODE: string  := "NO_CHANGE";
        PCS_CH3_TX_BIT_SLIP_CYCLES: integer := 0;
        PCS_CH3_INT_TX_MASK_0: string  := "FALSE";
        PCS_CH3_INT_TX_MASK_1: string  := "FALSE";
        PCS_CH3_INT_TX_MASK_2: string  := "FALSE";
        PCS_CH3_INT_TX_CLR_0: string  := "FALSE";
        PCS_CH3_INT_TX_CLR_1: string  := "FALSE";
        PCS_CH3_INT_TX_CLR_2: string  := "FALSE";
        PCS_CH3_TX_PMA_TCLK_POLINV: string  := "PMA_TCLK";
        PCS_CH3_TX_PCS_CLK_EN_SEL: string  := "FALSE";
        PCS_CH3_TX_BRIDGE_TCLK_SEL: string  := "PCS_TCLK";
        PCS_CH3_TX_TCLK_POLINV: string  := "TCLK";
        PCS_CH3_TX_PCS_TX_RSTN: string  := "FALSE";
        PCS_CH3_TX_SLAVE: string  := "SLAVE";
        PCS_CH3_TX_BRIDGE_CLK_EN_SEL: string  := "FALSE";
        PCS_CH3_DATA_WIDTH_MODE: string  := "X20";
        PCS_CH3_TX_TCLK2FABRIC_SEL: string  := "FALSE";
        PCS_CH3_TX_OUTZZ: string  := "FALSE";
        PCS_CH3_ENC_DUAL: string  := "FALSE";
        PCS_CH3_TX_BITSLIP_DATA_MODE: string  := "X10";
        PCS_CH3_COMMA_REG1: integer := 0;
        PCS_CH3_RAPID_IMAX: integer := 0;
        PCS_CH3_RAPID_VMIN_1: integer := 0;
        PCS_CH3_RAPID_VMIN_2: integer := 0;
        PCS_CH3_RX_PRBS_MODE: string  := "DISABLE";
        PCS_CH3_RX_ERRCNT_CLR: string  := "FALSE";
        PCS_CH3_TX_PRBS_MODE: string  := "DISABLE";
        PCS_CH3_TX_INSERT_ER: string  := "FALSE";
        PCS_CH3_ENABLE_PRBS_GEN: string  := "FALSE";
        PCS_CH3_ERR_CNT : integer := 0;
        PCS_CH3_DEFAULT_RADDR: integer := 0;
        PCS_CH3_MASTER_CHECK_OFFSET: integer := 0;
        PCS_CH3_DELAY_SET: integer := 0;
        PCS_CH3_SEACH_OFFSET: string  := "20BIT";
        PCS_CH3_CEB_RAPIDLS_MMAX: integer := 0;
        PCS_CH3_CTC_AFULL: integer := 0;
        PCS_CH3_CTC_AEMPTY: integer := 0;
        PCS_CH3_CTC_CONTI_SKP_SET: integer := 0;
        PCS_CH3_FAR_LOOP: string  := "FALSE";
        PCS_CH3_NEAR_LOOP: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_0: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_1: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_2: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_3: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_4: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_5: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_6: string  := "FALSE";
        PCS_CH3_INT_RX_MASK_7: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_0: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_1: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_2: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_3: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_4: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_5: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_6: string  := "FALSE";
        PCS_CH3_INT_RX_CLR_7: string  := "FALSE";
        PMA_CH0_REG_RX_PD: string  := "ON";
        PMA_CH0_REG_RX_PD_EN: string  := "FALSE";
        PMA_CH0_REG_RX_CLKPATH_PD: string  := "ON";
        PMA_CH0_REG_RX_CLKPATH_PD_EN: string  := "FALSE";
        PMA_CH0_REG_RX_DATAPATH_PD: string  := "ON";
        PMA_CH0_REG_RX_DATAPATH_PD_EN: string  := "FALSE";
        PMA_CH0_REG_RX_SIGDET_PD: string  := "ON";
        PMA_CH0_REG_RX_SIGDET_PD_EN: string  := "FALSE";
        PMA_CH0_REG_RX_DCC_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_DCC_RST_N_EN: string  := "FALSE";
        PMA_CH0_REG_RX_CDR_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_CDR_RST_N_EN: string  := "FALSE";
        PMA_CH0_REG_RX_SIGDET_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_SIGDET_RST_N_EN: string  := "FALSE";
        PMA_CH0_REG_RXPCLK_SLIP: string  := "FALSE";
        PMA_CH0_REG_RXPCLK_SLIP_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_PCLKSWITCH_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_PCLKSWITCH_RST_N_EN: string  := "FALSE";
        PMA_CH0_REG_RX_PCLKSWITCH: string  := "FALSE";
        PMA_CH0_REG_RX_PCLKSWITCH_EN: string  := "FALSE";
        PMA_CH0_REG_RX_HIGHZ: string  := "FALSE";
        PMA_CH0_REG_RX_HIGHZ_EN: string  := "FALSE";
        PMA_CH0_REG_RX_EQ_C_SET: integer := 8;
        PMA_CH0_REG_RX_EQ_R_SET: integer := 8;
        PMA_CH0_REG_RX_BUSWIDTH: string  := "20BIT";
        PMA_CH0_REG_RX_BUSWIDTH_EN: string  := "FALSE";
        PMA_CH0_REG_RX_RATE: string  := "DIV1";
        PMA_CH0_REG_RX_RATE_EN: string  := "FALSE";
        PMA_CH0_REG_RX_RES_TRIM: integer := 51;
        PMA_CH0_REG_RX_RES_TRIM_EN: string  := "FALSE";
        PMA_CH0_REG_RX_EQ_OFF: string  := "FALSE";
        PMA_CH0_REG_RX_PREAMP_IC: integer := 1367;
        PMA_CH0_REG_RX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH0_REG_RX_PIBUF_IC: integer := 2;
        PMA_CH0_REG_RX_DCC_IC_RX: integer := 3;
        PMA_CH0_REG_RX_DCC_IC_TX: integer := 3;
        PMA_CH0_REG_RX_ICTRL_TRX: string  := "100PCT";
        PMA_CH0_REG_RX_ICTRL_SIGDET: integer := 5;
        PMA_CH0_REG_RX_ICTRL_PREAMP: string  := "100PCT";
        PMA_CH0_REG_RX_ICTRL_SLICER: string  := "100PCT";
        PMA_CH0_REG_RX_ICTRL_PIBUF: string  := "100PCT";
        PMA_CH0_REG_RX_ICTRL_PI: string  := "100PCT";
        PMA_CH0_REG_RX_ICTRL_DCC: string  := "100PCT";
        PMA_CH0_REG_RX_ICTRL_PREDRV: string  := "100PCT";
        PMA_CH0_REG_TX_RATE: string  := "DIV1";
        PMA_CH0_REG_TX_RATE_EN: string  := "FALSE";
        PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N_EN: string  := "FALSE";
        PMA_CH0_REG_RX_TX2RX_PLPBK_EN: string  := "FALSE";
        PMA_CH0_REG_TXCLK_SEL: string  := "PLL";
        PMA_CH0_REG_RX_DATA_POLARITY: string  := "NORMAL";
        PMA_CH0_REG_RX_ERR_INSERT: string  := "FALSE";
        PMA_CH0_REG_UDP_CHK_EN: string  := "FALSE";
        PMA_CH0_REG_PRBS_SEL: string  := "PRBS7";
        PMA_CH0_REG_PRBS_CHK_EN: string  := "FALSE";
        PMA_CH0_REG_PRBS_CHK_WIDTH_SEL: string  := "20BIT";
        PMA_CH0_REG_BIST_CHK_PAT_SEL: string  := "PRBS";
        PMA_CH0_REG_LOAD_ERR_CNT: string  := "DISABLE";
        PMA_CH0_REG_CHK_COUNTER_EN: string  := "FALSE";
        PMA_CH0_REG_CDR_PROP_GAIN: integer := 2;
        PMA_CH0_REG_CDR_PROP_TURBO_GAIN: integer := 6;
        PMA_CH0_REG_CDR_INT_GAIN: integer := 2;
        PMA_CH0_REG_CDR_INT_TURBO_GAIN: integer := 6;
        PMA_CH0_REG_CDR_INT_SAT_MAX: integer := 992;
        PMA_CH0_REG_CDR_INT_SAT_MIN: integer := 32;
        PMA_CH0_REG_CDR_INT_RST: string  := "FALSE";
        PMA_CH0_REG_CDR_INT_RST_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_PROP_RST: string  := "FALSE";
        PMA_CH0_REG_CDR_PROP_RST_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_LOCK_RST: string  := "FALSE";
        PMA_CH0_REG_CDR_LOCK_RST_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_RX_PI_FORCE_SEL: integer := 0;
        PMA_CH0_REG_CDR_RX_PI_FORCE_D: integer := 0;
        PMA_CH0_REG_CDR_LOCK_TIMER: string  := "1_2U";
        PMA_CH0_REG_CDR_TURBO_MODE_TIMER: integer := 1;
        PMA_CH0_REG_CDR_LOCK_VAL: string  := "FALSE";
        PMA_CH0_REG_CDR_LOCK_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_INT_SAT_DET_EN: string  := "TRUE";
        PMA_CH0_REG_CDR_SAT_DET_STATUS_EN: string  := "FALSE";
        PMA_CH0_REG_CDR_SAT_DET_STATUS_RESET_EN: string  := "FALSE";
        PMA_CH0_REG_CDR_PI_CTRL_RST: string  := "FALSE";
        PMA_CH0_REG_CDR_PI_CTRL_RST_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_SAT_DET_RST: string  := "FALSE";
        PMA_CH0_REG_CDR_SAT_DET_RST_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_SAT_DET_STICKY_RST: string  := "FALSE";
        PMA_CH0_REG_CDR_SAT_DET_STICKY_RST_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_SIGDET_STATUS_DIS: string  := "FALSE";
        PMA_CH0_REG_CDR_SAT_DET_TIMER: integer := 2;
        PMA_CH0_REG_CDR_SAT_DET_STATUS_VAL: string  := "FALSE";
        PMA_CH0_REG_CDR_SAT_DET_STATUS_OW: string  := "DISABLE";
        PMA_CH0_REG_CDR_TURBO_MODE_EN: string  := "TRUE";
        PMA_CH0_REG_CDR_STATUS_RADDR_INIT: integer := 0;
        PMA_CH0_REG_CDR_STATUS_FIFO_EN: string  := "TRUE";
        PMA_CH0_REG_PMA_TEST_SEL: integer := 0;
        PMA_CH0_REG_OOB_COMWAKE_GAP_MIN: integer := 3;
        PMA_CH0_REG_OOB_COMWAKE_GAP_MAX: integer := 11;
        PMA_CH0_REG_OOB_COMINIT_GAP_MIN: integer := 15;
        PMA_CH0_REG_OOB_COMINIT_GAP_MAX: integer := 35;
        PMA_CH0_REG_RX_PIBUF_IC_TX: integer := 1;
        PMA_CH0_REG_COMWAKE_STATUS_CLEAR: integer := 0;
        PMA_CH0_REG_COMINIT_STATUS_CLEAR: integer := 0;
        PMA_CH0_REG_RX_SYNC_RST_N_EN: string  := "FALSE";
        PMA_CH0_REG_RX_SYNC_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_SATA_COMINIT_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_SATA_COMINIT: string  := "FALSE";
        PMA_CH0_REG_RX_SATA_COMWAKE_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_SATA_COMWAKE: string  := "FALSE";
        PMA_CH0_REG_RX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH0_REG_TX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH0_REG_RX_SLIP_SEL_EN: string  := "FALSE";
        PMA_CH0_REG_RX_SLIP_SEL: integer := 0;
        PMA_CH0_REG_RX_SLIP_EN: string  := "FALSE";
        PMA_CH0_REG_RX_SIGDET_STATUS_SEL: integer := 5;
        PMA_CH0_REG_RX_SIGDET_FSM_RST_N: string  := "TRUE";
        PMA_CH0_REG_RX_SIGDET_STATUS_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_SIGDET_STATUS: string  := "FALSE";
        PMA_CH0_REG_RX_SIGDET_VTH: string  := "50MV";
        PMA_CH0_REG_RX_SIGDET_GRM: integer := 0;
        PMA_CH0_REG_RX_SIGDET_PULSE_EXT: string  := "DISABLE";
        PMA_CH0_REG_RX_SIGDET_CH2_SEL: integer := 0;
        PMA_CH0_REG_RX_SIGDET_CH2_CHK_WINDOW: integer := 3;
        PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_EN: string  := "TRUE";
        PMA_CH0_REG_RX_SIGDET_NOSIG_COUNT_SETTING: integer := 4;
        PMA_CH0_REG_RX_SIGDET_OOB_DET_COUNT_VAL: integer := 0;
        PMA_CH0_REG_SLIP_FIFO_INV_EN: string  := "FALSE";
        PMA_CH0_REG_SLIP_FIFO_INV: string  := "POS_EDGE";
        PMA_CH0_REG_RX_SIGDET_4OOB_DET_SEL: integer := 7;
        PMA_CH0_REG_RX_SIGDET_IC_I: integer := 10;
        PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N: string  := "FALSE";
        PMA_CH0_REG_RX_OOB_DETECTOR_PD_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_OOB_DETECTOR_PD: string  := "ON";
        PMA_CH0_REG_RX_TERM_CM_CTRL: string  := "5DIV7";
        PMA_CH0_REG_TX_PD: string  := "ON";
        PMA_CH0_REG_TX_PD_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_CLKPATH_PD: string  := "ON";
        PMA_CH0_REG_TX_CLKPATH_PD_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_BEACON_TIMER_SEL: integer := 0;
        PMA_CH0_REG_TX_RXDET_REQ_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_RXDET_REQ: string  := "FALSE";
        PMA_CH0_REG_TX_BEACON_EN_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_BEACON_EN: string  := "FALSE";
        PMA_CH0_REG_TX_EI_EN_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_EI_EN: string  := "FALSE";
        PMA_CH0_REG_TX_RES_CAL_EN: string  := "FALSE";
        PMA_CH0_REG_TX_RES_CAL: integer := 51;
        PMA_CH0_REG_TX_BIAS_CAL_EN: string  := "FALSE";
        PMA_CH0_REG_TX_BIAS_CTRL: integer := 48;
        PMA_CH0_REG_TX_RXDET_TIMER_SEL: string  := "12CYCLE";
        PMA_CH0_REG_TX_SYNC_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_SYNC: string  := "DISABLE";
        PMA_CH0_REG_TX_PD_POST: string  := "OFF";
        PMA_CH0_REG_TX_PD_POST_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_RESET_N_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_RESET_N: string  := "TRUE";
        PMA_CH0_REG_TX_DCC_RESET_N_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_DCC_RESET_N: string  := "TRUE";
        PMA_CH0_REG_TX_BUSWIDTH_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_BUSWIDTH: string  := "20BIT";
        PMA_CH0_REG_PLL_READY_OW: string  := "DISABLE";
        PMA_CH0_REG_PLL_READY: string  := "TRUE";
        PMA_CH0_REG_TX_PCLK_SW_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_PCLK_SW: string  := "TRUE";
        PMA_CH0_REG_EI_PCLK_DELAY_SEL: integer := 0;
        PMA_CH0_REG_TX_DRV01_DAC0: integer := 0;
        PMA_CH0_REG_TX_DRV01_DAC1: integer := 10;
        PMA_CH0_REG_TX_DRV01_DAC2: integer := 16;
        PMA_CH0_REG_TX_DRV00_DAC0: integer := 63;
        PMA_CH0_REG_TX_DRV00_DAC1: integer := 53;
        PMA_CH0_REG_TX_DRV00_DAC2: integer := 48;
        PMA_CH0_REG_TX_AMP0: integer := 8;
        PMA_CH0_REG_TX_AMP1: integer := 16;
        PMA_CH0_REG_TX_AMP2: integer := 32;
        PMA_CH0_REG_TX_AMP3: integer := 48;
        PMA_CH0_REG_TX_AMP4: integer := 56;
        PMA_CH0_REG_TX_MARGIN: integer := 0;
        PMA_CH0_REG_TX_MARGIN_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_DEEMP: integer := 0;
        PMA_CH0_REG_TX_DEEMP_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_SWING: string  := "FALSE";
        PMA_CH0_REG_TX_SWING_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_RXDET_THRESHOLD: string  := "100MV";
        PMA_CH0_REG_TX_BEACON_OSC_CTRL: integer := 4;
        PMA_CH0_REG_TX_PREDRV_DAC: integer := 1;
        PMA_CH0_REG_TX_PREDRV_CM_CTRL: integer := 1;
        PMA_CH0_REG_TX_TX2RX_SLPBACK_EN: string  := "FALSE";
        PMA_CH0_REG_TX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH0_REG_TX_RXDET_STATUS_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_RXDET_STATUS: string  := "TRUE";
        PMA_CH0_REG_TX_PRBS_GEN_EN: string  := "FALSE";
        PMA_CH0_REG_TX_PRBS_GEN_WIDTH_SEL: string  := "20BIT";
        PMA_CH0_REG_TX_PRBS_SEL: string  := "PRBS7";
        PMA_CH0_REG_TX_UDP_DATA: integer := 256773;
        PMA_CH0_REG_TX_FIFO_RST_N: string  := "FALSE";
        PMA_CH0_REG_TX_FIFO_WP_CTRL: integer := 2;
        PMA_CH0_REG_TX_FIFO_EN: string  := "FALSE";
        PMA_CH0_REG_TX_DATA_MUX_SEL: integer := 2;
        PMA_CH0_REG_TX_ERR_INSERT: string  := "FALSE";
        PMA_CH0_REG_TX_SATA_EN: string  := "FALSE";
        PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON_OW: string  := "DISABLE";
        PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON: string  := "ENABLE";
        PMA_CH0_REG_TX_PULLUP_DAC0: integer := 8;
        PMA_CH0_REG_TX_PULLUP_DAC1: integer := 8;
        PMA_CH0_REG_TX_PULLUP_DAC2: integer := 8;
        PMA_CH0_REG_TX_PULLUP_DAC3: integer := 8;
        PMA_CH0_REG_TX_OOB_DELAY_SEL: integer := 0;
        PMA_CH0_REG_TX_POLARITY: string  := "NORMAL";
        PMA_CH0_REG_TX_SLPBK_AMP: integer := 1;
        PMA_CH0_REG_TX_LS_MODE_EN: string  := "FALSE";
        PMA_CH0_REG_TX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH0_REG_TX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH0_REG_RX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH0_REG_RX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH0_REG_RX_JTAG_OE: string  := "DISABLE";
        PMA_CH0_REG_RX_ACJTAG_VHYSTSE: integer := 0;
        PMA_CH0_REG_TX_FBCLK_FAR_EN: string  := "FALSE";
        PMA_CH0_REG_RX_TERM_MODE_CTRL: integer := 6;
        PMA_CH0_REG_PLPBK_TXPCLK_EN: string  := "TRUE";
        PMA_CH0_CFG_LANE_POWERUP: string  := "OFF";
        PMA_CH0_CFG_PMA_POR_N: string  := "FALSE";
        PMA_CH0_CFG_RX_LANE_POWERUP: string  := "OFF";
        PMA_CH0_CFG_RX_PMA_RSTN: string  := "FALSE";
        PMA_CH0_CFG_TX_LANE_POWERUP: string  := "OFF";
        PMA_CH0_CFG_TX_PMA_RSTN: string  := "FALSE";
        PMA_CH0_REG_RESERVED_48_45: integer := 0;
        PMA_CH0_REG_RESERVED_69: integer := 0;
        PMA_CH0_REG_RESERVED_77_76: integer := 0;
        PMA_CH0_REG_RESERVED_171_164: integer := 0;
        PMA_CH0_REG_RESERVED_175_172: integer := 0;
        PMA_CH0_REG_RESERVED_190: integer := 0;
        PMA_CH0_REG_RESERVED_233_232: integer := 0;
        PMA_CH0_REG_RESERVED_235_234: integer := 0;
        PMA_CH0_REG_RESERVED_241_240: integer := 0;
        PMA_CH0_REG_RESERVED_285_283: integer := 0;
        PMA_CH0_REG_RESERVED_286: integer := 0;
        PMA_CH0_REG_RESERVED_295: integer := 0;
        PMA_CH0_REG_RESERVED_298: integer := 0;
        PMA_CH0_REG_RESERVED_332_325: integer := 0;
        PMA_CH0_REG_RESERVED_340_333: integer := 0;
        PMA_CH0_REG_RESERVED_348_341: integer := 0;
        PMA_CH0_REG_RESERVED_354_349: integer := 0;
        PMA_CH0_REG_RESERVED_373: integer := 0;
        PMA_CH0_REG_RESERVED_376: integer := 0;
        PMA_CH0_REG_RESERVED_452: integer := 0;
        PMA_CH0_REG_RESERVED_502_499: integer := 0;
        PMA_CH0_REG_RESERVED_506_505: integer := 0;
        PMA_CH0_REG_RESERVED_550_549: integer := 0;
        PMA_CH0_REG_RESERVED_556_552: integer := 0;
        PMA_CH1_REG_RX_PD: string  := "ON";
        PMA_CH1_REG_RX_PD_EN: string  := "FALSE";
        PMA_CH1_REG_RX_CLKPATH_PD: string  := "ON";
        PMA_CH1_REG_RX_CLKPATH_PD_EN: string  := "FALSE";
        PMA_CH1_REG_RX_DATAPATH_PD: string  := "ON";
        PMA_CH1_REG_RX_DATAPATH_PD_EN: string  := "FALSE";
        PMA_CH1_REG_RX_SIGDET_PD: string  := "ON";
        PMA_CH1_REG_RX_SIGDET_PD_EN: string  := "FALSE";
        PMA_CH1_REG_RX_DCC_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_DCC_RST_N_EN: string  := "FALSE";
        PMA_CH1_REG_RX_CDR_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_CDR_RST_N_EN: string  := "FALSE";
        PMA_CH1_REG_RX_SIGDET_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_SIGDET_RST_N_EN: string  := "FALSE";
        PMA_CH1_REG_RXPCLK_SLIP: string  := "FALSE";
        PMA_CH1_REG_RXPCLK_SLIP_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_PCLKSWITCH_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_PCLKSWITCH_RST_N_EN: string  := "FALSE";
        PMA_CH1_REG_RX_PCLKSWITCH: string  := "FALSE";
        PMA_CH1_REG_RX_PCLKSWITCH_EN: string  := "FALSE";
        PMA_CH1_REG_RX_HIGHZ: string  := "FALSE";
        PMA_CH1_REG_RX_HIGHZ_EN: string  := "FALSE";
        PMA_CH1_REG_RX_EQ_C_SET: integer := 8;
        PMA_CH1_REG_RX_EQ_R_SET: integer := 8;
        PMA_CH1_REG_RX_BUSWIDTH: string  := "20BIT";
        PMA_CH1_REG_RX_BUSWIDTH_EN: string  := "FALSE";
        PMA_CH1_REG_RX_RATE: string  := "DIV1";
        PMA_CH1_REG_RX_RATE_EN: string  := "FALSE";
        PMA_CH1_REG_RX_RES_TRIM: integer := 51;
        PMA_CH1_REG_RX_RES_TRIM_EN: string  := "FALSE";
        PMA_CH1_REG_RX_EQ_OFF: string  := "FALSE";
        PMA_CH1_REG_RX_PREAMP_IC: integer := 1367;
        PMA_CH1_REG_RX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH1_REG_RX_PIBUF_IC: integer := 2;
        PMA_CH1_REG_RX_DCC_IC_RX: integer := 3;
        PMA_CH1_REG_RX_DCC_IC_TX: integer := 3;
        PMA_CH1_REG_RX_ICTRL_TRX: string  := "100PCT";
        PMA_CH1_REG_RX_ICTRL_SIGDET: integer := 5;
        PMA_CH1_REG_RX_ICTRL_PREAMP: string  := "100PCT";
        PMA_CH1_REG_RX_ICTRL_SLICER: string  := "100PCT";
        PMA_CH1_REG_RX_ICTRL_PIBUF: string  := "100PCT";
        PMA_CH1_REG_RX_ICTRL_PI: string  := "100PCT";
        PMA_CH1_REG_RX_ICTRL_DCC: string  := "100PCT";
        PMA_CH1_REG_RX_ICTRL_PREDRV: string  := "100PCT";
        PMA_CH1_REG_TX_RATE: string  := "DIV1";
        PMA_CH1_REG_TX_RATE_EN: string  := "FALSE";
        PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N_EN: string  := "FALSE";
        PMA_CH1_REG_RX_TX2RX_PLPBK_EN: string  := "FALSE";
        PMA_CH1_REG_TXCLK_SEL: string  := "PLL";
        PMA_CH1_REG_RX_DATA_POLARITY: string  := "NORMAL";
        PMA_CH1_REG_RX_ERR_INSERT: string  := "FALSE";
        PMA_CH1_REG_UDP_CHK_EN: string  := "FALSE";
        PMA_CH1_REG_PRBS_SEL: string  := "PRBS7";
        PMA_CH1_REG_PRBS_CHK_EN: string  := "FALSE";
        PMA_CH1_REG_PRBS_CHK_WIDTH_SEL: string  := "20BIT";
        PMA_CH1_REG_BIST_CHK_PAT_SEL: string  := "PRBS";
        PMA_CH1_REG_LOAD_ERR_CNT: string  := "DISABLE";
        PMA_CH1_REG_CHK_COUNTER_EN: string  := "FALSE";
        PMA_CH1_REG_CDR_PROP_GAIN: integer := 2;
        PMA_CH1_REG_CDR_PROP_TURBO_GAIN: integer := 6;
        PMA_CH1_REG_CDR_INT_GAIN: integer := 2;
        PMA_CH1_REG_CDR_INT_TURBO_GAIN: integer := 6;
        PMA_CH1_REG_CDR_INT_SAT_MAX: integer := 992;
        PMA_CH1_REG_CDR_INT_SAT_MIN: integer := 32;
        PMA_CH1_REG_CDR_INT_RST: string  := "FALSE";
        PMA_CH1_REG_CDR_INT_RST_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_PROP_RST: string  := "FALSE";
        PMA_CH1_REG_CDR_PROP_RST_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_LOCK_RST: string  := "FALSE";
        PMA_CH1_REG_CDR_LOCK_RST_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_RX_PI_FORCE_SEL: integer := 0;
        PMA_CH1_REG_CDR_RX_PI_FORCE_D: integer := 0;
        PMA_CH1_REG_CDR_LOCK_TIMER: string  := "1_2U";
        PMA_CH1_REG_CDR_TURBO_MODE_TIMER: integer := 1;
        PMA_CH1_REG_CDR_LOCK_VAL: string  := "FALSE";
        PMA_CH1_REG_CDR_LOCK_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_INT_SAT_DET_EN: string  := "TRUE";
        PMA_CH1_REG_CDR_SAT_DET_STATUS_EN: string  := "FALSE";
        PMA_CH1_REG_CDR_SAT_DET_STATUS_RESET_EN: string  := "FALSE";
        PMA_CH1_REG_CDR_PI_CTRL_RST: string  := "FALSE";
        PMA_CH1_REG_CDR_PI_CTRL_RST_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_SAT_DET_RST: string  := "FALSE";
        PMA_CH1_REG_CDR_SAT_DET_RST_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_SAT_DET_STICKY_RST: string  := "FALSE";
        PMA_CH1_REG_CDR_SAT_DET_STICKY_RST_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_SIGDET_STATUS_DIS: string  := "FALSE";
        PMA_CH1_REG_CDR_SAT_DET_TIMER: integer := 2;
        PMA_CH1_REG_CDR_SAT_DET_STATUS_VAL: string  := "FALSE";
        PMA_CH1_REG_CDR_SAT_DET_STATUS_OW: string  := "DISABLE";
        PMA_CH1_REG_CDR_TURBO_MODE_EN: string  := "TRUE";
        PMA_CH1_REG_CDR_STATUS_RADDR_INIT: integer := 0;
        PMA_CH1_REG_CDR_STATUS_FIFO_EN: string  := "TRUE";
        PMA_CH1_REG_PMA_TEST_SEL: integer := 0;
        PMA_CH1_REG_OOB_COMWAKE_GAP_MIN: integer := 3;
        PMA_CH1_REG_OOB_COMWAKE_GAP_MAX: integer := 11;
        PMA_CH1_REG_OOB_COMINIT_GAP_MIN: integer := 15;
        PMA_CH1_REG_OOB_COMINIT_GAP_MAX: integer := 35;
        PMA_CH1_REG_RX_PIBUF_IC_TX: integer := 1;
        PMA_CH1_REG_COMWAKE_STATUS_CLEAR: integer := 0;
        PMA_CH1_REG_COMINIT_STATUS_CLEAR: integer := 0;
        PMA_CH1_REG_RX_SYNC_RST_N_EN: string  := "FALSE";
        PMA_CH1_REG_RX_SYNC_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_SATA_COMINIT_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_SATA_COMINIT: string  := "FALSE";
        PMA_CH1_REG_RX_SATA_COMWAKE_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_SATA_COMWAKE: string  := "FALSE";
        PMA_CH1_REG_RX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH1_REG_TX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH1_REG_RX_SLIP_SEL_EN: string  := "FALSE";
        PMA_CH1_REG_RX_SLIP_SEL: integer := 0;
        PMA_CH1_REG_RX_SLIP_EN: string  := "FALSE";
        PMA_CH1_REG_RX_SIGDET_STATUS_SEL: integer := 5;
        PMA_CH1_REG_RX_SIGDET_FSM_RST_N: string  := "TRUE";
        PMA_CH1_REG_RX_SIGDET_STATUS_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_SIGDET_STATUS: string  := "FALSE";
        PMA_CH1_REG_RX_SIGDET_VTH: string  := "50MV";
        PMA_CH1_REG_RX_SIGDET_GRM: integer := 0;
        PMA_CH1_REG_RX_SIGDET_PULSE_EXT: string  := "DISABLE";
        PMA_CH1_REG_RX_SIGDET_CH2_SEL: integer := 0;
        PMA_CH1_REG_RX_SIGDET_CH2_CHK_WINDOW: integer := 3;
        PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_EN: string  := "TRUE";
        PMA_CH1_REG_RX_SIGDET_NOSIG_COUNT_SETTING: integer := 4;
        PMA_CH1_REG_RX_SIGDET_OOB_DET_COUNT_VAL: integer := 0;
        PMA_CH1_REG_SLIP_FIFO_INV_EN: string  := "FALSE";
        PMA_CH1_REG_SLIP_FIFO_INV: string  := "POS_EDGE";
        PMA_CH1_REG_RX_SIGDET_4OOB_DET_SEL: integer := 7;
        PMA_CH1_REG_RX_SIGDET_IC_I: integer := 10;
        PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N: string  := "FALSE";
        PMA_CH1_REG_RX_OOB_DETECTOR_PD_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_OOB_DETECTOR_PD: string  := "ON";
        PMA_CH1_REG_RX_TERM_CM_CTRL: string  := "5DIV7";
        PMA_CH1_REG_TX_PD: string  := "ON";
        PMA_CH1_REG_TX_PD_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_CLKPATH_PD: string  := "ON";
        PMA_CH1_REG_TX_CLKPATH_PD_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_BEACON_TIMER_SEL: integer := 0;
        PMA_CH1_REG_TX_RXDET_REQ_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_RXDET_REQ: string  := "FALSE";
        PMA_CH1_REG_TX_BEACON_EN_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_BEACON_EN: string  := "FALSE";
        PMA_CH1_REG_TX_EI_EN_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_EI_EN: string  := "FALSE";
        PMA_CH1_REG_TX_RES_CAL_EN: string  := "FALSE";
        PMA_CH1_REG_TX_RES_CAL: integer := 51;
        PMA_CH1_REG_TX_BIAS_CAL_EN: string  := "FALSE";
        PMA_CH1_REG_TX_BIAS_CTRL: integer := 48;
        PMA_CH1_REG_TX_RXDET_TIMER_SEL: string  := "12CYCLE";
        PMA_CH1_REG_TX_SYNC_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_SYNC: string  := "DISABLE";
        PMA_CH1_REG_TX_PD_POST: string  := "OFF";
        PMA_CH1_REG_TX_PD_POST_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_RESET_N_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_RESET_N: string  := "TRUE";
        PMA_CH1_REG_TX_DCC_RESET_N_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_DCC_RESET_N: string  := "TRUE";
        PMA_CH1_REG_TX_BUSWIDTH_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_BUSWIDTH: string  := "20BIT";
        PMA_CH1_REG_PLL_READY_OW: string  := "DISABLE";
        PMA_CH1_REG_PLL_READY: string  := "TRUE";
        PMA_CH1_REG_TX_PCLK_SW_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_PCLK_SW: string  := "TRUE";
        PMA_CH1_REG_EI_PCLK_DELAY_SEL: integer := 0;
        PMA_CH1_REG_TX_DRV01_DAC0: integer := 0;
        PMA_CH1_REG_TX_DRV01_DAC1: integer := 10;
        PMA_CH1_REG_TX_DRV01_DAC2: integer := 16;
        PMA_CH1_REG_TX_DRV00_DAC0: integer := 63;
        PMA_CH1_REG_TX_DRV00_DAC1: integer := 53;
        PMA_CH1_REG_TX_DRV00_DAC2: integer := 48;
        PMA_CH1_REG_TX_AMP0: integer := 8;
        PMA_CH1_REG_TX_AMP1: integer := 16;
        PMA_CH1_REG_TX_AMP2: integer := 32;
        PMA_CH1_REG_TX_AMP3: integer := 48;
        PMA_CH1_REG_TX_AMP4: integer := 56;
        PMA_CH1_REG_TX_MARGIN: integer := 0;
        PMA_CH1_REG_TX_MARGIN_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_DEEMP: integer := 0;
        PMA_CH1_REG_TX_DEEMP_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_SWING: string  := "FALSE";
        PMA_CH1_REG_TX_SWING_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_RXDET_THRESHOLD: string  := "100MV";
        PMA_CH1_REG_TX_BEACON_OSC_CTRL: integer := 4;
        PMA_CH1_REG_TX_PREDRV_DAC: integer := 1;
        PMA_CH1_REG_TX_PREDRV_CM_CTRL: integer := 1;
        PMA_CH1_REG_TX_TX2RX_SLPBACK_EN: string  := "FALSE";
        PMA_CH1_REG_TX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH1_REG_TX_RXDET_STATUS_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_RXDET_STATUS: string  := "TRUE";
        PMA_CH1_REG_TX_PRBS_GEN_EN: string  := "FALSE";
        PMA_CH1_REG_TX_PRBS_GEN_WIDTH_SEL: string  := "20BIT";
        PMA_CH1_REG_TX_PRBS_SEL: string  := "PRBS7";
        PMA_CH1_REG_TX_UDP_DATA: integer := 256773;
        PMA_CH1_REG_TX_FIFO_RST_N: string  := "FALSE";
        PMA_CH1_REG_TX_FIFO_WP_CTRL: integer := 2;
        PMA_CH1_REG_TX_FIFO_EN: string  := "FALSE";
        PMA_CH1_REG_TX_DATA_MUX_SEL: integer := 2;
        PMA_CH1_REG_TX_ERR_INSERT: string  := "FALSE";
        PMA_CH1_REG_TX_SATA_EN: string  := "FALSE";
        PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON_OW: string  := "DISABLE";
        PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON: string  := "ENABLE";
        PMA_CH1_REG_TX_PULLUP_DAC0: integer := 8;
        PMA_CH1_REG_TX_PULLUP_DAC1: integer := 8;
        PMA_CH1_REG_TX_PULLUP_DAC2: integer := 8;
        PMA_CH1_REG_TX_PULLUP_DAC3: integer := 8;
        PMA_CH1_REG_TX_OOB_DELAY_SEL: integer := 0;
        PMA_CH1_REG_TX_POLARITY: string  := "NORMAL";
        PMA_CH1_REG_TX_SLPBK_AMP: integer := 1;
        PMA_CH1_REG_TX_LS_MODE_EN: string  := "FALSE";
        PMA_CH1_REG_TX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH1_REG_TX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH1_REG_RX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH1_REG_RX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH1_REG_RX_JTAG_OE: string  := "DISABLE";
        PMA_CH1_REG_RX_ACJTAG_VHYSTSE: integer := 0;
        PMA_CH1_REG_TX_FBCLK_FAR_EN: string  := "FALSE";
        PMA_CH1_REG_RX_TERM_MODE_CTRL: integer := 6;
        PMA_CH1_REG_PLPBK_TXPCLK_EN: string  := "TRUE";
        PMA_CH1_CFG_LANE_POWERUP: string  := "OFF";
        PMA_CH1_CFG_PMA_POR_N: string  := "FALSE";
        PMA_CH1_CFG_RX_LANE_POWERUP: string  := "OFF";
        PMA_CH1_CFG_RX_PMA_RSTN: string  := "FALSE";
        PMA_CH1_CFG_TX_LANE_POWERUP: string  := "OFF";
        PMA_CH1_CFG_TX_PMA_RSTN: string  := "FALSE";
        PMA_CH1_REG_RESERVED_48_45: integer := 0;
        PMA_CH1_REG_RESERVED_69: integer := 0;
        PMA_CH1_REG_RESERVED_77_76: integer := 0;
        PMA_CH1_REG_RESERVED_171_164: integer := 0;
        PMA_CH1_REG_RESERVED_175_172: integer := 0;
        PMA_CH1_REG_RESERVED_190: integer := 0;
        PMA_CH1_REG_RESERVED_233_232: integer := 0;
        PMA_CH1_REG_RESERVED_235_234: integer := 0;
        PMA_CH1_REG_RESERVED_241_240: integer := 0;
        PMA_CH1_REG_RESERVED_285_283: integer := 0;
        PMA_CH1_REG_RESERVED_286: integer := 0;
        PMA_CH1_REG_RESERVED_295: integer := 0;
        PMA_CH1_REG_RESERVED_298: integer := 0;
        PMA_CH1_REG_RESERVED_332_325: integer := 0;
        PMA_CH1_REG_RESERVED_340_333: integer := 0;
        PMA_CH1_REG_RESERVED_348_341: integer := 0;
        PMA_CH1_REG_RESERVED_354_349: integer := 0;
        PMA_CH1_REG_RESERVED_373: integer := 0;
        PMA_CH1_REG_RESERVED_376: integer := 0;
        PMA_CH1_REG_RESERVED_452: integer := 0;
        PMA_CH1_REG_RESERVED_502_499: integer := 0;
        PMA_CH1_REG_RESERVED_506_505: integer := 0;
        PMA_CH1_REG_RESERVED_550_549: integer := 0;
        PMA_CH1_REG_RESERVED_556_552: integer := 0;
        PMA_CH2_REG_RX_PD: string  := "ON";
        PMA_CH2_REG_RX_PD_EN: string  := "FALSE";
        PMA_CH2_REG_RX_CLKPATH_PD: string  := "ON";
        PMA_CH2_REG_RX_CLKPATH_PD_EN: string  := "FALSE";
        PMA_CH2_REG_RX_DATAPATH_PD: string  := "ON";
        PMA_CH2_REG_RX_DATAPATH_PD_EN: string  := "FALSE";
        PMA_CH2_REG_RX_SIGDET_PD: string  := "ON";
        PMA_CH2_REG_RX_SIGDET_PD_EN: string  := "FALSE";
        PMA_CH2_REG_RX_DCC_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_DCC_RST_N_EN: string  := "FALSE";
        PMA_CH2_REG_RX_CDR_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_CDR_RST_N_EN: string  := "FALSE";
        PMA_CH2_REG_RX_SIGDET_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_SIGDET_RST_N_EN: string  := "FALSE";
        PMA_CH2_REG_RXPCLK_SLIP: string  := "FALSE";
        PMA_CH2_REG_RXPCLK_SLIP_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_PCLKSWITCH_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_PCLKSWITCH_RST_N_EN: string  := "FALSE";
        PMA_CH2_REG_RX_PCLKSWITCH: string  := "FALSE";
        PMA_CH2_REG_RX_PCLKSWITCH_EN: string  := "FALSE";
        PMA_CH2_REG_RX_HIGHZ: string  := "FALSE";
        PMA_CH2_REG_RX_HIGHZ_EN: string  := "FALSE";
        PMA_CH2_REG_RX_EQ_C_SET: integer := 8;
        PMA_CH2_REG_RX_EQ_R_SET: integer := 8;
        PMA_CH2_REG_RX_BUSWIDTH: string  := "20BIT";
        PMA_CH2_REG_RX_BUSWIDTH_EN: string  := "FALSE";
        PMA_CH2_REG_RX_RATE: string  := "DIV1";
        PMA_CH2_REG_RX_RATE_EN: string  := "FALSE";
        PMA_CH2_REG_RX_RES_TRIM: integer := 51;
        PMA_CH2_REG_RX_RES_TRIM_EN: string  := "FALSE";
        PMA_CH2_REG_RX_EQ_OFF: string  := "FALSE";
        PMA_CH2_REG_RX_PREAMP_IC: integer := 1367;
        PMA_CH2_REG_RX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH2_REG_RX_PIBUF_IC: integer := 2;
        PMA_CH2_REG_RX_DCC_IC_RX: integer := 3;
        PMA_CH2_REG_RX_DCC_IC_TX: integer := 3;
        PMA_CH2_REG_RX_ICTRL_TRX: string  := "100PCT";
        PMA_CH2_REG_RX_ICTRL_SIGDET: integer := 5;
        PMA_CH2_REG_RX_ICTRL_PREAMP: string  := "100PCT";
        PMA_CH2_REG_RX_ICTRL_SLICER: string  := "100PCT";
        PMA_CH2_REG_RX_ICTRL_PIBUF: string  := "100PCT";
        PMA_CH2_REG_RX_ICTRL_PI: string  := "100PCT";
        PMA_CH2_REG_RX_ICTRL_DCC: string  := "100PCT";
        PMA_CH2_REG_RX_ICTRL_PREDRV: string  := "100PCT";
        PMA_CH2_REG_TX_RATE: string  := "DIV1";
        PMA_CH2_REG_TX_RATE_EN: string  := "FALSE";
        PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N_EN: string  := "FALSE";
        PMA_CH2_REG_RX_TX2RX_PLPBK_EN: string  := "FALSE";
        PMA_CH2_REG_TXCLK_SEL: string  := "PLL";
        PMA_CH2_REG_RX_DATA_POLARITY: string  := "NORMAL";
        PMA_CH2_REG_RX_ERR_INSERT: string  := "FALSE";
        PMA_CH2_REG_UDP_CHK_EN: string  := "FALSE";
        PMA_CH2_REG_PRBS_SEL: string  := "PRBS7";
        PMA_CH2_REG_PRBS_CHK_EN: string  := "FALSE";
        PMA_CH2_REG_PRBS_CHK_WIDTH_SEL: string  := "20BIT";
        PMA_CH2_REG_BIST_CHK_PAT_SEL: string  := "PRBS";
        PMA_CH2_REG_LOAD_ERR_CNT: string  := "DISABLE";
        PMA_CH2_REG_CHK_COUNTER_EN: string  := "FALSE";
        PMA_CH2_REG_CDR_PROP_GAIN: integer := 2;
        PMA_CH2_REG_CDR_PROP_TURBO_GAIN: integer := 6;
        PMA_CH2_REG_CDR_INT_GAIN: integer := 2;
        PMA_CH2_REG_CDR_INT_TURBO_GAIN: integer := 6;
        PMA_CH2_REG_CDR_INT_SAT_MAX: integer := 992;
        PMA_CH2_REG_CDR_INT_SAT_MIN: integer := 32;
        PMA_CH2_REG_CDR_INT_RST: string  := "FALSE";
        PMA_CH2_REG_CDR_INT_RST_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_PROP_RST: string  := "FALSE";
        PMA_CH2_REG_CDR_PROP_RST_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_LOCK_RST: string  := "FALSE";
        PMA_CH2_REG_CDR_LOCK_RST_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_RX_PI_FORCE_SEL: integer := 0;
        PMA_CH2_REG_CDR_RX_PI_FORCE_D: integer := 0;
        PMA_CH2_REG_CDR_LOCK_TIMER: string  := "1_2U";
        PMA_CH2_REG_CDR_TURBO_MODE_TIMER: integer := 1;
        PMA_CH2_REG_CDR_LOCK_VAL: string  := "FALSE";
        PMA_CH2_REG_CDR_LOCK_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_INT_SAT_DET_EN: string  := "TRUE";
        PMA_CH2_REG_CDR_SAT_DET_STATUS_EN: string  := "FALSE";
        PMA_CH2_REG_CDR_SAT_DET_STATUS_RESET_EN: string  := "FALSE";
        PMA_CH2_REG_CDR_PI_CTRL_RST: string  := "FALSE";
        PMA_CH2_REG_CDR_PI_CTRL_RST_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_SAT_DET_RST: string  := "FALSE";
        PMA_CH2_REG_CDR_SAT_DET_RST_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_SAT_DET_STICKY_RST: string  := "FALSE";
        PMA_CH2_REG_CDR_SAT_DET_STICKY_RST_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_SIGDET_STATUS_DIS: string  := "FALSE";
        PMA_CH2_REG_CDR_SAT_DET_TIMER: integer := 2;
        PMA_CH2_REG_CDR_SAT_DET_STATUS_VAL: string  := "FALSE";
        PMA_CH2_REG_CDR_SAT_DET_STATUS_OW: string  := "DISABLE";
        PMA_CH2_REG_CDR_TURBO_MODE_EN: string  := "TRUE";
        PMA_CH2_REG_CDR_STATUS_RADDR_INIT: integer := 0;
        PMA_CH2_REG_CDR_STATUS_FIFO_EN: string  := "TRUE";
        PMA_CH2_REG_PMA_TEST_SEL: integer := 0;
        PMA_CH2_REG_OOB_COMWAKE_GAP_MIN: integer := 3;
        PMA_CH2_REG_OOB_COMWAKE_GAP_MAX: integer := 11;
        PMA_CH2_REG_OOB_COMINIT_GAP_MIN: integer := 15;
        PMA_CH2_REG_OOB_COMINIT_GAP_MAX: integer := 35;
        PMA_CH2_REG_RX_PIBUF_IC_TX: integer := 1;
        PMA_CH2_REG_COMWAKE_STATUS_CLEAR: integer := 0;
        PMA_CH2_REG_COMINIT_STATUS_CLEAR: integer := 0;
        PMA_CH2_REG_RX_SYNC_RST_N_EN: string  := "FALSE";
        PMA_CH2_REG_RX_SYNC_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_SATA_COMINIT_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_SATA_COMINIT: string  := "FALSE";
        PMA_CH2_REG_RX_SATA_COMWAKE_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_SATA_COMWAKE: string  := "FALSE";
        PMA_CH2_REG_RX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH2_REG_TX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH2_REG_RX_SLIP_SEL_EN: string  := "FALSE";
        PMA_CH2_REG_RX_SLIP_SEL: integer := 0;
        PMA_CH2_REG_RX_SLIP_EN: string  := "FALSE";
        PMA_CH2_REG_RX_SIGDET_STATUS_SEL: integer := 5;
        PMA_CH2_REG_RX_SIGDET_FSM_RST_N: string  := "TRUE";
        PMA_CH2_REG_RX_SIGDET_STATUS_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_SIGDET_STATUS: string  := "FALSE";
        PMA_CH2_REG_RX_SIGDET_VTH: string  := "50MV";
        PMA_CH2_REG_RX_SIGDET_GRM: integer := 0;
        PMA_CH2_REG_RX_SIGDET_PULSE_EXT: string  := "DISABLE";
        PMA_CH2_REG_RX_SIGDET_CH2_SEL: integer := 0;
        PMA_CH2_REG_RX_SIGDET_CH2_CHK_WINDOW: integer := 3;
        PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_EN: string  := "TRUE";
        PMA_CH2_REG_RX_SIGDET_NOSIG_COUNT_SETTING: integer := 4;
        PMA_CH2_REG_RX_SIGDET_OOB_DET_COUNT_VAL: integer := 0;
        PMA_CH2_REG_SLIP_FIFO_INV_EN: string  := "FALSE";
        PMA_CH2_REG_SLIP_FIFO_INV: string  := "POS_EDGE";
        PMA_CH2_REG_RX_SIGDET_4OOB_DET_SEL: integer := 7;
        PMA_CH2_REG_RX_SIGDET_IC_I: integer := 10;
        PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N: string  := "FALSE";
        PMA_CH2_REG_RX_OOB_DETECTOR_PD_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_OOB_DETECTOR_PD: string  := "ON";
        PMA_CH2_REG_RX_TERM_CM_CTRL: string  := "5DIV7";
        PMA_CH2_REG_TX_PD: string  := "ON";
        PMA_CH2_REG_TX_PD_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_CLKPATH_PD: string  := "ON";
        PMA_CH2_REG_TX_CLKPATH_PD_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_BEACON_TIMER_SEL: integer := 0;
        PMA_CH2_REG_TX_RXDET_REQ_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_RXDET_REQ: string  := "FALSE";
        PMA_CH2_REG_TX_BEACON_EN_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_BEACON_EN: string  := "FALSE";
        PMA_CH2_REG_TX_EI_EN_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_EI_EN: string  := "FALSE";
        PMA_CH2_REG_TX_RES_CAL_EN: string  := "FALSE";
        PMA_CH2_REG_TX_RES_CAL: integer := 51;
        PMA_CH2_REG_TX_BIAS_CAL_EN: string  := "FALSE";
        PMA_CH2_REG_TX_BIAS_CTRL: integer := 48;
        PMA_CH2_REG_TX_RXDET_TIMER_SEL: string  := "12CYCLE";
        PMA_CH2_REG_TX_SYNC_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_SYNC: string  := "DISABLE";
        PMA_CH2_REG_TX_PD_POST: string  := "OFF";
        PMA_CH2_REG_TX_PD_POST_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_RESET_N_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_RESET_N: string  := "TRUE";
        PMA_CH2_REG_TX_DCC_RESET_N_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_DCC_RESET_N: string  := "TRUE";
        PMA_CH2_REG_TX_BUSWIDTH_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_BUSWIDTH: string  := "20BIT";
        PMA_CH2_REG_PLL_READY_OW: string  := "DISABLE";
        PMA_CH2_REG_PLL_READY: string  := "TRUE";
        PMA_CH2_REG_TX_PCLK_SW_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_PCLK_SW: string  := "TRUE";
        PMA_CH2_REG_EI_PCLK_DELAY_SEL: integer := 0;
        PMA_CH2_REG_TX_DRV01_DAC0: integer := 0;
        PMA_CH2_REG_TX_DRV01_DAC1: integer := 10;
        PMA_CH2_REG_TX_DRV01_DAC2: integer := 16;
        PMA_CH2_REG_TX_DRV00_DAC0: integer := 63;
        PMA_CH2_REG_TX_DRV00_DAC1: integer := 53;
        PMA_CH2_REG_TX_DRV00_DAC2: integer := 48;
        PMA_CH2_REG_TX_AMP0: integer := 8;
        PMA_CH2_REG_TX_AMP1: integer := 16;
        PMA_CH2_REG_TX_AMP2: integer := 32;
        PMA_CH2_REG_TX_AMP3: integer := 48;
        PMA_CH2_REG_TX_AMP4: integer := 56;
        PMA_CH2_REG_TX_MARGIN: integer := 0;
        PMA_CH2_REG_TX_MARGIN_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_DEEMP: integer := 0;
        PMA_CH2_REG_TX_DEEMP_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_SWING: string  := "FALSE";
        PMA_CH2_REG_TX_SWING_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_RXDET_THRESHOLD: string  := "100MV";
        PMA_CH2_REG_TX_BEACON_OSC_CTRL: integer := 4;
        PMA_CH2_REG_TX_PREDRV_DAC: integer := 1;
        PMA_CH2_REG_TX_PREDRV_CM_CTRL: integer := 1;
        PMA_CH2_REG_TX_TX2RX_SLPBACK_EN: string  := "FALSE";
        PMA_CH2_REG_TX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH2_REG_TX_RXDET_STATUS_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_RXDET_STATUS: string  := "TRUE";
        PMA_CH2_REG_TX_PRBS_GEN_EN: string  := "FALSE";
        PMA_CH2_REG_TX_PRBS_GEN_WIDTH_SEL: string  := "20BIT";
        PMA_CH2_REG_TX_PRBS_SEL: string  := "PRBS7";
        PMA_CH2_REG_TX_UDP_DATA: integer := 256773;
        PMA_CH2_REG_TX_FIFO_RST_N: string  := "FALSE";
        PMA_CH2_REG_TX_FIFO_WP_CTRL: integer := 2;
        PMA_CH2_REG_TX_FIFO_EN: string  := "FALSE";
        PMA_CH2_REG_TX_DATA_MUX_SEL: integer := 2;
        PMA_CH2_REG_TX_ERR_INSERT: string  := "FALSE";
        PMA_CH2_REG_TX_SATA_EN: string  := "FALSE";
        PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON_OW: string  := "DISABLE";
        PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON: string  := "ENABLE";
        PMA_CH2_REG_TX_PULLUP_DAC0: integer := 8;
        PMA_CH2_REG_TX_PULLUP_DAC1: integer := 8;
        PMA_CH2_REG_TX_PULLUP_DAC2: integer := 8;
        PMA_CH2_REG_TX_PULLUP_DAC3: integer := 8;
        PMA_CH2_REG_TX_OOB_DELAY_SEL: integer := 0;
        PMA_CH2_REG_TX_POLARITY: string  := "NORMAL";
        PMA_CH2_REG_TX_SLPBK_AMP: integer := 1;
        PMA_CH2_REG_TX_LS_MODE_EN: string  := "FALSE";
        PMA_CH2_REG_TX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH2_REG_TX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH2_REG_RX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH2_REG_RX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH2_REG_RX_JTAG_OE: string  := "DISABLE";
        PMA_CH2_REG_RX_ACJTAG_VHYSTSE: integer := 0;
        PMA_CH2_REG_TX_FBCLK_FAR_EN: string  := "FALSE";
        PMA_CH2_REG_RX_TERM_MODE_CTRL: integer := 6;
        PMA_CH2_REG_PLPBK_TXPCLK_EN: string  := "TRUE";
        PMA_CH2_CFG_LANE_POWERUP: string  := "OFF";
        PMA_CH2_CFG_PMA_POR_N: string  := "FALSE";
        PMA_CH2_CFG_RX_LANE_POWERUP: string  := "OFF";
        PMA_CH2_CFG_RX_PMA_RSTN: string  := "FALSE";
        PMA_CH2_CFG_TX_LANE_POWERUP: string  := "OFF";
        PMA_CH2_CFG_TX_PMA_RSTN: string  := "FALSE";
        PMA_CH2_REG_RESERVED_48_45: integer := 0;
        PMA_CH2_REG_RESERVED_69: integer := 0;
        PMA_CH2_REG_RESERVED_77_76: integer := 0;
        PMA_CH2_REG_RESERVED_171_164: integer := 0;
        PMA_CH2_REG_RESERVED_175_172: integer := 0;
        PMA_CH2_REG_RESERVED_190: integer := 0;
        PMA_CH2_REG_RESERVED_233_232: integer := 0;
        PMA_CH2_REG_RESERVED_235_234: integer := 0;
        PMA_CH2_REG_RESERVED_241_240: integer := 0;
        PMA_CH2_REG_RESERVED_285_283: integer := 0;
        PMA_CH2_REG_RESERVED_286: integer := 0;
        PMA_CH2_REG_RESERVED_295: integer := 0;
        PMA_CH2_REG_RESERVED_298: integer := 0;
        PMA_CH2_REG_RESERVED_332_325: integer := 0;
        PMA_CH2_REG_RESERVED_340_333: integer := 0;
        PMA_CH2_REG_RESERVED_348_341: integer := 0;
        PMA_CH2_REG_RESERVED_354_349: integer := 0;
        PMA_CH2_REG_RESERVED_373: integer := 0;
        PMA_CH2_REG_RESERVED_376: integer := 0;
        PMA_CH2_REG_RESERVED_452: integer := 0;
        PMA_CH2_REG_RESERVED_502_499: integer := 0;
        PMA_CH2_REG_RESERVED_506_505: integer := 0;
        PMA_CH2_REG_RESERVED_550_549: integer := 0;
        PMA_CH2_REG_RESERVED_556_552: integer := 0;
        PMA_CH3_REG_RX_PD: string  := "ON";
        PMA_CH3_REG_RX_PD_EN: string  := "FALSE";
        PMA_CH3_REG_RX_CLKPATH_PD: string  := "ON";
        PMA_CH3_REG_RX_CLKPATH_PD_EN: string  := "FALSE";
        PMA_CH3_REG_RX_DATAPATH_PD: string  := "ON";
        PMA_CH3_REG_RX_DATAPATH_PD_EN: string  := "FALSE";
        PMA_CH3_REG_RX_SIGDET_PD: string  := "ON";
        PMA_CH3_REG_RX_SIGDET_PD_EN: string  := "FALSE";
        PMA_CH3_REG_RX_DCC_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_DCC_RST_N_EN: string  := "FALSE";
        PMA_CH3_REG_RX_CDR_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_CDR_RST_N_EN: string  := "FALSE";
        PMA_CH3_REG_RX_SIGDET_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_SIGDET_RST_N_EN: string  := "FALSE";
        PMA_CH3_REG_RXPCLK_SLIP: string  := "FALSE";
        PMA_CH3_REG_RXPCLK_SLIP_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_PCLKSWITCH_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_PCLKSWITCH_RST_N_EN: string  := "FALSE";
        PMA_CH3_REG_RX_PCLKSWITCH: string  := "FALSE";
        PMA_CH3_REG_RX_PCLKSWITCH_EN: string  := "FALSE";
        PMA_CH3_REG_RX_HIGHZ: string  := "FALSE";
        PMA_CH3_REG_RX_HIGHZ_EN: string  := "FALSE";
        PMA_CH3_REG_RX_EQ_C_SET: integer := 8;
        PMA_CH3_REG_RX_EQ_R_SET: integer := 8;
        PMA_CH3_REG_RX_BUSWIDTH: string  := "20BIT";
        PMA_CH3_REG_RX_BUSWIDTH_EN: string  := "FALSE";
        PMA_CH3_REG_RX_RATE: string  := "DIV1";
        PMA_CH3_REG_RX_RATE_EN: string  := "FALSE";
        PMA_CH3_REG_RX_RES_TRIM: integer := 51;
        PMA_CH3_REG_RX_RES_TRIM_EN: string  := "FALSE";
        PMA_CH3_REG_RX_EQ_OFF: string  := "FALSE";
        PMA_CH3_REG_RX_PREAMP_IC: integer := 1367;
        PMA_CH3_REG_RX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH3_REG_RX_PIBUF_IC: integer := 2;
        PMA_CH3_REG_RX_DCC_IC_RX: integer := 3;
        PMA_CH3_REG_RX_DCC_IC_TX: integer := 3;
        PMA_CH3_REG_RX_ICTRL_TRX: string  := "100PCT";
        PMA_CH3_REG_RX_ICTRL_SIGDET: integer := 5;
        PMA_CH3_REG_RX_ICTRL_PREAMP: string  := "100PCT";
        PMA_CH3_REG_RX_ICTRL_SLICER: string  := "100PCT";
        PMA_CH3_REG_RX_ICTRL_PIBUF: string  := "100PCT";
        PMA_CH3_REG_RX_ICTRL_PI: string  := "100PCT";
        PMA_CH3_REG_RX_ICTRL_DCC: string  := "100PCT";
        PMA_CH3_REG_RX_ICTRL_PREDRV: string  := "100PCT";
        PMA_CH3_REG_TX_RATE: string  := "DIV1";
        PMA_CH3_REG_TX_RATE_EN: string  := "FALSE";
        PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N_EN: string  := "FALSE";
        PMA_CH3_REG_RX_TX2RX_PLPBK_EN: string  := "FALSE";
        PMA_CH3_REG_TXCLK_SEL: string  := "PLL";
        PMA_CH3_REG_RX_DATA_POLARITY: string  := "NORMAL";
        PMA_CH3_REG_RX_ERR_INSERT: string  := "FALSE";
        PMA_CH3_REG_UDP_CHK_EN: string  := "FALSE";
        PMA_CH3_REG_PRBS_SEL: string  := "PRBS7";
        PMA_CH3_REG_PRBS_CHK_EN: string  := "FALSE";
        PMA_CH3_REG_PRBS_CHK_WIDTH_SEL: string  := "20BIT";
        PMA_CH3_REG_BIST_CHK_PAT_SEL: string  := "PRBS";
        PMA_CH3_REG_LOAD_ERR_CNT: string  := "DISABLE";
        PMA_CH3_REG_CHK_COUNTER_EN: string  := "FALSE";
        PMA_CH3_REG_CDR_PROP_GAIN: integer := 2;
        PMA_CH3_REG_CDR_PROP_TURBO_GAIN: integer := 6;
        PMA_CH3_REG_CDR_INT_GAIN: integer := 2;
        PMA_CH3_REG_CDR_INT_TURBO_GAIN: integer := 6;
        PMA_CH3_REG_CDR_INT_SAT_MAX: integer := 992;
        PMA_CH3_REG_CDR_INT_SAT_MIN: integer := 32;
        PMA_CH3_REG_CDR_INT_RST: string  := "FALSE";
        PMA_CH3_REG_CDR_INT_RST_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_PROP_RST: string  := "FALSE";
        PMA_CH3_REG_CDR_PROP_RST_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_LOCK_RST: string  := "FALSE";
        PMA_CH3_REG_CDR_LOCK_RST_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_RX_PI_FORCE_SEL: integer := 0;
        PMA_CH3_REG_CDR_RX_PI_FORCE_D: integer := 0;
        PMA_CH3_REG_CDR_LOCK_TIMER: string  := "1_2U";
        PMA_CH3_REG_CDR_TURBO_MODE_TIMER: integer := 1;
        PMA_CH3_REG_CDR_LOCK_VAL: string  := "FALSE";
        PMA_CH3_REG_CDR_LOCK_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_INT_SAT_DET_EN: string  := "TRUE";
        PMA_CH3_REG_CDR_SAT_DET_STATUS_EN: string  := "FALSE";
        PMA_CH3_REG_CDR_SAT_DET_STATUS_RESET_EN: string  := "FALSE";
        PMA_CH3_REG_CDR_PI_CTRL_RST: string  := "FALSE";
        PMA_CH3_REG_CDR_PI_CTRL_RST_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_SAT_DET_RST: string  := "FALSE";
        PMA_CH3_REG_CDR_SAT_DET_RST_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_SAT_DET_STICKY_RST: string  := "FALSE";
        PMA_CH3_REG_CDR_SAT_DET_STICKY_RST_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_SIGDET_STATUS_DIS: string  := "FALSE";
        PMA_CH3_REG_CDR_SAT_DET_TIMER: integer := 2;
        PMA_CH3_REG_CDR_SAT_DET_STATUS_VAL: string  := "FALSE";
        PMA_CH3_REG_CDR_SAT_DET_STATUS_OW: string  := "DISABLE";
        PMA_CH3_REG_CDR_TURBO_MODE_EN: string  := "TRUE";
        PMA_CH3_REG_CDR_STATUS_RADDR_INIT: integer := 0;
        PMA_CH3_REG_CDR_STATUS_FIFO_EN: string  := "TRUE";
        PMA_CH3_REG_PMA_TEST_SEL: integer := 0;
        PMA_CH3_REG_OOB_COMWAKE_GAP_MIN: integer := 3;
        PMA_CH3_REG_OOB_COMWAKE_GAP_MAX: integer := 11;
        PMA_CH3_REG_OOB_COMINIT_GAP_MIN: integer := 15;
        PMA_CH3_REG_OOB_COMINIT_GAP_MAX: integer := 35;
        PMA_CH3_REG_RX_PIBUF_IC_TX: integer := 1;
        PMA_CH3_REG_COMWAKE_STATUS_CLEAR: integer := 0;
        PMA_CH3_REG_COMINIT_STATUS_CLEAR: integer := 0;
        PMA_CH3_REG_RX_SYNC_RST_N_EN: string  := "FALSE";
        PMA_CH3_REG_RX_SYNC_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_SATA_COMINIT_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_SATA_COMINIT: string  := "FALSE";
        PMA_CH3_REG_RX_SATA_COMWAKE_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_SATA_COMWAKE: string  := "FALSE";
        PMA_CH3_REG_RX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH3_REG_TX_DCC_DISABLE: string  := "ENABLE";
        PMA_CH3_REG_RX_SLIP_SEL_EN: string  := "FALSE";
        PMA_CH3_REG_RX_SLIP_SEL: integer := 0;
        PMA_CH3_REG_RX_SLIP_EN: string  := "FALSE";
        PMA_CH3_REG_RX_SIGDET_STATUS_SEL: integer := 5;
        PMA_CH3_REG_RX_SIGDET_FSM_RST_N: string  := "TRUE";
        PMA_CH3_REG_RX_SIGDET_STATUS_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_SIGDET_STATUS: string  := "FALSE";
        PMA_CH3_REG_RX_SIGDET_VTH: string  := "50MV";
        PMA_CH3_REG_RX_SIGDET_GRM: integer := 0;
        PMA_CH3_REG_RX_SIGDET_PULSE_EXT: string  := "DISABLE";
        PMA_CH3_REG_RX_SIGDET_CH2_SEL: integer := 0;
        PMA_CH3_REG_RX_SIGDET_CH2_CHK_WINDOW: integer := 3;
        PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_EN: string  := "TRUE";
        PMA_CH3_REG_RX_SIGDET_NOSIG_COUNT_SETTING: integer := 4;
        PMA_CH3_REG_RX_SIGDET_OOB_DET_COUNT_VAL: integer := 0;
        PMA_CH3_REG_SLIP_FIFO_INV_EN: string  := "FALSE";
        PMA_CH3_REG_SLIP_FIFO_INV: string  := "POS_EDGE";
        PMA_CH3_REG_RX_SIGDET_4OOB_DET_SEL: integer := 7;
        PMA_CH3_REG_RX_SIGDET_IC_I: integer := 10;
        PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N: string  := "FALSE";
        PMA_CH3_REG_RX_OOB_DETECTOR_PD_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_OOB_DETECTOR_PD: string  := "ON";
        PMA_CH3_REG_RX_TERM_CM_CTRL: string  := "5DIV7";
        PMA_CH3_REG_TX_PD: string  := "ON";
        PMA_CH3_REG_TX_PD_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_CLKPATH_PD: string  := "ON";
        PMA_CH3_REG_TX_CLKPATH_PD_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_BEACON_TIMER_SEL: integer := 0;
        PMA_CH3_REG_TX_RXDET_REQ_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_RXDET_REQ: string  := "FALSE";
        PMA_CH3_REG_TX_BEACON_EN_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_BEACON_EN: string  := "FALSE";
        PMA_CH3_REG_TX_EI_EN_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_EI_EN: string  := "FALSE";
        PMA_CH3_REG_TX_RES_CAL_EN: string  := "FALSE";
        PMA_CH3_REG_TX_RES_CAL: integer := 51;
        PMA_CH3_REG_TX_BIAS_CAL_EN: string  := "FALSE";
        PMA_CH3_REG_TX_BIAS_CTRL: integer := 48;
        PMA_CH3_REG_TX_RXDET_TIMER_SEL: string  := "12CYCLE";
        PMA_CH3_REG_TX_SYNC_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_SYNC: string  := "DISABLE";
        PMA_CH3_REG_TX_PD_POST: string  := "OFF";
        PMA_CH3_REG_TX_PD_POST_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_RESET_N_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_RESET_N: string  := "TRUE";
        PMA_CH3_REG_TX_DCC_RESET_N_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_DCC_RESET_N: string  := "TRUE";
        PMA_CH3_REG_TX_BUSWIDTH_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_BUSWIDTH: string  := "20BIT";
        PMA_CH3_REG_PLL_READY_OW: string  := "DISABLE";
        PMA_CH3_REG_PLL_READY: string  := "TRUE";
        PMA_CH3_REG_TX_PCLK_SW_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_PCLK_SW: string  := "TRUE";
        PMA_CH3_REG_EI_PCLK_DELAY_SEL: integer := 0;
        PMA_CH3_REG_TX_DRV01_DAC0: integer := 0;
        PMA_CH3_REG_TX_DRV01_DAC1: integer := 10;
        PMA_CH3_REG_TX_DRV01_DAC2: integer := 16;
        PMA_CH3_REG_TX_DRV00_DAC0: integer := 63;
        PMA_CH3_REG_TX_DRV00_DAC1: integer := 53;
        PMA_CH3_REG_TX_DRV00_DAC2: integer := 48;
        PMA_CH3_REG_TX_AMP0: integer := 8;
        PMA_CH3_REG_TX_AMP1: integer := 16;
        PMA_CH3_REG_TX_AMP2: integer := 32;
        PMA_CH3_REG_TX_AMP3: integer := 48;
        PMA_CH3_REG_TX_AMP4: integer := 56;
        PMA_CH3_REG_TX_MARGIN: integer := 0;
        PMA_CH3_REG_TX_MARGIN_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_DEEMP: integer := 0;
        PMA_CH3_REG_TX_DEEMP_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_SWING: string  := "FALSE";
        PMA_CH3_REG_TX_SWING_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_RXDET_THRESHOLD: string  := "100MV";
        PMA_CH3_REG_TX_BEACON_OSC_CTRL: integer := 4;
        PMA_CH3_REG_TX_PREDRV_DAC: integer := 1;
        PMA_CH3_REG_TX_PREDRV_CM_CTRL: integer := 1;
        PMA_CH3_REG_TX_TX2RX_SLPBACK_EN: string  := "FALSE";
        PMA_CH3_REG_TX_PCLK_EDGE_SEL: string  := "POS_EDGE";
        PMA_CH3_REG_TX_RXDET_STATUS_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_RXDET_STATUS: string  := "TRUE";
        PMA_CH3_REG_TX_PRBS_GEN_EN: string  := "FALSE";
        PMA_CH3_REG_TX_PRBS_GEN_WIDTH_SEL: string  := "20BIT";
        PMA_CH3_REG_TX_PRBS_SEL: string  := "PRBS7";
        PMA_CH3_REG_TX_UDP_DATA: integer := 256773;
        PMA_CH3_REG_TX_FIFO_RST_N: string  := "FALSE";
        PMA_CH3_REG_TX_FIFO_WP_CTRL: integer := 2;
        PMA_CH3_REG_TX_FIFO_EN: string  := "FALSE";
        PMA_CH3_REG_TX_DATA_MUX_SEL: integer := 2;
        PMA_CH3_REG_TX_ERR_INSERT: string  := "FALSE";
        PMA_CH3_REG_TX_SATA_EN: string  := "FALSE";
        PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON_OW: string  := "DISABLE";
        PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON: string  := "ENABLE";
        PMA_CH3_REG_TX_PULLUP_DAC0: integer := 8;
        PMA_CH3_REG_TX_PULLUP_DAC1: integer := 8;
        PMA_CH3_REG_TX_PULLUP_DAC2: integer := 8;
        PMA_CH3_REG_TX_PULLUP_DAC3: integer := 8;
        PMA_CH3_REG_TX_OOB_DELAY_SEL: integer := 0;
        PMA_CH3_REG_TX_POLARITY: string  := "NORMAL";
        PMA_CH3_REG_TX_SLPBK_AMP: integer := 1;
        PMA_CH3_REG_TX_LS_MODE_EN: string  := "FALSE";
        PMA_CH3_REG_TX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH3_REG_TX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH3_REG_RX_JTAG_MODE_EN_OW: string  := "DISABLE";
        PMA_CH3_REG_RX_JTAG_MODE_EN: string  := "FALSE";
        PMA_CH3_REG_RX_JTAG_OE: string  := "DISABLE";
        PMA_CH3_REG_RX_ACJTAG_VHYSTSE: integer := 0;
        PMA_CH3_REG_TX_FBCLK_FAR_EN: string  := "FALSE";
        PMA_CH3_REG_RX_TERM_MODE_CTRL: integer := 6;
        PMA_CH3_REG_PLPBK_TXPCLK_EN: string  := "TRUE";
        PMA_CH3_CFG_LANE_POWERUP: string  := "OFF";
        PMA_CH3_CFG_PMA_POR_N: string  := "FALSE";
        PMA_CH3_CFG_RX_LANE_POWERUP: string  := "OFF";
        PMA_CH3_CFG_RX_PMA_RSTN: string  := "FALSE";
        PMA_CH3_CFG_TX_LANE_POWERUP: string  := "OFF";
        PMA_CH3_CFG_TX_PMA_RSTN: string  := "FALSE";
        PMA_CH3_REG_RESERVED_48_45: integer := 0;
        PMA_CH3_REG_RESERVED_69: integer := 0;
        PMA_CH3_REG_RESERVED_77_76: integer := 0;
        PMA_CH3_REG_RESERVED_171_164: integer := 0;
        PMA_CH3_REG_RESERVED_175_172: integer := 0;
        PMA_CH3_REG_RESERVED_190: integer := 0;
        PMA_CH3_REG_RESERVED_233_232: integer := 0;
        PMA_CH3_REG_RESERVED_235_234: integer := 0;
        PMA_CH3_REG_RESERVED_241_240: integer := 0;
        PMA_CH3_REG_RESERVED_285_283: integer := 0;
        PMA_CH3_REG_RESERVED_286: integer := 0;
        PMA_CH3_REG_RESERVED_295: integer := 0;
        PMA_CH3_REG_RESERVED_298: integer := 0;
        PMA_CH3_REG_RESERVED_332_325: integer := 0;
        PMA_CH3_REG_RESERVED_340_333: integer := 0;
        PMA_CH3_REG_RESERVED_348_341: integer := 0;
        PMA_CH3_REG_RESERVED_354_349: integer := 0;
        PMA_CH3_REG_RESERVED_373: integer := 0;
        PMA_CH3_REG_RESERVED_376: integer := 0;
        PMA_CH3_REG_RESERVED_452: integer := 0;
        PMA_CH3_REG_RESERVED_502_499: integer := 0;
        PMA_CH3_REG_RESERVED_506_505: integer := 0;
        PMA_CH3_REG_RESERVED_550_549: integer := 0;
        PMA_CH3_REG_RESERVED_556_552: integer := 0;
        PMA_PLL0_REG_PLL_POWERDOWN_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_POWERDOWN: string  := "ON";
        PMA_PLL0_REG_PLL_RESET_N_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_RESET_N: string  := "TRUE";
        PMA_PLL0_REG_PLL_READY_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_READY: string  := "FALSE";
        PMA_PLL0_REG_LANE_SYNC_OW: string  := "DISABLE";
        PMA_PLL0_REG_LANE_SYNC: string  := "FALSE";
        PMA_PLL0_REG_LOCKDET_REPEAT: string  := "DISABLE";
        PMA_PLL0_REG_RESCAL_I_CODE_PMA: string  := "DISABLE";
        PMA_PLL0_REG_RESCAL_RESET_N_OW: string  := "DISABLE";
        PMA_PLL0_REG_RESCAL_RESET_N: string  := "FALSE";
        PMA_PLL0_REG_RESCAL_DONE_OW: string  := "DISABLE";
        PMA_PLL0_REG_RESCAL_DONE: string  := "FALSE";
        PMA_PLL0_REG_RESCAL_CODE_OW: string  := "DISABLE";
        PMA_PLL0_REG_LDO_VREF_SEL: integer := 2;
        PMA_PLL0_REG_BIAS_VCOREP_C: integer := 1;
        PMA_PLL0_REG_RESCAL_I_CODE: integer := 32;
        PMA_PLL0_REG_RESCAL_ONCHIP_SMALL_OW: string  := "DISABLE";
        PMA_PLL0_REG_RESCAL_ONCHIP_SMALL: integer := 0;
        PMA_PLL0_REG_JTAG_OE: string  := "DISABLE";
        PMA_PLL0_REG_JTAG_AC_MODE: string  := "DISABLE";
        PMA_PLL0_REG_JTAG_VHYSTSEL: integer := 0;
        PMA_PLL0_REG_PLL_LOCKDET_EN_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_LOCKDET_EN: string  := "FALSE";
        PMA_PLL0_REG_PLL_LOCKDET_RESET_N_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_LOCKDET_RESET_N: string  := "FALSE";
        PMA_PLL0_REG_PLL_LOCKED_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_LOCKED: string  := "FALSE";
        PMA_PLL0_REG_PLL_LOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL0_REG_PLL_UNLOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL0_REG_NOFBCLK_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL0_REG_PLL_LOCKDET_REFCT: integer := 7;
        PMA_PLL0_REG_PLL_LOCKDET_FBCT: integer := 7;
        PMA_PLL0_REG_PLL_LOCKDET_LOCKCT: integer := 4;
        PMA_PLL0_REG_PLL_LOCKDET_ITER: integer := 3;
        PMA_PLL0_REG_PLL_UNLOCKDET_ITER: integer := 2;
        PMA_PLL0_REG_PD_VCO: string  := "ON";
        PMA_PLL0_REG_FBCLK_TEST_EN: string  := "FALSE";
        PMA_PLL0_REG_REFCLK_TEST_EN: string  := "FALSE";
        PMA_PLL0_REG_TEST_SEL: integer := 0;
        PMA_PLL0_REG_TEST_V_EN: string  := "FALSE";
        PMA_PLL0_REG_TEST_SIG_HALF_EN: string  := "FALSE";
        PMA_PLL0_REG_TEST_FSM: integer := 0;
        PMA_PLL0_REG_REFCLK_OUT_PD: string  := "OFF";
        PMA_PLL0_REG_BGR_STARTUP_EN: string  := "FALSE";
        PMA_PLL0_REG_BGR_STARTUP: string  := "FALSE";
        PMA_PLL0_REG_PD_BGR: string  := "ON";
        PMA_PLL0_REG_REFCLK_TERM_VCM_EN: string  := "TRUE";
        PMA_PLL0_REG_FBDIVA_5_EN: string  := "TRUE";
        PMA_PLL0_REG_FBDIVB: integer := 1;
        PMA_PLL0_REG_RESET_N_PFDQP_OW: string  := "DISABLE";
        PMA_PLL0_REG_RESET_N_PFDQP: string  := "FALSE";
        PMA_PLL0_REG_QPCURRENT: integer := 12;
        PMA_PLL0_REG_VC_FORCE_EN: string  := "FALSE";
        PMA_PLL0_REG_VCRESET_C_RING: integer := 24;
        PMA_PLL0_REG_LPF_R_C: integer := 0;
        PMA_PLL0_REG_LPF_TR_C: integer := 2;
        PMA_PLL0_REG_PD_BIAS: string  := "ON";
        PMA_PLL0_REG_ICTRL_PLL: integer := 1;
        PMA_PLL0_REG_BIAS_QP: integer := 1;
        PMA_PLL0_REG_BIAS_LANE_SYNC: integer := 1;
        PMA_PLL0_REG_BIAS_CLKBUFS1: integer := 1;
        PMA_PLL0_REG_TXPCLK_SEL: integer := 0;
        PMA_PLL0_REG_BIAS_CLKBUFS3: integer := 1;
        PMA_PLL0_REG_LANE_SYNC_EN: string  := "FALSE";
        PMA_PLL0_REG_LANE_SYNC_EN_OW: string  := "DISABLE";
        PMA_PLL0_REG_BIAS_D2S: integer := 1;
        PMA_PLL0_REG_BIAS_REFD2S_C: integer := 1;
        PMA_PLL0_REG_BIAS_VCRST_C: integer := 1;
        PMA_PLL0_REG_BIAS_REFBUF_C: integer := 1;
        PMA_PLL0_REG_CLKBUFS1_C: integer := 1;
        PMA_PLL0_REG_CLKBUFS2_C: integer := 6;
        PMA_PLL0_REG_CLKBUFS3_C: integer := 6;
        PMA_PLL0_REG_CLKBUFS4_C: integer := 1;
        PMA_PLL0_REG_PLL_REFCLK_CML_SEL: integer := 0;
        PMA_PLL0_REG_REFCLK_SEL: string  := "FALSE";
        PMA_PLL0_REG_RESCAL_R_CODE_SIGN: string  := "TRUE";
        PMA_PLL0_REG_PLL_UNLOCKED_OW: string  := "DISABLE";
        PMA_PLL0_REG_PLL_UNLOCKED: string  := "FALSE";
        PMA_PLL0_REG_PLL_LOCKDET_MODE: string  := "FALSE";
        PMA_PLL0_REG_PLL_CLKBUF_PD_LEFT: string  := "ON";
        PMA_PLL0_REG_PLL_CLKBUF_PD_RIGHT: string  := "ON";
        PMA_PLL0_REG_RESCAL_EN: string  := "FALSE";
        PMA_PLL0_REG_RESCAL_I_CODE_VAL: integer := 0;
        PMA_PLL0_REG_RESCAL_I_CODE_OW: integer := 0;
        PMA_PLL0_REG_RESCAL_ITER_VALID_SEL: integer := 0;
        PMA_PLL0_REG_RESCAL_WAIT_SEL: integer := 0;
        PMA_PLL0_REG_I_CTRL_MAX: integer := 45;
        PMA_PLL0_REG_I_CTRL_MIN: integer := 19;
        PARM_CFG_HSST_RSTN: string  := "FALSE";
        PARM_PLL0_POWERUP: string  := "OFF";
        PARM_PLL0_RSTN  : string  := "FALSE";
        PMA_PLL1_REG_PLL_POWERDOWN_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_POWERDOWN: string  := "ON";
        PMA_PLL1_REG_PLL_RESET_N_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_RESET_N: string  := "TRUE";
        PMA_PLL1_REG_PLL_READY_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_READY: string  := "FALSE";
        PMA_PLL1_REG_LANE_SYNC_OW: string  := "DISABLE";
        PMA_PLL1_REG_LANE_SYNC: string  := "FALSE";
        PMA_PLL1_REG_LOCKDET_REPEAT: string  := "DISABLE";
        PMA_PLL1_REG_RESCAL_I_CODE_PMA: string  := "DISABLE";
        PMA_PLL1_REG_RESCAL_RESET_N_OW: string  := "DISABLE";
        PMA_PLL1_REG_RESCAL_RESET_N: string  := "FALSE";
        PMA_PLL1_REG_RESCAL_DONE_OW: string  := "DISABLE";
        PMA_PLL1_REG_RESCAL_DONE: string  := "FALSE";
        PMA_PLL1_REG_RESCAL_CODE_OW: string  := "DISABLE";
        PMA_PLL1_REG_LDO_VREF_SEL: integer := 2;
        PMA_PLL1_REG_BIAS_VCOREP_C: integer := 1;
        PMA_PLL1_REG_RESCAL_I_CODE: integer := 32;
        PMA_PLL1_REG_RESCAL_ONCHIP_SMALL_OW: string  := "DISABLE";
        PMA_PLL1_REG_RESCAL_ONCHIP_SMALL: integer := 0;
        PMA_PLL1_REG_JTAG_OE: string  := "DISABLE";
        PMA_PLL1_REG_JTAG_AC_MODE: string  := "DISABLE";
        PMA_PLL1_REG_JTAG_VHYSTSEL: integer := 0;
        PMA_PLL1_REG_PLL_LOCKDET_EN_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_LOCKDET_EN: string  := "FALSE";
        PMA_PLL1_REG_PLL_LOCKDET_RESET_N_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_LOCKDET_RESET_N: string  := "FALSE";
        PMA_PLL1_REG_PLL_LOCKED_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_LOCKED: string  := "FALSE";
        PMA_PLL1_REG_PLL_LOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL1_REG_PLL_UNLOCKED_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL1_REG_NOFBCLK_STICKY_CLEAR: string  := "FALSE";
        PMA_PLL1_REG_PLL_LOCKDET_REFCT: integer := 7;
        PMA_PLL1_REG_PLL_LOCKDET_FBCT: integer := 7;
        PMA_PLL1_REG_PLL_LOCKDET_LOCKCT: integer := 4;
        PMA_PLL1_REG_PLL_LOCKDET_ITER: integer := 3;
        PMA_PLL1_REG_PLL_UNLOCKDET_ITER: integer := 2;
        PMA_PLL1_REG_PD_VCO: string  := "ON";
        PMA_PLL1_REG_FBCLK_TEST_EN: string  := "FALSE";
        PMA_PLL1_REG_REFCLK_TEST_EN: string  := "FALSE";
        PMA_PLL1_REG_TEST_SEL: integer := 0;
        PMA_PLL1_REG_TEST_V_EN: string  := "FALSE";
        PMA_PLL1_REG_TEST_SIG_HALF_EN: string  := "FALSE";
        PMA_PLL1_REG_TEST_FSM: integer := 0;
        PMA_PLL1_REG_REFCLK_OUT_PD: string  := "OFF";
        PMA_PLL1_REG_BGR_STARTUP_EN: string  := "FALSE";
        PMA_PLL1_REG_BGR_STARTUP: string  := "FALSE";
        PMA_PLL1_REG_PD_BGR: string  := "ON";
        PMA_PLL1_REG_REFCLK_TERM_VCM_EN: string  := "TRUE";
        PMA_PLL1_REG_FBDIVA_5_EN: string  := "TRUE";
        PMA_PLL1_REG_FBDIVB: integer := 1;
        PMA_PLL1_REG_RESET_N_PFDQP_OW: string  := "DISABLE";
        PMA_PLL1_REG_RESET_N_PFDQP: string  := "FALSE";
        PMA_PLL1_REG_QPCURRENT: integer := 12;
        PMA_PLL1_REG_VC_FORCE_EN: string  := "FALSE";
        PMA_PLL1_REG_VCRESET_C_RING: integer := 24;
        PMA_PLL1_REG_LPF_R_C: integer := 0;
        PMA_PLL1_REG_LPF_TR_C: integer := 2;
        PMA_PLL1_REG_PD_BIAS: string  := "ON";
        PMA_PLL1_REG_ICTRL_PLL: integer := 1;
        PMA_PLL1_REG_BIAS_QP: integer := 1;
        PMA_PLL1_REG_BIAS_LANE_SYNC: integer := 1;
        PMA_PLL1_REG_BIAS_CLKBUFS1: integer := 1;
        PMA_PLL1_REG_TXPCLK_SEL: integer := 0;
        PMA_PLL1_REG_BIAS_CLKBUFS3: integer := 1;
        PMA_PLL1_REG_LANE_SYNC_EN: string  := "FALSE";
        PMA_PLL1_REG_LANE_SYNC_EN_OW: string  := "DISABLE";
        PMA_PLL1_REG_BIAS_D2S: integer := 1;
        PMA_PLL1_REG_BIAS_REFD2S_C: integer := 1;
        PMA_PLL1_REG_BIAS_VCRST_C: integer := 1;
        PMA_PLL1_REG_BIAS_REFBUF_C: integer := 1;
        PMA_PLL1_REG_CLKBUFS1_C: integer := 1;
        PMA_PLL1_REG_CLKBUFS2_C: integer := 6;
        PMA_PLL1_REG_CLKBUFS3_C: integer := 6;
        PMA_PLL1_REG_CLKBUFS4_C: integer := 1;
        PMA_PLL1_REG_PLL_REFCLK_CML_SEL: integer := 0;
        PMA_PLL1_REG_REFCLK_SEL: string  := "FALSE";
        PMA_PLL1_REG_RESCAL_R_CODE_SIGN: string  := "TRUE";
        PMA_PLL1_REG_PLL_UNLOCKED_OW: string  := "DISABLE";
        PMA_PLL1_REG_PLL_UNLOCKED: string  := "FALSE";
        PMA_PLL1_REG_PLL_LOCKDET_MODE: string  := "FALSE";
        PMA_PLL1_REG_PLL_CLKBUF_PD_LEFT: string  := "ON";
        PMA_PLL1_REG_PLL_CLKBUF_PD_RIGHT: string  := "ON";
        PMA_PLL1_REG_RESCAL_EN: string  := "FALSE";
        PMA_PLL1_REG_RESCAL_I_CODE_VAL: integer := 0;
        PMA_PLL1_REG_RESCAL_I_CODE_OW: integer := 0;
        PMA_PLL1_REG_RESCAL_ITER_VALID_SEL: integer := 0;
        PMA_PLL1_REG_RESCAL_WAIT_SEL: integer := 0;
        PMA_PLL1_REG_I_CTRL_MAX: integer := 45;
        PMA_PLL1_REG_I_CTRL_MIN: integer := 19;
        PARM_PLL1_POWERUP: string  := "OFF";
        PARM_PLL1_RSTN  : string  := "FALSE";
        PARM_GRSN_DIS   : string  := "FALSE";
        PARM_CFG_RSTN   : string  := "FALSE"
    );
    port(
        P_REFCLKP_0     : in     vl_logic;
        P_REFCLKN_0     : in     vl_logic;
        P_PLL_TEST_0    : out    vl_logic;
        P_REFCLKP_1     : in     vl_logic;
        P_REFCLKN_1     : in     vl_logic;
        P_PLL_TEST_1    : out    vl_logic;
        P_RX_SDP0       : in     vl_logic;
        P_RX_SDN0       : in     vl_logic;
        P_TX_SDP0       : out    vl_logic;
        P_TX_SDN0       : out    vl_logic;
        P_RX_SDP1       : in     vl_logic;
        P_RX_SDN1       : in     vl_logic;
        P_TX_SDP1       : out    vl_logic;
        P_TX_SDN1       : out    vl_logic;
        P_RX_SDP2       : in     vl_logic;
        P_RX_SDN2       : in     vl_logic;
        P_TX_SDP2       : out    vl_logic;
        P_TX_SDN2       : out    vl_logic;
        P_RX_SDP3       : in     vl_logic;
        P_RX_SDN3       : in     vl_logic;
        P_TX_SDP3       : out    vl_logic;
        P_TX_SDN3       : out    vl_logic;
        P_RX0_CLK_FR_CORE: in     vl_logic;
        P_RX1_CLK_FR_CORE: in     vl_logic;
        P_RX2_CLK_FR_CORE: in     vl_logic;
        P_RX3_CLK_FR_CORE: in     vl_logic;
        P_TX0_CLK_FR_CORE: in     vl_logic;
        P_TX1_CLK_FR_CORE: in     vl_logic;
        P_TX2_CLK_FR_CORE: in     vl_logic;
        P_TX3_CLK_FR_CORE: in     vl_logic;
        P_HSST_RST      : in     vl_logic;
        P_PCS_RX_RST_0  : in     vl_logic;
        P_PCS_RX_RST_1  : in     vl_logic;
        P_PCS_RX_RST_2  : in     vl_logic;
        P_PCS_RX_RST_3  : in     vl_logic;
        P_PCS_TX_RST_0  : in     vl_logic;
        P_PCS_TX_RST_1  : in     vl_logic;
        P_PCS_TX_RST_2  : in     vl_logic;
        P_PCS_TX_RST_3  : in     vl_logic;
        P_CFG_CLK       : in     vl_logic;
        P_CFG_RST       : in     vl_logic;
        P_CFG_ENABLE    : in     vl_logic;
        P_CFG_WRITE     : in     vl_logic;
        P_CFG_ADDR      : in     vl_logic_vector(15 downto 0);
        P_CFG_WDATA     : in     vl_logic_vector(7 downto 0);
        P_TDATA_0       : in     vl_logic_vector(44 downto 0);
        P_TDATA_1       : in     vl_logic_vector(44 downto 0);
        P_TDATA_2       : in     vl_logic_vector(44 downto 0);
        P_TDATA_3       : in     vl_logic_vector(44 downto 0);
        P_PCS_WORD_ALIGN_EN: in     vl_logic_vector(3 downto 0);
        P_RX_POLARITY_INVERT: in     vl_logic_vector(3 downto 0);
        P_CEB_ADETECT_EN: in     vl_logic_vector(3 downto 0);
        P_PCS_MCB_EXT_EN: in     vl_logic_vector(3 downto 0);
        P_PCS_NEAREND_LOOP: in     vl_logic_vector(3 downto 0);
        P_PCS_FAREND_LOOP: in     vl_logic_vector(3 downto 0);
        P_CFG_READY     : out    vl_logic;
        P_CFG_RDATA     : out    vl_logic_vector(7 downto 0);
        P_CFG_INT       : out    vl_logic;
        P_PCS_RX_MCB_STATUS: out    vl_logic_vector(3 downto 0);
        P_PCS_LSM_SYNCED: out    vl_logic_vector(3 downto 0);
        P_RDATA_0       : out    vl_logic_vector(46 downto 0);
        P_RDATA_1       : out    vl_logic_vector(46 downto 0);
        P_RDATA_2       : out    vl_logic_vector(46 downto 0);
        P_RDATA_3       : out    vl_logic_vector(46 downto 0);
        P_RCLK2FABRIC   : out    vl_logic_vector(3 downto 0);
        P_TCLK2FABRIC   : out    vl_logic_vector(3 downto 0);
        P_RESCAL_RST_I  : in     vl_logic;
        P_RESCAL_I_CODE_I: in     vl_logic_vector(5 downto 0);
        P_RESCAL_I_CODE_O: out    vl_logic_vector(5 downto 0);
        P_REFCK2CORE_0  : out    vl_logic;
        P_PLL_REF_CLK_0 : in     vl_logic;
        P_PLL_RST_0     : in     vl_logic;
        P_PLLPOWERDOWN_0: in     vl_logic;
        P_PLL_READY_0   : out    vl_logic;
        P_LANE_SYNC_0   : in     vl_logic;
        P_LANE_SYNC_EN_0: in     vl_logic;
        P_RATE_CHANGE_TCLK_ON_0: in     vl_logic;
        P_REFCK2CORE_1  : out    vl_logic;
        P_PLL_REF_CLK_1 : in     vl_logic;
        P_PLL_RST_1     : in     vl_logic;
        P_PLLPOWERDOWN_1: in     vl_logic;
        P_PLL_READY_1   : out    vl_logic;
        P_LANE_SYNC_1   : in     vl_logic;
        P_LANE_SYNC_EN_1: in     vl_logic;
        P_RATE_CHANGE_TCLK_ON_1: in     vl_logic;
        P_LANE_PD_0     : in     vl_logic;
        P_LANE_RST_0    : in     vl_logic;
        P_RX_LANE_PD_0  : in     vl_logic;
        P_RX_PMA_RST_0  : in     vl_logic;
        P_RX_SIGDET_STATUS_0: out    vl_logic;
        P_RX_SATA_COMINIT_0: out    vl_logic;
        P_RX_SATA_COMWAKE_0: out    vl_logic;
        P_RX_LS_DATA_0  : out    vl_logic;
        P_RX_READY_0    : out    vl_logic;
        P_TEST_STATUS_0 : out    vl_logic_vector(19 downto 0);
        P_TX_DEEMP_0    : in     vl_logic_vector(1 downto 0);
        P_TX_LS_DATA_0  : in     vl_logic;
        P_TX_BEACON_EN_0: in     vl_logic;
        P_TX_SWING_0    : in     vl_logic;
        P_TX_RXDET_REQ_0: in     vl_logic;
        P_TX_RATE_0     : in     vl_logic_vector(2 downto 0);
        P_TX_BUSWIDTH_0 : in     vl_logic_vector(2 downto 0);
        P_TX_MARGIN_0   : in     vl_logic_vector(2 downto 0);
        P_TX_RXDET_STATUS_0: out    vl_logic;
        P_TX_PMA_RST_0  : in     vl_logic;
        P_TX_LANE_PD_0  : in     vl_logic;
        P_RX_RATE_0     : in     vl_logic_vector(2 downto 0);
        P_RX_BUSWIDTH_0 : in     vl_logic_vector(2 downto 0);
        P_RX_HIGHZ_0    : in     vl_logic;
        P_CA_ALIGN_RX   : out    vl_logic_vector(3 downto 0);
        P_CA_ALIGN_TX   : out    vl_logic_vector(3 downto 0);
        P_CIM_CLK_ALIGNER_RX0: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_ALIGNER_TX0: in     vl_logic_vector(7 downto 0);
        P_CIM_DYN_DLY_SEL_RX0: in     vl_logic;
        P_CIM_DYN_DLY_SEL_TX0: in     vl_logic;
        P_CIM_START_ALIGN_RX0: in     vl_logic;
        P_CIM_START_ALIGN_TX0: in     vl_logic;
        P_LANE_PD_1     : in     vl_logic;
        P_LANE_RST_1    : in     vl_logic;
        P_RX_LANE_PD_1  : in     vl_logic;
        P_RX_PMA_RST_1  : in     vl_logic;
        P_RX_SIGDET_STATUS_1: out    vl_logic;
        P_RX_SATA_COMINIT_1: out    vl_logic;
        P_RX_SATA_COMWAKE_1: out    vl_logic;
        P_RX_LS_DATA_1  : out    vl_logic;
        P_RX_READY_1    : out    vl_logic;
        P_TEST_STATUS_1 : out    vl_logic_vector(19 downto 0);
        P_TX_DEEMP_1    : in     vl_logic_vector(1 downto 0);
        P_TX_LS_DATA_1  : in     vl_logic;
        P_TX_BEACON_EN_1: in     vl_logic;
        P_TX_SWING_1    : in     vl_logic;
        P_TX_RXDET_REQ_1: in     vl_logic;
        P_TX_RATE_1     : in     vl_logic_vector(2 downto 0);
        P_TX_BUSWIDTH_1 : in     vl_logic_vector(2 downto 0);
        P_TX_MARGIN_1   : in     vl_logic_vector(2 downto 0);
        P_TX_RXDET_STATUS_1: out    vl_logic;
        P_TX_PMA_RST_1  : in     vl_logic;
        P_TX_LANE_PD_1  : in     vl_logic;
        P_RX_RATE_1     : in     vl_logic_vector(2 downto 0);
        P_RX_BUSWIDTH_1 : in     vl_logic_vector(2 downto 0);
        P_RX_HIGHZ_1    : in     vl_logic;
        P_CIM_CLK_ALIGNER_RX1: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_ALIGNER_TX1: in     vl_logic_vector(7 downto 0);
        P_CIM_DYN_DLY_SEL_RX1: in     vl_logic;
        P_CIM_DYN_DLY_SEL_TX1: in     vl_logic;
        P_CIM_START_ALIGN_RX1: in     vl_logic;
        P_CIM_START_ALIGN_TX1: in     vl_logic;
        P_LANE_PD_2     : in     vl_logic;
        P_LANE_RST_2    : in     vl_logic;
        P_RX_LANE_PD_2  : in     vl_logic;
        P_RX_PMA_RST_2  : in     vl_logic;
        P_RX_SIGDET_STATUS_2: out    vl_logic;
        P_RX_SATA_COMINIT_2: out    vl_logic;
        P_RX_SATA_COMWAKE_2: out    vl_logic;
        P_RX_LS_DATA_2  : out    vl_logic;
        P_RX_READY_2    : out    vl_logic;
        P_TEST_STATUS_2 : out    vl_logic_vector(19 downto 0);
        P_TX_DEEMP_2    : in     vl_logic_vector(1 downto 0);
        P_TX_LS_DATA_2  : in     vl_logic;
        P_TX_BEACON_EN_2: in     vl_logic;
        P_TX_SWING_2    : in     vl_logic;
        P_TX_RXDET_REQ_2: in     vl_logic;
        P_TX_RATE_2     : in     vl_logic_vector(2 downto 0);
        P_TX_BUSWIDTH_2 : in     vl_logic_vector(2 downto 0);
        P_TX_MARGIN_2   : in     vl_logic_vector(2 downto 0);
        P_TX_RXDET_STATUS_2: out    vl_logic;
        P_TX_PMA_RST_2  : in     vl_logic;
        P_TX_LANE_PD_2  : in     vl_logic;
        P_RX_RATE_2     : in     vl_logic_vector(2 downto 0);
        P_RX_BUSWIDTH_2 : in     vl_logic_vector(2 downto 0);
        P_RX_HIGHZ_2    : in     vl_logic;
        P_CIM_CLK_ALIGNER_RX2: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_ALIGNER_TX2: in     vl_logic_vector(7 downto 0);
        P_CIM_DYN_DLY_SEL_RX2: in     vl_logic;
        P_CIM_DYN_DLY_SEL_TX2: in     vl_logic;
        P_CIM_START_ALIGN_RX2: in     vl_logic;
        P_CIM_START_ALIGN_TX2: in     vl_logic;
        P_LANE_PD_3     : in     vl_logic;
        P_LANE_RST_3    : in     vl_logic;
        P_RX_LANE_PD_3  : in     vl_logic;
        P_RX_PMA_RST_3  : in     vl_logic;
        P_RX_SIGDET_STATUS_3: out    vl_logic;
        P_RX_SATA_COMINIT_3: out    vl_logic;
        P_RX_SATA_COMWAKE_3: out    vl_logic;
        P_RX_LS_DATA_3  : out    vl_logic;
        P_RX_READY_3    : out    vl_logic;
        P_TEST_STATUS_3 : out    vl_logic_vector(19 downto 0);
        P_TX_DEEMP_3    : in     vl_logic_vector(1 downto 0);
        P_TX_LS_DATA_3  : in     vl_logic;
        P_TX_BEACON_EN_3: in     vl_logic;
        P_TX_SWING_3    : in     vl_logic;
        P_TX_RXDET_REQ_3: in     vl_logic;
        P_TX_RATE_3     : in     vl_logic_vector(2 downto 0);
        P_TX_BUSWIDTH_3 : in     vl_logic_vector(2 downto 0);
        P_TX_MARGIN_3   : in     vl_logic_vector(2 downto 0);
        P_TX_RXDET_STATUS_3: out    vl_logic;
        P_TX_PMA_RST_3  : in     vl_logic;
        P_TX_LANE_PD_3  : in     vl_logic;
        P_RX_RATE_3     : in     vl_logic_vector(2 downto 0);
        P_RX_BUSWIDTH_3 : in     vl_logic_vector(2 downto 0);
        P_RX_HIGHZ_3    : in     vl_logic;
        P_CIM_CLK_ALIGNER_RX3: in     vl_logic_vector(7 downto 0);
        P_CIM_CLK_ALIGNER_TX3: in     vl_logic_vector(7 downto 0);
        P_CIM_DYN_DLY_SEL_RX3: in     vl_logic;
        P_CIM_DYN_DLY_SEL_TX3: in     vl_logic;
        P_CIM_START_ALIGN_RX3: in     vl_logic;
        P_CIM_START_ALIGN_TX3: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CTC_CONTI_SKP_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CA_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CA_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CA_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CA_RX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CA_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CA_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CA_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CA_TX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH0_CA_DYN_DLY_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CA_DYN_DLY_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CA_DYN_DLY_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CA_DYN_DLY_EN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CA_DYN_DLY_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CA_DYN_DLY_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CA_DYN_DLY_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CA_DYN_DLY_EN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CA_DYN_DLY_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CA_DYN_DLY_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CA_DYN_DLY_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CA_DYN_DLY_SEL_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CA_DYN_DLY_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CA_DYN_DLY_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CA_DYN_DLY_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CA_DYN_DLY_SEL_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CA_RSTN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CA_RSTN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CA_RSTN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CA_RSTN_RX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH0_CA_RSTN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CA_RSTN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CA_RSTN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CA_RSTN_TX : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_CTC_CONTI_SKP_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH1_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH1_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_CTC_CONTI_SKP_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH2_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH2_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_WORD_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_DENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_BONDING : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BYPASS_BRIDGE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_RX_POLARITY_INV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ALIGN_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SAMP_16B : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_MASK : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CEB_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_A_REG : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_GE_AUTO_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG0 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SKIP_REG3 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_DEC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_FIFOFLAG_CTC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_DET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ERRDETECT_SILENCE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PMA_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_MCB_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CB_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_AFTER_CTC_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_RCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BRIDGE_RCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CB_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_AFTER_CTC_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_AFTER_CTC_RCLK_EN_GB : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_BRIDGE_RCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_RX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCIE_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_PCS_CB_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_BRIDGE_UINT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_GEAR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_ENC : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BYPASS_BIT_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_GEAR_SPLIT : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_DRIVE_REG_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BIT_SLIP_CYCLES : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_TX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PMA_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PCS_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BRIDGE_TCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_TCLK_POLINV : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PCS_TX_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_SLAVE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BRIDGE_CLK_EN_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_DATA_WIDTH_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_TCLK2FABRIC_SEL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_OUTZZ : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ENC_DUAL : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_BITSLIP_DATA_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_COMMA_REG1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RAPID_IMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RAPID_VMIN_1 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RAPID_VMIN_2 : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_RX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_RX_ERRCNT_CLR : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_PRBS_MODE : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_TX_INSERT_ER : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ENABLE_PRBS_GEN : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_ERR_CNT : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_DEFAULT_RADDR : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_MASTER_CHECK_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_DELAY_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_SEACH_OFFSET : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_CEB_RAPIDLS_MMAX : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_AFULL : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_AEMPTY : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_CTC_CONTI_SKP_SET : constant is 2;
    attribute mti_svvh_generic_type of PCS_CH3_FAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_NEAR_LOOP : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_MASK_7 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_0 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_1 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_2 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_3 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_4 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_5 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_6 : constant is 1;
    attribute mti_svvh_generic_type of PCS_CH3_INT_RX_CLR_7 : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_CLKPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DATAPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DATAPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DCC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DCC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_CDR_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_CDR_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RXPCLK_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RXPCLK_SLIP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PCLKSWITCH_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PCLKSWITCH_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PCLKSWITCH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PCLKSWITCH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_HIGHZ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_HIGHZ_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_EQ_C_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_EQ_R_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_BUSWIDTH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_RES_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_RES_TRIM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_EQ_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PREAMP_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PIBUF_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DCC_IC_RX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DCC_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_TRX : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_SIGDET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_PREAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_SLICER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_PIBUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_PI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_DCC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ICTRL_PREDRV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_TX2RX_PLPBK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DATA_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_UDP_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PRBS_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PRBS_CHK_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_BIST_CHK_PAT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_LOAD_ERR_CNT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CHK_COUNTER_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_PROP_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_PROP_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_SAT_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_SAT_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_PROP_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_PROP_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_LOCK_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_LOCK_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_RX_PI_FORCE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_RX_PI_FORCE_D : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_LOCK_TIMER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_TURBO_MODE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_LOCK_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_LOCK_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_INT_SAT_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_STATUS_RESET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_PI_CTRL_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_PI_CTRL_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_STICKY_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_STICKY_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SIGDET_STATUS_DIS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_STATUS_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_SAT_DET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_TURBO_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_STATUS_RADDR_INIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_CDR_STATUS_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PMA_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_OOB_COMWAKE_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_OOB_COMWAKE_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_OOB_COMINIT_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_OOB_COMINIT_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_PIBUF_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_COMWAKE_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_COMINIT_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SYNC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SYNC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SATA_COMINIT_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SATA_COMINIT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SATA_COMWAKE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SATA_COMWAKE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SLIP_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SLIP_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SLIP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_STATUS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_FSM_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_GRM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_PULSE_EXT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_CH2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_CH2_CHK_WINDOW : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_NOSIG_COUNT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_OOB_DET_COUNT_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SLIP_FIFO_INV_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_SLIP_FIFO_INV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_4OOB_DET_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_SIGDET_IC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_OOB_DETECTOR_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_OOB_DETECTOR_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_TERM_CM_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_CLKPATH_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BEACON_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RXDET_REQ_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RXDET_REQ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BEACON_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BEACON_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RES_CAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BIAS_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BIAS_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RXDET_TIMER_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PD_POST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PD_POST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DCC_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DCC_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BUSWIDTH_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PCLK_SW_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PCLK_SW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_EI_PCLK_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DRV01_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DRV01_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DRV01_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DRV00_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DRV00_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DRV00_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_AMP0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_AMP1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_AMP2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_AMP3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_AMP4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_MARGIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_MARGIN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DEEMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DEEMP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_SWING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_SWING_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RXDET_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_BEACON_OSC_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PREDRV_DAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PREDRV_CM_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_TX2RX_SLPBACK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RXDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_RXDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PRBS_GEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PRBS_GEN_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_UDP_DATA : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_FIFO_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_FIFO_WP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_DATA_MUX_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_SATA_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PULLUP_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PULLUP_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PULLUP_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_PULLUP_DAC3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_OOB_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_SLPBK_AMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_ACJTAG_VHYSTSE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_TX_FBCLK_FAR_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RX_TERM_MODE_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_PLPBK_TXPCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CFG_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CFG_PMA_POR_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CFG_RX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CFG_RX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CFG_TX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_CFG_TX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_48_45 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_69 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_77_76 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_171_164 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_175_172 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_190 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_233_232 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_235_234 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_241_240 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_285_283 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_286 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_295 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_298 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_332_325 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_340_333 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_348_341 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_354_349 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_373 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_376 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_452 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_502_499 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_506_505 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_550_549 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH0_REG_RESERVED_556_552 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_CLKPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DATAPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DATAPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DCC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DCC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_CDR_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_CDR_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RXPCLK_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RXPCLK_SLIP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PCLKSWITCH_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PCLKSWITCH_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PCLKSWITCH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PCLKSWITCH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_HIGHZ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_HIGHZ_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_EQ_C_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_EQ_R_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_BUSWIDTH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_RES_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_RES_TRIM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_EQ_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PREAMP_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PIBUF_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DCC_IC_RX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DCC_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_TRX : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_SIGDET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_PREAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_SLICER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_PIBUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_PI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_DCC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ICTRL_PREDRV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_TX2RX_PLPBK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DATA_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_UDP_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PRBS_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PRBS_CHK_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_BIST_CHK_PAT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_LOAD_ERR_CNT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CHK_COUNTER_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_PROP_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_PROP_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_SAT_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_SAT_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_PROP_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_PROP_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_LOCK_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_LOCK_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_RX_PI_FORCE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_RX_PI_FORCE_D : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_LOCK_TIMER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_TURBO_MODE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_LOCK_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_LOCK_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_INT_SAT_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_STATUS_RESET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_PI_CTRL_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_PI_CTRL_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_STICKY_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_STICKY_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SIGDET_STATUS_DIS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_STATUS_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_SAT_DET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_TURBO_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_STATUS_RADDR_INIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_CDR_STATUS_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PMA_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_OOB_COMWAKE_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_OOB_COMWAKE_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_OOB_COMINIT_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_OOB_COMINIT_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_PIBUF_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_COMWAKE_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_COMINIT_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SYNC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SYNC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SATA_COMINIT_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SATA_COMINIT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SATA_COMWAKE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SATA_COMWAKE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SLIP_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SLIP_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SLIP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_STATUS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_FSM_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_GRM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_PULSE_EXT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_CH2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_CH2_CHK_WINDOW : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_NOSIG_COUNT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_OOB_DET_COUNT_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SLIP_FIFO_INV_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_SLIP_FIFO_INV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_4OOB_DET_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_SIGDET_IC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_OOB_DETECTOR_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_OOB_DETECTOR_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_TERM_CM_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_CLKPATH_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BEACON_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RXDET_REQ_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RXDET_REQ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BEACON_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BEACON_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RES_CAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BIAS_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BIAS_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RXDET_TIMER_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PD_POST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PD_POST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DCC_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DCC_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BUSWIDTH_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PCLK_SW_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PCLK_SW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_EI_PCLK_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DRV01_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DRV01_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DRV01_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DRV00_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DRV00_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DRV00_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_AMP0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_AMP1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_AMP2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_AMP3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_AMP4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_MARGIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_MARGIN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DEEMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DEEMP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_SWING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_SWING_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RXDET_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_BEACON_OSC_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PREDRV_DAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PREDRV_CM_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_TX2RX_SLPBACK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RXDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_RXDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PRBS_GEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PRBS_GEN_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_UDP_DATA : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_FIFO_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_FIFO_WP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_DATA_MUX_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_SATA_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PULLUP_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PULLUP_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PULLUP_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_PULLUP_DAC3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_OOB_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_SLPBK_AMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_ACJTAG_VHYSTSE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_TX_FBCLK_FAR_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RX_TERM_MODE_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_PLPBK_TXPCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CFG_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CFG_PMA_POR_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CFG_RX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CFG_RX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CFG_TX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_CFG_TX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_48_45 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_69 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_77_76 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_171_164 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_175_172 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_190 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_233_232 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_235_234 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_241_240 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_285_283 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_286 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_295 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_298 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_332_325 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_340_333 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_348_341 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_354_349 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_373 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_376 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_452 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_502_499 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_506_505 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_550_549 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH1_REG_RESERVED_556_552 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_CLKPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DATAPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DATAPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DCC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DCC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_CDR_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_CDR_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RXPCLK_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RXPCLK_SLIP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PCLKSWITCH_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PCLKSWITCH_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PCLKSWITCH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PCLKSWITCH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_HIGHZ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_HIGHZ_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_EQ_C_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_EQ_R_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_BUSWIDTH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_RES_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_RES_TRIM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_EQ_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PREAMP_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PIBUF_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DCC_IC_RX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DCC_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_TRX : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_SIGDET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_PREAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_SLICER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_PIBUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_PI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_DCC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ICTRL_PREDRV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_TX2RX_PLPBK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DATA_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_UDP_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PRBS_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PRBS_CHK_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_BIST_CHK_PAT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_LOAD_ERR_CNT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CHK_COUNTER_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_PROP_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_PROP_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_SAT_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_SAT_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_PROP_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_PROP_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_LOCK_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_LOCK_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_RX_PI_FORCE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_RX_PI_FORCE_D : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_LOCK_TIMER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_TURBO_MODE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_LOCK_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_LOCK_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_INT_SAT_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_STATUS_RESET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_PI_CTRL_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_PI_CTRL_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_STICKY_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_STICKY_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SIGDET_STATUS_DIS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_STATUS_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_SAT_DET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_TURBO_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_STATUS_RADDR_INIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_CDR_STATUS_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PMA_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_OOB_COMWAKE_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_OOB_COMWAKE_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_OOB_COMINIT_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_OOB_COMINIT_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_PIBUF_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_COMWAKE_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_COMINIT_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SYNC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SYNC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SATA_COMINIT_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SATA_COMINIT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SATA_COMWAKE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SATA_COMWAKE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SLIP_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SLIP_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SLIP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_STATUS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_FSM_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_GRM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_PULSE_EXT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_CH2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_CH2_CHK_WINDOW : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_NOSIG_COUNT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_OOB_DET_COUNT_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SLIP_FIFO_INV_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_SLIP_FIFO_INV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_4OOB_DET_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_SIGDET_IC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_OOB_DETECTOR_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_OOB_DETECTOR_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_TERM_CM_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_CLKPATH_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BEACON_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RXDET_REQ_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RXDET_REQ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BEACON_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BEACON_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RES_CAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BIAS_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BIAS_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RXDET_TIMER_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PD_POST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PD_POST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DCC_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DCC_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BUSWIDTH_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PCLK_SW_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PCLK_SW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_EI_PCLK_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DRV01_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DRV01_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DRV01_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DRV00_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DRV00_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DRV00_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_AMP0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_AMP1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_AMP2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_AMP3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_AMP4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_MARGIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_MARGIN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DEEMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DEEMP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_SWING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_SWING_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RXDET_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_BEACON_OSC_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PREDRV_DAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PREDRV_CM_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_TX2RX_SLPBACK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RXDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_RXDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PRBS_GEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PRBS_GEN_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_UDP_DATA : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_FIFO_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_FIFO_WP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_DATA_MUX_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_SATA_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PULLUP_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PULLUP_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PULLUP_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_PULLUP_DAC3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_OOB_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_SLPBK_AMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_ACJTAG_VHYSTSE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_TX_FBCLK_FAR_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RX_TERM_MODE_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_PLPBK_TXPCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CFG_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CFG_PMA_POR_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CFG_RX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CFG_RX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CFG_TX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_CFG_TX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_48_45 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_69 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_77_76 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_171_164 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_175_172 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_190 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_233_232 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_235_234 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_241_240 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_285_283 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_286 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_295 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_298 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_332_325 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_340_333 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_348_341 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_354_349 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_373 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_376 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_452 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_502_499 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_506_505 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_550_549 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH2_REG_RESERVED_556_552 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_CLKPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DATAPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DATAPATH_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_PD_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DCC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DCC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_CDR_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_CDR_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RXPCLK_SLIP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RXPCLK_SLIP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PCLKSWITCH_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PCLKSWITCH_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PCLKSWITCH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PCLKSWITCH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_HIGHZ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_HIGHZ_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_EQ_C_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_EQ_R_SET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_BUSWIDTH_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_RES_TRIM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_RES_TRIM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_EQ_OFF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PREAMP_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PIBUF_IC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DCC_IC_RX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DCC_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_TRX : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_SIGDET : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_PREAMP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_SLICER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_PIBUF : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_PI : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_DCC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ICTRL_PREDRV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RATE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RATE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_TX2RX_PLPBK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TXCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DATA_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_UDP_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PRBS_CHK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PRBS_CHK_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_BIST_CHK_PAT_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_LOAD_ERR_CNT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CHK_COUNTER_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_PROP_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_PROP_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_TURBO_GAIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_SAT_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_SAT_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_PROP_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_PROP_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_LOCK_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_LOCK_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_RX_PI_FORCE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_RX_PI_FORCE_D : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_LOCK_TIMER : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_TURBO_MODE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_LOCK_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_LOCK_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_INT_SAT_DET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_STATUS_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_STATUS_RESET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_PI_CTRL_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_PI_CTRL_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_STICKY_RST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_STICKY_RST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SIGDET_STATUS_DIS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_TIMER : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_STATUS_VAL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_SAT_DET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_TURBO_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_STATUS_RADDR_INIT : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_CDR_STATUS_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PMA_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_OOB_COMWAKE_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_OOB_COMWAKE_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_OOB_COMINIT_GAP_MIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_OOB_COMINIT_GAP_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_PIBUF_IC_TX : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_COMWAKE_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_COMINIT_STATUS_CLEAR : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SYNC_RST_N_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SYNC_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SATA_COMINIT_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SATA_COMINIT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SATA_COMWAKE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SATA_COMWAKE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DCC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SLIP_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SLIP_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SLIP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_STATUS_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_FSM_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_VTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_GRM : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_PULSE_EXT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_CH2_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_CH2_CHK_WINDOW : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_NOSIG_COUNT_SETTING : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_OOB_DET_COUNT_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SLIP_FIFO_INV_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_SLIP_FIFO_INV : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_4OOB_DET_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_SIGDET_IC_I : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_OOB_DETECTOR_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_OOB_DETECTOR_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_TERM_CM_CTRL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_CLKPATH_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_CLKPATH_PD_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BEACON_TIMER_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RXDET_REQ_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RXDET_REQ : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BEACON_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BEACON_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_EI_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_EI_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RES_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RES_CAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BIAS_CAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BIAS_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RXDET_TIMER_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PD_POST : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PD_POST_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DCC_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DCC_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BUSWIDTH_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BUSWIDTH : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PCLK_SW_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PCLK_SW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_EI_PCLK_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DRV01_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DRV01_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DRV01_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DRV00_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DRV00_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DRV00_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_AMP0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_AMP1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_AMP2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_AMP3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_AMP4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_MARGIN : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_MARGIN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DEEMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DEEMP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_SWING : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_SWING_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RXDET_THRESHOLD : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_BEACON_OSC_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PREDRV_DAC : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PREDRV_CM_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_TX2RX_SLPBACK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PCLK_EDGE_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RXDET_STATUS_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_RXDET_STATUS : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PRBS_GEN_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PRBS_GEN_WIDTH_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PRBS_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_UDP_DATA : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_FIFO_RST_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_FIFO_WP_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_FIFO_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_DATA_MUX_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_ERR_INSERT : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_SATA_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PULLUP_DAC0 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PULLUP_DAC1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PULLUP_DAC2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_PULLUP_DAC3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_OOB_DELAY_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_POLARITY : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_SLPBK_AMP : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_LS_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_JTAG_MODE_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_JTAG_MODE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_ACJTAG_VHYSTSE : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_TX_FBCLK_FAR_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RX_TERM_MODE_CTRL : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_PLPBK_TXPCLK_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CFG_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CFG_PMA_POR_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CFG_RX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CFG_RX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CFG_TX_LANE_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_CFG_TX_PMA_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_48_45 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_69 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_77_76 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_171_164 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_175_172 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_190 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_233_232 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_235_234 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_241_240 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_285_283 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_286 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_295 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_298 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_332_325 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_340_333 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_348_341 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_354_349 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_373 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_376 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_452 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_502_499 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_506_505 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_550_549 : constant is 2;
    attribute mti_svvh_generic_type of PMA_CH3_REG_RESERVED_556_552 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_POWERDOWN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_POWERDOWN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LANE_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LANE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LOCKDET_REPEAT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_I_CODE_PMA : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_DONE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_DONE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_CODE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LDO_VREF_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_VCOREP_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_I_CODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_ONCHIP_SMALL_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_ONCHIP_SMALL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_JTAG_AC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_JTAG_VHYSTSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_UNLOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_NOFBCLK_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_REFCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_FBCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_LOCKCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_UNLOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PD_VCO : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_FBCLK_TEST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_REFCLK_TEST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_TEST_V_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_TEST_SIG_HALF_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_TEST_FSM : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_REFCLK_OUT_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BGR_STARTUP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BGR_STARTUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PD_BGR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_REFCLK_TERM_VCM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_FBDIVA_5_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_FBDIVB : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESET_N_PFDQP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESET_N_PFDQP : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_QPCURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_VC_FORCE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_VCRESET_C_RING : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LPF_R_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LPF_TR_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PD_BIAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_ICTRL_PLL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_QP : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_LANE_SYNC : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_CLKBUFS1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_TXPCLK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_CLKBUFS3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LANE_SYNC_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_LANE_SYNC_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_D2S : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_REFD2S_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_VCRST_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_BIAS_REFBUF_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_CLKBUFS1_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_CLKBUFS2_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_CLKBUFS3_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_CLKBUFS4_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_REFCLK_CML_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_R_CODE_SIGN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_UNLOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_UNLOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_LOCKDET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_CLKBUF_PD_LEFT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_PLL_CLKBUF_PD_RIGHT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_I_CODE_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_I_CODE_OW : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_ITER_VALID_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_RESCAL_WAIT_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_I_CTRL_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL0_REG_I_CTRL_MIN : constant is 2;
    attribute mti_svvh_generic_type of PARM_CFG_HSST_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PARM_PLL0_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PARM_PLL0_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_POWERDOWN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_POWERDOWN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_READY_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_READY : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LANE_SYNC_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LANE_SYNC : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LOCKDET_REPEAT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_I_CODE_PMA : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_DONE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_DONE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_CODE_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LDO_VREF_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_VCOREP_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_I_CODE : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_ONCHIP_SMALL_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_ONCHIP_SMALL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_JTAG_OE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_JTAG_AC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_JTAG_VHYSTSEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_RESET_N_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_RESET_N : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_UNLOCKED_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_NOFBCLK_STICKY_CLEAR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_REFCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_FBCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_LOCKCT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_UNLOCKDET_ITER : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PD_VCO : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_FBCLK_TEST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_REFCLK_TEST_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_TEST_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_TEST_V_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_TEST_SIG_HALF_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_TEST_FSM : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_REFCLK_OUT_PD : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BGR_STARTUP_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BGR_STARTUP : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PD_BGR : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_REFCLK_TERM_VCM_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_FBDIVA_5_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_FBDIVB : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESET_N_PFDQP_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESET_N_PFDQP : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_QPCURRENT : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_VC_FORCE_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_VCRESET_C_RING : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LPF_R_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LPF_TR_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PD_BIAS : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_ICTRL_PLL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_QP : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_LANE_SYNC : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_CLKBUFS1 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_TXPCLK_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_CLKBUFS3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LANE_SYNC_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_LANE_SYNC_EN_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_D2S : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_REFD2S_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_VCRST_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_BIAS_REFBUF_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_CLKBUFS1_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_CLKBUFS2_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_CLKBUFS3_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_CLKBUFS4_C : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_REFCLK_CML_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_REFCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_R_CODE_SIGN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_UNLOCKED_OW : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_UNLOCKED : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_LOCKDET_MODE : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_CLKBUF_PD_LEFT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_PLL_CLKBUF_PD_RIGHT : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_EN : constant is 1;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_I_CODE_VAL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_I_CODE_OW : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_ITER_VALID_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_RESCAL_WAIT_SEL : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_I_CTRL_MAX : constant is 2;
    attribute mti_svvh_generic_type of PMA_PLL1_REG_I_CTRL_MIN : constant is 2;
    attribute mti_svvh_generic_type of PARM_PLL1_POWERUP : constant is 1;
    attribute mti_svvh_generic_type of PARM_PLL1_RSTN : constant is 1;
    attribute mti_svvh_generic_type of PARM_GRSN_DIS : constant is 1;
    attribute mti_svvh_generic_type of PARM_CFG_RSTN : constant is 1;
end GTP_HSST_E1;
