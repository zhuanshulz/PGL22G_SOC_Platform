`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CB+5/Q+u/PvZtBZ14y6QPg1zSAKDFm8Ll2LA1q44kD7u8TEeRdDmaItDmE5mQ15
1F4FARCR8CYytVlBWcwHZvjrkhVH3H0OZ6i8GWWFyZcECeSyC5WRqe28ojIcP5Pc
lbop8B8mOsRsRBGWk1k/mlJ54bXe4gExPj/zXizwZWjsjvfoX7Zm3CP8qL7ZDPXv
s76uNGqfXFKZNS1JH3cI6YPGuSPOwgvDrNqg6+RZy8H93WJxj6hUWrjT+cwT4bPD
94QQrUokOp538gEkwdL6uMbwZvqTrZIiX+epfNZWxKA/Sg4FqXJATGUznwHmNh2l
L4XRaQPdVYB6i7j2M1PGr+K1yHcYszteZEndOKNn5v7b5pQ1QckhaFUKHoJ8Zaol
b2OlM515H3iDSScaQqtu5S9Pq5Bpdh+vTHsf3S85GmX+XWhqwHgexFu6BIzjOAqv
KKPqXVAOWMBbI4MrrOcxxFLWb7cA8ImNfHzTUiiXej6qG+OPAap9spIJrh5N9f/v
mta5Iy8XSJVdWDr1w8K3HTrWDkCbAW7tOICCOf6BN9tY1MOyTK7hdDnetWcBURfV
6LLIi3+i8dQLplXKfGuIUFs8sFJJle7cYd8MBmrpKrpcDX5wPf1l3JQZLqL+dJOH
0VIAICQFU//+8yH5StxeCsYtM3SzXYRxbRrwor3sbunk+052GUYei9aiZWiLObYE
+qF6Uy3KvFWW9wrxrUNpTFPJKwQSvoWmSqdJmaCWXyCrRbPddd/yE4YMKo2T3sG0
6uxmosUGl1tQy/Vvhy5z5NYi2XKLzKqyLh78jHTlJ/dWa9/Hvb/dBz/fNwgEraE6
6FkHW24MdATgjxG6MqezvyL0Mxumo0wAnrsOCPZvcsR5jWDfPdoC+WedYKBWLqQX
EQK84kS8adFBudZU33iQk6/RfToPODTgqxC4PUi5iZmMbcWb6JFrfXWTvfk3mik3
C6fK2DX3hp+drZhKyDTTcXjDbwzaKtOitciltt6i4a9DILPQFGvX7Ro8oJBwEmyd
WADwckqGv+rE4Amok69jgboW+rrPr4Z5UIkgQ5E634ZrOk/jYeRPMpPKMHMhM+No
zE2Skk0Bfg+RHWOrdHz98ra8wOatrsY3ECWTHml94ybs4dy+wgRirTEJOm9u6a9m
YmiiBHpzW+EpKGID0Yw6rMzLuVlYREg6rIwDbxLKz9+LLCQHM+tHKpJzi+DDDuWB
dZnFxv6WFSs4MsLcV4d1YWdp446MU/uYvhQ9RA9UVOrUkgjtY5hiu+11uR5fzNeB
/pxGGtlHlLum+NAkEqd5UtmCfJAqIPDX5rj2YWeanGTlbSUTKX+lqHzWKnFBVsZO
fnsOGstiQ9dRB/xBDSLTcHgxCUVLZa3QdozCDehxieeQU4fbBIAolOhtenXqnKj1
cTQSPJlnT2T18za/k89XzHuuZtJRl1JTa9BIY+iTPvw=
`protect END_PROTECTED
