`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qUSSObz6UjIUNG2H3Xg96e32StyIeY1/pUR97A+DyuKbTznT0OFch/amikir0SRv
jmVvyfZUxWktCWHDzYB4D/lShOfl8Wg4HBojy8c4frGhIS+yLVqFoN0v1MVixrv1
w4HQN8n+1NYwTtnpyv0m41M0xkTh5YT3lbFXqtRte3SZIsUty/sw8KTwRxRRoW/4
jQdaZ9lAiBMYzn1FS4WJdjp3XZM0StSu6JwOO3JTtTa8sgtJqlX2qfjSTycn6o5s
IVF9ZOocyT5amTEpQDg2m7Ygj/uK7eqbPZK4vA3kIjuW35WvXSR94GgmpnDwWTym
mGr9KtypEJ5eAMBPxB3XQCmwL4fJKSCxr1H9vNlKDeuMfH7TJtenkk57S24FYr7E
3eOLddEVv6ViW9ElnhGpi7lzFM3g/JFh9XozgfZRHepCEimsGR157KQn18466Ee+
6ATzJ+KzO8BaeQRvXIWE2ujtCMQTyOHuZlJ8kWdfRJTQD6EcXUIUJdOqNQSJNWk0
rHx++qV69PHUUVg/6GcMuB7Ritdyuwkukx/voA7zky/zNiFGAgCpxjROITZASqhr
VgM9enemrpONb+UXLFgoHwzcG5gUqU+k80hRTqEUDQOF+LW3sAmgD2iOsUkD5xfy
/RH/wZ+ChCdhb173i0lvkzqFiEqF/BUBytwGawy3GiL3mBKAQ/Yf0rIbjvHmY0Eb
sW/ER9E7yEjoE1bJgCisC+guxH+FQT6lw3HdLDoTgQhd9zkQ0lcPgnIAr1WeagKu
FmBt7vbpi26MJuC8vbPgP/M1zWUVYzjM0xoMMTOh7nvHz/WFI2ySOfKelAQ/Cjbt
oz0bG5AgPPJDZIs+zGM/AyHlGd+eKrpX14Lme64N+23av6grcQEjQc186+aS18tJ
7iD6VpiTzx42/YBTYJpu+SFsZNfpckWm/r/6J8hY05Y3GgFQ7iCGCD539kcmWJHY
qVb3Hz+SRhvgucwg2kUbS257JOUlFi+GtYUnAx793rONvBIXN8/jyJk5jZsqBGtk
5Ru/kor9hq38H2gxpWscKLEYJNIJ+0uEWPtL7YoJ8mmRu+B0QFRWXcgvWajp3Btt
cXOxtCnMnrejuWmGgR/aVTqKX4mKE4quEFJrjbrWJQqPo5mq4hxgXykkah/zB3iq
I44cor13gCsa6rOCgCkWDNyM0eiPmXMdCupaUu/VEY26ZBHNNsKQEglfbsQTomZ3
HRO9UAYrvcUwEdsUnpPLAFll+l8jMwyNaNsaeUeiXrVQ6T71tiJNqyydlPNrrCzL
iyCbIfY6XIV8TfdGGuotDI1HmCD2Y+eiAg0yxj4x1g6+Psa+NHGdR2ZGDQwLuZ2k
lt2FS4/nNXZDPJsKHnwz71uf9vda4FT5MIdhmz/GQ1jAKwOuY8hHkQ5Nh8BASSmg
uKaKuaTNuZhm4rsxgYdcIDbHhP20gPG1NoV2RR+cmLcguesZMbfN4q2hXyXUp+bu
azZllC+WeS9IQ8C5yTKGKk9PE3R2kI3VllbqG3l0CGTEl5CBZgJjjGlDwcmkrdXG
EtTYkYZaqm9s66V0RQokXlY5N2O+bHidoET/MJw3c7ltQ8ETj6pVPuhmh+6+esF6
OpM6a+wTdqrV7aCfznRFb7zn8pjd5/kD3RbGnCUinA9cI2QmbfP0mTWHxaYw7bUD
LEeDfjbAnD6mVv86pHHf6k2BMVtmE0347uJZZzBcPA5bTrCR+ki48xen9s2nPJG2
mFZNAhaDvnMcGg7dk6EnQHfZkDBwqtr9b83ZOdzYzgTAwoe4VJv8rPqHyeY+Y50s
W7TziIwNO6eUh5ygYUFLHg314X2ipZFqjCovcE4jn+0iDcmJVkxHezvD59Izrufh
pnq9Eqd6tNHM/8fyPSJEQwaDYAkY4RXU0oESDHYB7jnAEZ2MWI034IPeXVMnEyTm
N/67fVQmpXWhczKiKf5Mo1kiA0HWo22iT5h+CmZY56MShFh3rz4ZbsV3B/RNSXtB
etNiDJIWGQHF6KDnWNcFVId7TKw2ur4hn7llYALSbwhxvunaeaObrO4r72/8Nkh1
NjdZpOtFmeCZc09nyRkDblLKgq2BBEnzxnVtygh7qos5Djg+S4uzj2p8A0qchTUa
Jrg5ELFRc4nXC6FHlBT1HixoN9GKBeJxbufvwvyfgmV033p/D3LXq7ybaoDSWW2j
aUiBTzaB98S91cu+zWPgcBY7lsHPU3BqPEUR+mA63ATSsEpiHqeB2Pabhh8tnlyT
MU8QtS572j45GAACLaBciXi03E/zdiGUtZJH57n8zLW5LQt5qpAOutdgqsUl1Xqp
H+zfKjZbxoaYsnfCZECcY3huEbkF3jvEVDeeYzEHA5pW2Ihj59EXjkNhvHzxKITp
6IZ+gO3NyhyMAVXzyq0bn/N3GRXIuDb+o1UM5e59a/mD5PSyiIXVDqssG+n8cAoL
oQWr5ZH5UnxdtV3vQw82EBf0wGU+iyNpM8i/y2U6yGFePYkKlgSS2+OExd+SfOLU
Vlk5Lw9QeySkyx301r07z3v/58BoFHbH3EajKQ94p0Kpab+zjaP1dCMF3n8RtEg+
dGjCN8s2fWZ50Sce9AekVfraFyCFqBQd3Kh76GbkKOXugu+0bzd6KJk5flF8/TVn
6ekyoWsDoX/YyUQ1uOteH6jUWN5cUI8EnZr+Jf//WjWvQMtmdVQsQgVQ81pL0JJ4
82fugY1PlFjQrf4y4aOUTbpDeQ9bUXfb8TmyphYDuUofj4/qRm13n8cM+UAaiWwo
3R45cxP6tw1aLOXtV3YckwZtRme4S5Lfq7tF8C/Gf/hXXYUeuoOv8IQgTbjYPr8m
Zt1erSDONb5srMmRv/ldcrhEPqweA3XDBy4TEIfq7HFxFRLxxBXKGFI4WRj2E1Xq
s4y+lMJ5G1bg77qiylWFS449Faz9Jf1dq5Jvgi3MP0U6+QqiXjWK3banZpbMwZGE
/jLQtYCMDRHHFsAAP174qnivVRyhZh93TSuvJMSk3RC76ZJEBUFX7WBk6T1//bmy
Ei+ryXVjnEMEnD4ZVq2GQVyTiC6PtO1TfZPhJUKai0C6hMy6Lm5eGdBnfxHSdq+n
tdZ9eoRBy8yA5aaxA68vxz+nZNGICLU5vIJBLMfpdJqLN5bm4s9h3c5jMQgO07XJ
0+QGsj98F3QgbRpvZ9n3DNDMQ67lUhCnjE8Z6M4f9G6V/Df+gjf0oYFkpBobSMDk
0sWhEzDof2V28Qwjm1xab5r+R7rYCyn43ESkQt88WWu2W3XulRck240dHBYpA/5P
Y2Zm0gDk8G47NkY/e+GQK0lQ4dF0ZctZ4R0jUnCcILYkDl7UzteunFCTwWa3wjXT
YeEZ9wmRAnm4yCHk0hZo/eqGvTsmGyusvMfuTQ8CeaY1yE3odaI/v5f/H/VvBMhw
FPdVzced0MFHSyzocdUPUIsHxhwjNp/qdBVHZzr9f/IA61HWiwScD/LmskUlwO/H
qex/lAlnWb70VxnXqcfe7mYcxf5uSFmE9OX785P+6tv0ewHznBU4T3PmErNqXCEb
Iy19Bw7qHa3Sawqh+HppX0V1pR3kNeUZPy9CFH/gPF7j6LI9hJCz5p44WgwlNyWZ
KUmIPB8TlrJDsFXq1iDoDJeSoDRBmpv2ISGtoQJdGtF6AXKIODSkUUNLa2/ul/5b
Iq3kCoSjD7dvsR7Kz5J/VpjPik8ZUnODivVSZ81qcOjQtgqsKIfEgtRZcg+CChDN
4al/5OM8zzCdJiY13y2QClvgdISE2cHvC5XEyyHkIzvyc3uRmlWeyL8uP41dDMw1
j9pGWovOYLGVh7Bf2aPlV7PJS2cMmPCaeOWyRK6n267/+odlMnfUE3i3qUA4cHst
JA2mKVMospIEHl8du9inACMvtzDgPMP2zB0QkhbhxwaZNbuZrBpyKpDwtYdJ2Wpo
PXAGU5a5JupalD0U3B5gUOEDkWZsRFVmBH2IcxiKVF1odmtaJl0TPvv6eaiOaYxo
cBXiOzvrAfF9+iwPbj/rk+zo7uUUpo4htw2+QbgG1VjyxwxSxdHGZBX7kZnuFUyx
aReC5WpAAtGSUJupU+XDAkncRJJX5UODk0lo0hLMBray5jmfpjThzqnGuqBpRmFE
Xk+6LrWJWAmQXG3+37nGAFZr2jnS5ByYS8/Qjb/UFzKskSkD6bHGGzdOn6rPY8ur
pU8wPT5Y0sj/RlroaFXemq8nHcktUEsUjcYuFwoR/hDRJ1ecXQhew5zeSzf6ocdA
7oZFlb4+m1O8S7HoKxWuVuPwMN03HbEJYOL8m6sZZFsnB7DIrI+AhjKEkve9dI0A
j7W1xdcMz8Af5dCwj1BSMweB51Ju/hNhnTx5jVha10UCn0bqUZNdIb+0p+iADXwp
WubTpugsWZ77mEMh2geW0fpDXcwP8TH9qyEdror1mrBZVDztP3F0Tbq/m89OExdX
4y9kKHrkt+z116tUhkP8rOQFBWd1nQ0RYjt5FziChR0ol0LR/4YmnvIDYUpa9Pz0
aaSZrAvpYeU+CPZjjYlJ6mjVGHOpgxDWq5H6IuVlFCL2fJkTXxoviVCHdpBkJFFb
yJ3EAgcpz6/mXDrZ9FuV6vapDMKANsGWFr60Qi1CUN2jP5cuOCO3ftI9hPUgBKhV
uk5gpPZl+NdO7kW+8rpgNKTOjPyuG+VW2SzIyxn3D8A463SWKJ/3Neus9qb/GzGN
kG+qKktNR7kVAHTFWWxc4fg0dXtjewRemyXMLCxyjVnrk/sgKv2IxX1JikGVFnUr
mkQdE0Br1jatw5cddxGXm4yBCmUhEugeGlLXZ/4RuJ3X9HZTbZqhH1qSMxHffxqG
rhDzpUnkjcp4AsOubjQrUsXdVsNDvAf+JYHm9F2+gimGBC49NtunpoQRjxEdZdyq
gG2rCtr4Xp8zC9UDOAHMNHClP04X/bAttCVqwDTS5WspnQFsKmEwGt9uX/eTQcEI
aN86qm5fCktM8kn4j+rJFqTf6D7dvRyO54pN9pl9gs9mJr9JDYa2uMoyKuubn7NO
Xmcz8md55yvif4kwn5FC6nyvMLQSbfq7lv6ZjBJPWO4Mt2bxfmAGaYz65hiQqy1h
xMUtAjCmNbTsW9aR6sJSMmFqFmMsyv4+bJ+fQZuYads2P8GCFDKGEL6w3KSvoVfP
kJhAIqvlW7tryds6yUSAnG/q4SfZki9xqofemk1sppIcbUnHbYKPK6F3yojMHSbl
IsqCQ0nFkmletrfUW5QlmCmv04W00L5O05SQBiSkmomzhBhQKd0pyPQ+k3ADKxih
X4LatnatYFVdrM1nObVhmWz5ZU6+qOos1aFE0Xt9vjEQz0KtGYdC5KF68kQQ2Ot4
lT5tv52TkjEMcrdtdrQyqzvVcw3Uq2RWBGVWB8uwYNCp7wuwATzv9uT8lL+qlode
L8u6rWWkTABBMRCeYKR+V+AWH5suGi5ZYdZkaY8h+0jblqhTsbRP0sbjIW5uM6/c
t02H8+DosnIfGtahGKKShOd9BTnCs9jgaUl/sRqKV7A=
`protect END_PROTECTED
