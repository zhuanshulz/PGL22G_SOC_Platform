`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sKZELWwKKk7WY0HFAJI2C+tpYcBnjUmXLa1TZoyDODrHAtSxe24G1xisNxKVCEf8
phHDl8M+qlxWD0241J4VEqWJ4uLJ35Q0ZsyIodZHyGUlsCz9Zy+V1zjYE3e73Cq3
a8PilL2I9ey6khyy1pso96Mq8XB939a0KGpygk7TuM8JFsHczFi552cYQgUdVLx2
tPax/9LGyPR+1XJHGjb7BH+K2W6PCDTN5Km9I2GxFC4KEGcEnVNfK34ZvxjvOdlt
D6BypGhLdkSghPMtmZ/I2HCDPsgq01Op7KiR6uto9Z5ZiHyWdBnIB2xJTSA5J4lP
qmPRIDJqpiorvcLHLkIIkAvzsWYSwDYwwh+AkvL+WGqiXHpe1fOAKtvT7Zw0+RQj
J3X6bIImoTQ6FRk4SuDKPnQ5cQIExJmnhtVpb/uK+gk0i7vLSElNzwna85CslwOY
W0I20FBnjBaytmKxmf8vRfl6Q4BZlzAWUsCU6egXJ2Xy9TGc633E4MDRMNADQTpH
VSfBmFG8vE1P4YO/fVntxyw3Hw7zU1KJNVR5F/J6v/oE07iA+VAAaa0TgxSyicNi
Kgfs5uMzDVAdlc0GhVMqeBz5s1GSMByf2a2r8zvdSpt3yO3RjlHLyOLATQ4g5dv1
najHjkrDomYJxSutmunRAa161ucZoIfg3CyPYrnb4h55WOM6wWWYqvQS2s2WpzBp
u7SwQlEEVD93DkjRE4oh7enrGRepAJG7QCHFyuDKTZX6+wkzu/rF/3JkPXUJsLER
0DrX7FOkQFSwbT6wb6HQFRaaG4bMaeXbxAl2HcEBIW7Q35lh5dWAU0L6cTf+r2pj
qC/9hr/zcLjWNm5JDy5+AO8pmOFi/d3v4dp+C+v/vGDxGDH8EXAYVu/tu4eUUdpQ
U9S58FKPc8hSI9MyYgSkbY1e9+p62TPH/Ss28equWaB/W+fhEmoEEg/q/tNGkWB0
+o/MCHZkfLqzKQu5OCX/E3DgvxlE05nBe26mHOIxivamXK2E08HgDSUhUrl/G4B7
TnEmE4xGZYOjNZ3AbJDfh+QhsEByzi5ImIbcSAUEp5YWrf0+X+jPKx4qojZVDsHh
Mhwp3wjRCmGJWxMye6AdjLwx15z/BSJ7EnYeET372wGzkKexRaWaSC7IgOWLwH+c
hDBcAA5cNVa8wzdfeV5T3g6ahYEl7Qz8d2+JplZXWhGE/v4GY85zG5mFLr59dnP6
TA25l4RJBRPbEdpDS/H1eMTZM/MyySsAivY/g5D471rh52IW5QmdGdH541eo62M8
YG6NK5rKvHJuui+IDdDwzkaZw2Mmye4P6lKdKrxuIfU=
`protect END_PROTECTED
