`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EolIvRh8jnAekCg3E8mPjXAOO7RXe/rVBvY8Aymgv/ErnBT1ntpMZoO2TM1qpUUJ
jP7wtaEx3gHBeyKVmmj6+TDI33Mug6tH8pM2To3Vo0FemRH4YrIS86l6GO5s4KPd
+u4Th9k1pSLgoNzib8hSOY/3bdAFV/mNCuEzyOP9dnSXwdUvlUgmdBMBSSh+E4Pu
bTLdWFc3f0iE+n/MB0Fv2kIRTryKNRiq1QrIn4qAGVLo7OofjDjDmCtv9yEeHclw
4DAYanhsBqTYJdC7AZv9z7kDGiFaOrElIHZEkfP3PWN5v7Uyfg9xtsGsxB+J+xNO
WbI4+goLY+jIShxwq9bbfrslA16bEV91sbTtKLzZLhRoKw/oMLV+Yg80nhovSso+
nRNMzUCL22ISpUyonMONk3CgaFc+wQyCe4aRaApeGAMxm+gXgfHZQEoLh7dRMY05
8u8GeBMlep4qRG5BRMY0uc8yu59W0DN7zrf7J4fVUqmd1Mk7/6KkYF/bklZ0IENS
y3Ev5pI7+sghge45PJSVqycLZ1Zj/1lMmS6mg6VTFUOblE0YMOpwsd0XutDBlwl8
Z8MfmZPkBR38xx4lF4QLMPXQ5Yo2SrjAdHMWxboxiThQr1FRjdtoxUQSM9flbS7J
/zFp6xQ3C82gUpe3ksWw08F19lXqF2ItEIbiSUWSpfUpCa+FcV9Ke0JlOIQoIsII
aqU4wsaceqjQ5AoHdmRL32y0ueeJExU2Fv33ObWHWo6LuXwe/t3aDSfl0eB4MglF
1oSI7qtCKh9Bq3UExjYexeBZOiFfiyiSS16hWd4xsnHs9qHOg81FvyK9376Jwe5H
Ci+y0k+Oao6UXd+WmCi16XPcwJFCrMZUh6n3TGx8gxURT8+2wk4nmWfwst1CDpjN
2v0dkDAnk/H9ucrzFuk7QhBVot3vviCdtpySG3KFuaEGNBS4WyAr1iv0+hcI16aR
N4XlaQ2sihydaDcmObjv0Dhl2lvQ4l4CtyMiPmCiHlgQ30Io1O7w4Uk9mLpfB1VA
P90qEPCTAfcXrxW6/tYMdTNXIFDkUvDwrzsoDvs/ZSeCJ7XckY5nKeHfSlGdjmD3
7XQiQbWtjB8DvL2jHQ+Olbxu4xU5l9mbi5O6QxN9GQlIPHxr+2qQfUESVsk6bP+X
eREIHHRF9/c91Z93ptkcbckMidVAEcIlwqZg9YYegZMm9wHpm5jmH6IKKFNE0344
YzKYk7XhxxvbTGhqfI3I6BUcq2MZdUrstzELu5QEpjjOOBV4uKlJeon4RzzGA3nm
0R/LV6wCI3Y6irpAnHqrmg==
`protect END_PROTECTED
