`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3gtig2aGU455H+7cBS8xZalZDJCJ6RQKCSuKy0F6J6foDNp1XPQsUQK+6KnN10z/
IjBJkEHOxmsk0cEPSziA10Kp+H2uY9MraxBNfQ0l6YqfrVijQsqhTooc/7CbMHph
oUlc4T95SyovQLXU0sQMEng+5I8R8dZOGlBLXjlN4Cii3stS/lbjE8ETlC66p3NC
6p3oraRzKZ34sNNqtMf30Cm8z55zIu9oF8C6DVV4VTMuYoDTJ0U9v4p4RRyKqkyM
iCuzrh7oF2muFr38hBV8SIA2bXD2mljoMdoTim0yL0NlEwzp1lyPHi98hE2HKcfZ
lVjJmUM3cJqS1mmoWFXDwoiaiRE1exhpl2I0UeunjOTh9aTNWpa8yQ82iNU6VqEw
nzQ7Qmhz1xeBkLX1t989NWOgO7diH+n3JsVFhsEMuz+gkWHxn6aFX0YAiR7alztq
Ihu4zgKhtJ1/vqVrks7zxLf+mqGAUQs7k6rDAaklwgr/FBhu8+fFNkvt+B+Pgpih
+5WO9OxPFYg9heKD1FdYrIwvqRL2eChTkuSWOIcIxAKiLSmZJwGT4Wq3+HnIf1Ss
VtGOSH4ZIy33sOTJSyH7qMrG0KBazWsN2Tl+tFzeclK6d2aBR3uOdD8fQi1JGRza
8PJ7ibS/vBZoMFnkiuXNsoEDbJ3pVC4ipyR8yKiy3Le2mxrOTzxGl+Cj9rjaGsx3
R5UJ7uEsj1gf32/3mAiadziy2GO0KiWwL+T5ihAnqEAEnmysmC22rBltZeHP+ySA
iN/zSGRhjVN43rIFr2YCJbsxVUp+MJFigmmGkgATVN3xAFYIN2kEa8EJv/T8IYu1
RBw5YVBR4E0l5MJbfMUfAX6VCJLAyDhkRDaDj+1AzDtIjAxjs6f23Sg9TTw6pwua
jTR5vScxI3VLxrdQ0swG+nkNmBcGa03MPX+2boXHmLernyE1nkk4B6oz+HpadpBN
SENGhD0wand+V/bquEujKyO87d3f3aRe2HSHHHr+gzsj0yfAnpIauXiklUTDd99B
bbVIjvbYlOBMjskNhzMvs9jv6WsXezeHS6aCfEjNvWEOZzLgefLdivVXrisRUOJp
f0DrJCWzEvF9+a4TEmUg9VySLeb690ILLNfJCGI/VyACmkrbjSIobpVm8O7d5UdB
Z9DjKnIuyCWfRTT4zXPL5wEq4g0JTXAcWNu1VZ8G5WDLV6rnvgEgD8eYrsnLpXyD
jSnzcmTz7ZO47hg9Ll2XVl0MUaQ79fF4pIKEBpnapih4N0z3ilyTPnYTO0y6zIB3
NpluzBB8Kebx8bdcfwLrbCaB/g9pKlnvQnyK2oNjRBLw4GQhYHrQ9Kbs5hc70Xwm
1WKaieeYCuaa/oGQ/8kTYimzTvjTjMOK50m1Ya9QfkkCuJbwpDJ8PXaWFJD/rk/8
ZxgRsTCsWPo8vK4Yhg1ie3cUPKQ6LrY6fcn/bmR9MciFe+jABJe+cDCWMg+1zMxS
TcYBbreWgaXVCQID9P0O0xhBctdbGvBnEKmWIiSJQR+xDpdWnDmTizubFld1dKH5
2AxOn498XmiCE/oEv32ym3OLxxcUenUk8luHA9YzZOAbR8u1p1MNcA1rZSdpGILh
XC2aOqKW2bPc+DlL5ZX1VSNc6bAW1bihgJu9Mt0q29cKaa6gB2dxK3SmTPIFTp8Q
C+MQJJK0KazUKSYEawTBP7fZ9M1Wm7+VnR34IRQ0fwUXlUMOg+k7edGoCM+uPODd
HhvgaB8VNQoeAWYApabmCYcu3xkt322r/B4vJYrtL59/xOJ8yGbrBz96cZpjot7R
9Vc6MZv7NVAl5ws8jnMQzJXEs2n11YVVkuDPxPUkRUu0ZUuhQa8su3wMsuCjQ+Gb
yLbtelWAfGyqzoaA4W2AdZEEBDUqZk6i8E+aQq7mQojw0a5sJA+Q/sDVwALmHAA8
AbOsaXqFLwt1GPENLItxzOKay2ayylUsg7qQ/qacDB3t9TJnnm8ab2tU94m7uAra
vdzzIXe3FLvI4Q+fOaEn21d9Vb9Ns3dUk26u2BROXjgrjrRqYggNdm7dUbelKulL
LGBCmL8gjJ6svEQL/Q21CEsr0r9p6aJkc1skYhTPRlB7gBzzaEjS+EecVETlHX1h
kjVoa32ndHrmDexdXXSm6dfSBe72gEnan3/Hgz1M8IUPtJgdfMlQNZS2PQdSwgFA
wG8uC14Ml/ikhioDIbBgVJejlEsrSCmhtWoacri5mcMpWBk1V9n+5HyaAfUhVxF6
NqVfIEWex4lBS437xHUQnTwbjRZdZPuvwpjqFmVvffe3102F742cTJPlA1T4+r9C
cAiPB9yFga9uUujF/9T1MBWa16HFIJ88doDcDiMxkzERiHZMqxyhqW2072KriQ6k
EuNc6eMLWiwpOZbVBlixQVdllco3aaR/YoP8DsFgfaE4Q0CFmbgrnDuN/D/JZmAk
ih2/9FW6zNDpfTcArcHz3DjVFZ6NDYzDPwNWzue1tZPzjcScjzEFxvFn3fEaVqAi
XHFrotVcWIVlw6HXQyPQBCntAJ1h2V6zACWUO24KEMzp7HEAsNZ8eDMG5ko9bMTc
J9ZCeV5ty5v3nesrb/lkLvv9C2so/z+35z/tEvIw6uOH2x2RmWaVdIwWnvpcxEPR
Pb4tycOl+JDJTT+04mj6SFCM9FWtpgK9+klJNzXlyglfuMfPblBHsj8U4o7Ntmqi
Em+KFbz09QJzTfAaYnT6u/RB549rUJ8UuyrUsi1MUtTwdOYTEd4qCS607C5HvIWU
FNjvuYsrRfwrDdupzfDGaD00EMiMQAM+a8KSyM7tClRfvs3RmLs44+neQCPZrdh2
8SEJ/aZyLMa4fiMctOtXK2plBCClvF1G+/KCrzSAHMhZmM/QIXnP4dFUrDvzF6H8
425smI2CwWWZbugXj4rVhOs3QD63gTNk87j6y0hau19/mWM/jZ8P49wIqibOA1K8
Ipkpw1UWDBskekFqJhqMxEekdz+4wxnxL+kKw5JiY+eFwHgQXdG2tBsLNNU5wVm5
3OK9kI4dbHop9UHdqSZhWM8pnjIeedtbqIbnBj+ofrfFS9JXHxirL/FuSRwe+6ZL
++cBQd42f4oPJeaK+tGrfCgHYnyXLQHMGTHl4HEoak23viz3wiM+Y5flH3FeVDLT
VzeKYPpYOn2o8d46KTG6mGPJ1dUpZX+1HRsaky/s7bUblwCLonvuO7RFvHZD/NfI
x8qVWznTOKvguIVf7yaCKZDU8b3x2w38Hw/gR+bSgXf8Yr/aXyj9wX52l4OSZjM/
wC21M4BNo9BJXa23WJXhr8+LluvUHaqyl7b9zvr+UgqLncowv9AAWHHtDf/f/hCv
AW8S/nLxYwg5Xi61bEaxhi5dtiCgdn+EGaIxRA4QBqiVhJj1sXKu7N45F7R6Fi+/
r8uOBTZw2DdgCPHoU7hzD2SsoDiUKxykd6wknuRak5BQ3LOL4GoeRXxQCiWBs9yY
3qKpi5R1jXWuCUGuj89zRiRHDk7qMBKt92ZKYrVyF9zXn6CzwGq4tq16RcGyEGaN
NP2cf+uuRvDrRtahIA0Mr59i5EHODYFHa8GPXc6xzB8jkOTBs2QcARyCksA86h5b
F1MRgzP/l2VQg7fFV6fgbqg2//s10FCjEGuLHy2IZme41VEGJS6TFWER02NDXAUJ
k1zTi8dgXxYfvWR7h7u6KwoJhlbbBge9WlxKOMknw7g8AQ3z2z9IlpfmePm5Kj/Y
1WNb24g10snE3HlgAU7MN26KvZeTEIn+H7Jlr6Yc8b+PxEvbUDGShqf2EP3fWZS6
1FzLMBgkZq/hW/6T0G94DYesptqVtZafSnPXhpANW/Lez1lyLcMt7iwvIxDXb0L/
kr5++61B0dN+kSpKbE/bC7dBoYPZ7wJwKxu9R9+okn2zwnIvtZbsnSCwY4TTkMP2
13te3g4kFYPXmV9BW7anJaMVtvMHz31dOC7aFSv3ejXU8n5Qq0XsG0ZhpcHKN3Mn
VacbaNB0ujwZZ5Yl1But1255RYb1NU8nQkpM17gJEFLOW5FtAWxbjyRCpg2y/ASW
dV+o6yY434JBD+L+CMYHmKGQLOKdOyTfl7QizJSnLChRQ7kXxdbsYvJdusEsGtJv
38l4WfctyUHFvdtpDxchJve2Z0sF4IlFeCQPwjp27wDXykSIZ9/UnUb5jehLqB0X
RLbny4vaYhlMz3B7f8O4yxE/J4Hsft7m04knn2WBbx9QVV+lcvjz1UySb1ArQruZ
9vMsd0kTJKhEtl0K0YApVcT07N/2QiecejA452PSddkpNjjtddjdBNSapy8vx4sr
Hc5FCLmWuiWHVkdTiYwSQXwQsAzZyRGkfXsSrkXvfqSjvWlTuKPFsxaVf+kjcAjn
u/i1K9qG1b5mSFeDyr8UG3ggaRLSRaR/3FmTSSQEKWYYo2pO/sKPwFGobwABjSTl
AxfbJGLM18VaJjzP0yH18QKCYWoV0vzJapPwvKtd69oX6ZzfFzR2iOAQN/D35OMh
5aq+SC0ghUQ5g48da1oILzZU/Ch0aRlfS3e+Ka/RXNbwl9SrSa7N6rZ3Fy/98gwt
W9uOJTLSeixYm60VAiOqlZmfH85I0nLdi3txsHZp9SWg8/oUcEVcVYWhVhHwQg/B
gup5e8klLl92ARbiqxM1tylhWVhxMOUjkTckncrCYZ/8k36PmN/4Gyxj8FLZ8l53
nfUvzdIlsW7ggbL4pydMIBURbS2twumZ4MlwxrUUdLNme6vFRd0mPtbR5FonDj3c
JdD5w+v1OPIlkkG1Os9m7OIEfucY1T1CCtsdlclnY3/Sq4k0mauW7JWN73RAEAoP
XQDXUm5M4RkJrn2+3nnyBNWCF6T4hF8LKNAaxYuMjy9EW0unXi/135q+957gBgng
qYIjQmDK7NKvoCK2906qGD5ZcVchYHhSpf8v94xK8ap1QvUhu57CoMP2fap0+4eT
kqsPRBkYTp5RID9CQ2vv+wRo5qVeSvz6JScwzqH5jTo/JNFeVVHrwnYvu/dBipM5
ZkdPaAzvD8GEkYo7eTd1UlksLz1w8fOboWnL5GoLWgDPAwp6IPnZpfVsnVMwyJ4t
60iXNzUWeU8ijaFSQxiZQE/Fyl0Ok5AH9YM1cZUGpOrex8H1syYVpFRD9qfaL91c
v8q1CI9YKyqiywx8g8q2JYIrWgHerKy2tsQj3E8VxtC0SQhPHbr/7v5D/hsepFjL
6+Z7TIyadS8e3w90FoJo54p56WBBjcrfThrO3YkRhaVi3D9xMp6MbW+YooHXg10Y
GtI3ZZviX3ci9rdYukNoz1tj5CjNWlOWASi1adGHBLcRXFnxWF8elipe1NL9mM85
UzLRGgmISpOBXl7MFudP09en9Syx0TJLPLoSfaoW7Zey+LcYcfsgK85XAh9I0V+s
s2RE5UnQ86jOldWFLHYXiHO2uAonQhU7Xlc1YQGWwyz67+JXqe0QQ59ABWeXgGaw
aj+fcudZrj1Z7GhGyL/IA/VaK2vXDYidOOq/P4fpeeWlpQSLpnKmeDpSW8XIzRjX
fSQogsvZDv1ZLDY/Yvlyxs/tXVxf+vaZs6IiPQszgbeTHlsN/eU8MuWS6zapatR0
rsCmMEnFTyB+ePqSjOwij7RRpE3q2byJZSq9MBfJPc84lP5zLBeKLQ5DxFjkDs/7
QofjWjGpwWFCMdX3PNRmR3o/Y5xDbWypnvbQDQ/PrMLSZdwmXFYogoLbWKTvVmUc
e9R2INyUe77VCgDg1MFEFvXGB/ME6FB/JcBIgDnlT+s=
`protect END_PROTECTED
