`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HcowWV9eYW7N8qe3MewWSEcY+gLMZhdKD776FayRmTBQRn6NdDPUgFN8bwbRDNHJ
DQke4Y0e5zkMpDQ7oMokMuF9NVmO8oT9/Av6wuAX3jniu4F1UfER9wIt4dmk+NOA
KIJImojRaXC4oRkSJUnnK9mows7IneMQvJhYMiDA+Gg4RqH9tzC16T0t2sn+HOYK
76L43y1WvV9AUjUreYu6FsKtKPf3tPDivPm5ZVRIePMCacVky9CAmQPNhQ4P3A7m
r58Az7FLKGkF0EN4TYmJZUzo9/cU4OPhkuLjBGq+bK8RiMAY/bSUcNr9ZxN3iRGL
3m764GUPSRKp4+b6CrSRVCHIQ+GvmPGUu86AjeNdC1lh6sNpqmOJKS+8W67SaE1t
125y8f874RCixMCcS1VDmn+oz+ud/drxVpTHNZWAgrgILGu8rv3bXa43MvhVHG0n
fhoDuwYdUleKZhYdZHR43n2akuNIVH51WwINZ1GWrrfYqzXx93xHQ2yMKYT0IEk6
L71NXwD4MqLCGwwYkdKnqpZjBpLtSkDz1i7xU9vMPsXCRLtRe9c9e7R+GnHQyvG0
vwYDf6AUvpiiSQZ4LqeOJiPLhzOie4efJ/jBGjcDD8HGM+jzF1ECRF2u6Q4bz5s4
9/etEOmBBJXQx6gLJo/e4D0bDuNtli0grHHZfL1eOkMMHNm2epf/vahKRHS0hXn3
a74nC50hLuHU4RiS8YP227NXgH/RXwxJ11TBqkzwlygMY+jOXy6QRbnRJOQM62gK
1njAHrBE8Rr+I3B+Amgz8utMtDnSGFXYc0SRr9+1k9/5x0/4BM06nR7XwqLx1Rxe
ErNSy59ZiR/ErZU8mjhP2fwEsQ/MdHxP0CamwZ+Io2bWGcFLYjaGtSAOPUeHTUuy
Ce9033f41TesSVuHVefVV9EBeF5utIbTE8fQoAh+f6QekczWGa80cQmMf83bEKSv
VE86p+z7ozfNUTKXg0T3cLJFpc55v3176ps8al8bdRsXsu/4W7WIVWK2QRNmALsX
govEdzwqrIKT33uhzzLBB+SQLFxHg1+gl5jEjGlngE9WZEwbB1sf3EN2Leg+xlhO
5BCDhFhW24qEjbrhTvuQMRSHOYg+VhpZEP8s9PJZ0VjSrUGgxy22D6eKMKy8y4nJ
G0u4Ed6mOcIxcXsEcdDRzl6HYxsxlG911X6vfTjnl3CvmTYeXgqyAUtEaOKHBZ3K
K3Gf6JzDntTw8heMnk+IQ6pDnIvbzstAM8QHtQOB2KJAu0r2II2ZVL+aW+CLwOtx
CYgoz5cRcfX9e8r/8WT7jU/ROU922MH8nuRPvVC4rbjxYpOUtuWxOkRZF4pHaIlh
ev92Y21Pni8fqL8lUzR6So7od6ioLU25Wa96cOMXMSkGqxoIWZxyV6aV1Z3i4SoR
vMT1galcmge8JXxucgxpvoVU3NOwK1lwb4/sc2ZdSS+H7Fmva8XzzAxTfOtkT+nZ
r0H+9j/Y9R6udl5oNnY4OPT79Jzloks4X7G5+iTdty9FVptGiHPrhfSPPZ+WSui1
wH920gIj2YmjwBbtlgO87Hg5nE81eqvwE+5EHj4F2F5yD1VHJ0WL5PJD2Bep7+2E
08c/oNwT81PazUjtMdyPYQ/g2nSyqeG5w5PpaLtsNuuSVMoDmy210H5SAQZ6+L2z
covPkeDJP5U3/eGHPGN0w4fnXQj8PmXzeAPIDeFH6Qxb9/EzrugS/Uc2LzWfCgNj
dx5nlwxEcIvmf8RnGiRrBQ==
`protect END_PROTECTED
