`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8ErxJM56FIfth0nu3gDDN3CXE+N66dPGvsavApRDS6mZqb1OkFJYrzv5ixMnl5G
S4FAHxZr5zABTMpUlOBaq8k2O+itU1J0VvhjTgPugCvZaW6ZlBr7t1jRFy5XY7KU
zv+xvhj/CnKca+NjE9GG+7Rsd5+Q/BZL9vPv5JsKltDXO4RD0Qe0jA9uhAlXo9sI
Cc32VMj+tYmW0DjtIw6CGIYG79ZCQIwDUOwV1qugcRwinRQfdnEVNoIW0lCQw9Ds
5eVgolOvpbOGRfO10Biizl3ysdMotzdLcpD/ePVKKAQtvCbIdxUzJWaeVFvBSYn5
uZVUgeIpibQHGZDSmJ7MxEmh/oTFh5bHmHb+zzZHMhWj+HWueAcuZ9MA33WrX6vF
ilD67ZTovjpXfgCCFwfUbPdk2tBz0J4JIrAvRMz8ub/aV8ei9FQyr81XPYR4vH5J
Yf6GTbchPbYDOE4HRvNTMzbsS+o2dw+Syu96QZwFtPMYZLig8NerrvZwDG0fMEZl
1DbWBz5im4dEhfkQqMs0STjigzAPgu3S2DX1D1WQ5UNAFO/tvPHIrITuP8mJ5lqK
+Su2Ef/Vvb1jWZgw50L3+0tVj8JEwFjsNbh7r+B/tuL0kElbOEnMEQtpymqxBVyW
OCsnlVSHsEueeYkcGePAQ191Bhzr7lFfoedTot5RhP62wqLNwbndsWcpb04RVkTA
dGMQJH5jaFVW73h2CXBFbLZaTTawFqRO/W8jjBi3yJYYOfaIJUqW34203xPeNP7r
30KH+qs+KgLH1wciRn/wk4R2s7l2kI5Vv8Se9THbsY7fvWmoHyP0dbGrIwJ4/Vrd
2yO/7QEf6ywC60h+xi9H504qm6Wynwan+0bBzn2pmOQw/n3UpfJvU5OBytBodB6v
KHKey1y15MClkps+qs6NFGGfTtXWTQNuDCExkvzbz07rSfPRwk0dbN5I1ITsLHQc
72gGLECOHmQb13FK+F419WudFM9wOnHUCbc9T9WyOBKXTriVSHjuBFJqjb6i/P51
M1jPJG7tvNviizlPcb56qvhg1LpPGTp3IycQgMp9Nq9Uel8P7lGMv/zIDySzasfM
+6smDJDFiGZMW6K6W5UeBbMDCpenTgORQprs+kJcQul18g4py01BbKw1ejEKL7A4
c+QQzz+Z20HHVZpxNOYLZ9oKFd/sxJUli9Nu92DagRue+dQLGoub1BZwD3SFTFUC
cXWCFTlUn+IGyo0X/jvxO17MkAjTVq63rZrapHg8o1/qWzGpCJyPEbewTfQt08Mz
wHm2mHKss1ZQTKbRvD3LfFwITvCDgo9Frjjx+p5mp64G5d9m9858dLcoePEiRvLe
FvLp6WKneHIrMLAHkU4AlMxJWrmBTnfB0aFpnM4Muty6Hccay+Dh/kzvIc6tbutb
qKsHmS40iRYb/I5xysAVEZ8R6BXGweqetqkT3vjVcQcP1Ue+IndtF8Dvkbx8RV5u
xOb9PoJJ9BWLN3PHqdXDLweGuNvVYkSDO21oafurpYWRYgB0wMVg9PacoihxbXPQ
gIVfQxHoqPHZFnHYeXmMH2y9bIEw9jZZ7ZJlG0LlEwyqanpmOB41goSHlnCOZJ7t
uxIBfSCRXC/FohiDKS7FcxN6XIusl/tDVpfnyDc4MyJr/siane4PyY07dx+sXp0M
LKYFeBXULQQcmDiL3FgOkMfgU8xz16dljXpMQAFZsmeasmDzpA9ET6W2dwMSvz1I
8otPnOgs0g78EXJLUbW1BBXmkPYJCCHP0VlBJ+szcEpC2gg2+ORsfdpjps/yaiOt
OB1IZhNNG+qdGKLzKc5z5PO0iOPoWVfPG3tqn1P88V2o4zsKDpDEuGB8VorupSA4
4qXGiMiqcQaAkbfrEeAqh9iompGV514RIRcXUJLg6H2PiuFpVqZ31kkys2agK3k5
pK5FKpGFuso7QYQHnOnRKERiOEqC9FbIbmDiHe517ZTTGBMp0zSiu/XrP1o3bAAy
2FuXK3ooplfeFQmtNfPIY2LdQcNhi5s4AwxqA9e2V95i+c3PzRg8Ej6hksm+K2PA
Er/NiUryLOoADx1oMv8WDMTdTx+ezw90QFBgW5M1nwL6NtsWkA0/6tZZY+1ITNuF
FByaH520/hW+6jhIzY4531w1QazO4B9VEdYQMVFyhQrAxPvda8hyCS0OAIaqcNV1
ibzoPBpkQVozGHuCEvdj9EK8DhoBFjFUhQu8Z8U869tPjhJnGaq+cqFbAVziYMAf
n/43cSQSGxuCERBphGgTqgVhB1IBIBE4yes8WkqGN0Vsg6UBrYCSKSa3/qKW2Wbk
kFFwBBrYRksC6bkxMcdUBvWoKzzibWHJYann8LqemW4d+OswgtQbDVQyPlDYEEhU
4zFhgOWiI7fwa60sJU3RpatwUctrW1TRLWsHCSnhki2AR6NYLHw714+dni9EI/Ej
mDmDLn62LI9r9cWC8TMMn/hlWzt/bdg9F1u9rYC15nwpxO8OOJ8tzDox7zPO1hdF
FyH3wz2a8C67az1y9+osSuM98NkEFN5obYr2N+WvHzptsZzqx+p8TO8T4esAxe79
oyYU6DqcGa/EqitnBKH2/qUXfak/7qe7j6CQu9wS+4r8m55eUE6IWdnZSYOGujN0
uJeLLIaHcdHGgYxHPh3fKaamK1lZZN6Asw7BcigCKC8c0eDX4wV4MD+/8Ei2ulBu
h41+gxmLVikJ34UczpHlSMAh95Mmznm5IDlWY21BZm/QPrz845nQIsHVVlwM9ar9
cHN//u9pE1G8yT6S2MVibw==
`protect END_PROTECTED
