`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lhbeoNxQ5kFwA4bPp3d1IZKXWcRGQw33X7p6/MCqtrhv+bXAiYyzVqIfxSwQEm5H
XBiJwBfpmJ5Frd6Qtk99KwXle592em8La79qOClPAbWFRr/xRWqHy5a1yE6I7Iv5
KeAFbauPt28ZxC8aKjFY/ZgDWk6xXFwsaBzXKvnTv1VTgQx8n5NwUqeoB4SaI9f/
q6lsI3L+S0UI1L0ljkF2pTdF3wGvXI5tR77nZrIJBlJQp8m6+nJB1Nena4tGf9FM
HDOsy2zwBtn9MnHYd600uHLH0JhXsaDwa0Ec9LP7EwaPpgdxJ7wkzeDKWa6pl0Wb
MAy6E2BhH7JQzlMPmsl1/miTXlp/Fw3/EeKbjxGO8ntur1js8YR7S1vj2dzaZpnn
HgWDUlmrPakhriizOMxrctYTTS5eiVWad11qAHIh8buw9Wj9XXA1Xve3D1EMszS/
QcNVSVFM6v3NzLXpAgwSgt20Jmz9Wdti4GUYxdQisVMsVqP0aw7ZXlZDRxNDaqyu
R8hDnxhCzXvjJ9fEbjWMl8XPqEmID4pxhspxxULrw77JeNPCCoDQHkmu7n4Jku/n
8/JFlTccPpeobalY0rger9WW0dEWGHxxgfmFwh+rNl3WB3kynOCOzD1kKFTk29ZZ
bqIOFj1tCWRNdNcS92PdScrlECb4Ph/y69kcL5KQh/Y9NEz9jt6PDVPejbLIBPc0
QTM/G3sD4T86kdEuAaZLu1bOURm6Ad7vYQjs+hpkrGogWip8T9fT8uJYLCxkYmJ0
PnXFWfJQDKaYVDl2b6eUkhqD4J71qm98eDiMbbu4H0qz+g4VGFLT7uNhWCCZappp
/bf81PCJ7rzgLit5UXXel0eDUefpYc416fZrj9nIy6JM5qY+RhtI85iJjHXWJZDG
FYryTdNMfb0RcSmVC3BPRzvI7EdmVRvUTLYn511crNpfW0YMwrx3RDGvk8D7B/Ds
uDDIAMa0elW3sZ5p5V7k5c6ce36CoKu1KP+vstGlJI9Y9Rm31XQ6KzOytguO8Re+
Jm92Ruh9ZR5p5awh5YWI8wFvfkPvAgH5z4oYyyy5VQOFWgCf8NOaBj5sVGYtGtaI
8ot1XVbNGtcw8iggsyDWhL7DsGRud2x01jqomznkE1Jjo5nlTwCxYiytVVCj5m32
PQrbDxeC5A7bkpZKIwa6O2/kxI14h+QfyioMnVBZ+Zle2jstQlzq/CuEHiGXbfPc
a1vn2smOpzyJtGEjSS4xpBnJ8VP5xnPDvq2ty9e+RTs0b4qVUfY8dcJ5SY+Xrr0z
s9RBDCqqzDIe73wx716bQ02FeUyNok4lrBCxfSWEKWhsIIPvT8P4KUQ1oBIP0vUJ
7RlbmMIQHqzmZ1M/tlersoGmrCJfD+SPI8kEI58enhCP3uY+T3hcYF1W8Uvk0gRI
8ir3M4rT8keVQ/ZDU9WLp9cW46zR+CfT14EdpthHLLHQxqPsbonBMl78o51DWYHe
u53MP2xCY4yulnSNIhrOdbkRVjj7l003cKOBNb/8pSJF7oWz5wivs9WHu1UZeR8V
hvj+ifooYMBewLUpRvQuAK6CiOEza104X7w3yUe0UUpVzPchIju0NjGao9reigTU
`protect END_PROTECTED
