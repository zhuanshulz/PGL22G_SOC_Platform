`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FrFhfszaJLkDJ7rNiRxfa/TTl5epEiFrBdcuQAUsszFRgLq8+pRi01V4BrNp+UWA
nc1k2NamvUe/ElrPC3hDOmZUBlefqQZBgYtc+LuQixTWFX6RaAODiVADtN5+u+hr
9KC4pjSSYjWhSkSXs98KezDgxyYrHnCYsVWf/F3ZcWKGHeDK4tfCxjjgQ/GUK1Ui
iQlBI1t28RQOgR1N01jaQaYHXIYDZbwWJBDyzaQBlmkcinRN481nonP2VsTXQv0P
hUNbXwULY4sfnR/OlNBD5ER/Qgd1waeJpiH+QLKJraHXhJubCJlTzObs66bW4Zya
Q6PJQDnnmXTioWaKkCmNjvxqtmipq2C9gEktud2ctBnugt0xeDhS7MiEIxfp/aLs
BDdOG13t74/UpNhs1l741Qd4Yl1l2xgaD+FNlEiu28oS8HI8na0e49V8ulmlusGj
`protect END_PROTECTED
