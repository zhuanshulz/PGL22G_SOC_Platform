`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EnVYopa+AI5PYG56veG09EvwhFFQm5aWzSEZm5uXzONcWaCMD9i8FDd+9CKvDQ2
SGCRewQhRdJyDN2i/9LSvDPMOCE+8h7PojSKfPI+4avEsKEXqimBUaQv1mFj1znA
0Ckay0ORnfOfURdd3az3IKwLU5le8HXFqhBUMSNMZ7j9P8jnozxcOwRK/rmiMQcw
eKXp+j2yqtq1hBvJrFRBuDgd+PuI1C6vFtNnPwSgA6CWGFgk5z7UINRJiXF7Cy6y
oAhfzyuVf2qAf9GsbRImZ4irI91xSu+g/myg05l6es3lsrTSxY3kj9iViwQr4o1m
efPNCL3M6nkVLys4M7aWXiRdhR0pDpgcyEakRIbIoR0VhxF4vF4eqSzKUigzrBYb
gHxTh0APXLG7zrHGRwWAHmTCedgzZZ9znZWEvjzMcOrZw9ktmRiRmZFWHbcTgi2W
o+Udu5YFVCeuAapkw3UiJT7Kk6yDpxdBfWdDxZBTFjJNvCuRCH30YU4Vw9pHOzf+
lPgmX9eC3IPn2MAu86qeT49g/mHm8IevTO86EOWkhg0=
`protect END_PROTECTED
