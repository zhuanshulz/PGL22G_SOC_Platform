`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZAVru1FsYiAA2eif4mBhpirvOze5IzG9exHNxLyVDq2GLVmfqLAFZGfrpTluhuLE
o1gBJuyFMrlY+RZWMblSgNPKi7Eg07jO9pJGjrcCrFo46MxxBMyI/fBBC/zwhtn9
eMuLxrgh0cpvLHujl3O3jdNcqOEy0SV0ZTQ/ziCIGfWgUzMLUnvdrbktbhNX1rVn
FFA+w5Ows6coC0xvjUPgTUKFClWfo1iTHNPoubH7AGuP5AXf+WYmHldIH9Z+fUPj
bvmkIyhXxzYVAjmtLngSKnzzwMQq3CJGZDuGLwxoQHP/J4LXUH/ouSDtMkGzsCm7
xNERH9wlJW5zgDmB44/JsUZbELshbLY5bjHD4zaKPjqTY5rz1vc+gj9ctSeA4NQ0
foVbOjd1l7IncT0rAaJxvXsAqcSpXIZ5JWJa08AKOUH23uP57LK7b3wFapPewjAi
/0brGghnmM7zUZjl1BfT4pRIii7+ZcwBpdU1OSdXS3X5uALDWk9eq78wtgOs/9iZ
8KxygLtzMbq4cSZ8HRv80KyT3Ug473McME9j6ZZqWqZ4S4Zm0RwC1bzvi5X6pvHS
c6xFUi+Eesb9M8mNW5rCeniuWg0iRRKcUh/OpiXec6bC7rJqgqXTMXOMtsRl4rir
PsmADjvQtXZsWqoXRgsilrXsWUkdgzfj+IW+ieKtbljDA80wbuuHzidoAZVNiIAX
SI5QDhP9/e927YeS5KVaNNrV7rGk3Kx0rp8zg4sc/GcBPXQksvtGB8ovwVMju6wx
xjeEjABrd+d7/8M23E0B8j0daUUKSz0DRyJzp1MaEKYOUEd5Lz0c3L1gy4z1UAS2
7bfN5zmaYlAvHS07lyWRnO/AiYNgOyIFOGqkS+JNjbqHCvvkaoPzOqdicSC0r8FR
0alcmUpMHwQWS3Hc4bjXhutpwu7lk+3sM7CGqTjplbUyo4nR3J865QI+/mfJ2Dg7
/NKHggBI/go8d9rGeM+nNfdpF9Q142R5tET+35m5Bvi4vfWdHdVE0zQOpXhuCqnV
zmPIBoaGW0N1Bhjx9LKDhhhcNMPqMQgkV1cf2xxLApc1vF93G9cWQsNPqAWhdE21
RBn4QTCWsY22usgJFK3RGZSlBY5Jbb/ixVpzwnFVjpdLZpa+XxuGKFfEYOZpA3/S
E/hFpGOlj1+nJgQHYueGfOLeEuH4EtS3cgPaDHi8M/gXjAbXepOhuhuSAsjQHQ9o
wrdcFiaKf7rdMDUTJC8J/+mJzHAc+xCizkN5Ac2nfZ2jJi25vgTgb2BgLBjZu8A0
LeuLW2hcaR8iEY1e4lBcK7U1OT9GvLzjLtZwXJdxvZiaWy8qcnkZBkpG+9nI43Rr
glVlXdERDBVqzThWxxkoXZMYb9DxCWBHNlsZhIxK95c3pSr67ZKREpt/odJtiLdn
S41kDriiBqwMvQe2G/JBWB5sjn5TlsLoO8Yv5wGNMIaCYUoD9RDoKqUuouRbxQ0a
wYd7/XdKdKwlYPNBrn3GwI9DyK6QLv37CThZCHlfR7xfy5YqvCe9WHWsWnICrmuv
O4khTz5AszmYHDBwE5Gv8OMr5tscg3WZDQ+pfvLzx3JphjvMrZ/fzKeXByRi6qHb
XiJblddvYGii0uKQCKly/u9uaDAXNjZQK9Q8dAmgQta7HfCHWDqUlcvaJb+6wYyF
hTKmIsFhfr3twgmRcEVfERZE8wBN3J/gbG8kO3eZWhVHvEw5rsnn3Lnor6/PKi3L
0ExlxmJw8a98a/gDPUC+kjEdjijglEJX/qJIVgtfu/JO1T7ZmqZsmLSfH0WFkuyB
fieDOXYvhU2GHMOSJXsjf87y24OlYyIDDROQ6mXTuY5apMt7XNKACB8ReLWvF7Fg
upq8iMhhHJKBLP2yv44XtTX+UT2G8qlnhutuIvSTNyQ=
`protect END_PROTECTED
