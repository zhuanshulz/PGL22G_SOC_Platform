`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sgjd0v06xMJkZPVc2/TPylfIaTXqxdkg9xz0Lm7n7NMdQfPrB6F+NCd7u9JhPOvL
lo5EfV0ROI91GPOpVNUuBzC8KG5uEGae2fT2uwL4DNFyZY6P7mWhoDD2tuKJJxKC
1rfC9jYW3sDMJJcb+r7gd8eNS6VrD7IX/qmuA4atq/3E0VyXyojqIsU1zll/xtR7
Ekaxxup84b2YjJoSjiyrAaQyLDXl0qMNgDrfY7nkByuSXUQ/NCJ8+dtqPewsi7Ux
AyC6FecpXDeZQmRwo5ti98o8f2xWEjTjTs9fLpF2Vy4AhBxl2onSfkaH6ojwDNbY
cFyo36OgJuTCifKYuqc8wo6QcHXNyvhJL8rRR7QMqu2uGobklXCP5wB9e9TX6q56
S0hSa/k2lxbafVdetAExDaBVzmMHeA4/30mv+FS4Jtzr+sm5QmfF1GQvM/YbXVBA
nQgLpluDwMtyJ/RETLckMeQGW1ynVq/L6wb9eP2HMjuq3AuXOKWJ7Bv5Z5YWinsv
stsb3hwfrzvsEVKG/r/Xr64/RkmqO0c0JCy5rXDbCJ7hUQkNbgAOD13creV8SpRY
5S+IAuJj5Be+UpBzjmoD2uf4YM27lkI/nleBwpe1y+qwcfw7sOYDbe9oSOlpTq89
9thRe5BjJT+1Px++N5WpttQPrs2hFkxaFD8hapHdcvrZllH37bI6SKHwFkCGh1N+
e28I2vjtogunjuiOogh/85mbG+dXqvcKURK0zt3YaYQ=
`protect END_PROTECTED
