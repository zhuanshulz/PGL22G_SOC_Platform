`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PpYSv96a95AEERgyNECwrdaEOmmnlkVMjPJt+gNkj2D/mGxqjJQ2HHn7FukjfUx1
wJvpfpUggjA+TuZBJH8KWboWl+p49KriQIH1pXSEgpfieIQ3pdp9EaZsnpzg3hCr
Y5F7RwfqRNnHS0Dm6hVLuxnlkguNnj2xpIOV3eqCZqtjFIVPEGTCuJrUNPqPZDdP
LZMx8iFL8KNZk8ztxWYy13/fKnRFyn10Kl9IuAXdOJyibAFqB+6ip1d59dGFDEj+
Y3UKXTKZFuc35qyFo0ag9iXSNRcUUaFuxZCbaDaEmApF0Q1KeslLG/aDEKjfSVCl
JEnx7hXcS3mxKracryAePns4S2KAxVAs4TcNLCBb9W4a0g0upR0N/7r97wNVUKns
kCE94CjGjTq8BKHZ9PiB8+oRdej62m7tq0ejRIv70Xi0WcABxN//IGt0cic36Dms
MVOQjWfubRS2vn46SEyT3g962e54SyZLJSclBFTcwk5sY/Fya7kwtMNdPuZtNlgD
6/izAPtwkVvQmDeuoH1lnjbWzdnQx+qHRb5RlG5V59JEkJPy+i7LcdxNqbSge6lg
Gi0MQGVeb1wHaxe+YCObkfd8M+PRFvDeAi9hksL4DV4=
`protect END_PROTECTED
