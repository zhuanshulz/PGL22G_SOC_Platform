`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZCAgh7PY1WUWAL4Q+p1NNAmZSIKWyvK8QzoCrRNy3Vn5pHbxuDs6pUaj6PwAqgUE
2Wq80LilnBm9xq1gKh8PCruZ73cuQGjmv5MT4YQh2Kd2IhsqvRkZgOV9LzoVQn3R
F/OpPU9HgJHK3+Phn4aGQF8AQMNVsIzhX7E+hcO4rT7UTTlZ7jYOOdRr2izGyAG7
NBRkbE08ZYrOiFYZiAXmJhne3ioGB1XFxvBIMb+iZh8LNb6B8q9ridT9x98viTzM
8JqrbsO3EPNTYzmvubqce7EX0MqfP0OUhCNPvbSNhNRXhzFAKQ6z0tJCTzwXQMbm
8CW1cY9D30AIsYxByqysK9Rxve0gt059dINBo/e+oNhFgSSAqodUnLKXWnhkfr+W
zlOHxqNK3vV8oiEtrHBFXTUiokET9gDm56Kd4c5BdaTl1gm38TEOyUrUiF4J67ev
lvz0dzKNjAO+9cBQMA+lDnIQd6x4LtxJRTi9wO9hKpN1vlGAhMx54tT2+wH42YHC
rbHdXA3LVCfMvRWzaM4zRGwVOMeYpTrNIUZlUKjB0f68kPbVfXqxyry4eeHS3Xc/
jTRwOI0Q9rL36ZFTpMZUHSCZXP/b4mwJM4y5VYHq4A90zH3HeEfjyaGigg8ZxgLu
ZgBAxuoEWZSwdl4HQIjteos9CUkc3ha39ge4CJPfY0zb4CddktJKkLgJNeciaxAu
S7L0nnRk14MYdH/IV8p4ig86yPUV2UDcr7bGUAvGe97IejWmGFhhctblhqJpXRcz
`protect END_PROTECTED
