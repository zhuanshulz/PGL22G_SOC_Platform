`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01OB3rJBO5y08CWLcOhkPxSxy7y68S0fgSKOkkhiTlLOzGN+7x38FK014dYECrVL
/xgc394DT3dvMZ61Fjr+LzMA/6zM/ptdj3NRKJf0lWIQsCEgAvLLaVdL1usPOqrC
4IjQee1++9ycTGHGyWX8SgYbO8g/5vdrpSEIW4pXYKjHxJbejA0JezUjXGNwN3fC
sXAIU7z6WYRxPpAAu/W9E+KMjm917Q6liDCNJtE2dVzAP2sfKxwkW8YgaOX+x9ru
K9UPXvEPatNonfX6nWD3kkI45BSzecBfZ0P6Ba51AcCIGIP3vgv+XVOfOWGLPKp3
39+KlvxSsk35mo3hPYsLmpQv8vhGx7Kf8367D2XwIbayb1CeN2UsaTR1eQC/Ug8U
IZn5hW4vExOPa6zSIA+gpCNJ2P6wTtN5VJprKnjJDJ0xJ1z127Nzuq6Yf+4mIrha
CHHhzgq+FQgWfsHoD8cBnCv86y3WJeiJ5yB+IO+s1DJXnLGHNI5/liPiXohDOaVE
My9lTJRaJZRP7Hb49N+M3w==
`protect END_PROTECTED
