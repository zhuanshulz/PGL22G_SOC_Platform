`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qP9sHkweVelEQ7ToG43jvpgnbNfYwyn4V7f2G/MKABJ4CPPFEafroDwwiMfnBm9V
clhYwricLRm0kvTOv3x4PaLGapYQsWmJFp5cw5O6JkpDCFdtKjEG0PzCIKXQCR5+
PiHiCAHfP3n9wk8gsjvT/qz4eZB95eg3MImsfzMC5WAWJtGmbfMD6NdsvPt5qdAI
K7j47MiTsmt8TKlmlanfdTOHtvwi+COx24bzqCLSjy8aj+1fsWn31Q3xP0rKtG3k
0m07Yy36b18+WY7ieTux+ZV32R9EyI01YV7V7dORCeCkU9r1Nc8OACg3wGnZxxbk
KNZgDQa/nUWmCvbz5WpAIbBHdfZeMYxsMN5X1zsmRxj7zQMWF0hAHEezkRHddmry
x6ad7qgkpqIPwDwUSG6KRk+nShfJe4VBJzHXi37ZOXVmYZ52H8FJJovwR2fR9EjP
CFkY6MsdufadVFP7TstGsixMCnjGnmsl/kybv7wpxZbzGbtt4rppz5Bj2maF8xk0
iQUykYlCtLrOWWrwpl9Ya37CcolqeBaMkclvnZjgddK90triYSl4kCe86VtDsfav
6ntEu6IH5OrunHSYDjJbA86aidf/v3jpa0TYGK8sbr24gTt5yBejxhPmoQEMeAfE
8EYPIVBVwAN9IFtewRhTfDctWyICZjE4xgvjdwO3XZBrqFhFIpJglN/Qf/Pe+90b
tB6GS+MUA9qIhIZZ4K9ZpanIdaLVzzFue4BlDU1WU94RXAMiMy1BmzZYcLsKHvTN
nc2sRwi5LZ3eRoa6GauKfTC2uJMUJ6AoLcA0yzJRAxCS14ZwZfxrU5EfbCCihmR/
jQb0Q6sxvdAvHZOdcTki6HQmDby/72LxfjkWvDYrS8K/SmppqMZ5B9gwURfoe+d5
IXqWhf2Oai9Kn50ee8aXA5lVNHTBfzR8sLCyTmUB9w/cZO9iYEEhxfBvNzMLejYr
fLSGTTpHo1gka1QzumEEdIye+Eoqjo/fPbcZyZP/uGrSl24xhqDKNFUIt4265M/p
gbxny3MDDtQPagl+MRO7zFU5cURM6mJ1RLJuG6Vyq0g=
`protect END_PROTECTED
