`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sbp0BqUQGk4VkikpKI4+b0EU7+KyFIEdc0dRHBU4sScleOKJJawfPre8sp1Acw5y
mu9TnLYF7rocgse2DXFxXxjSvDdRZpFzebWomwwBN1xNcaNFEhh0i8OMzwVVFNw9
eg/37NsFux/p7uUDb0FQQ8yVRHLIRbhqWTOi4AabGtEddnQcEn+OxvehdiY6ShyN
+ktWBu+D+dFhilA9DOdY1Pkjh+fOjvQp2X1/JyuFBJ9ADG3waIYi+1RE1jIayoqr
6ef0nUFfLKohA6EsVyZk5AfSCrCsezl6eOphwyGHewkaVewV1zbY81yrJjlWgyks
5J2P7tgh+wQFab5s5OoEWeQ2eWePiCSqeMRQsNWO3fHi1X+fswhP+4BOpV+1+9HF
/G/SXNkyj3em22AaUMj1rhOLXvJLXJz+DfVG0ejRjezT4kJAfilTNQS/UXOUeUN+
RpwQ1ZVch/h1tt3p2mC4Yn97R7ZWyGLH9OhdX15hYwVMaBu5J24si+e1GRltAU5R
pn0xBAB8n60Cmeo7IxZM5CmrxPjeWJDo0vxyiZ2t0tloNI1ySL4TASYSCxT38VMh
Rzo6qmR+dLhj04EfnMHCRsIpXlxe+VGmGV0Q5jB0YgjoJmd7F+OUjjuDWRxnIj2W
aUe7aojXrG7062QDGcvYR0lreXC859xSFtofeB6bcQQ=
`protect END_PROTECTED
