`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qitrdiKQE71rev8+EonGZe/cuOQOmddsJYxsdB8FJe85cOV6ihtatqclzN9iakqH
UG9vdGlcgl5zJtKZvK/jnAXjdzwvNzDouGxANxzh4TkO75eKkj52Iec0LxP/zlJf
kMh4sSFL2R2e+aOzzutg2ylsR7qOl9WLA9lBxp+mNQQWTEn5kWlAKK+fGJElkaQY
Ys7kgDtLhiz39y5EvNRLZR2dqctk+m+yLOI6O5U76imCai80rCGTuiToWzUVIxA/
0ylCHgOwFcVReufjw0Z/zRG2AlWeN8yamzZPoOWyMMryfljqKP0cmm3h/NCe7PYO
kNh56wP44iNYKeP4Kt1+u4SX3VvT26fJGdO/B+FDdXOAc6MEhSx90OEOTckS8INC
3Dc5WJae3DBzIhEBUAQPs272n64L/046BLGr5P2cDy0IKbtYe0D/jvhGJoAxFxHF
pNdUOCHLrYgf6lsmddVFHkmmgzvsoNk20ODrJPvhAnSRHMfjSe6GR2hOmmja9f2a
MdXEM2IOCze/Z1HygswO+S+zTa+UXRVWvDzfrVO0tD0u+rqsdrw5o/b7F9Km6bHH
4MwFo5Cy5yMMDJHyekepRg==
`protect END_PROTECTED
