`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ta6cebSRzPJl3noGbaODkqhKIMUM34jG9P0Xoq7sCN6RAloOabt/M6U7pNSK+W/S
G5YpRddZY3FK5R2GrSFePhCjBh8kvFyHe5wYTvA3OSoZobRLoq7JHfvO5mtcc6Vl
CJx+EabNR9Tfcf1j6secH6qB4fCxBgkCchLUpF6cSoDmVbG0z9QfJj6JdloDcbda
QI50RbdllSuEsS1pm3WyNNQqgLyoj3IBjpJY/gHA0Ky3vA+Uei+tjxHrNU3E5p0H
k0NJoTl+La8o/OQYTQwjLb4JI4b+Gd7ZChoxv8xMkEgp5D8g3onRzxvULwP7EuON
TMJSKrF5oqhLh0PvtJhQA7rV3C5zVwcMzdEleWIyQHub+D63DbU0doTD9GE9EmRa
karI4iS/L69F/F2THjCmWrvxlT0rHfxRL7VcMIPqgN+reFgw4ypInp9nP3/eG7vq
l+QFo4RFHzTVWSPDEFyww2OgCVLOfNOQvD0+lXFBOe75FIoWOXFgV05m7zMedod2
Skq35dmabKGIoZBJmR6NUhsRyMWT+1TmgKZSWamZ0D78EOWf4s2sXYXfijuxMlaR
t7gww6oJKIKj87rrbenEC2VVJmatlRbeL/72UVONVNY2nDM3eMsCVTJcdIn3Gl9x
ZsaHu+n/CsUFWO9IcOEfzGJMxePrcktBnyCbgvpoRty8KOOLR4FHmgO1FUItGFKL
GxJHBXfBy8v3k/+BAcN+CGWs7xkCUUuDmWX/rsYlA2CYBQcuaZMzSXCzbTevJQcP
EJ9Yn/HDLUEz980NUsaHNNDbojGtjlZKaqrM/votSH52N/40gUYCaUMLFoihp6KI
e3r73rS3qGe56fOPvfk+DNkHC1Lq+PROwlIP3KKSa+gDOtIf4d5lJegSjY2DuBjD
Fede3v2CUVIJzIxchC90hn0SRmjpF6rgCGyrpDEL0/Gif+n+p9Q297oZcj0HyaGW
mdqCm6SwF7efw3rAoSImkZEbud7gJ89W8HRTT1LPph4DTyElS0vZPJm3VkcUEAo9
QTCobM0xX4euaoXzXPMvIDb1s8jU0+diGL/JSgwByNLCWhAWUg1f4y+ETNeRlU2n
18gWg/brlUGhv4IgVDPKz9URKxED1i7mF7mf1B9WNR5+4CLfN7OBOEqqxQJIxDXk
q8BhwTv21QooAz2qwLt7EsVjuy3nSmSwnitORjziQnn0aRJ4k4AuGpjqvbB8A7j2
8LliEIDEMyl+0JWzXut+jtOGgRyLDkPiS7GqE10oHBMuqB9AUjyZEQFxxTGNIme9
N+iVPjUTRJ+RwbE8XOq+dtU3WHt0XniiB67OV7Z7TyZefmFAVnLsCgRX/CClUJqt
/aoVwhfWlRUq2B8W4Io2cgZYyVKwbjddiQAH9BOOnxLS88dIqr5Z91+ICBS/ckP3
U7kNPMdPbB2A7Q9XAZRVxfLFAV/ACV7QXvU5Fxy/IFfJU1qg156WHpv7XZFMuboo
kz+TAIbAhXoJp74C7cbn48qKfDtQ7WAm0wr12P0pacZCgsghkzS3RwVBJL0Q3PG0
EaP+y8GTx2vKFOsrcY6rhc0wBdGNwIvW4nBX1/tktV2DLVQqW1556EBqxajbrdre
FzSw2pts7z8M+KWXu92JumiSNqXds5yQC2b5zPQw5rrD6QSdykyDZA3Y+tI6LfUK
cvnJKTcg7Suae7ekmQjt5voUofAGS6OTbrItqJmeFAQt9tc40bSSwVknl0jv5vCE
QRCB9WOo4es3+bCUFgBYnBf3CpggkPfBgdXf5exAcYmP8xKZ1cabvHFAtTRztEr6
/tR2ccpn5htMSIbNn71JYt8XF2wqGMYBXLf+/rIBxhgwHS1g6lW6MnOEIVyoEXYr
vfBYpKLqYYOd0YAT7wF3/WSbXzf5tdavpi8xlOdSOYIHbINc/6G9h6zYugGOer0R
QU0e9ZoSDez0VVw/r7+YFyBRLnZ6U31twnbq3tz9HQCX3vUXRhsqX+TC/OLTr0YY
4/4a9pondn+utWqL/UZkODbJJffWVCyjXrUTS1tHk8Pm1AN6jZragge9YM7wogeB
Xo8Zs982E7LGn1SNYd9/OkDEYkFB2SpNBRMz73IpL9yXhpIG7xjpXMo3lLgI1N6J
kAOPD6yBTC9HrjaduytnbjiaN4jOutSsMZhdy3jEUuIuuv7/Ni9HlnLt/Inaoz/i
3eXhIEJJ1pAxfOH59ptHaRJ0Ts7Z976VIBXxBUeLQneTIa8hnO/IY4ciiXVyFTKy
8pIxPJVktMFjd293TU852GACs2sefYaCITYELC/cMdV/U4VOibXkw18q23ODIOmM
rbizxLZl4blSf0bnBO9EIn7LYI0O5hER9TvZeGMjNUeE3ukRuWyxbQmsdXkEvXq2
bEYqvnzrbp7NjbcoWzY80OfJR84FTdKhEHI41xQ8bB59rQrkwfAacKi3SpNB+/T+
k2+ge27Whxd7DenpGKbKa1mMO3SXZOmV00U881JD57H+Dz4k9qSFC6nyeNquDxYs
cv7hGnyOJOoLRmO2F8U9/g==
`protect END_PROTECTED
