`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Y2F94/A9GM6u7ZrsQ5ZuHWl9IWDpktzjtmvzpg3+gBMqYCCLKQktxoJ2g0QPDno
6n4h4mC7Qpb5jtyZWO2WlQB/UNVzpLYyEXAq0eBfKiiD38X1VjJer4x52GGCpwkl
Q/Y89Z2ThopNNchtxWQocOYMPLwbzHIYx6WK0br7VJEzKFQqnya+lwi7gMSDDOcL
xXB4x5tVq/rTMEZ/kELXf7dUA5zOKNxdWLw3RKkAMiIjzjA7BKHBLZ/aThhArDJx
G/3K8V5dBts5kRV9Gyp/NObaTbDJUe2O/8riZs789gprycWGO6gwiS+6MbKOM6Ex
S0Ro/z1XHMi8dGyuSkOQcK+7wx64rcawu8ZHCX4slkA2f6X5dzij70p7tGopZ/k7
Qxogjq7E/C1lQl+j8ky+ab8UA5Lcf9RLpGvtU6CX3Z0BYu7KDTFIwll34JC8jCYI
V8QDf/dlwAij5rOmPNTfIUBu+tQWXUP965sA+1fy1BmVe5BLcQS3mOOj2zD9xXuj
6L9bP7D0CS1k75tfziZ8TlnhCKO4PV3pEbkJmCNtY/AFGHTxgFh7SgYNntDzucdi
zfTj0MBWn7bM4JnqeXTZO9LY7yv0VujXyQ0a48Q6g//ajuAlIGKooVCUg2YBVuL3
qiHTTtqH99LbTVWEWErGQ4Tr4WONJzYZCVQZSHSqgD6nfnR1ulqLE93a2TKPGXIN
EzSs072+SwsI3G3bMNjmRdyllmZWa8ZpNCg9oRjFz/rNS2n6C980usbeleNHYNFA
R25LKGzfCD6xGYBwbkA28oJtpcIpndCqdNWLaENa0uCQMNd2oK2Z1S/GfwAcbE3J
AY+M+MjmzPr8tB6OT72J8Jxa7t/Nm4mOhNiwz3TII8tUnyEzuF9VeMdnraswdEjE
70wWegJhJ14XqQSulddufPVS7eDNy1FIUeZY84769FfW8k722ybFlA7SKMaRqEv+
f1j5Q1wtn8YXuEy8G2EMe1p3VuivFFFLvkB1Q2UL0wLNK4W2w84hT5LF6qNpeS9W
e/F0R9Wh0McgbR8L548J/fWd1+pDbAi/me51c3u18teBrfZH1wfsGCiUCUromxdz
9X69tR4Ns1OuRo1FtdbtXCvRRFPF4gJ4+Gg5xphptkX0+fVzJJoo2ST8os0ISq4P
fJ5hq2vRKl0WY8SrE/cTZJisDX2gaKarBJGG8cqvC1fcp33N+FeUCsj1zJOXDiBY
ns2M5HJZfYB5YMmA2kUq3VU/oz0sLW/2Z39ttv5ahpch1UV1rWfUY639vn6QDgzI
3D4Gl+YltVGT/PW5kNV8Pdd5+LETQVGL1s0cDEt2B1qkoYx1DYwvRxVEJCxB40If
wCW+/bQC2TWoEGsRHQA/vydNISni++l5dZUnMNRgSxoKc9gIhUZJ+9GkQxcWX5Iz
ojHDTRg6uAa1EvL3Ef9KfQe8IlnwS1Bbb65AR3pgx3UigNvKIo4c3kBu7Vv9mwKz
Na+y0A35/MVt/X9w6Zh1pM+mcM4XvcoCRTdtGIb1RvlPxu9yTV/0z3emSV2FgYn1
HDGS3ej5p1jE+RRCOUha0Z4oG47Sv6ku/3tvx59Fhxv2A/+pDcLk4vd3SsPKpvXy
/fJed31+no5bzZtaWc7Zfrb9mpk5G1aGMaM2WD3dPY5wYe5dweAw1/ALRQBw+vnw
RT469c6uBTKNQ/FeCI/H9tYaMtKW5AP8Ek0NIl+C9QdkXLUgZjtoWw9qFE9HPasK
dpZKvw81FiG0/rNGz+rozaoze8Qa/NRH6imnUoZvExUw++aRFQq4z7FkU2dKJ+8R
HRzLxxO7n1Rfh35daoJRNQd/dThpslycTO5WD2hw7ZpyfKwC9HWzXRfu+repGH+s
24+XoEC7+O93QzCQ0PhyzynP3Pz79az8kqGGiMXDxkWIx2L4NCEuR4VRO5LT/NHM
bJ3CtpcM9vaUVYoG/lLe0LSCKx/IprmehcP/erWDahoDYdhbnVDPak5x2G4e2AP9
pW+J/ZBtO3qN5f6+rcYgJQKUh4DIXsn0x6ncn4FVDh514AS2GGfqyDM/pkeBj7Ar
H0bzvsXrHxeW58ZFgQ4CKZgCGIv0hHOc4tkExIz4YsjalMNO3CUA3sZc7TCUY8zG
Cypbozd5GRuBuwzteYGdXtYFzuKdEwAn5RHSn+IukQYvCcuFHJ5Arc4gXl/FEck+
vkoPTHJeS9RRBJKfxoOL2zPqIBQ0fXEEKSn5u6YeAzAJhjMffGXPRs70gZFW0p9p
AjzmdzUbMAa5l2hdDzeZHPHzVyJq8JKb2Q2+nszXNDVWgE+l+k+yUuC8cbVqVGOb
cZ16lKS4TdIIjBJgtlvjTWPb0gKR53oCBmISTB3kiHw1BsHi1N+Zi/la+VvqI5YU
qSeE8HfY7dadCyw2Yrm7AovKuR+R0DvkFpnsMhSnve2xNRRWTvP9g4xkLQUrAjsS
Y96J9xOnCWkWyg5aUEnuiTPnx7f9OGSmUM6nnvnV3WA1MrmAX+v6vBP6xf2P2bSS
m1qq0byoN49S54YRePrC7IUM5SrVoOzKd/txUHNnp4ZTcotHJ90boIRuxSQy4TcX
Kv072b/8t6HTitJig9oNGeX1DRqo+GmN7L42aWSlsYX7g6XQloT6sLUsJAYwg+3i
JD/9f75PmUYte5mayVe1lYhgx4VM4XwRjVdGi7sqUHrL4LdydNDcShHzTt/ATvtR
mH9mP5BsR+ZgkA9Q+frBIywo9Vy1GepRtMx8d26EFrf1F3xSCLVgUyiz+qcRvo/m
mrB5Mb6OoVsGTb3kR3dmbg7XbiXuURJJfQ0LFv/OnGDemlQFpT+Sy16Ap9WZdgdp
RBR90B6YW7xS1qPbaVsuAiJy5tvEqvNP8KdlfKjWuiBWEBglm/aV6Xjv/GRKfNgW
qp8cuIWI5eMX1rU9zuDpgkPZonDzr6f6fwoKGoN4nQ8kOW5V+h7ajCJjxVnlm5iX
oj8mtlyJZNfUJaIoiD7WXCw+D9GaiqZhD1RSlu/sHsHI5fLY+6KR2yZmvAUaxwh5
iJd6FgS3uQYZEplgQg4ViKpwNMQjQnhl/nxPUJkYV4EEqEOegLzLMFq+P+LUotBO
nBPYM1SFxP6m6rhtwjPsPg==
`protect END_PROTECTED
