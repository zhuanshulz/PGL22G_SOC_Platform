`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFXwF0z0Nv0Zt0Wj4EdOaWT1AwWKL0XLWpS1qio9pyCuVsyK4yBO9n2JNnJ7yW5L
6CnFtO8wPSPdPLy/AExEQzJ54HSIoMxDKY2olXFLOGGDDuA7U44AxXTaTAUuOMUM
Th83DmHm8vlMbhLFna8r3p32DIKxsdcURrkcDLr/FrxESebG+g9UNpOafGs4erKK
z7szolIDnigc3r7Y9iSvSykmBxSmKZ6SWv+TJSUtARxhzJIJ6MPOc7hWCH1JEt1E
yX9y5WNeQtAkcQLma4IfPXyGmIMQr8jFG0SB37n42jhgmpScFfU6yxeWso4jULBj
PT+JrmQ26HGkbW79I13w2c71i/s445GmBXT6wajuw54Q2IVTJdAxvLFjppLmdScU
jR1lwws+1nklNuHfZCB1AdLY/gLmtj2wWakWpeDHtQJ6cUBnIIfhuiQm74l15dG8
30yLY2TJzmq3nfyjDJzAtY2a6OmkrKavAAjoSTqsTDocXcSeUhCBEh7y6Ru4I1Do
BULYE3C2+5oAypnBdqEvXWdWRErAFF3u3Nlqe7B0cff8O5zGXW1go42qidYnuXFY
nPJyvvGlrzeATYLnISMzvzKQXbO9K7OWe0g2qD16HcWkudra1wnE/BAlEv3tGeQl
TMWR6RO5evfUiuBycpz1dfK2NB4Td8qP3/MrUHOc4NxSDMjwBaJbfD8nufGy7eJk
9vKP0J42+YcYDn0IdPcMNTDlLtz1E/mgibzQb5+TVAh+OzaK/pzQyEi6I1A305mW
q04jr7SxSX7eEJm0HNcy569ZoJgi8QFEJQLVEaKJziAsyZrhummJY2JA/2+5/XFZ
9DmtblBPNLEcwaWibgmsR/Hc7P/FgsGKKzzAA5wSjfoVo5s/vBz3aDnw1NFJS6rM
zQZLDUSwACWE5JqK+UH+SL/TijKUXqVECdu0DX+ZCxzymzDW/zti7Oo24ycPTk13
YrY0oWE7ZkBbdYxp6RzAzU0+n9QDAKoTXh+81JqmQ+Z/vW2dYVxEnih/p1TxdC+K
z+r0JzJORlPpu63Kx1b1KiFtFI1NG78t0atEdebMv9mwD86H9J2k+D75WtFvkcHh
xzmmXeIoEEC54HSZonYO7TFg2fQV6A+A2NI9t3JzDSpVZVON/DiM+9tuk+gDqPPT
iisB6SeNrXFnN68OOO3NaP70YpJxAIr6sf+qmNCO74cFsSPJ4nbNkDjToh4DH/j1
jjBZbSnX8ChBjV/M8JA61dAJ3goj2/stlmw5ihDfaCd4INzyp9KLe6TMmbUJ9PTf
2AemQlsTcWLdcH4DIzgivXFRoUpDG3xJk+l7PvtON9hbw9qy+WUp+kJ6sSvq/3Ut
kd9SFTfw0UhkgVwtf43lB86yBe7kGSjIC9eRXj716DRkmSa+i0ZOauOS6JQs9Y55
aMKjJwBsaMo6m3/PAS8TDyT/vJqCuuBp8SViaMCsdpcFr+I38Hqc3L6bN1ChcFoj
H6gk8/ff93/CreIojbTuiDraUwQDQj/Z64yARWyrxSrSfTnaQUY9XC0gFNNwy8Wk
TRw6iA/Fk+RO6lwPuwd9zo399AJQ6ZFwYyVHSWnMALl+xs3GtglRFz1xCfE0+Mbj
0oYnYQD/zOarPmS5BjVBp/nn3iU9/tKVvAwJR5c6QedSRJxF5efODFlc0I6b9o5F
vOJeoF5M2xW5uAFlvXCu1GurqL8H70Nbh2+RecmH9wzH67R/cVL/2TNex6dKOO+T
JWm+YeUdQzv46pnJpeswfO7H3WTRNNzvmKXsbI0AtmXYnXwF6TTfiSOUbGqhYV+e
llAT+Y8ayXLyKS6Juqe2hwgaNHvLKh1lG0C487hrXBEbS4b1gi3yqA1f+u7PTyhu
CqV8MQnzS8Zjka0OGI32zLBug1IDkoNSOkp9S5/pyT94psjJD3qw07CnCk9u+qzh
Xk50moLqcYfZ0XeTsZRRQNHJsAyu7bK7+lkTrlhUdKCdEcOA1toxg+w/NgrnGxhZ
oSlKyGgomM28vKBq5QphR604o61i+TlkN26ICgzqawMPFiIF8MsZZlKbgj0Uopgj
Kvy3GsgftxCKAnEmTAMvw0He1lUZj9VIUriOW6tDCiLmRZ62/FTP9H0OoasTd2XX
yI6EnD+m5B8mcQyzodI+5zJVxBjfJTm0MH+Q0eMYoURjuHp5fl7SZfa+iltou94T
8v73+ybBK4XzyGVv67aPe32AtywFf7OvIl6QlHwYY0TuGwrk/qLytNM3QnaXf/O6
ICxkajkC21yD5H5f9NLQOq9nskXgw9qDG737VURjenPJqeazx1cdv9To+fB1PyXZ
`protect END_PROTECTED
