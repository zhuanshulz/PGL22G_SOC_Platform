`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNS6QQY7+g1e0O1Cqi2Y/MKNhfY0Z2Anvb3tByiMtF23Dbmi6i+rra6A8CTwr+4N
/zgHQyQjd6w/ebRj8oONM5BBLmSyhC4CKNdir6KB0N7rQcKaG6Eul3YAeosPBjoY
I8cLrOXZ3HWYw+qRzAr8khgkSHTnn6S3bk3Q8hB4hZ07NdgURbV7iOM3xty9VC2C
0Q83Zpe3bFHUh3WgvEAmNX2vcRxMMPYOwyg7tpPdl5exegLGb6RPmJVmHUihUKrH
eZDPzA9tBI1PQI7h3JOEaaRn3pFNwCeNPthX4RiqIxGiMiq/OCNgMCH9wmQzBzTp
TrMhE2qkXGvtfshe/9wHwA==
`protect END_PROTECTED
