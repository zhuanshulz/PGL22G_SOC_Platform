`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vQL0V0nUSYqxgXAYd3sflPFxY628uqUkB8LfGE9FIeSDm9oWyR3Zzi2WKUTHamad
+OtfnN+IiGP14dfjgWIL604kvUwiCa+ib+L1pgOdbuOvpC1PJqR6YgHP8LpJ6rRX
Vjfe3xysI+x+H/Ja5jFfjoeYhXylxPunbbgogmCmQ25z/K3T5lFQo409fNsNLucK
TXuUJpnL3FI0AOXeLLx7PgYePKQOv/KNWvtrkPMwNC88JJra17jaapvhugCpvvKC
WxjQT/oiUi6/PYnQ4KAtRX0WOV5B2EkOEiQNtz1XTu9HMmMaFpcwCXg6fO3+4yQD
fxQYRhabJcT39yf22nFrpR/o1kx6pY8TlssIEvHIOLpQ9yC2v0PNh8AXItKSBsLR
t3LxtKPxuy3FskNlkg4nQF7+pTDoJM0QQIdDuSzmzGWanwn4P/r/irw0t6CtHV3x
DCho00pZYAZs7RJVIuVRVxifXj6H6QraxE9RKaN6/Fbk7xwG0bIvvaNBTy96u2B6
/qG3LS9ghfr7U9BDc/C3BsWaRmvyfVGOgZBYlcAkKKjoBHhxRwjqWfTUD6Cxm2D7
uvktJ0WyFl2+2JgSN4a+Sh9pO8v0//BczpYSH6eUbdgM2UUahvZMQT3BC5kG5nFk
thIiM7weKCR0Y6MjfjtBUWYAcOLhS4VYr5kw30MXsdmxWoCnoka86GqyAA9483eG
qfC9BO/Dlbe3ZmanQoJ2+1mkeq9AGMD1DUJRAHZKqgWJK/8/5cpWe/OvK4o+bSw+
K77Hln6qP1vPrBYeApKCHvnMTW0yir5wbHlM+DMxUHaIERKeE09fp8Sw6Sotc4jY
oaceg9yUc9EmVTUZIrAwuRNwLlF7xa+Zx16W4mkyX7eK7+aKJ0Wneo+LAmKon4Q6
yBJRltdUl+2uv2A6gI1RQsPbq2y68bKpGadsTPCcWAp7AM6pmAoMJPPE0kX3L0Zq
BKsKZdqxsCcORtK/yQJgab3OyinOnkS58RO+jY2pM1/IjpLLq2qGiSMFFDXtNq62
fvwXWyWkYPZjttaz9T8XGTcC0Md0FqoWRvH06UpcVXNzSIFwbG4zHAriD6H1ZAY3
YFNXXRhiPAEkBZ1h1tZS2i2kH0qqWbDnbcPF4bYbdMcD+zAVk32CJ6sO0BTKssd7
tLo2E1UBhF1cdFb13CjXevQjVIOm2nVsB1P0eKSu+vd93Tk243ZOmXKlxrSU0vSD
cnxMWdTjkl/hNu9W8LN4JScbQ4WOf89qGSZO/bPSI0iSQwygd65d4VH0n7Z7W128
pExv0wsJ64hJFO/Gs7Gd5jxZbebGbWibkqNo+yrYH/ZWd9JAV14dxhV1m5gi9xwF
jIFdloNsAGCoyIrLgf8RcURTaaLzlzhSBMqxOEKI1jKUnxbC4p3+AbxKg+DG1soD
YeljbeSGiUaAcUdP70rpqdtd8OvhqGRDDu9zHXgpHqnjNm+ybQRvHoju6qglQ8OI
0J+7vFRyCMQv7TC4hUkdM4eAt9+w+K9q+NmHfw2VNubuBxGGUu8VgZz6thzPZvwq
W3ACgvc20oO8JeSDD3Zdx1G7i90kwP/F0EL7qtpi3R722IO0Aq22RoXaRf/d4pbD
O2iW4eMqJC6wqRjB6Ip22kaaYFPlxxvkA/YqSx828Zoz2+3fkNFjc0avwgAP21rq
+HwmlkQezu0eebRpu7+CEjMaxiRzTuWAEWAjEAQ+6/jBE2HCKEV6MOjvX4TFSZzl
Q6b5GB0lD98u5Jm08XZ6eLNNI6V2S6ekcFmrIhMRtEIry8ORa+q6OpDh7/bbb10K
vahaML7g7iHAW9AtIbexpPUfBlVBHI8UmRnz3ib3cMV89uWVrrjMSmdzAr0MkVmm
Ed51IgEPh6w1V0gZ4GPasFh7pS25u9a7URksLJQTuDxyLAOcEg6L6w1R1WAfgjt5
K72Rajt3DDW5CpL7eaN6n+so026lMhISJC0/VCRhm7WjOtn2LiVfhvhJlKyXK5Dc
Av4XffUMNrikjGlFbOnSkzNOqxWjfoDHIHp5vO5yfIuJwqPwF7CmWro2jrf95EQ2
+dFD1QW0ySGH2s7/Yw1a+IEV5Wwh4QlsIOfDoeUD3tw=
`protect END_PROTECTED
