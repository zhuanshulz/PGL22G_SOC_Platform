`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bBiFd4JO+0/HsUba0ZKSGJ2zSkBTscqQqfS2AheJ1jkpKOs/l5dMJ7sIf91LqMj8
JO54yFRzyUQ5Nc+P8QLtPHUyuWU67voJGuQyrwf8v4OILAibyIbuEiiw/z4+ypYP
EskalW6MqGw1c7eYiKBC6O0Ip0cE5lqsmDmXeP1/N6uXmpE/2yfR61hDFnGyAOyn
ygxnmF8yitenFx7nQRhiJVX/c+cmGFa9F9HzHKIlR46KHgy/j5JlnwftBacPjkBT
ouD8wMEuK1prJC7WUBuLDq+WjMbTcdYgYiSPm3XtyGkLP6QB6FGtnDiMDbb3K82y
cZ3DB0mDQLHnVVVymjwpOCZwDsjSoaEcwn8iUWb1SqvRwKi44lHd1R1CnrUAHlOi
L5+H7hBrITn7VfYvbvdBrMflJwFrK5gBjZZhxjuKoWlmCTEuXA+90cay5QpCFWBB
MeUP2RXbvS7yzmv/eE3Q/MAGN4YH2Y4fPAbNJ8p/FbNMU9aif3KkCtlbCTM0SFM4
pMcZPxheSDvQhWSAaKxWvCFAnssDv9fSc8ezcNbyXTIMqSkZnhtIl3k/HCpOV1+X
2cJ57vzVeDsZLk5/OH+fwEfaG5sokJO/bnm0oVsx/cEKXgyQLjnbF4OyIJy7ZbGg
PDMW6fx1KpJkT4ZwwWJjNgOSdyZMz9Tkdl2Pdg6J3S40BrD/Yp5CjoLZmkR31Vhs
4RsNFeiS8bJ0mHbTU4y2X8XoLbHzZfq13Dd/rdyAhNhRKzMFRTSLuL/WromPw+cU
QhdTt3Wa5C6F1oMjbcNeF30715NJYZuXHnTTRf8iojJOZVZ8o6pAR0eBVDwzTjEP
l6Wv+65gkaE8fwkX/ACLnWWvH22ol1FJteWjR+ajl50FlhSB5QpG6pzbxq27R1Ep
jp1Pj3QZeOXijVLAq56fbxm+U/4GWeWjg1s7e0wGJpS45awkj/uZR3+UM7maQZZe
qI18M7wn3WvhStPlBQ3nd1AkBuzJ/7IcAR8uI13YKJd9vYXrZl4Up7LoCUJdZg5u
7UbrYblbzSD9KjI+kLl3Kod7uS8b/J8DtXdMOLfGinpl1r22Pcunl+a+XrCyqqFl
if9MwUDuoxaInOhB48DeDYvjB+WyKAKBpNIcGonJkLosHhxwREgYbbf5rUpO9gUK
Hug606GC/VvqkQBnQxHGqifLjC/zcUrpUc3k7cJ9RPyEQ9VKdYuyOR2G/9S7Xszg
UE2msydOZlhnLGE2K57tfPIVq4+Ycdygulu0lMirzMtr3PcyUqpPeQMUuFqck+6m
dTvoOwMfJjHFmLouQsCy6M8hOz3DBRs0mQlXjChAmmiKxdThp6lBaaNXNzrEXXDd
ogHghiI/jYr61/QRIpuATFUTIAryluyo/Yd5xDkEahx3Wt0R6ciHiUvXZhqJogx8
sG/yW29VdtE22cXeSbb+7kPwA/YulUSxSc5ZO1AcIOJ5IIJGX4l+wbsM4VlINhST
rvqmm2AJA384buxc7cpb25uKqRiXJsQKqFCY9eers3GdpPT9WVuhCxB3juQXF959
KqA043gLlUQoy+ZAa+3lobzMS4HbWfGANf+DsvqKDQg=
`protect END_PROTECTED
