`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDg5QXGAMPCpXZ47rPu6YGF3ucZ3e30F1Oek6ml8o3nh9HjfMsgP11ZNKRmAldS3
P94aq4kJRJbu+jdCRDAQmaIW2se1ny489snXGd0LjEb0maUMBXYU4CwYTiWMh9hJ
eBomt/l/ilhshwMfWresnJFuKwdrQHjVNdIQLiENT3ni4RZmBEigVqw0yfBlk2d5
VE8/CM/H9RTbGd8Loa3F1JV16h8UFBgUr212zkwU7KPFMAb8RcrtmiDc9ped3Kcy
bga3OZWR/Tu3rqjKOcStKQ5xMlm1+XK5snHScdWa4p+DOZKGaqgPOqc9Qvw6Oxt9
i6M87Y2iS1NnaZ4adh1U0dHjeE2IDSpgWn7ZTwTHTz1LSLMj7zZfxOx2nzA5M0vY
tiWFmSfMZLbouWticCh4wcbKo4WHp7XBQ7eEatDkZQ+v4YySCA7d/rvK+abR5L0c
zlxkvThz2BFJgN3LXJtcdTcS/IRCycFDvxtwFLhsbG26XVAcQAFtib3w+2Rnde53
6OOllaHzjQh0KTiMNSihWaZorNmhRsG8AfgnxuGojFaKyGFavSK6jp//BlElTpLm
jg/FHFYY8QftvVNvb+IF/YvbtKcVmxpm65z5PYxmcPlDRdYEQESCJAROObolmWmb
SWPCAvt5TZd6JgzwIIYarim4rkt7dBJIiboNpuvnKfWviFilFAH5NSTJsn6MCyD8
mgk66XQO5OVpj3owlEJ8Y+MsVwBjOmM/nq/UpPd+B3+GKF4LQ+DHD0FLlYL72wpH
A2/GBT+64s/WZVJDnXOjpXwv+fmvBseLZtgxjHUmXGt8oYRqtFbGhHGYThpV0B+i
LUxQ1QmtIRXNouGVs3Jf4mKzczEOZo084n85lsqaikZVd/IPKPd+jFk8BaejVn7I
RwhMg2Y204Inl8I8QHHecSV83tDHm+RaveFx6gpiuj6xgyaZeMThTkZXgGUhS5gE
Xk561u2t5GkW6lsXAVgU9iVeKX5CxPLgrZgmZVUkHK3GErNF01gsniLny6vJK99H
O7Qqd7gAC5896asPHjlni6n1McUN7EcK0re5fCpEGlgH+vx9UK6+PXISR2eevLxi
kfYGeYyHNX1GWsCy4vIVcYKAUX11NpaTzibEERGnP9FAIlF5ZHKN7GbXlFNUjCZ5
1ERCSVWSW+UdcIgvepmxxdeZqWmbdQ5e/RCLkzK4YSMFPge1abUFcYIAd/zErwHv
bq7se6Gifqfzie7q6TP3zCO37uM1QrTQezmr720fF5YEU7osqcrWZfa00S2hC/Pb
Z7IuVWZLF7FiLqzhaFeie6VQyw3vhngcahYysrOVsgtpiTwn3UIO5pyIXUNjT2LG
0cEttPYzTzetGpRGZ/Yc3WASJortYRBG/GwpGj3kacZ00ADQkebeDITglqraiENv
gELsHQJSlWR3d6b0dEjJ5e8GiKQjuo6YuzSP/AoKUsXPXnlH2ly3t3K1faOv/jBQ
Rmbcoz+VzDsY/T4JD0E4Ee3bvjRfVxR5IykX/b+K3ak=
`protect END_PROTECTED
