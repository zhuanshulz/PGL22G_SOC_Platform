`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DA9TXzo+fYsFgerkv5f8XfZrypL7sClEmm1ROTef8RZm6dx8Nl7QtvJATC+NZAFY
zONAGEqc/e0lCkZfoW4+atUC2Zwp9flnq3SkV3vmTkiZ1e7JWa2NO1/QSP2xt2Lt
ejoRIFIdarGb74qWUZOOuZ3V6ry+7uNQr+I8EaODc3WBRsYMukzZ836LJp8M0krC
ubRvIm7TqFTt1l/jfFicNGn39raT42XdHazagRnQcfiu+6WCbq+K6YGebdViFZRe
5snM8NH1XFOxpUwsuewO0VlBl+FUUGH8e/JszjeCrniCUfXW/UiT4MMSKUHMZZSP
mzRlHc5KeoSW0spxvADhd04yQOxOSJBzLWXKCg93N/4T50TJpkHQ5CeSeR4vEHxj
hZaRk4OuexxnI+fIdy5vJqkwaGFatrE9tROb5OXQniDNVVOH/sU+t8E0xDMxiI3m
XprlZWBtNzYVW1EEodAmKTGosit/GU/XH40OE5QVDMWk8C4nLvoiav9XtgxdiZm3
4jVgOwblWoJwn6cRQPcCtJDuZLim3WnY19yalQJXbmynPTNglTb+42AiIWSNUN13
cdW5Z9+1qZ+i2fBeylLd0/oJ+XeRoMvfeWZ5f89EkvOluMTabnFduh66qmzQFs22
JB8GgVrOVl9HXvM+Ftf+LqpFJOgRag1n4LTycRhJS+pPqYEt2qLhdfOnvhhB8DDa
hZURar8K0SzKlZ3g0ccpBxznlAPzCfMB/YbCsDlHw96z7lsj9F1lMxuXqixtAc02
/df7ZDWjiubxYeDs40KSLL++JurbXn8KRUTYGpvJQw4a5ZCmp6oosHSos31VhYhh
WgTTN8q8XcWl9BKmAho8c0AhukZeoMkwmss/qtc3GiQhVkPAKVevGKW19Tp+CFDz
gz9Rusr6jMt6mnMy2VCH+bJoFSTe3HpWxNTk8XJut1I=
`protect END_PROTECTED
