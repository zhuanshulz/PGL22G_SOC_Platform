`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYsbwIazQJyRHG75i36AjUGctrCOz4fZD+dpiAwamJToG3r7V6yuBMOsV9nxwRsC
E1OZkgLGz2/JLMybZBhT755Sf8Egi9IJC6JdbmbQ1WPCwkmRU3+z1SFgzcunv3W9
XJV8KdbhBBMYjJYXjKYxcTkFIqVHyV+CABgnWxUom2f50pmvMADih0ay/kNwDH8j
liejohfIR/K6ou2IkeTzRJnGmyvIUJ+OlVxmsPURKO+FV+VqvIDAyPa0JiQYM1Pj
Ws0qJo9na+Fy3NelmMJ/hw/Irt1RjCxiO+m7gTi3kttsgwxScIbhlpQYbEJ+Ft56
Km0s7wx/aEknjwdOJtBkflrsOH4kNaDqEJk5gk0wc1AMPWJDehd0V/37uT6+xhHO
sdD5LN4BfhCdYYR5Ppz1k+mOD56TlTM0nM46eZ7TEVMJAIEw7G/MrtkoYikawAhX
bdUczgw2/slxJNu7r+zJMROmd27I51m+3fDlqzI7n5kwu7Mytieiobegnl4wyqM6
+bLEoXVEQmvd0j3QJjsB5hHJetB0q3uH2hcdQOYyOUp7/D0re3JsbgxnaA3O1DEK
rtYJbS/Wxh3Q8IKSmXcwX4qz9FRiUcTh1F1lsx55IBlFarjg4z0QVS2v1/ms7o/y
Ha78BxZ4SbstjYfPStFtRC+MDbqYotUoMG4pdQY0EZlfnv0vRGMs+R4Y4C1RJREj
Vm4bjf7dbhWa9scK90BpvAD0P39t/uy8MEe4y1n4M95LEOnCb8G+lP+bjFJaQN4C
z/aJnaBhrxWER/eWDXjy7r46O3bYPCGNFlLt6IGbS402ElNbv1+Pdc75AIdq1O+A
Y0fUlKRbeCR7f9d3Mc3VfZXCRdgW6amWY1W7Jwe2cWN3ifQccIxmzdvfU2LUANQF
nD/18he7fgRnfIZVZsckM1BjevjyPyqodJcN+Dsix3g/kP0pHK1ltcUIm5SHTC07
jAxrNmz+nRb3gzjj4fvB+DesGy4ktHbg3jFhBgQKRWNZbMBVj5PLyv3/FYbes5Z+
4DtxaUUr4IzLt72K3W6gVh9S05GqYIdKzGeYqhr4OJyuQmprf36emUm8I+f0pXUX
/3xmoqgeL8MHiNcYs7Tv25oDi/0LK0zVmzuA2QfiT+5ZakIpgouUTS89wpMPTY3y
vERQs3DNgISL8l3+ukCBM5dS0p3fMXYFj8mQFNmMtnJGi+dUB/yBI+FybXDI3Az/
3H5KK5cS5tWLLpqyN5u8CkntcuXG6Vr5qoxndLHwCQqjc7pfvO7IW95BUaUomg6A
Mjk3aAsroCoCJRlv8eacEoK3wXzIIPkISdkSqxWxt12lFIwsoyyGEgVX0lTQ4mDD
Nx/4lUi8lCUKmUkIH1/YO9kqBpZSrrwXt/LVTDWKMcAQVPmBOLlHr1tf/TWZqOWG
4eTf4ijfSl7eTW4E4HcSqgrk4gXQjoMIofdQxMERuDepdtwT4Lws1Y3j6h8ePZnm
oI2Eb+zg7ofX/O3WqVLNf9jwSJQaQFyD7FAXmBN4t3EmB884JgfbHmEpjo01WYKC
XqK9psm8FBI4C4veltoaByw+P4e3zpIy3dUPgNEOPIciYN0WrLhy1EeQlw0ZuRK2
PCTh3ydC1A94IA3AtOuzSZP2/TYkQrkROuQpBPT6s6JkP2H6Qd1l6fc+ULxn9NQX
xsq9UvULzx2VJVev1vkGU1Vw9aZcpfigYgJ6UyaGYyYjmjMWI/9G8CuLSt/535mR
od4qqAQuwcdUxSQ5yyPPd3iWAhi883AxwVG3+DkdeJaLAX8fdypvRSaJTVJdgbW6
8tcMW/ENtCeCuhUsfZ7yDaUR88e0icD6ruVu7p+shYFoUNPYQH34iLrcoNg+GPxY
Ovqny+TNmpEjv/W0mnceztg+0TmAYY+3gv9oeKVZCWWB+UlwQ4+55BoXGksk2t9c
WH65sH5QF8kBw+6A8N1g2A8SJj+swuzwkNurur0zxhf2uKWhcENCZO8qj01j6RC1
aPfC9vIQglNWkKf71aNR0xV3hEhYRKNLLmPDa3tOCHWW9YnG2R8oyVLU5Oc6MxFr
KoGP3Xt+lDsiH4AD6YLGJSPU181FrKfjr5R6rCCZDrLaa020mdOQ7I/Hv5fNqql2
8e0TWoUp4riDDqcy5jy1+SUQ9lB+/WRoPiBffha9VaeWj+SiHttFvk9DXGt2MMXA
GejbtyRWl/ev9b7mxDsO81Jls2AgdRE2MFZzHqg9RflaAbjhhGLuAsNtMxbSFny9
D1+Zow48u5HixA8SKNjJnzI/9xU4ZdP3gPZsVBH3+oQ2mR+Ghcr8JgaNsOtGV0Wr
lAwaJ2nposyTyoSWBVehiX//mUAIPuvqJ7kW7zQUFN9DAexorZWVCVYhGKbdxqNv
u3DzIyW+NQ54UjN81vF63QDtST35eZf7BIQl5toj2wGwBK1uWu5Ol5niBO9C0kCY
wQfy+d/inSRtp+yJ2PFjSuvfbeA+VmLUO6tX5krPoawsgItvXKsYjMA8ijm8WBzq
qQpzmxS9Wo7WD0zTumdLu75Rgiz/LMtpl9lE5JKRLGBQpd35dVzmmrj8I/U2FChQ
iP9ExAOwenBT3sqNnF9wXBht8WRLjjc018XygbHsmwAiXJKxNBF5tK1zdgOd1XnI
j1R00mlfjo11WvnoCZcuW+3wTOX4YFACBDIHh5kGG7V8o+mTnvSc/sUIa6IuTDSk
bXxdquW7fCLsc+ziwnnYpv+tzvaDIktFBHYnoPGXhjUH5L/P6fG7CXAifK0LKrgK
OlAhG4MDSKJONCjcW7IMgnfK/cawYG6DZtZ6F23T7n7gfCsocznd6UTP5tAjmZA5
XszTP2pOTmeysf2r74rhKiSgrT52rMTKzVvNi8MpjRiVPdRKGnxRpD+/nDFc9bvE
W0KXjOZxI8u66mHdMOPLnGqo9W1f1vnVCQexn43XUabK8WOZBXjAfzXpQ3toPIO7
GJy9x02ySL9vuoNSF8xD5Ru1oSOHjbXNS4rMkPVwGapZ2XunwsFWQHNl9OWvRojD
2zSBwRRAkmK/9dRnyWiu6Vrs7uqx5zmAU5YJxG1spLJG3MSoHRFFZYYQJKZWXl2N
cn6rxiF3qekMp85nyjWf493uEnohDm3Br/JhxvWsz+e/TlqYv+E4euot71l5hvfa
MSe64ViCvFIoS1+ncxzTo3QB/KppWeLAFG7yv8FeSsgg1prBJ7mhtDlO6Hry8Bvq
UfS+JqFSAbSD29RP1Bm4qvW+QLjg0CNT9X2Tp2OlIqGG4mDzqlZ4mzp0wbyns/Ov
PqvifLUzdDveI7WF25RUa/6tJLHcD/xQ71edPPcke/HrnoN0YDEzwfL21uL1PAt4
kkf0bRI1SzmoaD4dWtmUVlyiJK4X6Lyhe8lAc6EcH/x3eNdxFp39ZQI+sxPatds9
UA4SBk5XjIk8G86uJsRIeEpU0+ao4MQQ8nE6YIp8QiakQBRqVfK+V1YjRj/smHH5
kq+jsUkGOxMk6ETSipa0hiOlClw3vxv3AO/xZ7opyKdO0REY4iO0kR8e1EoY+AmN
qofMIm9dscUmqy2pyGOfzmagmTXc1qLH/AoTwmvUI47mCriBbvybT6lVtDZzx8gQ
uuJjN2PM1ZNd8REGicFV2T6Qpo23qFxJbuDmkR29ovmVH5E/IySOAnLy37ASir5L
qUU2g/DWsMQ6aijHGT5On5mokH0Kv7BYLNNok4SH4ZBuK6txO3DeMpPCtL5HaAsq
4AaY5P5RFek4ZguqUxrecJ5YpfA5TZ5s6yXSFFmD4kpL7QotSxPmccvnXyltBAL2
WogKz/pbrCgZ7XmnTENPhXFaEvVWVp+vh0eqAkBFsZco7cLnseS+++1nTG0GP6Ho
JgN0568e3OF2cexPcLY0mF5Nouo0RCiHNu1jjK6k/UKPADd8ulbQoB8V47KVlJEH
r5rnTO7aMe1YvBPNkJNoeS500Ohx73h534Fup0Mi+2Hh3kNadEITi1hFej75cvtc
jol6f71GYwMZ/DLdNW01IewRC23qFnIPpyyVZ4dL4m5Q/ZppP1In+qvO/LKgTS5o
cs2DH8v/rgU3eg2tp2ye5b2b350kS0ydloC5H57cXkN2lR8uP3CPHU0Xu1g8WYK/
km/Ks3Pz72fOLNHBsOK8BZFiFRPfeBXxz3rCsWzV0d6FHWRSbS7by8k8OZ1nuXzi
SBVf0Ubk1xUo1T+6sU3yvmexqsns9NxxJ5ZIV5iPTVOpiw/X7+wH5DywYcCHorac
DwXczBxJYJ8teN3iKAve3yZmGnly2d6R0M5ZQEHVVnQOomPucHQUrDV9cgWwd1ga
oT/8pAY55r+fZMbbhKmEIPfCOwjcszv5iLfGJdpCWE8+rxMHNbYqdGdtRW4hr5Ex
cb39VtdKcWm+89rppxG/FLezZhvUH5PwFVvw/3pB6sIQuor9mCw31kyx7QTfUwFG
IYj6qgXXp62rGXLRU5+B7P4+HQxUcC3eyHJQ+AmD87+7Prhvg2eYILe9nCGK7tJi
a02j9cf81uDLGsqRficJQMO6ZnFGXy/n6oTR7mpW1Ur9e6qLBAwi+FMLxJu7Ri7h
za2VLYbGwoaLM8fthtcgPVf2jjz3jq8Jessa7ADASNEvAO1BuHN1o5mC+7CHQx05
MJHjDfdAfMYjl1sUGU3FbCNziSmkxRuNgzzg9ykfAkVDzT4Xpqn95coSq3tvJTml
NkTMExmnqJVR2S2UGAPiFvyGnZqWJlEmJeRnSDubVileyvyV00CrRVyAAmLJaGxJ
BZR1BO53RrVFPnDF7eYnvlc10vlJuQf2l4WjVj++D8BxjkUR2gfLv4iCyOlKdtdJ
Oo4tFqoGKVxUJ649aMo0n6tXs4d388xn4FFtzrjHZPKbIuluz5lVRI55KXYMgsIX
x7VnmQoNGpG3pNKvfVxrD/T8ppScKT28Pqw9Tgkciut5pas8d6Ft8pbrzF5vE3zB
mSqD2S51sSkstlpw37ngAEQYSERk3E+29e/qYQGfUcS11hxGNQrZ/gWckHd2Zd3w
wH/1t30GFORSljd8c6xykOqLpWM8wCwcg8XVYcmWbxLJIhxvIYYZpE9Nrs+7XIWh
44ELcXeYaX8MLR+xvtuqob82WgtcB4b164K/JlgGKWHOV4Yho5OSMk8Zf4qTuvQU
jszmcQ65Brxxm0ENcfHY4+OSkcCKOE+11EemfC9GzEbEk2zLKmUH+WN3mtXLbyfH
+AVsjqdgWqoOLNkdIdHgw4uDcVkuxUHqbjk54kKqN0y1TMce30QEnfFu0jsPdfy+
Gpvo27K1GEwEG1oyV3A/zUNWIMGXalQF0Ao92HoJENy4Yl1HIW5laHPqYeiuRCp6
EoSfFXBBouNS5dh1/QklwMqXroqHRZEIbZXGmalCaARIiSj5DjZlZ+8n5piETYd6
28P7AuHFSGi0D4FgCbqLYv2pd2Agd0Ype9qEbO3fwn3dA93WkXVx4deoE5gQK3Q5
S3wwUPpZK/bjnB0aE1QL93EAQBceTwoDZtWVzPm8m41nOWmXPrjnHE9mxpCKRZqU
8ob90b3m6HESQa1pwnku8EQp1GedhDJvlneCj/LL8u+RVIlhtMvPlmgeEtcXCe0e
Mg5JXERRW0g1BeD5gpLD5heXkFdaFZcRy7hA3x6VBGpkieqkUu74N1nn6vAn1mYw
o6wejx/nZcgpefcOlXxFqUtPGnMkmCLYiaufMXmHa4UBpnolpnuD1IQUUTpIzVY7
MYh+dZfngWbf1zJuDiD5Dx/EFY4pp36PdPanRxLEwRkgh3OD2wp02owHxqQkqHsE
sVmBJ0/9DWbPDB46wequWC4VedcgcwZ8kpa0Hn9GUfCCm9rYVFuODNCHxpCRWXu5
kk9OOVel/oLMXwfLqSX/EQ9OgmqRT6rNBoOy2TMUVpZpqggo9t9w2r6CBua+EHVw
wNmImy+DhxeoGVqPYsLOh1CHrZRpL56kICUciaofaTNhg+CFdIY0rEqlT3htGHus
MhFcPrDjPU53klW/U/IN35bTEjCtYFXZpeZpnRUnLzCxcx4ATNyjr6UO2zbEpilg
3a0RAGinTYeeElhqwxAVMTvvw3S8gSaYMpluZkulBzBoJ8MfmqZuCfFxOoAv1k/0
`protect END_PROTECTED
