`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/R8iMFO5A9PqIgbhgHjGUOPjpev2moUxlCxbMoakL5wz2ylZQNYfBFPR6BpxRawV
JqBzQLRJaJQjl9kI3xgEhh9KE62z5ZYYFEsH+bWoB55+fZVYdZXn/5XEhVWQ80h8
JUlrkp+ctZZLR3DTkYN34eAW5CW6ZgEH8CBKCaRZzsiBNkdxzDGPWdLwJYcSNh1r
k1xJIK5ugD2Vzbh4f9JyYK3pnL8KiJsghXqWNkdLx4EyeQtOunWPhSz7Sv6Cotwt
yrP2K8uJ0xdsRsIBA/pukn8J/HWkf4RnU5nivLMW8E9qBwwDzi7E27nDUEc+yXxP
Zk7WVlrHbYWFWwEteSEmFLbmxaSd9MiceNMEUYwunbjsNQe7QGdWs+07kTIOJKv1
Ke1EJIolBQ8z628AxyteJgSmzj4PFNYRuMZqjPTDHp1YzHazYPOHRQsgd78F0uZa
7g1lVwQllhoCnSjGQ5kKXOwCPTvJEbMocLY3ZjmjZH5jLts67Qf0tJvFY8WU3Ib8
+3FCVR55FYo88VGL/5eQUW7FUbcqPMFRjoBZj2NJKxIIT0bkMoTM9HcI/pNR+52B
2SlmoFgOzjZR43lQWSfRes5oxVWmPsTAG16f0vXWBcbuxV+3fY8C4u/AEn312r4h
P3op19V56/ROHjs/8ACVr0k1We/+b9YhmLQ5lRAAtFxOerKm4S54/lS1WvpzTXxS
qSsAAqJCds6iN+s2ea11poqXZahEGFOgCJGmGoVj9dL/o2As6y2FzqsFUUh77xeF
`protect END_PROTECTED
