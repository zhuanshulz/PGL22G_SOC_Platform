`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A5ienlLF/Qm4oLMXyotI828Jz5QuSUDv6pF/ug3jUclKDF1HKOfV8paspcLkDMZf
HzEJTWoKBqHSFxuPhTqXaz+NarQA82ohcTfuuZZiZdGMmFmvt6gWKHHg6RCkEVlH
P/XxtnK1lJ1l3Br0x9980mm0CY3luj+k8HHuY/CvSjA8zsduUA6MQbdUmvJm3Vuk
V1oYdxYK0/FC9xBV08O64sJjVoB0mV/8xZNtV5Whwkow7oRg22JwTz9ji7RJR50n
V9P4hd2WXqljHVKD5c4+fY03Q+Jr2/wHQb4FwTTdwCV5Fv2sEhCGKOxZABze1FeP
Ilg3wnyRSfKQTDrzaDvJTyT2PvWeqy64q6PbdosCj/98tFz+LgInvJ0giKtQSL1b
Ze8giAURL3e+FXbrcwTa8egyl3GVBP3LuwFd8HqieiGOmIb++3QN3SUUw0ssklfI
BlZ2CXiayd8ntxqF9iOuUxfgkizPfkSPdU9SBR3MaK0=
`protect END_PROTECTED
