`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1MT9hxX4wmpwaymR6tqCOlu5chbeUO6SkUPNHlcCziN1G8ArxC3EpFBODlTEj2lp
+0aotcsgw1138rNyprLeLOw5wBliKwFIe0WSw/oe//KfIOm7/YAMl3hBMvN1acgd
YdF2cG332P94qIXw+SJgnd2lKEKBsb4MpMZW1NA2Xox/6KMrSkoKMHR3NS668Xln
hBV0PwH4MBh807GgOWH7AuUUHoNCqZj/BlNRpEHEuWqMIT81Tkj/MrjfYJsd7wmb
aiIBmdhaoZ5wVrUuIqouqqQiX3kOrGK5SPFEI+g046TWburAV/ueRwCqKGD6OWxw
CCY8p9a8+KliZzadsGHG349IKFZcDqUS3Ty6tobaSgr6JcwLJuBylA99N9s2Vr/r
5b7FOx0ThlwHNpW3ePdwoCve9XX4x6opCEkFG5MdQ8EWa9CTD66lHRgxuoSdgG3A
Va8P0CcWIhDwjgvRdGdDNnuXfVZSkjV4AyzPH7o3p/0eQpKG9B4h0bPMCCv150q6
RSedP7QdPRE/Rb3Qqk/D91jVl5Nexm5Zmxze4GYF1ojEOwzaj+rRhN1Tfwb2ZlFg
`protect END_PROTECTED
