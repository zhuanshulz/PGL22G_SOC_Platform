`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGcuKoq97knLZ8tpIkV9LGJo+QXMirJZdH07sijN6NhYa2JlBB1MDt3y75yxu/lb
7HdVXupYnGZCW4Aw9z9nkLR0B8pfveYgKg+tJSnSusei9gPeBfRRTJENkITchlhb
uOec5ihtYa4ZI8xbfneS9I72CR/X/8LDbjonzGi7elCL/pI2FAzgqCuDA4hTxaaO
mUeiJlBP0F4w2aSsXK5iafwKk7RxckCR4erre/6XD1M1dq/tmNaRrB56J+4BC9vn
rCK5a16YVyb6/IW5ECuIDuwMKfThSEssN3iE/a+aLpXZ+8xDk9nVtNzTf2I+GJX3
oJrgXv4RyK2dwQzRJe6THv7NRMQ66crmiFjUBSIs5eQV9KK/wALacOh0x0/DuabO
jQMx5Gugfrx8gEcaQkLT0w==
`protect END_PROTECTED
