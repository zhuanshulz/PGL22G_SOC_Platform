`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqXJaGJUqciXwr2fYX4oJbpmI0oZN+WI5V5qeFHhgt3qy0u+6f4bAxd08+ldH+rd
wUPFsJYqlTScPDdSz/cc5MOhaDeyVRM/krcxxbZKOfP4a0uWD9ZKlWfssWHYefBc
VKZ/3bvSnEUH2VzOe3PTNHfXgofeb4kfwpTaz9Y+N4KSzO7ZY3skI7eGV1+C4NHq
V3OZPi4gexHR3tyWR9dgDDVpp1EbrUQ4yNWWf5yA5WxbetE6y9xFqdS5gXU44QUJ
ToExd0++T0QDFyA/NyC9pOYuMB/2qQ0glvCbmYiGcGxuLpbVMk1MWb9b7DKACtGq
czcVJi3yC8gPVHt0RcAlNxm8eMAmtmjXZucNXqC0EPkErudq59EkfQZM3QUr739e
5j/IwTRCWjbImisnYhy3RZ06F4BWQAk4FSsrQCSBQxJTY6kpKx4dVC79nGiDBDs+
JKi7LDr8OnfdWYXbyqLfEVBmXoM1tEbgQy2XS43s6tj1aKE7NoXq6Rhsc5Z0f+Xn
Pzf1CDbT4pWUJd+mRAbCRxgASqs2lfBg/IEWsh+RcgUa826ZCcinQdrW3n/UlUN2
nL5HRWrsaCmQUKbZ7E6RDwtVcXCK/Q2+HmXaex3X/U4P38TupWSinG7IooraE489
3Ue4tYMnOnNw1axAiKmb9ATkEa8gKg7Ct/A9+oVQMYDExS4GRhPaJM12vSXrWjTy
0WvX2AN5t5JWZ/x0hgyTvA4rnktTVXG13kR4y8SjL+oQ+ovUW04H8Wc0Nu/hN72u
Pq6NK9KS1i9A0qJG9u3ydLAIomwgNs/QniAwHa2aqYF1gguAbUddl31iTtmgc3YW
oaxkWdTAugxOm0RKFGGe5R7OVB2S30J8G9CV6K7yEzYpudtFabuFel0c7xi8KAfa
+IYQJua1oHpX4ycQ44TungtwoIayUx5UA3usDW1eoeDbMxDBr63A/HNLF/qriwNp
Lr0FTPNi4475qDpkfWE3uq7tHxHpDAq2ewvGfrY/oTmvne4EYym8YlGFSmD6yBbh
3ZsOT143SV9fiU+B71QVhH7hboezBU6Je62y/Rh2pAMIG2JUuHEz5RN3bNJWK8AY
U2vAk5/USQbzkISnw46wCSY9yvY4YOb4AZK+kNTROTwWua/IL9j4WovWKobexdEm
CFbPokNYF5lIPHccb02dnlXtLWcDiLb3gYBYhJEVv4HMSD48gbXITolj8AUxJ2FV
hFP2LxOZZKwlKAMOfKl4bPJo2vauEVFrSVhZN2qUFGASn8MoN5Bj0GMp6w1DSYZy
bPVPZLdyaNNfstjieehsQOZZlJWiBbbRECzoMzPR/KlIgHPxkXHLa01r+L+46dfz
1Jp/lmIS85+ARM+mYoB0MTfOC69WWyQMerqE0xwPyJdKVenoTqIe3VW1fstrVSdm
wvoVnE56z3koSmr6rj8IAEgWq7vP7s7sNrYULoOuz5XT+UM3b8y5am8unLIWmAkv
`protect END_PROTECTED
