`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZq3dHwIO/vdVuyVughofL7g/wxR+LG0vJqLsbJmQHEE1R5r7DnqX8vL60c8p9z9
hrf9N7lXsP/WhabmwaMtq2ozxYs5CQx/C8WueWCTgB4OkVUqzHqvIgGYwksCseca
OlHFczALl6U8RhkQ4s+aeGYWziW+T/f/iCCFvcxBe3Lo3CbUDY6RWsWYwv/na7Hu
fbxmK7ontqfqBfn2CUjiaRHYuAr0BrwhY5tuH9tVZjRn5tmq0Cuj494eSQwjdAA9
4PKuIy2y7ifVzoY8kgK4t6dSRIY/TX4jzPaIqGj+52W/s1SD0CG1RSXvLS8DjOaX
swwK4dDlx/UUc43gptHtRjW8+Qjd4bR/MCh+D7MFNknWWO3YSdzC/vgSuRxjvxMQ
b6JrC8SKX3Bi5TH0wnT5Q+c4c/i/yMvrNKrm21qJev0WJbkw1swST4xDo4F6xJdS
9/ZLWXTVN5cfYRfACj4Pgr6FIhzPEgSyiDdCgK1VXlQm3icj5SPlmqnMGH99PBy5
azy3B0EAKG0Ccw2lDWiQyw9plBO1js5/6LjDoAQ1E1UkRuT8lrYmHVUfyZ5HcUtg
qKpauYjrX4wBO2obWD/CRZp2lNzK2wzO4bCm8NS+x2URcnYoUW8wSiMvKmbGdgho
GQotBE9oCls2xDAFoNA/g1PsAmX0hsoj/V+/D8G+w+M8z2WPpqF24841zuHOmLg5
j1kBjnH8Y6mFprF41VSGzSlkJVTNdaXOY0APRf09TmaJkEtzqjYCYOFKW7wlIsGu
ouDa1pZwZSL8fGFM6oKD3Vpecv0/IvKN8VVuXwoa+oPbDEXCb4Ai5RY1H0cwZ3ET
`protect END_PROTECTED
