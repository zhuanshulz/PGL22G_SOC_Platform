`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJJlW/37cqLznYkVRAoXvwm/1JMtztwzD5eJY6MmqpkzlI1QN3mQUXz7S9i7Sw59
/JejFfoKzw1zQC/IJXDrQCU+rBumlBkN2164+6riFUkfCsLaZ5cSV7gpR7NUawn5
XYp55TOZd094dMbnIuBhSeCHEiwIzDNnN6KAKbwV1Q9TR7kS8JFtr+mfluxffN6l
boqxcK7XVqpC2qt+qk9rT5hZpiCw78UsiGlq/GKvpey69V1zXmBg6ljj3hmu6mjs
t808BcFDz71qTlrZCEZZ5B5gfb1IPH9QsoeJ2137LSOYkZ/hETrSlSpD3Ow+KiWD
1jXUYGtVRuLlX3G24AtW53YFhLXSBe9dRPFGZd+MSgyM1Po9Mxsh5CMetRsKjTSg
TgrA5HOqqSwaewpEIRzk5uHlL+XYv7IAWAY/kinWQ6FUZWyP2zmhxuS9rNM9Y309
9DK4JvGRKsMwDJPpZSQI2QIiIh+c7pM+LL7y0HkJ6+x+L+z+0erCX7ATAgECLgQf
Iccen6eDE1jcbilEhKrXUqq50FR5QtuLXo6xUMvbXSvULF1PULQH2xS+wZ2Hr86L
xCgploNAvsYTgFfucYncWt7SOMjlTquloKWBL2oJTdo1rM5pkmRw3/Ded9ptbIC6
cDIBBE6DhtXZklETNjYae/qyJQFTmCc7FIC3vb9Pus8XX+KfRrmbTMN59Zby+u3Q
DRNrI7Ggc01qeDMZn1hzpc54uvfrI1LixdAdRBVx2KULfAYaEUIPHrn1yHaCn9hz
wwpHv5VKo0lKG4weMiZHuk9P83HLufwwvkvwpuAmNxmKeMOcUBZokdSb7AlMAblS
hNEtc/L7AKZ44uDpr+RVFrBvCD+XkuswO0Yx2wOAn8+C0MGPo8AyRCruqaWMVgoW
dPg9QGyLpoWZ4HiYGgPUY7uoS9G1YaNeBSYqruIVZU3m/bC8BhCN184IllMb4AeG
7o2LapuE4qwo/JVrtRG35kNIctq0VyKouxYHFEGyrsXti+owPZ9CSOV/yU+CMayY
bcSgtMPkmTGOzJUhpv6h2+WGc9HdUQF7A+y0PrkaZ00jyKa0EXjQ+Iit/shFUIDH
lRx+onl9L5Bj2r/jFk4owgjxOSs80YY01FtBbUJZJBsv/weTq1nV+d+uQHaPkKC2
CP1vq111oW7+haGeCHEy0qjKu9dj9KGXvelghRh/sRckJ9GggZcV/F7WLcbK/Faj
6dw2w65O6JUFPfeAdCvOUXxQbGayF0NL7PI5dnk2W4nz6NZ1TquCo81nJ6TISXDU
jj5WFp+4aOv2awfBp/129u13tL1A9EmDRDNVwwywRLzrJtvG/Pb5VYngcJfaCatX
OzjUBZCJAT5C3lS1u2WKeteEVZG1sGYkfBcbGwOrEB7O6oygvbIBcKq8Wtqqlut4
6fDvj81Hop20G+Mv0CFDgXA1URZtWSnC5ATLiKBhqwlVC2uys8XdoA7qBc+tR0CZ
Vaer7KPXSmoBcmN6o6aVj21lr6mSWgWhg4Tz8jHTX6it23Fdj10hX9qR9BhN5I6m
ZVV/uXEE/u5acpA0cNTGtG21IqjhzQZHygQNIbiOkPBwH0lnUDcwPIF7QQq8T70Z
5moKmfq7T7U3d6JkUm+b9zoSYWJtwfjqAChPeROmQpI=
`protect END_PROTECTED
