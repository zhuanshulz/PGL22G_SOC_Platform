`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
454BVIqiUVNP/FmbVmjrTvRKJoLHX2n806V6hQP3o+9jBSotsg/M4g5Af43NJd55
s5EJToHOQdFkg6J3gk2BjD5l3vD1+vPNe/rV8yUH7TEjRsJAHbnfIeZWaKMT7cAc
l4gectd1bYEZdaZwcV8GIYonjA9TUGv9u9j2QZ1+qAjsify9vg59YnwB7mTVoFOg
cx8xPM9YmMxD+e8nzWvyfN+VyhJQ4GMBW7z41Pqj3NLz01ELS7OBKQXL6zIt0uCG
lqKr2mANLhmE2Hd3WGrtjQHhhtDRsZim7SBMEJOtQqbF/CAbTOc8EBQmxZ7WxVM/
u396YdiN5jY0O69cxCaS5JYs+iLyDKYt0PqnHVP4Sci7CnEeo3xGkG4z9ePjPEU2
O60U8ANvZIBo1VI5W+uKM47KBhW8KA2Ea9zwWsxhY73DAkUrpj0nRCZ/qpp54VIj
M0hHNyPcZlsLWTf1tdYDiXxTk/8x4ucxd9P1hWKd+BVwEJueaD+PTXersO1vD+LF
MrvRaHBT0cMNqZVA2VoxN6H//3tMMoBIzx+EfudsaRtYOttdct/nuNFc2g6KyBFC
eG8WEQs3iuMzZmQgYsdApK6rnPwN1/apzEEPB11ooVyP/cvg4KnRkVXudySt0Q0A
r3qWe+1bxit6KzKDLcLBT3IIfEV5ofzd2MjZCtRenkI0Lw1lEN9XOTtoGOMlWEv/
nd1bOeOfInPEtgDUwE6dqI3CCYqyIyx5Uk3fw4hJxeKeR3lRBpjIKXJaU/H/CcRF
bE3tbkYiaYFc0eghTWJNBHgq1octS+/G1N0YAHRwouHcL/YaSzR3l3SW6ekEuQiF
BiEjbcCU00deUjey3pBNvOWpPYNaGM+emQxRtYQJC0hato88RHmLmYJ8/yYvFvzw
Zor89fKLLz8rKGVzAI2bqfFz+4kZ/d/m+pM9KA7JsBC+TCpUMJJzGYsZSpoSZfur
3D/F1vpijkES39ltbn3c/Fo4+WlIf5AyN3e33cBd2bG25B7X1VecUHb6C6Hz/jAD
UcDlxjbtQBrbAl7zsJBS+TZWS25GUBQtuQUxbAXG9Uc=
`protect END_PROTECTED
