`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pyil2C0GO9BJwHrbDylvzXS1Zh9xaqG1NZQIyiAt3g6aDlehV4kgXPqj9JPm4u3
AziOJp1BABbyb+4JEJs+RDP7nhVw6/QQ/+i8Ah/rpdOBYpabrfmIR87S3I+H/Xrb
rmLI9NtIjGuKBQEpVnEcosgD2GDM5CvCNwX9tvOJBstvBqT0iYKOT2m/eUWkz2Mj
aGzQ8C/nDNKfamshvvgfMQZZoyzIyMdUx0Kbb6GRygYE0dX9TotFldKVyWzCIwEP
NKDvPEyf4SW2iizugoKOPqtHf99QozWF/pHCEmzmwnGE/0cVhIynjT7pUoYjijQe
KEmIikTFkgbQaG4zfvnCvvpgUULRpUwLDDy0C7Pb91Z2/6f4Tbbe+868+3UdJ77J
khDvHjvIiXVuARghvqya41LF46jiZJ4aajpv/4aNz0iZWSh/x53IIZfM3G4eWNYY
cy6ga7QEtoLfISWYTUTQE5AtWB144TbXBOdxaFVsFRzqUpp9CW4A87Y915ypbogo
KDO5Ogxrsvn6oah1Nhi84q2OliGZayK91Fvmy2v+lwwcBqffNa1+9THgQmFlKr++
03VP4eQbX//VKyRiNWRmfzjqc6Z6NGmNA6vvxWSWm8RAUcZwlOG7dG35HEEWAQRu
vbXnRJG9sYC1rbs1krC59xPHe3GdA94VRaR1uzxUALR98K6D6DMPs2aL+8C3DpuL
iTzFqpSB9xR9CYWfHoxh2g==
`protect END_PROTECTED
