`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5I7wZXF9mCVOlrvG5mI6WuSStOevRAMVlSrc6lFF39JuJPVPpipnY4OBOwl8lB+s
bL8MvvLmQenj8gumCI3bBH85b0DffTJgDSR39EbuT7XzE+h3SMREUozAgz8cLz7b
fnPEWuQU38RKmDnNwHA2dA0vz1fIB4xDKWLVPsHAjPnLLBA8G0WzfAJSngeXtX0R
Lt31TMbqvMRmZiRxRvJVkyAmKCtkfIY62b8JDI1wEI7CIfeQTbhqiF9E3qpGb0SB
uB7XJqhrt3xmd8E7vOdzcIXapLKxDKVEQxuumC1Gf5oGE13m51oLE5RGYTTv3n/U
1+bMt54kXYar0FRHy2d/MxAeJr4a5vmVOGPcmDM+6Vp9B4+q1C7ZsKOMXv9d37Jo
yBcJr7z41jxMuWnJ0g8i908FwAxrio087hnJ+jfQ/nfbmTLARAXusrTsDMd4UUG6
vpDZzEJNYQW7PQlDyU6tT/W2UqK+X46Mud/BS8TtO4XRCS0N5JZa6veA9g2fgOJU
CMRJ+9O7M3tdrEzeFq/aBYmlMo3A82Nro2Z3bZ0lOroBcWBnCso4QlizloyGlmYp
/9zq/FvraAy8E/xubtpG/84jIQI6N5KKOM79gbC3DBXGzUNroleaaHl88hnM52PJ
VqhdPGpaw4/rrHs5rE/8p+oE5aD5fE0k92MfQ/+2b1o=
`protect END_PROTECTED
