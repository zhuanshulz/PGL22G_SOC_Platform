`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E4q89IKyEtRx+L/nEny4hjaGXQR7YzHcgPBqpRS62HKIF/5j9fGsTnY5oewoqsV5
bwnEgykTrOs44kHr5BR2CoKlzG4CWrxdbbgeQTYKVMaRu8sh8wXTjT9E7R5TdLDp
yE79x6KLI5kVXN1YuW40X+JQMdLvSG8P6DbEjHanfe6nnrF2IcgzbpRtP7cCeokZ
6PlWIDZR5Q3XgiBvsfh+5EitOx1+sp/z+ggTgDttwO2sxP2bd3AChZGhgiC2VDqt
hbDgLktXaWpKHL4GbKv3DRZkrm962qcD72Vis0Bs9TuZpGTKemQEDFn9oLsmYFS+
KBOOHrbNrcSRIpxLJQws/Vsz3L0PccQBGAUGVsZXYKMQ0aG69VJmN/I78D8s7p5m
OOsxib6gFEtNApBPDAUc+J9cebnRAqA40Uz2cplyE76MF3bfvm3c/icx+SGIS+7i
+L7lznhVYszeyL/YW7LT8rk2MBI14lUvXkt89tTeaHgWeNChaVT+u+yCjtJLHv2C
BQw9JtQGyDAQNa56NRSkkQ5MkRkXs7qNbLaD+RSEf/H7rd34n/0FqyA9PgacYLgF
vQ/oX6k9wiBjEYp6Z32jvJW0sX+zA2zKc18D0MSlQFFE2Pjg80svtvloneQs8kji
Xd7TauIw8SEmZZ/E3QfxwZcTSPqNYxu4ie0zppcZO4cnleyQP+gMnZaI1OhCQQHj
VMtx/d2/S+rglyhNkeQf5P8U9sF5uzT53zgrWeNAc23FZRXIyS1dWuzpqRw8P3tO
UFSxCh0NG7ky/BZXTAKY+pPxxdWoucK6yr9FEvclJjwG500WoT1ExDQ8KszYSv+z
f/UO8yDpNA5xv0/g7Mba4KBc3X8FT2L5gOz79Z64IOozhSllYyi1RthgmcyJVQp2
OYYUHPfXDdU9qsOZNDhqq1R5V4xqxvnB2FnOYy97nC2AKKQ/WbF2tvtZu8RtIk2k
iSxqviqi0uBNprAfOzo63Q==
`protect END_PROTECTED
