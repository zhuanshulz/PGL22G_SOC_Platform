`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NEpVPpa0ij/dRV/w1CgzfyzzXI6JhfDAgb2eEvZdC7dgnapVemPAJBqtH5xt6bSQ
bBRuLFFzzcSl/2kB/uSGqOwbVSQZLAUTU9hLxpcJFn5XE4/npk2Q4VejbDOfS/Uv
2xrOLuRCqyOTaCyvDZRp1icocF0fs+cZy3hJ0Th2yJ4Px6DhTkBEwnh9pFV/6/IX
XO2z0klqVgZrJuUohfAv3fAVCmVo+sBmroqaWQ1wUYMB79JY9h8HxQ4KG6RhvKMQ
95aozq6vniZW3aHRSxAccRiwrACT4ytZlJ72vVfgSITcstF7lIpfmBCns/TMJinC
CkQxDA/Lb14aSew2GsnQnTAE0DTUWXQV9Mu9hruNYtXrQ7jN7Pk0S5qgBwDaVU/k
cFRluVHfBVYV3uIeLpI9Xb45mb2OK8tcPBopS91eAmM=
`protect END_PROTECTED
