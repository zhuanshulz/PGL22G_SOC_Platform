`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OxiqKu22y4JnHlQIcDhZlMO3b8QfvYVEc9Pttqbl2F4ak7dHLEd04g7xHBW2P5t6
fY3FPgUNzKJ/CV/LoxbnJBcgWunPzJ5tHOc/K3sM1LUBF2jYLO2xpLHHxRu3ixmD
b91hycVZLNd+2Bo9TMMGYUqQPDX3mp6m0TfA6u8xKw2UQ0Hxm0vJfz0c8RAyw+8A
XdO2SWftivJlbrHUcrm7UuREeopauhg+h6YpWPf4YniqiSNQqyA7HihIxYiARk9v
O9x9I9QOZt1sW9/GICEmphpsFzoRFtaztvwXjnpgE7IYsZ+qfhyLkE5itzqMCPXO
x9JoC+JPsycgvCZ+KqcAdnRGmeSqPMtpvZwZ1M3LGjvmfpCNiU9640i6wp4Ke4Eg
ABKb5MAf5zYCODxXURen2kffBRLRi5s0IDxe/m6z/RbcT+IeeJ+lUzqIl1SomPx+
zh4F/nv4UkDcHjavfV8W690SLSgefn8ZIgloyiUNBBm1L113o97KhivCCdndXC77
OTpdrGGk1bSrXYr4Wdlr4t2T0DL67/2WgE0hJxmXTU8UCys6wQew5YkziJUNuGSA
5lxCUvKBDhaxkXVuiHSGDLnWYIdGUdKc7JxweHrYbylHoPJp9T6eALjzgCbaX9GY
gU7kdSfbGM2R8y2gdsSHPWI5CnHXyTOrDABYkQuzjLQC99EKXvjp5c7ZO4bQnOP8
yrogId1cTRs2bUmcrsC7rf4YJJloLgu7r9RXdzQvrMBHx//+WnEbBDJD9sGNUPie
HfLvwzJppuYJ632nCCJm3lpUMDQ47846zrpK2V5BQq80f4RR7tSH6h+O2EsJDkvn
S6LSQpA+N0V/F3ceVIVjoIcsOipJoYx2kVL2joViTMHXES+FEz9ScuN2HbWQ+6j8
QkSdcdNOYwpLPov74hUgNnPn2UADb4U8i4MH7b9Gi4nHW42hY6IK2SMwPCimn5r8
oLTNJcQhXZCweL23bSrxkb5J3zCiNd7bMF6+QW3OgjBCrlHMG6je6GDffZ8vwnWw
6Javco/iMTxbSyTl3jiRDk1zUD0CCwSVINcijAUHGMzIO2h4zYrFL/+NtePUmnK3
ZQBTJwIzEThfNKtsWizBxOyojLsJdH8e0AzcoiejcNDHy32LBFhWwKXimzi/wbyj
RGRe4xls8UyKigJmBhkHGSQwwvS7Ar4w3y6HwyvkLnkXRSKe6XFVUOxUkLrTFqWs
cq7Re5JKy8NuG+HJg3pEIQ/8saKzOr03iq4CQhtzZtZ0J4WiqSJ0YLc74GfZOwF2
I3VYT4Ql3jc3NcAsovV3pWLcu3v6OhUjv734ckCK1qIdWkXeax22Wml9yla0TA41
t73uw4jwO05KTofVFI2IHqPFDa5qum6Ex/Ld4pUNe/fj89pxRGiAUXR1sc9N9+83
UyzALEtrxyBLEHkD9SHhGq/LyL2s4LMy3pyibPNHtnLr+IjWR7oatBj3NJI0ucag
4UJxmE8PFvAOW00TN6adItszqcjgCeOLb3WXGx2vbm74Y80GA7gIs98xgNtLfVyH
DgiKLsHdFdx6s76peG7I9ZRt4/aahHEImPM+vsNUJpOTpVsvQeJV6+ZG4cizYqTn
HkCe5dRMGoZsd3CDeS3cOksf+DeI/y9ceYLpt+S/IK+GOadyDiyEvLzFVzDehoLk
rFD4mq3mIR4O6T0mafmNYuyCTOjwWwAWTfCJ5Ds0db14Afc4jEwnrT+EDBUtEXjx
iTsXoxnnpgBQedZAu2wEQ2Y2IFZkL21qTNzhmF33TxmRUN+y69cNz7OFYIb4Z0Vx
xbrb2WXjiXP777cE2aGM1Kph/Aut1YT3/YIu036xoekanucB4yZTyGPz8KqoDRxV
QzvzlaA7QcHUxtLNWPayB7Yu3xMyLHydj4Z464JL0sqDWzYiRYRQtMTR/KPbaqR/
2ydmcDUHeHl5+XqHbYO0dbSOFCCTN0v/H/CpTfXATPjryo3+ZZtqrxqjcFJH+QEd
1ii4dov/i4KathendH2sXnaeilTDQ3J4osVy6zNIHMagJAGSutQCV7/8h/Pa4Isu
kPKdITHNpaRqVVnlD4rrn9XBQEnSU+EEZmFFWAM20aUlLuiiGVsO/MnjzdC+JJ2K
l2lCi+ErYIgohYtp0Gp+dTNVmwwUQNNtFBqlPhQHw5ivflL6L0mZgVdXFGxJpmZI
iQCY5FlQI7On1zpmmLcgDevi6HS3hZ90n6uV1v7K05f6jA2/blAP7IWV2BklBxI6
ee+TYMQVCDdrt7bRjpS94kYVXo2tz49QAK1FzJniywFRphdMBmt6nTX8ctiz4TIC
hfBzRhHvZOHy6Nj0AQTsiPeDGUVMmtIfvhBM6MLWMbWTf8LJvm3/IWxLp6Y/5Kbf
eu8oQc7WJMzYBqNXqgvxDjPMiiUyOZWOEXH1YsRdaZxrUDc5KzzC3XU1llm1+eus
g5Fm1yusXCtpuAFG8S9w4hD6rhCw1AVsKFncr7+zttHkYI0h3hYKLGabcw1b0W7V
y3HGioUgDqQjvCMo/AX8fv897OFmqAF5H24d2D5r74PiFRxsELXDt56eGwmnxGVG
ld2vbckbMB1p/It87UPuyVsYYg3Bc72POZbDq7njYN8d5BYUQSSBwZ4CDEVCqwKz
QJbtm4LcRPVyH2ImBzrX04XqwhOYWy6wQ5kwzh22ttMo+KlP3qrXOOO+yEiZ2DN9
EfPEXLf0qEjYt39GvXxIpyjTnYW+UPu9uQxfCUejb+4QPH6v97ebUxxY3o1ZtkmP
dbO18dP5gFsztSvGXeTZPzAyCN2qkSWTbErnCbUySqh5r5l1nh7GJ/WSHUS9HDCn
i93cQG7B2GQckDJ6LMBfK6xtk6R75U+mAflFXwx6io4YoOvVA01VnUq0ZsxQ0VsB
EVaCs0vcpE1KKxW68hLuSBvQiDXSTigdcEQn+rt18O9zeZe4cPYvABnQp/67pgIS
YxowPuaFsaHaPOFojWByAgOxy4m/IppFUxIZQoDUs8yw6Ik+slVaV4upHUe9bg49
hXjUv01QMI18F7BIBKWcmVFIDG6aGxB37w2TAqBun9XRavpH0lqqqPG0yVXtiuxv
+ecmkRuNVe5LGTBWaA/0fl7Qe3HmuNQxIy61DFX9fYjBPJeETxUyClaXKa38xyEh
Vg07nH8MwP2ZysNK/pVEUkSFG2qFEfDO96BAUIM6uoScHsFk8pb66qATmX2Nj/ao
qUS6dlXUIQSPYeOGVLH6uPNbf6mc9gr27YNCKn3ZKIkl2QomxaMl3hR6FRsPWLTh
PNNtmFbUEcpufCNBp0xRfwzlFzLSyiPvcTrKB8+Rz6NbtvOIFudHbw8bah+AWUo+
85Fu6X8QBjRN4I8PeZipW2r5GSD/8KKDG1RAb8SiZx2vPNSN8TFpP1OkwMxsi2hh
wvzRrKwqWMoWa7SmIEH6pKbw14yE2CB+tRqJkt+CdA41KgH7S6aedTFG1aYsJpGB
V1rnW7qad93DaI9S8yD0klNh0CYWZqPAPmaWgbblJUW3xaebCHVuPzDDnE6fVWqq
Ei4/29dBqebukjej+6bWcdmT1f1M/0MJ7lRomnqezntNDtkqJAa2HUE0Id3p0BET
terGPEV/6Ch0Czb7Y4EIzvZtFabqVbo7lzI1Qqm/b6NnXvAzbGXmVVd2yX2QOQMc
5py0CvfhTu7IPlShQM3pPk1Lh7fTWiw0Jv8ZkKrCTUiMA9PVtTmo/P4YlOQ9W0Op
F+NRXObts2cVHtSj1ljpkcM/sru2m/nxQ+bEXzwfnMxWwFNhN2hhNbZFOrWXad0w
xwyLwULVGayrESQL+1tzaeLaR4bR+iVz0oTtJk9bCXA1cLdAmhXXC2l5L6BCCIOO
D3AZQircpNyyQabRhigFx6Qnvjd51rmUEu4SdR6F3Yo2lAV2uz1vkAg5TxIIndc9
Nu+OETYrTEXErtS391Uy4nFyLmCaaBBKNb8vZD0FX9zgCMv3JX+jgRzAVeA4tNtL
vUrT3DuxIXGt+fTfAJ941gpQkjAxfmPsHDZjPzNDRh7L5xMDImsDO9mcGgNcr7uj
eFSZbD86SP/oTh6OZN+CsyYy6RlvUer64IcGz6Bfg4ppLKAE3nCP6qiSJyepbDVS
ExriEberfQVKmpgIhWXcc52yUuOf5yMTaqkH8+xOhx+LCWVQld4mzyUI6K7v0kLQ
K3PBsiYoJ2bT9bxGV/B3Sf5k0VzjFrl5QO5cb1QSKmQfjhFc+Hj+0kersC1Dk9fC
3pzANFLmk1//XdusqzF5DQuIHXgEEyWXY8v0Ui8SMjRloQq3l1l/2G7EoKhlyFPy
jzlnf6ueOijHjoQvkRfXRNkcuJnNC+fKwjc6vkROjNdHNd42RS/ZXO1Yc5R8njfH
pO+5vZZ6VDNtdKM6DAWY4zpWNf8zmRuEwsCJcw4qCDwrRG+5fYkjv6gvx3+wXONf
GKujjcuPjwErRF5WUX25POboGPqjCvjs3lI4Kh0Y6PQ3QCAUaYbdaCL+HbKb2iOT
myytooB+GAhd1/3xlF40AaQdIsUQuUae0NvISFEqSJE0Sy3tdDckIr7KOOxTl2J3
vfv53BkBdfX5po8KnRL8DKl/2Ng4crZCUKIrn4Q1RuZxSHe67lB1LFASLHZu9j5p
Y2oudwXU4tveXEH6tZRqYxEEtsQ5Np7PTlJHrCdnyiSB5WLLqijQeI8cB8tFJFuC
IL3/GhVBQJuP7QvpQCFchXN6079Qx0QlcpRHtSvb2qPC9Uy2VZw6rRH4Xmr+f3GS
3beY8k5578ArfQcRmZfUATgHpsQQbbNKKl98Ln7XqETkggx7a4tct3aP/Y8fZavW
dUBQZ+8eRC9RXjvbGVcnruQFWVulNQB2Hjq5iYB+Nv2CoCqRtErbAnI8/CY5h1Gy
0GZ6IXyfkzBzTCKyI5j/+FJypeNJ7n8cr5Z5Zy7ZqeASqpvO6tN3H/Lauxdx1LQ1
vA++iESG3M6Qv+j3CAfhm73PIj0OhbsZwr4B+F2X+1bMaTbkMvj4qhtM36Uzhboe
/4JbV1rM9tmKYJWdsLiX5x/yKsLmkEqcSj7iH0WlqlqAe0jJMpPbUbyYuhe2Nw1O
XK3otZKHdKQtyb2JfDr7a7yiBBTlTVlpB8/wNhu2S83vrdN2Pg+mc7ydln/81IO4
yyV/eAVfZVlrozTHa9Rh841Qu5MVG4sewaHIhWBNtLazy82sa4uENn5nPeJm2Fjo
EqZByZ86ut5vL5jPIn8ltIvE+WasKDeZ2eYKOwQJ8vWg4ETo+fuS3H0IH0ywtjwH
Ln8cd6JQ5/DoN5aM/C0eOSdMi/6QxuSHdsEhII9En0vp15QE3dIAuEFexyUW0Lpf
87002Wf5SZhoObyaQ+OOVefV2cmQQjXWeHXNTPUZZbmFco4Y6w2Ci+2yc0yY9EVc
6Qd1JSUjOMKmNP6x0dgiiJHKe7Lc8xqRxgk8UxKCdNRBrHB70B3pLSAKZKQ6th1g
PxdsyDAzddy6BtvtT2TWxZov5tD6pbuFRTog1ugws1aDep5j77Gz0OkxtHRDvECq
9wljOdGHsG2CunBcbI6B1Tmen8Gb4bJ0H7m/yyzZ8wI4O+SKr7iy/5qOI1K1Q9uS
KzjCaKXlirZASzeW0hXO4mfhRUJpN4WV3XlTFdh1VS0N7Qiu9D6sh8+1G+5dfJCg
d6VeuURsk7uUqajEj3t+TmNqu4r1BSW4FGtgKZYKxwq29otFzMuYvuDzd9wiy5VH
+i42rvOwa25FRptNxLTPoBDWisaoOP26azlK95pbyTdUE7LZMfKOq8koMAIZZ/DV
ETjWOACzaYJ0BepdBzK5y7SVO40r79fm+6+APBpS+J4+toAHCy/RKzq1CIuxiokm
FgAS2UXDPV+8kff5zM6UyQ+ju7aqFuNvOMnJ9nAGH8/2zqYXuP18sEJ2ydb0LI6a
L1H6p3PpVJH+lolrvdpsrBiKcjLUrTixlAjEuaSAu8WnE2FLrFBRt6dd1wKpMahM
kWVXkNchcBUoAmMW6GU/+Smt84Ijtst1zA6G2Aas/unzcxnHHspaL6p9/LKtoRhq
tVpEiBD2GNMeAqeySzXCNaCmakklccBsrOmisFQQV5449eWqxQ8lvgxMHtjJ+Z7s
RCDvGnpxPrE2P9tHTJ7r5GSz+VwN2odkNEzkLCNyLo737Bnr7UaGQ1/NZue8Bo5S
pHKItCqC1b+PuP9hzKE1IQ0WMAeEOmsJbVf01lY5W1SwAndZEjlDKcogjwhiFn0p
5NKQD4j/kf/jJlrqu0eKCkbgclbkFN9I090a3bfAEgmIc3iu/eZH3i6UDtvuvR8s
y1lxkHutE5sS8J0fpASLl15aJTa76xq7sJ3AhYlZdobJATINaDoQUQ+WeYTR3dZu
rsy7cAPpsWSww1bBMVH8RS1L8t7F9POpt5VAeERoBxrcksDhWzu1hTghKZtQ7/jQ
rv0faEuGTWYdNtBheVuzadrvx3HbQN5zK6i0vc20w/CMXeqzfsnWtV0908YPN0Fd
0i5c06DY/fQnaB/lF27g3w==
`protect END_PROTECTED
