`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
po9ZVM/+je+ZJQprvcfJgSMhcyZd3CiZxPdBMxdK2V3X8Q+paczU4sGHLsLXh4jn
sabYLDOS/ZTi0IlN6lmkm+4DMtqbFvx8UYHk6At6eMdKBEHH6ohflAniuRCkVg0E
FS40A177K39toPgNVknUwF/WKgVE5k91cDaT3OX6YBQE44NF1NrmqpQMHAg9A4pd
u2XHRTBsTx6oSYOCig0aea8Tuv/KWCco4wIqbePg3zlqllGMfma6AKsLAT7bzN+K
1fXg/1h1aMmIa0dE0sUENr/f9LK+YwuoqxSXWS77dyCBtEgt1KBWIAyhoJszzlYT
CyihqBGVuFBCBKsXg4FSURmzCOBgccxUDGMqdGhHTuBuB/sXv36HX5rMr0stAzAd
79cmH3hsQDhLIztwLOBdBtcEv/CPCEkPQ6RSBX5paQDD395WfYD8uTxbyJ3r4PPo
r40MGAT021wjedyykqrTIjNtrEP8+9TaYs1ZujkQ8SjR4+dciPqE3rF6i0ZaphVf
q22dRr+DgQr3r9d3WX9td+U2pK9C4lAv9Cfs4MuAzkdekspkT0Kcssg2OehPB2Xk
y+F7/ntYOV2YvUd/jSXQr/tp/ad4wpiquS+U/SkpQz9qvttsoxkNyCUdLBH20z6u
Rj6Wvcx1KUhxdcdhPc+fhoq88ojhUawjS4iouMcIUArlHeb8djEO2b/HWqEZmlGh
ZcJ9ODKs91eZjcIVCbOCEL6PCBSRLw+mee+qo683LENF5DpC5/P4IWtc560m1BhR
J3s9aYUN0t2Xu9TfN/WFL+kfnfMTouGsf1E6ktLCARnvpT2mRkirEPVNA/uYJsfZ
mzOi8oKUs7qs7uRGhx0U+1DfR0AS3yXuV4xZqUrrMT8=
`protect END_PROTECTED
