`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ILWim9MJqz6Ru1yhR4x5/u9N5qOlZV9FURpfBneUBv60l1mWL0Ua4r++aMKLxhO
c9yPTcOObkuwZ+TKqIzP+ZVQeHJffwaieRMnFtubGZYhYq9eShFnnYiDUR/Llbc5
G8w0sN0NjhnUXTXOAodg09YuRHEeoMpYzvExDNaWZAxExkmwu8X0Zfhatw8l4cKs
EjtSNu55WAww4kQr9qWuZ26mLi57xrgicfDAq2Z/NSwcP0gv/LWZsgYx2rCTl50w
gmJ/tzYa19opEiCp/4Q3wVoWkppVmIB6XlJQpeDGjEKzo0926D9RwjHT40VAOtGV
Pgiz3Y+IsEdKmSloYg9udJWRL+pTolrBbv1zEb2DBPlJ5BW48S8ZHK6LWu0x+Ulj
deq4/ZCbOsXv0osN1FNhCkCLcsUWW73J0a4weu5qaSNnaACxjwSW/M2D/8NA87sv
pXKtXmFphn9NKREoo/aTpaxLpxpRdEZun0kaFuhpep3/M5vQE4CjSP8VN50Ajvxe
9A6ngb7FsvrVFleNQgKSntZ3FU0RJ2yJeC/bpFgauGn5eHi+RT0zUvlSZQ5LKA3R
5iWYegfj9u9LxfWa72v7pTupG4A02NIfcSyqkxqpT/yJ1PTmduIWlZ9C/0jUPKZ5
XDgLsfvbNt5r7GugRmx2n8C3THEB664TaGnjmt1w58THKpyn4xF5k0T52iF5LAyc
Ix9yVEl8FYREb/voqCj3WDCsYKm4Oa8e6NQOFit1lNNvwatu8UPpaqp34sbpXyXH
aEBYR9EAWIPl/hQtObls0HJASd8+Je1BHqUJcCyXFfCnjw/C2Vs5G+ix6Pn7zELR
yksFQpSfjzazhIc0KrA0rblsQSuSZYOJZ+zOa+fAR4YfjLBsclUe5MAt9+CsGmwY
caf8CilewjO+eWvJdk/4RWqdWSi4O3p0CFLITBeggHg8PnytEIqXnDkf8YgXGT7s
NdZPE7Fz+QXzn6Ry10G6JsxSaN9tJQB/sVjUMQ+tDHcOHNkR7sUA7quOWo+JWn1X
jX+cHmbb5BcIX9CrGjGs4A==
`protect END_PROTECTED
