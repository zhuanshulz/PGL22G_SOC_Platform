`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/77RzMrB78KqZ2obLIJTZ8yGwK0i9xk42VIYN8pHOGsW1LLyV+b5Dv9/phz7kDy
lQsBYgoGLzPH3RgSSFaTFYzJn3FzG/N45erzWuwzAcB8I1ePgcwtlcHORj+QcCEi
KD09FfSVwsbHPVzxPT5hPhzOZxXSZ/wfibdghdUvlaxn2jnGlfA3+X1nTKIX47CL
9q93TUtlbW6HMV7iZM9Gi5403cbqMwdUGRg6AASpgDuf/Jr1C/5+Y/OgM9kZju6D
k2z6hwSmNzjO/pSPUC9hYDnnvsaYDEmej3GEg6yJ6pBENwVSGW5AMNNjedetz+Pm
IXi1WZPExlQYXWztWqutmRZXTFwUSplPK1eju6YEK5MxKYl00oOkdU5p54fxojH3
Z5TXJs8NN7s1wgdQz9/+HXmydPlVM26ISNFehx9g70afIefWzXDWj1iXVVJDMyzx
oNEMk76ND0vZThCfwMYAtXfjnqjCgtq5ujO+qo9XuDCfg4a8JUgfTJtA7687gb/i
o9OtLnkKq+MEHtxnDwSt/wPEYXeBszphI2G1x6yO26yyMTAmvqkQLVeTbIbJMxLj
CEAiin8xgxdG+plk4PkghPYd/LA8mdKsgIVrKjnaFA2OgMO7IjQK36xUMg8I77TJ
cCUvCDFePaOAGg7ErFpt4IPiYDUoFcqhhONCfWkfCHpg8bDAfWddl3pqvemzWSAa
UKkQV435+t4rPO26hb3xr1oQ0zaRb6uuz+/MVtKFAIsSzrzVbIkMj1Tn/d4VG6xP
MNQrFZqEFPAAsDp6t0AKsmtOWcBqJUvfqJhEL0UkDOZ4iLt9cmDMwmpsQMQOtgAm
GY0sKrA9iMh4maguTNTdUsK2q9sRPEXe6NSwjXzGnw0i3rZD0bdIxdyqWe0Nxesh
4tMETcd+w8Z9RrHDOhXHvExswswhV07w9U2144P4zx2EZcDxGBD0Qn1eykJzdzPp
BvDEDk6wrjResLgAUMkvQrmoWXZnzQRX3B4eFHhQuOdizofnW2wkh2d9U355eAA0
xAksGrIJ8npf9nIbhnbmn64XkArmuBRV0vsfhgWDa+UNv7vU4e+6V0X15ghSxJxd
2WkHdXNBTExp16vANP4SJM4OcyiCYX2Kxle47dguvTX2J+DIZFT0xSCYVvJAqXhW
wpPvvVQcuxC4jsB10I48U4u8YcQQETyL/Z20YG3VDzzZeXTE0fBcxBODDGSsgAP8
OF5o2oZwqjF1jT9kIne88FpVc7LVOAr8QZ6DpiRgI5JzsjuvaKFQRUiuYTEVx3HA
ZWjDhhXeYfspxWAAoJ6aDyLLyGt7vuu2l/+aFZ0/JfZ3WDziZwKKmRDuI6mn5ita
d1D6EWf3+ViSqRER/4HdyUKMcReWA2wq0TDas16xUCdf1ptjrAjyzP2dLuB/05RI
YrfmOWxCaJl36e4C1e9kUDf4mktzQ2crvWVf1uKTy9oZiZA/ZrbP0akrb9svuwFT
6VqJA85VjxQsxQMfcF6TDSwhGKrfw84jrGxsqVdTdl1VH7fBJdoEKnJGiR6CVaMG
7Urf+q1iiDpVwyd8oDSoEDWoLWZa+WXx6Y2UGzw1f6uNRC+EOIULOlgHOqGlqvTG
Xzd2T9MCSn9aITXfobDYzc9IBz1P04YzAscSL/h41xRi/vol12kmnBUi2ps8M+4D
bbDvO79UZgPUym4ruvPCd96f4LK8UyCT/vBK3xljkjBpcrJXCy+WXdUldHDrzEbJ
gdSUzQIk6kYKbD19rlTztsmHFzjH+G6TwdL05cfg/NAtJxzvDUFZjT5sdABFQRr4
46th9Y0T3jK99/VErgYIcAbw6a5ZzSR6blZuGqsrJ17c9wSm/NmWE6vui4mn7a6r
ZaoSBWxT+3iqu9WvoeX1zVNDSBU/6HT03TeIMszV07lcJk3s8QkLxhMvLk45Hok3
LFvLGbpLaFH32/iKN6TlxJK+M9yeeAsCyigVTIJk6kzfJoV9gP3h5jpBRP8YpNVg
VFf49XodPmWOCg6G4UqjMn/i+eJSa0cdndzFAyaPvReGx9VIeXGTHzWuQFcQp3i5
vzmlARor3+ShpdCrCZzaHhawmXiTqbV6c2eHPLTGwhzgfeiO6yIXtOp9O8UJtrQN
0OWhLVfq3myo1XIsaZ5aYR/trT6Z56Rw++AfpRfAL36yNtU7zQwipBS0zdwKWxR7
k45I6G01WA+MbVAhh/h+K30ctPesuV1K14G0zOriqn2bbGunTL+tHFBl+c/a6HxV
wYHh7wmSybOLm64ESJmAR94rEUQZegzZXJMdvZU12WgCbtjre+0zw1y11TViEMrF
NnqTqH55fEGIj/lPGAXUL8F42xjoroAWqr4HFwNxhyGJ+lo9xrnatH9nCrzk4xNU
CUgjcjEjM8QfIPkitNhsAkS4q16wtKqYbbnolntMiKzzQaTJc5tnbTeCWYECiuXb
kgyL85m6QxBqoAq+dq8ckiZU0H96+J9jqnAY/sx7Z/ZyAW3EromrHWX8F1F+zJ9k
X2C66Q2r7pB3xaUVccFFUxJwciltmCj69wkFxt1Hk4Nb4B0g4rtAKUzesWKowTvB
Zlqm2w0FBl7hEbrMUNw3ny5FRfsjCEMBMY5oZgLVM4fk4aZNHka72cSBLgIFUeji
SWQCvg+lgOQGpYXfFphVpyrTyOrRwMoBPYs0WPyoV8v4PpE1N3pYsd7lw8VOqfDb
uR/Hh6+9Bz2eTceUlazTpppOT8lgZcLJHIvRKetq4g9lJn4jWdXEPWLYqW2ewvfn
x1RjlOTGJzvezvp3ZL/NfJDBJY798XX/nDQYE2LDIdj6uqpVQQWQNUIJ6vHuyKyR
nuUy/FY5IrP1rlZTI0kJ0a6d6Y5n/mPRUGVYuc9V5NPkCYQrffQG4vQP8xjzfk3e
/Zka1npkGnRmPLuXZhvkK+wYyiPuih6wPcDI3ATCO2jydw4Lk3h+O1+sxhYZFv+T
ajas1fiM/6BjLl/m7eh4RkN0rAEQJB5W8VCDpiyLdtVLHbvBqgYrgYRmZKkaxgc0
dvjC2XPBGVtH8mesGjfY4iPfCv4Gdxk+T7P9vAOSvDzzgIMHxMKFw9LR3l0qQUKL
yYz2sUJivCN/2IqyuZuEzsW1NYrcOVqfumJgr7L7sEGoXcllXSuzT2Uz/oj5wX3i
PyOHy5Nhxp7g5ap+6bV/aNgTgiddqt23tUF6vLpsZ+a5TKD6kgSslIvbfoSYN87I
EwHTvP/XcyYTZlO3Wj8QTMddQnHLe1FXDRRcWgooOF0vpg7o21CFu/NahtRJhkJ6
115dIyaj/TpN9sbh83xF2X+GWX5+dbmfuCIBB2ywRuRiVXa7q6FqlLOan33NONEl
LMou/TAJdDWbLdAozwNLQLqVn98+Dv0E3QUlw7lPlDbAFbef7PQpRUZbQq2F9JbW
HSs9UJ9lfnlhrxAHp7h37FGtMMoaBDf7NCOvftTvpB7UeelSmMjIUiqtKc+uXDjH
WvbNZ1pPot2AzE6iQJWIsCPnrX9MTXYwLS1D2BK3rcCugiIxgC/RH1Sid+yedvf4
JZIXkEGn+Euno+K/tUGfBUQ1JkXwb7S1FgJ9C5jQsqH3SyhKvCZOjq2XuZ32jvRy
0b2rx5A9YYZuEj8/agHt/rpzUTFNsMQxmO0i2JJl8oKjCwmUKF3F+felsebxzLrP
T6XL3RyZl+9wv1VWouFErzDNb8m4v62RdW42QT5sYxvdaWFlueDLEuTHOQQpRFI8
rFWy3b4wrtipdgRkgVEBxoee6OW1OW9Z6mXi8jrOVwzsoOvTb71PyPAoPWzUQwYJ
gU993HVqC4mhmLoq1CVkH7/6IAaH0K8eTNauquZPUWb2jrH+rF/rcyrMAmkY3A6y
jVgoizv7dBWd58Jzq5W2QO+LfYVa5+VfwzlcH793Onjlf6n9WX1ReCeLNrlPyJ/s
UKaSH2NejhWYobcC5+Ob4Rn8Zpj5ccnf6GC+0nC/QrL/dh6JJHHF7bQmrdlnwj9H
qt5SGzNCggYM6IKDKaEq6rqP6Vf/Cvi0WyE8BhKD/Y2rCNhlYTmk4oj9qDFK/rSV
EgC3CpNrMccUBKRxSKd1tBSb4aDtBTurox3YE/sOOtXOIQP7jUziDwKKsPHMYfyu
JgBOpHYRbhFg74KM8LMtd8AeqYwKca41MED/6vB1BOW44t2O5FwjDBgUw8wqfpFF
BUkFfRT47SP1TEqwdFH0jfmf+pi6dGWq2uCbYd1WHObJJfPSEaFMKT52veSV1Bz+
kunxRed8GIS1b7Z8MIjgDgnB4HSB1N7ztH7KmAgUYCNvneIsO2maxrwsLK5ZIffN
M6WPRjIqvbX1FlKI2jZqQJDd6M4YNvhZsqe0c/uB9cL1TTYrMuGNewbmJ+h9BgrY
9wXgEWYEO/rrkEHQwI7TSYS7EMXi3m/CtCgiB4bBppQ+Ep6JHhPUbufnIHvexe1K
2Q0GwjASsqrTi6Npb/5FNWJcd8etF866CcSa2WlfrWkjjW91KeKS9tvEtKH8ejEL
yBdFfbutxwn5XrRDBh9vwKAHO9zck7T6Yub4tRQAqdnXOXSj30C73PxahQwO4sSA
YnenokQH/cFnn29Eix76GeEddN1tcRQi4Xa3lOY9ZZeJhTZiyVj51Xi+UzHjV5Ba
B0nwD79iLlDcrutrF+4qjsA4ER9Uxvp5QPeR7EsjboKoQZFr3o/THvVocjb6dni1
R8uFLfK8CcJ076lLsBBgY7EbHw8PJ3awUME5OvP0F5Z+u3AHaP9zAfK+AbSmOBMi
EMO/17FG4oRQCgkS6cifD6tgwdHt9+8oQ54F+ay9ObVx2QOQ6qfn18yUIk4JwZLM
379qqWkdxpFQmh+SEx77fA46yY7F7GHNInoBSJ8l+01p42qxxrJCT0sQCNR6HKwp
Bz/BGVqQP/4XflarKcL3gqwiCc5mANvZ8c+XbtAqkSWf3JejiiR0yQg1ZAoZMFyM
tWl/N0BKtrjmPWtj93Scp/qeWJzbpqmMOicBWOG9U7V2e6pwK+w4ZtfyoTfHy7UL
7mBGiC+jy/g/jRjLG8yVV51xVXcWRzCaWHnD4avUt5v2BQ+g0DnVqqDoe2hbBSxN
NQKr4c1NhUS0OJ1qcFNPPlkfrcKMm1EOnqWeoDnQQz8RePZZnJGtmuW/d7RZPN46
MRFmWOjMaNJTbRU96uplig9puHZ6GgoTSVyTNAxTVRMbPyq6kYMTOVl4KZa1gkPh
4wSNxgalmwLACEPwshXkWSRR8C8hK679AKSV0zJ/kHyk/enHj5fVr7r9Zvg0AebN
mWEptt1qs1SxlEFPqRMwQmEComu3Oevfm+uXtQrkyaRDj67edE27m6TEDHgpRJtG
HrQNyCGepI6SO27z3li+I0jQWicER5aSA9R9UHFLlF3vsdwmw3sVbbqQ4eDaqxGF
SMwEmMmJQ0LQzXp3yWmm6l9rkWMLgxoIUcEGjTxzNNG3pvuSi4MDrUA2CcL4jNHM
bnT8NgOuSDeFg9/aI7iw926xVolEP0fShHV5Yzvv3rWsRNP7K2QxOr9y/PgfWG8+
6HpohLz1U/pTgCXe65pxPpEBfh+q+IjnmjGpr3jNIqkSmXOUVFPh+L5CFpvJW7Rm
X70uSw4uP2InIdDjhBw605/UxmkYZKkj2V4oCEjqCiXjGeihXzuxpakMacj34XPR
tJCC9jjn9d8Q/SKfheoS5c80rNA9hCAqv30SJG1xiDNs+NmVaxFZw/KxPszBAkl1
v1Mxflm3LhCIuSXGJnUVMSqJcJ0LRM1PMTV+SmM73+/1aWD0uNmrh+nPJjFGNbOx
hCSuMvVvJaw6kbWWGK6Y5Y+LbNRYECUV4Lj3o7xdeA88c40OvrvZTi5cKS7UD0vS
VsYFxy5o3ZyNj73Y95II7QHxQcIInIWSalGg8acbcILufB2NJQ0eDtZPy0pegAvY
vODzmNPhUAnFSVf4aq/dP5jKVZmcn/eADziS/UBvn6d847jTM8PFkNDkXgYqdbZ9
GemTmu9dAkQzuFk0F4VxRbOrYdXIQH7KJNPpQ3Z0fBnW394fzkrjIyEgX0j5WLLx
Cuklb5jSAkViXzmA0YOy0+4TSw3RoNkW1ZAgfqImGAYiDhPE/LKgqSGsqqvxUKyU
ZLdT24m/fcs6vfJ2IAaU2SQlbrmuw/1wr3KIdoi/xbxJ8pBkFkVBhN6OZmGdc91x
ym/AucYvVvhQeI1apLJpOSfCQHZ2RdyKAifZdpXPRBV4booCFH5OzRmf352VspIo
t06mKjE2uvAf+DbkrJwjpI0vVD5NRj/cP5JC/Cj3Iy1DYtiJ2ZUfkV5pBRXnh/5d
utpBypTLvXH2TxMSVb35ohGHSKYyi8JmR5oSJUHOTISqwRzzndQ0Sbw54mTNMHJg
ywWCtuO9X4xf9cQeQTHhZG+sfrjd1lZqBkcdXnWu6TUouXcEdyC65tDlaehchMJD
zlqsY8gI/XjK9FnoTlHSQqEF08ZBJVBTk8RScKy01EZwWqov7P/rHQEUIEb+zaCw
na3wCq10rMt30Mu18hEQYLddT5E8ODgenKVQvn9YZa3gfTtMZAmZQVbTnXGxaG+h
P67Z85YwC4lWnRlxVczjGI2vPF+8bxT4DkgEy/CgnKw6cIU/NrZ/CHiHVZkxC3+z
SI86NP+O1kxQuILOdSqjnIErcBIqrOe0b7Qm1EjYHUZXJppXDr/5eUbECnz/Ko9H
ThI8azBZ/iiQmpn8kdiJH3gRvRr1bvxKLC9ezU9uIWrfB//kAAUHWryM3uGCWeoq
l0GDReVyV3yAJbu+SrzVsz6C2tUxPamSYnAZmz14HaTfnepvNmmITNYMjyYdRd/z
eY4zE7JuzbLQxJTX+FIbnHXjIo2JDXO0LMmACxeSD9feSKTo1e3KcdljTXjPmte0
olP9BQnhxtalcpz2Os2TlMpbZHTOw/Vwt3wPwB4u8BRwBuKu4H/6El+fmTo9zM9y
KnWJRY2azBtu55bVHosnB/FS2yqMEbr46S283vHE0pF9/E/qH4SwJuIrZM17Rmfv
kyBz9wZDsMxadaELEoIdJRHn33MmF5LaMlQcVyc4b9ACYk82SmsTQA0EXQHTTupk
VOf5sAXbS6ZFKXT7bH/cd2j/w+AwwhEDp0ZuXp0dQF/yQ59QERw04W4wmhxEzjNw
B7DmD26aKYJGf2bM/uVrWOlXTauZ6BZ/zTSQBHBUTWOKiZfjecl84Eq2h3rf4EEZ
pbdd1z4gvNXlS/QPIYWV2M8e+yJqfmRfeJQbtPLwe4X+NLL+2OLjRYZPmkTVFg2f
o0WGLDx3+YSM5FbEre6hrA/ZJ5l6/LDzxF2K2TQxCfUtvbzDfMshmqGgeXHgimGu
Yi7BUXgeD8bEpMLkkcKq+0rEDdo0v8IP/et3PMhRKXL9IArmGuTJuF4f+qYoeab1
bjojrmfVOE0Wqply7VhAG/BoOCUwadf45QAQ3ptJPufaEZT7767EG6BrNFTLYfsf
MaJ/HprEkrGM6TilVwRAxX5ABEuOFpzv4xRn6CFTktszB+OGRSL250yISXX7K9pZ
aakJh02+qm3NJgktM4qk9Cm+0GOe8RnluKoP/7ROIhWfHuVyHcxdPKIKqeMUYpoJ
OWq9Y3iYE28aBxUrRCY+BXFUpMfZXs6+kLVgy2szbmwesLYODTsduM/x1X6lncu5
0VXejEHpHG3GsijUHGTyjBfIvHw1Exy4aLhO8SdNh1je4VjVIoUuxlq8PEMcwLSJ
4L7dBLVLrtLKTQ4sgDL02YQ+FgpGs/Dq4kOhTntS64Ynt8fHSXXSzWzxur3kS8kx
u/RfztkuP/ixaSfTX4Wgpvl8F5x5t/U80/aK4fj0zBrb3rYMwzAW/vX8pwKVL5eO
6HnGffL2EBT2uKQ24WOu1DmKk7pePPfbI6g6dsxkYu0U6kCEOGdYO69jPJHz9n7Y
tzC2JdX5CWTfl2k43rwzMKdxcUI/yWIPVmrgx9DLOF7Cf1EKV20t1EI380aPbRJ4
BmpUrKVPeMG2jgOfegMfx7BiwuXEvL+bhIAmRyF2QIAovGOOB8qutJX079Pt63Q4
OfjwPG9Tr/i93mD68CeLMUqwLGMotdOePnmScIoV4OQrOH2O735/1kLBpfAvfSE4
bCxyGZ73/JU4jEFcZHG7dAFgUh74NXzxEg9tZ0BDaCC+7v2yLCqi17KA/xlNS/AZ
j/tDyZVKkZv2qF9E+f0KfXuMfSvow4Jp9k7r/tjVc3PVkIisUTdd0/RksrHxibLl
bZAJrcJcFufibfVUiS5Ys5KOCQWnWen6ADXqVV0pIGv2F4bXO6sNr4+XSOj9/92I
+zN82Kkb1uFQdrdR2tTDaFak86n6Ugx490M/gpQy60tvSQH5C4K1j1+cLu/R9slZ
sYeLZFvNL2/MOgA/ptgQxD2dBtSvOMUtGhnYkjefjY7IVKy+mloBoPb6tgJkm0sa
kZGoXcZnH85JhH1U1/ow08PT6D4hS/8PXDGLVK5qOXi1lXYPoChV/mYzgdilnP3u
thnEe3nEs0ijz34YcSlE/FvSELrZr9DD5FFKeE5ZPIE2yGoPil6m6BcWl5gxnWMZ
xoQIhlsOva9+lVO+Hsm5cUw1RBjzPoPcxuv3L5mCS/LubWq1erVKEBeFpNm2Vi3O
iQLaefdr674X/HgK+UV2vzQR/ngNyEPM2bIzQ+h1970gRfb92+NRAoQFvQW29qCa
c/5UNAqCLnsxibuNQnLaAVBPlUVO/y4h/QWvnFCjwPmta7LjptGFyLaVVbzFViCP
f4vbf6SmAi+aNwlqpQV7vWNN7qGhj6Sky8+IWH+dm7VGxTOx141fH9VU+JDuvVlh
sscqxidwlIS24OTRIozQXu3EutE11EAOWOtYKoQOGHC083nVnp3uBLreTrSsWUbG
fdmQr4QSARGNL58m2VhvMgvaTHIcLY2vXqBwW2XFbwUkKL9qjaXEY31TgWQkE/j1
tz0AuomSFc/UzPgkYVbt4MiGyNAxr5uvDxqCEjT9FTPekDckzuNtrTiJ3nXbh/Ue
r+b1W7/fX5rWY6yDgTsLHgebAyQywAJ3/524Q5J6cu2uOO7Zn6glrsYwIkiXugxe
8tXndvlrHiKW/QYIqJg80wKze25SleIzPPiCt/eBQQpaOcyMjbM7+RTuZLiqfGl3
s8GT/fvuK28+hjsWD28JVIKgvcwnVhlG8j4AssLHciV5r+aKTLDNcW4bTVkF+ivi
Yxi/Wn4VbHTHkIDepkWz3hb1hb4uDWB0FnZv1I5KawWv/9ZtVYQHCCbQ01AJ7S23
oTpezGNe7NpsDfrHKkiUYK/5EUcDrTEDhQb0YpQdKPWBptzCmSllFtPu4SqXOPzF
4d57RUvodBQsiaNjDyoHJa1oj35kwMWrbFd+1aMz2gPHvvFciLKVS+dcIiBuZEgW
2HsveQBX3D8nSdSaq/xyZA==
`protect END_PROTECTED
