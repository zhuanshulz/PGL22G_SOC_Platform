`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXMlMHVo8W2nSV+N7+bMAZyLk5CroAQzLWJLmx7I5cCtpQyEjBHer3ZnRXk7Ild+
ezGxK/K56nMB1ykGRbeEYZE6ymZDUP+pKGYNy1CA91ttHtnPF1EoQ7oNO65Hig2W
/k/mHHgrfEA8x4x66M1d6KO8bpGlFBZGRt1jMkMOtG1nD1tBhULkOIawO+9BM8h+
TgtcCeoB59rZ9JbpBDGjHiPJMfm5tW8LWN7kNSt2PY4p2Ihf7htZd/HeInND2H94
vxg9j2FkbxpWHpLX3FijK/s0BnZXrg/RY0ViJisAsVtsKa552LpQZ6qF+cHdIiJ+
WHAcYaqVboPQNjhBKzBbCi6a40Dax2Lb1uSiHb13rWVt1EBn8BKTyMxScipPo9M0
rGYiK7VU/ZJoMSm3ovdYvcMPNaZcbBoih9goL5/TsYPTmgrNPEqB5uxiVkTYdu7g
GuwQytS1RrVYo4ezOsZ3lnMIIR+cOpVQzFLwNpkSBFuECZDAXrQP4Zq+iyzy64Ec
vUjmM73zuzqT3su8SgWZxKPHb8UfmjolfkNvc5wI6RckeVnqNPAP/gKt8q34o11M
hGTP6gVz5aVR20Q033gPbN2DxN3Cp90r5kdDcENze5+tYYNbuepDMDMD+ZoYCNbB
ziPb9YPuz+uzo+2xUB9YC/qO9qvxaoI56OIx//62aoSAES3/nD3ATKPGwXSMo8c6
0eUhNH8jyGeZ8BiQuwzwe6QZVGw1QSI7yMU3cIvD8ULTh7FxAZctfmKErhpL8mJ3
M/46LoJvNiKXSmR5hVRqgomqyVW1S3g5Fn50zVZ2orxS8ZF4wqFKN2DoLZcKVG+5
1xw32SF3k1NVgoX4DUfCbIMAuQN9LW1+viCjyY39w8UyuQCRx8GkamU88fL/0Um1
8mF7ZfVu6Mt6xaQPKyvep9GdWxCdbl2aKie47oUJp+cWF9RnweXHHlumx3pkck4s
qMO2jV1/npKIJD4qLQ+QnDYQYB67rw7MZM1rwn6N+has56XB5/g7++2EE6IrvFd8
M3zCO4g4VYRlpPODggMsjku3sa+6rgo1a6FYMh6W77zXDtrvuW5uwZ2OuI431InU
CN92A2m658av93SBpdzIGZYLIx+WpHn+AGzKFkYOzqhiFdmXrG3I6H212jT1xTDq
Y89w8MeNn3xtHXo/T8+2w3rhkOOeeAHYyQZleQPC0Pk+O+tH/rqn7Bb0T7OhmfJ8
BikxKFN+6N3Fn+cZFnxlTrBB9x09BH8FtLCkHnQPwSh5boOJ/FwRHXbbM6lqLoJd
N7Se0vMWv4RA/T5rPOS6Hioc865Q7sbJaStyMUpAfXlNWAe4m4wKoQ7djK6AD9KM
wIpRFY7aeJYQz1fpbvtJI9dKOb9Z5R4ZqiX9HvHtrnwCGxCfwggsSFZk+IcegScR
duLSlOFKgZtoiBq4wuW6CQBrcf8ybfigTQvAqw7znscFsXR/hV4jDi2SgXZtRSvv
f990/rykwiPd4wfJmElSMZ0nHZ1xBBjX83IqQ77BfMVkiVKI7gf20spkalgCFijH
xiaRGcfXrAZvtrzie4kcxmhSLNjNiYocBwEomMCaWUuSWxP8la+yqSOZ9Fg26kuU
OqnN5U/Q7XNWsbixcrun0jDwLwB4vLziC/gVCeE9sBriOnionD1zU7ct89I5416i
oDecy4Vkd3Rx65Zo7v3a3SrOdDJmCxrPlo1t6iUopNFFkvgsfQ6HtN0SP3lyXipn
oweEiJujJ7McGlDswuI0nkDYyJQtJzwMsZygBpE1WkHVVWerj6yoEeKvzM0VWGSO
qLWd1EzP4HrbfA8Bwx2LQHxz8gLNb2LGjwIxOqWV2NFM9E69h4mHTd4hwKlPREBu
YBPegVwqPuJdj6h2kcplUP7pHA3yE5lHtQqu3GbRrwzhLaFSXWhmZOKc5Dk/gYFp
01Zrl54o8+CIuH5GSsctBRaodHYnnOACzbM5y+o/pgR1zr7eSbI5Q99OmyyH62R8
N2qBjVvLAXpzdsuyndrI6l6OfOQD+lZKyzq6+vVyn3Kc+FBR5bWObve3tjD7eqjF
dzIY0g5bH3fTyaEbVC6M+uuIi+KfzLJAZzaozEyY6e90wiLJGoHxDXeyAQrsOy/F
UVjq3Qumy5EMhfeetcYkeI2QxxzP7eqBNPzjHCaoMAbb3jQ76yo4cugSHte1utTJ
CfbmkfZlYtnhBEc4hcutQAOYG+RSXLaufCYbaWbU7pq2gUY4KKbr+WWpknGzE5yh
5p41G4LpArJ74imjPkR9fP0sEq6I9VngDONg/a7tCTweVDKGarN5EKBFwNfABZ/u
CegwTHL8/HvQzwziEZFHFAXSu2szzxeduMh72gmlFT/gI4yuCA3L2SWIhOGSxSjf
faRogomwa4igEuEQl4aTnOwx1IhN4vjqkQCnkiorkiyIuHpkAfho20iFpBjJTnea
FKyD1XJ4J6m2P1QKnIGECUbEM4vgUrFuAhRflKOPKnuM3xSuke65XKh5dcfkYoDV
mljXggZDxDdeMN0o4yAwGsYUljmjCg+AdRhSd9hjLhV2jtJcVR5QLXdxcJWGhGNa
5x5L13mrVPOpq5YbieLKR7iNfnF4nP/2OEygrERc0Oq7LlzcQ+mVC0QN86T2YcJW
cA5u80KZK7+qs++S4Zk+6rUJqbfq48OZ26Erphs3rYOloscPRd0N//CaFbNKtvWt
hCNuuLgUok2zqpjQV7oiqiSiq6Zg33VtUci4Bournm8p7fy9epjwYQftwT76Ac1k
VoG2rBcSavDJwC2QA3eV8eOhXzGdsj4kP6wAsqrdSvbOQW8n6GRkmpmi93Kyaa9w
mHIM5j+AG9uuRnydBVtj9FKEhQb+Dnr2uLIyHAk65iOWbVGb7CRQGADrJBa9gXgM
8jSqD+u97bUhnE/DJtGkbeLvkGGWdOA8r+K9WoDBz4mDgzGKqnU1V7Gyvp/xA2bx
u70ZDkolaMvek3kfAdXlrgivWb2IyuzGeWwtWWzmk0D0pwLXz4TYerraYhIn+SBW
KTC3ylKEJ5LeQGtH74sd50+G13oblnT5/FAngmVL1FAHl+OuF/MutaZnMkR+/awa
8Zd0BC9fAdDHHgdBk3kAIN4juyxhce4//AL9P7OSqyvB+aWVPu592fZ797B9inms
fCYLDK0U/4a3S6LuXhuHiBg+O1KpVeDIyUC/tDsvHGxI7KEd3P1LwimFqbn57XLH
E7b/3HuH+AnJ82Lpkgf2q50x3vrFsOG6shWKajDjDtGXB3uNcIdvAwLrw8zdNT8C
ehOmu46utcE4557Xr7xEizfRc9KshrLY/RYhbbElAPrttBbDfBW4+0eGHfu/S40Z
Og3vrbyGYzEfHeGv0DjBPK0zMyyjQ7tVsOa7Be9LPmueLgZnJTQg0nVLLSCiSWS0
AIzWmVPf6SydsuslGk9d/6nf8flXSxplLCPAMXcUfTeAmS/1sGaHVxuTINev4muS
yC/JaI93eQ/ynsta43S3DMNvYcNhc/sdI7ehS8wfzrNOnej5zNQjiyYVNUhxfIC4
wIvVaB2YSbN1ptuDBkfVxkfce77GZM+vZYxhBiaSzcsF5Z5UVOJXkGD0xhgQLDiX
wnW4AmZurT3TsWt72A8e9U0cV6OKleGvWTIIjX3NTWwGh2oshBA/AzNLi9aZtgCT
yQpwtveta05rviH7+zMv3/igDftLYxKfqux19YZzYroApwY0WakJM87dx0+jOewW
H2Vehg1tch5gjo31oU6Hflc2O1qRpIwHb2cKV4OJ2kKWLcIPDPUA4GT42fvRIq6I
r+cSfqzUKRdk7XEMhiIVWxKEdCJsXCZnsWCPpaXqz1nD5ph00OlCZ5DAUWNbM5d3
HGJwLjh5gaQCVDm6qh8G83OpcVpQW2A9PuOALpxjoAFs4obp8PjvLj29p4mxmMEF
9SY/+V03jWRVhrAsbIhmGMf/4mhFAgIM/Pqkgd/moF08hwKpK4bOl2LEeT5lzTNy
UynmguFucWLU6BPqw5Xk92nmFiS+8ahz1ZWJbZ/g1LD89Z0u0H/TsGuZ9UIDPnxN
t4OAtZKygRr6vOHrjuK56+0mqElHRhRPVNzIh0ERl5BYjAC1pM/qyricscXH6EiH
X0xK0FBJjxvdkZSedbcM4bLhdH2CNgBObVjkxcXCJP83HnN37A5nV5RP6vRE06F7
kpTXkQdzZP5zGR2zBHp2YPoyJYkoE3LNqe1uwKBr4G527p6lptDWc8CIJysqgFUe
9Z2uH0dJKIGhym3FRjdUGl1xg+f1bVpLT5TL9SGQjonN4GpOxcueU1ewDRFICsTi
Qku8IpF418LIvhkHp4Dx1giyaDleH/myjynDnWOBtEPZGYMaBHRGHgxyaJJCREUz
Vsd1SlwSZ1MG7R5l24IbxWQPglhSSQ8oImM0/Mlg5MCj8BnTVU44rXLg7cNIOCXv
C1PBEYEbscCbsGwyFSUQopEs6Jp4joCrFDADNP54i8aieu/d2rk1fSxdG9zBPXal
OZqOZm0xjdn7qO6WAh8wYpd4Bm4he6BF/rh6JnQKmIA=
`protect END_PROTECTED
