`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dmWMSrTePa/hM3lRmuvR+9KZG9/eFCRXsRvOMXIWBLpvTvJIhVjosnPWiHpDY7g7
hu+moSzizFTrlO4dVWRkpN2bCw7qgx2j9ysGMePXz/xyVvbyc68EIvbt0viAdMyN
L1+c2OH7HFwJbvivHDJXg4M2oZIXed/VGrdodULTv6/RnCsFHjbE1Fr3xstoh1Ir
g+b3u+opJp8D3vbNkVloue0+RKj3SoEckRYqTDlaHIzh5ZssNOD9KVNhSz1c5ikG
QZWrnlZ7v2kenliB1+3UoudrLK9cm2fTnkynX+3Ytqrdm5kMConTyJVPq2fHQ1vH
LJNjKutRHTjGdA/mOnsU3IW5Djg5nTGmWZl6d8zqclCTBT3bGK2ChCbgmdOQo79W
8cp4iWZIrMyD8s3E7ufDi/kAmLxhM8n+69Ds+Onfo9zINiJo9Y9X4JhqnLuKjE0o
6DlksVmN9ZzNeA75ZdBPZALmz4gCIDSwar5NICz9+Vc=
`protect END_PROTECTED
