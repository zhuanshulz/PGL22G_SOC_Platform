`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V2OUR6OYAHwgscsXU6IKhsjJ0jEtluGySSSra41v3ITMdlCPuI9ccJ5Z3grV2qyy
tLPAX9brdJOfJS9ZHmBlyui8y2EoV1y/19O5GZXtgWJyl5oB81uMVHKh596+EmzW
VCEK+OTM8+MncxGDcvc1IDrq515DnlsQ950TfVOGTlp75iXx4jDByQYddPxL5kaZ
1kjH4TyrKpgtSYPB4h4PBN7OPgJvLm/LxCcKUKt+fmDO6NxBoXzcpQsPjHOLPkpW
aPEpz7tKLxmpHte00YTS3qjBjoZfq2GZD0Q/ery3TGGxSuNz3dZNBvLhR+fZPfcv
2Lxe4BG8q+a9zJZ0NtLKn5S0ogj/4xQlM5NCJY781FBKn9SrKPfi3VzK5DBOyuBA
wUUXXcQGf0yXvP3uYQ12beSLV01ULQ7MXAHkwXuSf9AeX/EV9kX7Pvy6pfURc0jM
X1n7oB3bklcgIneIlvgOI6GbPBycawss0rGW42GW1GvliMljkWxYWI3CWMA/zZCm
uZ152KA3XuT7fG3gUNvBfNQVKJ8+30sVrrQPXCmC8y3/aAqzmACmR0X14ib0VpGy
zRQTD2AyYfLMD+f5mEnEgQ92geyk+fWqjm3Ngo748wSSiGjcbJW7ZKsiVgIBlJ5E
JOYDH8daswXghpN2mIuGRxSvMXjJ/FU8jz+GwHrGRUPq/OOQZ4TcOoPXaNfaIjq0
elYAjftNz9TXfaOdgxuw4saXnsa41e97lELrIr2nKkbpAfxa/0IoRsOWxPCURwQ9
SbvpWMywByjeV1aN3g8Gvv3KyzhKPIiR9LoLV4fdg0cxfSR9fVQk4CdzekgtwNBH
XfyGBdAFTwXj9QhOp96w0z2GM2P325F9Cax538jvR6lMxfIuJqqRs0bFyy/4kNAu
nUVajm3PPRe6Sjqqp0BikUmfI40ARGcXxN6nAdjg88uhSorrh+b+0D6Z1tywRlbh
+0M+fsMcrMOPjZOD6nKBrzVphC3WM+dByKkSkyWMzDoyVm43IRlxiPW/nWZDAhxI
UmEEK3L9+BbhR2p5DXK8YoIcbVUlWiVr3IkqFlKKnbBrzit7EDGzydjqrYq/i6M9
iyCH9OmEVUcf4jzrgFIJ808rxpM3ZYFYhqG9uBpXyi3ekm6FVlRsTM9DV9opXsAI
PPf8j8mCj7xo6LuOInK36aruDUgGWAoJ+Nh7OppbJ7ptj53FGUcS3EtxtFBy6QEi
hdHoUZf55+sGn5Q4kXLNviEVyJdsEb4J+ivhuB8G5W1QgXjrN9TaU1sB+MfMHqGZ
fUFo+AOMB9lwhFIjwNOs9l0dS0Th4Jhk18h1aErHcF8Wz97vkoZ436Evr6GtUHQz
7Jq3LbBqNCURD4T0PK00vtkbmjv2IKrCTl9bhE0iu/fkjqwGxJA3rldOXF4yvwhj
wOGXuIQMKO6RVSlRPgUNMnkf+i7EbPrprglZcD0I8SHf2AJa0n8VAfLMMMaWydbs
8YKpzJgtL5KjJt6CdQejnAtmhJCSmSmncQf/5g7NiyjgGjBP5AlS80alUeMQPpaa
r9gZdymUiHPvExCyDOPb95yTL0iVQRW61EwdwOrh8+MJUKTZV1xjFIh2IXxTTaF6
lhM+Oyan54GF6q58xGUHuC+Ti8ZOq3KxQjhJ8ai03flqsiocMBMOncgdHg3KUo9E
p3YsBf3m5FMPK5w6+Od089faBwjmfuOgi7zsrXUS4mU9gm6mcV/vOvXV1kDp4sMt
GjCx/HkmDfKznPI02ePszMEiglP+2GhecpSHg5seilFgfhJJtKLMSIXG/ldT5sEJ
B6g3YZ+LKMVjkiVc8bHn1sy8JRYOwBH0PZuTh/Md+PTxLaaMt+XgcmgdszD7fktt
UoHrt0H4GytnbDoMNzTqeuazDCFk8pxAhI857unAjjPq5pN0Ajf7ufH934PSpGdM
DQGNHjJG6dPLPv91XcFuVRMLDh3Ao11uU/tqQzPZwsZ9PCsZz8DKt4OcgmGTfBqv
2SC1fjP9taNNWItYJxY1u9OdY2hC4ROFnH03qDzuiKH7xHDFWbfbwb2RsaB1jVR4
k4jswh88FmdbwIufOKiY9u8fgJp8mkOB0rChNjDXICjQmzlgpAaUBFdUbXYGi4PR
9Nefed/aKEjMHPXoKpTFyfh4MmgBz4ZrJ9Za8lrkoYe51HSp0dDfhzeBsPTPduSn
OitK7Wsdr+DUGaao1B0yRTYULPGQd4/3pwEAPmbx+xoHTvnGVuj7hyg4xQNB+mFF
NzvJ5FxffUPMrEaoVAjMXTU1FTddOWEuuao1zx2Gw/jMgdSQCTF3GPuhVXQMBOC4
qk3eZzpcVaj9e/qgfEzw+SszYv4pwxKGK7R7naWSDQmERwZyPBpNkcLUwXq/GLls
bE68Yk4QeV3HA3X/KpqqIngynnEk1R8U7PmQqKhKkHKyB0ih2c1twps8ukQcN5l5
ImwMWimhjRaJGPVKynDZz/XZdgLYRIt3hR2gkdzcZrAxbLJIHcbEpQR9z0h2MCoV
zQr5bUceMULCYRKbS8WWixbYSRhtHy7hAnpOht1Jll53buvxVAOeg4yBgifGyyE4
ke/Q4RfyTOoXF05s2eFH3jHd7HlQu2VVztWWRiqkgYwYvMcao+14pmMlIQ7pnJdu
6pvn0xCx8NtUzNMM9Adtboju1B6gYYDB+zLC7O0pNZjy8Z/4E+NOnWJe+KLAE7Td
DXP+6Xd2UDODt5T9rrp3f1boxlcfHGOjIWMXqrVO9tauQdiNT6L4ddJxiq7GF07P
PUOK/+PtY0AtDHpb3prqV3SUkbg4y+xSQfHkMIIClpDLQoOucVQjIAjEuHqGEn5/
FWQtCNO+J38F9XEzgTye8cWxYLERz8iFyOjzDRdCIRzXObtlOMiDflRBTI0qcaIs
63vp0xdOmGVBY90Jx90beE0KnW6hjBRHMBYPX6svgFsNwfRnNMblX8dYo6YY4UGI
z3SdnZbcwk37ptpEFyM6iXe3Tkw2rOTYC7bPUNUqL3dVAbt+N9v+N/9agON9UkFI
ed+ObBZW7ZOYbCkEPScTBYMsiJtP2EagcBcPuwdZ2g5dXoTG9DhXRcMja5TAxPM8
IxJk4qxjaWsAMxTGLq0/L0DuUSmJHWKORBFtEXJRTYOvxe/Uii5w712dvDCSR0RQ
oLjeOOIr9jZayvkPl2P5mKm+B0eSxDro7TCu+CAvEDhPgHfna4Gxuu5+YOmnJeng
/+dwhQUTi50Ostg8ZQ2aMtVnO2vmdp7ki65JS4RfAYhUyCgalBpaox/TI4eWaNYS
dMqxwtHVIZyaVS+ZhcT9MaHaNwBNxJmDc2eNXG7clQ4I8rfgSjFpGror4VXOYQ2D
aYUr3ETVzUOD1mKZMdZBkObcmX9Gnk8u/VoB3DJdiOFfD0t179xa1LO1NJvjHJeL
7cKhPt0ZB3vU8zdZwx07wc6TtjJYvq0b5xnmv/Q+D3Y6Y8OzUPyrH081U7LmqSB5
tcojgQUiAgmyCeDzH35xf+ydu+tudCk86aQU2aGPiRk1DyaYnl5BbcmOkRJMnmOX
UOOC4MnslR67uvXb1LRDxLoNcCdbyL+Qt4Jcqa3nhuloXkEkcZJiNcROlvoIjv0G
sjtpGZZ8mD6ZZj2FHM/oDm7JHBPpxJMRQPH+wbHlDDGITV2C3zoH3uesAGoPBXTo
ZNrWh10lZnGN7sTA4SiuFT+5Lv4jbRbadSB/o+2zFtZKflbF7N/xtVvVrXYG14Wy
n/RE45706I50zjbFwh/kNUAVPE5tvCACVUBREi07qAiMkLi8cqrAv1fKAZnHCza1
VgD3jXDZzV1RFlvuapR822DKY8jg5ODVkrnQ9vdyh4SD9JwllWTch4cO9K3jKCmM
yTB41akecoJbhSZUrxypp+ZRwdQrXlRA16kEye9Ow6rAAjjONJCWoikRnqx17v+3
MGUEG0V9iIuEEj7l0sutg+AVJj/iwZ/wGFRifUND4T2+23yLzfz8qsRGj1AuPKJU
U4o9NySb6CXXGeQxU7uqn1QONk+RiWcUJmq5IxkEpmG5bS6b5hYrqYKiHQYI0f5E
OpL1D60ow9w7pE9RZ+RqA+FTBiqDoukM3MO0APdhe9/BueSJByd6Mb/XspWeMv4e
5F1FGP++q4X5g7aJ3jewmhR/OKbsyl4cWOZwllzfZ5zBCHEnWbO2Ava0fF9KN9oC
tNfx2T4Vo4gr8FNItNFCQVp7aYxrCNWcUz8oB/vajaXvEr/EbX68PKdJod/SLygY
oYArctib+m0Fr6uX1z4HzA+9qdG2lm2iksCuDHngBPrcs+YUF8C5wAIRWFaIWJs5
wtDStm0IKh+9iPLvoajMjY1rzSGm4MdcYySxGKiLzTnYyZFbVtzxLmVbevU1ZnIM
aNGfEQ5cfmPqR6tv7Pu2kML46ZMgBdwW6guKIWRKiSZqGjH5YrCJuqg4w/dE48g6
ciDXQUGsQiLOGCjilBjjwwCDTJerpQOU+I+hbGp8R2Hd/3o6zJiDEN2g/uv5WRp5
WaMSXhzDQG4EcWZ6wBoU2WeimMDbQOz9YFogcdffsZX1d7tL2myfc08z3KnFXsx1
oHSKONJNBKLlrx4LOUMJLdBsGTRzayCZRPazhfV0KVB2ocYI5u6i261osgQqcMM1
DJVKh9cznQQbKYjcrmso255d5py+0NmXdQqxOuBw5GTak7+7RCe4ty9gKWM5wkN9
QEG/DIBPYkgFgMZrznlF8BjSAJ2qSo9eSXxlny51ybB7UHVQVGDTyoDVABBwzMmv
cYW8KzpohsWRHEPdyBifvxdQ0BGQeNN1akoiplZy6uNCDmhAy9y1oqe3F6ZI+8dl
NWmPpgBW9a9ZyPs58mStAOIRUPd0SRN0pdtTP4ySfSfXNBnnE0CvCMtH5Oj4K1GB
x6ukMoJHTEuLnZYS1D0KrXa4gF+iXDTvPUbie6899kYKhPQxyJ9No6nkDyxCBY72
+0dQPJVpXZPYS2hmOW/GnspMYDm9AWa6GgpXWnQ+DLJNqE3ccR6W+PSCdRphZyuZ
`protect END_PROTECTED
