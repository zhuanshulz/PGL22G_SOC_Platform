`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6/vLJBJkkL+/tgtyxdEdQTrtXAj4vU5OjBUBxW1Nd7vI0KJTE7cHnNdEvAIbLcO9
jnRibovZC2IHApgEpYduuVggZcg8wHx3V6Ud0gFVYSzzKdZEGOqOFvQYrOB8E1Dp
nZc+KaG/dJU82HqWYity9wJ1tcblDoH922mDDmF51+PKXJjnFkebZ55Z98qWNwW7
i1eAPNaT1+18Zllg1vMpO5eWjB9ox9e8CTSL2IrtE7sHqon0Ipvm50uNpvTu/ij2
YHN0wTYqo1rnB48d818KWvFa1xXzLEpWrYhP+EK1SXhKR2nYEgwmFei+zCLUFEHS
Zu3Xp3iemgcdIvWBVDzfFnhjU+v5dKhmf8/u6ziB9e/Net841N3p4R98vFO5VoBk
5q1U0FIWQKOL7YFKIcztMnjs8YEWth5dltuPpZcGulIyDjW2uFqZyB8SlyisYJEl
zf//fpyoCio+nrdH8Wl99jAoeSZf+6WQCCw7wJejBJ3feHLFsj56RELRJZNLoNNg
7n2DCbwt75Qz/E28+T3NZQ==
`protect END_PROTECTED
