`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
740lFQmpe+QriBDEDVoW7aUWWUYYn5wQ+tafU1CUlp3T6IEqyPPmpYGdvsaZISJ2
5JuOJxxSLjT8LOD0Nblwyej483h7M2cT1sXXs/lR4O7JN0op4EiRNQYI1sx3qCdF
3J6tJzHUUEqX7wn6+KpZWypUcKGyfT2U4t0Qa754qeQOilnr/aYOeOl7bK8TmPY1
HfMMu7Nc5Jl2m1Qlj71wakTsriwf0DVths4zaC966X7AKO58sdiV/bjbu5vnpL8X
gODu7KLB8jiwo+Z/ngIh9N8AuHPPNknPzGhyQQga8nf7k8FHwJIZl3NS2G+oHpH5
zXNxhtmrRMh+mxbo0oGzTXH3syGw2RY5NOGQEEmXM8LAnWjNAAXLzB+HwYO15zTm
x2/lOx7FjGFSFqAsu1ZuoQm8I8GcspLjXEnHtiFNZw+AtJ/jniGaU8Z8n/N0+AKI
krPtVOBXjRGeNne5k+XwPpSP35S4+sExaxaurZdJkJ30LsLWdDQQ1TVmZDghSpok
J7Ey4oj8qnRjnKm8gsxvaGmnCzTyvNfPw4jTVPqn7QIRx3w8oSQ/AIns2Cq2+zxs
hmp2wsHsljC+nQUHGjDaEDrTzAMIiotZ829zKBU9UHGN3wG3xkGgICb7bGScXuuk
GJNMX8CFoLCvyONU6msPQkUFiZJxaFumTc2gPJ3HS401kCf9G1Mbmoyi2jlaDhhL
3nv6K1rzYjErQmyoA8H4hq8H7YvmDV5ZZZ01VM5BTCNJmnd/DTpJ6WpeiW8q81Hx
sfpQF5hKMgi3JauqFH3zgjTbwNLrBxCvktuzpwuHIIzcZvYaXj9nGsjORQet8rqh
/WBaPDnAwrFvHlaO0hodYV+UEseCm4/Dnhwgok/k1mrzcLb8EIAsLwdDjQuARL+8
CTjSCh6C7Y/kiCZ3cR6Ir1yUK7INelH4t9nbhTht8v4NuGrMt2ZyJC0RRjsBE+JO
VizdCCVRatFaUUrSuP3SE1XbRrAHf40WDVfOcp0rMrxVihS0keNhgwIoqqwX6PcL
4scYBp+CC0P9r0/gxlodg9T7DxWjBrgdHAUSYlHtePvHmu8plCK2QFO9qV1Q46ge
5u+/K3FZyofOaPG1G2dI69vJaTZOaNWXAbiFLEHhJ1+T5jF/Zhi/LMyERmROJuyG
MTSBdc+TbV+74emwJP4UJyL4SHhBm9/uPwC9dCN/qoeDieKQxv29GXeHHUWn3C3x
qJ88h3klIRi3ESP6Yh0IKWxqPFUGeiOLV1m/hy8U4Eojgg+uHn/0rwhEL4s7UD61
MugDDoJiJ0rxhRanH4nhos6u4E+ba5RilmXOWEFvQCpINNxSvU2NiAxmXr7ghxVe
JMWhLpBoqtFUyAD6E8L50I6mhbnCHmL65Xyt288vb7e5O0ddfYDCf/Yzr+gXNaHo
ikq9lxiLw4ouVLoK2MnXX2RpMeUFo1eNKEG2PFfzEAEoGDn0yguvCdXmv0z85mBs
LOCahvqv9Q4abRpcT6aNmqI/AGRiRKGpfq6Anit4E2N9vAf9hwrwB3yrs9s37WSn
iidqD/xXh5+DECiloqFQo9QKs+CG3X5nfMRNyVjEnnkreKm9NF6m/Gypf6Z4epjh
ltX+YLiy1ykZOA7akmSGqV5GYEdT9QydEJJ45u1PWncuGYGwJKcCXlBsA7YquLOn
XLou5dKFMDEkE+UEgkyg8kcDB6S/XMPyiHVdBYpzsyDXqsdEByZ8RtWTFRrdi3So
5zLN8BVQiLg7sCZuBRlkG3Pfw0tkzlv423pFdGHXFHYuERIXf52fv/D9naTjwJIf
nAITnHhtGHXEY2JmLuBynqbxglYZVIMOoS/W5GwiZpbHrt7grSp3ZXr+hhN1gd30
MSjfTGLLVTxSJF1U7o6o/+RyOgkZiovnSWTuKSFM6D8NnszUAcP3OSbg393zTr8q
TnNlNyG1sy171OKMb45gEpaYs2ARwlJyOIAwjf0gkgArgHu32TfPtxx+Pf5s9B93
PTU+SN9vi3ehCYEvRP1xiUGvKm5CAOgBVr/z2VxLdw/wVIm8spwZSfwd0V38n7u8
35zSVve37wnyqeWsFLWo349vEfsGwPZXzujwVxGswGPuQE2BQREqjWmjcpQzHYWF
CiXjRzMOLANjMCwETLL8cTWTxb0oRyfVd8RLuL7gZifLBrg0vIgGscXbZT4RF2nd
M3plQZs0RbOU0o+SjA8EJnBrMwA+K2KNCJdQ2CwcXuJU+VO2W9BQ93dUNmrGdqAx
Q8p0+oZQiyjZeSd+GSgeORLoTOzy9xc3jzzH+vyT+mmiv9+A+qsJbQbUYTF4jRLy
XI4Ynt8cYhVT9pomD3LAOw6m9O7awhMIDa4RMKKRmNX1PPUOg4sQR/CdYL0Z91B5
UP96sA3kiqxiU6R/pqifpagIUdpSMXg3/sBHJ041E1EK+l+NgSJa+MahfEr4tArQ
q6TfUMIsaFljtGpZDjXMAADOTHnKHJSvShXG74qYRiSl79CZ8NLjALSpSVnBGeBD
zOQd9l1SCpICRl7LYQFzedSW6fgGNwWFJfV1y8ZRXTR3Tawq6MxqXIhlEFjGAlDq
bXeWlUNVt32cQf7z4auwUSF/UxdkMNWqfESpwQ6I5p7Z+YC/bw1ZL7lH7SNpK17i
rMyjCX4AtAiAILFEatdTiLuX39eap8CuD9UbL3akbtr1IuXolYvxGetjquEvA6sI
Pf+DHBaVQdSpllUdYS0dEdV7BrohTmO10AxQtIbd2VcOdSln0igByximx+ZZOq3k
WofT4s0QPxOs9X2CGdSq8foOtSuMbTAG0SiM/vA0S9hxzJPDLxu4qKm9EZ0Spdrf
2EX58larA0o/Y/IYcnHP0TuaLT/6D9SIgGTSi8q829dwIh/00CR7YDl9VwxkykAy
QIqwyC/PiBAjXT504xbHc+Cb8RNjsAAWB08c93FGQg8=
`protect END_PROTECTED
