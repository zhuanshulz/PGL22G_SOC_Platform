`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GO3ntlQgrH2/pRdU7exYbi7EmC6DRbkTIJVMB0pKS9yLZVHX3CIsGfmgOdd4cs2J
5ekqhHBc3KGWsFGv0DHJVdoxljG4jJ/BQ452KrVYXOwbehrHDkMKsHg31/K8YXVO
yjOfg2pSuSAmaDrHzcLAxftmtKDv85y+z260hknqAIzH7mTQ1XSWzd5HVbu81+Mw
AlPJtJT0rZ2hmKcsvobM+y87g8fOEgMeWdCJKPL1d/VwETNs3Nq42yKFK6be4FPk
oIK537w2S59KTuTS0SGDiUL0aOkjsfxexFGWFyct2WeuaX1traSYOGF/YcRw1jID
LKwDEcz7H1Zh0EZt8R7F2sIikaTafLldJrMlyqLp9ZFTy3jAz1/SjBMu3Qtw36tY
6bG6/0X2uRuYpJrge7TdceRsrVCytG8+D9QAnM1lv9taAv9YiE/yTnBZHtfZ2AJT
Gx8ciGggp1ULYpGRf0Fdil7Vt+M+8AUeXXHmk3a9Zlr7YyKGYlr0p0Vugibj+hz7
lhjceoaI/YGS16N2WQ+XGu0p1itRNaUYvK4W9uu4MHJ1YV/a36rrIFVO/mz6k9y/
fKiZDxWZ61Y6P3ztWnjPlqJYjK5WqmiADHPHvHGKFRT7gX0ZsTpjfTnsue74fWJf
eIG3zdrtZ5Z5iQ4XgOdg/33AG0rjP6CBvbdfsVIOY0oRlcb0fweXEmpakU03uDuV
lxVNjFJ288TpP0q8GQvluUeA5FYAX2BJhZuIAGvhGKhkujiGpzK9BK2lA1bZtw/D
zclctb2HazJl9e2u/8JWAukYOSwz2pYiHVq+hzCT6gkdsBYOEWyIWNDhOhct7yKw
+5UtT3oFwPlgumvzmnfYE7+nYvPoD585kC876x+8bwQMHny+H11+FKnWrGvT19R1
iz7l9EX8hrU3rE2KbDItWr9vZcnFd8Je4OC07yMn4rVbc0hMFfHgHNGaGvZIotoQ
GS+W8ywppBXoBONuZjPKNsWrv6e+x5/9INCKEqmwEtzhQBbnA0vBCvZ8x9KlkAcS
KoCUnEj31BCbfVBAposGKp6mCGA4qMWnzzefFqWns6N8AT52TppPbUrhlK6ruc23
WsENhdS1bYPyhN/iLh2ODPOhBw2z+YGt0KEwm2zNHTRSce7MwSgpZoZWW8UqlKmu
dCPrhasp9AbGeBFiDEkwxl6hvdOweDjS8oCwIpRLK0AY9foxqltJBuloBKkOuLLi
aft7HdJ+eZPeXXWb2uYjM100/imSW40rS/tmd2tGltSin3unwVjZR21+AHn8u4cM
PHldkiLSwPqYSAGjsF6JW2Do37RTedllBwtfNudFzVORt2F61/lz4EdUPtwe0B6v
MKLjjdEU/IQ1BO8TZqFzWSm/EsicnCeRpqkjurWkDlKTRtCYAOxn7C7w7CRXf/Xg
SsHDJf1MQqY9I8+sYPlOA9LPdsdJc0J+FrOi6jf8gSF7fcqX0AOJ6LLa/MnpzrH5
xww9PAL9FRLuqTxq8cpqk6AaoSSJ8OBx3deU9gUZ8Q6FfNmsYJAdxThP21cAsp2O
qaZVkOKgQw9pvWyX8JPGvnp8l+QlyhS4OiLk23eoW+F7s91iVX3G+EqWAMnEL3JL
jRtmh2C1odE6FRb2a4KcCpEEskf48Qp6KvvR7MDMKHcI4v8R27Cc1um7txt28q4m
JFIjsoU7A3cGpdMXtsQi70YA862IB7npJ9MIa773lKSeOD0h3vKaFU8IVM90yJKn
vKBZDXrCl/oZ0X3iCxPMDNDKJCqqj1KBqpX5GY1N05J+M3clahwj8gmjxQxXSNoa
WOvvl8h8neA3Caga4kT75l+A79Ppz2OzIGlXEFCLvYUAheby0UUacpFRr6kh7b5x
R1RPN2vQ5ZfOZ/OK9J8jFpjrJ/GcWO7lTtqCx7vP/IoPy1veGzJh3iQzFGmrAAhP
hu7ZcZnCPxU11X28de6oFWP/WYbQ2Gq6gTWvylBPfqYtSMwG8W4gVjstOsxQwvRs
REN71GKTRPEvw6dI0WggDMUv7fbDzRqvAMO11fNHdDWFT9PGr0gwP7sU0NaRcKf/
wSTJguGqy5iJscakA8wSrEWX8gxCqtSH11prexqdB7pPWWh6AfjOANCh+KIIrxq3
dq71uwxGWkIlvDZIuabTk4H8PMInaYtgsALZea6catZpptluMPGLmIy9TjZQuyUK
lPB/p5BSfmafRSAazimAWJz3hHcuGShKTE5QJQla3dgdoWsPQAy5H/LxsaqLtZOk
9gPZysXWdsTcFfVp/R3brbocOIA0f3OZdPXyatx/uU7EG79Fm19L9M+IPFUVhLFK
bdU24dMys9XWb6qWwd/6+vyzl+cF2/54/QGVkCDGlGCQ6wl6HtVs3hKhNGrzw6sI
4rsCNZGjYP7ElFlNogE6469JHVlsL4CREBp4yyBkvx5dBrlZmJ049jE3ZskJq3f0
N/dFNqHjmPvtGY/On2rvxJvstyrHI7si0zB1gF+eWRAhyxZtJwsX0zO2rsIaIJKk
c2srM8+uIMtnSMwLvW8WCeUc8IrND3P4RqSmcVqpynNIEic7qqFGp2BsGPKlOsNd
forh8WWgxIYni2R53wJ9Mw7lwYEtg46aFckRZ6XI2reEdadS6iMVfMytednynBF/
6qYbwoSYwxtZV0AnaLieiev7DgFFI3i/TYILCus0Vd5Gs9NawFcLorq/0//2Byf2
Bs7MegW615wu3G6rrLfGdwKYaxarqeOVy5qr4GaTkqeVEU1g5+SCw2pDIc+yOec7
fnikP6Ld+IR8dW9colfWoQCYCkPePp3z/Qq0hDXhBLDlajb3wswLtKisDtOVpSiC
mMQtHG0Gmo7MBwg5duS9WlrImtNBIh4K/UZKiMrV50m7z8uMXIlRssnsVuzp/XsR
mUC5+wtEqThF/q7bkDzehs/5mAgZU/OsFz/tyAnIHWuIDHj9i40M3ppZQwU4Ix9j
1/wNrW4Y/l8hhERAfhKtkhC+HvFPHcCglXPgOB3eW1msgfC9Qpx8bcH3l9iLrVDT
nBG/Pyl6JDEy8X6JRlmwBLL+L+Vd6v8Fg7Gdf6zb18twLgrAZdEb/zUMRSl78KEi
NV5sUdob8I0axGsA1aV28eI0W9+eBQHsRdrmVSwDl6xW9UM2aW5mGq6UqW8jhOxP
xQ4WAjFj4koD5vh6Tof+EsBfuNcI8MLYBxwGdtvs82UmFrySF/UtOVpkfRiDv8LO
omA1C6I8KkXiEKWt/C4qj2kyEAyNOfbShOKoCUNsc45PzPa00a5yB03n7j0t8aaq
WwG4DZOSIZaqVtyc/b+EFUSi0m4/UlXdtJxg+V9I/BKRpxMuioV6JmydWMpTowes
Gz4ySD3GFZDn86cB1DrsEOmvbSAaf657Vvb2ihnGG7aJmIQFzPHdKCK+jccZ5xZr
sw/KWuzfvZnapN5XiQjHWBdg7cCuXvXx1PFNaQyHKRd0Zc/TWaDMe6LgJdLcm8hO
0/pLwGb9ieDM08t1H2svwBqc1X6ZZ2cNKkquMGnOuaLnaxOJgRaCJrTyuSHJQfjx
x8DHeK9Dqvxri0+pfh8UdYCWByXQYbwrg7ImCihiFt0gEFL1RUVVZVVaxlQH6cSY
sy88EnnVog89ypM1e5sAKKp5IJNOM5O/oaaxt14vwDStrF7WV9dR/K4bfiKQf8bx
1Oq4h4vExm5XyEqyIAZosAquj6ucNEpE2S6iLZbZq3Cv6KTm5AfnN6n9yRDV0/2s
LDk/I3J4DIZ7KzFgA3jzovlLzqp1hYYpKK3L2VyaCLHZ95960Q/gM6RsmRXlQ4XF
prNzXY71FNRSPlw62B6AKsshftpcn9hsW/zmCTfWidSluTqn8RyL0y/hcaSfLFfD
4AxLzH7rB/0DgDDg+vBVOUs1XBzyVh0+LqA9hLADWQO7X1aWGveBmxEh5HduIh1E
Iu2IA9Egh7aqXDVwL9FLc6B0vJe9Lc7alFF3Nrp8QcrIqmgV11/Duw1l303dh3le
kaHGt9IViwQCoxbMcIswaKYysY67SKVf0CjEGLOorimdWNePMOjMFGXRiz6+2czb
Yis8zLJpqFcmt7udcu+hH9arnX+tquYxl8gH5hBb9crRvTljtrPg0q/IH9/7LQva
kJLU1+JFH3uA0sFnKJJTuqyTmkRniy9t1UQORjWRlgejDP+XC8SUETmj7mdFLmV6
GqnHj6RxEByVG8yFfY0IozzJUGLbhO6Sv8hYmJE952PSTXiYqLi1guJ4yJP7Qh2l
bB9Y5yVLVr3NKteTcTWl9b6QeeG+IXtCFqSKaKu8VZVD/UkUnKll77YjGka9BE3v
z1CAQEOtQTBhqNM2dNKIBmQqmE8SmDeBTzk8PhNFPISbeuO3usqYaxR5AkOFsUlI
Xk1CeLeFesjwVg+Bvvgk4rm0MLQQ6gK7H82HFuot55WpAKfRvEnNe4y39Z9GH+8r
+AAk2uNFi1WgBIx3NO/4ygBpJwxJeZkn93pTgLP23nM1M+1Xc0LJD8o/90k9W+Ks
uJp1IS1EN9Gl5ZemLpCYqTdrwbFgj6HMrzNHWtMrm5+QD9pAfMmtH4FhJ3cvLN4A
+C4L2/tj4niGkWp/GNagtHXoDbvUOWiw6enLZ4sO2wzPOPRQQTyOuHIkOxyH7id/
ii9H/wvL3SiRHXkvbVnSBwbQ08BHt6N0q9RPRxTaFGGMCECCFBzl/fMd3v93ThGH
MvwXVbjAW+Z3pmBhk8nDSS4f5ZhEJyrEXW73bNaR/6ojA9SUVDmGagTsz8Rw179G
gHwYK6bja5IAziQ3vIr/vgts9GYO4EGr7j6HKdMozinzRhZ8wjDtskrSttQNFycj
xaZjEjlbdzI/op/txWCpD7eSQWtfG8Ii2BbQs548LSQptNlbNhnV0I1kTFQ8MpZh
BWzAcjFkV3lyJVplCr//HnSN3RHJqY/pkY0+aoeRbtIOjO+aXU5f0ypL2lGQ6gtg
0My5szeELYOmZY4Uf300SQ0p5Pl3D4LzsWh/91qVTayKs6Dvpk2eHJps1AwI7ztL
`protect END_PROTECTED
