`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tCEd234rGPOtMNfDcYEYh9cPlR1lRKyYhpGl+56c0IQ3xjs5aWsfNGIfuGwhxY21
19Yd1u5KYOFjV37lLdT2OCEL6X+VJqwxRlsEhzFY/f4q0zHw6dRn6D2tj0sDUiy6
rbaRuEZ7L/vbLvCRKQVTeBwsKfNA4itR8tkgrZzFKrjNKt5W9JBNzlCjmap5YuTp
jJyzXU/AvHZEm32HpF6kIMOsGwdB7NEEJCTBELDLt2XXwUZsijk0DNhugt+V/HvL
YzTDB8ztnEl/KEeRNMxgRT3ZEvQf8E6IXYCCAMZzg6GUntafjb5odwSfaqqfXO8y
A4FFgIgINc/rbydbZEwe+1/TTo870fn0HwY1xCm2KASOO8wqzxPnDGbzuyfhcZKh
34l9Aomdp/tp5Lxi+BYakxgLNl2vum1SIBCm22rng2Fji0sTZFqsEBPScCPxALbN
zUzkqNN/IxvL8MhwWTDVHE5+jykQQbRIP5HBPbN+LM9gTNk1aUQdQZAQ1YshYUD0
uWUvvstfsynvDXiJL1eR0sbM7JmCzYptRlYXuTgmhPr52wI48dwbztQmd5qs5zGm
D1WkUd1jynkfAxMeONQu7aHMuuGw1+vbbiFi8omqK2p+1FV4zW7VaYdWlU7g71vM
3e+ohNVqouYhyMuap/YvlDtsjM2OJp3X3Hd3Ce5sHm8XZcE1fDCcQ++4tqd9KQud
7K7JdDhYcgdMcC8YyOswXNqUTz4pVdZ2REjs178xjuAgYyEDCCirz6eZBBcF9kg/
W9RQgkkw2VnO+oHxJnIDF/X4Wp5EVEUL2F6zIBUUwrBxiwzxIZiNMH7kR3hGb79n
xRnyotmvKmT+Zy7CpOXZ9/xi084e6BdxLOtzMEaNhKV2K25wFaeMRB5s0D/RFMjR
B5OKOsL1SWFRrfBVOvVkczmNUdUCWA+39wDEImJEMqtZ8EaSO/DLMhlVWePdW+Pe
eoF/yuc3HZe4Yul0gFudnpfh7jI5eorKt7jGPQwo2YucFT6WZABfkKM8PPwatdnT
QCTVsAjYKxeljKuv0LWJwU7kh+hULJK0b5OCj1tm6Y1H94lXjXG4jTGJFY+Q1g83
99gaFJ0dqc4O6I9F5Y8dIz+0Cz7lbSeEAOjtf5yLwS5kqIwkRrrikMfud5ujEU8D
5TwQtryfKKRtuoBekyn/dob5T3PjV+PBuDHV/epH5Wm5SguGB8HSEnuQAyWrGNeH
gNnyZwzNvhHgVYVEWe34OPuVTyGn3hI6hsUEyQIoGrP13Cj3ZRSnOuW45k3z86eL
Azc6pGWhzGJ2ZdRqG8IJ6y61Rq0lR+cqtF3Dh8w7eykWGN/goS+NMdLNEN1V9tGk
1AYfbjWLZ7sLGOieh0WUxQ2mYrbNjajBSdJcBMXrDbnjUfVSvBhYOFVtGNYhftgD
MlKSRO6HJjhSdOmQIz5NaACcPjDs5J9tuow6zhHJOv+59T24IE4OQKAHnxZXsu8G
wsGqoF8DUhHnJXjk5Ubcih8oUKzPXPLDrI+TIfovIx/aKaLZPwGvtnNqQbqbMHfe
6/r1+lbQt4RjOE7twwkRkPwYKWY7yOYGf6BF7m+PQwDOP2fLk+5BwxrjcMU3SepF
2ESMfXE9Db3aiD+7lKjb7h6CydebJSiVFTJbhRq8iXILgOzOjxep42/AGnwsOdCW
SpE3Z7QiTv6XNGB8vsxUG07YcErwhAF+XQT8Y4xLYmkFHVOExRhSnNpFjiNpaPIO
NM/4hGy1F5q7MWjCzZRCWCjjgDDr1Z8mJuPjukRqOLv8/l9j6eYPDIV5cfCsdv1I
/cnHq322xQCQqyZwn78B1z7EtO800DjH/hB9crBEcQQKBdWAfARjlB+ydu+fMbEj
vzXvK8+PKehqdgNsS9/M0Q4uzCGXeDJTuIXL9fbWGXUe+CJTcbMZ5y2I3plyC2Ds
qXqjTHh5HJN8bsFSjpEDda9t1tNas0mS97BNWCxpNySN6TvL0eNafqUN7gNm1aXM
39o4ipCDARC7B0x4TZm5vvX8ehST2stH7Iiy/eMhYY21kRRURNfvH5FmglNQMfQ/
z7TXd9g1ceGlyeYP0FFrKeG8QArwn/7U0lLoSlA8q101hy7mMxjcSteQzXZf/sQm
bYLLJmKD2Im9+z9RsdKhjw/mKRWMLfBM+9Zz0bl1m9UI6BeaUPT1TPgpyIrGWQnY
nV5vknYx7AdgeNOrZKP5rZAnRU/PiGNI/VddVDXo7qldZ3hDDaexgox3U19lPgZA
GXc1w2oljgRcANIeAQ/r0+je4SJHTc1m/RsmNq8JLPot48b/EJaC5hqjDEI7DQRL
yhAZm7bUl6yy6239Xfm5BJmOchgxd1QOPMDnMGbMDoS44GZg6AMuYbzibPCHPF9Y
iHRZsFkT8Jlt91FHYU4Tb4bY5Ns7xM/ZM8seWCYt2VETY3z5xsAF9xV6KUq7EUsF
HsYlLi0NXxmbNV7+irSwGHRakrJMZWgHi5Jwgo9GG8keCLnq5Dx2xd81juIvnUS6
J+ueslDKcnbg7GK707aTb3cgdk3INYuds6ekwO6YSfive8wgHmIt+0NrMNp+Ahid
6GH3IwTJ6UZ/46P5sZRCKonhOjjGTsAO1qO40aloB+0hosNvuDmOWeFFx/4N5J0t
zppFpTcrxBTdwEvxmT+m7ZVvAxhvJi6xwDCYhtg86vfxrur8YL+UPLgA+0EuFYSB
McvExiZwFp+AMPACVnlY5iyjXVhYNW1MIkdJvG39i/u2t6NwXDLYiRqHcuG2muIi
Qnh/JXOC1vDY7E645vVJAiT4CYo3Ku2j+5YVdbtKGDlOVsBfIryQ5guT94C71yhT
o/PQMJ2Vag15GHKGC8a+yhUw/+PPYjz0X7+aLwDkFnHVvUn3tjfCofxcIXmVwpyq
gThHydM7DRFrskseq+lQhtpzeLMOZ+SUXk83fBp+hLdgWIchxu0zQ22/9lM09vUi
24Cidh2ikBO4lGzqCzkr4fXTSN6qDf2dtZqOydbdeefvmooVa8MMMtewfXINGnsf
yFssLM57ImeUKjCUnIH62pl0XiouwxzrMVkycyGjTZiS+SwPUS91ecYxr6gmRfAk
E6Mgk+N0AeEdW5U+1xWEhN250rk9MjOvDbw0yvcgR6m6kYXWBH39OTDBR7sn3VNG
XBAJCu76737VI1F1U/zT9ge+h/M7edlNQIEWA5GIK//JS0jyIPHj68nC647amcNm
ralGsQ0nt6OEsH4AGbXzZtya3hA0WrN4qpmqqPD6Z3fQuuulnFitWx8gIEuc4ks8
FNFacz1xmCBivbhlVnVcT5wx2PC2fEki5Op78i636+AcrwNNrvgBw2aAOjoK9muf
6s1CoO2PtLQfSyhjlzx9T9DKhrJXrhHxt/8of9GNtvr+SAyHuXYETAaqCmArK+p8
7YiTUaszyjd2LW37DISRmtFJq2zG7+PyLqPzX45oXG3RFM3RmsvAd1BRCUxK7lc3
BmH6atm0IitBotSRIF/Gl2nja4EQyJo4pzQR4Vxnv86D27Rcu0LrDIQAq09hZ3BH
3+pJ86qItxgB2592xTqOA2w270ReoTQsxL/VowiV5MNk4v2/Bcor7d1yTOvAUhXo
ywQDlnB19JF9UCGSwDRRhoOLvFes/7ZosDH8s3WV23ywLRmhZ2DoSrHjyLu7bxmZ
cEupR1UknIO1fE5fMi8Je0WYilFl2wEUJ0aQAsOTRNTheljMpUWAnNgyG0WSaZ4s
WLZA1N8lyR+Yr8RchzPhkygkRlEgD/DMgGtwhmG93j629yP5Zil7bJ+mslShzBHu
PytzZogMF9JFkbh292z8GA4tmFtydVOhvbuIqcBeS7MA9elN+rA6v5Jz2XJghedm
oF7wsTZ4ltEYh0hvGXhOWf9UPmqDyVuxRfo8MeZexPMt39Thxjs3HFE6wG6lVoAK
TsvyyQhWjRX9pvi5oHuAEc0yRx2JdPq90tRFWiZVYhanWYQgezqwxlsLmokKP1ns
rDlvRWq9rI3sg2MPSzkGp2xqNJZswgtAvmYNzEDE1UMD0fTFs49PVuv9SHYJszsl
rOQzhbQNiE04U8JzqObyqyhCFEXhrXp9McY9bzhUX8gpx6qEl6eB+yROFSjZNBcR
9VUVqjaQzQuj6sWDimtRcVtLRAUKRzyHMtB+KGZHkJhWKzQ58yBVlEBWOVjHIm0l
EJ4vbed122oXGQqGMNNasBDVf5Rz1FQszSxrQNuMevCnCE5ogtGATpaQAqQ77qVm
xSA2QwLCdh1GlAbaz6G3r3sVb1y8ePa54NLfqiWVaP7t88mytpGXwN38JAneFL8E
ewhACtcAhFYPbjueGdQRRXj6cjhdYCxmVqaSXkPS780SMCuw60rUcIxzGvCSJb94
ybuTTF6ffcOJ4I6zAIauhQvmSjbvl4gmVZLBhUmQJ5P1vW7vDFpt15JrpVfp8uha
7m6EMvGSvpoSm/9MhucpK+fRV9Y4+FOLD73UHbQdC8knNS3BkKNG1E730Tx6UHIb
br/D+O65qajXMR1CYJnCfaFFkwZGGivYomVtaCHe0BZEIBD+737tVBGdcIOmM2Tk
FzJC5tlM+5mlwHsGfJfLUmJ5M9hqSza4chMxCWmYjqndv2ZbZ4jklNKZkpJv1ckh
vgRQ7/sFolCDgHo631fzGAwTxe/qy1UcsNokRZv0XpDGGs3Oj0lCovI4mA0HnxsS
/dEEjExa8szfvzehaz61I4Hq0MAr4aW4XRtWPci0LDqUkuVD3O6KlPXdFjjPK3zp
CDOpg/L1CLjF/MA6ZE/8zL2M2k4Xq72Lh1NCBtywkk7NDEAVrYFuABq+DMTabmmr
iyeosYZgEomEm0dROIuLJxqFqO5APjdbh0mN8BLZefXkdLXXfv2ssg5CA+4MmHmx
d4HwOqr4sxaXer/rbkYPoShYtsyijyaD2j/0QDI6eqAHfne/3K1jp0Pxg6MK0WpO
Vj7lz5NCxoW1e4eMpPNcPkvOzOOqpg/YuARIxjRUjTpDdkAakXl9K0CBiMKXJtUe
ikvoprm87LXg87JIBvhnm2d6cdQL6gRbIFgbMXc1CA5g3pYXRctQj7JRlrk6p83f
KTiVm5RDvlAmx/O8wQ1dLfDEl4dY+7rmbiM5HjBS5Y+tvS2sp17f61ndAXdhFreN
gTk+v+l1gAkgS+g65qDmMkoDGBATquck3QmneKsvOYulnd0v1c9FXtiSa877WBJJ
qdvIF4f5dnjnmit0Okj7HzlpYLe54OEryMwZ+YXRJJazpU4Cp+AX3BziHHIt1VGs
iw+Kf1AEVfeSO13Rvk/l/jXgxOOeiZESEjwspBYrbDa1nLATA6IW9O0CCHrO39QX
XNq+Lbl8xNrvcpWg969nWRzbmg4hGECkfWfwLKEixNeTf/YBOzimT6R+96lVc/1h
vREemeVx1Dmu0onHpXTA4wNtVCGlGHkng7tbJxQZQA9Q2p1m9tAvC2jV5VxtjjKk
zu3n6CSRnvspUTpUhq3/dnN6N10tvnvKmMivKXG3hxAbQ5lk2uAfcvyA1VHyM+Wg
DucxPT+CUyoK1HfwQLkWWfm9CfBI4lPhYu2xQ6iDUPxqnnZLwF7npw0TG8RXrRCE
QtuxTMrYm8n79pw09kQX9u4G8eSjnfjyEn+uNzO6Ib9tVekrcHOTk/Amj+f9VK00
trVeY080jyQy8Xu48rXpyrSJjUb2DXUajKysHWuRYFvAzHqlHfm4aDzhuBe73Rw/
/SH/iL+Pi4bpfQNCc9sj5gXKXK0pkXiNDreNIy+n1H9dxhhoZlGNxfUahGffLoio
kp0fgU7zSK+5zgqHuU40cDNrGNUSKH9oJg5WczusAt+RxSRkybCzobKQL5ID5avT
X0XHashWQDRM/YkKHrFXrSj6cbEjm+3OGICeiZFlpw9jvwil8L2L4cGutXfghUni
xhO6NijfDjTyVa6F4/YoEMw+mgGJ/pP/Ld9TUH+BVXIpdof49B9BU9dGudXX+ZYd
sXFWkDUy2+vynxHJ+YfN0Sf+TmTGlbjhwrPrsR537hWZjrEghlg6qN5VRQG7QW8q
cD3E+FzQNVwNc6Eim6Vpe9/eEwPogrP3+o1ePuVfKkj/X/KzCOXQ48SnK1J6pKgj
4jM9Ha2RNkW4rxh3UjGHA2u5OLwJ3RMHjLS02j6mHWYjeNX76yeVg19cFE0PnjYQ
odf7+11e7dFa4VrEY+Fxa5EIdkKuXdIGZd2BaAHSM27h+41E1DFpON4Y8D+GJkqM
h2gyOVYeTb2iUfrAnQpi+pwfgDvEw3TQOxorRCQ9ohRUXexK+BBIEZ1N7iToGy/l
UyZIUOiMqY7xJtgTq7DGAIn8nsW9tHn63Bn/05Xbd+64BF4aIDcwSGLcPti7q4sy
evADiGJ6Vs8n6jR35mtnIQqr3aIhQWXf5xweGSFyfFUz5C4DPWABitrh3p3otY1m
13kOdxwqDdxdIIAjHQCwiGjrmzFVklQWroyaBULs7EjHxM7pjyI9v56dJli6T2TH
YHGdgesdnTT+V48wJ/NQeFNyMnQ3oOTaWLg+JzJOxl0MO9nG6GVv0fRS+NZwF+FI
4T7IrlHNJ2ojOphxwtzG9SG6kHpi610XusPvdbaUgF5Fu86pHRekkexe7+3sntnK
ZICr+IReosVcTOiWl66ld8SfR68Taggx4+FilaFCquVE4GVHqWwGWdz8f5BmG21g
dvQJm2CladfIXHW+EI7KoV1zPxRlADwLXGien8oqetdylcekaJuA/pSIFLjJ2xK9
qt4OQt/suOExoaNWm7oC5z2iBf+kACA0l5wS2aCSamoM7BOlF5tm20JAVgQOMMBj
1OR659X450Hi7nhz64xEST/PazOz6VrmdwJRLvMa5db252pLDOz8Y1j2YCaM4HFT
vSkp9IWK4mP2cmrD1e00woep4cdm8X2ouB82QAIogA/GZ4f20xkw1MHIEHiRYK2b
1RPs2fhvFRF8HoCeBUAVjOpU8unAq4fFcZ0fogtkq3U1pxL+HUFBaIHQ/FwcGC7S
sLZk5JgM4jW+SDjWmZqOczCKzU2hn+2TqNosYhOJtXVItnxT0aAROMfEdV+keGGX
rkOMqB2hFzLqArA4bQjY/jw2kVsj8uGwxzD0WiY9Hh8=
`protect END_PROTECTED
