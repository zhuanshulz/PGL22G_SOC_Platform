`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uxh51b2mYan1GNGfC0tvpw0fp7CYIEdcLmSj5JEype+viraUgX485R/iYLS9DkM0
AJdgOvwXh7Njn82Nopfi1jAt9zTDB9Jp1RLJytbgVN4z2qvCRK77sfprcjyA69Ly
utuoeiHVRofOWXApU5c/DISMKSd6U35PcENtt652EKYVOIonz3xrH9O7dLToVyq7
vb2e1z8stq3CR3HVeYPR91WRJIR3qvW3PEQTz9RJrVjskWH4/h/D5IW8ekeYPRZA
fO0jw9qPjYeh9J4JYVF4/D6gFoIH0n6dpxDOgMTNYMgVO3A4FX/H3lDCqKVBaxas
E34luiDBCzopi1GHh13hGUVKYAkq40sxY+YUI42sKdyb4z+tzCXJzzic83348SnI
3iKfgJ/Sd/go5q3nolLPUGHvCAVswuspaPS0CZSVlCAf5h++dWeHXZCg58XQcTRb
`protect END_PROTECTED
