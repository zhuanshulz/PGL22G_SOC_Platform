`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBD7Ivm5NwNQv0EdJH8YAIrSBqAT8sW/AW5gwdGjCUYSZen+4eGOw2ZPpgyEPR6l
/WLO1D6eM7vmVdM9eb5spHZgW5bjHW26uKssuEOGijO9VcTvIKVfMtuJCzRZJ5FS
qHzmA+pCWRAR6fQ/EiUIdyzRgwAHQsnlEVcrO1unvaz4IewHv2+Ud8OuE15oNduF
OiqZJ1zBa2Ml5njqeYVmx+Hhh7vPUqLJeSHXcfTJ9UsXj8gZYSy17sGHFQ+MDDkw
RloIkrIxbFfSyw8D40eC5gp/OKrPQnWZ8qn/+YSm6uaZNXCcYgCUoYdAd9KCMD96
yHxLvcA7H1sInt4I8EMT8W7WNMxMEAjt4SQjQaF8PmrkkS5MYDK5hKFPqZqLugtA
bJVakSqyX1FWrfJEJ3GDVmsbP53TTlsFsgNNsdtn5v4kq/Np4IGzsb9bIsMN3OWt
7qUFW28fEQxDkCDnKhIOpUuYKImy+STiLUG5JUpNLXIo4ID7dsCRZM+E2N/2Pe0s
eNQ4jah0K0IcAHWI1NTB1ZLkDyii0vc9fJDzvenGFOF6s+aWGnMMqqphdm47MUbY
mSTIZCRqnzzJCem0z35OPfYlNZ3NyTfnmSiD3NAGSt/Ug+8NVG7paDH8rziIDvHS
TPJ9GdnTC3cTpb83QkWXpmy9y+/jeOkGLxaxHwqe1iIrQT+SECQ341GrldORQQR2
ZScOBHg6LlnqCMu9xPs0l9x3hvrhqeANtgzTQ5wKyxWcPYBTCeCV9ohZVFmZYhf4
kM9ywsjCgrqge7fAbP2Cq/b8Dy6KoscaKtiSNVjwZFt/lPg55n+FwdoEE+sd4+Fg
gm9zT0XYhfyNBOrAdaNGUFwbgMniihQ8CD7HJBNIRZC8qG1e6/O/tR1DYb3zL3fM
aHsT1mqRjWyyv2FUm+HdvALQ0u+XZd1GEFCLC+RxvYXd9RVs8cv1IKnmOwuiSa6P
dqt1xdOLSofDtKAy798GDA==
`protect END_PROTECTED
