`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1hj2EYerV0IdkZfDuq0c8Abkvzf96AFmWN2qDrwfucQOBKpCMZsoXU/ImkFVce4l
QBU+gLNU+14gktMBVs74KzJjrogCatyvfo5sF35wa0KkU5edL5Rku5LYWrv95dBc
qQ8ocMbINUcdxZ+m9eTBUggji2B6Xkm5SfgrbkLWvgF0wkI1UJer+RMH4bApjALc
MS1Zk4HYhQUt4Z56zWO0Dwtcf0gJ9DaKfp8Mv1Krj+6KgQUrgOnrUUpMtmsZ242k
EsYb+T1i6eurRIROJAeMxRzGiJ+T9sKNiC70N7RA/kJmGHdq+T88Bg9lK0srXGvQ
yEvrGRYdLUEYh1uGqLLhophORt4ABLPNgUoLtATyDj4kmO5WXXzOeMPa7Kf6gYCw
6O0JYozWyfk2goowYpwef6ItpRiayjP/kVstj1+f6f8jvIBfkjOBCvi8i/2oBWCj
6bwK7ipcm+nHLYs2lF42xn+RhClXUGecROlh6grSQboEKR3wncfaQLAIPi5nqIMz
dTWGXCRZbudLrsd7JiRZTqYcV+69NsovoIboDkeoxoqRlGCblzUnys34ehNVpkA7
h5aqnV0hd5RXrpbl533pob+nCx9YuiPUkYX+Z8aDmUzErp1ctRhuDFFD63p0fXqJ
IehMDGzlwCxAsQ0tzVD2jruVRZzHw6cpqIdDLfGXVNaqfqgDR8uxzL28tJ+mC705
NPJkb3MJvwUz43JjrQ0YTypyBHQImkCOGVoI9dFuVyjK5n/4Lr/hjYZbcp4Z7gdY
IkgQTH3t8mqLAuotUXaNQ2ifUrTasfWMC3V+5Sh5xC3Pjx6ez7ncR7JSzgDUCRI8
adUx5xc3qGcYWAMx/WwSGzQz/WyF4Q5LyvxTK04+RXIMY7hrdY4IYSVN7gEyZRO9
Te3jqy+jEbIGmXYPWMg3vvJLlVJR+fXjTN2gUK4FK7fMFj/JBBG0APAKvJdIq9y4
LAcTH6kt5ORgpHDy9Hw+JM86zEgHgPUx0iDPODKNve2bYTjNUVQstM/iBymDUoTU
qqUtxPzTQJKRyz3qeTJPoFz3LCFMOQdxOgEpYywpNMupgjyCT1kkgp8hc0SOYA/x
KR4wYpLYUxTzAN/Fe/Z0sw4ine3OnTtUvbDlTy9eot1F41jCWuw73jSEhnyyhKbS
wKCDFgT3vRjm20KASctEIjpZZ000d//oMqok0MTNK1VDXOPe0UBOvPq8wnTFuRuC
4eMHbR3aMKIyOo5tEoGjdaAGMpfLSoll/NTEyNnBr4FIRWejmfTThinvNe63x+n1
7Qz+YF2tqlb7y4Z8k1kBH4M+cEdrbQC/lPbBY1LlgkVJW5yqMBEn6mZMOtFDbdbJ
SPITog6DGxcuQVR6nz5LQ4Z6DUJCXsRWo2d0IAcJYwweXBKm+T6erKkUcWSuiwwS
x9RX6ozu9YdlyJHWbEmhlWPCP3SGfGvZs+9a2ivU8IkYMRpUAtAzwCJv0MihlwOx
Oxi//L5exPA4oi2lyXzZJhUBYIZWbJkg4Uy//bxQNPQxB2VD5qPH9q9jaeZLGpCF
ONXjGa0JXqVOk5M8af2AuIl2E3Lpl4+Fp5gIiKRm+9DX8/yacnV0bLrV78jijIE5
aRcC5HGZrTHs1L3stJcPekZENErU/PnHprRVXh2QkwWWW4fCdTm4MbWrGb26Dk7k
yhUWGrv/sEkeVAVbqhUADwXEb4h8rpUTw5iEEC/33sE=
`protect END_PROTECTED
