`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jboE5rJxvsKzVvTK1E2o4sfmuYV5Cje2qfD8M9li0PyB688PlbD9eqoGCFYVGZi8
IQhN7+blkB6SF4/OiUkwjpT1XxYHFWF7ueYxwiGOkXdrL5gCr22gH1OChCtltxOM
QkKyOy9VpKKATJchYBxy/w0O6E4OkzN4K/Q9EVUUOYMZWz6TWspNyusJUd40qQem
xly2dmyvm7nlebgne7nDZXbMZJJAwWTrOp9xuc1akfuVxG1H4shVHPnk6nis+lly
oDXVBq9sqUgb7kD1tSPy4Arp9wHT+Pl2m1K96juH2PDk1gKlE7rg1thk/WQQc9S1
N7ldpZFCnoAz1f27ID88Qg==
`protect END_PROTECTED
