`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2OhUPswmx3qso7h38LcBPgHhsHPY2lJnvwkd+yWhMTMha56NmBIJsRoYkk4U49YL
MKornSxfbi8guTrsyD2eUttO0wmW6WvIQYjPDKxY76XLYxj+Y0+NkuChoLhngZKO
C0TdCZUfJzYhzf/wA2HKBx9z7gPCzueBMCK4zncoh5LvQ/EPnnWTFeG1lDhDPiHD
sAYm5vI3LD3EUbFwa1+V+UPqy5KbqaKFPYTF4ouJOLyQ5XU4sevEZkxMkFUAJEEm
lJE0270utMAbUrkdVyNAOgxSBMFLMMDR7NfdxwdG7Q+UItndQq/u7AUrfRUBY8WX
Yknnbi9W7JhQAUOJPeEZUb51Nqkia1+uiqKBjQrD6ow7hFlzuZmEvxEM0oJtZrlN
YXNU8GscvWQVDDdLVv+E1BTgk2cRpbVH9JAB9T0Q14eS1jOBcbwWQkp5IYpxOmG/
j78knlNiUVuFQhvOavTMkuw2k4OFGZ/UJRFH0LjR9zSnh0llIL8yZ6t/3PIT0UKn
/GAsSD5ovaYoj/mlyiOkFGrxoVs89+AJgJ8RX+THv0cJSHg6cjcyDj6cYBKxFQpb
hTepdpXUDCIqXENgQ6Sw0xGHai7y70n9cQQ+uAugt+L6Adh35/D9pzXtpSlyLcBG
d6EgzeLbyOj9atfKCu2vxllzSMHEr6A0jchoAan+3eFiY9Pb0buleqtiKm0e25vS
0Ti/IrK/0o9QIV7PNeU6W/VCRK+BcIfZgo9wPXPjccC81vleVycws7CC2DayyF57
Vb5QOmKkn2XVgKCkqBw5tSrLOxy44k2uNbFqJkPDoF8F/9CsioySqht7O2mDYyST
FkdOsjbxkVICflfZpLjc82VieZJUztnPsuRyYV5ASjtvjx846XdBLnSoS8V15emR
orhgQ96EjhweS7f8124PLEjwqmlUGanXmlLqUrcO0lPC5bixEdutS7OsADBLcxY1
ax42HTIV1+zAX5zu05Oj/Fk4VwFwAqRmzrLko4Sdmj0lW25BjQq/WOnYJvsEUQGC
8kkHivjW9CuUTbWPMEQ6o4XH0+Dy1UDXVIYRJoap3v+uXlm365y1u/VtBYWebIDY
4QIrzd6ihTjCiT18dS0rc9dN4tZ+QdNNwoyO/vFr7fpmrcl/y9NYzUsmK+w4TZod
3X5UNYK9e4H8ikfoOP1NXacjsu5nYXgaWe0rIahaGhz3xIgkowkF3rMjEI9hVDy3
HjHWCaNLu2Hc/PacSHcj14hV0CZYDWlNQf0YASrJ3GCgCeAvfXJxVPJiMkcRRM/2
S09tkBPpwBuHUC5zLYwC66r7gmhQmYP6WxYSCzJ8mYAhXUNHepIwC396dj/UwgDk
ET5MqRk0STVBhKd/kxwCquGQcalHrB82YLUCpjTwtv+qKMuO/JhG1fbJYMZwbO5H
z2vdP/FySK8xWUaUUjjkG5vzOv1FNzJdAeodJMRoYjKsvQ0JkVAlad50/eKXkAN4
iJO7fDwPu6K0GVFzR1R/rHKTPYdFkefiSAycGjzGs2IFDYyIilDP5UIL7i/8xS0b
+sO2iCf2rDw2XVIWEdgLgacUd75sWviHWh/sYKn0JZKPxBBtfkOdyOrduhLcRafd
M3HHjro4ycUBh6yswAH/OcXJf5jYZan0LaIWriFCRXLFyds5bHJBcGgMHBIrq81s
6u5rHc9Wnns8BNGPmtBiwIvvJSHHBIkTwmsD1tGtKb3znroMZVDhnjJa5aOzR/dg
2ddcvqiKRkTzwhXmDSs+AXkIA6E0pwSFumKwGQSSTxFdcsS/WWbKLe8+0qxKzc6p
Sa2qCmkmjKbNvHSHLLXYcMPumuG+o060ArxXLmA4c1tW43wdzr6ApXyNQ5qQAWPk
nyHgx941U7OKsONYw1nsv30stBGkwC22ydYI4ihIt19e9dbZhtvigAq6iL4mXX1L
klFwK1tc8aw5QIoapTldtiA0jG+D428tnjTFVdD9ePiPea60Q/HDT0EFzZrusuqV
sNOL/Wgc2y4WgiGR748qxiyCF3JZhSxqYcp/MXC9uwVuthUBz4JIvgWn/s+qrvwU
4171rPXjACjpTAGDxoKhnsgel0LPcyZmLFFoTDFGhURx8mX+2VggMMDRmV3cFcHp
9C/fUgHifWSGnyd3O5wnNtGCmcbZUSi4XfXoFZl6dx+7DH+Z9/3xFNTmfNNGf18k
w/aTyncF1soWNJ0UtsfwPInuq0WjeSIk0sfIbg542dN6VADybSSks8AvDNtfbVOc
3V3ryzDxtaezkE2Ci+2SwT0s91PxE00GZDudXf1v0DhtWsRILXQDGnPXc3NZHz4N
rj3ITh/E1LdY8haztTRKJK4RkdV6oP5Ps4lKv1AvGg851rCxBqJRY0qxRjqHyKLl
ZYCHhYJVPR1gskvG8xi2xZGZF9oYbqdWkUzQRih7mtY4sjGiaI919O2NCukevNoh
YqeB8snz2WSz5Wo9bYfO6sUavFnzlSB+0qXiLBJqpvdZbYpVCYDUBzWAo0Y0hQ1A
WyON3DSjV8zFQUZbWFtusKi+GmJXok6q85OOtXew/4KqtSdl5HerPRGJMq7ZJGGs
eEc9ZGSeBnoxGeyUM7ppJDfdzPH7/hjuM4ok+AqNEfVNqQBg0gMfzRjAqfm8Za8E
mmgEtjOJYSYR37YXjh9HnUIWMxNQJLzFwVUQN0SNmvw0ftXJdLY5uy/rt8jmt6mr
hzxxUt4AK9QWPbUuUVaMkkFJ8u80o+25nSsWz7OWiT+/u4GGrPOVLc8eNU94hAqY
zz1/jqTmXOPbduhjWa/LDE232fuPeHho0mdwEqCk8xHLF5yI9updVtpTAmHurj9u
C5NMP2pxPocqoHV+tFsWBU5rhgXoQF9BfkTmMjvrW4vZqzhXz7Ld5UnFH3A4/bQQ
Xp4MME1ht+ce8G3RZ/C2h9mI3N+26N++rRk0bARpBakNESwC/iRugJMMgI6ZHnf2
2PVix3mpw00pQVSq3lBL9Z/s4LdcjuF8f6o42PCc4+Qu0N80u8zTby/ZcX6toyPo
iTD1zW+rAbtR9WfWmxfOO4qN+MCMcjyEaJWm2jUH8gejUVddgVGzYNUqZYnKh7L+
zdT/7t06T7mTVjLsQenhhGOxcW12z9YvnrT3ecrLYJBDkh6kQFmddsVXvYCMjxxq
yZdKRHEdbCJp4o8VXntCfe2j5XF3XVoHoMMjaV1ppkTaySbQSOTbUnPyGMz7Ttit
aaw7MY7KZkcct6NrDbK+sg2p275uR3Q9zJ7IMX9fcbXUqFIL35dG/UoK7LVdSZDF
/KjZucUsww0N/5EzMp7f7nj95ct1u4TdOE9YKi0NbAezx9MD7Z8nGEISo+bqZZgd
xZBD+9Hc4ZT8h9wY65BkggPDUKVYg2mjKzo4ROmOffKbjNnVhagHuHdKK0NupBDK
JYpD5GLQvPK391GTV7la1ZgS+1Nx6/TaOzytEaURnSSaBtSauKplscV3aoLLkiYU
9D+TjiAiO6X+m8+7UuEq38uzTqmtUWPC9dVEU0/kgP8F40AGGqbJ1cvkiNrKcRl0
loVePyvs2nZcOozoiDO4HkWFfxOg1CCOxfEUMEA5U8dUsW4LglaPoE0xuP3gdBCa
Bflq5zTn7uThKts6ktT3cpHWd20UFgGWtpPT8imnWDSMzRe9QYDSerOv2liJFVTN
XwZseTHUpxBhBgpbD2rlEkpBxVct5GS0MwckqhTWn6xYE8XwocTVpRCi46tKo0K+
xdx5plLHyAIsWRXd4a4ErikYY8EsXlPNr7wTiFNubEW8/IFplVb5+yH48rejFhsn
d3qR+Qe8628WqqYhjrCUE/ujqzEJn89IFXjj/Vpll4Z2PhY9EYe3BqBZXBtV3+vk
wC5HU06k2lWpZrxUJiYa/769+o8xee1T2Ebi/ool4Vdd72mgdA0mqpry9NrhW2Fd
ebzt5ffRqz/6h0O/PPQ6zlZw++o0v2zvYkiH0D4r8cKvoRmBEeG7FcWhlZGPMhg3
J4H9Nj0Gl1K3UaEY4NXB9cVG5S/pXuhzNFkamGhwHK/B57QXVUTT2EECNXZ6pd5B
rOJApqMzF6e4fw88us4/ty2Mi8NJkeDWiFNg61H5lx9keRtcV0wym/ESUzv0Db1x
dF1Wk83SSKfEGPy9o3a5hLw6lD7YNniSvnMeqSxNjWfNqWTPwlKiU/OqPHGARlza
ezgrKwR/Ch/Qr+H0KyGtPGIU6ErIWjZTy/tiarQyW0Q8F5/4TsOfID1FLxUcGwKy
uGx9k7hBLWGL9j8D9hjNrLCtJR63EpBmMn+BFvDdN3BmEJApVOP2ccDHN1SwU/zB
6XfWKjzhhE/Z0yjosFLwl/a3FHl0z3MC0MoU/hn7KpzCMYif9ZLRE+bIHIKJZiPO
PfFlFMdr92oaO5Xcj0umIXs1wbiFaPfYUKGgNahoctZ7FchIYUQl8DdTN62I1xab
Z7RiM5TT9re6j03zz6YIrdAafTXNKtVGM6lba69N9jbrCFcODwT/YyNhfG8wyhRZ
De0u+syxOVl4XaKzb7WAjJo+1bRFNWQGech4W42uzwbtHwhuJmpPcICaf2s2c6DF
1jNfieQCeNEXzysMzqE/ioMlWDL1nhRBJgZKH9JzienblLtGaYFiNL3Wr3r2eRgF
yrzfJjQ/BXOApkCb3cEwwfNA4fBpNIsO1SC1o9cCjowjbb4iKgb0oH+NLgANkmEO
daeM941ajUnbZmG5gQhH5XYTwPpdqi/E1WkvbPAgYwSar0qUTcUj9g0ZG6NLWi4F
UMXjsWGv/2h/pkMH8iBJibN8/rQydYHdZofQS808gIJiTtpCQs2IyIgZEqun82E/
OQW2LTPyWQmGs4OJXnBiIGyKcqpdj9Ge7i6VJElcTNdUNuxiBFETM5cL6513wmEP
5dKs6Sf03hx06fsA2CIgGQnATj8plfCHYWu6UIJLkEMefDtRsfKlTPl443GC7Ko/
L1GolXmoJCtXOquzfntmOvoL9xrs/9RSxUO1v9itMf0J0KI1SbtUMRO6MYkil9Wu
Ge8nBHE/j0iTxAJVdTJU24H7O2XdkqYYAYTBv7D2WwLw2JgqRJDgmTDVHk1iMQNd
3DYESjUy+9BKdxLVU5zaUauUGrIfWjoZ1c/0MEvG70WqP6GQiwO0Vm9i1vOWzYkB
CmJQZHEF0Gmz3otdG0NR0Q+5SAcEEGAjv2zQk1iXqucNVwRf9nlmR2o786DGV0Yq
1aHpGH0GSkk9qi64MRkcGdcQOWho88fStkJdYvAPYHRo3bq1+QFHpi94WKvCI39g
kLw/nQ2umpeEmXPKnmpTtxP+L5U0JEgj6BheAbRXEKouD2KNIRG17HCcAbHMs7xI
TXAhrHwy4o0MHauJdGTHsHWJJ1anVZxXrkoiNStAghHaJ2YDqRmvwCBARoDM96Si
xs+oJB2pVyVWtErRaecDkMPSFWzk/LFXmkAx21Xr3jzCHiBqPAsiS6B8yThYqMtz
Qwv/AISHqypSQ7P11wwADsAwf3rQi7xHuIn9M9Lex/eOeOQRf7Z/9Fu0elW8Sr/Y
yJ8V87PgU8ZUUOmK/zjB0xQMNvEFUzd6mYso81LdAypWEOMnrJX6e+Y6dOHEKfii
XhVbJrv4TaqZxQDaN83D/LjRCSUt9wLj+jPpNXmdfRO+6xeSzyTOgI7SBnrWTSWg
Q9Def9o7WwgkMTC8P+2ewi1Hqz4WEoe49tsDngntoaj0chwMTWBtACrL0/OaDLXC
8Wfb7n9pxm3ozdwZa0zg9iq6E1XQBsumx/wNkSqU3pr7daBkktTLuHYq8PIGByED
4rJ9FmbUZMKyS7c7BZm8CMoE+SIukFPVfoco4ygV/ykMnWUR/QDSUrhN48wZ1sj+
om2kmYcB3pobcaSIcYFk4wzTJnLJr9dDS8pDyju1ckj75Uf4xmEqEK4fZHqQ/WrE
FKniuXiXGHBnStk9+ycfNHGPfrdBRA6dkDtU1t/TPFgGgdak9gxsNgtn7frKSEmh
8cf2kdQ1vio4Em8GbraXahiBh8lHrZDCAwObT4VeJ1InLEcjk20g/c3Je1ct7b6v
J81NQLtDehp0uLPY/oAyHfszE/0gQVvfsHRIvIyPUMArSZ8NUpYkU1ItRQBwEtK5
5HoLaTVykF8JecWqXEqYj44oOCvjSE55zjYIy5qsk+iq8Bv0xxkg3Ph08uafrEl4
HmXhDGaQWaOju5faNeKp3NoydY5IZaId30NjLbR78VSLtTMcpLuSCLQxbROSJuNR
bHZv/PT8/1iFGjJDUYMZQFb48ft1lCb35OQMUYJv5HSWPD+fcfSqauEGZnWsfTyX
bPbCK8CsqbAgSpTMAJZH4v7o01ct3gcgFgf50N/WukceG0RJ/fMqDbK5eZvWsfup
mf7igSM0aJhqqAehc+4a1oylvz5EF56wxenku6pv+E7SZXabWj/2ja8S8Ymy4i2Q
L/KGF4FHxO1SJuVBn2ddiHIWc3HSMwRWEOVMy2qgloepFJIujl6VnrWWSSL3y5sH
Y8UKcL0MkQUNCJPIJRk22QEzQXT47VdilY9C+c6mA0HYU4YtJshLU+7FDyl9BI+X
4mx8LGbexw2yXqIBGCnilJ9u4mT5LoIY8v5y72mTJy2UWS4yZllwi45uxSezL/Mp
Oyn+sQECWsFTqvYcvm4bITpEmiDGIhZAaGRXQqgoEHa1oi/gUnKm6ZlY6E1E38j6
XT6vXNKxbGFC+5Rh3zx1NzJKxt/yAp5DsYxhSSh4GeuZC/gaBr0C9Fqu0E5TBy3y
a9ZXL8n+IDS+aQoKi/tuw4ziPXhNV+28UGrSGBOC4q/gBVCN9GDuF8NcGGjBWlvf
Ye8N41efSgj8M4WifmTno6IDEbjYeK23x8j+d9l13/Ln3t4+ZsFXqPMpJ8wOIlWP
ourFrZ4hr1G592NAYrsuHmMP6CiRh0v5MUfUdTXjUYnUBnRHN3PHfEKTgN92eImp
E9Yi+o4Q9f1z7zkp867niI/1ECJdCsk4dsKmIazjFYo0hIpgT+mJ/ERu27Gulvz2
ftfI3FT153TkqDxaQmVckbR9zQeh6fn2HRppmimbmMDTByb4NDLdIU4gSwjdxBmB
MUf1v45SmW39RCudxAXEfR4WLA5FxCKq5Gsd0epUqV313eZRWFOTayfwr2FfNOP4
SwhRgmQ/dqVv+UfRLIq3sro7SRwQ7bQT4iEECk+9SNBKw57qbfhVfaLb7rEjT/0V
DQ2fYwRpzNOKGJXfnSborUrm/nLHBxhWJbpNpgAK/XfhD7t984mcSPlCOX45y/qL
lc/CRB2P2ZWZu8kN9lFqHHpdxz/4/7EnrLU6eQf8snSc1ucVugISXu/9tMy8byPa
0wnm++4Gm3eYER970NHMi9iCibW2mMIrb3WadB8J6i+mB+XQ+Ltd+nceJHsOQvUB
AWtgLOGyhNbyLYqRCNTvU/PXQ5+AxacCRXsTp7MOUSx9/xE+FpK98W75lgEPQIm9
RpLFcZBpRorlVmJ+4gHR+6CJ/dhQdtSOAenDU/ibniDcr3VPz+Y+IQDKNzY3I/hI
ixr/q4HU7UhvUJbTihz0UWqh73cBWxq6dRFnHKvctXd4uWr7QlqaQqozfZlLRGm7
JQacCb38QD250X8a3HwXc0r3P2CGHo4vCcD1wL1sG+WfItI3eagSCSS2eXBUM6Gz
JvLoWfF1G/vIsVC3c+6lzrotwjyWFRnhKi0cIDCBdUwILnTW6fNmQXKx06bbt0Fq
AICaKxDb+LYK/uyGa0Z33YWuNYhgyidxVZPCnSDoz4c5FnUfqguE8jP6/TZBYJRy
ZAECFzxfXJ6of/CRmj6iLSUqVNYbVxSFVlhVxyBggffSfcwHts/6M22a+0gZZTfj
OI467LHLhb4cQFqGNtEUX2igEHyDzZd8LcJcaAcy5ccpA3Ok3oDjU2bnp69JusWz
QFyLQtVSQGrfaP6EB0blRPTobuAPX+OvNAaIfcPI035OcMRDTePp3keZ/inDjr3G
WVeAsvp27u4V5tJeicDthzKT6Q7850Zq79BZyK5WLsnCjMRslMGJtdtaZtKlawpz
5JVuKpP1Gy4nMVspMRKcUSk/brC5XanFsVYU2mUVZv+Hf7eeJ73hR0V1Fmqto+ZI
tut/2laLdfpXe+EmPQRCavDzUbFzffjZtGbH2A3tUiiwCMoHxfV2OXUCtGUTrveK
nmy2byhx7K8sIxdtA5+r1x6SQMdX07Xs5uK9HBYVOhv+s0V4aaLm7z2Dmaa6ns/b
lFp8/z9M37FYdWYTxcj4qhDa9ijDpzlhp06Qgz6n78cm6pNWGU9KxUy1NwgHzYRq
ucmfjTLwzWCeCMUIChlpV5wvFQDFkDTUJm0i48lysM233WO5U7CBFWJqmb34kUSi
m8HyHezl0JIW4vccViYUXSM64xAS5gImC+VfsDV525sTQfzHk1dUulyiQEKDvSA5
4iu7JlEZcwbmalaGiuZwTvI1UDqaeeKyRfTphokntKAMJutSiRi47L2IgdYOuzGo
th5cKGNtdSRva8HPEKK3/AJpCEpZc+r3LU9PxcZ388rGsoIVSgN10xeYcuse0Pw+
3OXfQ6Bcp2ZB/dXHvGFfov78Lm0VTEyQYHd+AhcnENfpjNiwaaQ5yXSO/y2QS5vZ
3E3JcIlokBIOZ3z4OAOAJDnXHQUPhm6teIcKiwQYDpq5L7+XZMEERetbq6RamLoK
LmmfFwpmkyDM0cxGe3aRxADG+pFXudJ0pEgUGVwF9mtQ6+4hCbAKLMBZqRWEj16C
+G9EeT3AGATubo0X19vuvKwsIJaW2tSw1u+EUbEdCBsufrw3VpFk1LnGnyBc3a24
AnoFmOj3YtKMCBAvUswD2eX0dEuxtWo8+MQ5+jrTFKqK2BjzmbEaChuL3Zp4yuXD
ckfOssc5IMXJDxS4gyMV1u/5WTvUAibLz7GO2v1hul9CzfI2GCgRD8PSO2YKestR
rsXV6Bu5pm5Pz3ZvQob1xqkghxPNAbIe6MOa2f68b+8s+IEADjW0lrsIZMLsjQKF
csr0jzY6n+biLL7fK7AWTGggjTYC71GFwcwYX59tz+8mXpkVl8W8Jo1tcgO6leCv
TTCatc99embcIFlnHrD5t2AFquA4Ce7Z4g/X5ENLrEJ42+u7qWiDTE4wxlZDgB6M
CyJsVTmxFXfgF6OVYBVSuevhSRf0thXweWwLoBqeXoD/nzLmHSeWrxeBDSKq6+m/
CLHTcgC4F2knxB3XvB8kjlczclrHFyhkuKCLAw3JgBX6/U4uIj+uHAeIy4LbuvQu
B0+a1hH2Ryw6rNf5mbm4ZZ3I4U4sVt4bJ1hrzFw0SnqAttVlw6Abmlzw5ZXpsPxz
wwGn5uE9Xf4wUs76yMdpFg0mJfulwaqX4I4lD9kkbqvw2dHohPQ2EJRzRVw7Hihf
DtvtVKf0rK/HlugzexHJSgCaKUg49YqZIplwurNnFOAmdlTgTPg90AljrGqT3woR
ueBHTonmp+8YO6vXEcsxpK2Eq7/i2/oro8QbF+/8auI07VFc53UCA3M057dEI2Bc
+9IPMF4PIGnKMemZJWcbTjyj+54WZX2z5QiZihfQsneh0uX2lFHGBEoMbnP0hUK/
4hix9eh12xkJFBX5cg649RaMF87iHITq41EfOmCL6PeyEekNcf1ZbkxMu7+i63FI
hsqHCZ4VINrPaX6K52CI7xe9m2BDJWgJDJe4pNqOVDAYONNXMNzc0s1cSMzWV9gJ
GjgEpytuWmynWnNsbzw7TO/YFiu/gg2DTFHdgT+71SyXhXZ4q5t/9el23A9M0Abw
WTp3y7Ryf4t8MBlDVsF9XNYwitn5AXvRNVbUHzQ+2+6gq4rQlWCOzqSm6TpbksU5
tmf4JTWBNb2g/LuQRpctw5KONsUljsHMBRC1Ar0x08rpw2kecvS32zbM0XPBgUxy
KIB2vrR3BxprtAxKt0AK5+e4Tsw2FBmwnSi8ZPbeGMVhQRTFUqx+NrUCOrJ12pVi
N6JG+CN2V6CU0TAPfqvQbTEuGm8i6yIXXJPutW3xxasFeaoUmPG8n2O5rctIcZbC
M93e2csjvbHCZHtomAE1an1GaxbORZNVW4y5Tyyay9ErsbxVTvy48JgD1yLcV6Wu
LfNxSqoNvumMf3r492ItGjiEuMHnUVkkCmGTgNQirw+h/kC0O4W8gMEMPLE+gmld
4fAH2k05xbu4WgfEiPU/efcDOrLayHN8y2YK3dQ+L/C4MVKKLivFqcXuhnaxTY4r
fdNNwXb3DAaMdQb/Hr0m2aN+CTZs5Zl3LrcN6x/L/GGV+eJFsiH2hN5EOBj4jRWu
VN9EnlyuPeigo9jGjshH0WhN3Nena04k6hlOa+r6NzqbW0t1LzyYLqdBM0lX/VlW
ehRxM+pDKyuk2+/Xgm1RNRjLM/tyVSlJub/keYq/d5RXX1m83EiJ/Mmltw/74b1+
ZCGO1EUEPnyvbqoZ7gs4p89Do/0kb4VLILeLRRbkJqE0r9pb2gwC5g93rkt5W/if
d4yYaHEBAcp2ZzR30cih/1Ls0FspLxKKOidko54F0AjAb4dEdjpkerj6MDIK0aCL
9jKvuxWDt+lMlNVJYkzrCsZLwgjcH1NsX/jXRRoBaS3FeiplVu1grnyBr1wsCyc3
JXB3YQQ0OfN0Pn6kSdwfcfky913vRnoswUrS/oV1uOXbiekbydbZT8/kK0LunYWE
Os9bW6OJqnbqLjpbIJfUNVIA8ZUSzKQ3rG9pROwr6pxQlewGusO9B/zKAqTt2azx
d4ktlZK+CTNa+8wxs04JOuj6Hfg9QkQQ9fi4jv2YcltArrA6dWmYGI+X67m6YbUQ
4btPO/TtzZaAOyoF0/kf228y3Zw7IADfgjMAiWMwOmBLzAE0E5oMKZSUhrji6D2B
lait16+cjIpgokzeVpSnDO4Z5BfmsXwV/DbigyzY/PVjsE+5+n0EWGe9u0CyTiss
ap3YbpHtfV5KmKEIdJQMGJtjs3TdpIv2CdvlGg/tG6cJyMDR5o58hQCyNF7cTmfd
Ls1j9Ztb6NF87dy84VBMNeDYEK4CvMrvN7hFsncSFSCpMcK5jrnqnYWE0JCNabn5
ZR0YbeIpoOld+VxzWXiAP/RB0VCKr17a0BUPZJFXVL7HFuZRcEHxPQZIhgCOAarh
eNMLGf68Pz0aoMHALS4JqTiPDh27RKqOv4IMpM3LkTcWI7RlEBq9mUYP2BRjLo+p
uzUh5M6lplbJCleTImM2tXYJZs1OGqx6xms3bW9ornpj8psAlHTV68QhnxNsWgrr
+FNiI4pkgLAOEEqWod6vSJi5htb8kH8xigZaQ4zA3fJdkMLNHRMgw3gWcj3jdYaG
wsV0IGVGtfFqi8U0iJv9GBYNgbRYGjG5+SnoGfU+kDd9QeDX7DOlBOO/twtdUye4
yjmbXm/CT+z0rrNARvKAyCD6gcpaYTBQAmH4LFwf8z9rLrmTH3ifRuX9zUqg4mXs
2MfvUlRYPKsAcAmOZXYOX0tTcQj9GH2SRuClbBjtyUG2zap2sUTuTddD0O04GF6l
LVc271LmMYYnYRxbwf562uzcdVB/vyiI6W6LzMeyWP7RJIIdjJk5zoC/Ax8JpO6a
hWQ0Z6cwCwdrV7ydANRZOiPt9wcM6cgCiri0pOGoaKH2Mq6VrgzLzhsFQmVA+qjk
dic6WuXIndffmsRp4GeU/UuQ1KUqdQoAFc5gseAzcDZxZ5B4NxrZUGZNZLPZrmcz
lZ2eoOibLtFsQHXNgHR959WX1qRRDLFthzXV7CtTVZ5zmAWzYBjq729uuRIqZTGL
uD5nXR9ubGvB+4xfYSyuoa/dpgu7foSc84UVHho7PuEqExIX43/Fki9WNaWZdO/a
2HBznHBt021cnb8JCfTqROiyri/HjuaTdp29/bWlt8hAGvoFYxiBG5chz2nLJi0Z
JXKZ7phNYU1Z+ahCAb9YcKgh/oIEcCKCqwYGdpGuJKxU6cuFqeY0tCO6S4dId9CZ
dJxzm+fnXIOGpPQiRuMcPaiqR2AiUbEB8NqgxMpTYD19lSMmqufD5QDtAyCq0i0A
AtyJj1PbFzd8n6CpGZyAtvl/DF6yJUGJWVUry/NkcF9iRgieCjb4nddyhj7CKHGl
xFGIy472Zj9ogb9sWhR2nd58S33ARUpl9lA5WJFI8oyEDxjM3F9HHI3sV281Ihzy
MIsTZrMhlJ8WEUwqXXm6/75JKC7+gN5amRjz1MtGPWRXlVoeXlSBp9U05ZW5bahS
xjdKWmMQNDAI7/tAsO6gshLpxj9li7KfIkVi6ThupgrqszV5SI9UIrFK0azIpfRk
A6DxXTh3k09QPsIorx43WivC04n/W3wgJWIVKyku7GCyJBpP84u+GDUa0g+kKgxe
QaEsmLI3bMEn8qVHO30z+WylesbwnqJ9S9F4tW7M5pH8L2A3i+4dTm+L3oDBXtNY
7/tkzqnMsDnwa/GcQzYxjS2tV2Khj9Vbbu4kQKWaGSTSiFuyTIVovVtysmNjhbdU
C2Ba6ucYfnThpq8E091wsXT5JmKtDJ4ukmH7DJGv56eY5EObnQ2hSZi+qj1LrFrk
06AKytgD0d+aAOJsESdHadQxN4noeO6yIvn/e3nqHoi1bA6fUw3fpeHCspP0KaN8
kpDyosZSP5UYT6uzqnE0Z+tCwmA0751W3xx3SFgqPp0Mn/UVxgN7X/htUAbbAaA/
Aa6cbup0+hIh5IZV8H1UJwiLQrx1OWbdTCWDjl6NS1IOj9bXx8Kd6XKzBm3jB79y
bH5jXcmbmKmy3DflBnJ8jK621K+uyry2v8FDY8yevvnJ61ewZkBRA1iH1CilajVS
OSzI9BopMLnK20qjKpv/JTDozkHEaRd1Z6emAGvki+vneHTsVEpRZEIkp08+JbP+
uCanq+wMpAz6l/2ExzACvYX6EovMJNwctS0miVZ81ZhMKif2fAsg1nr0o+x3Exj9
Vjt07HnOirHPPDZqcC7V17vUHyYEaaXXY87RePBX3Q5v+VNiIEyqNLM4tOs+pahe
xbR/3c4SclX1l8oCi/J3UPMWktuB1/vLJEKJ0v3v1Mq5NxnindSUQb3uN+i76Ypm
Hqh78u8DFivG7X4Bw3A4fAVHtcBQRDm8voZm8fG5gb6vMQL4za/1POkcxVyQAbRQ
0tpFWGOfcOXfGkGsCJQQRLHMObiiPPwDK2K8qW9uIcCzim7B5VNpn2L8h5eutx19
Fuq7j/LBGoLTU/jJ9XStb4x7tVooiL66d3E2aLUxQcVualSsmS8lKAYzBViK7YtM
SV2aM0oUiLFEryQtzHtLA6h3bvumCFBR5lvDVmzfqPtYeqh+ZmzemDK1MGp1m++M
0olW5iOIvqnm5A+PqlSk5RrfeW/fxeKWBy+OTnDtkxgdlYmyj6mohG9bWcbYLPgR
pZJlK6GgKm/TBjhwpDeIhgvV1AhD3P/Y3IuybRN12+qkfA5GEU2lOlaY9OZ1EWX5
2MKF4yfBzUhYt8ZTahmP6jejqiD/JjJsX2mvT+EuHyPJ2tfIezvBb989m6UUcC4/
cDDUkxy8zA3/E9ImNM+CtgvnQThUU6swk76/16s2F87IiysXgEH7Wq0yo2dti8jB
ZqO1n7oXzz8ohmH7xBahIZUl7A0u+pFlX3Qyt3B38m1tzMLlzXugo+ub2hQj2x51
ctYvbAjZoljCd8nhkOJ1OTpPQT0D8zqlDBF+JqK7KJXq1hhTuoZ3Ear4iMVDcIBJ
3Vh+KG9Ay8s3rhDyfedDT8n/M7zHwUTIm4m+GxZRPqyQPOIAaxj+M253cTqR4F7b
k+XN8+mkBRWPK51HWtVgTePdaYJPXLvtJ0WLElZbDiwb7kXjzhfleG5400MtMvL7
gsGig8tElUrd9T7JeAh+O6ry5WkdC/8kWSy0nQKO3x4yZ9qA8UDy3vIUleCNdP+P
qztqDPnlQeyIiRpzUdL7oqfbGAZ7KG96KiDthUM1xfXNzd9A98PSenHhxsvTyiNW
USnUyi+0gqI7TW9QzMhPvFe1liUXbYd0WGY9CothU7vxNj1buFHllnGjdRYqysPB
LOtgKUCwvMPWNdasw0+OAbnl16kF34tscZevAtIkM+D18UhhAwp+IHBz0UGyXxC9
CPj6kCtuDaKPE362AnfMr0hXhMp04jb4cztnMzMdWtPEJXYfKa8iF+X+/uLdpC56
g+BYY7tN1YO6wVTFj6gS9fIMJgQxZH5x61zRgvfDo2K3GuUliFngdKIAeNammSBM
3QtE11Fr+26Aoyq1gGcxVTlGNy2IrGw3GtfkVvs3P5dzr6t9mJ8tLKj/qy9LtuPP
6md4QRYfOKnRy0EUA3qEpjHEDnFOxH+cdShOJjfpYljAhucsS7R/R8ogs1n2Cb9D
UeWzUhcmK5GubZAHV6YDnInJM7Ogvsa1jKEb2f1ja9nBo5zcSCpZsgZc9O2GtOmK
CQNTLVw7w8K7uP3gi/8MKqV51Sx05yizwcrhLAW52aKZEnQgmOxfGH/3KgVFboC3
8yh6x9xLNwC5qHHZM60YWXNwNoLMYs06YPn7VRc5ZqHl/sV32txZ436L6Ql5g9fy
znG+jKi8Xm/yh5ypljbuQ/31Bfp3vFPu8cDBHI2DG+wpZpgdQwxblN1xm4VjzQsY
4bY0AQ/lBYazF1cjRJ5e1k2IkQ62jqmauWlhiNqX7raUH91RNjcs+ryQyljVnN0A
yQND95pPGtemw5zb9hsNGEFROvPQam/wcbFQ7hY5HU3mV0+PLochuTHWEi1rIcgQ
ZdVz2vHpf/JZXfZjVZOLNIrWuc1S/VCsij5AyPnbijrh92gx3VIh5p+BgDCGcxNb
kntcVZ99MXkZ2k5dNRXaVoh6lOUL0RuiwJQvjwdztZ5dyK9eB7OSu3Db2/oQSWKa
62o0hBKszCeEIRm/AAGYU6BljuE7PGx/hvmaoQb92B+0EWpyzPmiRcAPzC8Z4G0u
pjGX44uO8jpXtov9MEVOeS8iVtVNuFPao0/8xDcI4xngMLCUHaO2Thnltjdw/l+e
DgdW6ddCZgxrCWyDYN2eSiP13d7S3SNj3z2kxNZQD2VQb/e7c0VcqeoqU/jK6vQ8
ysX87V9Ta8yy6OnISHwFV7E5MZmkZ36nmFiTLf20B1SEDKN9aVI4Hft/iYcZljO7
bln7lv8CUy2poUreE4SlMHhB8Y6LW+yXuxOKL6pkIDSl8diIHtBd9Cjz7yrX4E/k
IgwRa98X3r3miCKYX5HmqEa6zYX5Ui6S5H+catbcYL2fm60vjcepIOiqZi/DEgaD
DqHyjzOMKQkevQAzjHOq4LxAOk2E61qyhJ4dj1Ob3215a2cFlUV0qf6L67jKdkKb
RXnArKfwgQV4zsehFPPwT4Mq5/g0JrkV6KFDFiavquAbael7kyi8dsFYx10PeowE
QO5sl/Cf1YpHvYVxtcIGXU1IqVfmWMhKTz58kK+BO2HDZWvvyirF3EKNHrk8cfef
oPfCILnaL5Kap15ACKS+ocnAfDKV3UHPxyZcihh6Xmp2cwk9PrnXbsFaUVntp6Fs
CqdVOF1qxOJzHw4wfhduLGfCHpCTIGtorhFLsGrzJBzCRc8GgBmUC5ndemISwVmD
h5ti53RGTPBSuLtLujnXGqZjms1PGLnl8t77hfoUxc7gzGRWSDqdd2f9u2winJZ3
aUaJtBiwtBzNZ/rwbkwt/MJpUTlet7fM80sWTv4mqEozfTTItAm4/M/KqA6YcPyY
nuk1D427cDDMGYeRqA/zJ35Va4cICtemaa9j3pdnWZt5+r0cJ7NUGQb27yWt8xKW
bU93NsilleJ/3f/jj7ea1PiEJPMN1p5QCR+Aa0BulYdRcT3SiNqZVt4+QVDrB+oV
1lYsefJlEDPqmPXt4LxK8scuCh6290LzoR3dHGYFgG9eppR731pGWhkPd3i2pkEs
Vi66GCGH3LXBdIwmlZqCwy6khmrNwSSQEYhSVVQlj2k0V1iCBNSCmR56BHTFEeM7
gQZET77RZgY2ns71/WT/eI7SrigPTnBeduD1QpVP5d0wJl7DUAWV4F+wdYwG8nDT
SnS5RnZNDMY+OaKSxJ/e2uECyXkUCQCpxpAgpCPgeGi1lGALdPLwixBDZd/Aej9e
ABaZDpJCZMJPwSgJ7zdlV0X0gknEOpARhzQrQblkj2gvdVAXdo1OZnL5ezB7b3+S
SbklwMCWHbN+MUv8kMl5+YMoX9ibVOK6+tpTWc3ESUmz7m+6AwhbBIGla45bOpE9
+B0MhjAlUBy/rnRQZxzvnVRQOTHhg1qYcIkKtaWieEL+AOSfxCSaJJfDLjQQjmYw
eGdjm2DpO2v//ydfcHd0QdxeJPK1ZA89ZwS0b7BQAXa93JJB9y6ZmiGOFEfKdUW4
8+anRgKXmBFeCHDWvPMCiTradr0PjEwF7iSYF5qZigKm7Y2JRfqVd4uGrEL/iTpv
VDAA6wEW4+PpVNHt+fO07Pz/aW/qdp+TmwOFaGWA/cVlLn1nl7YgLNbpC/thb+A5
M8xIT9j7PWbb5fmHjHpchsWC9UVSJdxTXymPbWGkK5+ictTLejDXcqDU68EI3X6t
0AXHKiyflUMab6WHIIuyLHlaGIv4cHdqZmhtMgls6tMqd6PioKIwHaEuyBSzAxea
bvYN78+4gSJkKTKETRfzSdGN1/hEtp4lF5nrN5SiNl0wukWR8FktkpON6KWzBMTo
wJcyeiOqlSblsw3I89JpDPsABpAIDn6jrldk5RI6lg9k6BgvbTTk1C7/IYx7AM+w
Bzf5ZTYAgOe2XgxrJMhahWphEisabO7YyuRQRvUWD6BZ/23aIVvOVzu1CBD3JbLf
t2PwJ6B5dotxdLfCl8m4osVoGyFydgmFio9/Rc3CgReJMGLu6KiPDt1I0rzlXA/r
OAoM1I2hAAErDqJelg0Ov1glaj15QmBARHogx6I52sjM8RvGy/Ij6FO2CrmhcNZy
ryFDoFIh9wGieNxtqTKAtE3Y/d+gOHQqXH7RRSoCqPUPsh4FTCSfWdxXXm01QOTo
q/u48BiNNyu+MtrT8bErz91k648rdUHdFnwij/1JOSbK+izdpCuHK6PL3xw17jEX
5Uq3TZmP25MuLDjMY8nC79p6FZ/byAR5PfYPpOZxps+tWd3SFhZ9WqVTfFpZDXJs
me6LWtdzFxYCL3nJVXKZR4P8C/tPmRE26FX431jlyvgGYs1CrY7Vsj7ii5PhGr6z
196JC8ERJqrQzvYO33a2YvA/UF12OWB5Z4JJi2KCqRZRzW+BXwI+iwSexAXLEU1o
pfzrWRftT9FxUKnkNMBGaA==
`protect END_PROTECTED
