`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8GoQANUHUqCGUP7I+ChHp7jouhXTnEI++DoDvBxACytB9iXESUxDA6zfPMSdf5XC
9Z9azWIThx05djJZnAK/ul0eG0MvoF5PekUCQeMQgT9ywXH35xYkgj2GOh+XowVk
e52SYVqPvJzQh4WE852TwJjPJDyYG1O05fRsgFLh0lijqPH6n1wnmcm+n+0bqxHf
jkxLYHDEH8zOehjVo9q4FNtUnaYilLp7IIkBZf4WwlACdyEli2U8tDqA0XRlW+uE
TToD5nHzpe0oJWSAnPWmj59Y/yRLNIqPossYc56y7FQqo1kBM1OtKMLlSs9iTGQI
G1CuCDoQMPo4XsXCWUfkOEc9D+D4oEcIFU4zK8Eje42pc026k3/2L5ypnc8FQKRG
S7l1R2iXNsjPz19+bRkIL3TSq7gzsZv9MAkiBHBqojWRDATFwwc1bEG5/e3d5tBK
VVucBPAz10PgK/RsiI0mX1C//DyYoeDrmanFYMv2zffQMh5xF7qoW/XXzGfAM3GY
AW8uYk5HDgkTkVkYWTyPSfB0EwVISdWi0evQEYriWWl47rHN6YIz0tegN9XueAqU
raTPf8gafbGo9fhVS2M1ZznkpCFWhKvKgpR3pHUzSK0cf40h1nE4VOct3p379KWp
Ddep86ZfVrnkHCQvtma5gx7DHPffYUe8+yMtAqqUBaX5qQwGC4WUtF/ClwyRe09F
EvBon1apHv3+oQJWBxna9xflOctg6rIFDeYXn5yjmVcHz1wfeXUS1zZxBJwaBk4y
u9lPKc1g6BYdus/5+/saLHLyRx6lXBAIhsMQbT4tCErNjxqwGZJV8a6IW9mhS1sK
mySf+PjSMhAogeMfu2UlBBC4ip+c1+hdbVa1GennY/Rg8GfR1wL27yE94EODTYoG
Hus87iRFDZVqermNacSwgdUeBg5VC4a/37sTfUImixnWlF54E7ZPZta2t1KCbwwv
kWCgsd28c0Xthzg0FXRrEJGXRdsVEbXwE3WHWR5mx+AzyYDAmvFeGKIbMEFkv6nx
CuyhHj9U+2RDLyfNf/c1xARnSe5q29XB8etjBek3vhyp7/cBHgaH0QWdXLGvofB9
n3nPF1pnQMA5Qox0DXY65iedfQtNcSV/w29tka9zRGvApwfjBZ9KGNHo/Kee5ErP
TlUc5ZT+lGindHN5tmD0K6PfyRiwUtBJYKsyUznVCNi21msFgwTJszwhaqjlsTEA
psJwDBgQCpY0qV7sSkzCfOJ7h7Ys+wXkvRypIRiI4/0IxA6LYyEo4IfonlqIXVb7
oDWdDnpg5OSa6WCsgNmXwwWYle2TfuqCbNb97U1l7iSNNZybUAOPYC5YhrhMYFxE
QRHA0Vgr72V0C4TVUsbBGAYpHJCenWYz9JwKe4BLehH5jZeCBOHkLtZn9dlO5683
70kxhLQDqZsHbnzyV9zyywSG8Sj1cuYLJpz2+q/GSlDDek8zDLuRdy3bjVzCgjWh
9iLC0nh708U1vbz6EPGBMz1DPwu7YS9tbDAnTn92+m0X9FWikyr2FP4fEsC3XWb7
2JMllOJIf9aE4DIL1EYND24SL6L8k6NbK8uWxnAy7Gis4/chcZKYoTRkDC7crx59
dWVRLEBslyatl3hoRqNUWIVGtVjCa2enqtZeEoeuNnlKubs3QJ3S2gpLcRP2u1dd
Bmj96IITSD9XDjA8cOFDxg==
`protect END_PROTECTED
