`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6LndpXTUdbXMJYYK/w6KJIVjJuD51iwSUXmILS+4lci/rKMT/Kla/gREVCQUDog
mWD4WtxrNLfv1T+V/u2Ath0LEUd9PoBduY6rBPpuuIZY9+aqzZr1hmV6D45KIIwr
zF2x7Ia2yjDsVs52eaZjKXx5xcKhO379mr9MXkjs3d2TlBwRD3j1KSPB0MyRLn77
jLX8FAPgj345je/xYSL2hBhj+So9xnszHXF/m2Zc/jmPlPnOT9iG8s3Yd2y+ER9K
RFlpvKGiZKV79RjKMtopvyQgFLdwa175AzvEOQ6uhqJvHbbQY6xKJ7jgETiVTgWS
qBGQ7l+C8G3EJepu14lSvFXbPNuXDLfQDL0rQIj6Z5qAr1afwSoL5Bg1Vmbd/tuv
/GBoWbEBroARelk/EizpGRi+4q2YwtY3rUBwb9AbhI2+HErIIYsYUE4rvO9Dgr89
PurNRsH62o47YuQP1d4c7arB01FxV5lGLqIEC9P7kAqFGFQW84Vhcfv5Iwx8Mr9z
r/6iV1DFeeEBhRkgQTluZ87PjwyGlmrhPP2VB+/7ucUC2/byeYcHZCqrsSF29DqV
903biJarZMlZSDGFlveVBo3saO5tArVfDE1XBubHmC6dMgV1/9uH6fbLeQSt8hXZ
2e55vchYrJz6OxaD6jAaKFjsEOmxWDVnztHouE9iLJbAxTKKj4ikE0hx4hmALqWW
ZDlOaamlCQxeawQPkT7ue+E0pxFxvMHD4iy2ry/mgmmIyfq1J4kL1QuyRuwz+hUv
xqTmu6v1sHOvvglnZnij1YZWn4+mqXVOl27TFIgbgphDt6AMDHCgk2LciHD744PW
jCC2k83AEOMHe1LxpzRi6ffAhzMvsmUvcNAiaNlQ2ik9wtSVmjdsEVo1bbxtMAcZ
n6FhJXZHGLggv7kFg/P8ow6j8RlPniRhLmR0AHXQKULaREBUJF+lhLmQ9ZcG4okW
G9tl6Av6MFGGU701ubn0NXmbfWXinTnpez/U64uuVYCuqIYTjCqwiZjNNPXhzP77
`protect END_PROTECTED
