`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vJYYKkOGXfsoSljsgqwcT6lyJgm9zNS41l4VFHgH1ev75KOIZL/JxVZ1POGIU9fp
jaEKqLeIwbIOeFE+VXTmjt6TqyQsuiONxGMMIYunKNAtfyhXuT5ST47qqNnHCHX2
+z15nvtC20Oh16vg4UCR/dUSKAo34IcutBSZsNWbwijk2+zJVSEwJjkYvkKzwQT8
uqP1Si0akVPwghlV746jn93zOSeJ1yHeCQXWG0r/V7uFOqn64rk3RyofnUrSt+Le
w7gAzjVmDwLDhEokzmOqYOimyDHgAnO0mHIII1h1BwV1BooMcseWaejwVAnEPUJP
oIOwPiBFjjoZf8l+ANWrrPRBgwjSTzDRO5zGs4snJC3i1zL9ObJmVwYE9W4fq/33
`protect END_PROTECTED
