`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWvk0zN1Q9Afz3/NKFIJYaL5I0Vl9OGrZR1C23RlYGO7joxipImjgLOX1WdpqrTg
gSO9RV/EQno55sfwmsvoipRYG9Uvft+gX0F5f7uRQsH5AKUfeJcTsYz8M1Vpl3uI
CLAKCiKlZW+lq0NjA+g93tSURcGnjQf/JWkQ13UaIw1XZhY/l2Q3AoGa20rNjnZw
mnPhvanL40fJ9FmPOW5gWwOWNqBuQ5WVsF5sxIy4pt8GSC32FOBYoUg4anP5E2tg
2NGPyWgC2JJmlecE63k7rnm7RcJX1jk39ZRsGk3BgXR6mbmGWMeMMyv1trb4HPPl
M7NxFne0L3A/Ryi715hDEJobpaHWjPUbiC4b0gWmsN9JfsUnVMq3IjMxh4L2X1h9
OeRwE3gtp/lZUKt8fxoCOQa9DhKGGbj9lVLQRP7hYFPtrGGkDuW830FpuvHA+Y3T
gos3RhlwVCd9rtUTwJsTYA==
`protect END_PROTECTED
