`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q3HQNkn0DwBsI7M6p6qEYAR1RIWVlPICN7TePkFwZz8Omg+3PcntDbPoMWk66FQp
JbPfIokLO3eu/1FfIlSCuOQEX7ahTHjb5tP5JXCGAPAmtne3ag6AqVt4gqMLG5oI
eOKApwAYuZ0udK7/xYX3opcPeZNy4hQMOlTq6x+y7Ll3qn/Nr+EuE4whVQA8Ci1P
X5vW5QbcIb5fsbc/X78JN5yoXevDYkaAQM4E9WbNh4IhC8xfQUgeq4ElwEVEEwsF
rwacHDndIG1H9uCxQyBFLzcD3fmruimeDOP6lOr3HMHkBrHy14QXkzuoqaje30Yk
mHlYMbMQENbeCeR9zksAsrtb/x3f4kgxvlYsDL46ITfXFMdUN1eMBZWp9VapO/79
qv4IVsiPS5z6tNksrZw5cNzuSKNZi/ACVubrHx3HUfb6gSr9DvT8F3fEx+fHiaL0
EgMza1SqFFMJDUNecexBMzgVvcxl+/P0VJjKImdotJ3hPjgKl3xm0o/MGX/z2t4M
OnvN62+zHzUvi0VJWc7fKFbaUTFNK5H4QCRdwqkoLl0RtlIiSqYp0AUqydQujlsy
Z5WW7beFiVViAlaxEh0dHTMDAaOYV37Y/oX6KHa3tEw14Sk4F06NSb7amNFwdC0V
B+LR2d6OOhaf9pvD1TjGwxGVINXY9K06y5thhC7en1EV+jx/fC99j9TYT1Xof6Kz
faBWEuRA1bm5ji6iICUMxv4tAVyqCszifGY/r+dJz0EHyXjM/wCZzk3BvUkiCYEP
bhTYdRMEi+FA/IIQE0yn8iIQ4IyH/DyJV/qI0u3OvZsePzRbMl0h7jRkQjFYGQjN
Jh5qW6U1IfNBh+qio8EMnbYuDh8vBcMJJlRoqpuvae7YaaGy3XYDfjF7zK7eRofx
+5lOFzS6UODmISSjC5g4e3kIjnbwRWpLCdSV0KowCiuAy3gNipFVr6ebb/RFW1/f
nEeP1R7i6lmAhw2/GGrQL9sVajP6lJSlZSECSMj2x+RoHFTsiPmjSGptHUiW1G2Y
6q+6kXOXCAIjRgKY6l/nSi7Tnd9/IaPBRfTKWVlV09eHFJ79Wgi+32Y9AEODgouN
X1IBAG0NFVQQbo03Pyp8lZlZZlVBQ4R8a37O3TI7iUMmpxhTCOdbLJ3xicIX+1+i
8kaY9R54nhW/xTEO875lIb7HhmXb8T+q5I60RN7zMgBQnwUajOZmxP4x+4aNp/Xk
HIN45jJ4TRtZNXGmpVBC3MgBffNDf+djCaKZbcsOpAEZJREyhdviQbvlSWYgVPqM
rcnPjfyDac6qaDAqWFOnCtg1Y/fWBdLN2KP/fh3tDmk0VAvyYy9SQq0LLkDfAe0j
L2fNLv/PBLlyPSYfOm23rW5L1lOme1bKdwB4J2WNdtdY2osFC386RFv0K1hiH9hc
lrXlnpTprio3rCGy2kveqqXUq9taXUQk3fE3LN4/rMfaTcloUnOCe/NKZAzTDabs
x/LB+tu58zcmsBjvEfFnrkpGzl5+m0DcLDxvGh0b+B1DY3kToFpzDpVUOMcB8cxZ
sojostcgouh9MZWxJrTfQyij2n8l6pQ5d/X7CXAOrosqDptZS7AvAjJCmWQs7ibh
Nim98qCj7saz/KAppHiA1bZaE3RwJcEMIv1SpDtXUfimWruXfoNucBxY6pz+I38i
F4RaBOLO6ktxE2vnbIIFXBnUPUu/cMr/A/z6/cE1nw5JKSglHmze8DGW36BaKGpv
5gafpRfFkZIGGsTfjb7hqpGY8XjhEKRwUNBVOYmbVt+hG7plaJ4jshif78lidKQf
HkpM4WtZdwxKXHoyAKUHV0RXQZTVyGnC9gn08Yy5Zt2K6cRGXlYeLgqFxNxs4OWD
+nCKN4N6oYk8AbjSU2T/A9EfDbwsH+DJRgUjTE5MplzeYCVTG0gAZocUNI5Frszf
kKaKKrIHWCJJremyTXHCJ/Nv4XOPLuJIDVbIjdNgyK3go9XUKf1yncM0FV3pAMfT
8Myr+Z1UB2uBYFgyEjzdzbwaQZp009VrnJf/hMWYdDf4W2ijCdRGXZjnFMs4fgB4
3MfIFDCg/CznhZlze+3KWD69sOA/Fpkl/Jo+Ut/GcfzG4pEMIXPb0g4xYpNHYB2G
9sHfZASaL43ECfZs3+Pro5B5dKEmCIpQSO+xbm6AUnBmZ2A35Y4FlhtVE8GD8RgQ
`protect END_PROTECTED
