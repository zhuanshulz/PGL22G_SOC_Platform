`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
REnfbA6ehADdS2u7QMaZ3iUnD6s6zNqflF5TlXSdJnWU0P3hcSdy48CAzHltMAey
ZLF3cSG0pcFUV6VGLEg/MulgijkZAKYH/JEsOnsw76ahj1wu0VB4oasVJNjy+ICq
VWAOYT6o1rQVCRIxIaLw0rNppgb5B3YSFaKAPdUyEvI4OKsC7ZFAluQG8iyvOq8r
qRn8hOa5EhrOjdIOnpe/x91HVvqNgGanx1QfdP7/LS8ThkRFxymh9cSW02YJrcBb
ZnW8qPFN0WLX7x9iRKwva2TnrVzTQckKTf7X7g2uMmG7iQJrdi4IpozhOGo9bAkb
zO3NZSgH8JgLiF9TSkiZlz2i3SbGxUAK8xWQRJ9YsxHxKOLHOFxV58dZRY+7sBOs
KVYLHFvjAlsd5oDW585rUR6tzuan2tR7Qdy43rX28rlYv6UmizesMQxxNWlruyyQ
UhpFfauAk7TUiraM9T8rfMt2elkzx8bbAzNsuhkDDlvFbnVIONKid1d6wR0ce2nn
2yHlDE1RfjAk3bb0M1Zu6Qvinid1cQA/DBxmb73hjz10nd/Ac/2blkOdHMXVHBV6
PrcjWx1wLMKLg/8YlmRWOUubpfOoElHOG4AGH0mB3pJWwqAdaP2kc8UpKPeRdADO
8fcoKr5CICX57662wbQPJzyaQgYChus5UyZJyyKGAcrfDWH5R6AP5Uq+W+UXRXma
YKsrvzFA5yrQlTiWsJRootbh08LVlmeC8PTWfcDT7Rb+PHsT/4sYzAgyw//I/Jfr
VJ1LkaX5u1FcCT2Uxf98vukLCGCBfedMv7/SSAmQWbGULQOyZFP9w7fY9Lm2c8T4
RHWhlYTeiYyS5ZsWqMzW6HjGmAXfTUGkIRQOWLPUN5DstIeJ7tPap1+pCwtSZetQ
djW70kGe15Xgnj7LiyWBGbZ/uYn/wX+FLB1b9NSlbtVZKTrGV/PLE8hI+DT2E4Wl
Xn0snYpFY9E5YR4lKt90sW7lTavAgdzaqSBRBd5hWnV3pQjlPo45tfE/TVwovKSe
K+La2ciDbjKkKiBRZIci6at2lLTpAsSOrEtUh+RnoE80LsLMTgEkm/8WExGfPowr
bXwLAcS5A86psYubAOUIlmK2zH6QE+qmlBn6HAurGFx/r3N4D/k6iOf+/S1SUYyw
cWgo86J90jL3iYvqD7chSd4xWuS/LzevvTZ6Ph8VDOew1lusQzG8K+heEsuD+rVp
zKaXqYGMvwBctT8WYUOUDnDOCy/XvqZASoI6UN0QS05McuJFL1w/UuRaCq2YC/9b
CUjwiMKtTFoJDXSTEBZjsasi3ubwMJlr4oE7ilts5lMqy+DxKbWHm+2AETAiMAs3
OeNGTpggsi3B/xNCpm5UIwjoYxYLv3apupqjR+BMN95cXI4Xe8D2W7af8UKd6Rk/
uJ6uBFi2iAWa8+mYox2kB41o+tixSpUK3R6hzUAtsT3XW9MxdpOtbgP5vaQv/abl
zVPg+3FHY9JCRig3QEhFYcDBL+LFcrYsCwFW2Zttc6XlSma2Uc11SrZ5XIOUYOWe
SzACL+u+dKgmXVBj3wVg/fMKhmekgtKvU1jTxgXEfvLm1j0Mg9SmMztziHJFWmRv
L9i24ydh4GwZYIDNkZIvDjWOoq+PKmLLlV7N6OQAeO6491bijPD2pkszHzoJcUxn
T9HgPOwvP+W0PFr/aLtha4VQDsvLy36QQRNYQeWPpfAsgsTv4Km8MxG72aU1UJlP
ylQqQb/3FY8j1ieCARHbI9GDKtL0l9mNJoobS14enNHJK63wCPKvMJHCit0uqf5H
`protect END_PROTECTED
