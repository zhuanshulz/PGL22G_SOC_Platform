`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ep/v8Luw8XNZ5zvAgHw8Rj8sp19QJ0ZqHZ9Bv1W+IWDzvhJ8ziEKpWnKWgDoxYyE
OIF+emwWGaMfJ14nm8rsDOu6wAx7w3lixUwLeJPbxlgP8Th+gvZy0eafZ2oGnSfG
U1ZKu1EBJ/STbRQHpDp1B7gEoDMD2LmLcF5jrwjovAPuY0nFB+HHHBWs+cdqS/D9
ioDWJcck2dbUPVE9MNjRie5lcROIEIsS4rzcZm+vlEj0eC/K0ayuMD+xxdGF6sOm
Wry9G/rreofkeUdbZO+UXKeM2eiQaeAbikob0lLOlL/U3oAImxAtlBBLaeCXzuMg
asXoxHEO+BIFdHycaWdD8O6sZJYR/8lRKyAs1HRiyDLZ4fslH9hRfuX467OP+g3a
9B2cFP1eAvP4R8HAHTEc2YUxTlKvljEC2pTWHzUKr+1Uv+h+ciNMwX1Bh/G3vrHu
1HvOxm5I+/KjPG9ih6xwHJNXU2fO3HBnJXDBwwJLU2jekS+jcGf546YrSVqJA4Er
CjhrsyeEjX22YTQsBeWHI03fyvJ+uNsbROS286cKVvxpxlEVc94Ws0GM/9/dvybL
y0fxj2X/A4T78O2zeQlvssVMAiRhn6RHvaf3HAHgangw1qY0QKanvoteldX5hjVZ
LslO5tSjUTKTwHSlE7Kiuw==
`protect END_PROTECTED
