`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvFtvcGlXRNc1/gIHbZjrviJOb1EVhrKijE2c6YfFM4ilqbk3iG4e3NS8SWDYpGd
WNWsUacRE2/61Bx5XfBAabcaGLXO0sLJBxJQeqUuBkvZFp1fzF7Im1gDs/o96Mf+
1zJOdMWnLxEtrYQtM/ewyZbALSpwiIs/k42YM3T8eKgbmyZTWPq4NL6iPs5r4H1R
TY8bu1CRaj1fD+Rw/IV5BOteq8hBdq7Q0zTzfZoFEwSIJ/bTAKEFNBKNU8USP0j3
rhgsNF98kQuGrRlwfc+ziUBdrDpXqpXRygisvVKeXM/Qj2C3PGM4jMWP2aIYuuYF
yzPrga0S/vtCHHPzbRD0Nn13TS+gkqtYmLmuYN2/xcZ4n9YRYJFcbkuwVjdpCu2z
H/VkfJChENQW5p7irJKqpZaE3863NxPFUHpKIfaXqXabpLPp7AXbVM1J2ZYzkz7b
kZG/Q2VbYpfaKmA6W0JO3JuANPP6qSncNtWHcxK5iVqe1zKYXJiBD69lG4S32I72
/6f8wGDv3BXWBYZBTfAyhaKINYdmg5BSLyP4PrGDXWR5UBBi0Fq8U3Tz8mdz4P4/
xkZp7LST8qxoZpktrOPqdPHzI2v1eu/eSR2nI/EqPy7Rfm+HMeqw+Wu5JKWvufC0
luDoPZtx2jWvxnznXFI2Ewejs2zooDniRo/9oaLC15ko7tU7ynGKMOooCffjbfrF
dbyMYacLquSTnBD49QcbK+kijWCmBO9ruhjtuWc7PKj3G02ZaanzciOQ1lPCfCyL
0E3cpY4CU+uvI7UCc8ZyAnA4ZY0MOdP4uZu/9ntm86V78ETGTsEaINfWWN8dMcx4
r4PVvfLjYpXAJxoDq/fu22DxXcRGsw6T0XeNzu+P7KHka44WL48MDdwEhbhGi6kj
dhQ2e6L1UQh+7L290N+2+XN3FlUK7bk1GP57r69/HiEE8QwFTOoP6VtRfYgOeh9z
aoNTq6Wb6NTrSVSj0qZh4cpJq49P0yP9+Qmyecghk6q9ORYqvXiKbIbVcwCZyLld
FQeZ5Ac4HfDYzzp0iBVtlS8onvN6miprxz5fGRdsyFESkKZPHKhSuT/KqIfuznYN
qe/LM0UyV2Kq3dYFAafbYry/1NGrCpcFoM3suSvWsEkX+qcI4/Y+u5tLZX7WJ39R
DTJGQAiJqt3hq0RpP/FLssHiG5DZnP5h3DtU7dCGHOTaVMepsZLhX5x3G9QUsjPg
fjAXPAk8zPP2QVpnaKVga0MEv02hGVFm1UjrKG04Omq310VlY0RJ4p8yfUP8CF4s
qQjrzdH8/gM24PJ8sSyXnZ+JC8HtZLsULAJSceLqYSXVJRixknSRviqHVy+z6YCA
Eekb7M+XqiySFMsojs4LyzoRhSBCD+qNEYud85VL2jIi+5jNE7hUZ+rKY9sK4gwf
4HRsVsPzTcZlpMNBhyC+GpEnbV/2IyeTfrAi7Mb6xljHz7+dPKHXS2Ykrq032Rgm
oTMxyhjkPLObjXrXZXnhV9/MyF03t7wbJnRkJIuLTl4yuJ9Nv/vthvTQKe3FNDLQ
RXTgY7ataEG4Ai3SH3pW9tDIVSwQSNV23walYV2RfgIhx9NuUD0Lau7imkUPPDmD
yqjaaQ8UtMEqlfplmGtp3EpNDvi3Uwr+7ND4mJcE75jpxsfg2F6toBCIasnZ4JXd
8lYFrutKB1+reu+IE7pUcjjraObi2oJRUCAaVj1kx3I0bQKdA7cNsqIVzmvmFhAr
FrADeY8m+QTy8ZFDtHJiaJHkaf+/uo+6ZT6KxD/fQY+eeEL84kgHgcQ+DdPYlPe6
JPhn5JwbpYIeFtCfCwC5KGaNw0vp/8YA0KC4r2JfSGXeodKInKerGCRam2OmJjzN
wsuQFNiLLQW5kbfTIDv01pAUHmQmvvB6NmrUpvihwb0abxPm50Kd+536QVsIr3U7
eLpI31+Hm7Do0tl3xWis46aKiqZjv0DVX6w4ufG2pX3rrgt3ctfEicpGqz0bDBMv
Y3F03TPPlL8F74Tn5Rqz/5qZ31IRnM2bLYkEUVaotZQN+Ck5V7Sn3BeCpw4w9Bm/
rnQXKYwV8wVO7ruWVr6uUanbt+yuL8HzPhLP8O8mzAUNG5wJwCiRK5uduNF6DK74
lLfzl1dXOzGvMYwr/hTcAw==
`protect END_PROTECTED
