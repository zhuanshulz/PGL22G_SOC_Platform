`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZAGOlbS1+FOVBxmpBLlIEk32zi8gLpP53bHP/gYooN1o4GZYwN59N8OUN6+nz1m
TMFSWStFCDRr1iAEDeXqqopo6ynB+8yEaL1o8PBSrAbQ0WPPUfUy4d4bafR5KVig
JDDCPrTOf1XGe+veA/LjK+nMlXsT1rMSsQtslL/4r32YFxBo7dFFAvRbFKMWrSRI
j3StvPwHIWgaXGipMvzXKRZaQ+5JSdLvi3QnyzUpKMB6QF9pPGR02ArXV/JWXjP7
kg714ZMMzVEMlCGU2sDc+mIdQgnttKk/ME0BEwqn/ORTSH//raB7t+vwTvrZa0Zo
c/OzDv8DX/pmywPdmqhM6W5tUvWfqiStwEapuzRGy61SdoXl32s+VXYU/pjqPFe/
J7PANAGMsnkbgIs6q6gFYvUZ4rF86tSsnnFL11d9HCvF7Gi8yRC0i/d5qXUSpdOK
+KmXDREaQzAqcrFJOFHElvt9xKLgWfdvcrxKsyX3oDJKKVDIsNBemvdMi8PSU/0+
TVxCCrbgTweH4NxJpIBueug0hYMvNr+w2LGBtWsN1aFeJX9kvoX+hZ3PYjwUnLCZ
wI5DtUG/C/NS7ER15rsnX60CXngzkPPotqg0KBan9nqixaFa6Jla/lGEZekz+Mqc
BONvLLIOFCaUDENhDt6jA5Mmb8sZb1LbpijbwvjgtM9plgcUJJYyudG1PuMZiftt
6YuKN0LIA3620lvWbCG/vf9ooV6cOVs2BaqUt8FWpWkfju2G+4Ypk7WK6jv4xMYU
GhMi9wX+o6siQ1tpxGb61zvibe6k1yoHENULBxhHtwWFtqn0qakW8QwBDW3esNB3
wTm4n1kJJP+lPo0heVGAbW3jrUgO7GM6EUxtjENnLW5t5wZc/unhCt4GVQw5Ulnh
Of2wqmzVPzQWrKnJj57JvMdpOCn6ud1HeAMXnn7GxKc1YaBJxFR9qI0l77iMfpk7
Bsj8HsUj3h96h8fi56/RVh0rkuKhUKthLWLX+69MX8wP61FNfJgt62G1eeTnvx55
4kzRwiwJN7C17dX6CjUBFaJYnFQlqNvmTzccBbArDp8XKPhQf1zMgNOTp3wZGEqw
W6uoPUgBgU3U5jtzt2xemKEiAnor9eiQqjxnS/PhN/rayYfhf+c8QHx2n0uvJ8NX
B7JMNBaIDiSxHWTXhYnx/E5MMIXIDYAbnFiwj65g1dKe+wkczX+aWAfXMICeTxMj
/WKP/oVuKFW7aVF12otVe3nN/CtGP6HMWa7mchpxhmaqal1ZgPjIFlX3qEpq1xWV
gvKzsvHir4pOQ4KyKlQPdJ/CvaMqhjt94UaaHp9laiE574jdS4XVfCo1ZZ1kNk1t
LbsZUmlT8xnxLOU7AZNyKa7TjzD0m+wKvoxb+0o62UHOR2CAxvEth2XWWvUGMbxV
Pp4nDqrIu+ONeilyO0wY3b3QNZKsRamfXVcmcKaaX1AgmFmkz+2hGDLxu/56elCX
sm2iuSQB5Xvq+T6hRGOME/n4U9mhWJxEauoIPrQgADJuFHqQERseygcLnEJ0K5jK
UhJpqVwoo1ZB2o+rNPohB6q7NK7c1YxAxzoc4d8Bafq6TJiI8OZQAYtP67Yxgz5n
MI16qTEWZHQAdGZA3hlhSc/zF3AzUSCKe5AGcOPubnbS4Urp4lN4s/NELcT0hV10
ia5tOaVnKD76HhrZP0j7QfeFbMTF+KbujqsMEUFY3uxx6YBsnZVxXVt9xYj6OmZy
sETcBdvK8efyyESkmC4B8h1kysXwHgx3KGy3b46WjNHXLzA7bkjJP4fbFEQ39CoQ
YMty5l4fvXI0hW7enzXl4uEVMmLj2jE+uqjalLhUcA1TenPKWhSG/JP8E/lxOmft
R+ccx1xj9NT9CCz4rHEZc7OBUkEUIth1+Wh0+nNIUvEEJsw5RamGgQeq45aDz4Jx
X9lAXN/P2wYpfc6PMuzZ+S48ufoV8l0hBEiQW/hxqPdJSZIb7e6tCAiQgYNPZ0Jl
Icm24VsC1kQ5veAqJGcK9eD/S/nke7KUeu+lwJvRm7SjejWJzBPqGkwNlVqPfCzH
RM5nb+DeVbMA5RYyM+Ow+aIsaG+upFUdY5V9suQAT+O4rKnSrQQvpnQ/hbQoiOLu
VVZTY3X3Yh+N2DrNT75NonzlzDbvE6lUTxSsz34NY3qfO9FtEbF/K3FpiWOXpjV/
OCnRolnip0jOlCkBVxOoN++N0hGnnNK19Gvb1vl09jV1vpABuS/3KtTP34EJzz8q
bXpQF7xaPP2ug5cdQ8C2BYnT8mmudacl/uSkRmyCqTOl9d5e2RQ0NKmhrEau7yow
+XF97fiZW4HLrvJsaPTS3SWy/3tff3K4RAkPqER/svi9jLTgvGpXsusZLYskqFwk
a7bmp7ID7J3pRfBVzjI084hzEmYhq1Ts/xW2icV9tUhin4NQi+N0r7itPgvwmN6a
FQnFq7D1415f9yXAz2o96Tl6dyO3UOG4nbNAYR5a3TiyEZsT1+IacjQ1U4NGRtZW
RGKb/b0LIKesNRxJgxwleBV488savWBjQVxArxAfVgTl5w//Ra9bYhp+Ecs94vt5
UYzIdso00k16ylNAphf+AwJxsiL0dWxp7Qs3vhUNcsuE8b8Xo0IXJF+rMjm432mr
DFagTEK1qnb5OUqaCKwV8HXOJGZnqTXPB2p51DAMveQe5aMThRnKZk9K4iu4xZ8Q
5Y5J+9sTj12ldpvKn/FZX+Nifid3IfZ1MikD+jP2jV0iJxUkn574aj4QaIqHvetx
LoKpphO3v/HdLXoJp+jp3TF8+629P/7SXKvZhh+ct+ogBysLIIH1s7wNwDqZVWG/
jpnIxIwqRUYjWd1puzppuFdh3dcTXYQuA64I/en8IcsqtFZjYMq9wD+AQlW1l0Ez
`protect END_PROTECTED
