`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgMisrJSvpnVm+ZtFbViHmMDi3LB953YxG/anLeq4Ea9z83Wss47+zaMWlObBAI7
3TjTqLMCRe9/2wtGlkD0YNw6M7/4Udp0aE8gpHnXf5TxIAgKH7T13vCYj5Y+RghX
nnM5qMWce1RIJs8+KurTrEckTJjRUIbhgy2Y3WWSSe7LlCrIE9dhpgiNSCDGRodS
GzSv7u4eEpdvVpAyucafiKqpNEEU1TZb1RMkFTVUDCZvpj26j9f51F/YMlys8J8P
Afdn728IXPME0GjMRTLqpm5r0x8HaRxmiqNbbdEWJ7rc5sJ0jXLcL5zHHgcZptZJ
yPi6EIGduJHymYkTkfmyOKxQAC3mVAHJfUV2gRjpdadulIqvwtCt9c1yJ0HB0Y1T
7hhs79lO7TcMA6JNTWwLyTujW8SNCkGVvYTt/EqEgL8TMjh+DPEpvvIjCZlzbD8H
LILGS3EUmSs9ASHUKDWkzzF8qZldWoiaGH6L1KlT6qImGz3z0nWEbA5ZAGeh58iu
18W2ovj0qNtHd6Bpm/KDNBBwAweJcDAIICJShZP6m0AH46TO6PCh2+HzXF3V4SB0
zTAk5oMElAlXMdX4S4Pg10RT+1zOySEeJTRGk5LW1MiqNHh9zq1ktxe4u9q+RS8y
s/SYcAPD6zFqvInXawDAA9FhhmscZqq46YFt/68tM4LzTGHU+H6u7uZXM1JtetWz
DS1wOsLLWo1wKQemMH5QsW2QAm/sVyFLzxyH/6yy+Pz4N2goBDMoMs4t8W/TKXVX
+l33ubVp0dfAlp/zxpQJ2YnG50PWq9rAe3U1Bk/RK0uzqgG5KZrYeZjT7uqPJaKy
Daby9YLwhYRRv3R5w04JV29ttCzLyNKUqASfifR3z5Xh9Vb0xPXNDa0zVrNkaDRe
s3Oz26EcYUEG+4hTFIxEM8D+Bi5NMXiOiDJUjQ3dvhriIuf2RGX4OwklXVVK7fDi
RwEULVUe0czVSNnr6rVB+BScRfczT9ljsS6rFwAoUX0rZ++f8j7x8faNHZtmouje
USFBgKZJN9O+fFUagygaTollMaq2f0wopURxOrQiY/FPd2JkBojjlygHJpH1KgtY
JSVwIllIBOdyoxs14VO+83FZtoo18Zk6SvUxaHmykq2cytSZKiuf0BOmi2KOwpB1
jcjUTDZJIh2Uql3ObRQGSO1Ww26vHng3P2818+3QGFVPc/hf0mLyM50RpqE+j+/Y
L+gKfTtnBOiAYBLICYgMazycGlvOJO6maRMA3lJbVfSsSypfMpzYp3wV9KiPKpKS
fC5hDSDahCifqBveDROGzBQfqyjyNxsxVK8YP8rsmcrNVoX+5K8I0tOiUdUbVLCI
HNSywYdCfbk6cOtxIXCqqhv9viNwxwgQHSS7DazYlVDxjOngp/e/8nTtrRoD3+hY
m+slq2TL4283tVeXCqXC5+rGuJkHh+P9qI2uRj3a7J5ZqDnPrqKM8vvehhHQcKPW
1QdqxOOTZUZdwh2rK8yjH2PCiEsEjmN/Lolv1zbAEp/827gvEiRv9SYpXKl78KSm
9GYsVGwpz/fsbhYIkuNlj/bOw+++J4Hs3xnkT/PZYNznZyp4aJmeiR6x8ttayQMT
8vVXQRXtg5XKec0Lw2z00G0rfatMuEqFBUw8jW/bKuQlktX+4HMq2R7btHuNG0Dm
vwbYAZ4U9LUnT3jizYD1y4+NBwsnMxAUSVhPgItv4HOdRgrVSlENr9akPwp8flWx
4+pRVMOLuHKf7ceBQiVL0Fc8dy68l4e6+PSpsvaOMs+K6mWncnxIybPU3arg9Ca3
8d6f4eg9Ix5fYioEyjEPvRQCIylPJMkHkPy7Gu8fJgnkLzRjmz/DkgbC0OUPR1v+
h2cCeAEd3k7puWNfIRvFEt55L4s+zGcztadZOQ09vlHahDv2R9PAEuhbKtt/3SBW
5dE+ujikTzmzRFX5PqCmN8wpxoq+wpS3rsih8in5Gqqb71apom39lBagNCVil4JY
PGXCHpN30Y4sCEDbfZDkuCLOCHCGy4189mWR0aBgCvFCPOeExXU9w11AKhiB3gLB
VuCTjLT9t13DSg5RoIVrCTlvt1WzKz8kdjamTtCLaLltkbIXmFuom6W5MaXf3jfo
pOZHZ6lXk1h6apF+24ymp1j/tjhCTdkhHqkCO/HHk6c4EqkLjvVf3dWTWiVMVUNF
hqlTzG/yrXR/LULfwg9uFxxqhMyrurJ7awlMBZL0vZQMv1B+jcWO4agooyfEZjRP
68bv8Nm2vqQOfL/ELLCN8dV0Coa9PVkffY4L34Db5l2pK9YlKRuLuFeAcjyO9rVN
kIcGJlWksGw3pfwBYL5LMICfj+VBTZbmS9gtPrJ4vqxAWYmZi2G17y31XaksY+6H
xxZ3n5B5jOpAyRFRwqhUkwPC5516pZ7mKi4OZGRb4w6Sev/AQ4OCEv6Hva8LQ532
VcRFqq6Cjr67aWSavSzDbR2My1IFH6wVGevUm6sA7TtqdWI5SRUeOU6BOCfeHXsE
sG1PPmt5YrFEGs0RP4FotPcCATzhdWIEcY3xppqp95Ohu3DcCpd5EwADREGzjr9/
0HJ4yGEsMrjk2wY5VbXt/+wM+hxsnthCveKoP7N9neg9RMS5oXuhndxMHJrYYzqD
Q3HY2MnkvP+tCILaE9OccvnS6MI184DhZrVz96I2Uogvtrf9uXIEpPXy3WBYAq8d
mfmGMH/u4yf8giwdvLqT8fz1tUeXSLcF8+4UFv8rV9dlFI2GL7sm4zugVpu1t7UK
J62KviQWc87JBy//OdUjv1rwWyufT6yu8ZDmXNZS2q+BuUNTvB+ZNgCkZJ0N9IxT
As2t9XZT7aphVOe/afAVnzLSce6kGoTiKJpXPMTU27BZweXKqJsuP37X3Q2dY7DH
FAHEsWAeuiLTlgmcnz+al6fsiYKLX9jesciiTqzHlnKJw2y69J2ltNaZt8Jm6zWD
PAx4Y0SpFWoJcOR8jmSI+B9BF5zSsYJl6poEFJU1TlsMAaapxMEKwaLbror36jZN
ny3MfNSY5afO0qsUR4QFZVlCxF+N/pOGhWWUxwKpyzRW8TG61mVM+7W/vmXNT4tn
vzyNxsQfmAMdMs9YSnGz2lH7/N2tcsufdIlY6+z5LjwCfg6NOwOTVNOJmTJcO4dF
mJ0+YSMFnCMBnxWwWH7wh1kObV006U9fxvVqWJ9d1TCyDVNz459hqduSvw93clDc
9mG/jwnC4GczLOWG6u49EW5QtiylxlmITW9qzroUNXBHtV+uYtJN3VZ7Bc7k+axO
fHa7jDgLsGEZlp5Np0Whu4ZPlSb6qjTgNk2/s/jIK76tbciPc3HfEIo1Wd8vOcbC
u1Twcm11wb/KAB9nlySq/EtXptzICWa8+NMFKPl5wOE6aAdMSzoOhW+rIuUqEfgq
2t+No3jhuGeAFn+u1lVSkEUOMxlxuF66h6Xea509/S7qMRz14DTS90qjgl6fMtro
1k18Yesw2zvew358pSrKYo/AT2e5s8I4O5dFJP8yJrvHSlKwkeuGYfivsudtioOf
jC87aYLxW1iFn47h5xxso28BqtQOXZvt5QRV84Oo502rAVFl8fqdooNEaR9+AGCB
twna5u7vQnQSIxEHDhH9Ie1fLbDgTwRnUhE1EHTmx9yBzPE+7LkK1CzUafqzSwVq
J0BfWj97QOXF63B86sftMEnSuTNfUE+00S+JQRKU0l2RoFlYafROIVFHGrr6v/NZ
GdvrpaDkRU4PC6BuEx/g5g2uG6yuiPl9kwj4pG1gspFLl4Gw8xPsW1HaC2M9SXDa
sNeU8sUSaZR21y4dZig6/9yRIbV7BFbPlpiiNV18kDY3vTC7/fKV7huxPec/sf4k
AlXjhkgR5/6SxRBS9x6Apn3G261qFKIdcnsRiDfXtlTQGRXpSMQ0byht2Dypns7Z
H2twyjLVdbSIfum69X3KXsunyvN/sChLyAjM4bzOIeJvrVbd7+rP19g63CTRwkmM
KNJIyO0NymIaMAbmGezUSWdThfpPeBoSlGoYX2Bb7PaRBMRRW5WPT8gk8QZikoud
1aPM1Pi5Qo9NjJCk1DV/+X4VZq7xkEpxpOZJShbrnzYuezdl85asbMcQHeWVmmFo
qoM9QBlOhMfnUIlzMSxnFGW7FHGgiDklFhOuJ0KGmFpx+0h3i7bPz8YDqfSaHUSr
j7QFoBCDJBNRMlI+k1BsZdm5GajNxm+Cab19iqW2+qxGJ3ymIn6aV9NNSr3v3N81
8lRplO1869G6Q44zdmLDQS2p/FRxrSEXL8R5EuOyxfi4gDPY+upC6ZMy/dQIz84M
puC+wvXwY3cEO+APSTgyueyzoIJFuF7vv994t3N4Ej4qQ9Ylhr+ytJQeBM+ZVgtr
tLhqiTL3H/hXt+169j0dcTsm4nt8eFclVKMXPGuW9WjZHY/kdoYnIVWYU/+U3RUV
84Mzv7PlQEH3RBxKcKbyrpk/Rr77nPAGaNIWMOIMQH5wQ0aAj0vqf48+hiZzChcV
9hipFeT5lVqmm1yrAauUMJMIAkzSU17hDmCaye3xwhkjAoZPQOa4Adx2SFmnGalf
qugD22MfNr3zVe37xT/R0ZppHilGFUOt7U285YfnRk7kTmP4Y3OaEnjRTS4ZwZkY
Q8o5VxA+lsO4kyf5TWd5MEcfLEdrUQzOxMbwARz3If2Q9JoMIyL/jbwTnZXD4QgL
hzp3um5fyjAc/SrZLBzbEfqlv4E7ZK5OhjWRI00n6EwSQD21O31IGUjoqfmWutPK
unfIuq3QK4A86lJAqc92NqviyvSBZkkAlETKUv8jN+yoV3MkJtGpQjwTjZp5320E
YgwMtVBoRTSNPneqZNXXSltneVKK/xHvejNnPsonFUnLYz4IWXLFgPZgzMEpPu/2
B1e5UecZfclg2gYDFsN3c/8kbGG7QEqzhsfxsZwB7BRi9kketiItCWzAQfJcX+87
O5hQRaAmL17XjQbfjvs57Q63kPNiHbyiLLOMPxlcrjSgKoweNwTOXG1gGewV6LTW
5Lp+aFk8MjGmfVPJnvZF1cs9gSbFaahuFRY9hlpQVICVQoBoATkCC7eSp2nBpRIr
PGIZs6Y9nKW0TagqMvRWcboWThwUA7FBLHQz8A838UJPJ5Tq+v3V2faW81+qco/h
nYYhPkOeAketfa5eEmXydJi01YI0QdfYDtVcP/seD79Hn9U1Zy7vhTqutpDENdSb
Aud8b5O6CkQBCpmLXKSSu0odemuyrAZzdVLRRJerGsqAlSftfrNcsw5YIYMOgJgy
RrsXIazcU3nRmzOsiqoKsovOIFpK6090LFZB0xQeYL1An9HQ/7ibKzuSyrDrF2qI
cip9qYwiEeBIEJdXFMBYRClGwCu2UXdmarOeDfJWjgygOHwmoREPsHcn+jBu6PnY
HuoNJnm62IkPKhB4o2l6zlO/qVRl2jYCjBIEmrwmgrYU2eqeSGlb65wcfbyVt9qg
WZLd7k5I4KVaK73gVIXUIu0r5BcSK4v5/3xyL8d76hSC4XmiUo0LAuPme9G9YTa3
WCPa0m8hxakVrN31pXieGDM+5Z81anoEEqmd1S1M/84vZpuHdrUrMLa4eUFC6gcr
+2Y9hP67adeYKLqLAaabDSccvmGGrn+Dmja3Kl4X4JhukF44I2PXj+1XYu6HMka5
S0n81nCGm86HizmgubcgTaLxof495v78b/cfW8JM8paXNUd1TVYPp2ljhrRlgW+T
wZF1228CBpggvDJBQLQ6jDerMtqiAxDHtWJ9EsoiEa9eMOO+j/0TJRyajJAqydo0
0OQJVAni5DTuFgbKM+W++dWQ3SHTfG/nDb1y03W4QuC/780rp6M9+wiAXPWDMzv2
A8vGRjizm8rHZUWFdic56cEILXNNHOANgLK9jRGeIWRuA9LiXIApqu02ReWtELGd
3eLF7Ly62Z91J95IsICmTweLe6IUEsP0Yb/27v9Ju423rWWvbrR8tSDJmoXkJ6jy
UNyIpWhlcqqn183MXEhMmXnfbi2pyYreYBlaEXeonFmpaqMsydq/hAUoxb/r39AF
xwVvWkhCYEemDgGTJ+CWQ4IWKmPNWpz9mDNGUJx7ZUrmBNkJT7ilJb07VvFegQ2j
dtJXUs/vIdqiue2vMO5/QsmMcUFZI8FNQy7hVvCKrWKpgeUPn1S2SGO+lTHHsqI5
1YfbqiAh/RgvTnNHwNunaxneQDbQRHX2dvF47xeDsIRuTczRJWqEdTSR1/hrRkhG
ln7ylKOkmd9VI1EsK7ildYtqY6rWR34UGtbhUZdb3bYxIjbzIa7qLgae2BD+kJOH
qSmWhVqZdOKX7Rupd34X8nIVuasIlbmNClYLvqt9bjZSogonhbiWjkXTM8bv3gmU
SyE5HOoAFKq8K7MOtkGs13ZoV8aShb/jWfJWylUfv+/UBvqJqt6DdJZ/NgzUz27K
dZGSP/fl2gYfPUXOD1nnJ778hrdCMIhXOiiNHngoKsH7KohKnqOH/fZGFHHztyfC
AeEcBc6ZPMuLEWJ/qLDeVpKjikZavzb1cgM2NS2E74q+J08otKzYFCL9/TYJXxhj
c9j3EAPPcR7Xv9c4SyG9MSaIRrXpwHIs8Y0t+5hFVmq8UuUZborgAPKCcr8JsiWU
DvPp4FJi0KMYWf4h97Zmmfvnj8e3pQENne6qkP5OBGN1TnTUp48i4Q/W6z9Lm2yg
+8dprWZxns5wG36UFRjnIoRgaYu2QBLa1g6J/2byLchheTuiLzk+froGb858OqKa
0K/WAwkKD0ABvFZwtuKa6OR2Lxi26emdZK8NIeQm89+I+VEPW5dHMYIvPRDZ12S7
5Na80myYeMrCXfyWNv/VFJEvFJb0/IPh77ibZlrbQEMK3OD0N/9Gk2f0f1jxReZd
zvM3STw/1AyEqAqt2R9d654f4n1AZ+q26DKrLzZWHZqdzgV7g7DbcVI8GbabFAdt
8rfou0VI8+DprfVPpgYSxZeLIolo8bldauRiQBnimNiGtVD3OOR/ceXLPbblHqgz
2inTiCYxcFLhdIxlUjuGX1+sEw8z7Z1IC3p9eiEldhU0Zc6HAOo8NTk94sExqZFD
NTmT3C4ffYMlidhPlI8lg14+6co8VqmC6wTfhsM0McMRH69qG8GannuzYfKHybgm
TeogJejrUXbgSV7gwKukDquJ7Hyupl8vEsoO8HfMjKHeRBT5O1fIH8zi3hYeAAK8
2p4E982AKexny5STRF8JfdkmqKyZSms3mwE2CLd1ZX0oS7+Q3Jms4LeI9bre2U/K
3OKkw6H9PXq+BYb3jeaPLAM3PJuJh7bMcKJ+qhvXSZIkF46wz66upG8zoPKV++wJ
HozAzvLuVBq2AlRLp7S8gYvE5eAbo6AXDKop5rO9Wrvd2kQmJeHn8n8VZvWM7C1Z
RLnIuit8PYCGE9jyRnBWCnigi0sflfFjfys9kFWaHz0BPwxcvvd2s5EAHejm4jZt
ooDmDZVAaV+7mmdN67vmCipxjUoNLrYNxXNoZ/mywrki3mp9cXf9jLjdtEPNe4EE
MGgAlMc+R1LwSigacLvt93L8vZ6okqm7OtGMBsqI7rS8ZDt4g3X8LS4gZflRhbVH
Ldbk+5ae5DMEO+kCr8LjIaV/17LsJs1r2sBAzhdqEvN1owErEEynVz6XWW2aQBXC
gMEraXxDDGU1JeINPxMjdz6nRA1teyKxFkgRhG2XZhLPAer2pS/uOkng/RkK4LM5
5vIztGmyXhgcQN1FpPi2TN3T6GSAdPYJVvB4qRnEP5OQkXA3UXSKkLbpo1erQtUJ
n7gZm4TeuLzYVdTbQ6Ftqj4Fp+38gyxFov+HY/kBT/gT26bynHEeorupBcuS+0Le
AX/RQGi/jtFevFPlkTxlq84tsUfj6ElXUuQesPOwCLu0v0/1Ry6wbWvA/6Npek12
Gclw8YRhhLSa9wwFP4LKJ+3tDi2sK/SOOyjZyfUsJFJ9pe3OTaC3h3NQTxgCocgv
/heH9zDArkBdr7AIgxA43bjZQbBQn1u8Qk50PE7xtZPh3SQDvDTV9CvyvFU7hzcr
Wre1Rg4nTMenZNja/Duj4tWoNQVfLvLtfhfEY6wrf0BB7C3Tqb+9vm5MOza5Dg1m
sO0MNhfhKCcpQLxoWf66QK+MN2yp8OHR0ghizAO8hWGlnavxG5gEXcFloTw4wpyq
XzOV9e8EzPN3ESYZePl399FLPiVohZN33rUVxTN3Kk4zgxl8XOyM+g5mhRCpE6jt
DBG2JFaPMBSv87MJM2PUiIYszmXX6LYwyIdwnqbbeHgIPZ9BSzisFe8eSdnSfcjk
EZdQufXOJyqlLyew7l5fSz2GszpoUVP56B2BYkozCCzlLN54V4FB0GQGfXafAW/S
VS81PLdxJXF5jsdK6WuPRFsCnXgAaf9dfzRLGo7bU1GoeOEQgbf2S7Fhew5ddEpw
sjysZ7phEFEmA4dGb4Esi7IbJlQnHW89CwPVPagrNW98AIqAxFn9lZWQIHc7B9st
HTl71c8d+yD0Dc1lhwU/tmGOtr0FfmHhqcmaFHRtDToKJDBJNGQjY2IP1C2kUEGt
/afk4aNCewygKWcgP3U5F5XwzgJeLT1saVOFbfKB0hg+97EKGihqdCWG8R8i1aFt
BBFaVDYYzs8HN1tX5o7jwFiZCc0tiFCjfZ8BrVWFEtba/Y0Y8ux+BQJQ+sFNoXK/
CTm6REUhQOoPoHCy+grEey8Qq/IAA9qS3s9R+P/a9Wmunlu47Q/bB5tzn+gTNzcW
jQUnJAn0B+8mKh7/A7h6l5kCLE4E6DIkqxkMujPFnzRaCBzHldT5wLbLtodnO34x
cjjBFLY7TUDqDwMXcjI+7YoOyKEJI1rg2bmqdnDIvz6EQ4AgEhNIyBsxZqIQmzyL
w477bUV76aS/wEEC1hmNg9fZtpkk1A4PzWwLxUeto39mH5xMCutxibSOBA8Fe8nh
jpxQgDeqGtN0JjjGL024hk6U5MucUZT0b9adFtMPcHV43FThsxERRCzpjCs4KaPF
qRGDMHaQUFfoFrMDFbZTU+COXRsgCsLLlrzsl+xE4t6gw6g/k4I+iC4sl6WZ4kqs
x/Icu6XHp6hD8pttpvsQVYBU+hiZGQnMtxsD1GeZ8mrvB9IUiyXadHtKrKDvum8S
hIgN4BPZVqSKOMLCQscPxuRA8ncvCZZJd15sbT1PPVlnQWlnHB1SY4hMCWNCkK8H
oUrUFDiueUNdDWUDCoPttD/SIGV1iay9XbINWtB8TeINCAftWHuBXVsZ6E/9dC9Y
mnCSh2J3IEYCsHCd0j7uBGnHakYfUwO0ief6dl9dBVNkD8iv1A6aTerMCMLJeS6/
SgSCI9c4IQN56xbp4ekMwCYIxalJ6aB75lHCgo4qetfMrkneISbH81+5aq9cB7zZ
l4niduznj3dH43QRgXcEeTmuf4PwSeN7k+alcQDNMgy/9+nvsTxe4Ubhm+2rvNaX
eRG58kKZrvJAU2659lvpVl1blnxbVSfhdcJOsbf0vZGW45YIY7iOyNMNxlRZfIN5
uuu9l+z9evrlnxJatYxIlUK6Yn9LvWvNl+o1T3NBP5rZf6ETp8swRsMakr15S0d1
0HDODLmxJDWT3CAxa6xX5CrUG2TrwsSoV/jZc8RfNqJKBFq6xmo8t3Mkri2iyi9P
NMLWPqwwgSvOqHGb2cep2g==
`protect END_PROTECTED
