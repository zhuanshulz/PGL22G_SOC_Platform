`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxHWHRpwFmjhbEcMqYgwxcYcdyD4oA3m5hJu6/z47stxWAE5uYvj5L1PpoVS4ggB
+XT2xle1KwcshTXlBJeYGoWxmJ3rTszSP2dTTZzV1ZvPubxpnBlsjsxMagszCAnL
MIORcc1hD3evhHqZcm53qR8wXZ0KZ/ni+nb6n0utW9sOvb791V5PT+90YiViCyra
+NxnXXDrAgZMgViKapcVMSbI6YnyzLQbsBQpjEOtQNtbY2ge/Y90Js+Gbf3xZwP5
qJwywGBX1x6yXoELEXdqF1Sn9HSSuGbMl0mNoYihKooq+BU3R5RO5nVYDKBifoNT
QBT64Px2/wD00ochgP4w5ifynkokadErkrvgrVOjArm0rcEx6gTH/VwS1r8CIY19
YFhsClh75c3uRezn69XE/mxALcLjx3dVsDfr7BhZELVw5IkFR7G6bBUAEkWDlUPt
CDbN2EYXd1r47WYuQo5FKt0pXzo7ffUvyJgR3J2s5NFdcHdJ5AA1omHb3ypPlwbd
IQ0fcrdIW+8nYMqZ62Z10KM8BLKnxNYndqTxswijhR8tYiqXQA1HFHclys3HOPe3
1uuFrRr17G1cb7bdcKXq8mGMCJ7FuqiuKq3Txz98WwAQ1OhfisCmrtytv2U67Juy
OIS4TbH/7sFrRYKsVu4Bh3+SDIan2pOyMJM1SJv4bkbSvaVEY6k5NbsDX2cGmZ+a
3dVD9CzZkBID7LUsDKJYVD9bqHb2/K833uuUlwg/nkA8mKbYbDEGdBwt9NHKU5wA
nicu3MOle2EpqfX31NwqA3iD5B5dUsCYiPlCrK1Yrk+/cqiFMzuYCyujXDF2JGgI
eDgHyEvRYkewTBqLUxrvhZjFSsuFrFAQgAAtC9chUwKwI5lTzvFPJ1A171dpRV47
8Kn+3ab0a5KlKOOQJ8h7w5X+e6w1fVc/45BKuBYmLWGzKp1Yb4WvcIJTXqz5O6f+
UlQabApgp+em/BGXdRCH3NHzHtgnrCfUgwwUrx8SkGbv9gLYCPaoYwxDMUOuqQr9
Nge8QivlMo9MSph0BBLeIGVnHVo9UAzzlYCQG5MHp48n3atAnI5EWDznw3qoul63
f8Xai9Y9QjO0CMDVht25G1KtrGt8xfz3aNWQdSWzkRK2hkSXOMO6Vy71CWN5SdgA
Ap0vgkebr8SefygKfrHzs4HH2+7TxPKwYeedmese/V9El46+1V5h6u47O2WKjNuK
EgunZcpX9Uu8BE2BkwGhIZZEj1goVB4dwbDY+cbgub8k2Ki8fJ4uGEbgzLdXBeex
bTM/XUSr6SKLerwzZWgi9UAxUjqlZ9lRMhwegrcrLIPSuqRaplHSzANRh1yocMtA
/FSMVsBDyHVWnNfoBgx44zTCU86AxN5pc3COaWFc8N/xspzCycn01Qjz6Dhz3630
6myKlOLPVzmEUNHxW9LbIVcCmdhJ+Pg+82xlGSoFpiu8Swq47wCGKF6MLWx+B3EQ
2d+20sAHdTvklbCNpfgOOWIHb8DQONGXL+Nlb3o7k3GUkXA77Wq0U90erFhkuLyJ
mRF6O/XOseVMTl/vFyWDHeVh6xRKDhEYC+QTFubvFO98fZsdYvoQMPWfXiKQf/5s
MS07WmAeywU1byaMTliDak0mOZaW/7MFiLY505AAKKbMh0NaUUwE0Iz9Iv7Vqmba
QXaeLjq8C6y3xokRabaJLmGB5XQAdxXBi6RAmYH7NVbx0Xf4rrw7CGfLUsxJAe7I
QlHPYkf7KyZ6kjKpnJjPml/n783GmUTuBKSxHWWnaMw2f8TfjWfcQ+oSSflfeC+p
3yQxqlV6pGBjfxSngSjcEIBi/gfz/JvzLysdsH/YoG+kg2zjcQHYjZta35LrCYO0
Xc472VB5sOYfh5PCKmhcnsHTQ5diYLb7rFjYlOH2aAW1ymHhq++QQa5FnyT1LvD4
J4Oo7zMTkPimU5GBx2AXIHWh+sbNYcswQIV7dKnPAEQeYy8LCowkzs5ZhepOO3x+
8b0B9NJ+voRjtAhZwkD87bZOJGi55JClG3Nhw4E5tYZTsr+1yNITtuxAWsZf8Btk
BB4MusE7EYP6h8h2Wp9W2NP7/WDhGjkyLwwK0e8g3F2RtlLcpoio3lyYZ7CJY2re
kJoTiVu7c7WCVsr+gqOK/MkLBK4fFNLX+MGx3hlcYOXovBTvcRZ+1lkXP76l+C8a
kAnF9cHnCe2TxFcGqFQIM69L7zDp3Jzoy5inzs3Jq2meW3eNQlOzGHF6p9qsxJW8
lWBiLBJ8JRyCjp1rClycgMs2i02ZO4VABgozlDnHjYjZPBkOu0+fgdzLptMo03JZ
0yeZbeFDCYIKFV6eNW8asHG78K56ALQWfXNxj8IgcMEN5chErdh0xJHkwBMEmfJf
C/n8JO8bfMlPpaWohCEEi5DtidXNJVmQaXSsnH1h1YHTam5mm91UGBf9yA74RVTT
6F/NhRej5JNySR6hsLq/3jgA5EBdDIzpKxoJYXMhgFHW8KFa6K/eGgPvkG+g2GEq
r5kAJ5d5LebViz5/Qd4vKBjG2PbtrC2wMri0nZ/E56ezkvpREpZO37raHgA8KqlS
MA3u8fbJw3hXkXIDdGXuUT92nyEdEtMaCcXem9vYc6KstW92xNp7DlazLr9753ME
u9tPD+3wXr/IMtQ8rl78M9m+npjiySKAfJsdTb3amTbDxGYFpXjd5OkGPCxQ53Nd
lvduz7AwhFym4+3GUFjrqQBoEXnV0NDCq33YbIfjty/CEapnQzw8sbX029xDih/W
OrICjAK/wlYnuSHfhW5Ya4pRmtv+7SSlQfIX3rRUdy0kvTNC4en3ij8G3CNSHsit
ea3o7Wb5B3ETYO+od+VwO45oa18G0i9S2uEkX8kKQWXJT0QFVmEQ+AAZceL8BBIs
vp6QGgyfnlaPKj/ogw/PPblDnpsd4EPmC8Cb5DzAjS2yYhwRJWmyBWFLbCO/X3u/
WH5r+elXE004aqGEYYKGuPr7p1jI2Qgdtl8QPKwH/oWaYb27lEJH0i1UpVQIpNEx
2VhKzt/1XfaX7uFbuRLrhChhSMqg/QyCjGRiTNNxJPEgwn1vlueDMS+8Tj84TwZu
GBbHuNfL0IL4dDLWhVEArWTezvwmnf6xJjCLjOKfv8F5LEYYKaTpOCMrT2pZgdPw
f3n+2R27nsYgE/9brs5ufT8uusXcB5cFb3p491xhgrUjngbtYGvp92WWCGLtxDpI
8i8ENq227Z/seNJ8MBhNBVGmXo5Fq664svcnFVV1ezHa7XENY+5aJLJcLK66VQgD
M9JYxnneFtvxJu44ae5oA/IPKNTSN+J6rJx7/Dj8kSZ8wdS6po4CVNTyGHgOdTMv
FLo961gNON1e+0I+RGizxNVocc/t9lzWjo3qmNfC9snM7jZjQ8yhxWXKjPa/VVga
SW5Sx9U2WKFfLIl6XWFMDSljEX/ly+V45ICZfjDdkbosxYYc4cZpPck0VTwYJTtc
F/0WoRXz01Y8EtpKNe2yw57KGPa6GkbR2y5/rfCewYWey8Su/DSn/yfTvuD2ys8j
xUsjn/tkSyTh34tXWFskOLsaoqpdDJ6XebUb9w87ZtQ5EDqrcOsjy2AbTvHbypwW
/HRLTjv0lXiaP20KqFGl5eFtjBaaqnCw7AEaQHjjiisMqnRnqA35PfexOTDot/uI
dRq1y6K6g4rkul3AiQU5VecBjbqJ551kRWE8JmVIr1uJboSKfgKAoKDPKCzJNKPn
fWLWFGuXxTdk1th87BuJWLVsBAhOMA6hwcbSO4aP3KlI0tNMzT+Ti/kvcUH5kqPV
xvIEoUM7QiDKlbVbEaTV7skX8gXT4B3d2MQuoRw3wzimTpwBD4hIJ48wNP1MMQnB
ew5PX67dhLFQaMWgmqJyiCgaI56ohoxGJvdFX/1zRmtnyQuehJp3PbQfFb9m8pkt
4fAVs8kZRW4ohLOVx0nc7IHxCE7Snuyc4CDyOrrUMZOwfom1r/XVOazO+brVWe8s
5Kcdc7z779vCIPNpvHWS4JJfabxGXJkzIHRIhZOyTsR15o9X56Dh5qHfW6DBxqcT
7eMW0TihoRG+hSEB3pidwogCDpmtUM6HEt24LUNfjiaIxKc+Rm1PMJz8BBTzYVCQ
wIHr1ASBdSJlC4J5DLkNWczrmqOS3AX5IJmfP6FvFnz823+028tDCTAnNcgo+LQu
R8J8X4tg4meID98JFdKRIIuJ7pOpx0b8Cdltji1GyGCBocvjRAh3KIb6fwReuuPb
gRjHYcxhnZrb/5t6V5TqkAi6Uv1L06CG4Wr503Me/qJOSmJZe+TYA4lt+d5W1SM6
CuZ/ZGlMztls2oT3Sdk78jg2DTM5kZXx0ul4jmXBqW+qQTNiUehi40Xgtjtg1EJy
wTs3sq2CokxCmSQHx01FdebD72R4tagS8WL7090BUzVSZm/kZ0auU9iK1bSU9QBu
c+nteVdISJxDO8AxC+EXlzSSliyxYP7ikxb6joDXDnUVZ8QTau1NXlAoF988ThBV
xwbXa1RNmTQyLH0/pANJwM8ls7n2IPJ1N4O7U5sLBfWGuBGTEguKUGCL1gDZGplb
xyBFiMIhqPpp8REkN9eGdB8RPcXl9C5x1ftW3HL6A3GAYFxCU1KyA0UJQizGfX3E
O4L7ZtDopBVPg5yftWJRNv/+OlWG/xEdDL3yePNIsKA6uR8wIZN0Y26sUNKHHI2m
9fcPtZge+H2RPPZ+kHJIX2Vo57hM4363jaEV5dwUvFHWlD0qHJquBLlytyLktL8j
eKtwbkE8u6pccyW+z9DzpwsS6PnWTtCJrWhW3bb7ytA0fipFpF+b5eFhkJjoO1Af
Wz5VXDqBzlWM3kVuyslkSlQM35WvL/SF1523VMvZWGS8R+ebcstLAfQmCkpwBCls
dENKNUtbbtJCAkdk/Wsjf33lJbBLv4qS885dqDQHyuQVqFY7ovtXkiag1gVHAJx4
nTCRzvEifotrc6SH26UfID04OtpJWqvOtmnvb/+IW+u3oIh00rEpLLMfiTwJ+Kqm
Kkq0dIoNrJSjTVZOARQP+5yOKwDb6RhUj+6UhNc5KGMHpUk+QdpZZ1z697Ah2ipo
aMKSJ7Avl16CAM+2IKt+IbkJEE3DYopgUYx8VMHIL2WxCobFTIcIpIFG8QogmLsV
s1O5ou68us4bVIh+tjAnpjx11alSlzYdlSg5wku2Q9xzZb3mrtsQy2kag8oPFlOs
Yjq5s5n+pAu5OdfLkauh+BrQpyaxirPFVfkbdcVvPtwZexkFCFTmhuMw/vrJ6uU0
6EYl9kUeFDe1SWGLt/EzMdlimDIazEc1rI0dHlRR7dG03rsxXfx8TWHsEAIgFK1D
a4M1CobeCtFCpC+pvUegob9ZIUgjRRtacBH3hVTUYCAQdFzN8wB6djAIRX8E8JVm
Sm6oGY+U8GObRnYJ1hyLh+MI2my9SQY7AqNkgALRy+NkdBti1HEBoGFVOZIzWA7C
4/Ud6tIHpT9gcSi4Y0J8eUL5U7JuS2bzlq7qkUMvFPDqVnlm+ROCg3FS++q1GnaN
4C4CEfAmvr6bZbRh5S65+WVvjVHre6QlCDpnpOeaU8KYvg+UkbzsvFHMVsjRjo6l
rQX5R+eIltUu4cB9VSlQy2S19spH73nBD4IX6pPl56x48CCHQIj/R8xPgl4HpXpb
NNvEuHpUU6XCjnRni84SYJ83VUIh6+3fiTwGMT+BZi+kBKqp84KG0+JBGijLBMWP
We+SoS+d8BhCa0oQVpKq98acJaWj5GR/L/AHHGcehGNpXBedq+DqGgeSkuHF9AjA
LUhTyohukUsGoV1Qh4zZ7Px5zHmrX0PfyvAqmHQBeisIVIm01YvlYPO7xQPwDPvX
7rsu7qvlwco2LW9DhZMEl/fpDt0kySJMe1I9u8WCU76r7jxB7NKtbYAx6+61nPVc
a1cMDsfITKxf6W/JB+jbQ/X39vTEVXrQlrAAfrsBYL+dlV19a/bXdt/nfahsJDUL
jBbXllvpM0DyZby5fD7iDPdDYf/hklfa+gtYT/BYv4kSHaaBVjVin209myRcTcyw
P3zkYc317gvsDaPegURGn6t6dVuXNnw9hj2i0IomXjoYWXbZdPDDlkPT52DhD4lW
sXdqunnuNdTNwjvjTbYLHjKdFmj9AP7ATXdBpD5eCBHExjCdukPcJ6lxCJfIdlLc
WyiIVsQKh/yM2EYVcSZc8o8IPaTRVurj0ZoO17zFRu9j2lYDAjyMrFPN8DWfXBfO
9xcxyMwrGmb3yaCAbuyGj/P2GJ/gZ+cdVjRvd8jaF2nyQKpZveFtdGbfhETOw6+0
k1ffXeLBRM1b1cIXv33J225GH/dCR4HPo2S77q8Tszon/jf3XUXcc+uo/iB0jYrx
ijRyCGHU+av/GZSylb5EE1RhzkG/O2fd+MQThQdvDJau5+wKe92qvDIAlvuqtg70
umxvhqIj7925N739r8nL+k77py+KEOdgK21cWWOviJzZOd7+HWgll1Hn0TFdI2u3
q31QimW/0wcBLua1LMl8444z2qQ/47jQ0nqg73/YhuwZW3rXZ0GdOu5ZHeZFqaKG
HhhVTpoGu8M5Rh5mZRvXST0QFFsF3Q5Guvnd+/U1+XgylvV/36p7pi6K8eG3cACc
XNeKYqLG7guRPtIQeUtxqYw/8MqS/LXV7hixUo2gCVEYoaczEj9SxTkqz/YROj8h
T8MMDYIzPvLAsiFKju98/FCwgt/iuDCQsnJ7eTtOtcT/eOSz1K2aSy/xet5i6Nsj
+zjRp+yPo01/iCUsNiWV2FtL9IxWfe8pQ+Wy6Ebf+T/YJGseUyZgmKqSMVEjM0/m
Yk1ZAoJexOzYEcgDgoQLgA+ydPThw1BP6y5dqcSaDeCEKHx9nIyoM5dvAa/p0Mdq
kDnt7WvCfazSw8ol8x/2uyeAC52BpY3HeRdRuVU22sstg25wD3cOdCti3zw/z2Qf
ZCvLRai8QwuPclUhP0DRV7HDg5z+SyDVLL1O2NxiRmvLiZozYZrHxGv2MAeMWGUl
YGj0Uo6pJfYRkuKqragPbjxgUGFY9YopQmw+XTWD7xShhTNQV3JqTR9Se/rvePvU
0g+1goM+QKtqy8SOCz01ZAAH6OwBcJSn8BHuXmUakAeHjj5GUeK4xKWDOS/o49GZ
63Md77iGJcs9yEIYYg1FMpk7scOXQL1Ba13x8C5i9mBSQ0juNVcF3uaO7prURQDM
x7wY6TGG621VugXvaU37Lz21+l9WhyyogUjenxXgOYLq9vFBGbwDPjXHjRWoInKw
eTJR54/i6R2AiUk2/YHK5tcUsohZC+vEvDcAxvxqGUDn1+hJYs2Ctso60zKr0kXR
ANhAyWNRVp9D1VB92qAaJi5/cHZSRmiFCnym6c80ojE9tkaI71HlV+DJvp7Pt9qi
64FjsYevZRDtcZoIEPumko+XELoZFfHvNx1eQrDqA2Ml2q1ffB5+QtrHHzsRPR4b
2e8i2/xnLdvOXdSLGuUjh3rCr021p5CwJwgTPIyYsfGCennR6dQhhH3rh82cxYNs
x2JkRoaPKT9y42Ms4AUA+grMUF+xLqMnYgPfOrKxnoO1/ckkjThYeIINGmc/4tsq
P9+WiR5HXWeoILxGYPcaU9nJr/6jwhjjgiAr/8F85ELhAjBDbL951Ge6jgnZ2hhc
zZ3ab05TXVWPPXOvzXnxmV4lDYMe6ZQ5sgRf/kjdiFLPcuZ1gVj/GcwQzV3Tos2/
XVBrm7N5lTBh+lVc0X1gNOPHdIQZTHtCFpifvt3Um1obuvP3sBAxGt8oLWRaNG+r
WjYi6yBaObgJnhdQapuHnew06hjDy53jsWKiAImJN8jjaL7vJLGXnsbz4vhXItXP
VYP1c36Ury5JZqQXiWREE0JtvNJM0/6oNZysDS8/jzTWlFiE3ZcgQYmX7nhSn1Ws
Nt5hSs7wuk1yO7jKKnGO4I0Bf8HGuBd84Paj0bkYMGuLVLUTzrGX2Bcl7uZ3yWTh
n5DbVoVCRq9pFx1E+3kPCUHHf0llKKQI5ni3NmDBwelD9A/qtCy0rm08Srpa+Ejj
+ALQO7Zd3qzwHm+kodj7C3EoWP6ylF02w/sAUjClwusC04RFprqA5Ndzm/5Mzd2r
j/J/Oum2/0E86u1+JWrRZcbdLax/JfMzxoVf22S0A0lGLvCpK+mUxtAoEixLIBAw
lm52RkWW9IhIcQRP9iUvBI3BtUKrjc1+03mPcbyyiNAvUedebm86vSQvwMHWKJXj
8uXeaT2O8aZanR/L94gGqcr1VAd7sRovehWmMpA9IPyjIXnQ6Iwb0+1m3ruEAde8
TTpl+e/OTfNngXSBldRhKVC2+b2x0U24ygNkwIx0u61NVKKPMCoUzIaHFWyN+se6
8mMEe1USa9kemc2TlG1AKPmYLOzgePloaEAK7SmbP5Me2Mv8aNzxCBmAhcpi92I0
qc3q+IpJknYwnVn2qdme0Hh3XOdJfjmxh0vxE7PEB3CrIByxOgWWaaD3iEFaMU6d
Rryxnrcdti1TCmqEVNudrwrgUZXsKAp5LYD41a05QwdvL8r9OS5AGdzJax8/Sj47
9Km/dZwfNhHonz4EkyYjoLa1uXBtbtZRfcqvfPIIvtTz42IWylJPCFzSSw3K7SbL
92JvzLoa8qjtoStyCUu7YdXqdUZA5+ov5HE8w8yZ2lu7ilhffiT/TQQtWElA3yAW
acpuxOFhrkxG30amcYYBt2CxvHYDhPIctoqfACmEzrBo9JyzwY6chQhIx1b8vRt6
c3Czn19rMjlD6lFSmxrGMXyRPXPOMo+wGbaf0YVbAaSpL3LKQE3+ZqxGdsqXZR+z
9kGCfqzR7uJdyXUiSSB+IIINfXNNWylIHExbFm5knf3fIMs1JPKfPknzbTIx38k3
PrjPAQLuAqvB6uuIEnFtlrltaFEJpB4CZdvlgYPnz+dzZvKJTJ386IsmDgUS3anY
D24zStqvjaPo0DocSwiDrk/8vOHeJmB8H7W5wg8BheJTIWlalkn0JIbvgYn6smjO
K78cirDWbxKqlsyOCUq6IRg8LGr7r0vsJeERF4vl6fLUmU8wIDQZ7NUM+W5l/i78
0Qt+dpv+sxPxy092+UvruO9PribTHmApOa5Ps3BToB3LJtTx3gr8DKo2lB5I7Ot1
lbebEIETIEslGqVSIWqO2e277IwQjCZfWP2FWxsORd4sH+lFC4Z4jNMC5VflEyuX
OEB8z6/KHPVg2on4HqostZg7fF1pTirg9lm+loz5MTy9Sx4qdj0YaMNldTOyGC73
OvP6yCLA2VwXI6+d2V3ldud4wHcGSbPuR40crcr9Nmh5dE8MLlwL9DCzdrC7x996
YaIkfW1InUr+O15Yo0c8/AGSEji/qofLj7WzY7TeZRXGepcUQQb6gS8j615KadsX
D2VQj0La4TVEUw/JpYqXmBtSy3Ba9zBKoNgqX/H3vk5zJxzWwPFQoCl72+XQloBK
jCTMyCQ6WDUFbfqsKphMTIkO2L/WNbNb0Nj9d2Owo7erymWzeBRxnn5S6s3vo/Ug
G2gG3AI6Dt/d3rGQXQfSCRAUd74a3RNMHEo/7bI1G8fhWttPjrHJLpOEgQmSLwjV
Nimoqij1W/U2GPgwfBTmoCgY+TzYVRt4dnUT1hLoRCAmsPjc2tT80lt0bYeP6RmJ
597LrTkd0QJSq3cGq6se2O4NGD0TI2BMfNxt9YSj93teYTxjebj9dnnkM2aavyfZ
+LneVU+LQnIi2dk0KbTuVQ221OFkP4juLyMaT1xkoVvs6873JZQcHlv5vB80xH2k
pgbSZi/zlHN6nBSvd6bIBmukwYHyKUza3yIrWKfU3iBa/ORDb0CJLRJGj9Q7p+P9
YOwqcanBxFWSZ9SeDLOkqyPM/V/4pviYD3uV07fuZRu+EwZKcG+hu4YyP3/rYW6+
2yKvtyaEdWsqRviBdyVQAYDvhwDFonHejuwYBtNabVCCgwzlTJZ1C1z8DDT5vzRJ
s3I/MWB7LI7b4O40ZOAbPf3JuqJjYCHo5hM7aWoodCbQph5Uy5/l8IAgqca9LfxQ
3E2FLw0GueuA3nXOlCo9SmQNI/lN+j8YvfFiipQ9dBy8+rC71Ao/pIvKEdivuS3k
Z1QDYW9TjIWfpN6/O2afHXWfoE75XyfHIoFTOXnVmXQOs9rf2yqM43EaTnXtsXUu
pmlepyDcFEWdd3xaMot637AcaswQqNy0UMJW2RUTfo0W/U0lBR+sffIUsbF3rAhK
1xw3ecIk88HdKNs75dw8cjLymjjdZ7QNLtvzzR+wYFzoTfbIddEjBeQQAhDBRJNe
UHvGZFRUic/imzKClHoE44uJjwdN+/uR2VzjLZUocwGmajInTGgAMc3MJi97FNC9
LE0/D/weMvcSWGZEad8NadRgaQvoWyZgWqnkDLoVD1yWjPwLtPbunOe0xTzrTuM9
Ew0uA0d7B3o2kPW9aN1qMMlM/WXe7jNPpG4fbrWEVnMKh3BdAZ01/6g6b7czV743
XJDCJ5QUzPYSV6cqbp+qFu83Rlx5HosTvK+09/gnjCTnJl7TTfP8dmJhbOlpVDIc
fdC9i8RCHWpwwjEljkp/OlSASYrL6VobHgENGaI7JyVsziyAvgm0aEMrq5A7kyNt
8+/KpdtGdYfdPl2EfGzwC9RMi2LgNjn1lMmFTI5A8i5ViDh9wLhrlw5I1gr8cfGS
ErkTKheoodtOE2VJ3u1+i6mTga4y6rdntInwlkfh3ssl+EiTBG0yfadS1mNZxoiD
KXdEVYCSy5DyrhZeau4hc2DixkgqUcU0tM59+BTfUNyIAOW3OR9iRkR8pg2mSh2V
0H83eCmhZLIyrwrqIfzcgxbcu67wn7QWvWIFxO6E9RT40UZ9cI1V5bUL/GNblybB
nh+EgwQsqYUjLcfoqMrMf00T+3ckkICdDMVj/+Lp92h7Cx0PMaEBS29WUHHJw1Xt
LaeKaz1+LWOW0MRd88LuV7lDxlSpMq+pOG+uhYfNTMVq9svJyb9Q3xQUZe+4/SjM
Vu2WIYBKpl2nN7JXbc7HsYJrOvsbg8foJcLVEMHojt27Y9epYgzk/iKof3xTT8n6
ChniNBB7RXTvWYzLYh6gNzO9uj4AruukS2zB/0myxb/cwnq3T9jZ6eRK0UeiRQoy
JChpvTfTQhn7Wep5B4Z26UQtbiQh9VjjQDQ9qsE0aNUqB9pjQi3M/gtI4w/Rtdmd
rHHphyeMYIgOieJCP9uaF4S7vmn92IzLQRaaE9QgfVHBgKK6C6EuWMm7m2W4HVgc
pLx6DPJGy9L0uxA/odRtdHTnuHQJlOdL53YPfDNn0++tf0gD/ZJilZwzWvUcnyFq
UxOGoQ8CGPDMdrmZ2BsSNqOt5ShjMSl1Unl3YM389izi35YSAhnDSoyQqYq6WR+v
PWGHRSLtA/iiIZdfk8VLz4aK6LF+HkawTPfTZ1QxyDntg060Gky8Qo8h/zIUpL40
mMjGAdMC6mwtq5EcUYjW3ReZRhrY0/IvL5JGNs8kVQm7GKEj0C8aHM1vA4WSh7Wb
/zcfJyUrj4h9n6segjpfLDv69ntuVfqYmwifBw472RTeORMDlWmxVmbitlhiu158
yemDKYs6KTt+ReVTebX6R/RYR91cul9rBJLOb7nMV9/o01uMSuZm5D86Zw2JhHve
KGvQxXUKxvThgM5Pj0zmlZnesCRTLbwFwVdnYORUDbcP93U60a/mEaxwPUJHVnDq
/Bx0rJDfDGvX3wfxJqJfF5pAHAUznn/I1pNdgPiAIlD324kpPf0aws+jeICwci8k
dK8019Gg3W44t/3182eTgyyVmazT0jBQfPFVI/AwqTGYeP+OMu5W0fndFk3UY8jf
T0khOkDgja2HrodrE24kAkCXluGnMWS2hIPW6reS8PLg8UoQ9oMFl3J8otYqfaJf
P5m3SpknKbF1k5gx3czY7QAiJJtNglsfpxxWn6xWtDcyeWEuG5c1nQQa1ZhzI0tI
vUe9EgMDu6V+AjVBJoYtcroW4nJMUlg2ENv1J4ubDc3u8HFz+v5T/tnRc+fj5XQx
mULb2dIDoymqF6QhsF1CaKgMlsqJZ4aBWlyzNRSbW83PbLEgcCguF0CQdnv+2eiS
YOk+d8eN+W3EsMzFllmVQDD+BWKTLSTDDsC00ET5NgKtD9Fr4i6gxcNbzQS4dNQp
SAR88mfsrrgz1Qo4NnpOChqE+7O6Z3yPOHkrJcSP7WxzCFqSB9sAuHgZj0vm9TlJ
azhD8wjp9myERw1Mxt23mXjdsmA13bIx3yisnXic2kJOBoPIIOHHM7fOx1EgtYaC
VB/Su8fnhE+VmOPUfoU87DH+b6lq+jFtOSEHi8uzq2mWJx1Rr9mw9jEjdczzdqQF
DbKLoCrnAv//QVRN4/BZjtPv7B8b4ScQn5vHMqAc6peZ1GqjXtJIngYavpQ2fRn5
c37JWp0qOnYZl7TbQoycprb+h5YU+lJDk/Ue/qrEvrNCTGholEECxyLDOTF7k+rJ
6QxqHepaP0DyxHFY6j26Jo91D53iyL/REIWP+rXF7lkHNhLuWnjvi8cIRtaflFSG
Oa34d0UHd/+XikNzQHLajwVyFMAMxk6Mx2DzqovGxA1u1IaFdNQIWMTbyl53j+bg
voqSPaZTbcWukZmxvVPitkw1ELjBidapgY9AxCbjzqStWakbkeKnqiLHLNzm2XZA
l5W/7JPVkuq/XZmZssYuWdMKW4/h0HzH17Kz6R+EJqSYYnnK7jJNTKHSIF6AKZFH
BTP0MDh/a/EKx6QFwsMTe8rQ6WNmsAY8apS2AMQ5VfL+p/zbnT5y+0/D9MsjeObO
RoTnrHRngC354vUA/ziC4VmPzeUkklKmTUG/XI5ZoSvWdfbmwzz11peWe6jePlaF
2ruANQEfy+fNscYoUJg9nZQkK1qqCJx12aPf06wlHX8CXYRTxSDx9LrvRiiC2PXr
CKmNtqkKltCP90ihJo37xJeol92CV2V4DySDV2MbWYzq8hgHCG+0L0SlJaOy/XZs
rflyrNBf3U34DrR7n10XTBe0nN1cNn46k6slXyNLjaOA78ZzuFb65HAHG3QhtzDr
fpquhucbu4xtawIgR3NL8BH9sWL8I7ajubM+erXB1URyU2dzzPtB+yJFJ/VE8oaf
+t6GYJCWHBpgtSeFXAalD5q2OTkiTH9QiR6PrLsn1HUF3E59yTGKywnJIZnNqXpm
AK6+sZnFKmKyTqb/ActkrLiXJ9COJqwIV/mcJXvHQCxkUDzMETJ6MzxQnPznPzxj
2+QFTDKzjzDmJzzhkRa9QFDjk6qmE+WCh9uvmz8TOzW/zhG3do9Pxxu7i81M8BOi
fFWKU34Fkv3CHms14lDbMpW2OVrLR1hbxu5lxOBmboVzvIVsYBnBiwCRDBDCys3/
gAEG/nI8budZ7uyg7DaGr6B/8RiCuvzgNmNoWC7rUZrAWigCErqeVrxKs0ZzCBxt
SIrz1Q30r2qkdK7SVAPsKmMBxs6ZnZ1+MbFDjxJ8oXwMh6AvmVRx21XJlYGwliDV
3Z60UJcEFt3auiyUKIwYvhjzDLHGjazUoOSVPWa3MAMtd7D/cO85F76fcnhf4rwk
AnHQCmeA66QDzDcjb22Kpy7eFL0DO1fELD1SmORrwKqhjtSCSP2Qa9ONgec49+f2
2Ez5BIK5uHO4HuZuna7mMzVwQTMZZvbWRR19HXrZrcHERK2o+mWo5zlmCOyMc7Ps
6Xh+7g/AmU55f7a1jEK3A+eRsp+uGux5yW3V/whhY/ltmI2dNat8KWF22KJoN2aq
EihDaQrlfPVJQKr+1k6bzos6zH8DgDZO+w1LTmihsOQnGmV+T3PXlk/afRbmn1L9
hJg5WuT9o0Uv6SUXxudC6841W06reZtkNP9YouTjyjkQl26PovGlXWmN8p0Ej4Br
qrE79R7EKiG4a06jcvsGgGdaQ4x26QKJsxD3+7uhIu6s+qYFtFoUHGceejmSoJza
dXoCyrsOKf+sRtG2ngPF7sjyldA/8LsS046baKI5FD/3cPh1KsOu78EfdRJFNczn
DdJOVuMYDDzQDUjgf1BdRE3Rxi93gQQiIgf3rFdR2QWak8HkiBUiDRtr0a9LtDBf
wlcYFt6fYDazqDOmreNfwSC893jDlKq5D/gi8VPbT8S7KIva224/7xHjzF6ILVH8
YBFO2lKhPD3wk8fQZTiJj3aZV/6LpGM7/Xh9O23LR6FX5e8nCFzCTrjZx8XGhPIn
ka7IDMlFnrm7I02kvN5jTa0ax68y26FdcB5NwH66Av56UWbyxI7AlrneeXLmFtDI
tuvdka/iOBSaWsz0hSpyyR5yE04ZjKkfsUSyVhx7ZDxOhrrzXJ+ExMG0aq/QgZ5S
trfx8+roidCJ4sm95g+auUq4IAnvkMYgIxu9I65tXYsMlIGMp/lq9eA5Idbr3Kha
TYKD2d9dRXYp/ovRbg+SFFSIF56ZAJKbwDjO7k5Br4tuquzWwsf5BYrAkHEVsaB7
21J0OT7C+/IiOXsim7hViyLfjZZeWPatqhIQR/oOo42dDYkGNB1NyDF4iFLFfLdZ
/W5oVO/p/MA+dpZGhngdu1f1zlBiplhwMSis7tLAKffk5yCebQDi7LZofBREBu8c
sqnP+jA8lQibvmA1GuxGHw8uXT/+O+crfnug02W3cHOnko6tgkdo2wshHxkJxQAo
bHHfRe227GERE8yeh+hDw8owH7rqjnG45fntssetIL5H+r/IHGusosxp7x36ehQg
GAZ0Dyp4u/9pcjAmxktMuL8GR7ZJlrApZ1SbHllhuSVp3Qk4Rmu0LCLN5Thtj3Ol
wkuz1votgnVVXTd3PlKH2jXA6YB7AsAYg3y3hNOwN2J6vt0nhKrqQBEH74QjhWbU
hFQrz6fMZQ566A+zChj0Y3jm9AwjCtKv0odAd+/Y3N9osrmNRQqTfeVlLnKP38t3
FVUTXaLzDiIsLOA4+YmD69Lydl2h5yFePCJk1LUN6pOQBOWb/CevvgnV2oreI9Cb
OwSd4E5vwecu2iYIBevPjD0nov7Zw56NpOKkVp+r8WOok2tS4/D0OM1yJEQOC35D
fkBJXQh81HEu2CWdySX0RwvWm4nu5F/OyU/9uN+CyZDCUGuim7W18XS53JQ/NDOI
MQCO6bqhsVvYyhCQCYnj4j8PQO9IyLlWN04rTEbyNEYpGhU0Ow0oOUjPaJgyAwjx
yFtJneNQw4nSuz03FzMua5zqakwgxFi3h4m4oVQLJIiI01iH1FmDpk0O6u14Po9u
49o8nm3O/DGgFmhGHzF01VL2i/5tLxc1C/2UvyYl7yW5Fa+5h/w0sz017M4mbyxH
MnaTVECED1WwOOyQOwFR8xbAwsjW3FkAj6yqr9dYwRiQ0s/5xBfwctF9VdDC77XW
rurBfbzjvfPYIrvXKtX2zggGCCQeD59LLRArtvvSep9+r/Hw2lc5YDMEuvOIB9CK
YQA85kfUu5zftmS+Pajj8ruSCSYpsAcxAjBXsqUu0SXwkmi3uzt3LziERGKyb/Hm
euH4b8dQzHh7jR4e+J7MgCJ+s8+VdGPS4qPDiO5BYbI/HfwmNLD/jqyKkdA3YieP
/HGOFf+aORJTSl93knHFGVk0ua2Tu29xKvFrhBs1H726rIAv8IAY7Z/kcy9CgqjO
Bg8OGN6YgUUbgw00MUIeRtaAOivBA3DKfXA9X904RaO+A578+xX+BhD5XCaUncE/
6HtIoMIZRPqlN1Tqt7cJfymWNuxYAu74BY/Nx8Kssnw1W3TzAtSarIlNdZFuHCpi
hfHYUmCH/ewK3gg2igcnJeKXmLAEC5g5cmrROZjeVZp7KnS3XaBuoHMzDcO2CG7k
/bLjeq51RMSfv5Oio/3ttz5y5YVR22MzMrssUH4821Uzm2HBET8l6+NH0WskX5RC
jAiEzQd3s0yeeFUNtNjl871sNOxrRPDvnTDdruEvIgi2vkAonftZecI8QCrEiYcp
FM5UgzreN0FcL5RnskPxJ385EYqr7KUst01fVF9gPSDIixGMmhJtauyRzUJoEedX
M5M7od70vM/Q/nm5LV5cZC1rc5FeQkZqH9gYznV+EDhSxCU12sDBDmiEe3bDm1Ai
4A129fTLD6FMQ2E5ElV+9S856xvQQfVlC0SUUjYx+5MqKRtzt5n9RsZqwbXdn+rM
3aUVD8bnVfE79lIDoTHETtGwLJOSmvJaFvpfSHJ37+fv682u/g5Ukg7pISQEq5KL
RSbicwA77Hx0uffBbMNHEt5eCv7sSPb80TNz2zyNL/2pz7ZQxuKt1VmjxnrLfLw4
DBI6gKTKUo/kem9hPj5U64SWC5X6eMLvHB8qCF9bshfQL/D7s0/XsOCmhVEqrDpU
gh3DEt0/NTSTE7M38+y3MMRq8sMRxuVLv+I2oWFn0LRuzqH+8prpCW+/hB2mO47k
Ettlbsj9YFB6MiniXsjaDtefh4krC3Bxmjmdvd9Qb09OCd1TTBg7tHjzyAZQyHIU
Dy1ImQxZYRVTRu7+LFg9B1as43sQ/Z7FYkH8TYyiwu6nyCB2pAy2sf1rLiC8Z/PW
67CzWWaMLUdEoVw8KJLqmjXHlVBfuavDptqcAaqUHfuR9ct8R4ZqzsoyBYXqJMBP
ydR92ibkio0N4X8q4nCfcj9fRfchihc3WNusoGKhWHHhd2VSicZI1Cw93hCKlw+p
lFidPLNSNWLU/IzGa5+dR67I6CEFFW1NJYpdBtl5+F0zq+0IWgdHlCoRSzPEs9BC
zwDcnghSMf1z8+jvuBrHJOCx6sMcEh+VnvmlshYQXJIA0tb2+YSBN+yg3/KzIF0X
KzWQZB8+JKzbjPv8/nV/Z36AJjO4zkH1wV8lEJHSdPB4ZsX7ewtcB7fh5j/c69Xc
LSDhUvoAVVzxRrVux07+G0a6+xEzOK12wCNv7QGTaTE7i7Q/y3NxWNYyvcatayrT
KIlGE5NKgt0P2+kjPpPiqgQWM6XmPBhFHg2WyHHMnjakOE2UU1TuNWCGsa6dLZ4c
kXRlHkjnQQQpl8cVpJamDdONSWyL8/86KZOZ/yHXi2jbrSMkJjFA6zW17+ITRt0r
0hcBIgodaMWQ4BN7mwi0Md5Ab6s+dop+INt5Kd/GHTs6YGU+XwURpaqhzMJzdsb2
OHRRPgEoeapQ/+SNdGyTRUzEnWjvy4/LD9wFGimhAJPekwu8H/X6g7PM6fp4MBuk
adF79bktuKnLkfTaw+gQVNl8xupt5FPaBNjyTZ5at7jSNAWMp23amv/E7SWhvVNa
28+pzCB54nlv98jst8+GxCNV4bHzdflpLSnWILSTi1j7C6Qs0nFxfubcske0bZq8
buqT9kY9SxlOwjpvdmJZ3J9n4DB8oSPNRDKORrI3HJK1r6GVBb2hR9ri3JxrI0vQ
QHnz1A9hqgcAYTLA08AWCdsJP13a7TDg8l4aEzd6W13R9mOKFsobOrG1Duy34StN
/Q9yDPXX5yR1T6KQ1kIRhIOqE34g1KaZR55HkNMJGFjZjYbtBnPsA8mQHVR6uaRB
0Ya4EeZTPK9fvo3XX6YVIyEbQqKzUykmtsCWubXOAPI9oc0EKVMFaAOSl6d+EGlG
hMcCaP0zM6OF2ASYiztLhWnUVU7d3GQVPyvlSJ3NlMd9YcELVaiCmZdE6IQfv/yQ
67Ilkxpf6cqSrCQF4A/uGCBXXgqWPi/IyAoL3fMqcegYjVzfAwVL2OqX4gcoHv6K
DH3c/LLk6OZs9/MrvdKuhyqnEaf6vTxRFeGoAIn/NuS/1EV/Ec8liwVZY+jRK+uu
qRFse2gkcm+tqJl+mmSBF6gjzKwK23MXI6f+D8qiEYh3ghIr5gAezM+eTbtoJzOu
EZ6x7KZOhPPELvpY6KhSQFKDAHpVfWTXtcIZd9WdeDX/k3+0vRCxObWeaL6HeuR5
dNkcWOHT6oBfNrt0wvEUnVqYYvkgKUPmR8qvcyUBjSzdxCIgkbDcAPEbrf5nPuBZ
z+LgO/nLBQOldy+97Q7FZp2B/8IHC+H39X0oaVDEUvVt5T7zrp03ZhSDHmH8XLAO
+zCzq75KAJ0MS7P3wbYOKCw9YsbJegHgVeAvPmen0UpYshvFhXrULYban/gsFDgl
qlsZW5NVFPsh/P8eATpEdKi1VvggKLO9uqwp8ZWJdtPGIP60LuA4d483ksvgkXo/
/tkDmilv4ebFAj3ORo0CvDhRDXeVb5ywHHjafIlWoykKXF2mkMY7Y+UIaF8UnqHJ
F0pOcP3WFL0CVUjVze9fFc7vkAxMeWI6l9SVi42eyuXNvyJysD1Pqg+Gi25DmfUx
7qNdgbp71GpWf9kUbhs14ecNM5CSRkdic+bbv9IYO3nCrP0Ir+IZNdYwnmHcdv8r
Nfsp2HQgys3ykxK78zv5MF49s9leYI19jyttXsZ6ic3MwAzonGLM3HUuClgsXU74
1mxiqLTqrBoCT431qzmCovLw+YCX0VXwQNsgksZluO7zLPlGMYE4lfEsoZdahwBU
rEpLVE/4hinuQASJ3pitDDb3Lr/f7/1xVo+1goTi5QWPKp43vOx09mO79YeGOul1
L7m4wpqieNSRKfLluTgmdhuuNmosEbDKTXJqgMW7etJLFCDXTydarhc9qzCQgZ/e
23xsvK20bkle4AnmPSLXo2y/pxnytGF1b20gigKurHwZ+alXTHNlJ2mGUQv/bZzh
t5NMLe6edSfg2dXfO0nSNgdYtj1bRFkWuWDeF41TkECm4UCdUAEqxxxbbM7o9yGX
0RSgG5WtGglswf1MyZYFbMuFFCl0UVe+rRoQvHNnHxCYJ7Zg1EZfYsdPeFU6qraO
DSEueTeSVFjGtAcIN8OEaAgy4BGGQp9wihGotezDSSGi9cgtdkZ6njCbKf+hJfr5
YXVpuEg5xeDMmJFpWqBzXWDqmCVNOslrPIY3T/fZidXNp2cxVkwo6b7LKDaKYny3
XfaO60fLMQhTO6yG+1R1gZHSDvbb3/Yf9j0x0MySvvo7uOdY1t+1vY1aCwrLLyLs
wS5G2rpFW+1c+FY3E+kp72xTtDIyVgCI+gU37s8nOaE+T+NjTSJ0G4B/Z14mtQci
NgDY7bnF+yiasGNw32ZPe0IWhlPriU9v0pXoN7o+Anz4x2FgXthiocBO3zhc+vhy
2kFgwxDYiEzMon148JjySX1zkq1qVIAULyciDHkv434j3myoJPwlzahHPadyktkP
TANOtK181226JjwMG3Uf2uGfJGP5eboBhJRj7aMBEJcFUJs/mnZTs+fbSTuA2uHS
8hT7rjDUCP1NDQBkTSHV+kdfXjUVOfzekghgiyxFzUYWcW2+LdR7UufEGz1v0V7I
AdChL4Ns8OhB9blqtR1Yj1zE3zsNMH0RaeldAqFPjs4qo31Zqfs2sNMmyUWyCpmC
sG9fZumPu3iy+ywUA89C8u6SkR2BjL5bYN0qaLUWB5rhuPS7LcuIvxcrmLIXAsEt
X3JMKIZGCralE1We+d5ekHVtyqUnDvNXoBWsybNxrr678iTrtTg4TF2eQUs3bJpp
/g787sjsrfd/SSuOmEBRagYSXIVA8jc8sKTfbFfNnVBnSQf7CfVL1dBJy/7w/v4N
tg0wODB8dESMtkF9/BFpx85ReUz8kfx3bBPCZRIIIyEATk3VCJZcLakVhSMmKKxp
v6d0UCZ0lwONIendtPL0L7jWBymKuFIKKiWX80HWxoVPzT1SBj3g4k3rbxGrdbLF
4ouWeL5RmpM633o6mxixyv0P6vLRIZZMynxhFGCanJ/8bDNtKU6S/Qh6z/ntJpVT
fVsE1QBx7JqAp73wQQojaAO3toZj0+guNcG/U6V6wVi+rNNtEbTXaZsJKd2viZ51
sTPJJdWO7ulVBcertvnGWJyMwKEtrkziF1Z627BJVGBZSHpXMUWyXzsqNLMHvwGY
kzrN2SML8F2tH6+bLAwFuApTqxWva6wWejZZexNeLfaxv9dbrLMNqtGrYZkMXN+p
lMgGlysoFikyiGikx9tk1ZMhs9yPTO2Nm08/7dFkTKtaa9L5oFuHvS+nfyoToz6B
AUZTNOnEauoVaYmBv7o7zZ/LCdfVHgeblZ3sk2nbuCKv2Oqy9xTOYcsLzBwrxtQ6
8QDDcrQMOTL2lMKgv+bKRY5EkuMgfqHAdFfmsmUoA1FMt2WDqFPcmXZf/Rdhx0Bw
oupXTJPzVW71eBAY2Cjrwc5vp5g4jbZxnPfHmRehhFZpcmxlUjblhETaLHMZZiVM
jtncDxGfuF9RaHWI4i/OuPES/3uj/+5nA2L+d9HJsx2+VNZveF0SZglZypsVRgPt
ZL53s4X6M1hh0jk8LkBPISpRLcKlmREfS9iyLB7ygPaNfSFCe5kjwcgVHEYfdPla
59yCqhG39LDgvoP2uUExDtDoz2vPYEU//4RSzJxTd7IBZpiAyL1cat5uZ/relaUB
+Qp1p528PAya2jI4LTh4zQfLhNA8FNo+XkEVwoCIAeUgIq9EM2utid2EnQ7LNnAJ
qATF28H6tXC6w2GRip1GX8tukxY0nE6ihE457qSLmjtpdJxrhwjLcbioFzlijKiy
/EklWR21CkERhqH8PekQM0D9DWaotslcyQdOJ/8xFXzkgwPCDAgn2qaHk73R2og5
f5VEAR491qwBNp9hk7p+yqhBULXXZlKCrb1vtJSpq8snXUT0s6LzPB+C8Cst+FPH
rLR5P3XvVOn7KU5Za+p2dvC+etWS2QKYoAF4BdSKNWLynv+DyONZNOhNjA4Gfz1K
EAbsmm5SNG6xshOhp68Hy3s3IcL0zelYP5MnzKT05KFQLAI1IBi5lBu1JgPv0/Ed
RDkOAXVuYwIKwvv+S/Vqnc8+N9d2aRYfS8EYlR5T97BTE+ID/pnADiF7AOf/uzRx
5MUtdcrvsqUOpAriFJLzQTbdvWhVzeoXMforEzmcCJFBNF02HXN80s4P3iWgvySO
NV/7OAKvQfxhVFD3FngVpfE9qPaU/W+Eo9XgsvvUMtgYVVoGlpnAlT69+Z7P+iSZ
pRuBw9CCY9j468RIYPxxEkGQGedZZgAFg3TPf+YYXyGo77dvUoQQ67p7Ca5nBoO2
tyQHt9RDKf6Uq3WImhZd8A3Uo4+JmLiYUBeQt99uEYap1ePVIGxHhCdn4tteLOZi
Tm/9c6FsTqFAWf+Z9Y2HceIdEKz5XYp/91lIDJojv+GCfOLjsdt8AEdXiuW4ch0H
b+KYjHhgonTfWDe52u/BxkJ5x8L5W8vztziHOtgIu7KMx/pYL18IPZAZphMS+uFl
locVZpdPwPMx0fHYrAwYJmS21KCp5RLUlYTiQfHOYi8btSoEXIT+bPiEikOvvbp9
fJEmpVjkGOaCQua+Fdc/7LWHZ/7xMCXIQX/BzAljKZQJCyXwMcxAjfR80yOOtQer
KswMC7WsY0g8Fw+o/YeQxVIDqAtSb6PnSGxBkH1QImF6KoIBOgRE0F+GqGl2fH53
jTpm1646I46p/prr2ouxlUf474RNN/bOTnMTPWT6KG0//Esfc1cvOZPu4WyNtDOc
FaT/0ddpShEntyH4bPS3MNa60Lf5NvcgEnFSPmXj8/0jxoKeCe3edVYyYahM75VX
ADeopCTf+9/YSJC3X5gZaWqCYxo4GdaA564PGk9KFcPLuabDN00LOraG3WoHLK6/
n4QG66fLau/5aDcvk+ypu1nFPptTiSBN1nKfOoOvPhGzR7Xs2qbB61zPp80PhRs/
HrOygYSqIkSzIQ2KwM+5wRoJGbmM0xlFMaNOFgwTsqjn7sErIngs5D3tDLfbl/oR
vmCTancSOzW0TOPWjFTwdl4qYw/dX8UM7Js3RQqF0JtikIU4A3D2oio4LnP4eqTN
PXvyXZEkNB6Xk/5sspjBjM7Eg9YCuE5Bf0ZoKcGe+T3onhOqjYCUYd64tmLaiso7
4YWSR5MLSXYctaC56eY3OdtOskT5s9ZMAK1aiIBJarqYf3kSnm3GPNDGHTAcC4kP
HHkCuaSkzbSib43WBjB+kCAxdbJj9rQIhDDhv7xajg6BkZbXjyt00jh/9PQ40/mN
6QVjUkevknEUGLfaE4nRglGCxIQzkTnoHQO9frn5Es8GTHqF3KbmviL/UDzFK4Kh
AJj/NVnyJsDjOpXvj26K71C23/cWwlkMSSkF5YKm04H4KgY6ITr4mze+sxDlfgf1
BV8BZVT4x71rP+Ng1hTFcGnukAg4yL+5XAi9euPUQZUBTK+1hzt2TVQCui6ziK9d
PdUrkrOIVxd7BvOGX5iodfWgnx8cZv5DBaxRdpXfqoKttQW2Px4h84SFAI1L0dO1
h3g0URgv5jy1qQMC3WYXtgk0nHPI8PdwvIa2Vhl2Pk0ZshVnIhSIvD794MEofETq
jCtNMqxKTq0Y3Ca4RMsd9pwb9rAAGMAfb7XQXgpyMUkDdXAAEi13cGwCtWcAF/Pa
//j3i/HwxYxg1W9m+9gCRQqmZhApIMBIAA/R0559W/d+UBtTBEISQdCiaoKmnkrf
fDQYnCo2ILeOm+oNoiG14i3kUgM+50JkNcQFpU6vLu1pp1wFSf2NufBs2Cs0RX5o
p5VSwDuJ8Io9Gik0R2X70l3TO9Avbros5+DPAW0qAVrUoPso2L2kpvhP1G3ltYLz
Um9+vbjJZhSn0ODwrWwcpZgwXb7mBtkwfuBDXYjPFN7UHC/mG0JH26HKzOf3cW9b
dggMjlUmJAXhwDgLK/7ai2ccM15nmMCUc+6L4euF4+1nCSx/Clfy3vDYSq13qe+b
sPqeWS4Z1DXEV5+TZbJtOG8MDU8NEnM/l2beZDtgw9STiJEfn05AhiHW25GrKeZg
ijtsQCqOKl6fQLX55yZuGBCoKGgK2QsS2L4vgRw6PIxKwHq2X/1YSp1FzBRUpi66
ulx99mtnoZpU5ohs7dStEczxdR6d3UcCMxbwFPYuBVfSGI9JUPQj7FAzaf6fXjyz
1FBeqeZ8NgSfMqUSEhV+fJb/G4f3P1Hl8WtWHKqDIwrffNv318BFUK9sp9zhusLr
rDBa4awp4dsKPU/idKn2mKp8Y3PJ7tv1hmwx296Ps/ePk4fNT7bF5G7fnXWcI2B/
y21ktNAqvIYfdi7DTTYcnDqTCWnl+M1SpyjkIKTiwVtG5wBYJbzJSzEq5oMRrlRu
v8pQiNx1J2Ux/goyuNeGmDOyMJ+FnwRoROUi9FjbrXVv6KEwfjZB59g06vvJHqqc
828IaoxCpjV8iQbPVhX6HqQVA0TRAE94ejy7ZVKxvMyUx658bnjL9IcWvEcKpFEx
Iz66J/frs1UEFBpritIKwHAnFkZVQs6qzvZQZrg+OKs+fVEP7ECxuotO9WByxavD
39TUNN2mvo7nWu60iW9w//mscPr7TvE+hIUBZRDVeeo846HP+eVkBOUSFS1isHve
fR56ngNu+yeJgiIdfh5uA3mGW+Zm86Yjt+rx/Gd0A9V4QQ9IELmWRQU1W8kgkauk
80lVGsTS68PxQizgxLjo7LOEAKGIrW3sGR4yzVXbgbZ90F7GzDyDixOt+iowYr1t
s2Y4WOs3jT4SYirpJyCuMgWHS1SjPhy/yWXzH890Cv3rYn/o3lLLcunUn92LdW0U
8VGhAjNeXn4LLt5TEm3p5JMmUBHw3bLJwrbVpQzoVKMPFAQAXiHshGvdq/tzPDre
mtgmJsfL2+dGjbnNLcIFJqMyoeUKeGtVc9CGvhDjsogoe8N4hoaGKx1JGEmbhz/c
cG58ehzFi7ZUIxgHmmgxPTMRnQ9CkRu1k/ExHfUfFsuF6VhrF+0fxgwhGS+OIPHZ
9RYeB20bfClOEG/VKI0zZZ67g67ZBFd4LwyH6Y6WS27Q4Cg7k+VA9BNI7boRtu1J
gZHZ4YGAZAjvLNpslcE1AmzAz2cbrZeH6cWypnatw81LSex8mRLDiWEfxAygw+tq
eTYBANGrxDpoR7K4K9okEH6zpObL96IdEBUwtL8TP1xbh88a9nhg22b/jCLfEA7i
DyP4oc7/XyeETMWvij+048/uwUY+1dojOz6x7eLAXOcZALlMcWPdY2l1whqpCRav
kXqXa48MVwj88ks2nwCsXrRSyOmOqQAr/CGB37p2JjyfbOEx1T+fPrILqgiS5VM9
TfkoiLPyCUzuaX0kUCsw79GwcbbYF4Zyj3pqHPm6FAxjzj44/O9ueDi0+Hg3qewh
JCTUGtF2zZeDYwkXSOu4a8v4Z5VT5vSWbODD0EBzrVuYhZxlUL7vu1uZwx5tLupw
9DcumYcr724SvQPtnQRTQh9FbideKDgzaMlnNcTO8cHLqjTLfOEbG+COSTqCJizi
+xsgaT8uLE5oxUf4IA5mzhkryK5Xa8y+3ebFhScNOSIam8aU61yU1d7HovsfnmkX
gHmNLrVTIJ+91vZkL3anLsEL6ZlJQenIwmYInMAx2VsbxHPxPBqPPwOLciiXRsL5
IYGtVq1T1bUWJJpevRHJrYqIJ8pCV6nJSB6zxOrhG/+q7YzKIDHdH96fjUS42kyg
dbKBsfTKGaskEJT8pHA4fJdMTry8zSl9w74HUdcSH3T1aeGxtEiMBqmnXEqh6Uig
J6vBVxbZ4+IiKh/u/VkmXKPD/tG8Y57uV8ekWwsbS3BxGuGohTcyYf2lYvct+JtM
FZxvw0Bo0hbRtBREZlsRPyJLYtdUCEZ7xyFBdDk/OuZ4FnbyMmCMtMgk3pvragZD
iZo4TWXCTi/qD8fRNFlJnTWT7zyYL8EvaQRw885DRMF2Q3y4zGAnZqnbwyCekuO5
gabtUa/YyKBUgd+oSuUdwPPnp65PTAYsFyNfpb6Qxv4PToVQba600ytdeC0/iolV
47uDVjQKorAKG7+1fdq6StS36OoSlKFWmVHVdf/ytLxXzNw/hapkjBW/TiNOlqbs
IsIAWftJxZZAjMB5HZWZeBRZCAkymbKU7vO2sEOTl1BT181uJhYQlYDcueM3FFJS
q8B/3taxernKPEbXDOVF1E6v+EFcEbMwDnBxRRz618SVIygYi1q7k4kt3IMoGues
YQaTSJhPdzzm99IsWOQ7Sus4pEKtzshOU5oFl9dEPdaFq/eddoqLjZVp2jOw4UK/
EfeHEs7f+WdcvRsbeQrGZAYd6D79XDrlTPHp2CkGm7zSkGhSw/cd88dSj/nyYenL
0yQb3DOJAwY6w+lzLoZTh69ZqUv7piim9JTzERhnOR2OzH50F1tumYk/b2oPBe1K
bi0NSoIeQ31EBcOYcEVlmCWMcgQHSAecuuTHoNHqYwZupvbnq4RdTGz4gYaPhwAc
GQExJqoTLHiysggGIPEAbqXdSelp4NqqCB0SaUVqyOZNsahyIBtLuYmbOy8+0kpo
DZxEBrcFBUkZLZVKO5F2MHmtfEqHa84m37eDpi/Yha2s183FkX5Q/yhFHmSPHI9d
mUSroomueayMU/SUfR88AmhM4KzGONyK+8NxVIrVXJYyWxXfJ07rf/LwFqaOpQ1d
YOWdcjZooNLeIz6gszSZ3ayilZ0Cv44JGPKKohRZwUoMJNmYou3qzwbFQT+3M1Xw
GfhaEpy++qLc/AJuIjwxTPQTiTcOcwFWA3pg0FjN4TEbLpGb/25uOb21eKiLGNoj
8v7Ck9oGC0Lv/c5qIVI7k11YLNkgW9hPtyYbzD8EZtx1RG1f8MsRrdRrCbdQGYmq
MutkVUdVyD5JXT9V+QjE5ma0ch5z091GyJQd7Z3y1OmO83Dld/ufR+87Ux63qExb
G6EDf+RWSAZkdS/k6ALXxNJyOe5C0Rlqv5q7nlcoxPCWVwC6yGGVgJuIBxsgmGIK
7wihdhvoEcQmUq4TKhY8PNaYePZuoydM23rXBTzT0Vf1u/k3XX4kKE9cMjKyg3az
uT0+I9PMMyhvps0rUhUh5tqfMVf7vphzPs2JvRdyEPVik/bzQBh8c4dNWJdj8kA8
R6W8KS5YXxoQZTjqO7aEgRTQlvlBjdfuZV/xuPDpXZVBKzECGR7RTlnUHDRs1e0/
cNRFW548f9/Um3gFrFA142C4X3BDPG+nQtBlIg9OFRNWA1K5SN5t36O6sAXzAgnv
Y1GW2pKEJ2xBFvD3GvQAhP26h1Zls43qs/vdMIJNuyzKfqHQo5rnGwqKJLAWm7+o
qXdfaqz7qvfePqG2Hbmq2D38Dp53wYABT1XHb++N3m9zl8YFhC5u++N47DUWz8zu
P4AAVyXIeUto/YqdkrRc3x6X7mxdeZ/g5IqFi9t2F9rFW/xaAbaqPlsWGLRnjk5t
aJBIzT1e/aOc56zX56QTP8n8EpGUoJha4qgBB17ku/VhVefjtsz5lGKG+k4rXk1j
lvZrR4XMyCz6iRIQckygkxEPnv/hlLu4u8Snh4FCfOvABjYsY5ISHkQJPEA8fe8Y
p0/dupdHFk6C0k3ejQsUljIOFJF5/Et7QjKvhuVz48OARdh3wjJyWV7oC9ZsVmrn
nydKQskeLaeACLItFM1Z37bMYzwXk5Lmm5N2jwGh33l5H0YaLmmTUgElowQbil/I
M1wDrT9ncSMxsPDWW8i8NAX4mr8W77cNDSasZ2eGlwBIkW3XG5+oys0e89zktya5
ASPIPMosA3BSPFGbo8OcnT/9CLdIsrAgr7Lm3rpnBiYIqktMs8/UgRkw1bHMDCG1
NHbhc66V/01xsMZuLxy9kgcKnpzT7scmrfTzScebMU7EZ2MpFgyttLfwNoViUyMf
cm4xhvVz3l2Esu14UsrzRCNWYuGafxx99ImRJgsRpa8xRzw4FT0EMKC3vtSW+Hif
JHoO69njfgpfnT/bzf7ELgWTlxiddU/WtmWzafUHeuqv3rEUrOVi9/Qv9xSqaBhw
Yb7iI9ERumpI8E6zoK7xzayfJRD4AWz6T7NeeL6mWx/1/CjqI9TW+DPfB2P01tvt
cJk6N4O2J18PjroCxaG2x4XExM3iXveGnsW0+sTGcWlIPtDciYV80ugPJyFOYPxi
LfMuKPfBmNHEYXlovl2ILFK0So2uetlTXYe/laByi/X1eY2bDp7Uz5sEyRh7DL2g
xLVWyw3jA1nZn/PP1y+bQLFCmrhX8sP5w0JArY3YwXP24h4008T9yMqKzVbEN/Fm
h7+3EM3RfIuXOtagrx+tUHf6qngnXNpn7C7T4d+Yc+cRReZdEPDEaY/VkQx5sh4S
g4oigq1M9Lie4Rq9TMz82Mtxp2mLookHToKb1oY3VWzjD3rJaQD3NC6UOzq0T7Uf
fF7/OTzuCcfEwBaq8t0XiGhVa82+RU3UXjRBhvM/b7cGJtrndSKqS9NrbBC3Na4P
jQvz7eKxGe5XS7QpRcXIXdcUsUpafD/cI1xTyT4wa6gcUhgd2bbB96Vgkdl+NwUy
vTmQJcnms0PRx5JYzPLuu7nuAEivTfdhcCOyNVphC23zVjLQPF6ZDvPufkjF9DFU
31Ne/VkPbDMvZrn/2iFttVfSQhPN5E55FP3nkiHMsiKB9t/qqRUv5fFSAt+Q34af
1gZH1EpS9W9UhuGNLiGK7qEJZPlo2jhLGq6bewPjhtYt+Hru2H0d/RDGK7gs6cJD
6ChQTiL6k+eEULa6MbBrV2kp05cA1dI5NxrnXooas2ApbnEtIKYp0vxb0r9JjjIc
7WVI+VKYr0nANZcOp5lEpSe9fKILHsyq+m8qe0y8qAdeOg3QmcB7JZoPS8LzQMqL
jkQNPnozJ/nx7ly2zZRMyhwb5+3oQ5W2X2I8AjdQdRoJiNEGl2aNAySAl0nvMZ9Z
G5RDzo7ShwADPqRwHlGF3ZChPmItKaO6piFTWlFmsPEaN9O9orMdBOrLXPQM4kW3
zaO5r/pXBI/emPndmudjJRitLf2MSiEVHT8+qvPFGXEMxcgLn8vN3+6aewpdpRCo
hC1pC5NtOzQt2RyD0TJW45Vq7RSiB9WVgLsHi++uCYQvGz4mrjMawRKlZIv20cqO
Vy6gw4o7maezYPuWgfqNF03KVrftlryuVb8jMiFrTP+Mkd5T8S+oQ3k+9m96E8V2
MCHUXai4Z7wxzChJFexkHww+U6VFVlcgvc0+XCVshZuVJcwzlQVRBQCf380s2j2s
OUoc/BXJV1pbSSTZI/+EixpbqUDBMRuJ77965y9NvVm/0Wbu3phbnndHaZxU1bQJ
mmZqEl00YcYtasGv9Q2y/iMWJoSKnWtW5ronuexSb5a3Z5iQNh0X/yc24fw4/zrN
8+X09hT3Ng8hHSE0fxeYajVfiOfNQ9RaU0OFOgVBHaahvbxRBR4FtIAbQ45PvckX
u0DQ5USFDTkIoQKR6vZoT4Pyy3XNRuYw63bhpaJpAc5vsfQPIHZdcRnxXKckjtg+
eCncKpFAdu/JRhP9qfNcLS+5zz6ZtOe9vspVzWw3XP6usVE1minD7DTEZkZWGBAC
DkRiw1L/P4njbtKC8T8mqoDhOEPBrXeJ+S5wv4Vjk5+NuQLPA729JBpN+kLomvSq
acYXhHeUmhmAzz08dOeWmNIzmtv2OvYGvkZUOZH0j23oMjSWJyvHKRM/22ABCZYe
RWWQ95fMoHxkXcuByoUJiPr04X3t8IKHSPfhd+Fy5BL2aKabfxaWNuOKAGAPexxx
rj8IJlYAZs4CUuWYafkIkooaiPErg8gTkc6//T66hEJB2uF+INL3Lm2WlFx3be0l
iI0NIdkgU3RpTzOHZxiFDCBuZILQRlEJyZgt5UB/XDuJ8Y+TfsIStv8Du+sgfL/1
DN0zIKom1/sn2pmM1yzPRd48CKhHCWmLY1jIBEq3GweDh8vFmDXzFqQ7pwyxOE6b
Dd6mCS7hh2YUvBcKjKbTnCm9rz0g2qU1cksgfCF0H1wmFRivkw9xeqkAAJ7l6Ebb
cX+/QqJtvkY126aGN4p2tKbKI7mQRumUuIevDm7UibAFAWZluNRfYsGMddVd8PCg
JFOD1K6I1dKQSd0O6md85N3ocYDfnL9IW/lkkWdUrsXUzBkNn9eHp4EFce8yC1xV
/gD4aEUVD5vrVt7LXtIiDozQ3/4J34fgL9M+aUOdh7M3arxFBwxvcrDfBTDfDLob
lo9ke86atzWXiQsJnG+9wvYdd41zKxCm7W/EUS3azacGsi55RBbecMltpnBpvYHb
uziVzvDZNlYfQhwUuigod4ADMnE9exfZW47zZDTaqjqx8ATp/JeXD2zUUM/JGWIi
csylzE6RQAZHysTq97qWipl308dxM9rkeQsafE0vGgd6A4V63LQFe505KzWX2Pz+
V90CT8U5FUXsHP+Q2/qTp83ze3VJjW3EYDjcSmAo06d929ZRBF1VSE+q2QllrAFS
TujvWZfSkta3vgsgBGCSCf8ESEjZAEN08ug6vS0daD4FjPQMdoFNSvXbMqfYL+R/
NJmkI5tvIi3nke04x2pYWBnm/LzBSpf3SYDbe9ckUKXCo2h4IQFl3F1Ubt6ZONUI
zu5r95RDX08eh7THVFrBqj9EBjbBYo/sd3s7m87sLlfpRfyBC4FtgpAkLpfYTPbS
v4y/b/m7MxDOcA6JdvFwVszb6km2lFx8yrVmEuiSYzQOj2XrMd5tCYEvflUw1qXr
lsqNQWy7Bq2H+dzyxImaoz0gBnw1dIbga2lunNn4jyCgOPaUFMPqtq1C1GOaBReq
SxfycYtyv7ke5eDf6z3MvwJ/aEpLeuQGVnmowoTPluaE5C1JnVHcQD3EOvagfa8a
2Q2SOnXDXwGtHSZseia8M99PMRLdCZ3Pb0u6/sdhtHA2Qh+qDZcge+3+wl51MpVe
ptruvRh7o9v+cFVBXRmTO/wi5ENf5eSN1pfO/sCBME+hOnVotkHHahrtClb0O5P+
F4qg1K5tQ+wAM8TnQ+AHrMoO/qnp90QKzHg+7XddOx3uLXOlC2pS7AJaJjwJeLBk
wcLFd4lYqhSdK4MO8rGUWJKIi8j9Uycgdy7L7KB8fPtLHuS1qQEhIyvvsVDa6xgD
LPwpJSHQS5cAz3Ctr7p0+dylvep8D5wn3UsnIbl/2GcDm0OpziwOflnv05ttf1zN
YpDv7b9jDS7LJjJo3+5ANQemEOfwFdgYyTWvdgCjDU7uWxSaq2ghL5iILoyE7EBj
fgBWSsuWrgyEuRvSiOF8nTFGqKWiJWSHel0q+R47IS2nRXE3zKKVVKfz5Tbv3N5I
RKDDktBEe0r0VqYMbt4/eJc03yL4HukJHYmIVd1QWy/cMSQDeooH2gYsF1036RVU
0ERmMJsNCZtsAWvqV8wJOZmpu8bOFzvo9KR9lj5lkyE8RqqzXGb4Pam+xdT09Mcq
tpnYu0poOa3ItFrodcSS7VuvWWS5hEPThsH8eUOcnLB0Pm5YcpOQvO4dtKczfeix
xze3sU+BbtdII8KZ/w4bY0Agezu4YpHJAkvPiA9DmK65oXM9AlUA+p/s2nwfqvAq
mjcKgGncyf1F0DNHMLq/SYkQ5TyUZ9us0bqUz5TGVUNOU19i3Oyfo7WsDApdBdvT
w4hxRDDw2Qdg1OZjQMeJC37O1sy6uXtqqJEzWaPRIsEP4O0VudpOp3rfIrZFRP1x
5tS/LvG6PPPz6qXR271wJsFRztr87L47h8FFr9jDmLXoM84ICHrLUzMnE4VA9QEW
Gx6KmGIFjLOWOAVOTBxIRf7i4iAganvm0IwobE2wDMQvCkOXjgejA31E5PbUee3e
xfhDbjieg217CwwrMdB8fZpm371MpJ3FyKunmb/mZWURLx4SdzhvTndwU0Nmazbx
BSemt3VeLg9VKH7Mw6ZhS5/IdNClq1+5pPP0AzPSevK/GfIFfiCmweGvzOmpmdkr
t4XpeVoyzQAUsHZrF+w931Y95RBzjV06AQAkTE+IJe5hyXaKGmS/HWzBclyjMnnh
5WKoZCaxmqFv37/O6iD7MVlBn0np4yM3rsp+yasES6vnxTuDWvKhiK383h5kOFOO
gWOTJNiDEYf7AIqiA3g1nQiKwXzfmgZaraM6F5FeGzlECbrj0KuHbvKILQHasWV8
yZProASJRrg/05Mz4sfbFqcfYqC7bo3f21WHhtk4sUw9yrcSOi9EPkypmXWTVg6P
5hvnPQd9rcuaHtKXkxQo3OlFB2ukAqcHVWdSfqcLLo93HQmhcbXXoqOMQtxC0BfO
PhYbSGqNbgcfZbsaTM1WAHeVoUG/RrE+89+XJM4X+S4O4JQ4B1oBK4eH7lwL85ID
3qQWnOFRH1tkJ3Yh1vaabi2KAWuGZu0jReLmdaOA1DffRt6oIscyv4yo4lhG6Bib
EIzf2Rr5UVIumPQ+WQFiYT1MiyEZw4xg9L8piWjarZWZVot2qRe8eMefITSMliMW
om58ZJFH9tLpa3LscIojE/I7B2DZ9r5Iunfp8JyB70ncYC7GMwt8/qkfNWg/iXKL
5Ll9wDokwA7+qljyWPB1qAVjfuukb1GEAAtyM7gpCWOS1lTcKpe6us28PHyX6sa3
aknj49x7NWHdXLf+SGcIvGdDyAgX+Z1MUmIeOUov6pf69ouCo3FURWcdicdBKzkF
gQawiMyndW+sogsOuDTztwmtXUL1jo3XxJkKgCwDsda1kWHgg4msqVYajb0qtCDp
6406cwo2IErd19C1Zlj4ASbF/31Wy0qHeV4/VMnfBE2RGkCMPneYgpuV+8Da2Wg7
D0LccWRLAQ/8yPVt2FSwPKfciT4j4mjWHu3p5E7G9evtRiTbuQm7YLSx0xhvGwvK
TDrLsRME3V6Sn/fkI2GCtSfVN1Gcr01U8U7p0s7LMm218RU2qL6motXTbDy9XTxp
JXtcB211zCNTeFVMMsihVy6UU3+U/0AuauCaJNnqwI/bKBNE330x/KRc0+Up8INx
RM++StiADTsZZnwwRN8gnxQbcOtspXJMLdWUU9oOostlq1HGlRHLwJQQR5gBS/VX
iFUZ2v+T6nECYiGQy+o/cdzfIJMtwaIfEgiOfkegxBq8zJBRaIkVPigqxQsiJUUT
tsqIvGHj0U8z5sgLDoe5c3xkgkQvclBf2Y3SU2Y8Z7jT2aOtZbVyvek4gxHUIngL
lbSRH6Ro6PVlMeoMlb79WopSTom4BCo4Mo3uElFpiDRYlf0+AZzw+mRT/XUxSCbL
ul9TAiQ4U6PcyhTkMy1kiwahrY3dzsZKtLWIYfrp/ol/tAw/ywSysDd1nLFBuEXW
t2zlo29uhxKxQZoVhufp+cujEKbpj7k8lZtEsAh2QpsChVnVd/A+DEM7A9v8lcGl
BXGl9mNBhn8/NfTHk+VrWPnZ4amzQNsruv/FkHwgBiVMilU2a/RWxjX+BZWsEGrh
es+9BAE3GlYeeJCUkG3E+TdW0sA0pRdrmIHer8tbFk2dUOMJ2Op2BE1RX+eMKJMr
eJNDnibg4jt02ddXmP8BReYVWp/Lm4U+CR+UrZnuXnZi1DluO+W9ANE5qWZPh3mq
J0VdHSheanpYWndjxd47qE8cCr4hXEpZIol/lywjUp86OiCBBkAgtqWD711oO5r+
n6JTUgDRkpOSHO+8PUuAKV6b4LWc2wYxA5zw0J0pfgWygX92pTJNLr/ucC4CK994
QQdHS9nC2XKvuE4WqjBmwio5Dw//y6xToGVB9yXjgWs+S9co1upLBuedP7XDxg6G
7pA6OBdoAugNsDBDOm0kHFS9zOvrsMrNxmLVr2y1IMun9cK3f0TWznKgJMytTiMG
3O3as2SwlSfTl2r83wmmbQh4XOdH3TvG62i++ZfseqvPN21E0unugKFQhz0bEGk7
CT5p2273q+cSlCOMogVHaUOR8KJGm/2UYEd3R5WZqY6AtlOAtsm4VPLz5AWTRQ43
cRiPBCTDOIpnxiLYYp+dYQODHK0hX8BdhLjhD0+TujGs/j/kIKWk1YgEK9K0+DqE
kiV1e0JkieqnIdK0sxXcoGjiugjIwFfvNTlvUcRIy+rG9DhI4uVLcGfSXCF634MH
PG6diz+f34c13A5KVk+A2BAcx+sBxhDvNYJcuefGn8Iw9ttSfRGJ0Erp7H+n8SOL
1DN0sRr9rtrxSVkNVxB67dUJgYNq8MEFifGOodMklwh/eglL7RXQr0H6D+BYPP2u
VFaFjcT2ilr5MJuc59AAuX/G6iQjsJ6flG9gP/RaN8IOoluVb8crizFPLI1S0SX4
i2q7h/EjtiqWZuFXTrqDxwO5JWBU+1xNhXtgdwaCQiOKVOiSnCxF6l0wTd8K/9yj
75Ggvwz/JPRPPNqIVFYrNXS2BJrG7EKN/p7CNp7cu61jnVSI94Zpcz5u2+Qv3ckl
Y1yQy+a3dxbECAKu/jvM2Bz2z599js9zHUOTqiksgzVLuS/N4rTvLcYSJwTPSRDy
FHy+ufCnSUNxNPaZs+3QMZSfoUuzLTmQEJVP+lkmqOroZgbsJKKCeczrUsrqKAW3
fjXQa/v3hTyZAVJ/dv7DzMqZ2cjQdY/sfv1WUlSk6DEA2xom1CHhjPTqumQW2u1F
oZhHl8EwzUbsBrHe5n/WkYJrIcrp8gDmlv1EFzV9KjGAGtmF7UzE3GDyTwbBJOtU
3rJx1cIqeNZJQBdU3kiBokuJ8vSO45XziJVWdZiLlnzAl1aq2/vsSoa6ZUw71yDW
IMejor7bKoWqQIZ6KW76sycJkNjDZAsyV40PPOIRllpG4l+QSl6ObVj8KOuh4bB5
hm5GubAtN5V7QDVHG6tuKO2lWT5433ipw5ec9nvJtIc0eFPjaxU60R7/HumJUyWQ
UQwdlWX6SLHBqKuf2kEiLWrLbzU8DNGlvmGlMlM4k+S2gAkeE/wOEVutH+6rdy63
scBrhWYHLYTvl7w+UI+tEmG+ThjvPk405OA5PvqQ/bChNbjYBXqhY2im4CoRqBKm
dfXJsO2q51tFzxh/lXZKviaMNEW2vNyKEH4W4MTlWcjVNxNF48rlFuyWng7SsXPY
FGVbFqrpEZxBa5/TUwepoOQHyKAAo07AeYj6tmMUZvbt7uz48Bo+oCFzv/j/zOTe
qyjWqw/s9UXhGLc+VIWiNMbBp5I5gbll2HQqpAVNzqeYhz0wg2PxoX10o8GXw1EO
GcKSmBvRNl4pxM7uHB5tibTv6rBuN7bm3eFzGChz5AhRXUvbk6OArH06ngHNmWLa
qWP3MYQqi5Waq3/FR3SrRjYnBDEXudeq2v088FRTdj2i0OAwbUCwaYk4fSdniOMm
52LObVyKJCZkO2+mevEzPE3R8zzkezshUokCQRqZesQkW42KQ91wYxLwCPJaKO5m
jzyl113BRErsgAzyXRVhDE6opZjgTGp5QARlrp8J39ydFe1v4FhJwy6BjZO7MWm6
YWyCgPoNRpjoxqIO9f09WPHChIlZ+panfZkwRAByB4Tgc4R0d9ArA2OL0lqEFVR6
oK41wvfUyXwfQ1IXaZ5s90u+dI//ObxUtflJJ6IkbQyfgez9YMjzvpuMeWyeZcS1
dujp2rMXj1gJMhXu32aqcrKvijZWJE5amzQzj5Xf9U4lz6MFzOUPL1hrlWtEZOKB
gRIoe8EEtLjeKRnQ1OzOhdEeVbe+QaV11fTqObaVhsMhxoMnUmmEWQSkfz8GkWRw
1rFytBIkSlTVxSC0Ukifp7E/hLjAMSA6LzzeqEAt7/Mvy2wbQx2R/1G3qPnIbfl1
rL1KX/K0BdNel5TX5puA2gKoS0Zj7P31c1VQrcaYS+MZ6MMzTFPzcMF9HM+H4fCi
1MqtH2B1sFkMyRSMtoaCf8s2Bo+YycfgssiLrD9fGd70RDS+UFHvJzIOdf9m7cGi
MHuu/rV0JXGukWbFo3iRDxiguPf+uejOOiehBix9KnJmiiYmlEEMDDFiNWTE/WO6
imitXdPyMVZ9eQn568q8e0p6CRpO/OYezenJMpH6CIBSAI3FI41R+2IuD/81thwU
dZTmr/q91MovKmEuDlaFwblYI9OvnutAHvjT3BLp1n/GkBQntXIrs0On8MIB0rUy
6zJbdMBCvNJRoHv6ggg/Y6GfsSovsFuiIHMxnrMWAm/+qI7rBMCHpQ9s6g6Zpfyq
D4iRATWxyiHQF1ymXUwM1f5WPwrVKOWifeoqTIEuG1PTw6HiyDjNFxCCP9VLX/0i
7OkHGwPCiQOQTIEuMo4O8/7b4DISO0S8aqhmBc6AAG2vuoJ1eAip3LqhTEioqAcG
qd1D3ytongeNTdSTuNoioPSb0RxDflpSblu7cc0TH3JTYs6TBo3qQvXBg0ph6BsX
0LY4wGGai0vsM0AhmTfKDgLHy/qH1vPQCQ2g0Lc+yFQk42iyXqZUgIGn70hMciyc
eRqicBw35Uke5p73ggWkqXUvclIiMeWhr8FA9Iwr788EUCip6en3V4CVQggsLTdu
Hpk0OdABYS+NMFPDlwce0d2+L/cu50HCMo3NpLYRir/gvL1oVZMSpMXLrqgdxge0
3W3Jd24tdRd8vrlu3PaDfaUMk9mu0XmENvI1JWG27Kj8KK+Ms9KgQBvUzggqjCPL
znDvPDKLX3O427hAvNgZqbY3UqFZY24s8MfnT50eeXCE8OPJB4bvhT/yK1iBC+0o
SOiCXSLEfnZNDrPOBgWlI81HvhHF8IEIbSIqVJ3Yh5A3DutCm5Jb+/VKBb9WtWWN
zSJhmq9YWlTE/Il5+7aBAL3GpOfFuCF9xCSke600hNtEDYpaWxXQyLukoWAf6VWD
yMx74VWqAePszDO3u+oIv3bkjJcyP970v5I8GMCbjJX65dtvgIzQQ04F8v+x6nwj
s/GGlltYsHaNYMKPJ5i2w3n4FA7iGoW73yF1SFuo/LSnkSJfK7/G1M6E92KsNQb1
rSns/NjiR2ZvkoX624kpaExhe6iU2gLB6EeALjctvR5cnxgkxESrHglKexDhF+TX
MFHmPRCp351hO5kauu0uimQivoM5soti9qKn/aq+01Ur2t1Gj0uZL5OQ+l8w+A1c
1rQ6azlVAuI1h1zT1tTy8wyfbs24Zb0HCAL3K5XcoCWARXE/xpKQTATezH9j2USZ
hYvV8VdfgNHa9RsjKfHnGwxoyXqf9qVx85X7ZXWX0pkVfi/7W27FHxUQVR2JXH/O
caXQqGJgarGvb9gxIoEz6JrmU3TgMM2ZHTmWlxUqLl6QcxwLS4Uh9411LytHH7v0
Lm3acAhxortQoK9HneTPlHN2Bj0whXaOHyu+XkX0hi+xsQc4pQRZP85PiZCI6phu
savcmW10s3CJv4uKn5np6QcKap1Q4U8zpmuA+Hr1p/YiwBbgucX9iyuYuaDNkEh3
X9lUjBGy8Nc7/Ue4cxLrcnKLZsxIaZKpIlUQMFvrlgRPOdcAqpXHLff9CBYdERn1
IGHOdtWzy6J+XOaFbstyY6Td77a/F4GNdrr1KaZcotfiHXde5E4j/Mbjgmslh5Oq
7zDrovTW9K/7ThgJTdhnlnM3YejQzOoR8osfLG2qAOS/O2qEniKB2FUMfK6TDyCK
yw93Xit6zrCNkr/JKmcCwusfEird+Y4qnMJO0Vp+Wjpxs9ThzVBqaIVSlvn1y1Ro
iKNHyNIlVqSS4YZzfLu0daUCnyWTb1GGY9pjIgImQ/EBhBGDYst3gk5uEoBOipUx
Kb2J6uGWUCOe6IuHVzAmlRDEVzlDWPl8Ija4EHEH9gzzv65WwxXiTXcApMB8Ba+S
iQC3VbFgKYaNDflzArC8KLU2yI3p6ewOAzQ1M7uIxi+mtvwrQfzrGKrE4FZeydL+
tORQ1TqteU2QyP7QPXHYemUfeMdRXKAp2481u6yxr/4xCTNwTgYDMmL3LRveUVlx
0+trbpYtf+wsU0zGBMZLodNegUvvAwTenCHuCRPaqzAJkkpUQuZGvl78OvMsvQeN
nFeyJ7oQtELmUeZGgtEOnsvnAkKvrK9mXr62fvklq3nQ9zS5bB3GiyP3ofFJhv2d
DiUDCHIGooxquiozCA6O6/y3iJBffFU7o1n4pmqUkJofJ5fqlJRrgZorOjlZr/qD
68yhFVVGBLS/hrjg7zLshcT+AQVBqjZM/HLZp1NqXSEyPe1JD/+ZQ2Bqi5yQChHM
JIU64EP3ENi/mjJUzkGWZg9SKGcKa70kd+rkENQ9Yt40km2do26u5fFMY+ilv+lo
cieaW8hxgpQOpIvigu74SXrgw8+GOFFfGNVKeF0T9VgoW6HLdBo7nUHvPnmnm4pt
d1moaB/5oyBcDhSq+iouloTXEDtm3qMD3bD8ZE5ir3uzRgbmKMl9rxNbJmYAx+gs
Tdjnrnwgb9vIXwzUBij9afEOKx00Ky2KQ3FRuOZLhbLVGJegzewfgVSqOB2tiqxx
xAPPgr+fb4U8offR3aX9dY6tsobhC1n/Y51jRdXocHsxKlKAw5KHovhoZsyH6fAH
/TTAhTzPFyw1/BwbiIqbgyj1zffapHQ1X+1KdaYfHz8zJWoKHJ2/2P6pWCMaI2Tq
Qz4VMqkhCZ82hnT6TH4ZTjoReZhG0Rk7yUQDt5P+5p7WyFg5Qgh9BmHmiLI92BQH
0c+gykDjv6MQTN/+V1BwwBM5s7vNJkMpuyq9uyLQ8Pw3urlwqkmUAOnVsduwarni
3YHQfZhwysEJYE1+bn6KkQFmY96n0njjhgUXYBtPPBfX7KVzyFiVFJdFC2wXFzAE
DbId7KWxESM2P0OSXqJbD7t82apKiBdniqt7MfaUEEyOTldH9yjgFqkyHo6kd+jX
qOnmHtE/7UNpLRnGG6iXQKTgzWpJRte5+RUucetmmik/ofUpkNbmCbQvmxNlqjhd
AE7KRvjlpjE3q6I3ProBLo88BK9PiRhQu195oog2wTD+dUGTawMIObEnJKtutGXq
EnZmMW/5wvS95GzIPfnuimb/XN4HQPvUjZ5JG/rTLhlyLS0f8izXbuhH4jd99HOW
SaTHGrrtxoRP9jyswMgbzMtpi5S9dxSBOZ3aYimYblpi8hRAMEOVX9zYSt3pNnJ0
BaIdsCtSz3oa3Eo3GxK6LXrMSoVd0gg07KfYCDjAeQzlpx0IFRSyOYrC6brz/6Eq
SHDM8Qi98g7Fwq3xk563znLK8TEJLbqfCuZvwU15RJiulQt7OZm2+wfjx6mYnm+k
9PimDEoIGXzoLLiAR6MobU+jtP6XtRkxCILk6lqJJ4LB3hcFYpjq+CczZq/4OSvj
0joPoKs/EnIK3lOrZ9P2kHXfOHdEf1q4RpIRhjqKJgjIv/iW83maPxLM7gzYAPhI
Tl5ydZ7I4YxdObM4jtbR6c2c+fDNg0meAK8Pvfv92q71nXBQ0k+u7YwNn6yEI7AQ
I97sFkOC2K5gaakfj35GrHmDgwDDXN38Zsr7KGd6xWbNYb9FhrW/SuLvaG024xqp
9JQaIUQndwCjgEGBd/zoOQPEVfjhHgNfsUsw7oMLRIjPHTCkVlmNzTLRVdiebmOI
MpU84OQNL2+gbLn4hhs393k85d/1qxiyRYqbUCYbiFNHpGhFfKO0zA8Iwdu3qtiH
arJl+s+4ErY+dL6V6/xOZqwzUCSw2O5MToRX/VivdC4VSfQdtSepJyI7vNEWRHC9
QgSvhsLb+5vSFdtKsdx7RF5aC+4+Y1v2+oYpIcNgWsOZg6b0awT1DmTXw2BUwTlq
8vwHTyAWpbldgO65srdtmqNIY5Rna/LkGTKu4PoWrl0cl7a4uTulc3hoMFcjSIU6
WKZ+4Pd0Pjx6+4PbwDiigbcHqiVnPIELBtWNhI8gk2cPTBJuFj7VDp8ZXmdHBB2G
VARNcILkQPMlhjem2wewD6j6DcVn7FHAANOhmIf54BUiQjKHqNoMOuq/2VrfP0eF
ckWVZL3R/9MAm2Wwc8xT3qp+gARghzcAShr7IH2PeFP7ycaSTIe8WGRD0P6iGNl2
FLQsCYdGkjafFnM99O3de0rEvw9mGmLPugM2N13VZGO+4akQzzss7F6UHPnG9IrR
x7REZPjWRmHG7Kf4TEIl9avZPvT4pqVmcgOwg0/n97Tb3dwQKFSictkcey85FqU7
P3Hs8LHq6mxTKUujBy7lKizkBOuFIybLVED8gY00xmBkKhTP7CyZ86wGFPL6Q00V
VexkbsPabpOs/PUXLQRxaac9p5Uo44MnHhVYwR11swwl0Gk3A25NWnPURrWfyd2g
sggbO+2txOLEJH4foDIgidp5NpNrbi8uQyrRhY6CGOg9E3e3IJWHO/kT71PfaFgL
JsdeH0F+j4mFt9BfW4yJsqTvVbj7GzMD3BU5bGWedV5Mm5DzOQm8QQVXi1I6xBqM
75CsaEYS3H40r0bYzrpGvMM5w2SAD7N/UYQoUjzavE//4459+GHghQCBUKg30hpk
V0s4Sof4eZlYHv2ExkQGxXPQ/weEAXsexKe/JrGQPpspu+gHCwsyJLIhIgkuTM3x
IoO0Cl6M5XxuZcqeTPlp5GPHonEcnXOSq/PShYl/DJ4HxQhXP8WjzrhF82gGm64e
4sb1GUmnn5zB+keZ/uZYWAIYegvviWHFnfq9UsD0V/ONJ/ShFR8vA8oO07fjqQDg
Mh+reuty6vkGKqfK+T8C8ph4STWPPGzQCwOFA4uWVHaEj6mvkAgPKcWryDEZzVMu
NI9L9pptSMEr6dS/vgrCvrx2TDSfiQuRoE6srwKjxE+LbBqaUZbOBsgADXGxWkwO
Y8QdzvzXcz82to3qhAgbU5E7P243H/B1V0yB0uCilvQNiMgFlMD0XwDW5BnQeGdZ
r2dpo3lZcRSMPr68nwUKJSJ1W/JolmpZ/fX0jRWLnIaYJn+S1UZW+gkHBm6Ye2G9
1pDKSsiy3dA6nsPkLlzAoRzmMAsi5/3mp5FiSDc5D7X1+F0gAQMkNPut0jaFt6BX
BsXeRxR/s2vZObZ3LXnpK4fEVwbHhsQ/x55qOm2pj6iwLWjd99dy4Rj4oh7zRnak
AIap1HRSU68nckxnwePPH5xDpKPXX8Dilh07JsnAm4AxV5ZLL+4hZv9kerK47tvb
7/RbsOKWp/D6fSGDdbU8NLN2SH76b4weK08rCBlLyZhuNyzobx7JEgLVQYUaOHup
SX81rPGDIjLG0qICg+hXbglXiCx2RZxmsWjQ0yFY6uFlmd7VaFUlETFoTNqO8prB
5jnJHB4wU302Z7TdJlbrdOfsegOCGr6HIlvUOg5e0OBx+mLWpz4OOMPJa0hH/LMH
pV+inR7rWmzm7HQfjeMf/I83vp0AxNBaLY6D5TNDprL1uoCqrBafXPu/61WJ5BbG
jwJY/CiETEp6cg1PP7sK5/yFIc1E2UsxEYDRZzXu2p440K0t1QUUIBzfl6bCmBO5
CO4gopaXhu+69ONOdTZZckqic6NeDUEaU1SzZiqMYgdT2wAbD4DeCtIFuXnTjDJx
4dOezIuYwh8SYI1+KaIlJ5Ei6az+83kQEAOj9RXgceU6QEcSqpJK5ZaEoHeCRkj+
lZkUKjrRYSUYMhAjEMnv4XrLkkGLZ5gnLyDc+XdHxOXvz4LgNIrOUA+hzStI4Rnd
SE3mwjifHZraOq+d88ZCGYGOeRBu6029Qd40KUqEAWIqP/bq1iU1mGXfOWdcbQLL
2eACNj0eLCYRCX7Qa9So+3wUvJ3uli3ZOBOE1mYQ+8XjdH6VTIr2jsjlPPzQ0ti6
PzCQNppwTiuc4hMzZNKhYrETLKf12EW+TvQU+b8DPBM1qhJlp+IjUbDG8N9uuimB
gEseJnLYwSPzdSt7qPbw1XjyzxC22CIeMlXHvx8caoVvv14EO2apINdA6ZXp+0Ub
G2oUWVfqERBWexr70Yre2UiUfoj+Qmtv4/oK7xz66KZGnPK3014afhPN04jv1tLx
DagamV2IsyzEXweYxRY68bRe7N42PdK4fAbiIeK/f503zgdh0aVl2SwGxRryYJyB
NyzDjvJ3NYW9Z8MfudJrYjqpWnjd2rFUd8shBxvdqbISg8KZ9lUmaQj9OSn8tNSI
W0EksQvD4maUAqRA5zGNFXio/QFIJL5+VEAFyo3t14yjo9uzTWmrS4aiUHuoAAmp
KT+PaZtDe4Bu8daaCu6QoNIi8onYoDxxNnqJDfkXzHo9LHGByIkRhtUkYc+oZ5/h
5SJoL3ZJ6eWIEcwCWtwu4eANqVkYxef64lGil5bTwdFbC1i2TKruLC7gAsZspZKE
cQT97v5zopNeYSA7A/6saWxXcFc1Cyly2N+dCuK6JKS40H9X0mCbjJVdtaTovvj5
DmWTMmhDhbntG0cTpHxMTEEyZ63WYU2xVEmZKxzw3vsc9osRTuWeQOXLVfw8PBJF
MZOPgEP4jFcM7dE2/ZwUUgkOqJihulxFVZkTp0vi6/zPL7uwtttu94bLKpR/UoiY
mq3Gj+kYw6fxs9hLWSgVkMLZiWULdZ4dNgMx+GDruDma95e5nOEefJ5tRtm6bs+7
FfVGnmxVOroPmVthv201UpDarNveqLQqqUzkQHk4nejw8r1S7jrOxRzSbTvSd8Wz
hbjP+uClnXCuWb0rp6upFeRXvqIjIo0PJrq498cat2crNwTD7o9LYE6EXzkDJ25E
Uy9VuvPg83UEDe6I2U8BbcH1fGKDAZgy1/fCdEj5ylyMtq+7Qs+DTIPVHnUUAg0e
KJ4rmP2DfskMC0SJFcPMXwf6M9fgRX861khoKMDHkpfw4QdXI67D0hc6RIbPBPqK
t02DLpzXr6HtMmvIks7VM0wnY+NJrbjytZPlH70nmSPLqfdXwCw+h6ana68dnD0r
DcgWDV3tLpqMvQa4oSNjcQjXrXSioh4i/gQdumhZd+hcA+okTs0uTb19akbO880m
zXjgQ6ES7lRUe4K4lwah4BuAveA9hWbblAACiI/WGajrO4+bKVDpt8qxE2vu/r0M
n3XQtuUhDcGdkK3UBJnDM2AjhJztbUCLYx5tdYnFW4d/D5Vhikcz3i/F7k9aWHzW
E6FxEu6ZpS0ps7A8ZFuCOmkbR4g0RsnaE5708PjIvbEbWQQhL1dnGnLq7qyOBxpJ
qZRguAnX9/Is2eIAKuvVBNoFjN77a92F4hPXVdh3RR2sMnq9rIuSpnKePXDHQr1Y
I0tISmi8aNNyylxrYCGE3x75wouJ0mT1PWb5z3NOobNL389CfKpIO4uIdLXYviWE
ftIedHwptNzaP879VSuAPbQv+Oz/CkU5dzd3Ba9DRMAxHIICQOECnmMDlyiLnAGI
AUzjRUwZQbONSxc1aaHp2M0Ad4KmKZQkoK+mMAUy7ypZRpj0GzcpsaKjrgMLjotw
V1w0UFhSO8K7dUrlEeRn3PykPHiQgwe+LFrT8o+Vm7EDAbOngJbHz7LrqNd+co6E
IyVYR0oAQj9HS39c6HCYnQHxSwc4WGXb/ElHCDn4pmiBQCIdF7maIWylTm0md5Sn
n+ve2LrgkTGkK81pWYJgTyuAmzMQ/AO18gakvmnv9G3R/fUnm69zDwCc464X2s0+
8mYtw7sGW/YX6cUsQcCUFrYf/uA2ngyCnw7mWCsdEst/a4Iv3R3Sl3MVjf0nheXf
pUG+HdYAh0jWr4mwL+xKxdRbXLojyQB5knGWQ9pskt7jA4Ks1SweegZum23hfYtz
7NZVrKYKdSdjkJyyyI50Gp+MSPS5hpRLxm9+zikyqgFehZN94vrUS0vPEcot0tdX
8XiX8vjpkZ7TTZc0PZOwneB3FWuVwaRuJyNIpv004DvGvRi9RFBjXRT+KQJank33
mCrQy4dBfBbo/25zJfp6zVs07A0ZRXkYak8n12WQreJX9MS31qKM1a4+nnvakjxK
TcOp/zDaF7gthBOshD9Pw2nNNfUilnSflql47XrjyBuFMeAzkASjvstEWyrBB7gG
8rn6K5rj5IHRsDlvHTuY6Pk8igo8v0SW8pB6iz2aCNBEhtPryMCha9IUoVm/SwAm
XamMLEQE3XrDjSngAIuJZhw+aOfW5o2sGx4mCl+2JUpdRByOjXgjs3VU8SyA7tXV
yCfpPuhB6dbt//rrf36mPJtpu1iTvFtIvwLRXsFfyAxcd8vfxDAN2q7jpOHA5svZ
at4ekzZzHz2/RxaNdnm3gjVxwmtihrCDrtc1BAGlwotNU9MsVa/UeasMuFzhfXXL
7IX5hGkpzhUMaA1HBdT816GI8oJGXMSPesRzuNivfsDcoPhKAoP7cjIlg4xyVzkl
rMGFiqfT++f3XKECcYUL/AcIQQLH2Ewp4wQU3T/8TA4NWlejLjO9W2zd5cP2jnzg
zfyOCamnQyCg8fSKPjgOEuvHnWfLgJ4KegFzNZubWkNfo5oDUHydyE5rDktdsCoI
OkmoiB3Ho3ALZjsaOPUIzrm5nqLlZh6WoBlKZxRCyjdpPAwVzOUlb/ZCkWwSsDw8
sUBD+xE7ncof580Ykmkpp7VvE2HqAJyKmgnNPPrmfUsTAPawLt8rFS1o/tOJSRBQ
prKUvEGCoNLyVRn40HCZDpLc6q3NfP8F/mvFsibO15i+sz8duKod7i/Moyp+VDc7
RT7vSKrRH4EJa1qZS4ONgOay7kVCf+TrjYC0KZ4QNpZtI0+NU0R+/vDeGuzWm3cN
5XhTAKCAqaCz1HDMy18dz41PZvFTydfVkWGjNL0yUGES8DExrNqz8akjmjrpR53+
QdF82F1WsM9f1zDGpbpXgHNrnHsHP5fW7VVyR3HVAhytO0VxD/TBXheowSJipW8u
GdBaaXTCU1ctA3wOG8RQq1kS50nvn7ol578rjukMCqKVUdXJc+H7uG/e/O5vkgeH
65mPvOmGSl/bFhVFR9cUh0IcTHs1pay/Z3KBAG5Gw2cYeeno+0oSMxG40iGx4P1g
yWzXnJF7pIWAhFR9VJYKrB3tPIMe4JcCpcO6hYoqFjFDVeLZ9vMoGuAP8QBw0gI/
dysg17PkShKuMRYRcCiSfRwgSDW73PMrR1a1ekljsm+THEjMEqZPtOxYDBvnkCGg
ipQlKh9gstFYMAkT3YOLR/sX147tTHeEOuICpkPRwU7ktGdb+nYdsRm8714zY96e
MFanFMp5hKiWsCqjOH4RyunhiLJeyv8IMNiMIuAgLjm4SPGdyiI1mfRQ6us5WkoR
TZJw+LM1PR5IgdoyXi26FvIq/aFKrGOd/8QIy1nqzN3pPlVJ7FEgX/wrSEXQWV7O
OMQX3H7r8NJzx8tIsUdjFYlKZ4EwestpcOqoDDPcuP8G0ig3dHaHATk2UB76pcmC
rYtsLNt6DkuWn2KzYoQaNgg2rgqW4FXMQ/iP7+sknI615xX3Jws6XujZisA+lZH0
02DJRlwEEyV/1SqCFJOIDRCh9TSDgwjLAylNRYr++5ivk2JOR7Upy0fIQgnXUP73
I/60QhP10QJSMvy6YbIjsixG3KmRfvsLtjSyoXSH0rYkNp4EqtAgJVTjWnjeB9Ie
hW1aZIVK2bq0ZKzNJ9Kb0l9l3jptCReNXTAQJykqpS24qbfmSas1c7Qx0ab8K7Kk
Q5KGR6e3sAneQgMoUtZ9SMX7Olyps7H7pHF1xpNNjoGMkqBhMk6wCrPoK1YqCUbb
QuHL+bmriLf4EkmrNiwZLFFYxKJ2ZvK+kn6qnfhoOy95Iu2wrXq3Bw48csE3CkuX
Emv4XnzRFtBwrdPsj0aDpSp9WuVuJ4JbQRZeNhVrQcAGl1lHcNgvq64VifqB5WkP
WBpwEhg1IRD+otF0xKZDl+xvWXRQcm/GJ9uG7hRlI3fovVrXd662NWHd/GXL3VAD
Dri5lpy85004LdMhpOAY6l3INEiyonhc8ARkhey39GcsO6Xs1f+JO2lACS4aPy72
Zi2I1ppBy2SEbhnFE1biOLkt1OV7yB+6dVjPjokZARVEtFSxfUrsUggTY3tSrEh/
gFc4KQ9cYSt/SjTBgXiHPhQ/s3fgwXwxrXJfNWaCjrV8li2dfiRJG5B/pS3EpdEY
oawy4bK+wPf6pGt3joqNs0WrWPni4zq1Yiz3jOUdDN4xQUIKrxXCGqXb/+XX7L7c
BuGIA0LXJFxA6CmvuYG/AMDkBBQvJGhHYrDLPKuKeKZcdBykmtp5oss1YGDcvETP
iOZjr3qo6URfKTom9yqtsot4kpmpdDMmMKIXGGYOk1UrD8U1IGII+d0ieoLCRQHj
ye9MdUuFRd2hKG7exIu5iry82mUAsnKZbz35kCrO9SME2rrNnjkSDHXH1Z9MUC37
9AmaR4g4lIpKuCGLJGeH+UAJAFuvAnRBAa6K/Jff2kskBwjibFadNntLnzHB5onS
eSDjnjSUuTVceGxQ3t4FqKORshUjLlBOrOl850fIvCwzzlMnICX3Dsi0DuU8+2H3
7Q5jqHj+rZbVPCeDWr2NawR+OoqOtuKaNs5pKJVUhdjSlcQBdaSRDO4K5bwR5bd3
cApHo0mE86gT82sZyyumCQuu7Ruc9BJN78z/7ytJ1VGVOzj+b6+aQQ8Da1k+tJvJ
w6v5I81C++8l+M52XrQ9aQ4U9D0yNO855IkhEm4cEj3H5dIGWlvJclYfo0RzAW/J
SQ7aBUT6RePxo0AaV0i873l2mGVWeCSRqH1uYcts1rymOlyE8+UHrDr8KBkBfDst
HWjWmwwMbfsY8MDU/puxG8b8Rc7zOvrgt+pxcw6NGkVrH5sRdLUrYwBcYDv4+dC/
jR/3O8NyjOYCI8WJ5lMoqn2yYllqN+pnFAb5YfQV2g2da4hyaybe4xEqEDojGEeE
uKE90QaMTL9BuuilGfJlzSLurh25ImdZgKZvygjF3WHasduKme/gRK3kv0EX74MM
8/59f/vwhUj1wsknv9k2hj1jsNMXKPKVTCj4Sd/xHZ6ZlU70j2HGclagIi/sTwgZ
QTfJF9vKwLguDOHc4suV8W7osy8+jAYsvecNwmzxaoADRi4TRzGDiGgF1cOiN/8V
a63bi2v/VuW//55rgZfWvh3dI+sL55PL977fPDbLufO2N/aD22WUXq/pxZ0wYuIJ
5RWHSGIpCGbHnh8+qtcrpKfy+OkUZyFz4Uqpxmi3GPVuRKAHRR03to3nXELkooxe
+yi12YtSWOTcaO17/HG3/tz1IKqeB7XE7lQHevkyTXHpdqUcMRBqw5Uvsg/MVt+D
Mm5ea+mf2FD2ivPgGbrApG+nEKhQZ4+xuTKX6SrcpENlARbaW6ya8bjkDAtXHK+c
zFFXM9GHfu2GoK7MKT9/dIaDSqJSUNbjf1yRAUNKkkEC40klnTuvf5dHoIGWY+Y1
PawweD9R6umXLP75fmwgguSMGtHJM7p/oSEFSxssyJlzw+MFVMW3Txh9fNeCfpyK
nr9cANgAJNsPzyahBR4PJ1kZ6C2llOUAuMi7/90rQcH/4HKxk2CzuC+uM1RUbMMm
agyiCK3zyBEhm85yrP6VwdECLxywkbpJ47NpZxKlyroUj2bPJ/LPVixUr0Nv4Hce
AFn1c+cPeGpUJZ5RaK3HvjW7+iZ2gfmmoT9ODmJ1IOwf6fWIh1KQ1/f94fICzZ7D
fE+On3UgZ6dXb34z7DY5ttHAw80Q5NHxcl9iplm2c2ahIJ2vbYI7s3rak24fqjUH
DSfcrpRIInhhnD6WIE17dsfPc1QZT6pogBwfyry5M6i4yMjujvRXEOc9PdyLHYQc
IzzrU7um84VHU0svOfO0QlqurUAIQYBOLiXQjjLqjQ8mzlKOBnoxrDadafjmFLXE
KJ1hg7xil3TgiecE5BfD+1m+j3gZMlzxdJnCx3/xz6HhEYxfS5p/gm88FfdmIpum
jkszpDZmIMmDaxQUg8JYg/eGV1A3da0CfbjOzy/ydlk9U0w0kzIwgkoQ9Mk6nfht
21WGeaVzCVCYdC7W8am63kMrVjA5tf/dZzWIbwRUrYHe+wkEq+9mwnPCITLS8mOS
3CVxz59F/bXD2s4Gx7jA0f/jNqSFac0OeBRq4PkIvZvPnB6JXkt2/KoaMJjHyoe4
1juhSCF50Vy6+V6vVz8D7HC/P4nz69KuN8peSAi0VMQi1ATiL6YKKpE1TMkLN4ot
pa7LzVCwoOl3zoXmkB73+mh2hfUrQw2drkozGKFHYAjoUIsgC3yJSo3a0ibWEeUW
AhB5Ki7zFJzk2L6g+pyoUBvUqBk/ke/0JMyNBIM/d/OPPMemaVizH6TV2ZNVvYa1
d7odFFK8sSwpWJ3guMCGwAhbdbsaI+vuLSPsp5R5lJPbzfuXbppRu4LwsV3hS1fN
sUJ+uIjHgY3qIkSMFvkMrjjqa7WsOiT/HdBkxXCYCWIM9mxgDL53GDh1SzgFq4ye
paH1muzkZ8tilyjvryjxiVy5vI/qVMitpkIOem7y3UwhBV99Uh/2+0HXlTjzZnav
aRMJeuG/Ubcai7q034I2/XJk9ziMa3FUIQI9r6G6PfZrn6w1tHIMAjzy3ftkJdZu
+4NzYcCTfH9GK4y21loA0z6SZ83ZsnU7g9OD0LRzh5b7yna+YE7xLX3MeCujpZA5
Z75bNvN/lSYPZI5gg8tX6BXHVOKLw9TmouH6Z/uxibwKyd1FFZBu2A2oybA6sTNn
xA8ZNJdDoVLmRFICx22p1yXpPo2k+MFhj+ip+N4qEbTc4es8hN0lcE0s7V2RCAS7
hEQVwyVcuQ4/byv8qXfUFDyqH5U3/Dj+JBGLakQ/HkxYHpdx0Wu18ZydLSAEtCZp
Tgxg2SI29zPtQ8ACO42upoqpYPAoC0Yg/3UlDZe62eQkMMut+yvWUli5xhEBCsu9
eqSFUcW5AeL3XxxhzSINlCkeokUMdD0ZAWSGfHGXUx8prjHZvF7ce9J2N+2INtZm
N/W4Gj1EvyGtJNERL4Q5sN0wu9Ys0/gNzNPKoTYqtjMVv23FpGlhoZPn/qeYayrF
BF/IycM2j7PwSi9uKMDNa9mtmebRNBAWi03pZQiv1XetpY7Ba5T5I9gXsNj0/BQj
SagP997oLw3mA08TpVEQCJzp2L79W8jZ5RXM5zbq4UEnHIMzgf9oazR6HR7mBY0p
RaL2Wo8BXWk/ztlVG6mQSqfvQ6Dc4HIhoFsdrfkUkm3rZnV8yb9NMzxjXAa78MH0
plmiWGrw6k2PT3+8UI0BNwMydN6SmpFTLejPljS0dqerqbrzOyLnAcApjPxhPUqW
rXIYz9SukL2KGx8jd8q629BIcFEtGNw6ZDFkZexQZbX9R46vRe08uEgJandWgw0N
tbq3THy8Ll5cI1o4JG10sBR5uuAkfKXoTuOCcDYqluExJWdi2KXM/qjkcYFFLypO
SylY1/tfUQa724SAGM+F3hSjp8bkjXCh+PULzkdq1xPzvHPqyiFRGI6M2qDQk8P2
K3c50qTqoDYJseqFrdnb82BCIy4yziI7hLaoliVg09jXVDLt7tsnlwx+j07eiiIK
amorOHSi4XOL9jlfsxRUQjb67dWsHlof34U1h3yIapkwzsHG5yJ3NRjTz26GG0gw
nNSCBHTXh+nwFWR7jt4FX+CEywVgfh7V7ayHpw+aWBMLKpljWilqCHTIWzinhY9X
VDevhTaBSTFjC4888VxyvQnu6eLD2K5WVGN4gcuyMQ1aSYbBKtaazBS+etqBKgyZ
pMxhDgn5om405H+C46o02+hXWduN1eebEQMyhC8VXviQSe7VZeONaHD38Whuab/D
eIqlAXDU2LXj9T7BxJBjDgDF94jTBJZklhKXc2VUXqaeg9mwM9K+uXrUa/8BchOV
QYvi1J3MrSIETaw/5htlgCyzvEtapmFj7ZhnVYJJigflK60rhapCnxbbS9r1XUpd
lff/gemrQvENv1nH29sTN4c5nKTi4BVCsDD+78wlMAO5jMdNeTOtP/6GxgZl5zGP
B4kebywM+XFq9NPlsDw2VZ6ihPp/Z/VBifSqXNoobMigCcsfawUFu1i/Hg35SDBD
BrPmA/TLBs0Q6hcZThmIzifXpPeY9SHL7KZD6NrCDuGhD7yeqoQH1xcIDaLFjMuR
JqD2+XXUtPRebkXt3ELt3ltXP+s0OSi+C/yULpIcfWqJ2YJhz7/Pyv9BQpxQyABw
SNaCAsQvtaoeoL5yBaeZmBoO8lNGTKP9JNHwalc/9YDD2phO8DQiUR9XYrg3ewap
eC1AYnFe9aqJAVHOtwNa0RzGJ4I1/U7F1UxUB8NCYRPBz8UG6SkeuNSkHeXmpMIu
y4etrX7UvKCL06rmofZzAjdmOERhm2sappWXNh8oHQfctQDds57yaSl8OV3B869C
jpNbGFeNkdkD0b9dmaASgOqBhi26G21rISRLBRclgQyPXXO0l7t+se5j2NF9skub
ektsq4IR/6+wroNMPXy10ukhciDcEYkMRiuufLTg/CeqSCEJSUOCfY3bw3VoWakB
0FEOPMuJFA2qs0ayIJo9LM3n8z+J+yf4i3cZO+8pbGvl7imC2vvp0ILh8aBFE+ey
u32qK/Vv7I1tDJKYa4FkAizaPZA3tjgIUpJ9RY3yLZYhAErpZaCfz0jVVnhpoufW
4y7DJWrKXUYmWZFVXDSavzeiUL2gzQhBk+G2gsl5eXRNpRPvrPmKdfaBjtPvhpAC
LFhy5JhX0OtbHf3tQjlTi4Vn4iUkt+PLqIefKc8V3PbJXK3xAZIGbMd0NQacaW1O
sm+C4gexIkbq2mW/4VVOgiPE+b4gjyUb3pm5mKzQJrPy9jOVPlX+UFdLregBTJUj
vKi2HSvi7wmNhTtb7JGK0f3CwO08776F3SbMr51UcpQaqmJ9tzFMJvxGctklFVDc
i4gpeeEA+iTdJyKmXXyOGNysNEDIiOejOpZWVkjNViBFqMfXxvS5vqkW9CQqTYK+
FaE0TTe6x0x67zZXKVEOrf5vlJ9qULnjcst6pbrdl4KyoxcrSe1L8gzt8wUGDPc9
GWL9ZPi+m6Q1eB5jGk/A+eEejQrG0CzSjyydDMccENlKCAwiqUPpyIsItBCad1sN
oFIvPkXNm62pwY1LHjp2ac0//6va2wHcaaO7e2t9aEaiuyRQBHR3XOJ6LHC04Nxx
M+88+jiCUwERba6Ni/iYupnuIbjiV9gCONytF9ojrjlCwif0A2NhacMTcYWjDj+V
5G03kgr39vExL66wHu8NDWhh+6AqL7Hg4xJX9Qa+tIAHKr7bBpiWjGdOuQAm+9XH
vHn9ZVBz6YNv8olU8fQSRnXMfqTu21dd60WwS4uF3EtwG/6nDXHHW9JwCH6NQN3h
J9La6j21HdR8q0RW3us1pgzOOUgM6AFW02K25+L1N2sO1yFiuwoCPU589jZTDhoT
OCP8KYib/8Ds3BAAvPjk1iciEIrbmd85aHiYvqcU9NmjG6F5G5ygl4Nwl4k/kPW5
4ccMHNX197+4Bt3jA3xdm82Q2Vh0DKck60C/AbxoZyiVokyE/NFtPBfrCFsjY/Gq
U9dDKWbX8Qb08dtnN7tfEEev8b6Lj0VNOlLx8fWfvpvgJUYT3CyKspe3w0aEQu/Z
1JfI9kbM75m6RsJJBNILaplvBkVYA0MwhYgJcqaThU+5LruqtRM8hve8erarKnYt
snf/XRydoB9L8ruiA7akKQiSYzMZ5erppapnnFp9v2swhxNiS9kEp9NPqf8Tqo0B
EfOkoYibG/FK2WXC6g1j2FICndFSoY9YTyH33ZUuvDosE4UMghYIod/dOl0RCosh
oD/VrKkoELUqpmE972G8xTZSHjpYq0FbTtZWlUx537atk3cPpPz8ONvV43v59883
Z2jUdk1PDyr/2Ysfit1SI+bZcgNHrM0qkSfmHuu8Ew/A4FXo0kKVaiS9ynTxv23K
lJOBiTSw5XEb8g54PoFV8Jw7EoUQw/LzimeUfsgMMjXwrkchJBeaiy0uDc0mtjeQ
NZTY+PX4QIaNcuwX2opitAyEAueODSDfVrJnJgDbN7drsAAG0ZS2Raln0E8mZzqt
+95b5gFLfluzRQuNR3dZvFBz7ajxak/dd2/6GBtZ7QMhi7OKuwrmVBq0XUZ/Uud3
2aTDIZx8SAVZIeToHoGtab0jbzwlaTMP2Q+WctIhsMLDraDBg7sEPTeN7wzRsh4p
JGi1OJFl4tEwQejQlniL29JEADrklYp5ZaJxHblo3+tDqR2uC8sbqOrbBIeyfUqq
ChHhQdId8IXoaGfMY+K93xvYu3jf9+N3s66F2Xa1APp44TAbEcGAVRkNU0aRjLUo
WbkXEWPPKgqadEXEp7SZxf5FiJdzUDxcA44r5tRk2fCwzdiQa2qij1cFu6p8frk3
6cMzQgx/AjOMrfn62Q8NHM33bhNorLYkS4rIgdJMhM6JjSJdq/4dBVjXY/HQTPwK
hzPZn08WMFrnXzszIKSnk6UrvGyAqQxnUFrqa+dj4d0tTJSS+DzPZRUufFpeZPE/
XHcUxKTLw04g/+gFQuxi7Hf5bUvafrQb3oVAnbJWffEPesBRTlMTKOMmSrD507Od
usLe9bdYSEcKO9uJBgH3ThrKtWZxQyt2EhEzyNg14coV+3pu6afi17MO2ES87C0s
0vr/EEBJ1OQisPjr535tN1zADNwCDMkzIfuQC7zRPygn9OnS5sy0Si+YSV5kriQO
Rd4RjeoQcu4Bp/r3hlQ2EPnMcJIG1FmuMugcP1XsKF+6fBOezqmyRhkpO03SSFbq
awFf4RQhxZMqvzJPCUY8vk89JAHrrzxT7OtjE8LZ2FrZqUkssZVGrruRaAk2lEbM
jro+yWt4PoHVayfZlNQUSvQmnt4QdZl0Ec4opv3xkEU7QMHLeKp9xIRpaF/XUdC9
ADihSDSKd/GrRZ7El+tarln4/LM7pkM7FJu+V1iimIBqOTxXY96nkWO262ybL+sE
KqX4O6VPuqQVzE9Pd8w3LhdOOkawzWOIIwTHxL7eJdcvg3VLM7GX3Dwd/7saZF+/
tTFQJYenZjlH1HwmaakxtMP/sTsgaxHpnxhaAWFptuGJivyg3cRzXiWQqyFsAm3v
3k1jBvhmI+KO+4MJqw/XMQ7oYN8DSMa8kcjkphIos3T0yAJcPhNbcx56ggXk2Sj2
IFQBcTV/KJA2GtrIm1rh2vr3+cqUBKPbRwRGGkmrS6GUukLnw+oA1iqKC2h0IOst
WuintyEhthapPnYAV29ontSk7ZK/6SCoqcl3cWgzgWJ4d23MAQBEtHbO2kI33gcB
aZGrRyCaUz01Vcz+CtSmb2Mtza5E1Yd8hJWky5zyJFKLhcmFT+b3fDkN8DaL92LT
UWUXZK6dO3LXK4g7fGl7f9iT/hhGQKc1GTxRrkwym1JEvLOkv17DHthafQ4Go8lN
8CQs6vuUhF0IqEqxuf+4BXMUnvwQq5ov8OWA2q6h7KrKMfDCRcn6mhgWRn/cWtCm
BHExLeNrWqXFaMchZuZuQBxUFmuvuk9TRV5HizHCIGZEMWZvPx00mkH3xCbVXdQn
2fDqEafMg77xTAOW8gcissuy73wTXM224o7OCYlTZ2+UJ1gtFp1benzQwckuNoBr
tX1j0AewY2r6ctWztqakLyChCUD2d8g0pO+Bidj0nmCfMGN+uV6FBBu1jjO9knlC
QejSNjchRC2Xf79PIL4Mt6JKJhw0tSOp2IrOMHKx/nKO7Hm9vEVFKv9jfUiVnLXD
kCnbPIyKH5wEWFllhSdbTXusGoYy9nGG7agG4w5coxg1uhWKh0olTVfiRfLL+36x
bLZj1tFjnuBsxGkeq3OU3GftGVaqRSrlRLaysNRyJcf61O5dlTdJb47qQ9bXvOCU
+AfYkjfhNABjSx8GPcHpPAbIYk5kzGXlNUo9y1WBxM4ePaNeiLKZ48q/0eSnWgRl
6QpFK6jQF8z1PqfQSmCUYY9mjex2Auhfoi2MhBap+TEqV4PFTJjMG46cO6Evwpgt
RnjxLPo6PApfhGCBDAxvZfwdgwV8pIo6h0r0EXvbxpkOmn1SoeBCTzK8bFCqNntC
Gy2r9Oe4NBoqURwm2Yl7zBoEHdGIFZQiZoiG7uhIikbwvw9LpgFerUs9jSObXDBP
yx8ftBu9jemajc0jDe+jYoqaQt2VNALHnvaNJGq9YwQT/KKgb2I9RrJyPYkkX5Wm
Um0kkBNPXog8nE/Rha35M8QsUbahu62ZMLLWvV0kJysmyHQjwCGstsIgDND5x3qM
zpZTEIUNP8fxzwTwD+/sSiHYVmnkdCBXj83x+NOleCLoLiIlllcMiYMRqbSnIeFf
xEJfUImPjt5p9FdaHqHn9/jex3r+JCJ7DlqhbYBvpbtZIN0bX94a9wCR2G1s5Qbr
irNszYjCCllfETL624bc8pTzhj/T0kTWbuxSnfxoWiFnX3Ei85Cj6vrp86ZxZl+m
kjGk2EnInXtbRq4PGbeqKrQrusFIaIWUu62kFqFzJt8LnPmn7QJSHvi6GjH2z27c
rQS03fVVhbEF87sTyebGGNd/OVuW2WbNc2Mh9eKYGxJLm7Wk8v4pRp6TZqsOs7AJ
+FMiDmtKBVQPLIMHKcuJpy2R4bKMvybxOAmVbSA08206XZ0x283VqaMMtGaHwP2G
KWwHyW/tEpznd/n8/msC0yrM2jOogmWwmmS/1d8BQvo5cSbhStSGePJAuvxkhxef
jCMHdeMMtSe5B1OUZUtmJ09tJUTQMKiYe5FWFaVUQzNbArZq0iEzfRLrT+RhKSiw
NOES02ruqjviD05zXMWtGSGxe+Xf5M35eb7QBOWshgmOreS+9RiUonVgt5vnqhSS
pq/qtSvquHAp+ydNUNT2ydtXWkVUCEzvIYrvmscnDkCr8+2M5lQKiilSOeU6Di2j
S6QGX0UusZTEd2GcF0nuAjqWUcCTda2b6e2hiqmL1HzZLmDaDANH2+XxLUcSdqcL
/yVRKZ7t48APH6gjc0NFI4SNuHqVFcpO3qscrTZplCFIH0qzAeXMaSZ6F4RLDm+e
yUTVnhUMlQR3+p6xIu5De/yzDqQeyRsFOjGHagaImC80hoNcF2XNUS47ZCuWbuUN
DsZ0CNSB72vJwDiTQkU+cov0v1gCt591FFv3cvlOKaelo0fB19tqcL9kq0uICH2l
kTDvz4pqeVz9Om2qC2FlzT9hJLY96jkBXr/9tAR4h7UFGS5RcRENYDzHfvtO4lZz
SDi0g2wJVTVYNVI6Rfw2iPv2yPcC+efL4dsp1wR9MszEUVwyIYePncM4Ghz/tfVJ
LyE01ZBKquMVJvZEuvYnQhQOLQI0I/6uap9mMclFXYiwDETgLKJbigtZ/ReXTy4l
Jfb4adc8QNnxGr6eHMOs2LyxVt2ZudWFO4AO0TtwKBaG58CU9Qdsnw5esDpl5YTn
PWwiL9oKfBoKY86DA/FZ3ZolXI0aShks+WXhSB/JsczAzaVBpAZxp2+VefJmG/Hr
C49liV9E3B2Tu6TaoHaP/i14VydQqyFJzqgrG+86X4OIi2oOOocedOHlJTQa/zgx
FjUsAHbDO9BasmV2DgCX42MjkpTpjcL6LoJ1fOBzZChSHt0yAvzuHKFw1wfox9Pt
9DSV2jRIESZtIhdNhX5xrVxokdbW2vfhc7OlanBk//Kcx98jQFu7B53MLXBzSQ/K
2Su/mgmm9qyTOpqNzZn6D/NWoaCsBn5h7Z4ZlKilvs9VF85+QIZ98j7rjkHhM+yh
QYFQuG6cAsolwfUGrp3AVR3I2s/YNRVyQ6NlxQdRJ9R7ad84syGL2F1qA4+5W1Bi
u8oXXlICpPEmpSVIRGjpV8+BW0+C3MmEVNg0GltAqG9fdEdW183qQdoe7TCH1rW4
A+fUy22J9y68U5ljqeIZC8tZCqkLh1sThPcNbrf6E8EOtL134RlHQEyETURnmJfH
VhWCBS7JCQBE+pIJLSgEfDBgzBePVVaCQSsU2pxLlr/fnw57bP2F2FlkiMzG6LKu
9zVufeDE+8zX37MLFOLtncGd3D5/VWX9mxHflNMLQ7jd8xouVl1LqhdpVh80fNz9
maXOmE2Jd2VLXFGu+todA96pQsd9pNppYCI6nR1Wgqe0AwBe++LvzJilibLmvX5H
4OP2+15oKWuh9okTw1n8hNHZ/jNo+JIxttfHsaSbYIBqW0E0QFv8x7lX1wvcl/bQ
SpuhGUhl11+K5xFh+tborKQfIF+Da14gkUDNMZhhRe/CpsvhFho+49SMkpq5BfVo
4804nk2PfT1cspyuNE3CMjVod5aWRsS/N6Ln39ge3y+aKZf4vTAqbAq/JgffJiu2
gF3YqhitfGFkfBKkC/Snij2GMHpOIAoIfBNYK0w+cDduh6pd0x28jFpEY3CK1W9e
sczGnVf+6ecC1c30NCnMeCm2NtejbEXjxkBAXqXjfZaxLW7ecC/RJIDIQb8wGsJd
MmhqO0KRUpRcTNMWq2J1GHR+jpqWDkTHQYzjMUxYk6JyNoqok1IfQzpabHUl7WlD
xDvwceyYpyc4oJiKXlgkB59hlv69CauMomgHbQVo8zdFgvNfIy0HlwYzdoueI1Ob
2tX03HVs862SHuAz8dmJZr6A+LN4Q7Z4uOAxmTxiGFBHjoWkpIlARAsAep/Ls6ya
7+SYlPGCmcj1Ff0X6/A7lxRutnEQUhJVHVXVa3YZFe+3bWxqk9Dejd7BZDWVrQ5N
fJGQ31BqjsEa9LhcGlC6CSWMRl+XxyQYIjcLkGQYGZRaSiEShVDqgWLAIzRmuzI0
O6sijpA6xRzX6yR0CJBOulxrjz2rguK0b6vhi4ZsVDxl/xdhzXKXWb18b8INjP19
X+0XMZY6LCxvv3N7w42dXU9K67QfBefGt85eyFZw/IxtOZWplGWo5W/VtRo47EuB
fz/8BwNMcdieKAuj6dbEGWqN+iIPL+XTwZyA0juvviVEmH4ObjVG+7Nrk6AujHCI
Hff5gRM+VQw0JwvgKAzVa+3cpIrZVetYh2L1MtrAsx/LHYRzmwg1105slyvgOqn2
IzPHE6BqbzHN3HGgOi5/mAR5k/d8OBgsmWFRqZdCLqzL5xQy75SbpFCtN/NtbOoK
BKgJbO6o7LFsbz9k9BNy16+PcGnsmRvG9rMSXjg6Y23yLaoxLwmYaMM55qelsCID
yfYQ3I6OPnjkHPD3YrT7aGVlniMDii/05u1LuelZygShOx6nCDJ/rpPPF25fDDJE
qyInMG4A1OGz0Ax6Rr2Pjz4nstIvesCKB4QEX8EAw5RCHi0sgsTuyEY9gU7fr0Df
HbudelNYxDLNGayiWJMdgRQmNn+XnsEqenxjM3m2Q3Z8C2M5OwqZ+PsAbcVhqbat
VaHzPatnPuL5EnOayB4813nWm4gMLlRjdXfi8g+voNnPD4etB7myWIzR9ifP9L5n
5bPCabE27iMhgns6yKHNTgeNu2e72LdwkTCQ/5Xmou4HPhV0SbYfXxhcz6Q3uYk6
/cRkmujYr6nxdv+5x/jwP8fFCisZXTnNrEePChJJfuN+5DT82zqGzGx9LZimM7ai
JN3WWuKOi50FO7dwfwzXmEhMGSafvVqqNM2bmh7+ulflBsvrKnIEm5/PAbWgqcLD
cvmF2JkLxZ/wDr1v4ql0MJd+txtXK1POfr0Mh0Ej7ZzWSg4YElKCRkekxrzXP5zv
TB3lvTby3Y60lGJKHX1wY0Vc3dU2zfq4VLCV3IA+nSqZ7b/RoOx8hmUrGBufSYIi
ZDSQSo8/R9nerl1X+6arNyf509EQHJa3Umex1PhnwbO78TDnFgcrDAwOuWltX7rQ
PLFf2kB5IrdeqBadA/NO+8gpAhwVPCctzFxzBLol8WVS3ak20hGSI9hculJERlpz
eEQ7ETLL52byJMVCoglEs3AQHS0rlqflP8PkDETcp2TM7k3Ee6u4W39mvgFlA8jB
9Hiq116ngN12CuIf117dDub/CLyneYCgARxM2iTANVNgQsWsKPVwQmZUXLTRL0yE
uwEfBp5Ap38odPBOEh8oaXogcq3sJI72UeCasvnHXT3UrZZPyccHGUFJdbSk8pfq
khbEV0ic0PNKEMT/fvsj9HV6Rk2V5NiNWbTIrcSgAFIjHubAdsB0dELgZPMVv1X0
8YX5Z42P5t6V74XyliE09jRJZoUdXh4LTM5DkOPFz/4DdapMzNOgrF8Zdzmbk6ca
drlIm7isdtOFerT8ZZ7S8plka0zd07FUa8l+uc4Y7jAZ3m7GSp+s8qCeJoifB+w5
kZi4/7/gOCF1yxoGi/UYSZlFFYS3+tih9XUhSmycnyxR6auyimtoh8DXux5FPxRE
kQkewNEPtx8BLnaICS/hPqnI2Jd1rlqI71xpHDpvVkmt3PVBKuHESPhBA04DP26K
GmpykYB3qOBzdz8aFKztH1ivtw+q7zdy4cFBDKEwHSrG1bSVD9iEno3TkPveXWF6
SiHMuxdnhIy8LXb+n2Nku98VWWPH4tH5H44Pa4Sew3/7T3s5eo7ATav0ZgabFbI+
rO34Af8h9kh70wDlJZOhUjk92yrzq5CqfHSbR8UMqAYCj5aBP8kznDFCXp06V4oK
2Js/VsbSfSAkvZWuEI535sgQ6E/oohqaes30WpKjc+x6X4WrgBJbXYCtKkJ0yF9n
BF/bz+1Oe+pIuPaP+Ylg5NSEl5Lk/UZlj9Hx3FeK2xEF0n4MCykRJaORFTt7PAH8
wdo0di094a+RuMWBpUgQgiQgS3AUnVMpFulN3m/JifdW7+alnXmw9AO4WxkSoOQl
Ls3r7Wl0q/vTrrPuMknEOytPS2DfroP1nu96akLEq+dJwqyv7upf/tZSFKcuPvxd
WVyTS7Ov22M9A+NTrjClBlH94bsf9gP5V1NnZlVzeiVcv3IbBUHCViIO06mx+9BX
DBUslLlDFlArQtZDxiGn1ef+qrUMtilwG4sUa5KTNxjN9rk3dTuCaBaUckArJ5dw
r/YPtbjr3avzbYCfRH06OaoJPlK02WJ32MQNbnpKlL9mxKaC4PJsgbbS63VHnTYB
68x/RvzNtGmueVS9snheEjnrG4p9jzdUkxs2qvaTXU0GNILMqFj+GDaa66o6lhoq
AALvo2cfeN/sWggVQiQheoF7hMkWlqJrtkKdWdgPlxTPpxHZqi+pvEMcD7b4Q9EF
q2lavbKo1BMLoW8EVr2qIg5oKHC3VlJksSogyBcraXogrK7VH2BGp/UmZrCv2LR3
M6r9XLfmIp4Y1SN4Hy+V0v+Q41YAsHEPzHM/CKEd/EXVVBg814Jm5fZfu6wXEzVg
OieRPblxxkmR5YYh1j0yK9FbS7zR4Vx9D2wIhdUSIlc9/ggO8zFTw7dF5HASWHBJ
IOUq/77PYbqFo6nvkX1K3HksKWYeyX06vbmDgn5BXGW4L6a4u7qX5tSxG1fz+jxK
q2lwvf4blPjdcKLIZS87tBroEeyCcDYZcXwL6Ys6VWdUQf1xl/I26IVN9WVEyaL2
zuHECM80myPTTL565gE+qyPF6psIh9az8/oLa3lMrFiYPJ7WWSApOUFMOj1+59EH
vePqwPNDeYoss7LQywnPhotArg0AZc2BeHGsI+JFIOMoBcqc/xjAAIlqMRUQJmfq
DcOxw7QiOI1o6eGyevp8sW5wkUfGY3/g48cpwoAxbhrQIIJAh0djKob3gM6cdCZy
I18VBFmgVJT9MvHBR2b791agd+OkNniFolKChcubkAeLE7dbpzRW6L/xxii+PN7J
AAg70iJGG+79X1JrgRqCxNhFeUXYrMrCw3KQGs81kGtTsYYVxnPtBeU2rpPnx3cs
0Qh7lgdwB6oaRnKCQof/UJRK4W26qNaOPef24QukK5wTL7m0q7Tv7uAfucMyQyEP
WSOsKJpGYLfaXz1u9Pkl5hBbYjy3uGZg6zqP33yGXvqFDzossZ45ve5j5fTXD0w0
koc5mM1HZZXzk4lWJ3NHzPQrhs1XdI+QmgTZT4N1u6FyYPpCHyTLU61Om4uZtDLl
StN5cAl7E2LQiIAtx83J9tWLsmtUB01GltHXsuXl10+BI1v0Z2vdXJIz+1KXv7na
QbppwIw8GGdkFGXhLQfQpJGXc7roH6jztQqUGKX+YLS7yU7EqbU+8ThAWcSb8fyx
Wnzmq9leS+YemkzD6QaD4qaU3wSnpK2kZv41U80x1NeExeSMdica/G36PtOXtEif
SUD5nYT3KBM9o0S3OsFuMj9jtOJy1+Enbfon3rWqZYbPMmnkC7R/EXJPk8W0Y4kb
zCfoynFPXUX/PD94dliiqKO9QuPI5eB+jz4SiErR6UO38riuhJeL/RbLzRC3xnZA
iYmla27LDeIzZXkOBDIFcmFQGhEb22QIH96jJZJd2gAqz55CauJuvA6hPaPx/suA
okoc6yAAUg9qGyoUGw8WeKNgIOZ6NhRfKNuf+nqgvpSX4mdhZLKBPRlImAF9G3wE
Hro9hZOvAKEgMipGd3aGhoGdMGf5g6ul8lhzsQqwCFGkUhnTuhlS10yDKT/tleya
Am2XID+YEsidHsS/gu6hJLaChGrLTTLRyRBnDwFM/vfpWAimVtyh2gj9mnEvIoja
PlKBLAnUxrLAV1RTyEDQjHd1LY5dJkDIcLFk0SJHrZ1ISoKbQwl3/gry/queIVNf
Gd253bztlDq2GCMt8mAvaO49sp/AFDVZbCJxg63oTK221fyvC5m0PdcO5jUaj7V1
UgVv/ZW68GPZAsjfguqE1VDuVhbMiRAvJQNwpTXBc3zlOXD6IfDMyxpOtHAs/N6Z
FWKSJ6KFaGkobadXrtHtWuXaRtXQ2Cxqq+ac/qOoU//Iha9c2TehF/M70/mwwia3
gwIiiT1b90NcV8eeH524sjslBktGlRDDcTvo008aeMPHzFp+f/DMjw3WbImdyr3p
FPFoIZueKW91z9C2Gm59Hs6ZALlUG/noyCAYvmpj6Ib5HU3C2o23erJBiLtFftXA
gLM9eJpIWPmDQX58mjQxFouD1hLF08tlDb/fZg3lJEBsidknTa0FY08PyDot7tIv
42fQYT1TLjTs8MOxwBvL0qfASYhEn19meR/vBNobXNhJKpyz3JLIiXQsSVlorK/K
4/iMgGz02U411v/qlCK3KIDFAyN4mhRCr6ghIv6d7kwUu+G0BUEDNVxO3MUZX4pr
qSozmY+yukpNyL45iy5I8pr7Q29rQLZBMzOMe59kssdHrm80O2fLVOZbfDpygeLd
2ps/FFsV7zwXrGx5pUicKhz3OXqM/DmHXjCqaO7FETxXTKoGue5tQkCHP3e0T36s
yQ0gh4ZNjFjB7Rh2JAi9LBxjFUBcGyLl1v5TWUh3FRrlV6Jct7XfU1BzLfKP1B+C
cS4iVAbhP+tLCaoBlv+DTRArKrE7l4C4hui7dgXJvCFwizUnvTSLQH3fvYg5Oa4v
9DoJjEciTKNNY2P2b9LTHfZEzqEse6xZR5DRo2hN2vrD64Im89Xs6oOWut7zCqA7
NdAOtHhwRXKCHPcu45M8tao9mQYDvoW3cFOm0wcfh765RYdLkbD7dQQTKNGGyXCt
VQPZWNtypajxi7GVhf2nWQdZgKBQRkHlF3GD6koA+Ca30pxBmdL47Ui6kcxuDa5x
CnOL5SaECSUpbrjh2X3vc1w4p40IsdUyQi+RaV8rAIYnP/0TV2V/0m5OCATXhHhA
JxkTO8GaFYjKsJ1TOG/uBKCNX0bq5i0KTOTlp+NTYTTjVFOw1sc3sEd1TUazACAq
JiyOqu1nVG/0hPERx5cOjocK9glIcXiNtbUjg3u85WkDv4Iohu/6fTKI9Wvsy4TG
hvo+kpuvQFvjNqwkryl3imRWKbrcWyk7GOZVitOkUnDH+0lZfFgqhShxEvEgzYqa
DknWqgm6Pzxx2SZCR55eiN2ml1+9dk3jbAu9DaIMC9TR+UZ+0D8goUOcNCge5Aud
nz15yYsKUwoFREWbAs7FNkiBFD9gwNYjpaIhC42YWfSKkfFglAQsGHg6rCchccm4
AiuifDCHy4hnFU0MMgAyD5liHZpYtjYEtPBh4hTwNl1o2IdFLhoqO3pA4SkwEgYR
3KMGslve5Wn7ze6+66UuvUks9jCI0cMbg+IFuw6JKKrfO2o6tpwmDkOHlOUfWiqb
NGoRS70HeZAJ8JRP7yny4eACQ+NZXDSFQPoBmJYB59WtGHx2X1WapXVpOuqnkk1s
fvwZFCmoqQMpuKPVDrS+GoDnYWA/L8+N9N1nWVWoNXdEpc1dwy7uR4a4j0yHbyDR
6qPK8Wy+FDUu+4znyulDxzIHCW32KoUgxgCNlAwF2SDeZXL2JH1h4//tDbX1gQQs
rJj59jJomeA0KdJgw93CwGNrl8XStAJMhN1goBp/SAkoAt/8AxHaeo3gjIXfID2u
91S3YhZ1Lo0ZZIca54ZUpRkANA3j8NJ45QvT20hgHCVC0I1FjHIPrtlmVg/ldIrg
qonQVEwz+LzmPqXBugNNtxujK/LZY5n8l8BI0BsazscpqAJ+inDN48I9NNzPmNfo
H6RkdoGqayO+WWmXFUnv/X1WHz/kWPhZjjYmUB555AX9A4lIkPDtftFXcPbVPCGZ
QHdFR6VEr5zFRkSFNhi0FEKjiziMleat/A5ZXTyWdVGP3eXm4HwHuRwYt9cZ4LUM
m8Rn3Qz1IAlvqVHlB1X+F+6QKbF++1Ns+0lLmz6kU/5ALNn6VbH2afY+cG6vNSBn
g6YeSlc30KeLsCvIonflLb8IcT9voW2TlHQwfzi8lxe9N3npINYuWeiTU5Oxxu/V
BDOylD9JXId5z6SxT29htKZsYgUqQDzbt7SxGeLd/aPDP/ZMwb8F6XtMTqdHDFVA
R0tpgthF7kth/L+PDY9Vlwb/pXyGJOo1CX3haXgy4V4/ENKgy19aA5y1iqWZuuNJ
oJbV9IJJ6PUY2CMsZdu/+c84nv6auwaOmEL+KkebLfwwZOqKXctacMCFPpSC1nLo
G9hIYGuOASWv/G5R5gVtjzMnTY1QRIUir8mGhbiQlpOa2H6GttqIYaipuWGz+MMy
jRtKgxfocfSS2mr4h3wLQR17ZpjGzDmPf5HocRxH/UhcYW35p1pZQ9CWhXCZTvPM
nZh4OhwOXgwxyeGB8NNwQZ+M4434kik7lqPMgYdcFB3T8RRogkuWnUSReEqAUAVJ
CnaGrwP2vUaWWnEfVa2sFICLA0Cd7W+3JUpI+jf09IEu/Gg24V+QExkl6OiyZbk6
rrNLRPOg+HPi1zZ9RGMb2Wiu6cP0+vLSjHw+SYHNY9u+9ozZA+zRau52iJj229x3
EECKHHEZo/4xQNuDtMyDRqysRwlUV3azEKGMS8cBaTT2CgRF8SYZHQEiIDoyuj1B
+F2T/MQQCtUaHwg25Ys2IgiuXJ/Nb7SLc5Glu1oVmX1spQ7FhNjoKz3cDq2GokAU
OKt6g90OPayU6Xa30o8Bkn6kozeuc5E+jWbKF4bUu/owKFDaZBI96Wv6J7IRO9Wj
M+xCw25HMDBMkI3riN/MOtjgB9V/UqwX1lLdfV6XVLFy1K9k5sDaoM/8h0/mzpzr
vvIqmQfKkOSrRvNLb10E9FwB+dgx+Cp3gS/0lprinpBBwTrNcVK06YbGLjbl1RSN
o0EqLQpw0eHaOiX69sS60Bq7XXELQ+Un/rBUV/eMGdqg39Nq0EWIU8ppqCVsFb81
Od5wH0XFCNHuDKVaKYLVm/3dm+jFd4pFKC30dhPG82kkxpluRAhnT1NGMWvngqSN
QHK7s3Ux2Qkom+zNAFXjlRDRB21AOtqLyjMZaPK3QjBi96zr9/QZyLST9Tcf69aC
+9/xrf303sCGx0TlTzKkk0i0GL/PkNNuo5SACvSpzQbL6QtrslCzLTKxBb24ecCn
QywoPptrBbgt4hElMtnScU6aLC/OFuqYqocZtCKP7aaSwvIpID67ZZVDvUIwq0oR
eV0S6VPnGeYoT/VsPiNlVe4/eVSegB8+ujz79UFVFeSbPU2mUqnKI0liFzSjXmaa
f0OcDsX8Zusi8XzQYxEvpCcqSkp9oX2GYRH+2cWbs0cltloHGyPq6hM7iXSWeFWM
nkpsXB6lCje57foP35k7AgEAhOkLtxZNyiy3QUQEi937cHnv78nBdVINSfLMeP9B
sdeMrq63ttoi+nKh72EwV1i9N233s7K3LOf8f4ZCDAPvJz1HMiqGDgaPt5beVpGQ
gclZFPbfpwrsqJsLO8GFnfe83/stICx0e3BXwiO7Z6TFtovQTQOQJdaoLHGfU0Ih
l2EcAOAu7Fz144zNygJE57Db1EsfOiPP2cNNicPV8ObBl/ZqNIIeVMhAz9wdpYez
OCqKWuZI8A0QuDoSrspYa6DhMSZmKo+XOLR/pa17cRj0KnlqmMO0UJBJu31y8W8W
xOgZnP4fYk3+Dk2MH/bNFduoSHvbG8GugoiZqXQcr9ssei8wM+fprFD8/mtN8Ekz
eyrdIFSkaboRBvGrcY7+8lw10+bPJ6ov5ep7muchog0WltjsRQFdt0rVJa1CeGEb
Lyjtg7EaZM8NN4HIG+e8GZaeDLQjgGvHGxIyC6E1IPYMdfftCOQA9Rj0isim5i0c
M+gH78YIUekN6H31bIKtgQAtD9rE5KMwEI5N1yGVlkaovOiBdjcFxIMW4nx2NLXB
rHSRtjJVLaAGxCTldl/FlTG/3Xsn7zt7ehCAVdpWloH/39ciiKgQxgUvpCwOXr0F
o9KaVvILSybZGHzWZZh/a7rOOmZH/VTp4M8mpcDQkl55wXmkDPO6GcBODJNSvSkV
JzqTq3zQYeKmNUnc1VM1Q+ceB5EYZT5vF4ibO76A2dYLrfeLupUA+O6/ysE+HGo4
WnvrTOhD6HmqL9O6Mpj3K/Sxx6Ys5YmgXgP+Jn7jdbKN0FNXtnPmu0xmWhkh6mx4
Nt7pic/J7Yaj/ZTbYk47KoT/J7yaayPctqJnzHEjHVTodrUDSHtagYuNu1WlIrfm
lfC6EDLBBUSZF8V+ODw9DdG9Kvop60r/0HPocifqti07JtoeS2499roUs8kifpDV
Jit4S3DqqE+lwX+5KnIAcVSzZeK2hecz0SXkHAjqinVj8mEpZPMTNqalMMTlt2bo
xkYqWrCbwGz5PwJkvQL5tWTBUZm7D1oiCV3UoRvXKpqrB87r4qUrFJhWW363vN5C
2pZYcvXuW4hTf4qAaPD6Iwmb55VINtuU0eRVV+Z4JMWs8isQwit/rRZIFb+/TTzS
H69DTzL6QflohqaOGr/8f4KHut467Jtfdm+gNRsnPZ1UFh1LOTg6G6v0B6newdwg
wenjX+2HOJAkrJ0sUBGdtYp5hE9XTfXFRseM3AEok/eMl0ShJeQxzaaXPVn9zMSX
agb5hyjoWI8AmkBa+Bri9gj+LsvL69X1oR2RzEb5BoV8mW5sCTgiUiMbo81Rx3mN
oTUPSOf4ERcCLn4cef9s2sFp14NnVEpV9cdmwQmwpB/HxT2cwFzEN+Wr1KhAOObP
HWLQUReZz0CnVsostkttJ7fVGIAdYRS3EkyNuDQJQ3AzaNgp/THj0cwhPMkd4iAS
w6x/4YbDy47R3dhSICg/+AESdAd3A9BBI4xY3YAVZcSMGJ0HkLAFWRLTqA3j9OdF
tv1Wq6ci++Elq5uNL31U4dERnG0/A3kjxB/iDtYofn0aAOk3KmWns1u2B2YjldUh
GvYmYxjBlxa5jWKJyBu99UiCb/YCecn5zwfYEgsiaaNfQME295wrMjcLpmaXe4ae
IcSQmSDX6UjnqiwSdx83zSBlX3q8k7MtyC9PRNQfGFAQdK7soW+SV5FfdXHbB43A
9DmR3iGtwGkh4Vaq0DSzMTfdH5DBmZBlkfE0ShrSZXW8EN9/a8GaGTn1yM1RIir5
kW7pa1ff+UsXE2npZ9QULCJ4c4LZFWp52Zlf+YX/qMQh/iGkrOF0/BnT1PWPnrci
4obQNmHXZvreEpS5ge+7HUSsP2RMQU51ZY0Yz/P81dnO4AZqt9Kj326GKcYJMKQT
QHR9knyaJABhPnx8yq7Qx+gKGag7jeAGmmCNes1q9+hprjCgp2bZoiM2Qh2i8S7O
0JjrjrRl4YFe27VbYI2yneOojVHZI5FO0EAdeJDIUvAci/nlsrio48MZOcwgeQke
DSxupIgAWs2sc9qieGql4nTIBE3shZxetCT1asHZxAKRLG8BNjOpLv0z7n+3T0zq
/Z3unMYiaaABAp+H4FPWcwnhoT3YmP2gYVAPeYhdF9eOiTXL+EA3gTKJvsXpvcgQ
BHl6KyKPqsZnVs00/jWNKGaEW6WciZ67GLuFsxDY/fls8HSoHmKtC2TbzvUW/A5E
7Fnyrc0kgBLDqSrSn+TV8E64gn1ijg+y7zDm4wKvtv8ft+cjMgsZyZkTjR1dZqf8
HYl1jGHzWRx1o7f0xx8CnLiUX8rSIDAfmxSgWc/Nxa2vtdFydDTdl8K6KQijT8g7
JBZPtnJdshuaBkQZPvtD0aPzimVDwv9FY13UoaV2fJ++CpPtwFZyzz5IFKgtIcKy
y2AUCJ2230RipCGSMSkmUC6Zj8B6NXReQ9xxvj5hCJTkZj3JpShEludGtdFEB6Vq
CAr5MDxuIQvM5F5JHMPbSfRvOE9CMjWP7PqPi3MUlQkiBWw49zeUX2AWu6yDi5IQ
MgL9GEMWCZG04f9CwrKBdMlIdJ67r8Ju9OOyZVbY6VG6twE1F3djPmzBvEzppP4f
ReX1id1dNVHCsRcfN2Hy8T+wWNTwp13IP1tJWZyQ8/wVCQ+gmGw315ywtULIr2O2
b48XbkRYvbcfZQ2S5EY+Ki0hizv+vYUHqBOV5jBWGdnXi1nAQT8p0SugVCg31VLd
+FZOjl/y1ur7yUFgbij6p6a8bb+XcuX4HE6MQ5jN+TxRCPV4jTdsj+lE6mZmxzEa
PujeG0Ulbo2e/bRwA6hrsn0HclH8k9iWknWwdE7lXq7FBvto0jy7T0horhn1M30I
uFxEv+bnmfrTiG8Dkfdz+rQGcqC8saCQF8e0ZLy+7U4DSHk0A1vzGWjQ95xnrDuz
cJUZLRPyAHFJPJVsZi5VcHiLJw3eQ9z0I/smD7tr8ZNIG1eeiUW8SIaVxXnJVo6g
sP1tPwlF5RF5Y4uQRHjoyfhLzy7BimYgDuhuly2HzPQoBtlCsT9e8YA5JgqFTe7p
4B5EM2ppJDAdMQ8sviSm8xUPPEl3Wr4jWDdYZ1KT99i80v9Y20tEphw2H2aONtns
Mw9g3GgMihetXpxBdnelJuAIh1GBzs81cwaGtrzSKTopzHbGNimp7oTZQ4yVD9Ei
ndAtPVK2LSDON2vttGlqeggjtH6826ukyvfQu0GxmhX5JNdFx1NdP4WlGvXQf1Y/
Hp5zjrZLnnZvXzxPojcend2gW8PQFhNYhFJ6X4fqMEmMkAK6DrPLxa0fO1apvu0H
qXn3u++Omoaoh8r4FIT3T+CEcGguuREPYt0fOQvxBHeMXBuf9Sc8HK6JWe2a4VKe
1p1k+/WakL0n6+P6vVZhzX+3l+ZmRmTbxfbbqiv5j5HCJlDYzcK6jcboXVx/lr9/
gMJ/zn5VK0qJ0npWEdOwq7Q6/b0BX6AONx/6pys+MGoX6EMpmMQkpc1croL8Zl9M
ivG5pDz7TPGInryx1juMZhCLxfL9avbuAja3hS2qkE160AaeVhsBQi/x7/lFO/do
okSbhjF6sIRdne1pqjr0aAKMkjwPOVHwJurwXsk6IClZIqRliXOJ2Y4WCRtIstW1
aQAGmo5YXduqR+0AGgiTeeHogtVfgs3QOCtMunfk2/OoU1NmTP11xaFGHmhzUp2N
u8T9JKOUIgC7KozMAKg3Ofr0rBQO70zbjJWPIIFPRKr6DFsMj4eJo5+ZKaVsJW7f
Jh/8QtSI5b/NeYStASPAtJWF8OXRvakuxUmCXaU6mLVZLXwh3lEZoKXOwyPGv1sT
qeggbFjRSh3LpH2JXnFy+62ROgTbzWaoJDz3rgNZ7k6bjF8cB4/ebiMqx6XKYtOU
+QDyoaPd+Ja5lyfZFZnMUMgF66X//mNovkinpA8FTwXTsx1ys5xZMccfCQ8UClvI
z5C4E7g7G+L2GQAGO6OBThcjOpgGcehWL7jH+9kctOIeNAOC8sBRpmgFKYQPagLk
Dl819KQS7OLNEqDA1tyD7DXVUNjVZOnyStGz4f1j6rqp/+ZQQqUzcQ9f27g6eV8x
OZqeXdd5EBsKQTC6s0Ee8QIz4OTlz58rzOCd1R9JAtisoW4ZNylwvpC8+BquMnKp
m1qWrrQQg3vGprA5pj//9VBSbGgAWTd+Nm4QugTg1kjMfOmGSZ7eTwLgm91qZoKp
V4eSniDKir3//N7hENbyq2lvt3Z9Ofe07Llkzh/QzoRiW7MddSarcveJ/tEA//nS
c1PL9/sdFnDYA/kjepGUPShDSElFjbCV5Jolnt8fAG/ULepM99yRAthr8Yy916JC
psON60hwaqOmNvc7EeY90yw43rsSRQPzp0D2TBrX81o299Bk+8mjTmxCx0YZg0jE
KnuJsJM6xhhYwWOeSgBr46gMXXMdDdpwAQtaIDWk3wBfbcLbCedx6+hnJB+p3ws+
lwd1Iwa6QAqQPoJA2myBFmdKsXRri2tlx9/YqYIlwhgHTfhXID4h6JQJROlAIEj1
TJ0Q7iPj5nz/nBP54dFWTD1kuYtprRXQMZzJeWCmHGaMnv5/fJNET+Oa1GTm58jl
I1H5jxMiMm0JN1oXTx/Bplz9LizE0SxpDeseSA2C6uvO4jTABcaV45p1/uAKNrZd
cvXNmD8EVf25yUlWzy6NiODbPEknzXXNu9U0pyb/BOiEnkrqtApdvihivI87TQ3x
vg76C7IlLIJ9ReD5Gi7fXeBP2z8ciKoy+WUcptfzGktn2PqKZlpq4v0hEywYZ1Jp
167sm3x5yonfcoh2BojGaU72KSMcWiE4LvXfXo7SzMFtzFv0ZqPtY6FPA9sJ9dJj
/RU6YNXQ0xvi8HMpkppFFEmA7Uh9/4ARzptXSTFPP4s8c22JMRsduBLL8z/5+Uo2
+8f0uYU+vXs6vIC5L+ncRBpc8woGUa2e4JXcMwOo1n8/tn5x+Khj2H07QK5x8nxq
XvSHaTpF0/hUzB5rlsCbBfNBITDvpwghZK/peO1CtJv7eQ2zUygz7/7HfrWxojBa
Y21CfqmkNFJLscu7S/kytPvnUNrAEze6wHRl0fgn6CcADED1XXUBN5PTu2OOjBZv
4aoXGdQDHKNZvR1N0T6qLy6KbPLzBBu1nuMqurOR0pD1xcmdervMIW5AJbzKEjJ9
W6kNvZC71J7ALaA16WKlcc0Crc4KTLERM85RaBLSr5Xy48OrWYSdOXFTrLFwUH4x
FOTMvSsuSsgBHqxLIQ3ccNG7B8gaaeYAJm4X1giFUjM9g1Cj1nQ3HVMuBbtPia3q
G0AGHL/D3tkAhLIl/SukKLSJ37zCFCB8Gbp7LIUAXf1Kef6558D1f20RUc1Mk+Zw
TFSAQzTcJMB6XHsQILKkVP6NkdS++NkdCvAEkFddNg7PQac0LOLcrIR03Mrf1gWt
D0S8jA/qiALr2GoevwBgxEQxChonelJ+smbl+ayJ8eMWvNjAj99JlJRkaNCTpf+3
JA3Rnt7NxAMRj3gqviIDgMLrgE3pVdrLGoOPxFeYukuPDy+mHDqTKbojqEjCcLmS
0ikR3Qj4/kDgg8M8DcVhGEdCNlTOse2VMgMLQEaM/74K5UEUHlUdRHRrAZe1S8IC
p3uU9MNSYSMo+4LZpLsyJ6UPUZSFWHEke9i/SR6FADMeSLsIDAKvg/p3zFqyfsGx
/IrMN03GIG69B7dQYJI3ekHN8V7gvka2FHJJiVMlxs+VzLKnOh8CDR0tvQYD7HaX
2PXFeAbNvu1QFDln4NCY5296OTcbK6XR6RQcxw+xmU5D6S+frRLJXsIoKzISUbX6
usEY2H7H6V8BiJMyAPXmVNeZhNO6897GvxENYkNhvI7VUsc7pE45znxbe3k4Lppj
j3Uf6BklaAQNkKyloDl2hZNX2nDGRe5vsOqCc0Hy9HgNhu0MjCxkeFsS71YmFJMN
A6/vPeQ9kJZdDKImUdHJI5q0KIdGWCED11MG/lVaYa3xaz9puPRqqYbpJ0BZlREs
Q5hxVbkC6mtesymhjCxGjLT7I3ej8sLquzSIhCXtUAvcn3tXlH/lDM7lo/g92P+F
wKLA3ufishHvFmW88jeMsnLT7tThCtK4ovK91ANx05ptz8lBd3fC3A0jFOSMWJ8v
OtQuGjUKh1xbQnoeV1m4F/eLUNjjBbjPiX8U0Arl0rJbko3mCsyShhCkUKcjoOhr
ZbFrcoRq3/RERo/QM+NtfXbtXj1oGeQRpBXfxPac+fmR6sSGuZKMAIey9UzWGoJq
Y6ECUH+ZujbCsB9TNfsOnXJJdt9vnXQX3HIAqwgfuwBTEww1bdhy9IvPiPmNCDs3
an8GGiEbNz2MBcrVgAgS6Kqkwo/4sFBBh6VyNhUnKRFz3iDjZDBo9Ay626sd1l4i
7b2BMfvuFWUC1U21ZbbxBnk+PbkYBFpeUSrzm2bgkgAIBPfC9MjcQi8JvS54UXaS
kf5eBLHwqXcS67SPTZvNYVwnZw2Hpe6kDtq+lyrEdoBSxckJbU1w/nkMtqqS0Plz
rslq+koO1/zRlIgnX88PV5bVKHNQHdELUWdH4bD36V6Om/sFFZALrM7Yf/SxuojB
VRZF0Cmi+dU5fwGcjVPC8A1cjODgJjmYI3Jh03ujWWUMJz7pxLBRfoSDrtUer4T6
1QkoU5isn5a3ZAs4RjntcI2oR2w83SFINVeYW7Kq+3AMGgeHXepJ6HxKmuG8sjWS
WQ9In6eKMWZiSYdRvTJ7es3jRO1GQUs6Nt7wqeBta1ukPlKwMHZAhhGhbl76azTJ
WlgM23p0Hz/7H99dUz2XOeINeoIVK9PGbRZKvo2HFQqQ3toj7qOVXRO/pt6KnoYV
icXq2s05LW2ga6pX/shl03uSRyHzEfEER9I1r5G9hJIIe8qo2OmoDwEmMSzFwncv
93ktKuln4mZNrml+xUnXsw1LnsFu9BR8znH9vz61heI7qs8TFuWFawNin0/t9Xqp
ZH+koB6xkY6mK9dH4pwAQvnGDKKu7VX14s1dtR97Wug1YTpCqzPVPIq72tJyC/ld
GFJy5rLwp06i90FxfFN08qhNn9THJrwwSGkoOpR3B+haMZf91IneTGQcEsDZj10e
RMxsCX3BCwz118SbzFrNbW8Cwm0WsYuciI5SXmuFglHiET/D5H7bD9WBpCr9IWii
FDyCsxClCfd2UzOb1peNnd8YmuGZsESUywTRH6L7t4eyL/YmD+X/M7HWWDc6XhYk
F3nTLArKTLENQ+MCg1q98XhPH/RnUahHAuApvgRuh+pJ8OnuJuOtxFYWfIQ4TrUw
B5Cy07QeOlkBFiK2ZwqD5fPC+YGqZDo6DytqAkOTDP/E052ejBnU8PSmIoO7pJvD
K3NObgJE9Yw/ym56sz6bVecl58/S3QXVbsQyFL70ZwlU15b4/8xL2V1w9rm9szdm
WpMkctCx2OhTQHRLmod4SfAJUO5HUUtxKUm6mWEdYCwK74KDpOSsQvdAPJwKhboo
jStnOCTuzH4BuLKvJUH7XTyUhZ9J/tKh0PxbPehGnZXcQI08TQj4P2WrRqxEChbl
GG+ndJ/ZEJueI9a9Nc6At94XXzpyQ4g3+KySmu+7CRcsMZX+/ymWZesrCZ59jPCK
e1Tq3ljwwLw5FwRxXIhAss5xkqtgGA6A4OXXkckgVyMDC0ECOTTbcFOrvYZLbbkA
wMNC3iQJfeKO0qRb78y+VvJvrPKLhnD98+1WskiDkoER3mVXXesu9QOKqK8xbVOh
PdZCgvcfGkMkfePcIqiv4Ji5GMLPVz8EdML7xrN9GZxq054GdvPG+6gW9rNTUCWl
hazPBjca9yurSu4pg45pPsMDEafGlFNymHIuMw2QruC80gfUCY+7D61OAgVQXgrf
hptikJ/JcrppgU9f6pi+pPcsotdSVjmAhsXB2WDgwCHduf2p9r+3eHwgeguFvxut
YLvZnDH/mowPKYb53BEyj3XW3/8Up0i6CMZEk9bYXEMeYzh0ZjQDE+IH+l8KIAl8
1Mthej6G96xdZHls1KQeAMg5S1jhMDQ+MqzKvrVpchE3TsrplOpJTF3JL1dZM1xH
ywLkcrSfJ0GA7UjF2eV7b0eFMjQGGduHB0xsQNfLsGu8SBKHcOjmeghWm/+F3jJ9
1lAlzmfGaqtZNvpoF9mvhVWu6ztoMxVZI+to/yTMGK3PjlNV0tPHzAtqdh+sUr6r
qt2Ka/XGINhaM5tJlKeyDokMr9VamCxAwtrbC4iAxs8Ql8jkS8GNRL7oDo5xsYuW
3AHtkqvCGn+lRH+rXfGpSrj4PMqMftRcuLlKihYzLQlsT3XHHKkxcGVbs4rdvrat
sWpX7tT6XFl3rjOz5IYrkkY8Qr7GB6xV/3g5SlrtmYe2tLJasivTT3annUUPeuJF
6KzGGIC9kPVzbRsT6bNoa3kl1T2JttIzqJ3EPJQMXHmRMwhK62PcReOfW0IILdkN
QlFGs+8B7dg6j+N+51nvvP3hlQLbgiiyyE6VC24TWnqAD2fGMEIikI/uUqLx4MQL
JuVNZOsRdb0tH8YiiJn2KsbWoagfhOewNSqDLuv8/OwcrcRjZQz3skdMRVVgOMKb
z6sCTqLmM13qK+arQ6eIHsbc/vu8/EITZXsotrOU3tyREXeK1SP+9uof9137qZvT
xKuHphMD7TlVqykkUpIN3aLt9zBzW0xfEY8OqnjFq17QbLFe6xTeORXWKZX6TJXV
uAn5YQ1ZryIJc9mDXmvCyAN9Wei30XOMKOVyRwQvsj10oEEtkCUXYmGOJy0VvNvT
E3zHMZVZFkVA+gegZC/iKqyXRKibQNIQqBfj+uheVUkX0Paa2BzuvDHD5ACwmo3n
63A24tPHx+64YU0zFfaiyojd2Skq7iFdOOzCUPXmxtxhHT7b6VY/02BsHwruxxYo
VscM5s7ipNpaxKNQbXAXQ6FP1bAmNFi0VGrIh4zeg4yV42pXG5Dk439j9wpAuKtG
NSfIeZ+vGZO5z2Chx/f5aUz5hFtFRtyyyS/aTcevqsMDw0hoXq0YxGw49oaw19Gf
rZR7fC8LDMC/2bSXyoxG+KoiilswtRZtouTtcccL/Hb6kvKp9rfYJhXuokY30fso
xVRIZ4lTKS3ESvMlibBN2toH+dPkbB2B0Ye9UnNiY3KsOo/6/oiaI2HGtkajFMmr
mlXvN/4l749rYoY9jl6Un2LhP2xMU42+TRo2Xg6/6yZXsHZOBwxgKethCp05XJ4a
hNkWsz96Ge9fpofDnkmi8V8/c0v5g4YbGOOvOAUW8ayai3EGIPjwr3o9p2Fvc7vC
OWw/XPYbLiyn+GJXupCM7XdnLtT7SbQimGt6LhvGnAKjmeH0rk1lHMW6vFzZAcny
kKvm7mOMbXgdIZpWL8uHoZoCgBu0uqgI9QEB0OOlMVoXd5uAk81gu0gacwk/uHSQ
7iF3G62Qoisga5r9vKMT3eu5KLR3jsxamW9AwWlHW53hueOHasWYxhXxlVpydtlg
ZqyEb0twkNHWdQGdtz8NNtucJwasOypvTf1GAStRX855U79QFqn9zDothSDlArmr
pejZ9JxFNK/RmHS4e+rMayn/+yw03VMPlknJveEcMkTpmUpND3M+VQ+bHjTvEOCc
v/lHr3PevdTxJ7QlkRU4ksvoLvavR0d32xPV+lA4L+3PuBeJrR9SK6QhgyQ0NrzP
zMUh5zkEljpyed9d81yM8NKm4TvCkRqgCrAWYIWYFHlahOnM5TJFxp+GKw8J5Kup
hwmXlYDly/WXVKWop2i90qN+Mu1hBrDln7AHRr4OUDgm6ehNikssk6S1EMkNMEhd
qmhoVmepwMH+wRZU6TkGkfPsbiXQ8EJN49DJfeN4bHeXG/MnTeOKQJpbbJ8V2UI6
nk6TNWqE96fLLhJNln+P5F48Fx8RFAlrNBpI+f+0yuAusekl5hDPVF0REgsY6uAj
2U8VuyPOXYi0TZOtcHAtsqbBxRH/+ZftpQHInM3JrIbfAChsabLlvtXc+pa2FN9R
ByP9kULadcX6oEjp3CCWJhI0gepgIWJPlpcRkeue2fmP072Rs5ig6wbNZpMZwD1t
gC53i5REHNCH3wVvne4EaYP35LdmvtpN5jT6pt8mWUqokcG404eN+EoosXeWj1Pf
HA89s88t1ux6KU53RUaDEK+d81kQCve03Rf0j77P8iI5U8OOAfx9RIhr7HXgVWRc
aO51M7RkIdOFhg6gMB8js819CQEWtA16fQ+d4G7F4bd2c7PiN9a0sbrAT3ovUcJh
cKAtXgt1eJmMUOfvrj/N4L5hqEqai78QNlyT73FBpT+1qkQBAkMlg5OzJR+YQNMH
CcD/egZf/HvQtYngxK8pLZaMpNC6uWIiPGHkJCJhZJgejCOsKFt2NPF/Q8zNuaiJ
NmZ/HfvWga4rbjPkL0jFSdsomI5mLGJipWZpg9eeOnz8xNwesKHLqJXtgYkkEKax
O4ECPGGnQLF2OBtqlNRgm3zBiL6fJs3XuuaIQ6ZHGEp6ycsgTYQFQTsjsU4nS4+Y
cx2K/60mb/gRx4/JJSM5xnrGnwT8lWVgK+1ScN3l+5BCXEQmMQ4rIR6SHfbXyPzf
8Nh8fnOQMO6ABqZHENAuWNN9aDs6uIB4isXGCGUQn3lx5O0fkdsHc9/71TqEi23H
AZiWLxFs4K3uOq+GxMYgyXHKAONm14xxKtE5H0RjCDQmawV5txNNVIiJPgz7uJwb
T7uVF5A1KGWJK6N7tpChuYpelEmvCNr2UV78s/8vItaGGSsgP8aSXlmyFup+RvBm
nBijHgn5EUTXkexNlKV0iu3dXpJ5oxbUQ8AY6n25tAK3a4ykcRB0PAJKf/YmhLqy
R8ZxPHSIrxnobCOt3XKvcIKQJ/8jn3gPUoepS5mUyXtQPH8q8WjwDHzjq2lQE/vJ
eNUzj0R/ciDLH2x68Pqt6Zo+6X4VGKM5w9Za2MwZCYsHfkBaxj/NyNI9aIx0TYx8
p/LVg0QL2OCUMFPwzlrfT2J4dLScUmon3/2tMMhyEv0elCEThUzRRdUgpY9FYG4r
+bnCA7G+22vGfa8szzPz3uNVu+kiDZqAyV/5wbHOX2mBmjMEV6t4hC9Fi0Qrzt9c
SJLKLMsoCgGF+INmyodma9+Yb/MmM6785J/O4NyiCqa+8uKiMPrM0eAVwPY3YO/0
9i+g07ghUzjKMl2bdb88Vl3m92YIKWsWrvEctnhHs9t2ogP4mDK9z7f07J3REJDl
WJ2Ov6UUrc+L7zUNhEsk6csuGRy6okjrN1W7dQeT+73hyMCsjbWmNxFu1Qtw2VVt
JSgJHvRe7zjJgjUDbAU3OObzChBCAqfRv5Krlvpcg+nuuSENskfFBEBrywRN/pD+
x0vlZzL5++PzqREdkwNVL0vmOJEi5pGkA2+cKK76JCUxBvc6WFIoWhnfU2ccZFb+
1iaTh96SyTU1xL9W803OTmDEjXAggYq+58mqdEBiONaNm+BneIRpWpplPVP6nAuq
q9VVUNzLgxHOBwKhtC8Z1v2euT0oRHblzCNI7Q2FNzwxO9QNG3fCofimsQiWOhx1
VgR7zZ3DG5IJEwtsk3+w3Ue/CQZIfcDLNkBbrDIumyWFTLQoaKlgPRGIn/gfoWnY
fjRq/HkLPJtq6g7oI2BRfzis0jSkw13VjSMcxUf25+hXxdRfPBoDweaAewr5EnLQ
/wZi7nNkTVOK3P+45aFEqsQomdHJM6E5p1j1A57exm0ODL2g7/6MyINMxRp4CTvp
QZI09rhP+QQ48dQTSU2XaMP5XnQ82hvJWSzUiYtAP1YfFA1BtW4XhRwmbR7qvvUJ
TjI+/R+7kheqb2bXTp5xVjdsiJoX8lTXnnczntmb9urOeQpgC4yHXtv14t0ozjm1
6CEhR2ZMDuzgXKeSgDa10v+eOvLGQYMz9jieIIehpRCjvRV0v/+GlYVBSfKQzClt
NQIY3WLDmtWfeH1l1cn+OzbUxIN9a5R3OggDEZup06kN7j/BqmazqINXQ7trhLa9
QtlHHdjY15hiGzyi8qNXASOB3CZ6KOK3YmdlEV5nSuRTMELVxQh8YNHpotsmuZvf
MUf/VM5VTjPT1Rux82LkzN8aba5xz3gEdLczhBv4zOXME1eNBzdJ6/WyvkOEs7Iu
uzehkzcues20Q7da7r2l7HyVpGL9ROwz2i8Gj2xcsKjnh9HvFEKvRSeKQ1cCmyYT
f31yjrRfPPQKdqtykc5bvpetSHxuPvMagdM2T78+BDa3JVBvz7va8G/6/rKCjffg
KYwBkATgqusPhFfqWnjGu1AleebMEQTbLM+RP1DPh6SxOzFpaeBjtQ/aVpglMwQI
008grGS/lU4fbdf5LdKe51yN+JyT/p8QCP43QPdPgTfjSZ9YIGJ+kXptsNpwmoWU
WZ95QixsnNsODGNndAjIa05akbwVg5KZphHBvEV1zGGAa9Qj/oJHhhdD/0InHZgk
V/RHJEBs+CsS92lGjau63Kk2n2yh1QoN4cD7KiTBTCFNh2E3q2gH3l8ce6tFTKgI
3oyzY9v3/2LERKnwtmf2YJjgbVreQvBYP1lOZtDU/vupxmITIodmZwXovrciM9VF
iUHxmkOOKUXAYydIAFDDE+w9h5AvVYlrW9P/67QWXWg1kejKMobvFwFkaRCz4EUM
8e6uhQDHSgchxGjnj3ft4QMzunze4LmhsiQn1nBi9EGV6dIMLHUdf7AOCeSxQm/1
yqBgsFYWE65/3dw/mDu3m79gaqrOxuOuWFtxeTEyMtc0wmPYLLowjeie+hEBEGfm
CrCZzox2N6Vl0/d/oW8u5XIIh73i5kZXUEsdkmYwtNQ+Dw24sCZmPKNY+BFeIdSg
flWnr3CPvFrUdh4IiMuTMIdv+MhsufZvIj65aDU1u0B5L+GIDwsYbM4te4zBfnc1
jmv3DY48I7KXbLlhj2CzXJ62hXdzOUOkdJlfVnN0Aie7YSBuhQyMuT4H1gjlE2pf
9vdWel0j+ADbYHpgCFCiZl0iRdwcXGeszsTEVl+4JkYMVes7WEQVjIH8IspwmCnY
9wmcPj9OUZibcSEMqmLEzLNY7A+AlzYEWSfWGTa0vJTrtK2EZb2DN4mkInijdBCR
W2+bA03xXcPnKMHI3djVWrHwxCTtC7D2yWcwrWESQZXGpB5/D53v1DEqSu/bEufy
JJaFplgV8sc6MXMXPBUngzexMoTm4YdtXDaOsmvJTLQSg2TZCllOOQ+7KdzK6aMl
/pNPys+4Yb4ZuOjLE9Tc/59F4v9y+GXj+sY2S2iBtTTyT4tESDyZXOxxl4UeORwO
IowERudMQemhNGS0iWJUiGDjEXH63FljvQLUJDtW1u2C4DVD2BDIptxApZdRlNrJ
WBIpCrzAYH4EvZOudsSNCJrf9DP7Jrg6eBSfW+sSGlevfcTR73+v1mY84O+M+6Dk
i2S57zxF/kINOvR9JWXt1p9owBS7VSxobsVtCqpgjHYqRt8Z75FXFN4zJjCP9Lw9
utYMmmElYZGQr3QqDUwlTvv0qQqL/O/YETTuyaVr21G0NnGgiTmOhRUlAhHO3Iv9
yUkQ0mDQhL3joBC2TfWpz2FuxgoRDHde39rOvO0BZ/yWSBZtemjp6ToUWwVZdGeQ
Jz+F95ZaakJdnAcfhHk7i1CrilmPTQnAlaYgxGoVRjib/WmSrvjS2mwHMyeeR0ae
WzkhnpeTgDKMkJUBYxlVYuKcn/J6sAKsJSKzfHr5mhqCDZ4C4WzI28WKDS6y7R3Y
rqDZImWXH2nJkbHLuvSl/hCk+05ag+/KKUjd4C86/3a05KPfLa5IgKJc5eACSM3n
j/8yeYTEfm1OxssUAriPClxAlbZ+Fn0pC2ERgzCitl2tGFghszUrkVyE6VUaphXH
LhNfBi/PcsSFkSu9xY4M4xh13G7B68Fyvk+WKEz1XWCud0er2w3ZMEZj37qOCyY1
qXoV6xU2fYcVvGD/X9rfGJTimMawp3+Fr9s3W4lNhVnwOsPyGugnghggBDFHdBHU
YeMHUeuNjx1x2WkMWm66R8gqfxZ1uutlXUos7C24a3DoZmMckQVIrMxtM/FhzYJs
zPZu3fCdHOrA8BtqIHJtr+DhetCmPnrqvWo9u66fNbl8GIMxbDPp3f6ymFUb6qSM
gBip3dzhHNmmDPe6t9i2kd/qL0/D8aedOvhIz8KwIOOZQBAa+zisY3UToGGQK2M9
QCVOCbTwgeMO5tkuKbgbjbwnIIE1ph4kTiyNcc1bxrr16g9gbbYbadh6XM7HHh/T
/UonStsKSCyJGbz2Npy7pzRREkH6HUSscl16f/H43yCwS+nk5OSbE95robqCinP8
4izGTeogAZ5ncjoz/3k8bA9YSK5rDNXTRtk0Vpc4U3zn/0Qwvlh9qBCaKfw7x8Xp
3ap34ErQwDSJ64ke7k2liE0AstKDWnOBDRVAWT41qA4apbI6S429VaiaWvxL+zWa
37b3apnahqvjwtaXF/Yzmz8cNR5TbNxTXBTp9nGMnH4ANPcESLgPa6KIfimtJ31Z
KqLSLTDn9QJuGFRmFkxmX6Ieg1H6iXZa53oeTlPLZ5DjGVPFZXD3o7dtkVDrx8Dk
YtiB0YB0mKV94pYQFmU+tAVbU72FMV3yVYiL/ER1xcs+/+3pewNTiKuEjwi1QfpZ
K3J3tH8VMvmiS0JzrduVQx3hmGXm9rVRMv39S+yILRECD2dr3PC5iYckXZIgm5rR
rThwbnLoX/2ylQpcP+yuNANAeUPEE64El3bOU3RpatbdWpgSPelhNGN5jdSezZUR
EjFABKBWbfYgvPzYUF/3XLbbMc32oofBhiI0+CxhRvjI7/b7cp6khAo63OkhUyAE
9C+SvPEC5g2TlVpyEEaQR3m98bK7ILvMfaiLM+DoJp1Trj6TytUAqd8EzOICG+en
h4xj8VnxX3az0iQL/RhP9aLP4g/jYezX5SOyoukaTw5hP5I7zkoEoaPjZv3/cQf5
USWvQ45QilpjNQiBus7DtEtl90SSgVlxT9qb7sZx8BMaI1sOxUN/2hPw6rMoLMoW
nY82gOzIXH7o2f547k4EWlpWtU0PN+/XJWqT255kqYBt/JAyeGax9X34rnLF3+k6
ShrzriN1+I9KYrYatgSsMlEHgyGPPZ6N3YfQmx/Xya8uV0zVNCyjHySsBfllJsGx
m0wHq9X7F0TAWMh4e2qGSDj2LSgCP9uAEwwELwFBlbyzP+oRWI5KYS8SUkw0jfVE
98Q9BJWn/nhhcuNPDztqOy7DbxDvOw9SRcp+uKig69z/EtFjB0ZRanTa6cmVJjOQ
cUzX9lzaNYrcoZ1bvg41F5sF7LfxvCzCgE8EFl2wF3JUS99pY6vuL/1pQSBiaktE
UtV8UnetOznuhoXrdsO2mLebngRTGJiAXQCS0w0WSCuc3SZX13vr9Gy+s0+YUQkX
ZrL19dU41dXazgFwNENZSPAQEcMIICz9+PFxqHVUt3o+mQBq+4A0VePNnruG9kY9
lwrzRQTr6nBi3LxHLICB3Qi09i83gw68BEgYpn0PLkPEThcG11o4tW9ZriC3dDr1
XPLBdAyYQGvs9xVbto+L+3O7peBAL54nYGQOIeNX642eMD3pKoD/WTXv5/PJDers
WrARYOJRTVEOWdlF1Lj+yw+AZBYbiTQ0uYaMfMNrEmOmBQ9IpOT6VXNQXdCxG3lW
wmHTwTVpK4dEjS99lLveQVhYGj7ETxeHWRkGDWqyQ9JVkOlLuGiFtKDsoprfjWp0
HlnzyEaq4ncpAWj5wyjPO3dLZjLp6HQao94CsftHJgEDuIaqVKqYreJB1yxmb61l
7XCzpsIv+eBLIEbDhbwWcMllypOnzs+fpavQenuoaQgoQC29be0LhZ0vvMmGhwM8
ZGKIVyXcEhOOwm0/4axkHFisrxWxpd+VRZu4cmAgKausv75aKXSx9Ieo8DQ5ZHvw
6XWYVPFGrORgkii62aL3kAIq9YJl793do2F1Pkdq0pWzfIUb7Pr7efukHgh61/4P
ChuzP/MTZ5L59lIRnqPyCgWMnzQLPi4WqmkI7FehGLXJQNaTz/PX0w8lx2zwo0mk
OQe27oE0zqr8GJTaA1ex5fv0go0dJNRd8J3/AGzpA2ldrBVs3k5eT6sde8luSOqc
BNkkcmzusV1yqO6c2fpV9veAO0V8c0Al2a2AnEPjdhxHrRAqmqBVMuKrJ6uVbGYj
JE6Gtf/PMaxDvkrK69OHRmvrMBSu6nRNMOZCuhK9FCGUhDp5Li/6yTWBQNRFvDKZ
ztCI4Gr2oOrPY6WixKi6JCQ/aVsKKpKUBpq5ebi14Lger5v1iYlfTNTL7+OjV8Rt
96RbrBtCce6gbAzkwU28gSGHcQMt1M1ziqs4LGk53LSpL92LHq9fRnUZJbCrKLJk
w4aLrO+8YoUOJGdxgeRHCgMiK4k3ch04VIW5vPeG4sZRn2xmgxxeqvuS4U03z7mC
fZxgQYAUPfDX5Vjw9CkfTVJQtgkSqUj9Hn4//UHMR7QuTRXCu43gRCzDzMEXCHPE
8BmxRpTfGJ4HxxwFdZ+WHdz4+kwH/4mWy0nBZh5UtRmTcnPStDYgCbo3b5szM3mk
OOsyujwGpp4/H3pcL1lyzMK7JAanhnuERL44e1EHQjgjqykaJnTo4ZB5nftv+ULe
a+mQdoySYM2d2GoTozo2Erc8y46dN31T/dFPqZfVHLC9D3QlIgqEcI3V8IajSHaX
K/Fw/XQFDBCvMJTlfH/Z2aqv4eMFd12tpvM5vEXmwVwOMRDrc/HPMDXvLDkZGcEL
qjmIn4M6pynIlO2OiahLjq9A6SVWIDj4TJwohFxydz62uIZgGqswe7n7R0zyrH71
Dyqy0+HS0wugebZI7rkUXIXW0zdnRM7cpiIl8NyWlVOFKnQ8MEvMwJ99JDR2Ljed
7+2ObaqBg70cBgApN8XrhVDPLZ1w+e/R7apsNZnkaRPXy5k1E/aq/r21bwhwdWYs
Ln7y1O+OHdZeTpm+YI9DvwQ8xUMRLZuPY7yxO6V+9ypsK0pZmyKGDljbsfdUpD52
j0hMcT3wYGzfcCHktaHO79JVCnW8woNuJF2xyGwk8NLqrXTeFl2denqK0juJn5Lh
okTDG/ceLE8Ga3w2Wix3vpYUVKUTA3V8HBBDkW79ejVXjhlYANH4Y4wOkJXocHC4
Ky5rppw8NNnjE22IjJH4pbftCcmDXUJQywrtZTVrFEPS/q5UvINmGiHmiZe4+5Oz
AJ/AC11lvpGyz7+bjlJZn1kHh5ukVtXhKcpCHgiOEzQ7fN9Qi6aZn+6u4pBdHzMw
hwLOw4PXeMd0nJqyzgf+tLFPMIfzfowzimlbsWBaHH0awIfaxR0kRA99gYMK8AbY
8sZLS9Ld1hrvicnhN/40lCi8AJ7kh/jxK+bNwVE5jII2/AuS1Rby15h+0FuE6occ
wAWLKOZB0oiN/I8BRmggTKm1tWWjvz/p6RRJ43Ud3v80HsooL/dVc4pUpzVPbtcK
lOxvshz0KSrAhYZbwS2EA8I6qJdHVqCpU8vhxAiCOUlqp6l95hQk9Zgign/KkjgW
m4g/noofPsIyn3R0My9PwXxJ6nQzwoaIEbggx/PGXEvsISDQkmTmauVJ2W98euvZ
Xjcg/pqMqk59+eCa5bkoIfAnk5tPsqUkh3LHQibpggfZMc3smNTwh8Y3ADEAwh8W
HORclWLdVG3v//0MfNUSqgzGz9aLO+TBmB0NEzvv5zA9mqFtBYS5N18STSMQCecH
Kyy2avDumYxk3Wf3SUqingc5YipShgbDmMu8Ga3jzqxLShb7x77tZcQ3JaKNpQse
dXCqCmVH3P1uBVsHCqrDxKlqYmQ7h/m7z1KxLQ30F2vfEz5DBUB7zhHeBqKUFsQu
Htj1gq4YcyMnpS6fCT6sG80PRKQtHni3IvTWbI17Q+/yZmqEliuZyZWLzqCrd56d
UsF/N2VbtF0dcFUji8hDHEJaMYeG9KTTa+aRGCmjv/mGSocs8akiv5FAcyfdNZUS
08Ay/6xVv8rdJS/JvpBwIE2kcUYzxZ4RtN2Op4tHGeY1G5NSrK07ZzR45htkIVwv
XFe4Q+G1HrQHto6ELwD5NhQirs+vJO66VsCe0+clJoTPcVkXNsIxNueLUk/0DJ/r
SnR+748OiXi6votqzLbcyxnKBXaW9UykbofxUZauHs9WqcKn6v857S1Nl3qRWWXt
4zYQiVpNKFvlPN2JP2tOf0W46C44jExoWUe/ZF2vAfhSFpBCVZFiZ2qIaq4pjqqv
iCDbhwniXeE8oMYP7FAeVceJc/EbpvTlGKLqXXVD9AgeRecqhl87UuLV8n0jWbf2
1ufvVEwI5oEHOUbDkfAfigP8s2eOI/MWdVIwtv3MKfcqmnR/Gyz9H28dNXwhjJVo
8G68IUgjGiY+uNAkRxADAl5QU1AejzYqWcTiFtxsSIihLtrJLwfIN6Na/bJGcF5E
PCJwFK+FG4vgIX41yNktpp9N2bcoOkdsIpeu0RFLG5SVBsM4mpc+Mewgfq94rT3U
RBRZ9tWz4fDbnLqPwsD73aL3q/sfBUpKZO0IuI1HOX5A3IXvEnxcfjQat9eMdCRz
JKMv+owLdWfBJjc4aLjtInuf5xDeEXl6hYN2kFY1OXOZx1ryK/1T5YB8ZhEq60v8
MmUJiLBSppBmYbobvTobtA4SD5FGwjpcUE8XUzKVO7RFvEznU8iEsWClWWns/lyb
PLKyrtG8U+cvfMFWl9Wz5Fb9rho+zJGq7H0/CrfaZ6JZOkOr6CWDmBsdIsOcIdyF
cvtKs93cwebz2QM8MFlYqPc2fuAw+ArXK1DEBQu+c04WK3lnj+Lz/30AgOLIStcu
xI5RizVb2nwHzVX/ZYlSpYdp8cQ1Vi/s6lnYgtkFNa4gz2cN3KVw92XHBApHQ/Ir
a+/AOtMiH571x/eH2g+Ng0gqx89KC5zxApXh6+epMPMEJ6DzdvCmuoLn7Rp3J/gA
IQr8nUorigLvAQ+NlWcA1cq6wGlR9semeF1LY3PJPW7ZMaAeXDCnDZLBvYqrdnX2
86Ilkijv4uobL3siytX2T0Kj2CemISYO9pVCgXE6Jpd9RYDbacTlSZj2zZvr9wsQ
GVvKFFAccBR4S/14DSzfDh3PknRg/5iIg95rvalu5zlvMyF/zH0ImvKVZt1WuYRO
aZ9XZnXeuB3iL39MIOklflb0E3tGQeC8VRhpTOal08exPBPUH+JYZZsy+nDUlvKO
JGMagg/Lj3v/VRdmGw5Xj5gBXQ/9Sj4JWuUpquZqq/L5nMVv2UetSlne4cvTjQwG
0ZoOC8CHSrMD3m3ch98Z4IiGpv2Q9ulFMS9hZ/Kl8c9zCwAiMmZgzHhR1Ad/6VuA
fKMlKZPvCNrv2UesNokf2ZvSufJfiU3VD6O+UPe1NBJOGBC0YEBz+mfHDqk33MxA
H9uvwU3aeNK11/DNMJ9aISkqHF7mM+GhLwqlSmxtECzrxj77W+CxP5Ud3R2D56fQ
h/fVdqo0SBHFioF8LMjjWb8zu4nxzIFimk4ZqjeUmXiHj4Mbhbq16S7CP1PLGLpa
Uuw4jH62Ml6HDzJ64u/1O33aKGoepRFmRFCvaZFglbOtl+KcegyvWXSvPKvsMbyk
9gQ5tZDVod3OpXiCVnqlmrTqq01teL0OtIFt8Xxxe7Ffk+9CtjsWzKno/7zweXwg
LGjLZhc+HIHWwh9nRqEm4qa1Ses/0KlG1I6Obi9ikE01sfSwuglhrAc2JvQ9YCd3
ynslvSN4PGetgNEbcEWd5Ba11V8TshajO843WScZ7GMn8Pdvqy2wLnj4y5WCovue
2yPicXXIW7hUgr9kGR6J4w/gr+gFeD6vB7nFhJo+ZvSJhMv8qcEs+nB7/Z3bBPmh
W23wCzebChjSXmrVrr1n+WdRgCdui5F43leofGVKPIAZufRs1Uc9dRoez4geFUu/
nj1ZR59In21eTMpZfq8XvF6XeL0edxVLtP/SQyoeWXQpPwokC4OHp42MFEUbi8FT
kmnymbcGd/TiKd5Dr2xXUIHP7VWV9noy6kCftoKHaRV9eYXgNpQiyTxH/nrv9EJg
OWjb+cIsNKFOapmht/JCixghMdpVIQkxj0AO1BSdOIsRL9njy6WdtlMnxQFvBMOV
5QKu7aPC8VnOnyykV+mZgtchPuYP+wkD9uzi7y1cTedm45p7yZ+x1WFWQyjfP/Ey
zYRYaHxZFQurXxbWnFApD9RLWzNPvHZFQhozRrme02ZEL0ZX7FDFkG8GiLCUR2bM
OUTA+/ZVbcUuStka0OQFMoQZy47G3rjP7DRLAf5uglYTWJJKq52kPaocI9+ePjxT
sik1VGnoezsgNgZPAgKIU+g9O2xEAYDk1Ozp/G4Ib94tgAa1WtQjYC7LrLepN7SX
C/FUKxmEotHdEJYoeu+CQGaijUESGQxY5P5vL7WWAuPUEivs8IPOEs4XkncNhndq
Q8hI1ioIz4sse+P/LpF1plVvk4bkeSXvukhSGoOvWMTa3/xAFEd9PoOLx4Xf/Tat
If+YsJupaH9yq+6A9dGkTUGFSNC8u0BHyFQ00ElJgHSPCFKv8W+SDk/sGV7egcf9
+OFc7aszXwcNNWxOKS6oW/ptVMmDpj2GNjyje4mPhKA+ur4hTTXE/ISry9icLRhF
iC8J52iCgH4RUuD09oJRYerdqpdobxen6balLyZ1N4XbaY3dIkxeZOBOLQyLrRIl
866Cr47A5pc25Zmmmeh36vsJoHriC4YekgWrjO1S92I00fmSUcmG3D5kmKd+NPqs
jhyEzaAvF6hcBCd4utLRHHjqEVvFLQ4MF4ePPLOST6f6WRoC8hQZVEDqweax00qB
xItEv21Xg+DcD1LMWmsbDr1lYeZbXCgz6U6hwqvHC7VEXm/PkR9sUJ/UFAqgdURz
zA776wYSyMUwejqhD6q0IPSOWvMKsReXM7dhfQPoxCXvx6nqfB55ocG+FuurwcpW
qRVvYfqfv7jGCFt6xapdMyCAHJjRVETlvAOCzIcAFcDXZ9LcnXvdWu8HikUAg3/c
fRN04wlSQWpt8ANSlDvLVgi7uY1T9vOu89ocf273xSAyYpjEUoS0KHxqUzCdsfwC
95xSyaePhZESAIzTXvJEy0b+SayPsp2D1hFivGNQSZ8m/9+SjdVnu/hIPz+DnWKE
IJ3Gs7fLbze46/uPINUBZ3KsqLwnD8akv6HDIWGKgkfMGyQMewT5LWOrfL7v5Fxr
0rzb4K3CQ/vYa+pm6nI3zL08BDDmulYiaTyUVOi5gGThy2L67u/eo/yLKgzfOjTE
K9uJZsG5DKzEcrNxV76HkgrddWU0lpV9p1k202mWWCqk3k/15DlWxo4gXGJzVeLU
IxYM/AqCvzCjgvF4A9gsUhTTBWKzYpHOOQWOJyaA3dM/Helk28PGWl2vGBADfKWh
SZEzoGdVPo8EOOdhI9Q/OB0AndreqHvwh5I2ZW0P9bBHn1mQ7r6/Hg1wFAg6Q/Y4
wotk3t9BdZNnOurqh1zmT0qMqrdTL+ECxvvLE1rcOx53tvSfm79H7KBFlE52pkLs
dL4xCqHGRqFmVNiSfbywK/VBV5s7c63GOd3UEcygbc6Yh1tSp/E6rJb41wUUYuh0
DQFR2QILHPDJ+71dQMGOpb+5YK2MCQuZBkkImO6uH8VACccTBA3vNpd/ZSrLGPb0
670iGSNT6oFzVWQrJMSM3q7hvf6tZSp7XkJDdbvk5+YKLwN+lCsO6OzuEo2ibFx1
bRBU+09I8m2qtKUAYTtC0WCzruXKjj9YRfnS4EIqmjQipubY9K1mKYdq4u1U3cdj
21ZHJFRq6sZdDH8pURw/b4wz4gH64hqU3iexjkkI89B/UBzrfxuXPNGOwR4+yImI
2St+iSaz/q3owzfvgbSgygUtiPENs852UmLzamaH3LtwZEtPUJ0FQgThggrB6Qzn
uDLm1gZdcLX2LaUHloW4wHz0Bl2TDMNfRZQ4ApzsCvmFNBZ85qiSQcy1Ne00B/Oa
8tjqj4SRXemu30a1vrywa/6BHIVyLpBBZiRb8MqYAI+NtoH8vFwYxW/dagfnHqOk
5v3w4b0RBQwdIdql3qqPzExSeyFp+DjbGpOTzLeU4rmG4SUb3yGAoNCiAqhdG5/A
jZbpjctz+mkcj5a/smXq3df/FKpgcgXoXVvXhc0JeDlELbTIBDwL3Prr0tfwaBo2
H8W1ZaT1nzQcA0/68YLc7PjlolkF32hC4s3wh8AbF7oYkLMpUmOke2AUHXUxHxh/
qBYyfLw7f9RphSNh6SusT0xRj6gSrAoMMA73WFFG7wbwOpynRt588d0XeyQtt1AU
ZrOhHkNPd22Vm4y6f2e0RTFrf+qegrYfprGNs8iwggvEUJ/3StK69niMo25OktcN
UxmPXIpSOrm/OoONJFBT9/WJr4thUASy2CrfYiCe7A5u6g1axk0NvJ89R6BgtwaP
Wz9YsJFE03GM9D9G5He/ProQ8hiG+DChMP/c87tnxmwXHHja2h+Cz5mOaVbY7lJs
hSVgMaSg5OYLmC+kP/XkH8nfmsUMx8hKNmoEX59K6S9vX1pax7EBJLFuVUUuZMQf
DnV7w2vFiS8zxBTof0D+thr7r6DiIpRTL5iHMvTutZvobuUrbFf36N69n/XwULbx
IWdMnMSIa5ntKXNufqpHQojJRdhfspTIPWjJjflv4oY5pUzGurh/Zcp1Za4SovBX
CRdaEViGjoy+L785AMAsZhbxsm0dduUody0Xx9Ijxh+y4jZuKUtdyqhEKNwhG6gm
wQzdWvZVKBw3vhnka2vcuNkITaCHaMsLNCyEyy6RNmlanscwez6+rwPGQzjom3t3
KinJsx16V27mMgQVHNjeCSQOd21xpbASUfnTJJRRlLBPVYSjXWHbRdFvmo7yn4c5
sYmHPEJGSf3rfrcVEn+4KjK/o+sG6HXLDq33eSvKXPfT0qNlQwR+xXcuGLTdZ4DZ
MtXAKZQagu/UgXfdw7cWyJZxT0Ypfq7p8hzCeTSdbCyEti5GykcbKLiUAb56dDYs
2Z4Xh7FyGrP9onBSeQwqJJtIlPEq6IfmTLzaKb0khbsZgJuPQr40eqLguO91JWwk
DKLShM5ZyXJ6YQ/Ha3JpBAioSFEkU/j1OQOabZG8VEc/7wbo+ZDRdYF8BZCv7JTv
KzQ7uLkc5dnqqpyolqB/WEDX4yB+litYXqP+4E7Qsl04mBumiuL1U1oG3V5d6AZm
++kKNBxWh30aukT3AKjrP2ATeBo2PH0eOwmx4bHC2yOTp+ndvHphi9slx6synPTl
XouHIbDNYuqfd3iGFMj/z9WnRdS8tkx2Krcrnf1Dg0y8cBe5vXvaeaDvcHa6W3wT
qCO/oC4QvYPUZr8zlfQUZfbSj9HPEEvOD3IEyxaMv/B1zRNiax1LMjYNWUEP2dFE
PbqU+xe2vtVFjc3VJfUaZFIzgRT6CmknYZk6GaGFwMuqQjnsKK5UHUozWO6TOhyq
xotQXdNzgLvG38AzkKWUbaYosl1gWrzZvZ2f78utiQTYNN1QxisR6lXm5iP4o2IL
FSnyfIG/UeXZGC3iH5P9jUMn1ygXBp3xdzZW/Prlazh8X+eshw067Hw0WNiCRdgV
k7ZVqvVsE7Vccw63Z8iX/+Jqm3qWDtQEqzPIXfi4ikeUdoYV75ONdAWfrM2z7Nmx
oGIAIwIMqCYwDLHUfP477sEHAGbWMVtT2zF2d5gF25xBL0qvsD1nZ5ERTZMajSgb
snZ23qepY8AJGkFxG/pmwOpf8GsM9g/9Rad6T2KdM2QqnQL1lRuBrHfrzGW3engU
6cFfDtrd1WUEvljlooa0WqCobyay+V6gip0sd30ktcI9jej5gtR/s51mMfIT2kk2
ZW6SyDW+EgxWyJUEYhbHCQxjZSwPQ30RvLOp9PSgH/0SAiRCtYJ3A5HGIxkjtACV
GYERWcMw7iAEtOTF3BX6kqeHXaAQHmyLt+AAM6T1iMB/OM3GJK8P6gFsx8pzbBhk
Qyf9+y4oXvoUWMJKpyfaSPmTggtFc1/65Ho3Odpvyh5SiFERV9LVlTNtB1N2bDnt
f+LGDib9tMrynJ/wWBMRwOitAiDs9sJPBHb+owj1C+1DMP/GKcu94WHk5bPfnys9
aR8RXbrzR/o6vmfBS1G2QAKddrSLsQeg1YbWcvBi54jgzqKCBEExTwHVz2Hs2BAU
a4j2/SBO4e/qGLRcYEmqmFINXQTdPYlQOJ6tORfaHWxMTtSM1N54Uk7v1ua8rmjt
FY53lJw3Nr/705Qei1cA+jx3qvf48k/fHX5YkxLJaTOsmX0v9alhvv0vUQ1PGRoQ
i8jxhLNUmi9Wj2vzj+8WWIfPaZE1f1lFI9T2tdclO8S1xWCUfYxR+XfV4JJy/fP2
SGON269RExPgo2v6gRXq2pw6/aZk0sFcVJS/JRTKSQpb4EzdeiRh1kMH10p8i90v
f5R80gOaa/7wf296HLzjC+NBDPgoaDqLGZlxb0cu1MOujl8KK/lYlKg0NxnX927m
EzIJZv9Ywza6phnkPKWC8b8SUySMwtMjVah8cnMix0rFBvNOkkEpRkGAJtFITpOF
BshOnRq1CtBE/SkJMIm55bOdJvscF8ni1Pxfv3zqblxRAmeIrsVxPMzbXU15IIx5
9WQTpsDiPTwv7rzln6t8EeRiZZbPopvdDiCAjlZmbio8bv86RlxbN1idi2eUD7kc
nAiZr+VX50a16g+/P+dZVHbehm/bVGyGlyitZokag4hiRSlxP2rtJFcMjeyiyI0X
U3Okgk0BFB5S0pIZIrKB8fDQ2pYUaLH9EBofswpl/pt0BAoZ0X52SRwGu9pwzcm0
1urEbg6rUPsbXNMoePRTslAES0oXWxJ+gfQGP/NozFTX1/e/nbyjC5p3PgvDtfdY
TW+PxjcyIEsnjtIr/StlVKQ3f0yQV7fuZi8lMWmnR3aceeyDL0tvrmw6PaDU1tsi
ayyuQLceZlMcN3ypkteAhwjOElCxhFruHjyau9wsQhjLAN/4YfUAKyVamyWqbX/I
Jbqryu/MuglDpupuyhe3hlgXBrCHApkSgJRRFPAf6F3H0XgGbFiZS3Ziz+xcy6ue
b7bC1DFlTM9qlmQK03Xqh1xcu9O/oiDEdwmlq+n3MN6x8Z5TMsFbIlltAE8I1CQW
X9zRla5F/nqK7UOHQNq0np8yx7DRd7vsoJK9vmaHBJ/xPk8fTIFtTzKGiCZskHGO
4l11tWADMeNApZjAztbWAqZ/VrQnVccGAHaMSuM1oSil1zSZrGsUlOJUDe+mGHrQ
oD4t0NJNFB0CoHQS2+Y+PigrjkeoJg0GUILeuO7eMYbr3w+uTc8mblKV9yfCm70h
XqndNFtKIocsxQwRJX2O+bsuKUXXraxicpVzP7bRyeixMtNRKnfYEJCwD3p/e+J+
E8fifDiM6Zg2zBCkYVwTlgknEXBZ7oMS1XZCYL+5YYgaq4aCaPD7i/QkmKoSnY7t
ylCQEctSgxSVZSHFTCtDS3uYKZNs95/QZMqI2gThFhWiD81zKeWLbWPFLdHe9stN
hrvt2wVJy1r9RGq8acIS2CjWsx8Hhe5UHziqtaqIX5ssd2yhIBMswRrxHf2Uz9gK
EN5DJbrFMvgctvB7HtrW8Rg7YnCdn9RUURpj3vbA21NWn01QSg8P7vspFkuCCoPB
NwprfTocEFwFVjWsOSjqK2BlCs2OENFSQ2HVs6qgKYyC8M6r+e85+TdgtsRWvHHs
Y81unWBhkNggM7XTDmKRfJX1gltIrXXKlUSiUfOJP1kIn4y/Ww+lSsCvMktz18Zb
tBNL9eLVvoN9KE1dr30CnrDp71JmZAe5R4tr/M4vhRE7A36JTb4YPaJ+tG3g5KPZ
j0elrq61ynNo6r9peRN1VbSmbl/VWsX2IozkiNaJhnHY/y1zcgWozHq+ZpLFNqHh
R5c5RsRPxdhfVZJH4LXfeQHqHD1UtRgZE2ILPvwAPJry0joPgao4ym5ZkdmjyI9Q
XwINGYVeGkiRPumCjOb/Z7taebggL7uQY9ethWDqAXvysa26HgvyI63G5Az4/3Ij
t42koxLxn1jCG8RPDhalRsvY6c8+P2Ta1je/aKqIqVupiFFV+Thrgfxx1QDWyrEN
j/GWaZA1FSkwJClThrZSBWwZhm1H/0DaPskKPdkaPofqHqqQvtq8gzuuvjgwJw5B
tyIfYqkaNpRn/gJXYsLRvDjqrqXMazHFsw9BXw7NVtrPZJZcFi5/2NzMkp42cq7l
1xqVAHlRk8qUIgPB8848QCdpFiXLqWJ7hrYLaiqiGSUe8HWD7lHG61cDQ0c/XX44
komX4TG0+qtE16h3HCgihm4IxxJ/TKeQYwjnsOJob1l1OkLPgTpwjiE6FeApJ1Y+
+XYDiKjdwdiM6+vX6/7pjKwusoAh5PnNrZMTRv0KhteSinQR/g9ziajpqh1dst8q
MxlYeIfgwsQ6Hss4GLRb8s3el8SG8gCVHM3ohfA1AAkGPgyJOOr/c+kXrJ59r+j2
pvZBnMCKDmAILysG0fMMZ1XAoK43+YP63dEnc8W5R58amtqEBPawT9F8JNkF23zN
pX2p2xJdumoeUifVzqj0drKxmDHYYBPzbKLTICod1Us9usCuxNl/0irP8VvjhvHp
fTwkx9oSthuOEhqy4sgjvOViMlfIW8OHN+ugYYcdwI5Iq50I28lQmQ31qPp+5Ypw
cEp/QrQP1Kxj79+ppvFIZzIhVdKWaMkg9EwoE8itB60gFtW1kIIS7bmlQifxvimL
D/ij1N4W7v34Wv09AaQeAT/x+7A1In4W1KH4Iq0OsQaMEVzOgWlH+XDuzL0AWiP1
ZM8FmMTzHlBaWSS6Zm7fxRkz7MyLkQJrW/kItLBT3GXZAfPn7qF6MYqVfAFeDxUp
EE24BG2V5O2Zkz3XSRMT1Q3mrjnBZu4UPZw1/1UWsoUBOTVLrjI7Krq3/khwa3H8
7Riq0LStESfY513nPeBE+vmQVseSiiGAS02j3bSOztIAa+OEw5uV5Enm3HDala9o
1ttQNdpEqrzb23XcrSz0h+jZjUqhvI0MX98VokvhFQFvaWMdum+DTcgVp+0mqEcz
MxQkFtQ35zPGGrI8XY9n1UGEHy+4QWuB07RdK7bATf7N8fsczkiLJjz2Z0NTTfKN
dZKkQj+MWPSZvuSFCdiE1BcqLGY1uyhFxfXmRTgVPWItf7ZtEFEsCwg+aoqW5rAX
7C8garycqyYrSN2NkxEiikz2XFktHmsMd+Wrvq/MzzlBf6S2bXU9Ztp6sExPnMBx
koI6MxdDQ/22AwU/b8sA/OhhCzFF/sgOvqdSCJJDPdql2/Qb/VyjmoUoB/4viSY5
ADc/qnasGrhPKyMtC+lE9tHFdy7Z56SC93GZwX4u/ZGa/DJUeolORxBBf8fAGp6y
z4MjfM2xhRJfr2FRRtzH7y6A2Yc7IkM9qILzojS07/753P77vSAnluEy3KUmkEMB
1CElT7jkOmYqdERwW1XtX7n6+5ee9DBHKXf3iL+aHEQkl83dG99ZDQS7ZAmiwJ9N
KY0f6v4cK4ILIKQEZq0DE+j/S96AlFyXApQH/sdCq67P0xKOCyXIS20KH+JwbSfn
IN+cAu5IaA/LuXo1LfLV7t33kN1oFjfO0gXSaOdCchnyxb5AuAi4V94O8Yedscp6
VjHOU1hcKUe25C715uEFjIgEaXqFNwskhgT6tJhUn4AL/o69BbeSKcWOTS2b02DH
rIMNO6DPYDwLsM1Qa8WxxkSuPMvm48K3wiZ/KvFnA/EQjsmhku3gtKZ3Tw8OpaOs
PmCfIBardDldY7ZXX9Gy2STD/qti9q4A8BWWCgcSJxCxiyz/iRXgE+Ub9VDBi+Pr
H8X2bsV4AE0xXvTHgo+FHr2n/Lb2CKBReMCRuJMDPt7h0oEyjJBj6IZ0dQ3oD8LW
6YfXwQSkKC8TWz7uCKsv1sFR3F20Uqa4wdiQIAegT/LvCn8pPIdgPj3XT4TNZvOp
xovVfiHbDMjs5Dp8XTvEgSSEp1MF/zBbkD2V+JIBpa2vMhM+EiMRSe+ugEwHygl1
XWOe3rIfMqjfF/Gh7iQtR0lVCmCH69gOE8H450PK/KOFfGLHWVZ220v4ihghBF8W
gLYikN07B4bgR3i8SxpWiJatGo/yUlN3OlSPDLHJBEJh7YdSnmjNgbh1dI65ZLxO
MXZ9EKVH5ko/YOuUM8/WYkDdCLGPi+9lgkFRPzu2bdFwt1zKguST9jfIAr4iDYFY
wggyx6hgyUJYtq8mmrMxGgnUsR4oV3JQOnVAgJ1+yPZLQZzEND3HtTBc5gIphqYN
9adHNb4TeX5xjsbTFoNL7D1AD4n/HH4Z8bLK/XCbpqeFSZ4lTB048fYiLRwPrTul
njhQIKryU2FdpaoOcnY5kyYkxXInG0GYO/PwGjs4j7o4ATDMI/VhlufuGklxMALt
4/87UaHESOCJu2qxSakO6B+2KASJSXqZY41qgpCW2sUGxg8VGl/9/G/APkzXx68n
KKTfyAbehf+2gvpnodRiEJHcB/1Q1kZJrdcnkPy/LCujW500FTq2/MC/1/X1deJB
/Aaely/OkfM1ehvGOaJrVH7QFjhT+crWs4TPhFv/vAcgiyrk70YTvYM/nitNDxpc
xIfQIbAhgC+57e2/RFLkG/n/Iy04kZDuiwMzyyRTvhFZK9HteOB849VwfoP1KCH8
to2+dxj0N91b4JOWRiFvQ/M/cOCxuGzbBxgdTRuIKZ6bQexMNFRvVmisz0JlDdmD
Q+zWzpvby2SN9LBz/L7wthLnpmrr/r6SWbyB5ve/BpLIcBTiHA4gNYEotOtI+nfh
nOTk9yPWqcnAkmjcJKainCnc0hwrRipQZTqDecsKdRSFII4uxIX45EZQ9+kkSplP
7D4GQ5LVg0JgwjrEqME+LMNNTNTVB9HsTygx9BpHcz1yaoYmCtqHS/4eutwgQKCV
UBuxNOHEt1piCzvkxyvEy2TCcTMPVYxo802peTxqDVIxykxtesHcBCTcOe79xvxF
82jsAEsvnSBSI7mNCpSSQyBP/b+eez2+bKFKaWOazyhnuGor1CVkXdA9co/3DWiC
t3rK/u5hRkJyu//B2nAyx55Xx+Qx6aDkmp49fxj3MUBgvJHwGY+6TWUPV8YpiCEl
Q2Hbf2tFXBTLKSN2Ot7N0ywfzAxNFZh0HNGhBgfMGAnN9T0cBEeCJr12c8b3/foH
UqtTF0tx3NdxP1jtGddLzGdm9NzRMhbrNMHcKRvsttNwSciriG2rfATheWw9lRER
TyL36h6gQEg4Q9C2QaofIpfH0WQ7EShWlaZCsGBxfO1P8Et2cRD/3JytQh8JJGjw
DQm3phP/4dCqQ8B0NK4B+YPg56OcP3LuK8XzgyOri2KU98bdwXdwigOleGjEbV7C
PW53Bi1w81uP/rEiluKvMKAg57+kwUnZE0a0yr7UZ0cU8pR0pWp+gAnTGio9LD1v
ZL+V5lzhmajsuVloeXmlKkfnyL8LzAnDu5nQLuTEpYn5Qp0/hG/vA2DZrraSZYmS
3iS3YVycw4KPofNIX1WX0uvgM7vBTYm0NrhIN+Vch+fHD0AHBfZwDkACP9EuCEoA
oFqIJLMqPX3DBQPYh3dvVNcv+iilskkbAwQpIkVChuo6QcePcj/w7S3VgIzirkb5
oHwz+k5ywiGfipA6cw82NZ9qoszX1XKk/u25/lqz69BmabJysmOEFYRVjkMqLSvu
kb74GlWy05hC9YqsU/zNSrXWbaT3PGg02qDq6GJXEQg1KCS5osiqa32cFAAPswWD
96wTBtLG8i3X+KkOrih5hVC1oKY9nQ0q0z4UebGFphMjrufNZtiS0NCk7EBisN2q
q1B/iW9T61/BX6DY+wvHDmFb6orvlmACS6LRcrSuAhbOfgpbxAeKs81xZMoz8D5j
r8HCCiEq1b68hDp/ybg18LdgvUiWtYUQhy+qC85gSWcfRfQSDre1lsGnOmBARKeo
s21GixJFCD4v1cRYPOMcAc4DsPUspH7+4YRFjMEeWde+9bolz6qSU1n2GSIpzw6m
J8Bmz5MWDRKo4Lz+QJl3/ui5H0DvphNkTN5wd/RSC3qbdEh8JRfHn/dPoGsPZEwJ
RGtJ40xvjKi+/mFa9cE6QmFqlcFh+7jbchT7je4rN35IdV7b8qF8M+DZUcr60Ofq
EAsITwNAoHnUHljHpM4mDGhYerf5g2zFTEg5hg57muChVCozWu+HPFgR08lLEzxP
dXhq5pdE1Gm5XBs91Z7UqyvBYdmgYozNxZGNCUIoBBPDDpmUzLCnKdKG6ez1D8hg
UcD+mAjujDznmLlj9X86NEeSZc+cc64yrZMMJJDLPTGxq5CxxvM7wLB/0Dmo1oLn
Irx8H9K+kbiLUQDuwJn5JXcS96goUEUTPccHDxU2m2U34/PYct7Cp1ZHjAd9I0zw
ru3s0ckrm00+gWG9PXRhKDsuXbTCEkvlwlL+rjPd+vFPNswtyMsYHZ9OrxlQ8zZr
sCwxwJUwmSZNf/QyouGhuw1eW7S3/QiZPaNIrwTqfChtfcLiQvb2pMLmWxXOkFG8
1Ai8GPLLOuEpVmM1nRTqKimOOfP/qllv//GdsGLDTQ0Cf6Rs2W1EcShS8+zEwwvM
NqjeJ5pauEjPxhl2aQKar/iat962tOxHt3FSjrJK4D7eOHiWAXpi3/vFfIb2FMcB
9LfzevUztJhMuuF+Ro/4HoGxxI/68BvU1ujK18SVgUmZCR3Aow9fLeArOOMj1FdU
gReYfDnskUiN+eGBY4m7atDELFClWl8mca5DlzC41nhIEQIWES8pZWb3+hcoBM3j
fQIdMbrg6pS4/NaUo6DCZwcFHgd7Nx4kpzM6fJjdLVrr80Rhe1b88EToh0EFkNyg
Co3dCcJ/rvs/dr+mGrMxJ2IRH8ypXdlT+6h9xsidtp2zlY+VRVShGLEAZBaQNt/d
fbIqHT/Y5Lqccwow2p2xeFHE4tHGOZNKTBevNFzTmz7jVNCDispfBYnJENZwnKcB
h+kzwENHeowcHNdye6CgCwqIGWVvRN+TmNfBo2KC6Rq0FjSrqb3V+coZJ75l2Oat
zegEs/9hAJ/XJhpVGQ0nrFsSvAGp6sAAWidwmwwUQr6xTpNZGEDlWFrtt0R92uwU
hyvFab28kg/EzRcO3kyzEPMsnbHwCHx93Q8oNPloKQmd0j4BN1iEctUEkIcrssJ0
cqRsC/a0GMMQV8ddRkXxPO+3MQWgbJWuI+1THxTYLZJHsN39IPAD1TaAy/0qnCDi
ANUH2fhKZy5C9intb0V2vR9hj84t4Z8T+XPVHGupXFeD37ovIg9gxRFptDwJTgVU
Xr+Rt0jRtkmdFWurqrJJQbT0ejKqN/jT88AC7Q3J6BgMkxIXHt8Q1BHblgKRNIuU
x81wO60wODxLY+G0O54XW6EJUOXfsL7v+QMcv7lDklyk/y1jcuXVQ49IkkjW0XVt
Gb+9aJJO5/HGfTlfDJwR/yw4iOnkBSktjaJGsZokC0oM0C4efAs18yg0PVxWy5gL
C6TM0fh9xmiYVgGubs5oLQ==
`protect END_PROTECTED
