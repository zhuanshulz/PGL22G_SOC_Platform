`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0k+imr+VwB03ommtx7FSL9oxJ+u8m1kg6YiyTDPcNcaIp0jFnkVgODVBGV5sacPv
Tci1NV+VyKL42o5MO63SfZkEL9CkH0cH7TvJ33rN2O2Drh8JHmSmp3JLW2nZffkR
FlCf1t8HxAEvt2EpkjhefMl0RbxNxJuNgYEPIQHeybRSnGGO0OCi7eWwytUUCoYY
4rZPcBLj0Xcnv04oKHu7eab6IL0U435JBxQEWDUDakzSMkRv62z0sl3xCDhzGn1y
0WpVSO6ifzsLQrKyTiPoxcXyjMavw8uJkR4qgqcwfvJqAVTZcV6J/LvonA6NQKaK
BHImFvIpsTUB7WJyL3fQ7F7HqdCSw/lNIbRGapAQeqC5r9b252JrMKMrg9vRoscq
6Oom382U+f5/ks2yGHGpxHCAyfgag8QVutTdqRMxfmdbdpT1DLIStBwhYo7fsCL2
iiSnZc2zN83vyPynYCxmq8ga6oRz4rOia697rvWuc/fqpjtx8pAPWbpkoXNMFj7Q
aDhZqoRQe+1YrrTjzcuUrPym5ooylNc0Lh6P+UE+qoPlBMLk6c/vYqCKw5aiIEmu
5xfZ61U/Su8FOFZV3w9eBZ2QHa8HjqGbv/DcM6B+ouA+mS5wj+WsS+cqPYLHHcGH
TJQP4v6qeeWh8Qc7sPZWVkQU2IumVJn1tbBJzSdTGahxVi0nHmKwm4UTM0n/Y2KR
ycxpLvhO2BqHFRhnhE4NqzdTgY/Xm4AEoHkRKs0VccMucetPleOCBt1XQuGevu4A
mD2VxUzH70YmtLI81iwhSTBpPBBy1fkoJy5rwJg2yKKYWzfMpjwwo71wDyxLtxQX
Bhj5Y7WKNKjvqgtXd5GBiPGsvfo7o4SlLz3BmNYDKmiZnipUdACfA/yI6rA2jDdu
HNJhKuGe3FGI3JoDVoxDhgpyDd4b19ypvbo/civIkKVylnwFNKqRCSQ2zMdaqkxf
n0tahDPqunwldJkXlpWaGK1C/r1tC6f80Is1Cm8alAmyGdNzuCOpHikkuQo0vUAR
z9VVT460cspnE8MyXZQZ1Gzr+j/xxQdMwCfe7SE51q4Zl40h7MLvUyIHxqHz9ZvK
l+/P/JUCNPqYbsES3AKveX5n3vVWLqUHVJ9sdBs7b9yEQZnvzq0ACKtBNwA9nsOV
JJerUwf6YcUajm0sygFuCy1ofDrix7zMlmkfzz5JxFbFJPo4rC5kyyCOW7Yj932H
`protect END_PROTECTED
