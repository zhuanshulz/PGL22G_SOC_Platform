library verilog;
use verilog.vl_types.all;
entity GTP_GRS is
    port(
        GRS_N           : in     vl_logic
    );
end GTP_GRS;
