`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JZuJ/RsCBf9fNAEbh3sR0/TNWhqlaFNa8la7l+l2hRpaCvxuuO5OOWZtJ2Vul/C
JyUnlPQWp9MlkWKDqlyPCozRhZFjxPDJN2LiOh5SmaQk6qDaOBgJ/7YkSVw6RiCX
I4Okw1i2/4c2/Jug2Jvnm6/JqLk24bdhuzrdm5FXPC0W+IPe5fC+NZyu5klSA4dy
zL4FiEe1KzewNJdAELj6A/zHC7JrEH4+zz54apl9DjZtjstM7CR1r39MB12ux+7K
zCLyT1PixBX4Uj8jm3onAaboh42VFvvZU89YTqjbEjRTvCR1+/J5/fNKmTo23UYt
wj7yh8q9ka+5eKbhnTAT5FfxEqyEJQRAbf0WxnnXXDbfG5k26fWoTrWrB+LMGdxZ
XBMgC7wxevoH7XDaiy98jlXz8FwTARsXRTF1dac/qDkf5Rz4A5jYb7h82AICJCTh
r8cUJU+ZpxG2zWk26H/t+nniliHkwkGhCDIB1e52gQob+kw2Lv1aYA01Bf3GLuu5
BFQQTggJ2hZsuYU85ZDwQ99375Ju+8g2EZVWXK4cnfrORpjOvIrNuCtemFgJJI+k
d5GGiXbHg9/LL10s2JPkbJeogTrjmPNC3xyCLXptXpE1eHvysAGv5wF6FJkfnEhR
rzWwZsLjr/4sFrdMwUgvSuxtB5ye4h34n/rWfnCT/wiCiFnuXq1CCKoIFmSiTLsB
tbrSyMRj341GBt3W7iujMSxXrqSp4OyuE+Ys0HX1j12iLseNSVO3Jx3awL1HLQjX
6YnF6TW8BvGTz+y/cUPVbs5IrfmRYNNZOZyrDpLWXmAmvVXIZ9JSpEJnIHK84XzU
JTUxvy7BhhHi2+dJhFqaoT1CSn425YDaWI1TYu99BxFWAdPWfb9brK14jDPM86Y9
nDXvfPrdYuiPrImAZ/KliGAp0apOxPHDep+JAs6pwLJ0OMCUXtqY5sPXN7eUDNAV
dvf6/C5EtwmzUlH4nQNJ7kt8T2rzykGdDkfUaeZ+KVng9bpw3x+BqUII+pc82+cM
zuNKyNPcGNggnaC1hqZoS+h6Z7T+8Qao8C/vy5y8wm/MpRzwe5NWBwzTZZqQYvd8
tTeH/NdHrLcfeaHzYux3/+Ke486xXKMbmSuXnV/9lNWhew2P4PFWzqDNc/Sea3l4
Gwl/IT9BYl4WGJ7tm7uJpN1jUEXsmHmt9nMJHvL9BFZiJ3UI6IGofAi6NPzqgTQz
rGtLKEEaTMJlhdh6xmnjtG7KxUsb8Kd9gCk111TDIP7XT307urj8aoZ6JXU9sKhg
jrWc4ytA3BCI5yGPLruDb2bm4ZufS3gb3BQzwGTsbANkKDeapjNECAYkigPZNG4J
49pX9sQgqI0GItYKKTC6KVLtYecH4u815brN8Y1N7+9NeIUnNMJuNdB9blrxsMSf
CqNssJ/zpijIC+bQjRfcSqf3gWjzFBNtX5PgB0RjWERGKhtRHBPLBxNsUq33Mh21
scNgWsEvW1cyn5fYVkD3ZYlUgCw9MeeRhbxbxuLKRDZ9j/Vk5VDGhmgN+DTHQXvB
EjBGPFhR7gWrMa1bUSTYdS/tC1vO/a9kEWcNIwm6MxD4eNyJKT6OtYcjksVgrsLZ
oz1PFEL42lyBR8s5lehobNCNCwbCn4yA0ymAU4Ym0+pey7SS7inSPEK90BA6pTI0
IlWwDTzbz9gGTlKfFCNXonZfV+ynB3A71RNtDSHhHVEzDy42sqprdheiV9a6YneC
p9ZmKKosUss3zM2ot2Yi+GlPQ86dCgIeUYLeJqbuv+9V4EFb4TkMWMtgDt703pwP
th+iPwAVEPp//YTMapmP/Syd0T5ukKMPyb8jpk32+Z7zWTacRGYopw0tJ/IM4VtZ
5BzzFhuToWbbRaFcay1BNZKYYsokLHDNnQ2gJTjAR7+67kdXXcGWMiBF3x8HVXJS
TmQLxp2hqMk5yKgKVjo9oGwNbP3diJodtYpfSM9kvjchp/syYD87UiB1JSefirU1
QzwSgCejAwbh7EOMM7SkqwJQVMWFdOnIpSELLPcr3nvyoXUDJzNbX8Jd8FxJr52v
cB/H050KTahVqOb4ZP4PgYQ0YsXkHBHrvoVAD+G0CcVAbBJhHSUwFWmrm7AVna+N
XbUS5Py30u6CV/scMIhpM+x9cGFcBpCVJjCP5OHx0DTiEu4mLFkTaoN5e1nSd8oR
qouZkRUuYiN5Rr1ZI2FDtIuibIOaqJDK4OZXM8HatvwRRmUdRR4Wf5cV3g5qIbbm
7eKAvDFfijZtgn6+JNRZ1l3K/HI75PyQKwhIA8TRk3nrdE/0ZrLAXGmpASgvXcIK
3Bi5RUtumGj/M0uTIlDTWOXdz1lQbfEoNJofiSbihUuhGOfK1GTWkNzcsPLJYsrC
uEOxH3cmYMUmX4tpUw65oLTbGAHQiA0Us7Gjnq8rAfyTbpMqZo8Giidh6zSmlGQr
tBAd6rNrCBm/mWaowUUEvM21glDGyB4smSh3XSfGcQGykEzLRa4weu6Xn48nVZWf
db2f90rCweMiFJqlAyPKR/Sm0N27/gcA35nOC7NMBWmmrfIvDkfMOl8c8uaQ5326
CP+iwwjcFuOaCNJQMoCcdNbzRqk2OFyuDPtQRVHwBLOB7A0nSNhBiNZwbFR3Focg
d269h9ZVVc0CiCL5hTtOKZe4sBXEeGhNx9SKj5vx1hjNFGlrcCZRhCsxdSpT9863
7zYdkdzKVLywWAvwN+LPkaoFPbXAtvIyC9hTg8Gcj3Ln2ZrTSyPSFGClvjWlQ6KB
N6BTLG5bIDJR0Fy7tkqpkaoSEiNZfCikxay9eGnO7JYztvdJL2WESJ+H4oFCpWMT
6vPyurzB3A3WxHN1jAH4ate7CkwrD9cCUZfR0pRhvLEjynK4zMaqRFu1N/WWbvkQ
BiZqsYsllrU71XgR9zkgSqnhvOgbFFBsU13lMZ6IbXNfNG46Yb9AZmneZEhThKbJ
GMnh/gyLercUjV+uaaSfTVllKrUpz+YCd07WND3/uGVGIco1pU3N5fAWF2nU0DSe
rO6BCGjYMH1MT5ApyVXR3ZuTyssIMmN4Jn7mnDy2AsO7XjKkzREo7vyqwZ4rtvNl
+z46l0MD5CuHyUr7J9k/xxrce9RyqaAu83Jg0j27sp2BbqnbisMrDN5m4ldG3zse
oiYgew8yfZRC4SXrFcxdj9ZlOS5I76Q2LuAX65I2bctkaarXtqslJsm37duC1e52
n6GQqx25e2aGFchaWR5k00Ee9tP9fMVKbLVD+sSL0JkysZ3Xf2rYJsmXjKAeccuQ
YCtr5mRCp7pvkuZzwHrqXlHkbbcbaie+0MvBy3/cRGfCwNllbBECVccv1HAsYa/7
wWMQzG0PgtkE40ABF+gkOnxQqGepGo0vOTdk4mULvd4Hogn4WLghjl6SSJLiOe1F
yMCNGZZK52Axqrxpo23vtTM76D/bs/kt18UHv5D1nKTKIs6wNmI/NEq2SrWiPpjG
+b72aaIF8Z41dBZR/9HQgiOSigl2PvH0ei6pFzhjFqBCAEdDxQe1RdfnyhPIxg6T
GgpAERsfavV1i1yB19wjjpEBA78Bh31+wo+w4IwVqvsCY7+sPt7XQEdSmSY1+Gc1
1qUxd2UfUi+qqzcur41WYdSOJ0eisabADFZs3yw7pNSNN8nq6PaGjh15Lx5DcuFg
DLFFzMCYG3ao2Q+EdzvOr35/h9VkJYET44tmGQfgPJO7B9Oa2IjQs8vZATyvTIGL
t4Qp5411BTxix3NeLN7D8jmrj8Q9M1F9CDVMXb/V58aCcJom5hVLb8CJOJVKQ/Cn
zdj5lx1F8YcaE3a79KT/YNKtedLHQJmUqHj35gZRAXYg1J3bmAUBiapzOAAK72Hs
T/STPoZXjbrc7R2pFD99YY/JcyCpGyltBn8Bvw5Di8/2i4df9IALhLPE4mGACfSr
gZ3AU1FBc1VUbKFQ70biScHXHWg5zNgpkdpSmHvjGAqY6bVaKT3h3r1moxiqQ5Kr
1y/3Ix/dP/EeVk/qPM1c1iaQ592AKQvSKeM/v+HqSMk0SYJalVMg/A0cM1u5kSKN
epXkCWKJIGxL3eW3m14ypwOFPgI4trEheL6bZMtmixFikiS1NeT43r+29QKGGVkV
zzJN75mYDBmmSA6YKhVzLBnlJBNIb0Qo/71ijNmXUNLyoex6vzWxllxZibwYIQgn
7nH/BMdK+qB1/kz1ZFkrFLnFRMf9wstOvj7RRm2xYHCrUCo2qZDpZJEqgPCnTmiq
sp5JZXXrJIucGnLdkJZLS/1h1yZ0myxGRDgJx626hv2/WCoY2U2U8z66x5AsVmMp
scPnnTEoOszju3lo8LsvQlTtgOa+25PIzrQ5YToC4XviGl0il16Cga2tJg0K1Tf9
qMnmKK/hCJF+4ovjF71sVbAfR6A7V3RDxQVO5mBpd+FHSGJhDfIekU4gNhioTM7X
zyq2Zyiwclvjxl7l60JDuSstrT44clpY2ZR+IZQLTGh8UtZ/eq7ZILfr6JnDIvLf
9J/vIQ5Pae91hyNti59XW5yM1Zwqn4qg1C0Kdd9drP3NJAfXzuAsjzmAL1MCmVZw
fu9oTCOQiUqke6zxwDpgw6irQnHBeaGhfhPlcpK/ZvZWkfuPeSkQkxNNz0/k2CUk
U9ZB1w6zgUuSD+Lg83RPk9EfRwjRUv2nswf+GuieJmvSPvvuoc721a042b/WIaGn
ZwtwLOrKjrWhjxz/0UXh4Uz3eyBEpSQ5jGgw9Midt/lJlxiF6IwsAc5J3g+QnYue
CUPikrE08H5nAlgJIBN5oTUSiYHp/jCAqXhjWcF3L2M+RDB7aV/QH5elFzqUAJeT
81VDetb616s1nvkWYuaf//LI9Mq00AtytjK52vPhTne6iMNPEn/siSmrbpdczDaE
ToPJ+wKuQ/fixeacrHwWCFbAD6QHjcvbOgDpgcqze5X6YRoQRPRYth5TGx+Qs6Rc
T/eDLUjNexC4uLPn/CTohCemQugfhKd2vlTOj62v0TD6aX8T2oDWsj6F7xTC19lx
dwqdAf4O+/J1XOGjDt3ipstxYZZB0jCwuSH09860/ckwGo+iy8XzpPYOAKg64/lQ
NtB80oKYXfNRufyI/h2wenoQvzyR2qYJy5D2GvmY1EqnA06Qe+ZdbhijrbC/Xreq
0R5iHzyKKycCYmVUg1uutq1gL1yOCWOo2wQi3IaCojmfqYx8bqVP7I7PlGz0Ok1m
rFqAIBiv1BuZdlLlcPbNEwLMq0IIkGVep/iv6TLOcRXjumheSmwQ/l8LMcxMHnrn
jKOjTpHZDFnqwRH08pZpnLcV0Sc+pBOJYAdU6Q0todgcfFRYQ61rwzKxt1iUmD6w
2YCNPS2Kwulct3BiepWPrGL2h8idmfjTRBBMtmqx1tCBwW8P5cIK4JgUoZmHIazI
2uBEybxiIRu44NU/xlKRbZIYqrqw5ldN/XDittyLhnrHfyUA3rIeg39fcvBvOu+x
Vj9Q5uwey+ALm5jrNA//BOU0Iv404oGgBvOQ5xcXYX4KIOyidO7ToaG+bUJKUiTE
ba48KkQ+lmTQvmIzCBUsdkI2UhuJz+qH+h8It1b1EQ8honLdDJVHxXF9jRLixFnj
9+OCAxnZC0TzfaaF7fXUL1O3clZPE0X9KXVc7ToSobwUHL4n5b9aE8w0a6cVOuuP
whKYW+cr8FLXYTyAwhcbv/3zcBDVOEsuTNzHOBppiYPyTSl6rHqqdMCjrkj5IC1L
bwMGiypALf1NFdL1ijGTMCN6mNSsFGdTUXvAOlBXWB7VI6M8aH8dOu5DhU/cTfDB
t8fd73/RcrOGxrzbwCGZH03MmOiLv2QkabRhFoRD9iPdyoktMhXzrIq0SjEJzEIW
X65sDcx4j/kUDlL4dC0gtab0BdO06VSKsG+PTCcNKjtXJjYIJ3Hqr1Q/LBcBDdgn
KgV14f+ykx0ERN22MjCU570hI4uUx1L0DHc4Lq70i/3PGJjD2u/2utMzc1daAeyf
NY+5HPiwB45UbeJ4W1EU34WK5dmHFy3kg0aJY8yqwB1Z3zRc5fSJwRTsOwj+GWzt
RD0u+mC0zBxNOOldPprFkoi2b6BZt2XyHGdrgtW5Juidb+bfd7R5iU9hjXbw9nkN
vz/YW03MjyUPi1i0F6sU/sY0bJGrfSxW6WDMHsMy90zOcC+MDRkoqgdQ76mxabyZ
5bay1hS1e5jOBo+iK0uRGhZV7gLzW0QRHP+SH/9LkwoDYCn9hTCyTP/yPtG3JbzX
J+fHOP5tHK8xVTOebJzTX0jpa3NNysZDllHUsbp8UF05WGezpDHyOZhMYiNsTF8A
8gY8wsxpSubJHaKLVr56Hwz9QA8L4X+SNJ+05tecBj6RvrBasM+U1HbYdaBRZ855
nGR+Rkpt1QXXuPrmN4JsCq7KAjWX/etu6OvzdTgZXUdTJU7LIVWyyJ3QMVx7LdPL
2UpJt4t4KnQmjiSfHKHiMbwlIfV0wiVfDOLYQ1CCCrYgJ3TqTEc91NEidMH+r916
dxlqaHkVEJnnD+ahnRT87B7bHT9eSJkMSfmQ1jcTqv5as3eNJWnRTf2KwbqMYInt
zBO6SOp58aNe7RptPlynSeFwCzf9wa6mgLVyfL4FIbvcmOK0wP/3J6/qOVOA83TF
`protect END_PROTECTED
