`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
54KMuTjYdUsa5Ma2sdplqOZSw6O0x05nKvUwHQxM2Tdv+0R+hip27U4p8m05MiEf
rRmQEatA0cpGZ1KU+HibRdXTsVl0eSkIK0cMu1zlyqQboaEooc+sWyC5NOZcB4eS
f+4/ppOgAm7Eq+Kn+eX5njatVVCClR5+69bO7nzJPVcbmMwPI/ODxVgfByKGedSu
7zuG2F/zmd3DQNiJqt0EKvxgRdgiWVexO1ukLZgF7GxeMPpdSo5UpcF8vKRo4f7n
J/jxPoTVWjpS4V/1JM/6RQfPJFe1TFjRRvw0KClATlLjhMbJJrbnFDIdAiFuB5xo
HuCk92KHcWT8jJojcvXfo2tAfXX+wC1d7aQbjfb5hE78w1+/P90dCreO6R5cjzLh
fNLEdOVuJAJfdm5eK9sueelCsJmexAooTjA5eoA6p4cIMvgn6JmFWks//PRVatNY
I98FBbLQdEQctTJCtxsaag9OeYYnlpb2PuN7ceoZsE+j5p56LthbZ5WJXoGuOEPE
Q+E7ap52JYcH4JYF2XvcawgN2SPsPB4wGMg2Q9nqBq9nk+O9f7nBsxaaOLZE+8Fl
dJgWvoTfvl4VQxBKCIRaYOv070/1PCJWz+1G51q1vHRyIud7bmKwIQ7NO25UP4ZE
HwWrnZF7dykMiI2RdfeXuEvY5YpuKmnOsHIVpxiOz6gv0mduoi4f2DLpVdSZwLfH
X2pVRYAgDGf202oaSQSOT4201Jf8XDdhQDBhtxgtL4PIHNFYd+zIBZaHR3fzrTAB
vDHhB1lWxFihaPOFi2v7q+HUXrdCb3Q7/SP3/kZNnz7n1HYMDaN0lJnXBRUXNuZf
obKskVdmN05BBFtju0nv2kIEaCrLEiJQ7B1GTeYO4wRD6b92mZIeM0MCOxsE7JtL
xj3sLne2YREzUQiAXeT6nhbM8JUiFTa7hCg3sCwVNJ67Lytws4CckimPXRPONdeM
XMRciGgfrq+kjAeXhENuljLihO/5RsSnvJ8ooCsZgyBLK/gzx9Cn4UV66HjgxsBq
ri45VQRx7K7MNGB+eO/HCzM2LZ4DrU7Tlg8Q4agm7/KcsNgYSJPCwzsXAN12f+89
vT6KB6DimLTcU/o6Xho10P6CCsj0t7fk8coFjd4skjPu02QavQ8dKCyXdkGe/IK+
c1jFhQHj5AIr6KlxLaxj/hXuqKB0l9TymJCSmq4XCMwqY5/I3HEJd3yJ+TkwNqdP
rCH9gvuHfeA9ltFF0ZCHCp5bH86K4S/XYeL8ml46qVjhooSENyt17d7oyKVBKnae
+na6FPzh1Q87BlTd/QvKQgCjIWbA4yXKWFzQaaCXlGBJLZ/dHcaWE/ISJRv6aLOC
T7dQ95YGK5yBYl5rV7U4LcHRkJjVm812mFfsmnU5AtCkTJEYjPc+4YOwVpLbmq8F
BeWKNrkvtemYY5uRQWa1vcD82WxPltk7LnFxug0yEAIob1Nql87IRGw4rgyyO2CC
1P1hBvKkf3C6BJ69baSznsZjUPtlpKHSb57McxfvBGi7ORTqOBb+X+P/AKOQsiLT
p4TXwOO6N2xMnh1NlWwwCDdNw+UvOltjueoqtP+uBIGRILqr+V/5kA/zGGtSNioT
oDpYvhqo2fD1270aO6hBmGe9G8SK0LY70onWpek8Dasn4/oH8IlhFGhZfsja7shL
e02sXtIiZJ5wyR63DZ2JpB6zJymLd+e3g/i3OohlqZbscSjYz8P4Riovy0w+78hv
C2ohq1Jb1r5UysrlC2ZEB4aaLPNIUE9HiBtE6pBWsKgJPNDkD3cmzadpVnss1Zow
8dkdJ8gCX/aP8nTctfmTELCOzslb1AOjSMiVotUrg/yhg2uxPFkFi2VfiLnUaDFi
fp7TE0VTK2We1zvSmcrvr0EBdDRKsDKqsMn0s3fHC8AH+OQ7GViHGgGaqCns2Bgs
0hr6FDdsHx43M067s2QWUz4yL3+diQdQA2sG2AcI15C7ghVZyYmU4XNNoP162zCP
LX/izfeB39VzCo9YCFhbp/TT0tFx8ULdD6y97BXOllISUNZRm9Wde2MrqOWetp2K
xEUAaFYVz3KT9IlbZ5WRqQqcc4vuut2T+inrv2Rhhl7rEfXqq5m5LjcUX47ZnWJs
VrBzlGNzvUIBHLZVM784HkGlYjBE+5o83SbBSdOwfKgVyDfjOirNbeAo0SQx7kVj
IjVESoK1scm1eyE3wD2IZ0Jq9/4QMl6HeoVVk2MIBok+LE+rAKr5mYCISaS1RoaY
B7SizicsxQHQkfj+U+YV6AgSx8tOYdQfkA/ODGKgX2Y5E6GcfrqKagCWaUW+HVQI
fbWoAX/UCbBa5VhdKn3vTVZOHBQPvkIT3hUg0A6Wn63Zm02J5efmGvFZ+xUPYz+s
lHCTE2zKn0ERwWGdaqvrxPSEWslG7QDqfdgPUJX4SD0txdCyksl2das9hINi8hLc
VssYAV5XmBEmF+c0vM+ssSkQrpgYCW4IdXrGbCYJW7QU0OtZVNg0cy/3fDdyACAk
4egnDUBQdwYeFyFIleBUuAgtZJxIlDWvCYSTpeltq99RJIkUMt4z+z7bm5JilAAh
q1KeUwloJ9C02o9MMsbcHu6iDR3w8uuPW2zyueNriOvNRIozABHPvcDoSpwIaVSy
3UFqHeDn1won/AighSdMkVnes3HDTQJ5ODXoLlGgodlUD6YL7vcYM5NmjpYFnkjW
Riych4VUF/eoCTKjnRP0gJ+0RjdqxZX74ZZC5PDdfVivG9wblSaAOl2BN1GWtgbI
GHjbPPkKl4uEXDtodM7HdvdMeZSk9AF0i8ldHku0Vo5Ev7aqRCKQ9T3aNWpclnWn
/P7PFoCQr9UXCnv4LkmqHFqjGyXwIJL8JHz72/ozfB6b+nk+vwFUuBCwjrWJRaa3
Rpmkw4l8nwX79YDTu/Q5rsWeYJ0l1ed1b9YKkxZyHVYPKQQfX41GgCEfE41etveJ
3N7HHY8H+BQyuSmvDaCXGZHPHcabskzGmNLFuqmoEA/ZeWd61jcwUa8jeN3TovAR
wjEeift5X/KOk4wRhUHp9fwqJB7pWQCMdWKhzZcyfuauWzbogARRHEIXlbiu61oO
GXkot3E9RNQMcjh5kMGwbQU2NbyPX8K6xdHun/0L75wDDqcCwQ6Hw3wWEnJhVACT
RVokmwWcbHWeR91GC5oVVMbquyu/tQRTckcgjOMeku0e4wk72rTZ2N4pFMWtoaue
gh4GEkUFqGwIn3n2r0OznNe39RqmNV8iM11AmjW+s2D/9s8Y7HG042hbMj9ohQbX
`protect END_PROTECTED
