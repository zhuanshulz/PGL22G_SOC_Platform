`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gXUrtLzL5EbE4qrrPlU11d26t81rymUZhgx8CckT7fTaJUeUt8hCdcuNQu7qfY7
1e/kZLf1rkz875CgquSE5Zgxjh26kPs2mTfEK/wuin+aHJJvGM3QhSf53Ei/d3He
HyT2aRADvwQG30HzlFj3Zw3r3I7jPGyE5SCMeIWyNHSW3Vi0dFBAj4pDdVp57p6o
/n6M/GnhbM4GgTGjQ/RVuJ1nJ8UJo3Ksc4a5DEOXyvZlBCYL4ktkBDXJAnApzYkT
NWjFuCJm0v2as+452WUGlCnDjccTJVmRYM/FXlnHN4Bu+Zx8PEjg2fM5kqUS5PRY
x7O2wHsBfeFePSeKmEy7Pw==
`protect END_PROTECTED
