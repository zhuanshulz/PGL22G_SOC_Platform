library verilog;
use verilog.vl_types.all;
entity V_PLL_E3 is
    generic(
        CLKIN_FREQ      : real    := 5.000000e+001;
        PFDEN_EN        : string  := "FALSE";
        VCOCLK_DIV2     : vl_logic := Hi0;
        DYNAMIC_RATIOI_EN: string  := "FALSE";
        DYNAMIC_RATIOM_EN: string  := "FALSE";
        DYNAMIC_RATIO0_EN: string  := "FALSE";
        DYNAMIC_RATIO1_EN: string  := "FALSE";
        DYNAMIC_RATIO2_EN: string  := "FALSE";
        DYNAMIC_RATIO3_EN: string  := "FALSE";
        DYNAMIC_RATIO4_EN: string  := "FALSE";
        DYNAMIC_RATIOF_EN: string  := "FALSE";
        STATIC_RATIOI   : integer := 1;
        STATIC_RATIOM   : integer := 1;
        STATIC_RATIO0   : integer := 1;
        STATIC_RATIO1   : integer := 1;
        STATIC_RATIO2   : integer := 1;
        STATIC_RATIO3   : integer := 1;
        STATIC_RATIO4   : integer := 1;
        STATIC_RATIOF   : integer := 1;
        DYNAMIC_DUTY0_EN: string  := "FALSE";
        DYNAMIC_DUTY1_EN: string  := "FALSE";
        DYNAMIC_DUTY2_EN: string  := "FALSE";
        DYNAMIC_DUTY3_EN: string  := "FALSE";
        DYNAMIC_DUTY4_EN: string  := "FALSE";
        STATIC_DUTY0    : integer := 2;
        STATIC_DUTY1    : integer := 2;
        STATIC_DUTY2    : integer := 2;
        STATIC_DUTY3    : integer := 2;
        STATIC_DUTY4    : integer := 2;
        STATIC_PHASE0   : integer := 0;
        STATIC_PHASE1   : integer := 0;
        STATIC_PHASE2   : integer := 0;
        STATIC_PHASE3   : integer := 0;
        STATIC_PHASE4   : integer := 0;
        STATIC_PHASEF   : integer := 0;
        STATIC_CPHASE0  : integer := 0;
        STATIC_CPHASE1  : integer := 0;
        STATIC_CPHASE2  : integer := 0;
        STATIC_CPHASE3  : integer := 0;
        STATIC_CPHASE4  : integer := 0;
        STATIC_CPHASEF  : integer := 0;
        CLK_CAS1_EN     : string  := "FALSE";
        CLK_CAS2_EN     : string  := "FALSE";
        CLK_CAS3_EN     : string  := "FALSE";
        CLK_CAS4_EN     : string  := "FALSE";
        CLKOUT5_SEL     : integer := 0;
        CLKIN_BYPASS_EN : string  := "FALSE";
        CLKOUT0_SYN_EN  : string  := "FALSE";
        CLKOUT0_EXT_SYN_EN: string  := "FALSE";
        CLKOUT1_SYN_EN  : string  := "FALSE";
        CLKOUT2_SYN_EN  : string  := "FALSE";
        CLKOUT3_SYN_EN  : string  := "FALSE";
        CLKOUT4_SYN_EN  : string  := "FALSE";
        CLKOUT5_SYN_EN  : string  := "FALSE";
        INTERNAL_FB     : string  := "ENABLE";
        EXTERNAL_FB     : string  := "DISABLE";
        DYNAMIC_LOOP_EN : string  := "FALSE";
        LOOP_MAPPING_EN : string  := "FALSE";
        BANDWIDTH       : string  := "OPTIMIZED"
    );
    port(
        CLKOUT0         : out    vl_logic;
        CLKOUT0_EXT     : out    vl_logic;
        CLKOUT1         : out    vl_logic;
        CLKOUT2         : out    vl_logic;
        CLKOUT3         : out    vl_logic;
        CLKOUT4         : out    vl_logic;
        CLKOUT5         : out    vl_logic;
        CLKSWITCH_FLAG  : out    vl_logic;
        LOCK            : out    vl_logic;
        CLKIN1          : in     vl_logic;
        CLKIN2          : in     vl_logic;
        CLKFB           : in     vl_logic;
        CLKIN_SEL       : in     vl_logic;
        CLKIN_SEL_EN    : in     vl_logic;
        PFDEN           : in     vl_logic;
        ICP_BASE        : in     vl_logic;
        ICP_SEL         : in     vl_logic_vector(3 downto 0);
        LPFRES_SEL      : in     vl_logic_vector(2 downto 0);
        CRIPPLE_SEL     : in     vl_logic;
        PHASE_SEL       : in     vl_logic_vector(2 downto 0);
        PHASE_DIR       : in     vl_logic;
        PHASE_STEP_N    : in     vl_logic;
        LOAD_PHASE      : in     vl_logic;
        RATIOI          : in     vl_logic_vector(9 downto 0);
        RATIOM          : in     vl_logic_vector(6 downto 0);
        RATIO0          : in     vl_logic_vector(9 downto 0);
        RATIO1          : in     vl_logic_vector(9 downto 0);
        RATIO2          : in     vl_logic_vector(9 downto 0);
        RATIO3          : in     vl_logic_vector(9 downto 0);
        RATIO4          : in     vl_logic_vector(9 downto 0);
        RATIOF          : in     vl_logic_vector(9 downto 0);
        DUTY0           : in     vl_logic_vector(9 downto 0);
        DUTY1           : in     vl_logic_vector(9 downto 0);
        DUTY2           : in     vl_logic_vector(9 downto 0);
        DUTY3           : in     vl_logic_vector(9 downto 0);
        DUTY4           : in     vl_logic_vector(9 downto 0);
        CLKOUT0_SYN     : in     vl_logic;
        CLKOUT0_EXT_SYN : in     vl_logic;
        CLKOUT1_SYN     : in     vl_logic;
        CLKOUT2_SYN     : in     vl_logic;
        CLKOUT3_SYN     : in     vl_logic;
        CLKOUT4_SYN     : in     vl_logic;
        CLKOUT5_SYN     : in     vl_logic;
        PLL_PWD         : in     vl_logic;
        RST             : in     vl_logic;
        RSTODIV         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CLKIN_FREQ : constant is 2;
    attribute mti_svvh_generic_type of PFDEN_EN : constant is 1;
    attribute mti_svvh_generic_type of VCOCLK_DIV2 : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIOI_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIOM_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO0_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO1_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO2_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO3_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIO4_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_RATIOF_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_RATIOI : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIOM : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIO4 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_RATIOF : constant is 2;
    attribute mti_svvh_generic_type of DYNAMIC_DUTY0_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_DUTY1_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_DUTY2_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_DUTY3_EN : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_DUTY4_EN : constant is 1;
    attribute mti_svvh_generic_type of STATIC_DUTY0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_DUTY1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_DUTY2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_DUTY3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_DUTY4 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASE4 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_PHASEF : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE0 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE1 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE2 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE3 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASE4 : constant is 2;
    attribute mti_svvh_generic_type of STATIC_CPHASEF : constant is 2;
    attribute mti_svvh_generic_type of CLK_CAS1_EN : constant is 1;
    attribute mti_svvh_generic_type of CLK_CAS2_EN : constant is 1;
    attribute mti_svvh_generic_type of CLK_CAS3_EN : constant is 1;
    attribute mti_svvh_generic_type of CLK_CAS4_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT5_SEL : constant is 2;
    attribute mti_svvh_generic_type of CLKIN_BYPASS_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT0_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT0_EXT_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT1_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT2_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT3_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT4_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT5_SYN_EN : constant is 1;
    attribute mti_svvh_generic_type of INTERNAL_FB : constant is 1;
    attribute mti_svvh_generic_type of EXTERNAL_FB : constant is 1;
    attribute mti_svvh_generic_type of DYNAMIC_LOOP_EN : constant is 1;
    attribute mti_svvh_generic_type of LOOP_MAPPING_EN : constant is 1;
    attribute mti_svvh_generic_type of BANDWIDTH : constant is 1;
end V_PLL_E3;
