`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qTlV7ZzWZWDp6ljRxKmOmu5e0PrzXAqrrXy/RoEmq02JiTEbhyR6Ypc8k6AQdIan
Vf1Zkk8IxKF2WMXEpB8PienHbIyKGFTlz9sgI+CT5kHA1UdZBfIllUioUnp4ql0t
gfCZiR81+omS2Z3JB3B6wl+CdPQ8lwp3oa/S19COSDWuOjSNn1BgQW2BE5+wKDFB
jE22N72GA2KLbJYbxXmnYQH41qJK4sp1zWlUjOVz879tkzbDKNk21+l4vqEyNvSd
/zdOjfJzBhwwQsspNwRml50t0M2pAGoJN+vo3OGEYkKE95I94wNWzS+gAskLPfOw
ldMr9k3fB8rXOMBdQYq6BBhlRbLL2G6a8AmG77GFBHd93BdBiGuJilqLfKXrkoQ8
8rb7i8MIl6G0KFfut/+mks1RNMxtI8XU16tFBVSZl7gvrIyLYJ769P6/MBX+rRmd
EYiVfX26Sy3p3SyX/FlxXNHg8Hyin4IqQ5WQO6n+YB3NqWdXv+UaeuxO9vnBfjd2
HXQQLo5ZTLtrBVotmOZfJSAanOK1aQcJtQp4oiQF2B7uKlvVtasjhX4MqmMtMA1T
WY+7GtlQ+r+WkVCsjxU6E5CrAtZMnCTRuoTLPUI9MiN29ZCjmWVVZgaOWNPY1txL
JGb79QiP0OQG9gmJyyZhLlB3yL1NWBb6ACktP7oRCKESI6QeKJcY3IDatHVEpkw3
oZ+J7IVNLJoodAdw0KUp2E423Pu9HwHhI78VgfkUil49wmjHOM6ZTvD8xVp8vH5j
4V2Tc+qO314BFX3oXQZLkxfmm8/IecZbL6OtUS1UlyOZSa4XCgOBI5XzW7KrRDVl
idh751H7TkA35oCHbH16SNtTLBUueELE+0/Ji40JYPGvIzTW0uS3e4UuorHJEDAM
yEDNEj/HjCrpUxLMZJpoCOpoybG3tc53bwxKWAUfSzc2/Kl0BgHmEIxYsSDf7xH9
ebjlFATANde1T/T15oSn1qeq5Edq3pmiNDiNSynQfbL6CyOjJDOrjuNBidIjdCpA
QfG+JyoOO5uDKOT4HjQpXwtzhbdgrU0+Jn0hCjYegolCX712N3XoW2TyAbvSh9Zh
dWhMZ1UlmwcZXnzSjSm7a9sMfw3SkYpqmUI/lNjcdLCkMUMVIVqy5lRepsxmV17Z
Yggw2fx52ODR5oz3XZ/aRHzNyfUzNQXegis2bVNvr7z+SqFLr240nyDt8AwPlGDf
90YFXHeVWXEFkn8/6R5pIDeCk+vuynX3rgvnuugv6Ckzb49TMK+iz+k3qzDS48Qa
MXxNl4kY2rgxO47kilV9u9IuQtNRmzxshuuSpjGBb0Olfscme73yJW9vsqmL/FzJ
uwnJIKvbXvMXqFQRKipyD3CzpIcpNHxVcIVUKrXnIaNliyAX2PSQRuiz1jHMphCS
upbIpbZ3+WaFpknBC0QXYhMpxZlBvU49EcGayZwrMUagp5ULR/S+sZSDMPUld+As
M95wZ1ExX6RK8TW2quilH1AAoRzre5S5peKudFQOAXg1IutGu/ZiY8LELK45HjlL
qG2Z+juTmXyUVSJYL6hicgu6GjOqS8SNGoj07+bn+MGIdyOWWy+/hDzQfEqZpCjx
3PJJ9df0sl9yu8yxdw1RBlna3/mQIUYLqIfP4aGPBmM+9pCUtntjsDJbU5FMMi2l
LGfcpevgn8Gtnuz7rQltBLbaG3KMJzqrVnWba1xGH05yoS1ea+TcVXnEWKeAVPVB
NTWYomkUTp6/w6/ECWoWApfXmSlobzQwZ6KlPgP8FLU4vv9pBU49ayn3pVDgJc2f
SQ20E/hX0vCD3MJFWsuDfzJUJFWHqEKl3kGtOLHkaTpRYZpUWhhS5uuK6lfprasN
mxo/NwpQaJrBBf9sgVMU5zKrqHsi6E9U734p6TxcGbKYjtiiKGvqtgnBbPswF76y
wmSa/Us83FcxJHBENMO0aev/G7gDrzzNGAAsBhpSU9LomzRVPZCgfRH0Vmx9jDVe
iFIu4mutrSRTf4D4a6TI6DUZ6EKJs5ZXGQvxgBo2cX4p6m/SKHi2EQcDI0vUYSZJ
bvgi1x7aUyBe5J6Qzpz/3QybMB4Sbd6TIcHUcD6GAE+A9MJJY/V+WM5gXFEVGw+E
8lHxjfcv19CoGoe55HN6dat2zMEuZNDdf+G3olumQ5Y=
`protect END_PROTECTED
