`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkl1igfgPkswK7QctIBLNXL7Wgt1tdlyS0ZBlUOD1g/jR9fQ8Bnz0BrTDhxYhu6w
veWVG8AR1dxv0drHLWlepgZBTGlg3asEXGDvriqYuNsHZaNbt11SpkH+WxcjfGrq
oPN9X6dfRAzr9AMd9JUZ+J0y1AbbS8E8JOWKJiLm3u4p5kTB6lF73TAOV9ha1g1h
2YMterJLsSOyMTTUvwFSA7VJAWo14Jziy7x2fgFuZCRc4c1rm1n/CxLMiOjP/sIO
a7lkBrI2HbPBEiSlRF5sTDr+E4a15R4kGlfP1Ap5UDsaic4iZWWy6qnBkry8YRya
LONT7ye1NLLxGPpyEVDZNK8Bc6zFoTOhv9UKnp0ul44crkFtYyAOwOqWGqVWiHAh
XSNA/wzorajOdSM/PETGPPwWTEuh87H3hxndxWSvTzrxyC3PBuQgnJ0MhYSKbrua
lc84zgiPvjXG9Htuj8ZzkOM2zSmaNv+pssgZZ16BUwEvQKrnRNca3uRf7XVcsDmC
9t2BgI+bw0CaRm6OOvIr5xZltEVE9yCvMdIUQVuL4XEiQHCYMAyWqw8WfinubTwY
Yq0tQ2v9ySoQWNpjtx92ZQtdJxBdDzzzfgi0vacSLio3zk9zDEpsMQBL47/0WufD
4t5p0AUzfhH7KoM3lSx5jnL69iE/6Gl10hxWx1Xf52P01hNgjesxuSioFADQ2Ja9
vT+HwZc88yguzkRgUx6iCwZEdWhg2XAo9OFTVJZ3W0lpQ3xzg2O3eAJs1T9yJGPK
hGXAtas8GVP32TBCcP1oLo3aA2/vUiVBcBjrewreIZg0jmsnm6MgVArkmbDX3lsq
ajJusYA7DQ+JtuVKD1NzwcXwoT3Ssh4+Tj2HkkUJmyv8rGj5uYCYqiAiO/vLyqcO
PHDEmc4MKF2w60V1LaHNfHDZElA0XvjK8RjiLqrncufuvecWCdKPpHuDcPS4mDkL
6t7pViy/nXFKvTlQfWDAuGPGy0RkpRcF9LVyisQtHPOkaKAxOKX1++vlJkA/aC3R
K2OZWnvpx9G/7sC3wzPHbmDxBgbSl6H0lKV0nYsDW59AsdHy8i8TTioKeb9Q2e82
KIuhiMT2uQKAR3t1ffNinZ2C94LTKdkfNcVMY1GEeo/ZXjx1YYlDu3Wc/YyjLeeU
DAn2laYWLl+T6Knx3yFAIetYZinYDB0VoP2TCSpMOzjliv0fzlcZwSbcU/loHFTG
EOEOS6yoKhKCoe1IYC8I76vrkWhiC/CJoNCzJy7iFiXqoVshaXmSGbH95KZZx4s7
+pdZRdMximmokPiUqxNth7kx8DqHF6EL0vMVGy/SZlp5rGJg3ckAL/IvMZ6mMEwo
gLEkCLL542TvodLjg8qAuZKigbEw7Uh+9FU1QN0105twQqW4WCNYzGjlhLZ/86Q2
`protect END_PROTECTED
