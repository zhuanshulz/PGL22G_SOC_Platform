`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4u+hgtfeniS9GuvKu2z+M5Fea7JMaAvvetyF7z0nD29kOnPXlMNeJVoy5UJJCexK
B8BhA0GZIWybrianr9QTjxg7XgHmjKmX+84pP4F3sLtcGcuVnUVR2YPCnBwIDiD0
bJC/GFnJqDw7nuagBTaPbqp05m7KWwla2zU5tHxVLjCgSemlx7p8nLYw+vo+Cz17
r47YqfDqSKDYiMDm/viK5Qx0SV0Uzq2w1vaBThCxc0f9AioLlXrUK9z/Yeuy6XLs
wrAGP9Foti0hEHk6D/3M7wrc6kuCJb1N3QfEd3N+G2K+j+nXX/0+vDli3Hc5CkMW
/P+pOveDJ7OVEsbBMbnkOh1b6biuFgwwHeF9nxOsyEgUIMELF8edDHAQD/TlrAJq
OOxVFLCwpb7KRrQuo6wNk2tEha6gt7E9MCBJBikiQuglsmNoe9fEcyK4dc0/+5st
87m80AEvt32EPCB+CgM62y2fJT+O0k4l/L/eo6QcqLzoWQAT2Hu3bdqOG/NhDdFj
IGAWTCwRnF6iUU09NjsLz68pgRfBYlmei5lvYWcx+NUUmEOKDjgiPxk/o6P5vWNW
LGwu0shMBUFiDYxaeOb1UPf3XwlxjaLRU99sUQfLDV1jW9S2G97guy0cSp7plc3D
HdlDOWz8aqf+H8qqpGvdaZ6FAyhvonl/EpPbZKqKmBENBpRJVuM6FxpiUFox7Cj4
N4buu2Ib0kvbIbbLasjpIwOqrH0tX5Fv10lUZ6FKLuY+GNaUOoZ81osrUVlC/lmB
uyFePpD4ms8veg78koY2NpbUYczNPW/kLOICeIJne1lJDMW5IksKMEn1Vym8aoKj
qdyLJytgpbtr38+WeMyOndd/eulA1EZeoKlVfQRCtHLC9QuHH44zravblHdxTf5G
x3YFFtS6b2Mi1t6ib6b2kVc9HlJ7Ypl00bKPSfJWHUHDdY2Pcp33SeWhpUi4LOFR
pzHgRp09HmAnChpPfABpn7TwUFbNEDO6CY1YFIM4xFmzHUep8/vhY6wa5ScZ1SwG
BBSp06PrKxFGLniw1V/mA/E5gVOZb1I4PKv8cojdyhonWoiCCww+gaTF1yxZ1jjN
4YBNDy+TZorlRIT2LtO8GG+jmYZjxv1P0xY9yPZZaC05lvxEYtWHg+CmPVXcNOl7
Dv3Cb+aUbgf15f89HACxbZo4MrVCqnmHyR3sCzyE1a3Y63TSn2Q/G1I7/Z3wveXF
4uT1mfB1Bb35fDA0vG4xsC6yZCXUFv3t3Cz0K0t/RfIwPD7XvvNQBWZ7UOGZTnTt
HoET7VXkF4gZZK0HiQJsVtcmv+tb5XBWjURz9t7CLFH5nr9uB/m7fTHexwZytuvm
tIsWvmvKKM1SRyhIM1mdWNf8ZwDKhdk909bVNzLDvzFMSE7wx63IO3e88jH09Z0y
I8/noM51ZJ3h4ba7sHfMdzExgg01aXr7taDrzlO+/z0DNiNGAHADCZSXYHQUPGXj
uZQUravz+t/FYk7ABtDt44WPMDjME3vrx9/rYxJqnHF1R7HckPHd0MXrRPecGjkk
p018gJHmSlw4ie/ezqRxLXeFrV7BuYlBE1FpneSLc+9VzOx6ij665ufYf5QcXn7N
Qf3hpQH6rrGnke+IDY99lY0tGN0Bl0qWhyuqpFaAPPQu0EgbP3f92+oJWRWn1G/D
l3nh1l3KejjDa68zpg7bG8J7lMkQ1F5YQSXE6DW1Lw8OUovjObW7gxX5dspC5zer
/oQUveaOMgXjaIx24SMSr4cYLTzghdnPGg3KHRyOtPG56wDIoFGxrbB79DG91/4l
NAPom+RveBrk41sL/ZTF33Vu2XixfcI6DSVDcxnIeqJ83fqgD/3jW9LlYHcNCwta
RUTODUHvgNFfL43SudliWtS0OJ1UHsYG9BaX3kZOaLlelkys7xCaeeyLtYNqaSIh
ILZ0Nmq4ze5vjAr9W7YY9ssGO78U8h6LHCg5VpkV/DQ+JAJNrn7e3WhLV6FxHj7Y
0ec7JcyZF9pG2ikmriUXad+vc0WJc17RK3w6PGPJQuZb6azfxDQbpkEzbPz5G3kL
dj7Od45rO6X93n5O9h5fB2y70ru/LkUBbPpHZSnZxBVSoZ+5rkbs95y6281lq41v
Z6KCRUW4AvHBmKDFNqe9/55mj1ScCLHgvQdcfMmN/F0TqFIHbCX4Ozv98Aij7Vte
aIhajGEbzvh4CMucoXAWKdNNCjyiR9po3urtHU1IoFUamLCjLHVwuVekI8O/tPea
IglAcNpXCPgt2RIdWddkxVjejX6OqUu+IxKiK6XwZg7c+9w1ke2iTjczzmSBtXoC
Q/T8AHT5bFnHOL4yZgXCZ9dMo0A0NiL9xUR7QV8DsoWsDn5oUEF1cTYr4htub3fD
HraOyc4h3Rheg9rszl1jYok4p6PYPIxBaQRaIKJgZQ5I0PphnMMnwK54s+r2d894
hubT6P+C0kPHU1rM3KbB4UD7yu48Okb9VsLT9ezWO9pp8tSmBKq4CbPHB6xgIwMs
dHeyVmZuBnb5sUFis7GpgZFb4zPT2QZWhEMNrVvPgYVV4elUA3GCJ65WpUi4VjCe
TOulVA0rzQohB6fJh0OXwr7MjMfhrPEV9iW59Dkh71WutFEBcF34DJt7a158O9QD
E8huWeKFlx3dPV4UjGs3MpqtbbvWfVPmJJjVJq3WBVLKyj2qIuzuQy/sCtmmotYc
rquwC+YHrCp9j3amClP+nrTxZmLsjd24g4neFSRLFJhnA7tTZ3u/yhZyX/p8/vgz
7Vwi2OGzmYKkInNjvr4WhfpqKNAr3/72rvpszCxB+vz9vKoxwCVlR7+QUUcQkqUZ
G/kxNAgSqGOVlcw3nv2N9C7RVjV1f0CbrZ09FyZ3yzTnVORtFunsze4135wQtAcS
FS1cuWXjavUFid1YcwwbVNJWlijvTRmgB2Cap4p8JzocX6NVSF9s7Y6izLH0B2OD
V1fUxTodmzjX5LdzyU9xh8LTVo+GP0mM3qvavDc8PH4zu6oLlWT0zDU30uq1SYIv
QNOBx/3cyyyuW+/iitxgBOs7NbrDNGDZmy4AYjruOQLmIgwbY/yx8SXN1+D5lnZp
I7NHQs3vcJSC7fdeYJgPJDYDlZBkOPWN8c1hcKNskWGSgZ1TKLWtBmZwlnwp08k4
KDkPeQGfAof5WXoCFmZB3xRFukIJxwDP+LKja6cLb8BrKVp85JuH90JNsasEdLoa
tTPXe+xz6W+2ZeDhj5B/+tUaRjIfCpKX4/XIU/7W9nesTIG6m4JoMm4ajUuUjPq5
kgJ+tBMz7sFqSRxT8Gg21xvavOPl+EHvJDyPq8LXGsbpYsbjbZFUmQfWyzcGq3H/
1If/qKLnTMC5M/g4v5p0vjVxMbxBEtC62WJLB0l6MAzHLWlqIjPnKF89iRymbxnx
XDqeDxC7YDz/fghvJGZwxEjLchbknTFMnlsFGZvwnbd6jrvA9qVtIRkiwc8Yp88r
mfryWXvAzwomZSb2OiiimPFZR9Kb5IVmbUzk9E9PFVd02tHK+iCZNCPBvgljmxBZ
CJWuJexVH/UjlxyTjEUMMzuVdYfGW9TyEz6nFCShcgJ4gOxdYBLWAjHEtO+U75nX
6HqXuP+yGJoW/lnKnvBumHAe1JZt1W2HI/gc7/fTukKzdtZQp3CbnJpvdNNN5+tx
WJWbQOG2QYRW/Sj2utIR9xQwgS2exylDAcIAN0eDa3x6bUCHBsCrZXpA3Q+MszRu
09umqNzQjSiDnQ+2Oy1y8mp+8BOJzDrif5qJUlxYyuXvk/beIQ1OCrKqYpW5QJ3F
myH/pxu0fgelxVk704T2rydsVCUvO5W+ID8kRR+nQ/yPlHNdZXO+eezajI4mCcq8
tRZryyfBhB+4Nzr6Z0sqTAKQKjqxFzJ+WBDe1JobObfQSREWzW7m5trNjOhd+9K2
eeG9xgrKt73cVXcQ91fsrX+rFA5HIfAIfxbhn1jzHvnn3QbGbRgvqp/aRWU7oHKo
vRLgldOBY/PKN/4OG7WP/tV9nXgd8hep4XGM/A77t6aJexDPFM2QfSu4kvSiZWuD
W2/wGFbIvFEf2ixpRebqCKwxfny9Z/EKFNXOR9q3IhyIUgSVsdPAjQ9ysEgQjQFm
Om/HHM2HaE2d2kjy9JsCRJqEDHpo/RdvcqQiKEAUi09Ajs8ZkNptfEv/J6Gj+X4b
J+2ogUCNoijS2ecbJAKDk+cd+9Fu1koy4il9cvB13yYPII/U4AOXxmjMj5Bf7Bai
86QA8vdqZXExoROUOt2VYY/MQFq3skUnrX6+sdA7L5SUgZzS3yHy5ejqheVvh/Fc
Pe9X2p2//MpJTr/zTyGkAyXA7DhQry8OUpzTRGzy9hJerzS5k9mcPd9N/U9xYuuv
n25mxx4WRgtL6xR6hyphkJz0RBfGDtVeRnBZM+oEDrmW/fqAS91M938FW446DIML
tayHXTQzULgVAVaJBYwqoXunWwFpviFJ7Hfh3sfmjlrtk+jY34AKgrkeNLoz9R3b
enTJPuvRmsri0r5hll3/jC5UKxFiV7sU29/vtlkQHpF9/s9ZJGtZHFI+QZQqX80a
hrO0NQjKIA74AIMqzSWCfOqAZVafM+f+CJFXanHqLABxPx7LeICoT0ZPM3j1O1zg
wjQsxRQAL9V7r9DRFAdoXCvBYIWv1bJR1vGcQ63Xn9f8BUoczY6E5w6r5I5J1pzr
xA83Vdsnzk9ixkgg/wkYly4t0RJh262PrZqs4JfGqTSYjF6Gn48gaAUwzYeOG37n
7Iry4vrVp3ZQFKr+AUUa6dEvJFIiOoIhfsLMBgOq+jicn8LBpmkvYBSMrFxtt8CI
B44libZgXAiZnZ11ZtRilafV+u2jyZbcMMboMGKrN7cmgUTY8MVuVRFQRVoCQQOV
2UwZeoUP4hU+PaOGZQLT6d5szSeToX2/x7zH0q+iWbHtYfxti3hmCScgQBydhwEU
dfJaCoKsuofDzeltOm8Kn5sy6pDXJsOgbUCzJ3pYyKqoehNWJh+3M98dnSaUkpxu
A4nCgZH+agnF5ViLAGcv+FbeFiOvuAPXkp13gzCzpjoi8Tl6btDRF38skTCw0rUu
8jRC4q0IEWG/OtWkUbHMvMaBaUUtdb2qMIv7RZtGuuAg3whxf15LAIunjYWVASfh
B+m+79bd27bNsh9QBK6aO1S+kZwiwEWjK1PYaL4GUU2mttIgE5tfN7IKvr7a2bAl
JN998y4SJwPY0nGID3KzhnktWt2QTjlfHEQEVk3vBoE71rdTegTUo4OL9XXxDcVk
LeXTQanjg8ycCEoH7dHAYDfMOmzDtMsLLy68+3ehzADqFtu7Y9l2iwQET/+8TRfS
HUKxkopdHDuAlGRurZHR0QyOwzM5R+H9jk2yoTkpv87AFXYnA1VvvmMNVDHeA3Zd
Mptb3sK3fTmEDRjEu/8jTrOD1cH8KOmjyGYE+K5gTGr/bSV1x1ADBUxnTfGw70FY
PuHgQB+up5oWAcp7BUiEAmPXJR0KSF/RLCTuN0kNTVga50PMBeu6LdoUybfoa9/w
jsNgjnu2t7A6sYWHEAmT0ZbUE411KjgYZj3ytK677JRT4peQQRuMYLvl/CEF7WV8
v+dFLJZozbjSrWv963XFUQs8+6R3XjeJK4tgprIhN4eqneo3YWvvbUs84E6jb0sd
KykkJks/PsjGMFGksk6m8chqcsUmhjoRyYm3wQ/1440iR0ZoZP4Zvg/G1Zlsgn9Q
DirMTS+OImw+H0Je80+VjIeyMi+TzJG90WPtWJsQIrtEnc/8PNGggP5rmy9n3wlV
dU/uo2sVu5fq/cAMSJSJ1pczpEWmMucI6W0vsdmruViDz/anZ2Qp/Hki2QJW3Koh
/BziJH4r5pyP1M9CtiQwi0QtZei0zhHSZ3KOkcKd63LF8VLH2kAUav2US9ja16K1
R6GvQ8A+QdMozyjQBmLqKGm9XuG9qu/CqRqitKBx9r9GP2UnMlmer5MVOFs99ksv
DItt59WGeJ6ncybecgPcYuHVTntIiAm2b+dLxmcqUH+8V0fks9miiAJ8WEvncpSw
I2BQ8SjR5vcMIR4LoEmqRRXmCyCGYwWkwdwOYkvszvOHouOvctGBjs7XRGPj1RGI
/RkvzfNto8/uq5FgpDJLYse6Bj0j6hz5UDKlMiWvkZtOfFwSAld+RSuhjAkdVHRL
Ww2knHOz9JM2Y3FQQzog1DJ5v1VZ8Hk8IhthyprMthrytwhf41sP373Y6ZGQyOm/
CtW3DvfJRuQuT9GphgCDHnxySCIjumksr9Gt7JOlNR0hm+Marhk+dX038hmqlZtQ
C71oTQqDnguVyICvc6JOmRKaHHirYzYTGW8Up65hXj69GKe+HO3V9N/maDMJES4K
rQmJAo1aKOY8hKDsEeTfHr9KdLrk7f7mDsXk+tUCufYBoemQTrzECUOCxEAy0Eaa
KWmFATf0W1X3PL4VOYkDvuzPifthQVtNxinb8+Z+IBtirgMymp5lU2YMvz6JnXMY
nc3lVPcYb2nLWCc5AgRBWyxkwvFbPWGOwApPEdYS/u6qySBqx4qxZsxcuvOCsWfk
vcySFs8Apxxrjdu2PiwktJH88TSkvRg3YWwus6hHZ5zOywVrcFRNXshkZzsx9/fL
joJ21/X6v5jIrYXYffIUjGe9nADgmTh3Il4tZSR8VKl/is1aduLxzOtackTSofq4
raxP2ou5QbfXgQYTNU+TzSIP+i3rzHKsh2J/VBQX/p2NlfcoVV+Os8KwkwDdW0hl
esNtpFYhEvvw9U7O7tFEIH4PPAhxb5LPKd/YFJ622TEVcjcD64MlQgzjj6XPj1iF
OKnQl9el6MT1OHmKTVR5EW62KxJJQV6LLA5ZATOUILRC14Rn2ninvQ0c8psP3e5/
KpX9E+Fi8j0ATByNpn+4e/QfSK7xvNPx0Ynoj1f/zW5Kk1mWnjWkBrZb9jQn4rq/
qM8bsZYx2kEbzXl04h/92dGn4WbOeCj8JDpFKn1SVBk7Btpcl37yQQhkYqQrSG+J
P9wIRcfu0+8nVwixisnjS9XEpANFHBDKnNdZQks/dmIF7wldnVcwzNWigeoEkomG
SfQ3WFsrd2cUOJ1TLeL20BWDmpMDcfcUUNGlOHd2cTBVedtp7hR7YOI2MDEDAbWa
t9cu8Ejy6m8QRynbN0U8DvQNUB8B0UC+3mw7XE46CmQq0jozhRhyZwX7Ak1J2QoQ
grNh1dGqGL1vALwKiG0AcCe6BAabMmvcWgU+H9KaTFOEMj4ohh1tFNjS1rAgGUDO
yrkX+LMdmIO1ljK/ckH+PL1NH90edB0O0+CZkKjTCLzXNQgImiAHD+Sleuq9TkvW
nbD54LDdaRwASBQ7+Q6hlWMLA9+5OKAbbH0tqSeynJJ5jSpWdC21VGdIjCrIMhO5
mu5GHK+lmTCPFij58eqrDyJmf3xBtciUI4XteG6kdbN/hcguaReMQ5/1sx2Qn6pc
imCZ9hPz63uHFu45VQDvYe40XBZDpemDyZYQVQm6vZyKe+bdPX2bK5/ctmPAyKcB
5OETohYObfmtmg6gi4wOq5/ktNlnkhdo1ACNmodPvVf622/JbpUKljKma3xooj5Z
h+am1oE4fffXicCpy9EaPe2w5extksrZMwQVDhkKXLledA6DoaOR/B57quf9dspW
7tRXgKkwG5PiqX3wU2ysR5MdVrWFy4jjrmKTUw/f8fI/iAp1/UYBWfm56uXT37Mu
qp89hI4v+Xxr/r0WckJrFtFmnW75aem3OxHOEN4AzOKo+nDnI3lBwDaDf5hJYASa
KalV19PFltSO6ZdxhBn846UU6jPdgcyicTF+3OGgMrK9ts/n7mHpRFpgDHv9vQvm
AK4OE8kmHUcDMEN+5y0mHcxh6u80NTMd9ZqNf3Hm9DrY0T143l4gPBRf+9xRlCu3
xphW0PnXDP/frHgyDOODoejFjvUbBhOXDxtftAZ24sSm6gj3LDToXEu8p7xoKHn5
1CMSD/SOqNKI8mcHOH3E9jc+E1CygeqeSsCDFD3DTsTtetB1hYd+biRTrL5GjSy2
FvS/5kLFWG7NOatSYbJ2Sc0ehbMJMfsmHhqm2wP1aVoxN5oVRt9dLu6bLAUlyjKa
XJa6kQVEhnNY2vMnBanMxy/7CxhVDvE64+ipL40V7nn6quNPEAncSeaMemOiWwNs
ScVJnX6ypc+iq1wR/09zPzRfDBxsA5wep611Q1JU7IFtKtY00DCHZx5LwmFvWOu1
NvZJmqrcg6SWVuPymPE/sFs8VEFCS0gT8PxvDjFc5Sspy9mGjIZt9tkTn0Q+UBtq
CnNSE1vSGNJZNWVOczAn2PJL6xgCt9KWvi3fSLqxKxhAq7+jkeuQfO+7rHR7AyTF
qLCGxSv1TRMiVehYlSG7DexEcJmIYdWBd/df8yx4qxCiZLNzHmqquDSNG4S6L0ag
ra+GhOIQakvjpmWQu4ta7sZRHoXKMZ4ZrqjptsLWJsq2qWFTjly/K4ftoHujKII2
z0G6xu1EExDHsLJ1TmVF8K6izrYagcNL7Dgi4hEvdHC+xTLgceB0lWA07cyjFKZ/
nhy66Gbx56W45SE9yL3eA+pfE3bB/28KWvZXDxy31YpQvB8GLan3BYrxWQic5nlx
ZnrPyxHC2RsQPP0KLGf6DheEu+RA6+GbGIYcTi6t09BCRGT9E1mVHStKlE15417y
`protect END_PROTECTED
