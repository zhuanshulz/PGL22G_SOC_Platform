`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wabod+DToxwaZn0dPA14keB7Zx00cuzWULho6hMKVKP7IHIR+3tg2QY2/mTOjVRa
fSuGi9c4eLziBGxuQ0SoJVtG1SYZIpNxNL+Io3JJ74FOGR8CLPOwsloRuC1MiPIB
DvlSf29rRBQ4HSEx4HcEF9Z2ROnx0of4tOPbdDCBEMovBrEdzbc6gCbzsWysCSdy
j/v5DGkD1rgZgL8FRNjlq1lwKananM9cVtfwwighQtxk7l2aR/c/BAHi3znNONdM
77p4Y9OhQXpdIVcXssvrMr0SekOxui1WrAHRGENQUbYF8yI/JE9iOVauH8CRlwuR
5IMQz7yhDT9/DfLiOeFXQc2JUUGzmIN5/tkLND8RnGue0cqxYr8+jdTVkKGeKNHD
4WQyTqa3o4Jpv2gJcMkB8G91xEbxl8q7uodBPSZD8y7qX9QqtmiywSm2e3oXPdXy
cGZ/bXEkAFQI9SaH10hypIcNIBWzygtRlDPfDQ3HLfH1BjGyh0WiG61rt9Re9y7c
+qXuo2SP7vsrvhGCiIFdaA==
`protect END_PROTECTED
