`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e5/X07aCFSkl9lPuhHHfhEKTe6zEYgi9lLBl7NxjRwPtueKb5YSjDBDAwRcqyANA
msj+OBrIJ2+HYd60jpqJ6RdLotZNWL8rJSva7jdSKtNeIKALXoDlIqlMeYgoPoVK
rOhSt1x96Mgr0rH4STQOol/EZwqk3lQ0ez3g8G0ht0lDZ/WuqFFxMnk/3gGodrw9
NfNdGj49OgJ4sHptTp5a1BpyA+/dibWWnZJzyvqGtwMMEM7sWBm1VdBwiqKT+7TV
+4XUi/R6CoF2gk9f09EAWlARVFtGtsy6KEggopBMA/RcEIO9gMByGsIiNn/7gYsT
Dd6phJMb6mF6VPEoHYIKGn/1Tdv6w0ODPDQkHnzuaovn/BR3ywN075PAJoqyEpiN
VLPwfqdoP3E/IVvoIkBI/aw0uNqyYGTnQkxD1ifuotcr+oAG2ITq7juG9N89uX+J
+ryl5HHFiZc2xZNyCyUhjD8J9NbCgHLpS2dgvrSA1+iFrEsgq5vkNG1o/a3ocdEZ
y2Yc+lTWOkB2nm9Ife0ukBBYVAGsSfHtGB66inSF0MkfxxrtZtp2gCjXri42Ktv8
kMSrt+tOP3zyVcEchcRX6og8s9YO3dqUSVZ/VOlrEysugo3iFJkvCQbTB3le/8mR
UisXZTsktjDoCLltm3InEixwjVf8gS1PT+smzpfIhanvGIMp/jvWNhzRqoFqaZlu
pk0fv8YUDlMRUba7tFnIL8XdY4T8Nqw95PHi/5C9G230xZyL075wE++r3f+7Xn1H
E1icUykCaiwxsWfNAivRm8nBNsvftvi36/bTIzPPFPTuVU/cp4DwEo/kByExHyo4
c2VykoI9AH/8CELr+YTmfw3kBU53ZaAmDrNWpwhRKCWyJqyRsfwvmByKXZ9wUnLj
6XRPjK2Q9JtVOuF9/e9jT4eLIratw5JD3f8tQjQB9BX7tYXxyVldwHbxTVr5aWRm
Elxp6reBR9JI8LnFCsUSP6Eqp3aId/Bt4qwfDFMJRdnhcpYtV3L8R+JAcX6j3U34
Wwk9LieaeR4mehdU/HWcTWG/erT6woLs6L6duGp0Kx0No95Jc7LTHs9M23+dGDCT
SoLKwEyS/aeQAHnimECxJIhyMyJO/L3LS0/yvJ2tEhg9VDgisJZTtOEHNiNPgx93
1KEYwT9kgoVJpvSmkzyOjAhlB7X2N5dAMSYTki4XPCdRZuPM8aGJ/DvuY0DQiWov
v2PbUY/sw2uXXtDWv53N1Y9LSzDo208A01vPJhdbMj9CyWNtmIom2fYD7U2rKf19
cfe1Gx21vtWENZgNdK0S5sEgT1oJ79/i9PbvXmq77ftMZuTBVrKLBMJnZ+rDnmBI
uD8o6AWZDSTsFB9fX1uT1tf+9RaJWLjnfdxRa1KYpNqduV8dYbwuMaec879X8jam
cM1A7zahCaReAOEi1zrq//aZuAT61DDh9DbXBZ/DcyH/+ZjV05KLU7P/y/dsuJD/
4rU6UvdGniT0iISmeybFJE9yamhdJhpcuJYjjsnVAnfvtb8K0bjbw3HEO5FDCmQv
uHnvhTYKjpGbh+UNhxJ1XUtJhzOhftUYRCKq8M4YTM4DNEUsghQM+M+MkcKmd95Z
PThjPKmBl0FsMvbN5imaSfQzE72uYXEWLszXaZft0nzmoBZ2ni48EEa+iQaGo9/E
xanH4SDP3hQUKZdX+B0pDduD/T7WAduJ+AAr7vDY5F417sEI0valKNdE3SNOgWjk
bSsnRV45ZOMPHp/nISrN2saj1fC3ZZ6XLTR5nHi2Iq5vYCDhjAsFkczc9rlEdh7v
yBhxqn3EiNj9PYmOWmz9qCTC431/LJDNnHhI+EgdHU+/XUIyM7ucmfR5DCxMqAzK
iihOkmDOfJZgS1CE/ubpjTpNRVDhB/Klv2EQxGEpWApz/WeGx1pH3Yvup93Dxo+g
HmHHgNUIYfZ3ygE30yMPiEyX7IwEV3x30/XPxlgEG9q7/0uSYqDkp3ocfjt+q+sS
5lIsYovgCMb+xMQ+3N8Eeotp9wAavMYypOdoW0RZFLyuQnmXsgcIdlZS9RZ5Fpl2
k2WdyjsgPd6aaZho+TXDpa7qxd8b/ZgCZnwE1jkF6kYXaJ4az4bxYyhI2uvwzX33
nEZIb7HUgipOqNhrmgLIh0LoG9D5bSOmnrpH0dM3gq+1kTc//pMwOf28eCvKQGXd
GQLBr9S1hasE4DRpRe9PprgxLcOUG5d4KOENRVJ72xSV0dcEqGFUssrVQVerz3lc
/d5kK+Y3LoiTznoBsuSmbsZphK8823Vi7nz7uqj/pwwS4Mv4WfygS9wfcYwfezdF
AHBrb7afjhE9iMqnrQcGtgKyYI2oQvgfajI0rB5Ye4dtSTBn7PE8fwzjplvIZad7
G2Edr/gfpn8SzxIaWb3KZ/3HhSl56GZJbOFBSF2STzXZcR1LZCmkJJxBEYfs1xz8
BJwyqpZzBmu/eWANigEzDzxwRa++m5ws4uLUNSLVwUIwWqdD0muydNJ5hBBVgtJT
Uzj8zxWYTk25NF/YtDZuBq44xdZcjd14AgVP2QJ+ZHTG/bUKLeJbnDK1IyG+lM4L
Vuz+yMhfnRSgKUBNlm/AfYCw3NasT34E64/17O3ON+FqTsCmX2n32HXcojUVvFPo
JXDnRU2C/Pgpap7VKkEob8hIusJeptjfsj/Owsu1B9zcv2kTKLHBWw/hClGNnHIX
FutPj6SYtH+bqmlVHs09qofQubzYxkVZGX/q+nWuu98akpdJ2u6q81cJX9wu6CC2
NT3/XTtGMGKeZIUOolCyHNSFKNHEdFasml7/qAkvYxFrBV9zmaxqhLZO/j9eZrO0
lTVHx8OSAxrqVcL5Ug6rXEv1klLf+iWbiFC+PKcQaici7Hkd/IF7iUkC08eiPw1g
PK7IBreKOywEmA7Ybu09fyNjWld6rcHOpvzappa6XrxZOw4UVWjU6oa/5MTvB3F7
XyVsc2A/dyFwmO0Q5vxIT5kAvgCWSMWG7+PZK0l3yfoxtPPCvRyP7vhU6f414b2q
8HAAjXk+QQdyiDwy/+QGkJTreKGMNLIaFOy8B6r89rgAbzkneYuorkGt9JnJymEe
VGII+dVVh9rD/ytjtHdso/IIF5ykWOumf1yfijD85mWUwSH1FqCc49F6TXQrzHPX
j7M5RCfIfAYPahVSe+LepZzRSVnJrKjrZcKaAzJ2/bSX1xCLWl7XPDeSwxK5mUdE
1yAjHcNK1WjfDe7fe1NlKupUywsnb1IxeoBM2nLH268YST9ZhxmHWo0HgBTinZBt
XnpSUxafMMhMgBrbJNG69trXZb0U2uh5s11onw/9Ws9miR/6EeEY+XvAi07eo+1G
ysQewyHR8LO51miNbXHNtRYMoSSsQasgqcl8KF4RXY2UzumNrzf2l3lf8hPYcgfD
ll1FmcNnPnWl3fz5nBKtn+exCCYWy2evAsW8xhWGzrh2REX5L+vHWq9M0ooAEj2d
wkTCUrhTDNfGfs62sdXewPK+cjaDLlmCWi/9avY2b3pfy8H0OVupj3m/KvzG8m/G
Eu1zobu9bibcqSjob2BSmdEeYpwFfaZv5Xh8q2OWqGfZudRJAMaMP3nbIihrBXdg
iSXQD3M4YOeJYiAIxhTqKLNOJ1xUzq3WgU1lrDETCi/RXVqH5jGdhPTgBSFV55pw
XUXFXyl0mHNrj6ICMcpa5xDx6XH3cQJvB84gATbg6VecVnNj17mgbEoUCF2gTCn0
H6y0k9Dv18IVq/7q8UDKhM3983zJKxHZZ/BwoV9X1h9Tv6dxfZJwkwDPmasXaABm
D25UO2Ff/m0GOfvRI4iLN04qBb9Ea5M4dlmTtkty1sqvQnZauBB4bDf3ia+cLxLr
m6RVkAYXXbh9HtW9gGsHc4ZSqsqd5W1HSbnY1d/ykaUPX55NSiMNASgRJ8rNvRBN
7BnCHDwQKzxd6nEe2sgIV3AmnPWUVe3g4+Wq6z2WDZWlIDZX6eFXrJ32gGLRKPBG
iwHDJoQgpTm6fkrd16432ThDt/bmSEF1MBBCuMthph/z4f8W/rERiIMyc6VS/WDG
cquNlL/vrIrJe5bW9EiKIZIUOOLk68ItoP+fl0AyhiqmS3V5OEQNJe8umJGeMNJO
0q+fUvekRkh0ASlPdV8BoPmvWwZramO/WhFtoDzvAGKacGqCE4KLqWggRPt9ivIV
PgMZokIpbHKVN2p5qLMZsWhbwKTdXk3ZTa95v4OxF/DpYuOdYCk9OE3/eb8/FMPr
YIIhKWn4pSKDuD6B/t3/zRJb1xYkbLlfp8dK64LxLhGnENQR4M7+ZZiMvRKmfp47
5YT5yaWLnkUiOfgvaYmO9Yy4b7esJfGna1wzUOBsm6qNEarWM76ByVg23jM8hsQi
tOFYv2sY6fZaVsWYwgxoktwmC+hI9McV++03ZlPrtke6Rp9NYPrhbHFmbIV7SmMc
PRSr013ilhOmxM/eh4w38ZI7P9uoEdd4ZMPt6kuxTZyrMOAkG/OJIDPmsfX5RjX6
AWKZkPolAJdGimgmvpcp11vaJE4AjWP9QtIVmPXCCX6IMh+64MOTFOB4bUvtjUw9
mXfknPkC0yfKuruNPEVWUSsHB5qQ81ou3s5DInUn2iu0oaeLBsjA3cWLOJHPklJ1
vJipenw2o29/Lfq3j/DSqPOGwI4MFXmfpEX7OlzyQx3+ocG+4D7K8dV9HpkzKWbB
/9Qry4EEI//kikgyOWG0eDYmHY2rV3VZX9i3e3qHmWzNbizbjtPPSiS+cQRlGUKW
ujAtsbn9TwXp5DrwWGq8MRf/o1Fqn0KmzXHRhPXbRlJnzVccVz03a5piUbzfsyKd
ShVBqkylCRTicJKz5rsWcx19sMRjJUtYVA6OWEnBpY6SYzcp9koU6vFNtS7we3iP
v3oHYCwGNAUKxn1D6uunBbppNbu6eku8ck0dOJdZBVDVolGKQ2h+SAFGpAllIB4I
rw7H9XJpMqfYYsRDJu2BVB/aCBOGU5uVuL4MYVPx8DC3BTVcpObMiZGW3Lg+dlSI
D4pgaQWa0ZS0rtKwQ0qgacUHiJXk37km1BZDlr2uz6hSEDGiwD9X8oeBVQ0D1XLI
8WQiW5af0E2vfATmAYazhjNSLiPtpXnqeumfwZO3saKyml4GH08Dg7lDA97Tqj2f
fKNGWhi69IJog+c4OuYA9PLh484+mTctqwXqW+ssd5yn2Xnhe2KV5vnwq4LfTF2o
MIrMH015EEJJbTyxppigb4GgnYGbkoL6UEhq5W8tMvzS9wFa/Fm+TRX3Y6tQbDOR
Fdkl7YCC7v+p4bOHk2feN2R3/KG05TRViwmkx4+mML4bF17uxn79aOmrEBrHun0v
ko9p7nL82iT8XGmTnaLIry04aAODAJrzdZXtmUyj72IiN3WsJM92CE4rfVs8llET
WzUhj6KHXGSJx4mY5mN6NEheOd57J7ZX583DZ0TaxPaPtAtyEkA6NYu7gnIvWc/+
j1y9ACoEp3qlyRU5nd1w0no8lRotFi717AsvJqZKlclwjUHO5iT+H/fvY8bPpl+V
wZLRDuqCD6PfQXHMqOjR7IC58FFF4j7eF3ZuodR56Os809XtkqREeVekQOYd9DJD
ypbfa2JmDAAk/UiiasCiBeg2Y2CJulSHht/awBSMqVj/kbJmhfqASea2Qs5/Nkeq
Aglj9fEiWnEWsFv8onQ0nJNthU6vW/ic3muKqP8O2eRD2sXU/AOA8Qb/3XrwK9vP
3fZRDVrRYYvjcpBlDmCACSWctqyiGH4aoiBzkTjsgzllIuVaUaPyoIQxoyVXm2Mm
a/wbNIejeyklDnEPgMO1ZJxZZHHY6kdXOfEKs+vOuSDaM+p5a2QvYq81C+TXrTOK
R58yqUsOXGMctvF5nNjda7cUm8Buz+WpEg6TZHB9ydi7iD1GGZRP38gFdo6WmhMN
TBOmmYvjbIsWvqB61vX5byAcOVDpbKIeGEPVnyr5V33E4XEKPaYvX+hjVyVy0j09
4e7qZ4Bs9479ozq2n5oNyoumEd1vO61ZthVInUwW1l2zHaxCjr8MhfLIwJvO07Zx
iqsheCkVSLF7ZSnKpA7PmZlk2Z27d//xHuk5eMQF+dnyZbcLH07GLI0HNGBpsj3c
WglATGLyOQUwax8pPg/O18w/02zA3mqpJRMpShWRowdPIUApjJIP8mujNnp0dGcU
HECxjdnLVUy/0SR0jnXlfFL28XRHM0ju7SHA1DDOUG0Bbh8AliVbKmfWkbR2M5YY
5oIBoOh5sx6kQ99QJ9gP7cJQ2GSgWCQ8TsHNmTcj6A+xohhiw1hXjZISMwn58+1k
lVarXoy3hmH9fb6v+hgsyZ8u/rKV1CrheF44B+cj4TYzt5KXR/stxuvNQZAPYk/d
0tinL/NLbFqlHWE82CacYR1p92q2E+oxpCepAnfn6vqKvjA7nNL40TqWc140Bmfl
RMyPS5Mn5OoGYB0cW5366U/y2tR4VNktLkhXUzoaNgM=
`protect END_PROTECTED
