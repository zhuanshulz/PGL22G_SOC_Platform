`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BXicWDZeuQH5feG9AcXrm5dPeVlvfTGEQlNIsNRn6R5/1QXaQZGxndNfbXXaGLRj
h2tKBanpQSvlyaMPpa36Tn8eY+swP+wCFRiLNGAtmMRpXRi7AT0jU3gPjgYGj3DF
PB/snSYmo1UZfd+O8gDThY1zHx9LRIo23JI5vHBYMOyXsX/ucMWziyfcxIc4vLw1
vjC66ftE8K4QK8Kdnb0lsytR/LYKufeIg2tHd35kVHiSfprG8ygZueGshvbIrFRe
8SjZQd6LVQWTBWzl4GAb/+pq8g/+zFy1nLvVwsACA+x7znvZ/G4lypcTUUse9t4j
vnGsubucuDVP8BIea97begp17t/JrGEGU8gtk4ZwTGRqP7fLRdntTYjraDpihuZ0
qEpD336yYylt24W2gyyOADiVQL7YrdjCO0ZMYlQTXivKWI/1oVJoqkWbuc4cOyXb
I2WZVQvfQqWlPvN7IB9420FQ3v0UEfr7O4J5yNyHTmrFBPFq2nqYXxrvZjQvMivh
BnabFyZfmXojNEDdBpuR00BIBdxNo8Deio3FDBvWPrLEOE8tumRO3Pwaqhqekx9t
9CcYSTaYHfpUqH9kYkd7FXoUiMu/qsO6dZuLB6uetWe9/c7vGDd7ZEkiu1YhPTrg
mi1JFeVCO5/dS3s/5SHYgXNhzJ3xCsphjr/C9PUoKN6cFudipw2PT1EuRohR+cek
cXWAZqrLsVaiEgDFaBnvC1ZP20p93OI0XncSj1kLpIr6yw6o6/kS37I1+oqdy3IP
2q6ENU/D9AurBpAnQENUyJ+2xOCs4XSho3dBebhAiXQomHVx/r6tQ6tSxG4pioAB
7QpXLDXFJhn6QG4bu1CVOOvgPBJvzMReMq54YTVQqcaO+tEqoxrJViWHr0QVT9g7
BkSiEyoxXGsfRMA+9tz27zRGCiFexzzAV1a4jX1i5q3X18dD4Lk4dpB6uvFLKJuA
cGbx87+l/pAnhokZvoxzupDt6reHFiu+KaXrhQl6sf9b6gelZ3wbbeAkwpO+93Xs
VAGilq3BxUzqTHEoXNbFm1i2plgUuEdeis7z+tK5/vXu5Bw1dwnLZR/QoCPlxJNn
hFhnbgWY+wDEK3Xs/x3bRtB7RzhlIPzgqw9kMfA4Kt8WC3oDpf9UXADvHlEYDNSz
ZBPqodVgJGBkHEC2ZeBQARnwLwJxlkW/PIzHafUvADMBOeGSO41gskuHOL/sbMAS
+dPOB3/AwjKaZVnefHAwN3PpyaxrHq61/yuOX/IvZ3dxBCeOh5T6j1oOIUbVikNC
47g1edn+3G+8zvR6P6RNP6OpRdyHqhIumxpfVOmVsBs=
`protect END_PROTECTED
