`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Va8CNieo8xDjwPuP+opKqPPmmC+8/D5btETSpi79qIK0sURbjRxNMay540XeXe5H
195ihaYigkVUHm1cx0gTb5hElyTx2lrHvlPo6woOZdkpAwjc2eJyPhxHtwiD+VTq
9gCvsn5vl4BK6+sf5cLCxZRr4Nwp73nWy61Z+/5OtCSDLw5oGaIt+yDrGIhtM/Ny
vua7I42sW5Vz+6HH2TBXNdguU9r6wFhQwl6ML+9OAYJJ6iNozG0OCYBgLbwTHWbo
qybZiW8lch2j1Jz0fKnsLJhXtbwwkGc0nNLT7UOOEnZg/IwLpb25wh5d1fDoEa02
UQfpu6tOK6u9wf6KRMWX23NPUE6WxEsHGEMavxjEwd9YeGg2hHAsLVVkBF9DJrNY
CIAFhmoCeQzOT30VpWVhC5Hip9XJri3AR25yLcPxZ5HkDKfzFn/G914O4FXVUwKk
wcy0FefPgSshgXbWajU+FQpzg4d+x1SlsgnJEqGVB58qQaoF9tVYxIX48f/xPdGV
3Fubb2w+wgizbNuKQPcE9NgHSV7AR9kdpn/Nj/FBNjKG0/HZZgSL01lreRXyZAc/
E8MiTK6TPwojqc5JtVX1Fd7u+BEEOQgA+GX05iI5kY9hujIAHWXBGWZlCc6IvIn2
u4Pkww5mQTw/BEzefLIGGMzfbbe6nh6WCK3bOvFGUjSHifk8ZZgIzmrimsOOGNv4
G2eGkrCjopnuVr31eGvokFKyIPJANDKZk+XI/+2caQuDng6PizFQHvP6sCKO9gJs
E4M64bsXqhbznHDlCU7Fw+ghi971GFf49mXph+msHPsO5XhH0Q5FP0CQPxX3jDm6
zxitZeftBoqp5WvLkTUXUYcD4E2q+xvxr5AA144ZEb9IVyxjB6VhLmZXEpMCmkBD
13MdVjiKDXGMLmNYQEnI/f7jqQ4Gr6cYy0ps2+qoSZ5pVBF7KmtRPkYyTE7TYCNc
dF1bBkAUdMN0Z7FLxy1W6psIngy5dSR9OUg0XwRm1o1dWovBtE0DX4e2lH3jLdic
6+XBN+8F2JyAgmsXGBOquCVPopWmeuEhZ0r5Wdjotg6vqBidPAZRWrUYBJCR7Ljh
vYMfVpJouC8foeswpQq55tnaVFAKnNHyPuWZtLek0b2JQBN9a4tvjVXlT6m53URi
YGCRhXRdFTB3Zgj9m/ag/Q+wk7JJXZ5ihOqBI701RCQF53Zwdg32szLicFZ7+cJX
2++O05IkJWXY229RcsUGOr321Cqp/R3TubTqhTGDv0LLrkXJfFboj11wPCqk6qut
ple60f30OpTxbY9+eHaVythAf4K9LByJdA4O6QMr8TiSX9bzzZTV+Z2Yf5N5w0vl
5LtKgIxDOIwqEYVtCkYpohu9LfBv1JNQMCeEGj9R8g+ijEypyZAqqmUHTFfJGXUV
6l/kVJBUYbEyAXyh0FcJIjnbtm8/gFs9MAMljRAAQvrxqnsDXl+WIHFoEj74/gx2
TRw+IqL4kWOSXigZ2/s2JW6vz7Sw+xcPf6m8cZ779sVQYke5Xnfja+El5aqKnpjC
EpQBwIs6BDXEXsHlToii49dMLAjhCVt+HKixz8gTOZ+9kLoYUZ+dNokt5mnNst25
VgyGeSlTU6IQKQJZJ2yb+XNBD4EY1Grqjxb5Q83EH1x/D+1aYW2w83b6RIMs2HYn
Z6s+ifQt90QdOm/BZX3vcpBWyH66jvTSDn/2AlP7u+0HMls698cEArCN3wswY7sc
gT8K7NKuLzmCyKuRASBAJH466n6kWC9tfPOc0jSoFxKkz7ExVcCGtxs4XDEda15H
15Ho/7bTASBsyxxCbq5Hl2pVX+LO8MJ+TKXL3RKlAiNXukO0hivF9pzFCAmaMbH/
4d2AczYYbK4nP/SD2wKzfFb28LTaBEgbSxthESAtalaTmoG3WDTwq3eAXxT4naqL
RiqbGAkWoU2h0DxBykUwIdbdc8lrB1THYKhFHP/L+kYc59rKUgTGW3HLKkZrHvZt
OWjLEcQGbSnCaCuFCmrRhlBwAwRj0LhjGafUagMaHa24jgr+891yhry3Wn2d2SLO
M96/mvCxwhjM9BCKXejkbPYJqA34gE7HakJiUiETNv4VurG3FeoGgBV4rZ8rGgh9
V4hT/NrLDwwBmfmxlA6t6JVYug+mM/uVsMVYHuen9zkmI+hG4tmCqcD2KWj6kCeD
mxNjrvuzzgTP2s8Y0ey7q3VMovU7GNNh+gufaTixjjS/w11wuUzD+HSQDjuQmNse
rz8DblxmIPTzikzr4mHJ2FQ15UTv1P5wZo+Sl+aizthBQg1nEI9n0J3fu2W+EdoR
SD7ofs9wPoPIaCIZGr/BJp8IQis7gO4aaTrp/MOyEJp1bhFPqCtK/Qe9lg0p7XTJ
VabZGCBI92SYYiSsi5f1ALFzNOxBC0OxL+gS14X+DWBJx6+nmMz1RHgFTSUqtQP0
h8izWzinpkTfS8DnZaJ5N8jTXmXsMrY75EPaWnXYZzX4FJ6lDKsymXyFiFYmW9+Y
2/Vd8/it9jZn1clsMgOUNJXsINH5oQ1W62NAymdpbPwyyfIDe021V8ohLGEWd9eu
HLyi5IWJXj3ep42yxF1JY04jYy9xGeVAQNFbl+Z5H5P4CMVf4KJVGXkMx/ZpS3zs
GLpl6DMCLMiYmhOkmx7ru1fXtlR8qnZdFcqdAVusGkt8eWEz6swOlRv7gvCtoWw9
do4jEergTWQNgP887Fcsed0NRZgxeGEnwQPr5NUKmNy6ckQz9rWNkv/XoFDAZF6J
oBCvymKTbpuGf4aNtZCFr3Z4enhoVlPweAfFKAJubcEGgMGgO1qm3QSIrZmr0Ifz
9Dqck2zOJdgcnh9Rb4cqboHdWIQ3dEtJ7i+nHffbVNgvJ5aWBEEEoUyWgEzrA0+X
olJM8+U9JX4rSqegp+yQGUV/0MZihSJl1twnnKHT5Tv4/XNJQeUWU+eOjDJBoWqX
5btduTjZrAr7tnkj8k3ZzSb6iN32FSHveyKFN3jP3bkGxguNGZDxN7q4jYcnlibb
lxPZT7fN0JiX7AXZE1GTQOGUPD2awqsYqszDwoSNMiif3sQ5y/nBQY4qPIIkO18M
/XkRb0L1uRbsjVeZhw/VSpuoOPj0GOpMuarF3wcdaYtCv3DCXpLeLVY/EPviyIel
g+nFuIsy2VD+A2P6OJ25LwrcMQvS8bTmA2Uj+3bf6OhWvLHKz2rsfrMSCBjNktB0
kMXagTW7tVkF6yIZKZVoZAPbyGz4F213sdpSDaq6oJIxfH7rXYEC5IwVO5gGtFnv
jFSDiOCe5sce32IY+REoFCx7S1tOziKV5LfVDrv+v2uy+knLEC54+zLv4rKXVAfX
seE1acaptkh8WjFhtcwEiyBcDE367WDSrsqQNKvobLLmQNlXM97jqiUpgqCjAwDw
k7K167U+aTv2y7xTC1X+WzyADF1a4wuPZA8j+YvPnKO/HCLPS85fVOIdy0gmGiC1
o8ZQY7p4KiKtcEb1pZhrYB7Mbc3kCFm8xcqkYCGD9Zs3Bb46fApb/l2DQu15W6fi
Z6FMVK84wyPG86SRM2Nye26VRzGiezmCsvnLSCjmdsZ4KmK4jji4PM9tNM2ppVdq
FdgpRg9Sipd/+YKwBfxSLeKwnyEH+3YZakAzC3B9uyO37JmwWKtPrfhpITOJeaKU
50j5ah3KyZO+gPjTnlKQ4zPyl3Mqtp54Nox8m9kQoHf6MNC5qka88MzAbww9CoFN
eMY7BcSGb+mx+fz45nKe+6IdiqyzK4OQIS3HrG34hmsKbZzx6PMDm1snfsY+APW8
AqEkCjUM8SWAEwZNrZ88PXY7xW2glKMsX8lU4H0TyNNYuTzZVTup/TeZcyNbQpBo
TYdC17cbr8WEB5xBpEZmZ7rulPmJQNWbiCWdWMH2qfXKISOxXFt3Jz/sdEEvcTyd
CXRWE0mFtSMY1dtioQZHVRWvCXRxg9wbHWGjBkB5/EnhQpJzunf5JqCs/04kOH+Z
LKx9csxtObmJgCEFzjuo4na+KiwqnR4FrfJ+eTBLEaE+MOs0bZG1HQv2LCcKfHt5
vgjp9bTgT2YI2j0lp7C1VxL/MfbP/aYtRbroe2Xo4D32uaClMY+XTznJ4fv98u7n
LzvVHb387TlRFaV0aj26DjZBx+4kdzyODGFIyTiICQ9J4UlP+gPOucfOILDk1kTY
eAohxj84rrM9rNP+IPU+Z5frT6j+oO2x4Z5y2rs8eFfNg15B1B1C0e6FKrppnxqk
VtMrriVHvmXx6Fy0IkMOfqaeAb8uLdlExGp4jIb8jG4+7zRzcNy3cSWKfnbTDRjY
8HYCBdXkILzQpTGc17vMA0BAchqYkQfcwjG0YlOMRn9p6KB2N4TZLL6y9npYzmSZ
xGXSZnSXfs2xyPmalFDIAQ9Xi4N/HanBLcxp6Pl6IY1bpCugsfX2gWSFU/IP67sh
pNTvq+SF2f3w1kseo3H8QPUMzf2sYmfRSulTOkvY5iynkzp79+g1b9JGrPlX5D6+
McuJuw9e0aan17v2gagHKZ+MAudoStJeIimGB6vZfR2OQ554EHm/7a6CN9Vp9iyn
prlQJbxgyaaisvMXb1pk+B5MEFkRHScTYQsYk7O4YDzeTZiz+C3ZKVGdEDT5T4m7
zRhiLIllRb+GwgEPSxJkZRrkTuaHiOAaSzjuPMuZMVXPatEkMB5wZxbPOG0JL2ZT
Fg4VDzatgFFz6L2wPr48MMexPFSxaO5Kftb9G7f9UR7+xk13iA/kmA6DQsRrRMO2
XKbghNuIFGH0ROgcRn1GeFlcRGAJcgVSyIMBPMqLuS9VJzZIMJ5OtCK2hxCYJytk
pVZX1+N0jcovINE2oHPYfwwTkP9TEtonE/9QtYJ+xDO3a4wbP6aFw2231QJC6sM4
MPimx7owqtgB5ooa2AqUztWyT26A7IbtADsKjMo/i35b6Cu5f0s3FK9XU1WwONYU
JUkNEo8KcCzMuqgXmb69CvRvmlmuT1lxINj3IM2bWlxz/c02cAjKJ1UIpK7O+u/p
W0+rIKW6rtMHtNEDPKwXeZf5CHbwDN7Y/sVEvsXQ9qZ/ZJmw18GHrZf8vcfC1xEt
MGsri4Jk/OY4qybm70B1jQrX3f8WQNHZXnbL1l4sNFtIfgszelW5QSGwnUtwq2Gi
zNqFpqz+dS5Fe6QZACLTFHej8EGM4cvTJOWty56XS1HL7wW+hSquWCB2funa6WSp
iR8V77zx+SN9F6DQ7uqogt4lRCb6x7gCmVGDNN+8QiQbtpYTVG626Ul4mOlcQ7j0
Oyr05XjesQWPyu76hP5EJd9HhQ+TYMz1W14Hcwoihc9lp51D8Nu12KBvGUHpwMSy
eJCnklNadV5MlmzcvO9QlEcHOZEgMkUa6xEe4YBc/zKNlZU6S7ITlPDZMcxIBhqN
0reOpWsnC7Fc1+OFdFJ9dyO6/ypOjP7tUkfwQ18j2/XdzzX2mhxMPrWkcNXCz4sO
NyKdG2c9ZX3lEVGpbtbd4P9r2TWcm5wdoQOu5oPTOZg7XdHSRYxI/Nk47MnXw4fX
i8zdEwxVLpQGqxQ9EZcMk1w3bJD66GJUbMWHhTd2yuFgSxy4mOW7euoVm/L9HTow
DHhRuwSgs54NirSikkBvWjNr+pI7coM/uX0mUDRQdwUbmewvhIMYUeAKWzljX+W/
f6NTijswYzC8jbzPYI4+Lq79VwxyahtRJypD7jXX9DMkNmgpTULHCr9Wg3vzThJj
iKG9slKlQyoIV5aOKbKq4pj8TiYKE2bkxmx1dTb+7s9CbuM/yUatBKJec2dkP5wF
TdvGOne4OaGUTTIb4zw6X90A35i/HA8MPDVxC4r0vP3jDj8QdmI5kogfdtIdenK8
e4Yy9N1Vbt6sGHi2B+KpTBp2OJWzuUe9UIaqHam27V+NVhvCcXH+VH4SgQbYJapq
iDCYcujU6zSt+UwqOGttOtNWFixujviu2qYkJwV/pMw3jJDANLM4+XjFzmftvX0d
GPXwNLAuIMjlCVBb4SdLxZJSHS7Hs8qwRjTOM9aOP4m9Xyp2wwrZwfMkAiWs+LxX
0/spEfukpfpydtG8FLlcJMldaJlmYpElTWrdYW/0NUA4392UzKL9Zv+Jt/gTfkid
0ZISHDueGrnrb7yZ+uFa/0TDZroWe8siaF9l3FiAaNdw6mrARWqsetIxdQ0YGjEM
NShwqlcEn/tf5zAn55Jud7ZrqTBeoA0ijtRVegJL/Vh740xTFSH0/X9dVLYZo2yE
FbMUyaCvnBm4XVw8gD4OuLITFrchRX96tIbfx1vKBKuR48gprKy9h4GLjkZBbtM6
cnalX28CPQ+Qw3Y1xOyqggIa2TcIjyvbNKXdKSt7cjeF/uAZebXllwHGiszOzNMB
4T0X4OOAXyFUBsCkp0g34N1fC9R1gAg+08EKesOdyOanfrUhxYada3N2xhzfbVUj
wKA27sllHb5Q1mD35R1J0VjGAFszv4zvLjqjneYvj5oC2w8QOGbiS/Wo6Hfm3QIt
F4i5O9VooPjwy5nur/K7lH3QLw4zFAWpmjGeAuE/R/yoRebPcU9FhWDOGzj8f4K8
oJaHmQe0aovx+sFs9nWMScZ35j9ESSYQXgFcr4hax8l0AUSe44R24MgUOp9EyUbz
EjvsHw2nX8OC3WQihi5CB8QTFRL4KCJ6GWv8r1IXb97e8XkOUeDyaoYInPAcpld/
Wjkf4Ttx/TGatvr+fD3tRPxGUiSoyU5FFedyZgH4361M2oyocRugLgb6T4plIg7Q
7WC/P1qBXEPtGzN7VD2l2SOxlTSW7QIY08HuKbKMZaSH3mSznsTeqfmNLfvYhIty
oLi8/3gKfDz5pmBXODOUzWiA9EbX7ol+4GvsV/FNeWXePx6iuapbDgrPZem+RD8Z
XnCegUAk5B596H6wJcGAvHpgcp0+bt5yVZeyrD7QQ3ILesquGu/xFekmNIV60v0N
16arY/TJi8lSZ1q9l6umb1DI5H9TfLGX0DO5ExG9Erbb/ZLaxknsBSXb0RuprZhW
r3EmHh8qfR+DuoTT19sADbWR87r10Tu2pH0jqUMHWX3mLOw5pHhOWp4E02DdFHh1
hGPHbIYoXVXeb418yyUILX4CXxtSFX5pvecDes8M1He2Y/1RbKBORcDeCOrz5lnS
vASmnoPR/hQui4mMemQNsOc2LM54hDAZflHzrds+0zD0/vYt2/XVWhqW+8Ocjeo5
7etNITazeYmfcKqWiu/8+aMm0VShU5n+0c2XtoJWCrLPghnS/8bN+qCikCIXVyfF
/LiChgLv6VyhGvq2EETEMOZ4ufrQjEbOKiXLTG7gGAoCkUctUKWMfyBL1jjUNveq
fXoZ+I3YxscKMxR97lDGe7+aSXwYlruA7QnY6mfHm3RNmx1DRWV9HayHz/yOE7+Q
jqsyXmfhr/1lO9a5KYAU0K0U9piTSWtbY2RGZgogccR5QWn4WgUY+h3MO8YuMluV
iAPzhkCwxv1nOn5kaTPa+HBeaFgDcVDgfueXcg0k8ItOHBDqcWIq1Jb6NRdMxOoT
43WAmcpbmCftM89aUP2ryH/gN/zbw0NHJdBGmIE7pGMWPqWa7nHR596+9emFP7Dv
+tc5iTN69io3hsaDJ3GfQatG3otafOzAdtCus7ysWDKKjjZrK6RdSPCv40H09A7o
pre+wO2V52OyPefZoPWcEgPK04cR6c8nsCOlNZxfA72kEujLMcm2cdtAmpGccFu2
w4AYKdH7sGAZOOu27ZpEuuxQCSVfiBwME3ImsnMzZPKGpLt2jt2nqGcjbXPNgaOz
fFla/jf+PmEymvUOuIVgXWvo6bWwEiwn/GpLw24rC/07Y32x247m58xLekHUC3lf
zFb3hI2/d0Z9f+IuF6eR/gg5WRsldrUro2V3bbNxGnLlZ9oVXikq/oZneyfFExdF
64N+AkYfRzR5MxeZF8v974IXog1f5scwomg05KBFCh+4pvjjsDia0/VmaXThnHCo
az7qpdsXAi205AkNs6lp4gzwYTs1V1q4b9Xyh+1Y/4vL2+zdJaD4X63GZY57gq8q
GrxbSjq8KaoQ1ATUMsZ2YYZGGfS0cWr+w2yUalym8kdd/9Oi1ZehukjJa4jCMLAK
eqdnLUmhCRPivvesz/kbaT0SSlIW8HCbXT5jHH/TCx/1fA+J1Xwj1zEJ4/Tkz8WW
ZetfAh/eEt7kl2E3juJlJ0vMuq9W1ROsIVc42x7dVcKILk8Wb+TW1zOUK44extG5
je+U1a3Rphk9stHTFb7ksEvxk1EFsgEe2oPeQttHWDOKZ09EwswBojPHDNtA1ufU
7AeUf9Ixq+TZgyfPGs6nnY6sqWmdwI5idDitQcnmDKXd6qe9wUk6OZyggS6VDGTo
LeozSzDmCIoYxEjE/CCrsUAjXbzOWXGWfGralgWqJIZNYsk7wHv/pDuwG+6HYvRH
OpP+siT7W/ZMjY34ItZ17TCXhDVLjQi7UXs+XZM3tTgc1+g9X97UCE6owtxNmnRS
3UCrR/vwntUPrZtnbHZ/66NtgtRO5cFSmx7zyKXTNHNDrKMmVJ9lhAfS58iSF1pf
4xiYuXsHrOO3NqrUAOnGPVVWIehx2GVk83GZiYqC62zFXq0s2Q3qaWGiwQANg6fC
B660aYXaG6qB+K76I3yCDbrcNIE2wt6vrG2XtITc3Rl+tzGpfc0zdr8d/118LTgT
27X1NuPCbvozF4wL4rfKdRFk9rApE6FBKJUWGj7llN1al5T31Lag2S4T93YrABl7
E6K4PN+fOg+ZbWxKoFG8IA6ZFLRzzTePfAU0WOr8TApNDaG+AGlj0Uqg9p6XthxD
pNiIFJyOvHVG5cCJ9FrFoblwboKfcvzl3j6nMvQmFXdwH8+MVIfYeEac9RPkyQXP
ndaQ1wA+jH1cgD0UxqNUW40c3ozrhOpouqAcNdvVtBq2SjLO9daWwulNJPU7H9+9
YgJUGvqeSg2Hq4n6WIABlCEXAjcyc8XyYR5Sd0mXGe7x4gC1YRttCVFOe6vOE4e+
AAEfLbKx8R01t6ouwgWzZioDgptt+27ddgDCoiWuMygXIRWNQivHFMoX3IaolwWN
skf4JohZJneosvi1Pxk8mjSkyzTyYvUikRHg12jGrpO9sW8Vjm00Jn9oNQpo32oX
ZOk/lncvE3Qvb8inpp7cBBtSxMsur4HgbMKSZBbYdpZlXdvua5VzJma1KWDS7+KN
wo+HQVrgEND1LL3gKchEBi7RPhiZ/ZyqOX2zdmpt0ruSFySPOoQjWRsYmCb9WWSg
yq4g7gSKXrcb/SF8jNjHaGOTUvqnHvhyfeXITNdubp0iw1IunKzcNHiVC/PYJsaM
xSW42vLOTFaMpa0/QUpB12twc2WI4xuwjk3eXSvs4vYi5Ym2Eq7fKr+gCIwOZcNT
K4LkczBhChoq7M60zxfEjhnRDAQlVnc/2gvdm0u7lL+0aiBNQBTUIzpzwVnF+elY
CGrPXZsoCiaR2qyOQAGyPk0ArgqXTNgDY+2wRFCofcVOtPB/63r1VdUxGHRllgfy
l4JaZDQKLJLc8qIgH8fNE/6f+fjeyAL0f+l4XW86HleI+bOkIZG3WNEs5cOYsOUF
hx2tyXqK4YP31KFXgDib2OU2xK1rnVb85kBb9VrIwJQvCa86sckr2DPD79PRGCH4
PZlffmABtiBslk6xgkDV0aXSHGaU4epRuTC55uSWHIK1fieMA/c0ZQvAAHP8srlJ
CkxbBrxghLjtYvJScLKUouHZ+TJDAypa3kBDY+BtAOtmfc+sgxXhoLZwTXyQuIRN
cVcVj/pYn5bPlHiTNY8FMdPdehwB9LFJZqDBrWuQ1YW7NIF//LnBN9lal7lJmghx
W/O0ptTneC7TdkqOiciP8s/uW4C7I5pRkWnB6C30kVO0KBFYhrLu3rsqKnrKVxO0
oBRg/8owxFDBS7+dCsm60eE02rMj5Ct8EtqCdoyIssmszjHTeN3bJzg7AgYfFSA8
bimcWYcW855e9uNXT7yVugpDTdS8Snsu7HWI5nY7nceC7unxX5wdi/7QGAgfFIsM
zjNssCqimFqDNO1WO5LSSqLaqb54lEE2WmVK6V7YwyfJbbS5/5n7yWeOExiSx9XW
EPIEUS9lGfZZadNF/SSMwnpC3mtAZGI9vNDmDoJLAcDgYHRVE4XMfAzrx6CLIxkS
o4kUiWaXNCCjMihkOeQm2NBhw7b0weslOdx/WDjxsNyGbmJ+B6iIBhOaL52T4OTz
coUNHUuJw4pFhXkF2veq5XJz/IZqijrHq+xhFeouTqgNdM16BJvy+t4eYBF/65RX
u8WtSp2cEqj0wAjM73kJKDmZORdC7AO/+nra2+zyPfz46YUN4ePIV7ojn4AUKzo9
LjPuXl8vw7qTEjeoxVFcY8lbxalTAg+549xxcoPHUtoFI8KKmRbhQcX08BpRuQdV
xPluuBC7FJf269xidNHK9C2Sf7HLsUrBW1387ZnZSX54YQsMsidWKGDKPEOiTl0R
Y3ShbRzUVdVbJmST2F/KroUnIoYWeDAuJcs5Xr0dqcHPbO08EFbIQWBbYA5qStxF
Pxo0vs5rm3LW7smffURLV8zDdst1u1KZYyeikS1Q8oCHpvuQ/6u6TsIvrXkSAZk9
x5q5yU1XOil2GM2G1h9WLtfkbFTuCVfjnkv3L+H66V+aNPEM3qIZe9bC9WuJCoL8
j67HzLJzpbDupb/Tf4WrwFrsgWdISBx4p1BhIgVxsBV9rpVmyvznAWzk6kwEWNWE
IA/XxCf65bMGSXDpWnyAVJsgumFue152jvHdzK/pDWBS2/142tqOFBLCj0dH7L1T
yfCs2SsxNAb3oTC20B9AtN6wCjbUR9kRhEa1ox5cowKWsSTtmWznc5TJoP/wQ249
pUBmONogj+o05BFuWHzX20VYDF1qF/n09gHhIxdPLSfFF1YMPKcyVRZTXJuegR08
gKDvI2w+gRdhMo5jeu1SanWlqn8Wa4y/z2WvMUrPlGPHyz0Phm2Lgn0d6IKydaTc
pG7nU9Ihy63syDSDQbJFKrK4zomnrSFo/+WYCj1CnAOgt64qhyArhRfR0fhlgZHy
WNxUQDMDNppLiZbB164LfKTKuzmZnW2GjrMafcKeA/LhNwtoYeE4d9HE+867efUL
fzz23UcxN+9uJ4cd3cN6Jk28MqN1bx3KVYa5wSvp6o7ePzEFWFpZIsuBdKqGC4ky
E/U6MBLRkKrTobRioIABZ8QBid9NnhjClltTh3hzCvTSy4IDOh4+EkZTLCFuW+vd
Bb+peUNcRyys7ih1aIk7jUdCM2q5iSCfYe7HP8AjNRsWe0QB4dIIZugv35OrJ1oF
vrOJJceuKdFXZDBsjMphjMLZXJiww4OtrDYiLpoVWEOzPEY5oOW/EUgHZhYPbmYV
8QZXHBLrhfFDIFPcAh8sAQ3YQvZRTs6jP4w/L+P6fw7DThblo7VZoXhh79D+//JS
UznrquiopLS9V5UImoJKKHJ2BEeGKKHzG5OJjk2nn+2IwBnqKolQf7+ROGZNs+Kc
z1Q5PrHmxUaEn1+AYag6SCyxiS49uFbUFXXGTjJfXqKgCyq99UrSDnhrChHN615x
mBnyI8+wrqxkzig9IH1O3uDtFW3f46JjL2iDUCoL9qetgycXYvb73P8xDW9UHq+o
CS52Y6iqTRIq1G3IkQbO8obDij9FXqoyfs5uwdoCAxTeCD4dRJBvLICF32Az5axq
h35XpxZ45JySPCloaM/p+s2WlJATIGEP+uEaPWDDNk7uQ8CBOV7cwHhwk8R2nTyj
4/rSX+rCLDjWQtJQ/4Gl06AT4pYsQgnDmqTwK+kIvKGgRTza4SZKzop4wgogekft
Vupogq6yqWZarhmFypzxebbQUCwuNfcV030sMeVfB16TQS7nHBpIJhKZKU9DB7Yu
TaVS5km19PAofDBqzmiW66UEQMee9aDh3I18mhKiaeLkyYRE01E/7wNHFn7Kwp61
JzTCnh9/kG+IV75+cna688bLW8kct5FpmbqDgUxwBl1PJaeBWQzE7z9bRqEGRo5T
9NLUdPbDbbjwMYB8vBn7bP+xMdq4kzSmj54n8SANqicP6CKtvnS3ER6DP7VOPUea
UVfah8leS7ocq1TP7DPMjnKTtj2I/iIlmf9EbHAsNOPOSG9N8i/zS+idXCTrjrNK
/U3wS6UQ9+he8f+IwXvPekeOAMZ9oixyZJGbHLqohiJhm8M3cjmaPUmjyrCjEPK6
gVhWaEm5TqWZuqQNh08BXRXgk6tsH0oyHcclcTo9xDIDv5E8ZGiZcAP32QP/HyYR
Ap2fn61PCmkeJidz0XE1F70bXeqFxTH7jfYbshpk6cBAyZKVBuJDyfHmEDq+tjB+
enGt2IG0Ry56YA+UyCIEahPSHz9NJC+e1dM3HTz6dk/x/iAbUUtpcv9GZuPpHkkb
ndYF8GzsFJkn+hkqd/duW7weFIl3lekmR5XI7vyNye0+IrREuGrVjWbL5PJ0QDIw
6B3c3ESO5QbCFHDzDO8poXTR5UMY4YX69c6YBTX07RwKk1j1Wq8NxwrFBEsDfPgJ
n9RTUAmVRe7U8b3jiB+LTcgbCTGWbji+l/4Y0OwM2klif/CpUJVMzFaL5Hav9+cj
rZ9nd0pbfQgOSnQ7fGsEYT4+Yf90sGUowqzMm322KV6VLb+HuRs943PyJdmNPgO+
dpLPoZWdNmV4UKCLbL1cfxH5zS/iRUo5alRhYapFk01LhHRXhrvh8K9qmTZPwswC
WObxa2R1Hd5/IL4Q8hlBhL3bmHlAk0E+MhpTULyOo7xlq5qEAjB5bjkybtiM7r3k
VSLXMku/RSe732jNlB/5JzghYOhAiQM01Bcz1Gh5GHg+nelu/j966j0F9G3vkzu8
m0JrZFucwgjSw6FwvJTxYNFWqBs7flxq5IDvoHsLENGX8j16g5MCEhR/PgZuRFOD
hRdA8k4CXmBhqsDMF1CoYLF5licAkXwFxa72chokQhJKUliZFOxP1mHj4/VwGsnB
UBCTjwpM6e+18Wt22ebuQQXGpJpAZJ9VEsVXvxSQ9CXJ4pBrB3fvHRbA856fM/n+
Q5Lfq1qiiU6KNiYRg36WJzEYBxWy+wl+GzOJoVdFp/RF7vNWSsXyDcfIrsDvpRcW
ux7IHUTE32BKp834L2y7JV8ZkJdXyjsCy1cWM3bLRPT/pl/Gcp8TWxgN2XH7xz4V
wFJxA5GMah38aK534HXyn62YGdW8IVCGlUZnKiSih0cAK+aNOdKIfNsRyB8XTnDt
9C5h4E1QjRRszSsFQHbmJK2yoJU7opsCZQpXHsc3JSQ71O6iVhIPXxuTQ7vIPYO/
87T2Hupii5iPu9t5/sAuBN4l8novSLCObhgwLURC8F38nRSSq0Ac8ymc+oHKXkog
z13Kd6xQiorzegBMWOt/YBmfTxCx7qu0B12JY+KasesXegWDMRAeqb4E58NCgTnZ
UXAHYE3qacLkQmC9Eh8IIgkm9g44gWzJ33wc455QD/ddrYNxga862+gvREW7SXcl
Aegvtw5kc0+8D2pKShrkjq7arfefUZl1titWDRwAS87CD25SGJbwICLGkPNy+/Mt
55W1ZLSOiVAOm/xa9kxgzlQCawavErSiafd2TITjw0UusJUcNEXGZcwiY2RoJwfi
l0Dny+1LfeZ34nVViyVLeAyC2vNfjA1JrCddMjqOniT+jqKvVa6IQvf2UJJLtpI/
FzHph+cLl2zi4gexiOUodDNOUBbfZfmVDtp1be+ZU5ZTQUE+f0+plagIPgboej2I
qOl8B+N8hSNFppHTOdowwrstv2gUjUFIjSllrvKO5tljMLLAqXuSaYhIH188XkG7
eUIXUcWZw/v68Kax3avUIFnThrVQ1Qua73/Rp1BRI/Cwmdt9B6q9p6Q0Q7qWkw4c
NgKtFTKQ8SMIb0upUy09OzknypBrFAF2sJEkalPb6r0DDSRRM0E1Jm+ZTzULUxnK
psqzpcWo9SnlQUSfwdSAD7TGLv46tZgoJY/Z1SDElENwcxeDBfSK7NlDT7EgpKdO
inRMvOsIdzDAY5s2T/R9Ro57dDMMTaInmiLXOcVYPwvMVQz3wjC2BblzL3RS0VO+
roef5ZhQoTOJLv78GsgMFbE3KIvuubT9Nvf/L/PMYyHd9nDPoqhMQ2dl1+Yp9SB3
FTZOfxNN1Bu9bqMm1q7huZuXireC34HnY71yZnQDf5dgm8wJd1GIqusrkxmLqljn
TK4tPJCgn6K0nEwLqVABb9KGD/Cyloy1BMchrpF+dFu+EnVnX0edfEucMxG0TXcJ
BuSd5iPrPH+UfVNGKuwDFRDDbrmSjpwXPsjjtPCiOye1i+S1GN5SWIT7/DL9bFbA
6sYv/ISGGm4BnxjK3EgBkF/PCyMa9TfSaboKAU/KkShG7jXWVRkyillGZk9Qhk+w
CUzStVn33rqxgTWUMIeA8+UcNUYIrLLWnZb01+EWj5HT/i6e9VenjQllYBZxOYdg
3FlgSEoVf2Gs4FtiqqoRKsRQb/8ygl0PP0xBCTQ/qIXNv77LPSzoxGAMWEe2ENlJ
kpU7sVv1fFFzrQwxxQGEjYYqT/NS86OcuEWyv/AWUYzyitVVOUQj+3hee+btyJpd
1wm15nBg8isk7/j7uj5L7R5td9zIdqgRPuC75Z448zf7CZPWGdXVqd3u76JQKN0e
5ZkIveJdLflITMSFYEOy4erbS7Iy2f36ZGjpYVepxWOz73SUu8WRa6M63mYVoAdm
yUoJCmMYeZqVWdt/kl/Zk/VtozLnXCIeZ1wTNffWXhL93CWqnllhMquEoQmiup31
Q3tnbKvEhV3lIdno1mrJ/LIFNrbDYGKoVjifjtHuWpvwT8aFQnuBupVjpyfukWOe
iBGv3yM+YYZLsNNHIKqhwvTeU9yOJKk/gEF16cQfjk21Gb7nKTlEiKqie2CRdtkV
1hgL5m2WT+xLyBfMHGKxjoKn2gwzMzp1jcYCO53Xf6I/YXge9nOqRAmVps7dyjb5
90DdaOPPC7Pq0Ropxa3m7EPTi+Cq6yY+OMWhJJDD28sEIg0TyrnJcJVJ2RUM868x
RCRDM46Ly0rtX8YtbJreHdflATGmcm/1LOWqz18ivw9BmeO2kUJmUz/8buJXRzGc
hS4It7FKXtdoZvH2rYw398tcdO06229dvsDzYn+KsRAqhsVHYzFqX+BvTQZXWUCc
I0OlVKCHbBczwyotQfppIUUOMHZ8WQ6aJ8EGWQJutbN/gEmpK3YlaTkyMdvZLViT
6m1fPEl5OAj6+PvU7VejIgDrI+o+tlx69qnQ5I+yeBdSMulw4BmM0Toh2yC9lk7R
e/XHpKGnO48JD6PxeRBvvEQl6EfQb+fNZWaeTKJYI4VVzOJVxY99TYSL8zleXhvX
/1GwJEyMTVnEJvGRNqouvmYwBDZx0ScFqFb6xybhEiPUthejtnWC39buZybq9XGP
ycwyRZ18igejX6PxlG5dTfbX2yQDZh5oIE8LakCBKv2EJiwfXKMoFVcxj4X0/sO0
Lcym/wuBIushkD6Wt0fHPWlfn5n8fiDScjEtAahERS3fv9u3757BjNPuktFI7qgF
Qz/1dSLPzoeOdqMPm+aOhaaUoKd6RWUsNnqNdgQiaoyBdWuRvbwysxF1BAjvvohj
wxdEOEbjcVu4Ug04FVGpyeFKQkHjvln0dPoxxzKfOuKfVl1ydSf6bZZtJ9RsDVgd
CD3B2V64auLjZ2iJAc758yGB+sTbBA/96DNxScNc516k4L0yj6fxB0kVsNi+at82
KB7OaXO/bfvd2JOWu+f++Dg1zF4n2DaCvUhD5RtEJKW7AaRlJPgbyqQfy3sz+Gl+
SEiQ2Q6OpntUbEA9OXg/yA15ATE0RiXWT8PkQbQNahRg3fSKkOSiB75yolYLav5Z
pFXiNIFstJGG8Vii165KsTRqB+dVy/JViN1aJe+rtKprD9BdA5cFAYjwxdz1jzic
/L+uaTQVNQk8BKtrldYfFbCri9lVwzyU7h59PY98caJsH5vwwpR5SlQ2iFfU9O6N
g1FAwhIsP2GkryI+LcF87FkF0+oRlGaK7BfH4H5Ki2orJ0BVyDbmGW16zJlYwZOR
QamWbQgQZVcqBgHeYUvdlRJtIYoZqEt3+Z97ws6Na0r3ULiit/X6CBxCI5GN5tFF
1PpalbeEc2j/oufvHFpe+xoSNEKxKcaaAwkhTiCri+u1t3YsiGC7beg7LjK1Rc7R
ENqZAj0jvS8j6gK9vuGL0wp+m5Qs74tCrBYStQ2jRBxzg+Z3V6XtDIjFs42dbO8i
ajSO3bHolmHlyKl925g8ZtJt60HU8rshRxJr+i5IzeUdexWH/4efBbv4r+xAfChQ
k6+F1excPh0ft12EtcjDeP5+yzp6y/z0oL0ODh7Yv52D6Cby74AohILI7qIJzHlk
iwS9LMyTKmOEQX2/HJtrySola2gTNJnZ+JpW8PjY4FWUjH4Ee8JTrvBMiI1s8ciu
j2jEXNAK6As6d/n4ufWd4pB3WCyDqqbI92Dr6EGPKGyyegxHetMp9njHLJzkMjzm
vGZZbBDRLXBzCBBjt1+4ADS/yg4L/eP/SJmKsgD0nBbbi6symmfAFjfcH8HNC+DK
N9H4ptY/5rJpT0giW1qVZyUVyooEEkdxQG2ORUL7xAg7sj877/RUgnpZmc0jbiHZ
VRdQovfwhIp6JQXUJQ8WjuWC+FsWcbFo43s/inZ8LviqLrGpFFQa2pAzVfEuQA0s
28XfwxH53ax/nzRVvxD3QpRps5jOMt/38ahkhAoZkaFli9rcqIxlfwaznXpxE2IZ
nIss7yl8kveQQANf+nKtOb8fJpi6tgEK3eRZ9d9NOU3ZqgYTWiiF8B5rly4q/cpA
oIgztM2cpzyZcgVujqTROx3JGtG5j3xY1cd1gzrsFVfEw4DhGLirAIVqVZUXeJAq
1/UggK+851207YgySBYJIjXRwD6+oWCldE/+HNRv+9xJ7tSS/i3jPkmOekQ/RYoj
cTJTrU/AXI0esvpRP+vXqSdyhw+rSNV8SRIwex8IIMsO2EdxhjubeeUUigeoQquA
ZIqGI6He3De27QywV8iFF59YH5eRufcu/dL9QLf3q4e/2KP7S9r4ZRx7O+TnOEy9
XkySvElCu4aSi8keQN1ZH+QAYI6BLoYFkKUs+wvB9LMyxUOLldYQjfh3zxBj3IXf
06tx31LvUbLe+Sv2dNzR1O0mGXFLt9Z5Sbi6VHiLJMs5j3ZQSPJ+xrliROJBnW/0
zvN+Wssge5hueezbf2WD/CGsaYB+zcKU+dvWz+lY376NB7uKpjMg+idUcGi1qfzG
59Cp7frFKnzX4qsTC6mrF7IJOmqwknlNZArm9fHeJYP6CmZ85jcfnIiwCnkdt/61
VgER588WN2dAuu31dofcJBy0sly41NtTjjzZwYpCG+eFjyGwO1jdzQKUwaCb6+p/
SuzDzDy2tCw1H11rlFZOopgZLPg4jiPWDSK3b8H8z6DVSK8El4ptfwmSlIW5k+OX
eHHGv30lRwHhVtpBA+XMZ5vkbFQ/vBmChnA02bWJq6ZSboJu28DIhfiTZm9tH5GB
aWR93wAHxmGlgg+mZDKUcpmzYD6YfVu+1keJnhkJpm9/LmTPgE1dYof9iwIPSFhm
VEXS4CrZ1Te34QSkuRI6n7LxXqCztOB9Y0bZUR2E/TYVVtAEwtJbD1napnnep8q8
FCo5gMJsP2/7IFbe4S8yuubDrmGyS2csonLYjv6rvsOl9T8gE/fF3E3p840EHHRJ
U/9XshS0rku7pZypMrPC6G1qAGuGHhIxCShsGsEf272fZbanaYIuZgPuya2VbtCz
Ta4GZUg+Nl8ieEOwx74+G7cPU23Ha+sU4deDGRS+5oiJP+ZDOzAdOaTB3cMKH+U4
bEOV2uvvpZmfnIfgCXa1DkD0GzO32WKyh5pQoV5PVgsknH+GiHfwXj4rBc5iFyEu
qEcRh5RryvqXIZiQVqCRgKWAwl318P+s1vujUKndnfyWpNLRuDCxfEGZliHK4rD6
d6jGFl3wzChee6tTtXeuITsDaSeqA4voZV1YPgoXxzcY/84SIlQws9MUw748ZvPm
bKheYajBiCfnMYkeFub/rtFFuTzMhkLQD1bZ6FPGF1P2UpdRLlO6yUDx+0r02suz
8xXXkc/iHIO+7MX/vZEyBDkfqF1y5W84BvZosWgECiZnX84zbmXphndlL/MJ4F6a
DQVTo/DDXVfBQ4919WmhKoDSJPaqSPUV4Ja+nIMgLB72gcaUX8uaAw5oA2gPtmvM
tINRcvjCTWTNoNL+Ku5X34i/cE3LvJf9l3DDf5ITvDHQZMaWZv1qW7zShGFTuUPK
Glu4eaMeY76zGlVZmdTuq4BjDM/MZfFlz3VXX1GjxyHU+LvSwHB7hi5HlRDjoS/c
JIYuEWZZuaGHIhCC83f0sdLS3dXGD+qbBdBKYBRbiU2XjnibHLToYrN9s0yRORJu
RyMT40QBIb76ja04ospAQC0cS3hbAvJaM/lI0fnkJiytNHBmEHTsd+63Yf6X6xd8
lk42XGqmAfKIPeWcJ3ehCHwsnHHmtpir+u++xMS6IWi+NFBAyYNOIXo+olc9PsKD
S80pYlWT7gKWmQ9RlbR+mFfY+0GJznZxCva3nnLnueTi8PYMub5NS9hw4jsQwnL3
9euyJXZ1UtxxhRVnOGsbDfJ7tOxtzWNLHIROrwdqbPUS+A445WF8cH9qbXrBPxFw
gc8K6M5rVEv5dWCVyWcD59NAYpJr6dJSnqlKqwEAvUOyajiQjxvOA83buenIPZ8R
VNM6C2Xrcnhrp3dAArtrwssJ/vdo2ERyujcGAaQsuy5ZD+iLCubDKiw/yqTwLI8E
MqwFKtRHSAO0R/hVHicPRNzbWG5NC9al3Yd/ZcuT+QO0yKzVDNpK96F79NUSgHYA
Qwq0nlpLTFY/F8WlvlIti1XyiOKEa5IibnpmYXQVzJJgswfGWk8Tr98p3GtoKRYI
L8HratTzyQYHsMiUdJUAROOTI5mQvqCmN2cmgm4XgFYR8Ngt8DF+4isjP5gm9mMJ
45J/6qG59OGyH1O9CNt6tQW5to+2xytbIVf3D62ApdHYBf3kY73b+/p26Du7551B
5DgAwhaB7kHYwzOToFH3Zd9AAa8peQRTI7R5AQXiAw+/7uhpcp/WHPyI9Kgssz0b
j+Z2APXYunB/CinSK3wvQP7W9/ZAs2DhyewMZOn59HFk+2NNG8BqWonq2T10Qvge
k7NXoMtAHv0KVld0UxhPHX03UZFvlddudxW7smwpNtLxvwvJCIeBB5c5gb7ishS9
gCQMd1/rr7QAA3mviVLKTw2ZB/7ftP5Q+pkrN76HgLHqQ+HwaWr0hPadFzlvxvGJ
hHbVIbZFD4Ss++Lxe5AU2+LLaz48rsST4OrvvYKNlZXaTvZpBAt0sZ+4JaQ+2HVA
EY0HmrZ40GUtITCb1zK9RUDInQCxlFF0e3C3R13KQfZ1WfV3nydCcHaaRAEUkYUQ
aZGJjnoXfzsuQoBujM4kPPFJ40g2qlrFjKINDaSEblB5+WayvY67blwrr4cYXSEZ
bTYLOYiGf95hZHONo/2csuhjzfsGEawWilCJx4fjpYdRcNOQbtpCv342EiHYnmjg
hATR8J9K96v0YUcnq9/LTXW+onXM3bBGxllqzWS936ocJC3RSrI+rZpmKub+44Ry
bLbnQM8g6z5nI2aourk/mewDo1leORMcyODWojnzCgzjuE4qqGTFIfSfNNATw2rq
d1IZvdBsVAYbi7NXRiJXfb3oIPZMsZhkvZXpQWNouTJrRNM5Y8s9meD/2OG3ki9P
RJ+enYmTWVe6lJwk11mbg9uTWPHQA6aNuIHKmNoYgLKZwU+r0zySH10XFI6/eIf+
woNmhcqVb3gP0d+oh1hQMh8VFT4f+jLuvrGfDnxDKLk0yKAFOQAFA1ixSRXdKFqn
J8H+hgIfIwB/VyOHXY1t/EuBz/euxcrpekC0N90GASJN7etZzfCO5nAW5u+GH/Ii
UMp+zxmDc/WP0KMhDRLtaXvZg3AedfcIQ3QbGW6y28EZACPl0CorDXOnpiz5i0W6
uFPquFvsitXPl80Z4BUrdKWGfwkvTqDdWigaTyO+HvYysOSs6l6MPmOyXfyHCqlm
6XV6M+jeSWkxZ8HLFohBIo9T7T1Ijc41PChRvbvAApzlW43hVJQwHOxsnG5XZh73
uquWFyOu6mO6vjy8nCrA8R0AIqRWTVfrgbvPX4Me8cekmJsxQ/HlCRIc2zwFom9F
x+Ko4mrskd4uUfmHMfMy0+ZswGBrCUO56eLn+qfqBN2/9QJtFG78GxwQTgtTQxB8
SyZRKSk285GQt0xaa2vHxOLv+8epvpM+GG1N2+sLAS1O5Ky1Qg4gMFKZOze0Pkxv
YN7W1/xMssj8DFkhWQkHRcgA+egfYn9AiOYlQb74HAAoPbDfWPUiAMd7g8mAaK9S
gq23CbnMOBRrDYg8bO/8EO26efvTzbNg8x/oY8NFWjEULHUjgEyrwEA6zTs4/wct
pFxcvDx2kKTuvFtp9Z7SA36P76Z1HGTV8mv21Cd6aaZl/mjNspHR5fu3bDqNbzVU
ytf/gccKQxjhhgAHuweZ8dCvq0KuLMhymIx+7wjg8+WK3ibxA7UYv5o6hjR2Y1uB
Ea3Shu5WlPohlQyqGvYS4WLYpokJVeL3DcSa3auV6lMF4NxrEpfzeTdEfxD+IRu+
9X9ZCtDkVzymjp5EZA6kjO4b83QNOrY+uWPJr0udeLAff8rLUwPwA752RSbYtRU1
vIqF0tn/vvCz7/VMLkk1HP4x05OdbDx6EfF7RUy7gTx31yzcHj8poUm0Kh/FH5jN
01DhcDnAAtAEYgkIjxyogPOokmj195E5iTgo5NARgxMzPgH97XlgT+UNCppPgY+N
QfeeIS0AZZRUarAflG+K8KcswQLJZtBaZDBZj0mrxf/XWwNoWqM4Y1nTb+vwfljT
Kwl7CH0lo+KGB3TL6v9yU5oB3r7S7EKtP5S9Dk8xWiXqH3SpS8j7J/9zeXWhJhA1
LWLVO5PqSRLluCuWgeixvzvt6XBmSvqRj9GIIVqAiMr0uL8MUttgHombpMj4TcV1
8vWyVa6Jo3q5wZAmTEvAT0u1QxIhS9Hpviyt89Fp97NgWJubO5zL5i/C2ah5Q8/A
Q2piA4pOcC2FzyWL/HzTjr3WJ1szMYKO4fh78AAl4iah2IhvhQFGgHjCNciw4rfk
UDJ1gFKdPPplkifvaIzfnXNx/Yn2LZQrZHpTQICxUt0G3xrQEL5xrwpyt8/GLIbR
Jcq+rqyrkmKYKTIEZi6uDiTTkOgdlEW43YQX4z/2aknSzL1jRPFRS4ZjOF69Zcjd
gPKy5+2RMPLS51QsJ2Itq1sq1nBFWi5d8UGui93dgZBSZ/s1VTkwiCx5C5iUbCgU
NTry3CF5wRB2hqApLyCfz48vQ6a0yOzwEv0grN8Nj/0GgUFoVnicfuNrozg3dJzg
ucv0GDTrhsvMxGbJjPF+me5qfF9Au8ro5jex29SZnHeVh9/YWvrDB6NRrKhlgB2e
ryPp2gjQjO+a4OZAqkFhypPEuq5wrl1+s0KyJfEmzc5rslCwRqmi9aeVlXWGG+uC
YZ28ECq2EiOAX4Fg/NHQYnzoQhmgyh6L/AjnrN8vfInaTha81I6ZII7fiJgJ/5dO
4GtS3mTjaojJ27Tn7x21qfYmeoHtXnMmXj8AqiDAZRGft9t+HfawU4ITLSYlfZxg
exF9t+bZDCWkhjv89RxhYuVvKWyu3/L69TRBfFYL1JhOsRSNU701W/Pny9O6i78J
+bwyUbHJNu5PC+IH1ysdxNFo7MLbCnmcJj9aJU/nCgc4kKcsBoyl/5I9I+RuuGXc
UCTfthyi2yko+dpswIrswyq0WR6lZwb3hetN4a5xwXqI/N/hib0SHBQZtCbZrNr8
qQwCOdOKQa1vPEbl3Pd7Hq/D+33WHBc3J8/I10BflFpXfra02E74or2EkfOutp28
mUdb0v+2t3vo1mCyslb1b4H8M+OYxEU9+X1JtMhvpHENTFkbC54GDpBxk1dAtBvz
h75x0QruaEBmO9GalmNI7maR9SwnraxnPfCO6e98CBYOolmJfeW1P98DH1wtgNei
zKq+fiq36S0vAf6jaJxGiYZ+RfEdTu1VVwqTTc1uU1GjilgQJBkISF35Xzuy8B6z
5PaLo8mWDcbzU0cna02zAWr4LqfcF70aiJM/+AsIjgGNb7dwLeMKRsen8uxElrWV
80ZpjA4n1fz6PcnTYpxv4yPzePS8a9NNrQIgFY2PGvt92zEWbSnCezeL9XpILWN3
v+jgld0KiTE/gY3Du797hyNpH5Z8YK1Fv4F2rUig+rVp5eC2wHMMD3s5PlYCzzkd
KdJoGI9CZ/f41J/IXn3il9utoegcP8/cOItuidvHyhtcjaO2sYlAQj7NOZMV/TCO
098C9owd84KCs8+5AoY1w2izNEgk/fIPIIqpMnUjSPy4rm2fcMjetymra3fbDjyD
4DebtmR3YA8C7bMLVopzA6SgtmMwZsAw1qcdI6hrbmxhxkL7bpe8l0RmzRNlAogO
0CvHlDlLAn+xyAMhjlePcDVcdts/7OnmCpY2ViKOElfb9PfV/htiPZneThKwGsfg
aegu5WOuPCSAToWNp1H5oR42s/27ncnkr8CtkRoNXGosHc+zUHQJsVE0cmIyydYf
WcxebNCSFyqg6v3KoRzCTX/YUfSjpGGLpNqNcYHyzi9GX2JUcBnneWaaVr2N2zvE
wsUUzlZ7mx0kmsyXJVEtLJX2gbpYQ7fgoXBCweTGDkNPsVqZ7v6L9a9177z734RW
T4w6mborennoeWMhjU6TVECKYqPVhlcF+V8mUWV0O8y3wTzv8Tu3lniMWVHJtZkm
M8hedQk/HJrxPYVeDdYv7Bd6KKDVYv1OC3pk+fxrUYt+lZS6gWz7XwrveQMuZ1wH
GMeP2m8JbTl87hrEhhGnxjXPELNRM1adcdtGhiAoFPyIi+a6jd/1HUt81xslLSry
D0Xlq00+lVPE3hRhAUa4MlVslvKoORc3XJd6SWQEDEvKf6xnOHwXApwp2LYNquop
/WAKjsg1kS7gIDQ4lI/rbzxela/R+1Bk2Xv7w2BVNpT0f+eIkX/WEH0kbMLjEHTk
WlzdYrU+G6aFadK7/UMr4YQWR5Y2CZX0QhBsJoYmRbRmi/pISf1cjnUmqRCrI2bP
ZHswmASRxLPuKJZYLWfs/YAg4vOIjdoQ+odz0Fq59CCFqM5uVuUryKGjtMqEjya2
gchhvF4qSnS3kPOO+q8drJKFUwl2BcknwxHQHWzoFs4RaakaEM2QXRs8283xcpd2
DNz7XL/4CAWoyqDJqwhw+2CGq7s0IKcNTLKGs5QNP8vlA1jqJHU1nXmF/eG8Vpff
qS0fSI6mJ0OkLOptYC4owiOBKCZU3e8j06NLTr2fln018eZe12Td40o9kG2c6M4o
l2n5Ij5q51IRxtRetAt9KQbh0uEsX+6lqe9MfXL+iZCYA9hVuB2g7hcgyFAtus1x
qf/L9AHu2fIdBhP9Kgc5Wfx30Sjrj0OxeUV4vyFL/08s1Rpi7/Akre6ilXUfYDcw
dLeiLc0PUwHNvNC7vm8C8GmSTG2kjCKHf6qqcLeOC24AeiQ45bCdOfiY0oIvm6Vi
OvmfaIw0FHemsZhiH8JchY5m/9F6RuERCiHnocK39BuBTgkg3Cuf62Nvs5QgZBib
VKTHKJKX4/ooNvmBU0ZAjfS5R5on1iaghFKLiM2m2UMMAJFH9VXEVLimANQ5qWHa
qi+T+kMz3dalDC4D0BL/LgkY4wXRRbdr5PXNWUaBMd1QPeyE4+bq0uO7Tj8DX9ay
elulech5kjF8O/NZ0PcXbrC7b2MiEqsmYFN81jV8ozfYPC9/U003mojhMpNUbMKE
n/GIDP3suiedPcFOkNSmmt6bYQxkZBPBYKcGx2RZyuLZsFbT9XtvBmYIlx+x8moz
4iBgHoeACnO8Bp/gls6k4fW9THRp/S/hhWUawWrXWWG0Fu2udYNXZ7+a96lIDgdn
Meldl9yibwbBzvmapR4Nr8YhBuRlLwzwp8S4eFB3CoLm8JddcxYLkRI3Lm+SzZs+
AlKZZxWw4UuyLqbZTG3s4qxUHhOJmyibSLLAuWoiLHXUL+lLmowUnL6xbGPB8BH7
8vw1F3hE1+rBUgOlgeudhZpgOmxq6YXSJPMXCsAmygL3rfO59XIWV/3aR8ti2KVw
xCYSyabgMHJmJ54nUhFLBaURVrCzVl6DW2N+OW9W/mPBHeK2hs5pMgvqphAfRyMX
LzFHVIJWZ2Pv1R+wMPwRkQP2Cyi0482IkKrluSQu4n208Q4zx0XO83MhnPcdAi3t
0IMOKp4HbYmw3xe1AU1hfy1+YjsD5h1cfNALH7gfEI+/cjygo5oCPsBPhl790SWe
FXs5pvoPjGdHkOkgrEbOarMHLptlv+gcrzkS9+U+lLBPdegLAnFjva8DVt37Nnpy
TEsXq8BQ8qr71akQG6SRKvqh/Pwr8kUa0gbFZ147FIIaQswlj+8KGeDF3tHw2zhU
JyR30pFjAodMzMWYCOirQhPf05mm145UGyBmpXfBPYK1I0OM8ux4a/nYlyqztiz9
5ppZsItpJVhZ2bzEh1UyFUo/mxuay2W56fbpT+SPuLs/i2BaPSJyzakrIzXWzD7x
2OdxmMNfk8mh1KWj606p3MITVEfHwFAu4MmLpgRDHdbDrcZKEFOvcW/zNaDFIRbc
WM1X2+yNBYGAIYruK7bwiEBR3ZqW2PBigua4Ml+6VxWBoxqC3e0AVQsRC+tFTA3J
m2OJeh+wXaL5IRn0qoiB5vpxMImR4pmfCGrQPK6v/QDqMJ+PhSQF3pS5jhdkpp8H
jx1IuO+9nSQlkkqYSML0UARzK7FjUoobskq9HJC7WhatRwarOwyf5VFiuwETlOjT
3NSwhr4IhxhiOwHp4Zo6J8RuBTjghhUshvLzd0nvMB9V7dHmnWQFHMFsit0EQoyB
aS8O9JjiuGOkisGwOurI48hj4+CJVfjq49i6ZYQzXDlFkDX2/T972UPup65V8EeH
A+q0W6mUQHn8Jg2e3pub1cGsk4C+CNqnL+KFiBkf7IvqPWDBkY5TOFtb3sbS/7g6
aDFFZE3eZ2YsW2TSmtN3+/RNquQ859ZQQTY+V8fzckAOSYYD+GH7QOzv1xVpoPCY
iQexDjspeO0W7TI2z58+YB2EZ0PcwOUotoDPFEP7QUZNnTj7Y0qOQVQMgMmiDYGF
i4MSn6LkEXynv3i0C589lGry4a634C4uFjWB8yxssZ8=
`protect END_PROTECTED
