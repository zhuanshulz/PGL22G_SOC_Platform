`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4zVXfCVWMHbFhvCDYUzEmOzPytbUopVyiTqVwUlWVDcbvT1Zuht1I5NvY+T5JWd3
/0XwEBdHkaTANIY7Yzbwp9+7IVKIzMxIM6pTl3t62fi8fljwmB2aBkCY3riFn7q2
aXwV7z11YLbaYt4EB03PnUasOX1TL7/W7cLrsLv1P8FOwU3mn4w6rEm4ltRFgM+V
P2n9Roe9QIJsk6xRbiFx0UQ9Q37HcfFdgOBlQI2VGlsK4MsvisOcTOiwIMjvS1yK
gH57jbe+dstkJJm8ndM0EngCkZxfYXp4sAdfafB003z9XgwXIbwZO4/ubFcudvh6
y+68EKfEQRaHB55Zj6IH3o7N0pcyuZRcmq5QkBlNJg+CLf1YyBMIReYeueBrNAhQ
NQ0C2dTPkBo7CjcVnaCqPA==
`protect END_PROTECTED
