`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V4I5JNmREwpOHG/HTlSSLun/+ZCYm0psJfrkycCdeS6spMcEqox5yOMHyORMoVjK
g3OmOz52SoYluiIW1VX7iqORXoeSymxYrgio3B5vbvkd3SgIC8y4f0FSSTuq9+CR
7wZbW4oZkd/YDi1EYgoZf+/fDVGkF7h2jxAwNq97mDETCvHj7UmxuHq24LN6ZPmW
H5zVcIw77n/hNQ5tPsVf3fYcBPNhcIcBnEDYnReFdOdovzrkBDgU3tcYrVB0+nLc
52D9SvImUOT5eEwF+jIDGNHNkFRUqSnFI63wj6VE0PDMFoNSUfkzL6n9aCPZniw8
3l4LxUeGa5f76F5xivdRRZc+/kOkRIYhJZQAWAX3p5hQ6gM9Obra9G9JblpBDj06
q9e0GWqgQ6lC72AnYR1nXg==
`protect END_PROTECTED
