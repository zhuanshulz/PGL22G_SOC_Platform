`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xFMgTahKWgfar/EdmXLLXJ6Y1t0pM/hAzUy0LGjgroXYNaWTcVxaQQvEOVydPJ8w
nZMYMmkGf+jW18zFq3KD4i4O/1k0QcfP6P0EOsBhwOAzIne2uVcyJu6evdmZDRWR
PnwiCsMM0oRr2ypimNd1+gnijIZjdgDj4pny5eZ3kEti4G4W/S4/UzhzxJRcJh+w
EzhalI/yt5kXhxCoh+G2zZN3+u3Xcp0uiXN1HyAGeRD6FYeaSRFTvVTBZcNQjUnG
3Q6cPc6v+x9kFozTD/MtFzhuVatbUm0LBRQ2byavJzlZ5RH6wOq//YmpiFVYwMmz
DJUv8jFaUfFHq6W/9Swqf+vvPv9mkLGqPh8GQyVftoChXWo909Bmqt1mhqfU/XZi
jFv8Iy/f4Yh/EeoAFtOYg1yxvz2XqBzvJQ3lhWrS5AQDMQBNoQF22KwpmBdkbaB1
/w+SKB+iEzrrROWy+q9A8wTmhH8u2x1CgK3/nlvrQ+owxxh6XYLKZypx4xWZQadL
0sJAZ8A1M2joGkbZiG7LnjZZ0NZTW7bwmBwnXdz7r5P3pmiEAXCGnSW7WhbGGrEx
Po1AZQ/fui5tEzvUDh0tTJ8BEFbwM9+vg4f/2ot++O/boB6Bglg2vA2YO9pk/WXo
2b3QNMghBB1Hdt2nsKQLN4i4FWrafKiduYCaVOSZ9S3+g4TMkiXMB0/D+ITu0/pG
IcDdz+TOjjWaHpBBvc4vDhBWlaZkBXaei1AhBwd9YLrrZZ2id697iCWF6prSiTNZ
ODC3Q8oSZ9hGc+8xZhtPblsBa7jFprg1IVtwx+6X9IXEiJLcNqmDWD/JN5Vjh27z
s2VLHxVf+fEDcxe0DNjjwIGrkrsLFAdrk8FuJW5noVmseHoxQxfTUvD48fqIiZJA
QH5OgNtub/YeKi8qMbwCmw==
`protect END_PROTECTED
