`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhFyOtUtyUC6EUT1ndlJyujkmapuU2ulGMYdSo9bQlfDGBSwAGOawfOEco1FHUZc
MTQWJp3E4MnPSo6SW+D/L/C2lAnqP5JwRCxYXbD0c093tQxPFL7a1bUDtH3ZQsAW
g2ww2VAgl22cAbRaKkI8k7KceHuTEviW7kMNqP/lbvpGQVj9ni+0G/ZG2t9uvH99
5zuvF/6qGY3J2CBRmI+OWaLUX1Qy1bhxC6xQ+SH4ZoHOAzdIai3rgAztJxx8JS2i
rmb/3j53h+Jj7brkq9TNj7LJOnZO0f0BmNlvLPV4Ob8ihYrqZvTg3PWG7CVhDFlQ
bFkLXPaohsVt41ehobWT1XOwOzQVmHgH8WUEsp/8Qf841qf8k1mc0O1f3r8vRtbF
F3aex8Xc2l+Fwa7rjKyMX8wxh/3ap4ponR36gpqNnkPEZo/xzPbpdTJ83VQZrHfs
6SIY8cYD93s4zZkZHZVHdVpMxi/1iHKI6e6va3BBto2HyUU92+FLkLHSHfhoN2W0
pTxmPWq/migweNAAJMAHiEd1cjUINHT0JHmA8k8QaL5DA0UhRuduhgS2N2Ar77q7
7Q0tyAmq0pxUIxyJK8AJsDs5YPJpvupNhlQqzaxuNznZuZj/w4zXdiGV17ExnhmD
OPjL9ThyL9yTk38JTqbQAZI/NKqCK5WQPV4NrL98rSJ4a7OeVLo99Q3V8ProhGb5
cy/7CHlKP6QXVOxn5O2hCKjt7pKx5PcRiXZ6y12YMPkkKte83s9y44HdTt1pM+jv
Mn+GLYdvtDixQ/voQA/6m6h3eTpQXAac/d+0vHSnVkxzk9fWj7viZE8MOpzG9LnY
`protect END_PROTECTED
