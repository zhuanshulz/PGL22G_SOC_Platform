`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GhJCLWjKDZ5cYzfPbkwLULtJfDRnFUbWkzwzfFnwxNXztPUIE+Mlypq88myE/h/Q
31bPRxIqM8emnDdYtDhn/HVFHrLQxU660xsth47Fvvprb2/GdCs+LnSf3vor4bLy
iLrHC1C2oV/CM79tEZlgEte79kvKPsmiCy7eqPBUPOs574agITVAAEpudqzBmf5I
KUiq2QR6HwuYE3E6dRJFgs0bqPK7k74FUgCG9u38CHGpKoyuu5Lc04RGBXkqGLMb
p+jWUjMNGRvBXMZ9E44cZssmQS4M7mC5iWhnwuPDLlIWTUrSSp55iYFX70rPla0u
CFcjt9I934S1qlqEM5ykbuClGC5eyxyr+UxXkHopJAx3MaC7vepkfcxkEIR7ODiI
O+c1GfrNqEADFfyDCZkUNfqsaHP4UESRY/I44MJ7dKBIKudq0t+SPWPykt9m028B
qjZ5jg5jpBxjg07r5c50Y5OfyRr80RpcLUvSOxM3xHcefhOqx+YJ6420pTray69l
TDa4g59SRAmSXcw/hBGEgh1Ui0LJANXJc3BIEVstVlIVJ7efeWUyRC18jJe4TrkM
3hkC0oTY0M1pW1eHmYgbbUBFDBzeDbdRbTxnxVzbQicaZKKSNOk6avCJg5AX18Y5
iNMS6eT8sWdwoAqR87i6ZnSr0RuVzU4fLcUgsJOmwZ6HMOmw3pK+UXrzwWjMftDW
wx4SM8nD5mxAJHdSfPWAb6oCvlDSty9rLF1e2lP0qYFNbHxeM2FSd/eeBuJiRP1M
NyhNvaI9cg8zQv9o8zwh0XK3aVOlJL5OEk5QW5x3Q5oBajt5WBwU4i+bcBx6doeY
61KvHdt9Ik/Y/iUBbmsDEax1AeNYvXyY633UT0jcJy3usIkHMdjZAmKA4TUSa7tO
`protect END_PROTECTED
