`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBISAk5f/XItvhS3Q3/G18QgQkBUoI7cN7AoObmFWjXPL1Ymq0WEz4bc2vkmmMSw
W9EGCjw0Zb/sWZI9tvjEqe2a8gURGmc6Z4aPFqvfOmxPE4vcMMrmJlgo4DXwdZTy
ivCPfKvFVV+JugKLycuoYvwbzIq8ERW5VKnx6bUGix6Ps9kr63dPNT8+GQnfl/hT
JBfPIbhg67cRlFG8co6Dsh4V9XGFB43VeYZV4b9ksv9PE/8nxRFpJ8sweL1ZNdCz
cmIhqz+aFZ1gwbxXAXxwcTD0HgZwjJqHyNeUZOq0ybjgrEYbux+1H55Dh4s++cWF
dEklACBPnvoJsZjMJiFWxsi3EGZwROi/aOajCPR3Tq3/IuzIOOvMnuy4IbG4HQUd
`protect END_PROTECTED
