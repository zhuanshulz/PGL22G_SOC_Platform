`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85dRmbXTRKwhcqv62yIE3TbUieHw3Ch3nmqcOp+rgXsxc26XzsDxjrtmscnqh+8y
C2a0WLK2XX/a9riTSWm7Go/ljcrt2X1mJ45oD9b4ew0nDDyUc+bs6mjmvrbfHyIV
l1S3aRoqbFDZfpci1kinl853XDVyJE6G0uCJKpw0JU/B1q4FKIBQna/ZoFUZZbS8
rV5EuiE+TeqP7sOeohnAmoaRIrk5KVlpguSDz0MTpxNLZMJW9N+K0wIN5weuF8eQ
MZqVfKs3S7QQCufAyWVDCU5jV7iMn/NhqjRJwEAk3gR8vh0aGqAOlZI5dmxGWF7V
/qWbYLND561XPuwEscT2VXzRbUK12nClcGxKE4d9AMtJN0rtrRw+8DycWjYznNWl
dQ3thkWe5Y4KqgkwDbdk4EVsiO2BWN4FXBUxPnzCMRU=
`protect END_PROTECTED
