`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m+qZtYdf0gUhV/sHI6ksNZsdn1vaiCH4JmZ/VjjO5GP4oBLIWu93CoQsqw1GDp6K
4lRnzP2pmONcAKkWYYb4nwfATJ/2clVOHhMoAohiQaj+LvmMHJdRglUFEbH3P8mC
OFqqHIr8ah4w1iFUsXSe/48BzF+DTIw2MrvG3zgykOdS7Vi3Fb073y99ZYZMNVZA
cvlTHOZ7PA818WwJ4b+MHBU7cK5m+8a8KrrK7X1XrZfHKr7cpE4tbYfLQATzN8X3
j0EM2WMq671RVwSy0pvgobSKV55gbWcPuwng3Vom23J6oZOyCKii/7juG0LDW/tn
ebuQCO8dDPXnMYVx6dfqnQE+QuEdaIDfTc4ZZu42djoC8oqKOnq/cdBxGtmRSS/U
yWzJbBAY9smiI5h4GbwZ6xfbb+4oRDT9vcPgYdFr0RyFfW9mJa5O+vDasnDVC9uT
oloCp6kvvWpKLRe2vPgQOvio0cuF9RQEwRPBi0Fvv66KQgzrIj6bnGbCqWkvahXB
+PwCIjIDpWs1/a6hR+Jeh6Qtmbf8roQ6vHj5mTV9S8zTvyhJpSiZhDGPu9DBMRpB
YUG/0Q4rx5Xr69bXJ/YvIG4JeHOzvOoav9bHd9U6YC4=
`protect END_PROTECTED
