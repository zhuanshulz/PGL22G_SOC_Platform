`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J5OHIJQA+m9edO3E/+Pdbf071S+uSUN4lMbVW7dm7AVuzL/pyI7H5CdvGKqaLPQz
ZnrmOdTecGldaWMrXh84iAoi5Tq1GCug+vdBk372Ffh6OVxgXARWim0qMESuNsUG
KZ4Kl8VeP16ZAqU/HIbrKj0D+WRxgPqOtZWE2L1ZLHIKIWWFbanRZ2lbx9rs5SBZ
qcYdqBJhFI2kKB6wtwBAn8PXzMrsidRSs5n7onjzBma+Bv6gtrjstkdvzoMKwNUg
QPbFUJecFvVzecaMKfIku8cY/XR3hPp6wJaKlPBUNX7tBrTMpK35bNOy2jfA+YuT
1mn2P6XNDmL4n0PWjy8pqy6kZHJa/sIO+AcC0s9yuTsSJmbAsC0kSDWe9JztjhxB
j66nBMTWzV2ja0uGG3Jk0hmeogmBY46rg4P+wPioK66YyfW2z0nfF8p7W8Tr0KmG
h/HxI8sGwfK5eglpZ3TX63bTLQiPsp90Scc/vh2tliVJnMPX8HvOLSRNlCxox1Hm
+b9FK9DFjSDKzgHAo2ccK/Sc8wYoMrmBRsI/YfNuPP/4gw1biDNXicrWo1oNlVl6
Kr9cGEyGHplGE5DWUq4iKEiR73YMv5U5706R7Hs08Vkh2t1dNKkX9kMJVEx6Aw3F
8Xvwz0eJjOA+3LXJhoFODFCR7ZBWBXkUjnH5SEhkYbdYz0sJPT2/zydxMDftdNos
FzcZikKctJ93ch1dMTDU4t6A+8wxgKFyNCsh8zNuX0pfJcL/SdfPFOATvo3KK/xH
S2JLLW8uPmT+34tFq6MAYviektfYxemGw4wTv9A/S3zquRQScelaFsbJzFMpiKkk
qXW7WfJclwMb4TeGzhHVDdb1RfHKqvjJKoMERL38iMJ8B9ZaVdXhFzc6+tLRglit
IyLElCt+RfV4e+x6hsr5COuvezNOTV0+j1YhJA6C1Sol/nOCnUf9Lkzryw6DC6R0
qwBAihi4N/ANQNocUmkWtiBifLoiazAMpg315CMV3yabBZpOCDYp8lrP2K8lgVCo
rh7T5j4IKw/Rlwx9ps/DWbLgwY/yFyGKOyaIeQXFR5tiAfYjdpmSIisNb7wtG6zF
IEZgh14CqqpPNp2/FDRJaTKtu1BGEbFk2xgEPjJUu+2jTdlFdeq3TAARq8k3w6zE
0ErhFAySxAABTMDpEEjC0KtlyJ/J4Vw2aAeWvtGBKwnY5N5g4LLpBPp8PAMQxjeI
XumGLsfT4OJ9AnsfN9KI0lab0a3GbRIVZ6/GVtAX0YqdmvFXZ6f5SeXez24aQxfu
T1L7c0NYh6nNY1iD+c5FwtQhRltpOzIKYicXkoMPr+rzzuDpgI+Cm36c+UNqUjrL
RcVkcOTLQv1L6O9nQtNKdaEsmKjjH+BKY80lngW3/sRYbgqO/nagWXI1nfqbmHN3
SBd48EtdBUA+baVRxwMhaMX2GLlhR4WDGnC1T0E8YqonAgHozGzwdFZ/S1NIxk5T
otm39+fe/ns1flLhfVsvmiNZXnhkESCSbIFadYJ81DTk2W1wztFgd2CDKPCnfx5r
b0OFJJNoe71fS9XhyF20ukWVa2QJlsh3wfSUmpwRt+HE2WW2GNmk3sncsBpRq2wJ
ZkVRL4YJGGY+ImNlfbkESOoLRuVhyK6Ev6UzMVS9SX+QOnrLc35D0047L6mlV98J
5Okw4Y9AhTnbz3goyenzvW+HVDJ/UVVxt6fOzvXZ4gcp+33Qj7GbWD1G1Dz7ygj7
8RaUOFLegc+bmzhvcERhDuXtB7TTHbDzWCX+9VGRHJXQtsaYmlXzLEC/Hwbp6miB
ub8oHZ4pEzyWmowWDzzWOgM044RfrGwvKRpoOdctUxLNKUFunBFC7Y3mSQd8KdRQ
Ub0CmlvXqu5n6TW5TAbktpcphFAt5qPXW8MpqSMg5GZ2YvNdHFOhonqkFDIRuqK0
cYbFyY3l5lhDNsXfZ4mo70BTRGkFu5NOMgyvxNegCJWh+ZOyPjXw92JR+dBaFmy7
V0HIoN1rRUMscsAYb34moMph968z4CLP7Fpzi306+ibU0dim7rgQApa+fg1Q/Rwr
SY5E+LbjJiMPgXRWKEhAQhz26txpsTcBDrYXAQ7KZFvGzkeuw1yUn4LsLM9/m1xk
S9A0D7r34OER9meL+cqjRX1ujfLOWmbH0y5JZYZnsWM9NZ5sCFzeueTB+0bOMJlH
LHCMmN+h/uol0fApLNfokztXAFf/uIZ4wp6xZZaxM5zRtVAxazCo2q+gFJuI6s5m
q9FOMrNHeDxWr7P4MP4IRGjniS8uDbdlzwulobceJl4=
`protect END_PROTECTED
