`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QhIC8Ifc6n6QKlFbTK1cJKs+9Qp2sdWFmnhDMEJepq1NhxGq88flpTnmuSVAUSJz
QJSsqGT+3a3TczPyHeyhwLymvmw9+dFfBAS9JrTJIa3aHaJZVGEKzKYo2YqK1MnS
u+YWeUtu+4r3sIQd/7bgBK0km6BS6hMHBVhJbX4NGcU7Se3az0eY1CiWRZA5qh/6
u9GrD1whCa+iyA2BB6kCCAe2hdo/XbDF/2CqFP2WlkxubWE0RcvuqDD7CK/MJOzm
tK9MB71GiNt2c6T/ySirS+0Hr/FJl6zJg09BX3/eDa7O2ATjYsZYMLYPzVHR3egX
o6nrnN59UXlh8C1MiGyo43PH9av+liDBAERIGwA/0AEDYdIYE0YBEUeiWPOBa3qQ
X8Jf62795hwoSLjNcZxRgia64bRZip1KC5u+PNSl32kRUnmihdHko8phOL12ptDr
tbDe5VBNk17YCMJPu98u3E9UXyq3Kt2GgPHAI0PgIrPwWgsmxhmgA/M2QmfY04qt
lqLbVOz5vCdse74LwH2PFTGE3qWccl4gTSf1T6kT0aQmXli0BsyDEB6EXtJxQpPn
fySRvRDyplvrlmLolp/8xhQwjbn9OS9GYyFA7Df1B+OMSWyvJSWWeZ7kkoBAlFqo
ZXNdJG9aRhpnGOVnvqfS2muea9dWqwq5YDf0ajnv5U0nslVlxp7CGtC9K3+ZRxRh
2xOQSttp0CaRQ06jmYYUab/J8nzrgUfVdYUowAXbM5Lt64Xa8ag6FZSjenHURF+v
+fid8SBY9vh9G7lslgqPh9RESFP5rrFCAP3220Pt8PFYJq7JaARJxz0yYOtBUPaC
FHpmmFNJgNkNwOFyIXEGwC89FdQkAXE0z/ZhFUXzTNujDkJKuCOWIo+ZtvQ+Q4as
zJ7N/cV+XebaV5LzmJxpeRSKY1lDTQ1oVwlyBb9hh5gqtCG4ayS801O+pur1xQSY
eSCEQ+zP4/FYU3Of+iagO4juK553oiKSrFvcGWLAMxw=
`protect END_PROTECTED
