`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33uGa0/nGB2Meqn4xEeXGuQSsQMfv8MNnpUdGiJZUbtcs73nNT8jVzWD8Wh/JkvP
IrO992m3F2+gO1Y0361Z6ShoIOm2niOKxyofgfYPozZK3HEJlfSBsqkvbRb5p1Dm
r22DK/pvsZzsaAB5yYx7u3ApXu9YirX4bqdk2iRjXjChrWCFe2OZNCsiLxadwiW8
fl+CwudXmKQT3A9UqK3ovqm8nvz53uRC7paHbuG7oNAyhz3Tt+MrQ3+AAGkMHPXx
ftq5P1HyWo/KT/1dmKN8/UZy9j7LdChisWIYzI9iHhoI0/6hsDLQmwGBUDR2xJee
Y8+iV8m1i4xgCOiajUqfPQeeTVYfPP+mv/WNsm39/UgEskeV2v20Zkf1uH8gJyh1
ruAiWWKjceFKHAAJbxkrGi0lnCQNIwWT5mUkGJQzkrbkiwvI01KwZxGuw40+74kT
PXfeT0+sXtGBNDDF8iRJDuilNdK4VP7hHvdPtIL8KzACFo7mCyMes6N2xRI5/AN2
5BqULx/qQ2S7zgfTcpcdzw96CGM74hWZiyw2/OVd1wkXVc7Sb6VlPGECZB+LYL44
o8vdPCRlDnFN+U8mCOXaIqhDCl6d9GHKYwOOdaASStBwMWHDBVes2ypFuE15TMM2
cacfNb1DiUHwZV3G54feQM6XXTYaz4lRONmPdIigC5wgsFhWtuAR7HGv5bbnQp6Y
Jot+s+j+YQfYG6rumfbu7gkB2+7INtnpEEzvbCZbkYw=
`protect END_PROTECTED
