`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTxzv5qwyu4xouVI6BrAX+XvbmwWAiqbeYV81AvyXSS0M9W6NpKwg4M778Mw0+W/
Qtzp1/zjBy7dVZu6K5f6r/f+J7gG1xXE0augKaANCHUDZJDbZ0x2cuE+uI7vZjXJ
aFXvJ9ypC9lqayd4SmCX72bnnhmL8oP1woelhHMCyN3uR86mrOwKjtz8RXaRHLKY
mpM/SXjioQO0HyiivNpbkaLEbuMOUPKRKq1mgDeTxMJbeo6vc7fAfqP7W5USX/WD
9yCQYaOnnm76LE0ki2ZQ4fgRKZOGbaZP/n856uAK2ftqyTQM8tx42gyUyYWbqpiu
tGuiIIBhvEikG4NmuIMtG8tHut/PUaC7rDzosVDIkEtaZvPgRrT1u5mXAynJAYMH
fALH4uII3fyBUFSVCgyT1e9dlYhnuNMpxKu9chwnIi1r8OH7ob4i9hIs631VATHy
iZAamICbU+tsYKDl/wt5JBJnaAE7kybkfwvkPoox1Pl9S8tYBIt67/+3QUbJ0WHs
ofPOmA66h4maC5ctM/lIXV03GH8PVObdpWn7zEYS4wZbe5q1BEyIM4ZE0QYJ8zLT
qwaiaLpr6x+oQntdS9dP1HVeXMIb/zVwot79oFzLF2R3ccGqg8IplJeE195gZD3N
mq/bp/UVYjfSu7pRsdZDMwm7vnpvmgPgVpaxUCDnFbTBGqdrn4rFf844BTp6R4YO
OIA+eU5wZOEEN8VUtUeA7PQpT08/BwsAZm+dZoUl0bpiJtu6pL7dnwjTTujGK6GV
MMfOMidETXhXYwAcWqUVCZX8NXlPYHy9t5xLSwesS1ZbRRg+dX2LVLieyDpXDa4i
4fqCuOvdE427ss9KT696U7uLb/8OaE/KTbkJoQvX6yxkhcwOahOVEFUNGTuDNZ8U
KrEF3/CXiMf65Z67MXJPbT/esFuLZsgSW2+v30qCdi3ByunJhX/YFWS8OqRMvFCz
ibgAN4SZaei3drJvFZp2Q7U59QfCMiVA87mkjnkI+WMCFxmFhXK7os7nSn96pKuN
RpZJQpBpG86kpa5p+92vvRdeSYf+YOGtVZ+nkLLC8iQc45hfH2cm20J3S19a1v4l
y5MiaHeK2gExXDAvD/8Hp7mGnwd3l6tkzF+tp7ppUDBwqV8wKFTekNgarS3es+xh
1AH0QfFGvx12X4i4xpDplg==
`protect END_PROTECTED
