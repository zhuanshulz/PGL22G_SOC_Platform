`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDB7cmnMLXwAEEZRW9tRy5W4Zvh0PtdX+Hp+R0OXPwQjCQcp5evzdIcl5+aHprEu
gugw8OI/BTiB4pNzGLvgFRL3YtnsUNMW3LalrcejyWNrNc8Il8Q5Aeii8Rd24qN9
OueEcsZp01GEko7Q7gHjRMRlO9kLMpWvXu99JIW9mI48Pzi+OuzZYnaEM4wLcz9L
cqBzWRRe2pr4loPiwDXkQIEQokGRfAX12y0QYmqc/1wv1ZcbdgdAxhFiwkHD+DXz
`protect END_PROTECTED
