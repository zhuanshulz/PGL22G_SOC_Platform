`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xo73GoAiNc86Tc2F02bYv/pHOqVQ88XbWfEjPXhn2RikvYrt9fDuu7C5Ut1skf1g
zyF/J7mnNdInt6VJ84QCj/HUtKAL6LB7OoOIeSOTzXuwKoMvz7BUgKf/iSYEH0CY
Uz2AnpAlnVew5EKwZObps7iSMD+7RvgTvPkd3N34e2V9vEf0jNfT9eEVBBgLYZTf
S2Q4vbZsd2NGA4kjSrLfj1ybUB524OKxoS9bcZVjSwXLXloFAfj5ALYujib1hBY6
QxcQ2lyc1QUUbNVkzJD+ZOev/m8BlhKhmtWkFUYrp/maw7vu7yRAiEyH8hZsy/gs
fAEAFTgU0jiS2ogufYS08Pf/4xzJ5HyYBfKUAuYnnph8KDTmhXgjIV0zIyG55wZc
1ASvXskNRmljrJVjDz5VNPqSkcaB59wK7yQpo91oPSPAxSTYzuZbNrjlTgVhWOaE
X8enwUcDBR+od/hsVm1jtipoqxX6jO5cff3Y5fWvMkDBsFJiCzeZdiVJMA2wH42/
gzUuFJRGFstEGOgeK2lPdc/qfOUzZ6s6Yk2J+cImyvQIeUb1vfQpkNfSt3ZsNEUJ
6OZ42sX2o94dmCSKDDuZGlttuaNzEHkcxl+vHBomJsHhq4dXsWAhsuDcF8gaPaZn
58vt09LvHVg5wyaXz97TE0EKqdCupuOKyETHS6hDNJrD0RJ+jO2EtnHEOZhvM69P
0xlQ4y0pf4Vp7oABzFu4iLicshroOzX1b29Ny7zNy+KyslqNKAKRZ66h0OAONn6k
/QJLRe1eehTbkFyX4fhNbeQFBJ/zVQLFQ1YfkTQ3GiS9/K5P5ytTM+97tZddrWBk
cPXf9eRax/dH1R4pODx09M0jMGKpEjByv1pz6OZ71itpZ2r0wsSH0eFyNtpVIwM9
5y6Y7tSjMTLfB2zCTaRlkqjDY/P3g4DIGBVbua0tpFT9Jah+37L/TA3KuYu7ZSoJ
Y/fLQV3hnmBHn0fCm2IpwDiTojx/Qfs7deUcqZ9dKgFdR407Fy9HV1LHzoi92ECB
W6JcrRnTgQJH0tbuLWtBWi6debwyIAiS+Fc+/xYDKV0p2siAWzxE64kqJFBzMdBl
lVbrgssYlFAeEy+4sstqoJXy09lt/J20RGObUW7/krqmXhOLPRQ527BNQw9diKHp
8frIcBEjqmkblt5WRvodzepetT8GoD/WGZLEDo98R0o0+437n2SAiFrpXEP2mBg7
Sm8SAzelvM3Kvqc8VS2zmHt4qR3UH7ykovhbB1sN4GDdmSQ11HcuYszTC2JH82k/
zKI+jp0COMqbI9sG7eJA7Thb1yktr9Q8gjG/HjvAB9WFYS5xH8E1IYpPb5bgPSTa
nyhR6CM2l4qZ+T8diHqawRqC8B5JoRv0VXa+6JlBBKsAdF7XbupAlZ4sUdbbapA5
5mzAVYFUvwUOVPtymywHwNN24Vb/H8p7DbfXL0sO/PeNKmgcFfcVorwtwbeTrygX
h5/o+ahA2PtTsr9IvLzyr4XD0M6oQRSTy8iyZuLyiWJI/T5LcyKHQqu6qKlj0Hs6
Yg4gTs39gwTkBWCe3/ZMnnBPz2obCAyowuGvIsdbeBIZ98rTWbVc1uNBPffeCZAM
kNNucafYMCHWpOD0sif1vcjtLZk0w3KcZQe+IRXn8Ojclkc/bnacddhlxgjslMen
2z4BZ7rlrqQdePe0lhHf6UW7n/ikvUxk7h/GyonBu2lWVzfAIH6bv8jI8NDie2e1
aFqej61MNxQ3Hx+RT2RmxrpGRBEskK44GzP8unSYIDvw4o+gFTPIAV9VyUR+eleu
T9tmDugtvkRXp+h4tnJcqz0rywnSrBwsYxu7cHDlRQ2Osf+xLtwvlhk1VUqybqH2
Yi27tUBpnQ9H7YkOqymalWuc+t0u8MZ/VhJRlfSW9o4nB23QAaRjpFTWtCOU3J0f
ECWGbJsyWe/qvv2XxSf1k9fi2fhMMVNpoLzUtcIRCeaoj1aeQxxriTfhH6t/a7zg
JIHCUym5LO17saEQ3yyLLWHlxBAT4018LTlfclZGrKQKVTqcZU1eGdS2scEhGHPb
wLZXwTFHiYVDiVOcpMixRM4hegWb8cDFBQSXWT5JHZuTQrI0ecVjeeJIPoGErEm0
eEZI9haMM/8uG4q3B1Ybhjj/Wo7GXp3rNjpfhUcki5eUjbWYirot3ZunM3ya1uOL
xG7op6lrdyciMDjvcpA4pkIzWIMWFQGhyVbWEc1dowqoTKBCrNvv3221h9j7NSfp
NJtFKqMntKK2BIk6RF1tGqhAE2lrSXx3iWsCiFrLSke6daIXVwGEfTrcLFFhsUKp
JDEfOaYApSFjVbYiXH5YzdPBs25BskLDROEI+XuYSNZKhugS35QAKwOoJRr7YsfP
AiEBJEI9YI7/YE+6TJj5gIg2/A3Os4y5waUpUmDFQNYgs5QrPcwQo+3oYl8pelCS
vR04sFA5iCi8Iixf3et/GhEW7SlQH88UnSf+x1j6QduL69lrBHVYRYT7N7L6Thmx
efvQrDOuPCuKQqHiyuGSlUFmzc0qK68NLokhMq6Iqn8+S8QQh1i3clNiy5o3hOm0
MUSi3JgOsNfelu0Dc4tCY7RzIkCTlCneXhFgXGNUiK0fZ9OZEOSV9uvB/DqlERwu
RtllYcmeDQs2wO4gzUCM0o87bS9TIutBeahcDEAUoOpGkvPbjRPB4QW3yrjFKOOo
UCUtlZvkmAN2RB+VRb87H/myvE92nbJiBr4gjOngvUkzzlqA79v/KwPvhPI+ikf4
T7J0y7HANrRncHSlDq03EFgzkBdx4B5ebVjsUJWnH7ngX+alMNyyPS7AAOsXYAep
b7dN1vXbhiefTixSxy0nNasiuBaTFV80+dMhPrMwv0v2iJNzzPT7+ASvdqTBrY/C
HGbsYO77OCi0wxoGGBFWkGCCSe42liVee5TIB4gix8vWch9vaoXg6VXWrvFYqDEq
ywPtSMccndiToPmpkwF8lpbWTFCVcmKq8mOiPLCwdiOwW2RhmpTq97Z0S97AxS1C
j8BouNlFE2hvZgPgwA3DqlPpheIeVTxPnP6ICLbhcvtUDdzhWJhUrFWZ0DTxLOOY
8MSMqDF+Qzqq8NE39BkBl9yPKXn+258QggmRYrkgKlQp6Wp13BLplA8+H21CFsJU
uTQZuLY9ZLinOznjTSKHjAzqRSvGgeKe2yfASuPXaCXA8/l+GwscKpwBQ7GeK21e
+gVV0crPUeMQu06otprhqAmrizPkhcCzajq8qS7hBSD73TTVwe6W6mA3UmI5kmrB
dbYVn1sZrH0fslodrGg9PwPnjsBX85V1ojtvysjeXtJqiZyShDe8NCfavQOvklYh
SH6dFCmpSg0G5lnKXDGB1vxV/qJZs/AwzK16F/0gJurncbCkj5Fx3+NQkNpji7BU
eEAz9OvS0+pivzs7KgU8yC41Iay7J99zcLVQXgP93hJzsL6W26qO4KjkQOvi5ItL
3Ou4oWV6D4SkJj3YCtDw+gNsHpreb90yerM44qIc1G6uom+gp7DgZZBcoprgsZ76
4rrHmdArYIMpqj6dbE4x27RBhqohZcG8fB1yLAoOVqCo/9CKpVW4/0AnMf/oaGmn
GMf7WeR31S10J7ZwXp/Ttr/0xR9cxwH2pkgXVPtJKweEqT2vO0bXQ5yrBbxA9UM9
srEbjYwxpnAvPHxpt6bbNM7Q+ZtTe5jPcdMohoy2VyCSVPJ/Z4qBATXlz4e8Hze2
8xLF9aBxxUo2YJTLMh6wxDarNTCVnQSbZPRU/K/9Utmfzs8EAW8aYxU/bUG4cUoz
q1rROYPt0GIVp+Q33yRu41yjlJufj6LW9QRgYHGMZGmvIBVn6QWcOEp4Ch/hYYU2
rbq5psm4i+VlhKhkJvPkM+9R7VJzCReSoWkoR3DZj0n7/HfzE7O/gmighPh3tQK8
jCUqO5GIexKCvmrHx07WMJqW8CaktMM5kC62/fdJljKjOaFOttePM3w6DFu+SNNd
rLZL1etEqiPdh87NCdBpWA==
`protect END_PROTECTED
