`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5d9oha2kJRcpbBl4OAjyz+PzmHkbfkLmCWxitVOiVuJpfk0pHMehYpbFyC4DgGgU
E9y6zcVCYx72kxdafurXN3QLb0WodKAl1FO9b9S8CnM9e6qV4vkf3LikuQCTCp4A
qhvl1eAk2rU+txfYNOEtKW7v0wNjF2eaMe5OaRUyWElgVUdMCNH3KWndZN0Fg2VR
CSNkNqTWO0GIdTGqXSvO348Ewrj7g5qobHm9yEaWqNp5ZzJi7IpxtDaUxNgEV4WP
+C0jste9SON9WXt2aZv3ywcgu/I784WRxNKDvEfAZiKy7fRp456E3diWn4D0wS7t
HVxV6LZsl5Q7hAUc1mf9CscV+ihO+Z2noSi1hH/V64mwmMNJXNU1umlOX3/sAwcL
npJJhtvphZkMTrVMwaLVNQRJV5wnyv4bJnnGR2bkz8xOCTizSnNRNWQQ5lJFMOAU
rY/4zE96KOLYUhcnu0x5QDQFReaRhtJq5PEpB0z9laQldb7mkH4IJFCj+Osb+Aap
E/YPZXls57r5KrGps7paOG4MYRFI/iSCwGKyGvmNBpsMNYh1kMmxjH8fQThW/IFe
+SMr6EnOGR6bUJcHtGhHP+flvh1tQ7JfyexvGUZenRb+WqHLFddTFOTX3jW3VDQr
1CwQy/zDrfvx97YvjkalBmPDY1Gpod2PpIbyZCtYzv063iBAJRUDVA+wPtu0edjh
oMjfgLHCFh03EwQaLQGqGP/9sKh4oelVQ+BY8ZhUaISLpreB0y7axkys26SVoDJo
ixZwt9+2mMhpBprI5PUJQsTe1hLfEPmYKE0HJjiWzx945a4DNbzzkH9+YQ2IHRWr
bdc18OjnM8okZ722N1mY8w==
`protect END_PROTECTED
