`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N3x26OeFBDH61XJaKwl0wSQgO9l/me4hvEOupbQNf3F7x7vnZpUJxs3TLgchnjAv
r6/baYsQypnW5kkkC/aeZjG6HkCHQY6H7CmdLMYhQX0MCS5VsGejmFFeNy+Rs+79
K7RISuDMcYYB/Mz4lWu1sp2t8/mpCb0btF9TJj3ukwB7L4x47hE7SA4xx8xpjBAQ
4ua8mhFf12ilB/iLYY0ekCz9YMB3YOXbDGRIYF1Jcjhf+7RO1/YcsZQNPJh9z9+p
j+cI6lItl471LMZrj35HbWcFbDJbYF9/N4Alca/Uy3Iav9UCDgfTfOtO9XMrOspd
cb3xO+Myqif1ojXpYQa8syrawPxwZqMbuGYYCza/TNNTMZD7LbozLoDwZrN+q+YX
ICNjl4k0RxRv/v6Ba+fdw/d11bjVYgXkep4KzJwWwpZcsJgrfUgLuyx7rKT+OP8L
XUOdzoFCwRcnGIIqb9WwMAQKDWw8abjkRph6mVhn/v7/4RD2KTXHoGxx+XC1g8NQ
m916Q89550ZHxTM9dlIKgknWc4HLR4vKTCAF3N6OiJz0dcYyhghxWLmHUiQ0Aaae
WmIHoQ0Y1a3cocy12+Q9Ug==
`protect END_PROTECTED
