`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EwgkoNmvr/NtZcdoR/pjYe/33Zjs4vZvQPeoZebXgoinQeP3dWC7oWUabt2cDJnJ
MuglufN0z7SQbarVkJcaSvNnheHyxqTSbJV2MHthu2kCANWh6CIMtm2/AEX7Ey2d
oQ1YA8VxNuQtRy8orv5iVLLSzt4rcgM6YUpW2O+RszjR1IsupsdtuU7O58iWZ4PD
BuYmh1dB+nHkwMz/XItmciOHBHn/LiK3qrFHbkUxAfzpjENArvQ0X4r9neeOV7mq
oimdIvNvgf0fJtc06tM9R1n8274lpNqUPcMtPCQg+kPT/nyr2MoDRaZPbPomVm4f
YMxk6oXUiGporORLzqPdw+ntZ0oWA+/BbnGGwqu6wMUNiCpWLiikMhh7ekI6xmOD
F2p1HYkXjxuJJHSKECpilIh2B/nZhFbb4BkIuAuhwqYr/L6FtINMcciU0onGWDMt
I3vOibhlhJw7DpxNsqCpUl5OK+SHh28G1fq/SkYO2tyNtkdztPEc1viLxBd4LsZz
47oKojw25zUiOTa0P20rz3nJ79buSnJIEBlfv8vppXSe/+JwbnhrU2mP2p2LUbjl
afFFF1kkN1+hipkTF2wlRWe8UdIY3av4TjKVH7WyhOq+ixK7JXz3Q6pEhsP1oj+D
ViXbq1Km1RRtM9mNlNPihhwgHmU89VjCu6Mp5VHEOjgMpYn3WLqwV34iz9/LKXKG
LVImCxZA5mI3G7BiQOdPENTZBJ4aKOvXxcLqV/FVcf1HQ04BMgPgRiELIKa7diwV
W4clISQhTOIyhU4sgPDRKJ2IhvGaqjTl0fRq04tCGHQ0FlGlgcX4sfkbILWioZK5
IXYJseBK7O1fFI7ZxnVMXYGrHKcN7QlLyxvXc2qsCAZY/qZy3USnUUCYW3xPVbrs
gj3fVmnLAWQZY35oprqH5PapH9e3kIMo9utAnszKikhCrFy0YE74gh8YNV0UCML1
tzJpIaO2HSI4xhSd+I17AbDDoWxANUFaNvOE7cBDxLWRzdY/NFSxQGkw3DKeNoFo
WIZq5iG3EgsRp91CHf7wixVVF9yxHcqSNJzRR7jTx6ZNFURP2d5p6MWY3bsbf3n7
ihTgEtVkw88ClRzM/gVbSHKias7IPT+cKIjuguKzenJPi/uGgHAH5eWoG373SfSc
82nJufFIJ5CWmGgF0qKqxfUxQpyswLmDLmZQYy6LC8UBIVVT7udUUbzFefcF4q7R
7+0WhKp3VHSubAPHHwMJiMlSRBblQXQA9aRI7AHhoHIpFmz7uDfRj04JZLvbHhA1
OZCRPP1/kHgLwJIDqjoy8JiGJB7DOWq4vtp4O/ahtoy1HlFPXMXHLbJkjoB6bloq
/H9XWN8s4kJyQFryp2rHCM6H/WxszdLdJuc6XSWoeT7b9sQrOeZmml3ArJwOHUKc
dkDjdRxSk0pf1r3nuAeSolpXSYOBkpGOxNhP2TYL73rTp5rnoVAofCzYEkNrYu4H
i+ennTvhAKwdPz9qihE0q/+jS2hAHViIgXlF3Qs8mQvniYYkDiQ2wPnvJf9w9PcY
x/cCYeWPrLWM+8kny7OSbZKyh0LXBQWFrZPHXSrtQee0xk026tfWC/yNp2qVSuuI
txm3YOvC/XzC8FhFXi2mVXIPzzF/dpabSmutWXHE2TfZVdGRCqUh3c9OCkHKSqX2
GlZS4LbDpZ+Ch/7S2eCk8jv1ej5d82HIwaM10QABDp16mZkeFOWvOYQ6hxY65tP+
3LIfx3Ajv8cIuVwNtvCIO4Rl7QRPp9oWb/4muSPM6s2YGEWgzZSSj6w+P/SDvs+X
7PJpTYlRdUt9cmKS46YWCAsVIaJcbtFriUbDU0QIhuwRj+wsfMDXlVWZ3vcxaOHU
IVCZdcaPj+5jUh1Pslc1OdOsSGC/EVw8muUq9BFeYqzE16qQschdM/+OV766/WHe
ZkrX9AMQa564LUfbOPBhZg3Y1oVeidH3xoAinEPuFWMX042wA3sn14CWZTKUcr0A
bYgYQeSbvuiVDPiuKru48b1yxka646nYcqqIT+ArjhBGZV7cSNM8RH55MzGYCoaC
JZut8uAiA6c4MAmABNkMsi0+7gaWGolpZCpUuc/sSvV43iY/H927Fjs0a0GdAIiu
1mH+ifB47xv0Q9mOJSgjxEYMmFwGq9rS2XKBy64zqTQ5hGo3xbuhB38wUqMFg/RW
PCXHw01dpAHN23w6CTaR8VuMrnnzKnn/jw+e82Z+SUcQsqXJGoyuFy38r5pZo1Le
Ea6vuh0UbYwmbk8J7Bzm8f08JSqr8EP9+vr+DB70tjONPYKWb++NKh/ChPZP8QPo
gTkocraUwmhkWB2yDDDcm1aiqnqsVd4rBqh5nKNUT3yJVsNSBYnb2HkmAWlwVh7T
KionZfbrbQWoN9WjEIYcdlx/bYw11vxxQPPzUgKGEnXguNiXQQS9+tFKQ3pUJufj
c9UmouZlul2UiqlXKs45A3tglM+dP1Qu48WJfWRRGZjodj9PIW9JRNCP7OJV5PpS
+LANvFLge39/i6GfUmVx0mY9sWpGxEiOeW9Xqh1tKRNu+Z6yhXfMogaem4mTaBfP
S8AqAIlRO5+qW7CxhcEDHQr1ROymk3B63NdwmtyDuZLzz4WN0V3cJW5+inuZkYvS
/AwKTtPGsistPQsLd7BDPAqPQVwfCVt9TTbtYQnAC2fdAyHlNVrQEUdnn79ZVeyy
4GX49iVEh9J7qVXQb484zmxvhs8ufxy/IWcKEeWCX5WcOFMxz3AMxwYUQuSt+GtU
XGPx3mGEuj0nGoL/d7vVEiz92zrfbXUpyjWFOQ+10wfH2TH4T7Cvjpfu++b+6a9Q
G7xcPcvCAEH4NEsYOwWOlnWZPNP2vpHX9qeXIs+aXVdimdbJx+Wg7tZTCybE99BV
g0M7RSNyo1deVZXAyLeOrs0aLJrRm3Ogydu/Fl8y/AgGlS2xCPIBU7+oQa4p+Acp
/ZeOXkppevrgZV8A5WztEql4YyUIKASFx4oGGU3pbrbysuIFwePI1xtY/3ZGFw2M
mpxQSr9h15NEUF+sGlhTR2BRp7lWYWC/j4KG8aMCvze0UKzWLfHUSqAMUj/6L96u
WydYH1vMNeE7dEaP+lWpbUcu+/Yf8L5K+EoFaChwEA67e9rVNUSrek3vwxcowViY
oA0SHCbM64OG2HOv/Naf7iB3ZPz0pQeC/qtGp7xHGSbYfPCy876DCSs4I6oljGdE
RKRF2HPg8qZeaGFrBIwNFtVfDAwPFynx6CVs5QcE/Te4bz0UVq/hGJVJ3980VZcW
nK1D1UgXtQlXThlJRA1gJU6CW40/hpElbr3htmejC0rqRvT63Slc32URSTbhhXAx
9w71fMdqbLo+hansQ2JHPHtW0k+8n4SP82LrVaHtU81iquiFk+XFzfyG4jmAyHQC
2xctDPSSuz4c1yK/HUrQfruea/kvD/AyaCJXD27MV2KmhvZLBpx2VY1nVtjhm8jd
KtjShQRaDNMfohnY8/5HAGDCupz+sQLQYSdJel1xnjV/5d1t60L0r5zJbb9rujIq
L34juQa5n+4OnRHjilMZvBlDJA2zMAN9nxgp7FTc+oob3lSgRxw1kzVGBJd39FBU
dUgUqEDNaToFzSgSJtpYFYelxKde6pp/9iI3OzWV7/tZWlAZJktLXTFZyhQG4cb8
Y2q2svPrTcDXK/58wN3hABypRzcYLoOTR0ujVgHB4LXyWAZuKHxRWvA7n84dHisW
tnVKXrHGLTD0pH0RduR9WyRn3QwK6uz4XShNV/IhAgXntTbc1hGd2SW7uwzv44xh
aU40dAIsTJfoF7CUkNIZWZf1r6l05csI7tB/olfVkfmQTL8JfgaVgAeQ19JBirNb
aqiVgPLDv3/P0zu6rTsIfbS2RK3hQ0PnZYGtM4pgEjMn4dv5/freY3P3vU088xkH
ISrHo8LrIAIc9TQHQ9EQJcFAW+BXO6n7rc1CNhHnl2WEajgHeVboziHOuNIlA8X3
/tATbQqmcG87cGBwa1+UUEYlENrZgiFRvDRhDZAflvo0ruNV65JlJH59kRmHqedF
+l4pOVAPPAig/4q7VuIBEuut8T0nPif/lpWlc7g9wTN3Vi+Y/UIQK37YC7QC4qOV
uCu9KNkkEl0K+AnZibvNyl7mbARt6W0VTlVeEklwlWudHYnNRvbjkNEj9ACzwE4R
EAlwLp16MHU8d9imnPIeP9bJdQ8PRCLNTHw+acHS29x+/JahFYs127vWHh1o/S6a
tj/TUYBe2P3/4IoC6YXVWj+SbNjXnnGnIpfKgn8GHKFi8H96KRPUlthMoeZjVEXn
LP9/2sNtUCYtpVmqt+PX4c3iJz8ywkbzt8pumuwJZiIVCEs75PRL3oflbOuHr5en
KlmvIGMEtSeeBEDd2DO3sL0hsrDNMR1rGOcVGIkS2CFZ71Ph5cb4rHgPCAjaguy2
YHJcOSpf3E7cQ3muE41HewBQV48btoj1M4Q484W7fMGAwJcQMnv1rxRiX9fsQBQ9
0+E2CGJXK+F8HXNkGOmHR10HCVHMfrQlTwg1ByiNSaNemtUX/BpbaTN+VoKRLuBX
O9Od5G+CJ47d6ODdi66nr9RbtUC5i4iw0EKiXrgXYqDwl35Cjygv+gNseHDYGEuT
sJVyD2//fPjtftxQH8zERAsCNpO7jn9hWP2xvhgazxVgf52kOWqMaaUY0yE2T7D7
jGCs7ps1KtMX4KzE+uxewetwt0IQEiMCucou3uG+qd7GzSbH4uCkLwyi7BR3JK72
qSMvK0u2uBDtSd/etnm5LUjPPHE7AFG1xuUCBGzvXVhJRxg27b09+wXVP52Gs76G
5AGSXUNS8oEp/lNOkx1L5iF7VNffYS/b1x3DnVYCLj6h37eBPLK1O2hIs/huD0fB
8FDNEZZsOSFqKMRcb3DGATdLpPLU22yPisj6VxxvN8u3TymfgSsB5BjL7YCzvivT
gHVVERcnYiW5MmtRFlYCYOhjWaCxCy/GYAltetuHb9zl2HZZAGAM3pVRLGGYdz9w
le2eMdh0lCUaY3XtB1OBXR2ptEWNxVbe6O7zp2rLlJBjqKj+IcC1kL0xzbKRVa8k
oX3WaFaa7/sgQpxiO7Kghfx8cqiXBMGsrMC4bj/SKW4bp5m+AS611PMGqyYnKT4b
IOspiv0J7D5LBMHMob6YzPh8K0InqZwqKYxLO0yAqrt2jRpbbj/bLvYmsQnihSbV
tDblsLsiLHodTetu9J1+OzJQzlUqqCY7fNlT+T3bC2OvtgPupvP/NzPpTkFKD+cH
Ahv9mZEa0DslK8ngt5097UHwvGnpJxbzPaZGsl2ClZJRCcjzofCaS0jCeov4KmkC
IOY9ZnqMXIQB2gsxe0PcXOwH3VRKBQxYCLig5d3ZrS+E0vFcant2sna/mO8tnCfN
HI4g1Z3ZYvz7K2r9oOOgcKRIF+P4PDAvUZGx0A47T9EV1vH+/h3FomeikpN3JJ3l
pZuq9va7167P1V8LI40q+d1gDZKkdyWdGFPsXOE343spqddYugEk7G5MfMHStu5U
ogfn1QRF5rzt//fcNO3Jt4frfCRa9Fm6+M6x1foQvh5aqwGV1USI6YQLPuDCsLfJ
wj4cquroS5Kn9bP5ZSrD7dGHzmhuGGqL8gTZ6X+SBp6Rw7O0VElsP9W/rr7lUmjV
sFw65DqBATveHz+8OMmSpjJTTZ48WltVFqZNRL1Q1ho7eeq7eIBR1cbsGEXQ7yzJ
37hD/wPJatCRdohhKuail0xV7VhUsiVD8YPPHLMSVRwF/a0HcTwQEmQFKx5YouuQ
vp0GVhT36XhupaGlEYvkXNKVgOiwHkjDriG+qMet6y2yEYhWqMkeZaQ5IOWWtcUJ
y7ygygRUq5Jg5t+SdSeWlJpmGtNsePFSzQh+IRfBapqjxQ+c4eaB3wnXfj9zkVku
TAGRhQCNXOpM/YdwGQ4NOIAIFanAKGzR6ijbw5Cm+9W8QqPU5KnpWgppGZdd0NF8
2c1Y8FA8QgDdKItF5badVdgY82H7CST3E1X9wNpvtriC7Mco97guDkX5eWS8wOgW
TboG5Yq0LghltQms6CaJ7jpGPmhDNL8CBkHJq1Pnzye0OzDiyNBMoCgHn5QYpqIh
zuJk0sQhL8ALQR9hc4QdPRKsGa19B6DmuPGVy5UDrgAsOq5iEbPeOz3bH95pm1bc
pPKM26SD0+UmUDjZBQ+syQUgD5UAbh1lZpYNzoAxv27JRrj2BKpPtqClcJfvaAnT
YflqSaHy/ldI6BfWzbA0VyvyJBfDcoWvjDsRHLvI32X/hBKKpYlRo4bXSS3mc+ON
TFdViFrbolCaca8/3YGl8zOvDt0HlsDV4yoWqcuNoJyyxvkPoGkyoVInhCOTDFWV
Odc7Irp7YvHuOMitb09zbnJqFvCSkipVVsJWjbRkIEoKVbPqzLPcN6B/O+hX2nJE
cKGAdgw4RiTjUWaEhXojxke6bBDPhibg4c9/m0Vjpru/iSurzPc+3Jvi1hSxgBbu
Le/zxltOEK0hzoMdSePfDqtW0t+/5toU1jyo+DCsGKVkMqcXrwvg2dAR1QDMI4nW
HGEJs7X56n5agpXELYCNHy5BM5K+iZMDBvLpY4d2SakM0/L1yNWMtKE8PmTfbZIx
JPp9T4JkBzxwLoOQ0kRc1uSX8pmbY7vRauhJxqvAcOJ+V0DyoMBXdRcRMZYQFvRH
ovDiLdwK2O8SvhXlh5Uqgsf9kmyE/jwaRXhjW8fEUovMEBwCauZURi2yY+LzJP/0
Nv0f5RBW5yWgw/5+F8kxNRqsLndhZ53/9NmySleAl5+PlszapyJYorFyik2qBsra
9JMY6IZV8osRaFNCXh2ikAJmJIUdxpDPwzLn2FXXjq2mAFlf2H2hvP0APT2fHhro
IbceKaiLpYG4l3nXcQ199kiP3UIsmOkoXCnT5BpFucQitpVBvC+6rXUWlkNXK0wH
owfv7pk9iSN1jPBtzD9kywgaJENfPOrZ+CqcQrkXnUCkUrzz7ublOisPdC3ojuK/
kosKFBZfFEmEFWZ7drXuRE074mWsydU17CHTVAak5NwTJxAQWjTlHkgZnQpcKQFw
TR+L+Sv49uR3VekmwWE1Upl2DH482a5DUSp+nR9R52eHfr5g2QciO29qDGvX/4ej
Re0Rwj3iRAg7RpJy0efx7FDZ81Xhxvo/Fy/rHCi/8gtwoHtpg4s1NdH9Y9weUnUb
+BB4kmMJS9IvgH4T+Q7dWoo/7Cg6ifssr6oo+Ev2wuxteSLJaT0XUiNprURsbo6t
+C1o4WJvLD9eZKeYYcJL23zGCerhFQx0Kxz7nQY9FUARun33LgE1yfX8IdxaFE9w
8GUnXYYAYrwOwL9g0m9bjeOe1P1Olw5HFxXiXFr8Q7uZmDr2VlqdjqQSJzE6RaON
FJkB4SD2ZvqIxJd2i17ih17Q/xdcvGi43+UMXqsEo2W8jjpf8RFayqfWB1q/MRUg
uwEZWMTm0AkbtEX2OZGeoylr40wM2bbDVz8T8yFMqNCqjuWgVp7SOqXEVMBYF+uD
aRZw00WChjq0dk9lGbrRnwJBC3txaOgICSVtDGVHt81vQN401HViHKiAtUueMYur
YNYZAIEeTLC2lmta0kEpfhLcaI3+8/kaCmUvIAYA1PkxX41aGwsbU7dE56Vkc+cv
goqJxZgUFoACcUSkpUapL3ObmUFMQ19gacMC8dP3FCKuuSQrvTESc1RfwA+I6uGb
QbnfwqUvkogJwCvW2gWvXun8pYcGQfGfoLaMYJmP7MOAhwbVcFh8oWTu+a4lMH2C
QupZ/1EPglMcT/qbTbYalmUN18kk4QJAf+Fjpq/qxC+XnaBYcPkf2BoBhhblv3ir
g2w/IhtFtDEjHyC2nGNxhn96kI5gfFeLqk3vbitXOHdvyS0bo0+Txym1oWPoDJGf
VJPOT1EQxJdLZjP1szqMqYiUewtmPk1SyeUVAszDXFNrlcKLk7yhFbKFPrbn+4qI
02uh14aHH+4LR8JrwrYl5DlPv1M9bvq2rXWnJlJxyniG9iIA0wZNkTvnH1GUsdFe
zOkLqJXTqrEqpenzEf4BlWEQIsPQMvEl6uD9tuyIdZO2bVcZCVOV2gx5PrEV6Bwx
cvyZElvOUH/yULLDBvvnSgc0B9a8LZ06pWswwJBvOTnDSZAI7Yb7dFXirb9rEYXb
w4+r7nzvFrvUdcfccVjTJeQb9q348Ceu+MgqGf/rgekWKofaIV4pQHMExScZk/3W
88nZaS7I89+fKi2KsNmcA2bQhxJLEN13xU1Fj5SAQqB31J6vSpqOpMnvsmlXl7mH
MNq4rpenS5iwl9VxfjUS0oG1yGDut3bjoMj1fm/vrNzpwKGKNBlQmJJKbBy8Oh2I
MNB72LoAPj9SKgx5o9wlTJDHj1EJadbWy01AvV4jHLv2GPpiAKue7mfS6KTbCAlN
97ZQG4SHlj0JjlKh0VIqqkyKR+Z0XYNy/iUl6vEM0fY+XB07bW8V+N7/6q+6C0yB
u219uAi2WYyXI80n8aVjYyAOJ9teGF8Wlamoz0M024Ilq9V2fRaWu8XUVz9GJJq6
tGKmXjRwj3F3w6vDpdmaAYhwT62QR6cxyFs3V3KHD6D27YM4I556bxDXY5tEJtFY
3bRJzGnYQxGTlnzL0y6GyY6G24PmtYUyG1UmrtYbTDj2N4o/kQRa1zWBTgSivz44
8LJj/gsICy2hl1K01QjSdP5fkaf+TDwHtQ9PLP1Z9hm8WTVwBPu0IB0r2VcYWEdG
Q+23K/qpEwxFs98y2YB7zfVg53+HK4VTTVSnEBM87YWLwTjcCTStGTr6cr//ffq+
gS/TcUDra0OmRWVY11AXPx5ja7Jrx33aTVXjfQzTyD0mYepUJrKTUQ+5fhAFfIBA
RiFzW/JvPCqk1IP0jXqT2SZyOGu6tWB5qweHnMez7zjYIdm4HG/EwQd9K9bU48eW
vtl7w/5vGBjF1FAspwRo/Kllsk9vAaQTvpbmkK1pJPjt2TKbb7JPfqIzKnbwyKaS
MYN2/cMCynCd6RN01tQ3PqF7pFlbPmEG7jceZuLJ4rvkI5r4dUSYd+LPnUnb9e5N
oER94v4eT7i6r8Tz94/F3D8hJ5CTSgo4U3JHPwzouyzPlPNwQfg57UInGw/G99Qm
FsKE/lp1889Krcjpo69mtzgqYGkyooN5rIzzrR/YKuGJBs+gBdgaj2/kmt6LaXhm
NJb6TxVNqfAgdEl72KVMeByKRfMMKUbl2wryRWBCPgvLxBJ8uC+ABzoWEUVCSJnl
NVtAW55UZOmBtHbypBSxApBOImkhezV/QMz90U3HRrcnICtAMFl4QN5ykRIsfdzB
Yv39a7y4Ph3x3SdSMsNGh3QdvoQi5AgViy1mSyoySt5jQKmdB46S+I0cuivTp0i3
KSp0OuOtlvPGhQzeoylt4Wijxmx3UJkQdmMvA8W1GNyOUMdeu/8Z80ldMxGqbkb7
6kFpPbM4cQhsTcM6TZs5Hh2b9AuIsAT4Tom+6kSZ6hWG1gAFXkS2Nj29F3pGRadx
dmHxK24behkRcwjTC84MSD8pE8jxxw7etKXJPXSCZ0SQFX5zUKd8brdrd+SrfEPs
L6zyDkFaQz873biBRj9it8pjRG9IxEPTWbHZOdfZvJkE51ihJX/uTuodGiC9W4jO
bEUGjrAHMthrxnlM3rTlgagLqHEiT+9qb56id/CK6fr6DSjfc3wKq/iDhZse4DXU
zGoOoeO1R2AjaIhqMQG+7VfPVWzJr2luYFHcTw0rwOCPhVLEioKD7eKzW+EbH+dl
rE0uXW5A2JotNSwf/DlWc4rCvrpUtUnLkoz+oOaT1EhBhTzoeb358ClrGMX8zIX1
w9ia2+neCBpSK2Bv9ilvPZF5KitsyeQ88zm7IQg/d9Uvsi70fqp1++STfvzahQ6X
Gcf2pbEGeive5aK/mXH1RtZAF38S20xkQaIhpbAHweu4Ce6LkTiDPcuLZlfG+1V7
yOODycmw3xEtprzolBufdX4d02MBbXZtebMwnOpKQ9aHNf9XRp4dJ25nE/+6dP+s
y8iVIxoJxfELNR2qv4RK2zEgVYraLrzoWqOuH6yVYB0Gj4p1H8Zbj5+2+TER1TOv
UAnY+FHCMrMPnTIuUnLgeX6TX+1RfJHFFTUndeayEQTkr8/gRgGJpoPTCauQGgYw
btyFLpXe+XERgU9393dtxLv5YxoB4DS30pWEE5A4zr47H3mia7i3d8rf9i6qvRPQ
MavX2EUwn9leO8DWpseOZbS6ez8+hH7sxVz0HadpM6lO5lQRNNLvmU4ba7FdqJlI
1MBApwbgXV+9QnuKsgUai8dbJFbvE9etUesrxafnFpKtU2KFupkXj4JhYZpLe06n
ccc+tIWGAifTJ4bn8ETpgO2JcxQxJwKYqFa8RsZXAKvmI6xt5e1RTR+O1x8IPzLp
gRt7daZkNHGnCjsyOxoNFjNJqCVH/VTp/R0XWUjxiwhcYYwvolnNZZ8aO8iZQhSk
T72Ay65t7clc4B+xOMcVRbPDcXn5ILxxtC0DDa6XP5t+h5xO3ZslKGNskDrwZlNs
Ld8ALab/U+tD4hl8Hb2Rp2lW3txO6WwEMlGSOUDpClbNhD6ibeUjSmKSaK7ozHur
msArAwZ3f/AzgsuLaK78prMnJzB0QnttJ9QFpurrv3MbJPdAxk+QMnF3FskBHG+J
LY6sl/2+MJGv22eantMUkLuk4oolZVaDbpWq49EiB3hIw0h+RUo0BCPykNxzxRSN
95cefgVzM31MNS5vf2dK8hv2Niq/7LMg+0XhJZPCsKqSdR+l1V0OPqpamAKdek5f
AILKrfIYqh8IunN3D7T4U497y41pwHqFlDm8FJOV8co9QEiqIK/CyZmDP/0Z6QDT
8bUsDTR5u20vC6/4iALfpOVk2SC95ginfo/aKp7DJIEt97euLsZ61anD8Zmzv+u6
luIQSK+OPkBXkA8ZH/+XYzjfXx04ANr1rIR8ljNQRa/4WbDMs6T0+sYYAtqnfLkI
9VXIIM1XDBk9P8krj4XEfSsEy+NzjIIm2Rlr3hR42zrSBGbGJ/XISZQUi6gScela
YE9DACuZdyNFa6p1maOBl1phsgrI5FEjcJf75DoXwEIUBP4fVoYa6aG7WVvXRVKz
7Tq6h3fP0QmKwg9oPmpcjEf2HnW/GiyBS/JRZlea4GtFSSYkWmu4pQ7t80gCPP7U
VKKavBmikTm4f9mnVTtemuayknSYWXu5ULalwckHAJO3pr5i7VEi2yTuOJjU8ePQ
V6le1hLu/mkqOdP7z8Mskn9QckKBDYpIxr1ikmeNQJwzhYTFfCkW6YNEnC2gxXR/
apTEvS6MYoyzwBiGo+u12dIxMKsrw7KlVJLp5/aQ0Pwb+sp+3MU+ytPv2Wu347i7
2STXkbQtINrTS54tjg0nEv7OdiALOfWMlAIMfhPeeQ0aXiMUz5G/coNyIdJOmGz/
eBvsl2fJ7huakenYeSmxWhewigsA4kwpE3vx5FJyBiBVXCG96ylEnzhX4o9r5riL
aeLKvVaj16knqwAr3TNJz1AOQQuL2x0fm3GPFof3pyWZ0Z7FCaMkAtnaRFjAoU+b
3Wr6whc/RQDjxTcTh4kcH0qGdpWjJh9L7gwx3RWfrj83PCwcUhsECqhuIxQH3IQ2
XPaLBDFqnRvJkRAfCSJJKVhCeKL1LToVOnIGjrBvyNjvFxNqtarneY7pfqPWhXCh
HnbfMuXDNb4NqYx6+KLl+TO+imJia8kTt9J+EcudiAvDnlWVHRf0W7cIn3gOLgs8
VKx4jvKGHMgdG6HrR/f9spifX4DNqqFO6hipOmIHi/uOkq8NifCqiDlf1rItF3Of
gxGCgcuoCktbqHPXYPYMGGu2eHNztr1UXRQi2r5VBLvDozGGLrzygaFljU9bW7xm
S9pKc+tctFDSW5DLI8WTQajxDvr1nHVDb07+T5A+fhayQpiaFOnGQ03S1bvVYekB
urfcBZaOL9vO2GYJuXLyxnGDJqm6wMTJAK69+MvHe3PfKqvHm3LEQIMb5He0Sufw
4XfpjzEn2WE6P2RNlUAxeHStlVtitCHJmEWdClYlF0D245folk/ngWjEYPe7XxR+
Ca3fQ+nmdl5l/4c35Gy5CGDrbuFh88UVssb/vdqENrSk77gRVCHak/gQHJj1rBj7
xkWC0bDgKNCciR3qYH7bdw17jYZIdgzmiJDCtr2JI3y9hwcP7ZldmSASUwLecOHj
UqNXDafu8UO1rK0MILp4qe2hw0ML/rcNwliGaLbul5nYubM/F2bXk5UVR8EDcqUk
iPu8VjkzjWW5UMwEGWRrQJC0siBkyIV7GQTU5AX/KaEd9zL93/sUbHBgv7XtC9b6
M/WjRf0+SHb4LXN8zK0vo524xgJvOnWmV/iHcYEZD8JwE+0bAbDHzUNWYPDSSYUv
Jfiyh6E32DB0N6my8mv5jJBn+xiD1izF7Koaw9MtFBafouBV8UVqQ9lwobxX5/su
cnZ8k6eol74No2JbBhioEL35k5NWdFQbwAFUgEOCEq3LYJkIoxEi6hA9unFUBIT8
np5pqt86b/8FVZ0LXYySuMkHjfHZJizjQyIayl3qjpH40Y3GxfETXY1cqIWzCaLH
1ONR5FEub/kQ6O7c+jG0vPzy4orFSPQPKmIQ16LT/eApsvFpJE/knrK3LmQ5rb0T
BfdY80rPJg9ZNG7iii5I+HszAwQvlcNwyBOtR/ERqon1VDV+AIfcuOcmg587DTf0
hGyH/XcR4vYKcBcgUYYgZ6OESZILGkfONz412fJDqlCdeTagYF7V7QzT6IB++HW/
xjZkegoIYBAaw7fsVbh6TBhHzDvmEE7j1yqhHTrgqz7SCdGaIUqGuLQyHsglt0x4
B5HjI0eyY2xZfSCTv8fzPefHAPEBFA6xiPOkB2e0rIT4C1NzjfRIG+HVmYqF57ZH
jBAZLL9YeSBbDdEa1KlOAidkzuVPxFl1zHQ2OXahrvLNScqlDFDi1wyvtFJkf7jR
gbXiGxyzGudyO/4NaCBYAGeMVd+zNQ8sV3tmZ70QOQHbvJCcf1SpC/VRu2phwW+9
koM6ifBtPIWTOqgQeDDkUAnDOlmgDTZ2pRnwc0gnKbasF4YcpB7tMPH3ZGMRqlbU
/6vT3kuqQ1MplqveVGET0plsoHW1NVZDT3C6w/zF2bwcq0FUjAJRG7RNK318vQP5
W2PG+Eld9ckQDBNoSr4XM+5RWplEg0Q4B4x68CLIH7F/Y7MPVObekEyLiOordvXY
HLD8jmA8Ek0my6kSESeM6mVEwzJml/LvWVvtMznnnJumEIXoDCzRdzdB6olO/sHc
xA3TsgR/0viSMYAf1qhEU6hbmYO+Tl4AIyeaNLvKZ0Rdqk37vo8kbvM26hTd/BBU
HuaA8xEWRX7ELevD0Obdi8r2rCgX+hAG1QDH90VxH+xmbecNGDOfcTSEIzDa9IgJ
biXkA9Y/Aqcbb9CV2Q9vengamaZl3B0+S+yM68kX+opCUVtkgL5EgqwZGojDQRnu
PfBEEhaHE+9El1xUD1vun7iyXPNsyUOc6CTotM9yjCQVtaPBJ1N/CBhB/v4F0uxA
PsnjRGs7R5k2W1O1BD143tt+EcBBZBmssxdm9qBrwVpbss8MDIkif6atU1pTwwyY
XzXQD3MQnkwHKbjiI9UzVtWsGpBQwEK2nT1ihSkcsYQTp8mcZDIatLzeNDVaokN9
UtXh8tfhX5GTmNqL7WAdXqUlLahqKiWrRjKATSZqjqRnNFNksYO92iB61Ge8+XYe
EtVXLDL/+zwXSvE8hsb0qlGnIkET1TAD2r7sLrr5V3cQ4Imop+3DKCfSV0ycF9CF
HUw4eHwURUQXDJEIhWe2XfT+ER5LVpYOBBTEdtfl3S48kvMbaDaxrJtVXaF6EqVo
tgT6u2CbWyEZj66pB1WY6LWPOmPcID19VbkhkcAKO5W0kACRKoImcxjo1oVVmJNc
9mUAZmTA6gElRpkNrd480CYb0qK75so2LshQG0vW9q1SHWrmjXQH3wG/LQPJICgG
kQtWshBKLM6XEt17jP7dE+IRxnFudcpGxtb4unBwdGTkGLZ5Bz25Ze36jzndkT7a
gBREv2DTQuVCX0zBqB2vK4sOwKUh1sMTxQ8F1SQ2GhT4FTepOgZvkATtP3OwtmXt
js11cvVjMt9YnEfY2ysFTkq2st1BscKDnj1jeLzey7PsNAB/qfjweWw8vObRbjJr
k0vj2UQKpljBCAWj6iNd48OEKiIGbgoOjzJQGC9g9WI38C3Lyt/hnmYU6hI98a2t
qSxwhU9cd6MZjkTDcL0yA+Hhusry8hXEYoQs30Tebdfsg/M7Nmuj7Gm9VXBMgaTa
GiiLj8X0AHQy6AHuq6kDb+rnG42vXZSHiC+Keej2La3hbUVFsyvjBCeepcTM9sjD
X0BQqkykPb87ZwvWxVCD4bvYh6yDgYypab15FuxznHXXtQefvPo+FGeLatQulU9C
+z7BUfZAXwLT/DY3v8OrHuwyym59073Pw7Al8GSSk1bypP7G9JXWUqFPR0Ecopap
4ZDgUtueytRpSwOqy6Y+CnSlulbuBB3gmXy6KKrGHkC1FRk+QkV0bLMj8L/mp6T2
63TSJEDMV+Fy+rLgrr+JItOJKtki5XJsrHUD/ILyAc5MRFZFIdUWXpYvR2XK9yzS
/WnM6vBp19sXtnhIcgWQJV+HzI3qbVSOVfr7X2gIYWhuQmhaQaUWZkgGQjqawx1+
yjIQJ2DDqe/WZA+AdfnSJYmkUd+pLCsd9AlJ/gSkRdiVog4idGTCw+sHRnYpD31e
lRQbnizNCZHgZZjiv+ij3Itd1rLwgRm9jlw1w0B3lDUfliL/rPlWVMhPqy46WHSX
F1O3nGAIXhKaGVCtSSp9p2HVKd/quOkI8AtC7q2ZHD9guMPtwDAX2svQT6HYScgX
48brmEoTQkq2oZi0kMPcaVyvJTuqkuipJ2mqpLhpzN2zbfHZOhgRQVBP1McAdoiy
WqmXPR28l9h6/2Vbd3zqE+/516yj0cMm4/WEhMHdWvZaG5imTVt/89z9gwHq7coB
hKvO/DhpSSwlsPjdGqDj2erIFXOObuNDRLUboh+aEybsCRnr63uPKTMkdx4/MXQk
yuVWtZq0EwGNUDLiOcZgehpb01oQmR4bBYDUdwrvvEkwG2gQ97GZPDkbxsAs21JA
yIziWwTa8zn/Zc3f8k9lFY9qlNfp61e2b9QcGzuMTFHnbwWSq26IfizpTkYyCmKy
gJbOAeZRcLgjVfINDP8pAxBZiojwG5zSjeIglv3Pynv0VLkWXhBnHUYNKoqJbgOy
t9RYrvQG0RE+HRoNcQtcMBxs0744a0YwuYH4Tsldn+gV725bxAHjBCjKtX0pFxHY
oroCSyR112hvJ8CRBmVYiGXcRapvvDKkD/atDtzcfvZDregjnDTFfJzOSxGht41C
yZjfesiBBAxOam95CPS2XflA7e9Cys8M6oWUx/6R2wzsgS7jgwxxXzAIQETtzwME
cx2JwngkVOXSQ6ysR/dcUqb+ujOiowprQ/UXJ+mofVLuKsd3hayry+e2ntPdXM5r
w2wn5Oaq2/zK2nSKsZOKdH+kSonj3jnyRGQWXkZcaWRwSMZWpAdnt48lYF85h4Nv
NexoxPXoqzvKEtwmI/nFlmEbasVzBWRTL7r1yUgMwmq+/RQ8k0QTVNETd7p2Hais
GXQWgYL3x2MH0nIXujye5HhiqbGmhJv1U8X+Lx7fOdQsDbmDE1b1Y90yq+JdXtfs
+bPkf+BfNvGHYQUXgIv4G9AvZtAp8FmsGIKLgUZc2HwR8dVXounjYp15dHj7FDGN
z4SKCXOISJvTQuJZ13JysirYuu8/zxL4PatSdJm/2XK0m/1p4K+lslSY9IuDhUxM
qn5P8LdrCbN86P1AQT+qpvjurTlYRaRrd9em5vZpAOcJTDrEG7bFUp005Sx71QS5
JAs6CYnW1yS3i7jBJETSsVMwy7vkvQ+p+xVXtW2NZaSdxfV5KxyG+jzypYX3LIls
/Auv9jp+PeDErzYgZwofd41LlbJdfSx75o/66/ruyzq2SOV5Ryfd27ec18g0fXXV
fzNieTHQViqcwb2ozs+4Rwb/yF7xxEoYLOpwcWSCe4axxhZyjl0Jp2/7WVEpQvWs
kW6gdh/+rGGgSWvJpd3x3uBmxZpeCT9wmUGCSsev0D71RRBLjuH3OU3yZg09kYn+
EZNOBfCrG1lr7E9gtexxdV41Vj3IosZKPfIdk9zR5h3PzGEwhnXzOIN5Vrx98jK+
j6uHqpFEzDunT1hEWkpdmFnB5FnXgJtmP3BfKEuQG7dlik7XSoTIGOcvX+yyDZ8K
8i804KKYNfaa28jW9jdd51hdWyBdRaVwX2LI9pJjpLiIiHjhxrWHqv5smFKXA9W3
qUkZZF9TscJorJfFG9egOgUK64tBiMmj0V16RiK8wDeVKuP/YaKDPfPI1l0I0q1u
LDYdJ0MWO5N8G5jmvxLTy4gVHEtZxOyQDTgJP/EoU4wzabhSci3DZVPjf0qeMKJd
l8o26yPrFc+NvIAni45XGcJL2PC03ZGQcDjHB17oJ1du1VFpJDBrDgvuM5PYjb94
qVllrD+xvaEkyJ6KTggG6a5gTyy7BY3/EQm2CqQOM5v5rMpsKzyKLhSyzfn2xVTW
8DKyzLAIWweDd6bpbWHPBASEE1c7VTP/FNyet50ciDsovEX1FLxK1M4ZmT7YW3S/
v4Rf4uPWFKH86Jpx++frVSPiqmu6bJBn/16zMqZaim5gSTHfCRBUlz5mSQTXZC0a
b28raq92WJjrMf7K1hnDm3b503xXBsodHFw6aYX4Q+a+uzuC/FOuPkPApdJKuAn5
dWkyt4jkBwDwiygx7xrYq5hqCogSWdLhvn8ZtJWZlw7HCmYZKYPrzof6wBUgSbUQ
5tom+cS1bD3Pj4CxIqriXaScdvtOzhHpcCLQyHmRtU93TJz0MOQftOd70lsLLJyt
fbcm2zeu+3b28875MVWwYbk60SmXoXzEcIIOqchJZJqiXBbaEZVBSwQPgN/TBJ8h
GqyFKw9JZI2ONUD7m6a6CItG5zEhYlUjy3Zo3YYawiYQsf8fKbXbo9HSuGt6Sfl7
983fAeooCOD18kKe/B7GaSi49IAk6WAC8DbrtFTkBNUS6WdB/Qs4KJ5PKf7OOYcT
1keDEGNUbuQ+fWVGZn/lMGBdGopNTq1W/U/Q2nNkXIyxohsoFomVwX/oIwEhU8OI
qU4xQ/ruH32A1dkfpuZ4jZ41eU7mALKI7AbSRBugORUuiAm1lCOB+UF19novWNMC
4pC+FOx2wbXforDX5H5kxW6bCoxkWD/L84qR9J7WmzFvlliQfRDHOigYXkaMRwjs
dOyDd9Jtl83qfCyuw6ihDKDsy6DFLSOkIhL06PKc06tksjIPX88rwp5mhg44Rs0n
AGZA8qvv1Ln6lJmN95dM8AW8dF7MLdJSiGWWLNjCbTs9BOx/A3asgj7HETAX13FP
+dXDYre+Uz3HsCtz+O11dfUCOZlOL95Q2gCUISKJOo6fm3a+uozZnrz2nkVKLQjy
AEnF/pksJUrG0Qa6mxdTD4VSafeuFlK9G36dktdl0dEMazwFWwWVYiKxeWBExnMe
pA8KuG+MMdGTS8GXhR6sf8g3rhrt2+8+j32tKvbxcFipwa997GtXbhvJjVu6NDb0
wLQ2RR/zgTD6UUnh0AHpX4eQS6Iclo8vBlMa9f4pqkizaONFXSKQkBvjAo2r/cDi
ykI20KiNvBY9lKMWd+jlsVhuZaian0kbrTbLB1qb+sQIXMSQDIer9nPlOnj4YPJD
GQYKOF6x4kYcVZbaU+ZivzWQcb7qa4OOU31vJbG3cxk8VRqBxxxInjP9Vgo6KymI
hphUMX06MCNbBbOcBxd7vi5CVoy7Prl2xoWJWZ1AtEx6GmR+YSM8A6rVUjd9k14I
kxbwNXHsAH+laV/03yLpiX107t6jKrMmTkQXopjCOCRa5VzIGyxhmccN5YMha7Tg
iVSx5opMV6rqiz9/ws0tDldS1EQJDcf+6LfnZlo8FEXs6wfBsfs1pI6aXfsniI01
0JDvPqDEIKgPm0O/pPyBXU/qAbduKPe2DF7kr0vSDI9JBpX8yrLOk7/1uTcdfY1Z
k9iJHa9zW81DOu/p1POYkVys+oyEu16xeMYzhK7aCxZax61m6t7RbLXoaJTj0dkW
R7uBV2wZmVWQuwkYl9ZORrZjarlipiK1RmOMzyk5l+IBSnqJEWPCK+sUxIfHy2zb
5T/31oPpAEf6sI+/Pf9M20UC7ZDapjLWlTekqGBquO/ntFx7zosW0mc39dSGzPqt
Tq8R86Oro3kLLnx6ZokxJzCGrpTZNYbcM3UyH8GDFWKZobPA+Vd9QDUjzcJq1c0H
Cyft4Jl8rsvcyI2a1oNxAU75ddBlBhAiI/ot57dnoyj+2+6Imw9OcmelW3XdUECC
SHysnNbfrxUUPYjCb6f9RpjGgN6ZAPTa6aU+PH9ZUNbtbockQ1JRRGfznGa3m793
IixRze7kt2PSa6cwLO6h7M2N8FFuPYUeDTf9pTYEhpFv1/C8bcX5ruW9I65Sj3ma
OSDyYdBeWCzCcehmP++Eofz4f4GW8bHQjhauO2rAtMYJdeJpgOAG4fqr+wIH5q/G
bxroxmiAUaNsvdazLBYzHbVGYmI9RhUEFWfo6C/TKa2Q3HQgKLJLuMjEZSqaxYIq
pJ5ZldfrZM0frAW4PduIy4IapFpHiEPyKoKCUV21835QzIZQnwfv3brvkUrJDOoU
lmxjTl5lSDT7SwYVsL+8ZfthXFyXRMIGRQ/E/0ekn+Afg/s1n4cL92zLw2wiGTBo
f8j7BHpm7ZsopFQFzWMZUDA9d66whEMwhJzuWdfOeVFRhiKgQaho4EYlhgxPbD1B
GzsdTV+wCetp9/HUilBzitvEFmedqv9rZM/+ymnpRW6fzLQUM9hLsg4CKoHlN36i
P9SeU2KgNSWDBRZerfldymnCx4lV/Wakv8VvFWlzbnUuxEAPME52IwqxHgRcUQpf
rppEIp06D5o/D4ZnATGrPziV7lKNxPQLEl0g8kyZ42FnOR5NM+qV0QstDchqfoxh
7PiPSX4ffZQ4qyzvBHSCGr303rgfHUpC5VCzhcc4gWns6D+dwSVzGbVot2rBhk4L
WBtshtTUOkWaLEq0R4yYA52sWZEn7k6nLwDEfLzE83M/l/O1BWfmUmEJcTHqurs4
EsTlXYm0VnJfMj0ro786x0u3rdaWibzSpO7tOdQXDOA3QcTu04DX+XE2Y3wHes+m
99DiM73FWIQHPbZCROz+D37dVlCu3RoWlRElTM0hkjCSTACYWv2E3NhdgeA8+zIC
QbfzcOC7y9SRgh7PYMiXt5rld5Lx4aXCHibWTic9OiTV5umGPtsUa1PdKz5+CYYm
Su3xdSLDYgt1C3aEKX3Qqss7dUr3vweZzVGmXL5zScoUL87qLWPByaXaLAhxMZ43
ljE1EEGidQJPZUYXHBNquumI57C+LQEFMJwBKyeK9jhbDxzkrh5V3LigotritVkX
fcPYqmLTKxiz6C6nC9PZKdmkDg3tKshyoOU8xN9/0IbVX08DPlJUGSC0O64a8ON8
YNoa+HUygH0iZ1DUs9fmcbXBGieF6Sa5fZSRkIc+hZ34PyddV0j+nK45d0UgF3P7
QbAB/VClgkefIo/b/GQ+iZesSlOOPoLN2EIthiUMOJYIf3q+brhhrTael2DiveTd
Y/R78UfyyQiR4IAmSuavawRoZYxE0FVndSuaFHVDjPeIislsLTysfgRqfDqk0ZaO
D/el2MhtSS+qVRETFPFhCScyFCltyDKNW/7PJ7BuRF80D/0Xw8lDbooFsG6pomVD
buWUkxX4AF+mKHyjZp0EEwVtsMpMdtqKVgYc2lf+7sF7hWBU4B7cR1Bs930vjcBW
dhbKNIUWeDlIxGGjixp/8H6vpr0/AJVk79TkOo/+KWkbQaVqIxgHtYzogt72oy4b
RtB+KXbljU35mYVstRjKqA+FnckKqQjzvMy1jbVwjOWhsCC25gIN7klXRep0HXqw
tkZGnULTT9lXCrftLOz0/ZkRmoKW9HLjOM22oScSegPrGuoePACVOTI5GdBzW1it
PXCh5kBxkrBftFvazpmP4to0C9RLHJeXO8tkdgZj+nhY5E0CU3g7nc7waYNB2MWB
QggE7NCAWEtCiqVISmfdRIpYM/nM+pI8jmxaKzsgiIkR4GouJYERlhtxHbBz/QBa
eLtYOM72hfS7iJROd885B+BrNcPp80EIuVYCSiYisp8v4g0lulLoWidKCUypBPxw
7MhPOBf36QhErxwdctLlVNX1Ag/zbusCsh/ksw8C0IaSH2H6iTWdh00Ly33tKtTS
e778A4vqRudrTpJ/jQ63mcjf1/QRfSoSZ582IF+zPAGx2192kUeHkzb6YJMYiHCh
Kym+ybauxyIX8dtzAuceKpDUPDFS0UetCN0kC9E8K9/v6YZCtjPDNlK00+rUcpOO
wqEANMOxpg9wrguSavbsivo5A8YN0Nm10ejpwejMoSHYeCbdXomKXx7uSu0XFBm9
iQ6NS/jZuDWQET5gWBid1El+tLNsTc0YMMcAl+fWG0UFC43Mhcexj6HfAq3KMMQ6
XnjCcfTB2pOGqjsgp0cEMry1H+wyUVewrGECMK1bDJ6JS6DN7No/SlW3UAZWwi68
r+YRahirqT0viFqOIRDdEs30lixvfyo9DfQdyUI0OvdffhqNLqzDh0qOxPGo7gFD
AmOZ3f2/SmCIpv2KRMDulHapOlXikUr5OFqhBeqzlLIfuWuZY8DT9ZIgUPr92gxC
twESfAmGovbP3EGBED5OdNWXhKXpfrcwEyiCIT4HjJH9+qEpsBTjX67QrLXHgYtp
8QVu5SNJpS1QaU38d3+w/lm+FRpQ+zTPNWhb5B1ZR2QP2B4qvBgOU19exCJ0Mgd4
K5fGpH4sDPlLGO2nEIAaRhDUdXbBjJcAIBBlzRYjCdFkNJEzwh2MFRUkNqgjtBn8
VFKnclI1VXpzbcG4hR0Bb8sDmqwJPQ7Zv8WmcpqfwNUSmn/TQMWjjqxIFNu8U6ou
9f8llI5xWLGypeWZzFVPogeqWCjBwa/gmyNRg+vt88YDe9MPlIP41lxiq2EHGkJE
jMpXJqENuP54TzMJbPXKPFO2Pwv/fqLxcPGKn+iTU31jSVEOKag3DnS5AQRIVmhH
6kRN4gcGugAOnpu0HixYaQrKPGjAtZXE4ViQuLkyZRbQIM3v7Tt2O4I200vovvm1
/GxyDrwp5Mj/MVU4B1lvN5lgUR01lCpiKYbcd/F0mtgYDJXMf8VqpAy0FcPdJN8G
mHODBfpjvvRmE0ctBUgXwy0js5MQmbi+W8AirEfWhbwmGlDCbT4WRmY8FwACASuI
jty4exNbKUXH5f7Krf8YSHk/zjIISNyY8+nLqFzaxEtSbY99KUE0pCsnPun1f/8u
QOLzKENoqomyKTbT5wIZym52sS/3AC9cpJfTkCfXIthNprO7x63o1cZkqAQBU+D1
3pPRJX2ssnf7Xw33WeE1RgIl6Iq5hUpvukMdCpL/2+w0M1nmhxT763/RED+9BirX
9OlKT72Iz6xxR52O2CdZOFuYinkeMTdbInsIdA5R3tB+7RV7R5MGRyL2aR8na60b
69r24QPBEUhs1/GtnWOHUpIWY9A5kJCFtcIZ+zo8ia2aoQIWLv9XIjP9s1y4mglZ
RKMPVjZ1Uk8KSVv3oK3HI2KSv0NLg9CRqa9frftdBH8REFLzDmAzgBJEIjzKXSPq
pjQwKEm7F5qG6MkFcb++P2ItrsHaIILcWaTob+Kck+QPwkX03Du73wZFVW+Tp6hu
4TAJU9yf8ciGwrzV7b/eWlS/pdsA34UKp5TvvR9ZnMzA8PlfSLoesvFDWyJIxqkf
rX3mbxKx+FOEyQp11dwqxaZkWth8xiQ7cb0BI13+pKoXV0n4gMzSTaxpkjnticLR
PHXneh2Rmi/3XLpzXDz9dhMkAZYWGhr+NPBsbADQlMYIWNQMiuPmD+y/FaAEI6wZ
GSOGli5hdBShlfC9GLxdd9gr64+SX/+KbmS44KGAlU+LV77xjgYzWcFLq3yd5N54
0YYC9m358Gw1ocKxkwU+Xsto9i8CAk43gw9nyAlZVw/MmOqV0wneiQOr3AhivvgN
ywoMRz641bK6+1bhkxF/gXGgTnK9THDuW2mvKXOILVL50EqTI5zGJu7t5Z/g3MR0
ojDl39NScaHz9Wo5LJu4DcsYv0W/Yvld2P00+a1pxQmpktQh+I2RgDe2w4brKfZ4
O+R2d8z6fdXoGQYEflCy2Dw/eNgGktBDaYR+W0TLjzcauuYJ3fum2l84VshYjfjS
GCj/G18sUjHozqGYsRLu6R30kcjSTfpfSweH0rvX+6lv3af3kQ+ubffUwUWBv29d
uX3U3eTdfNFw7jIgeYpunbVUT2uG/jLMY6jOB9BMCtSlrZ7J7fhg9tYw953IRmdO
KufIKUzbNqTBVhVv6b5vv4j0lne76QuljMivHhWBjYuwlBFMNrzucRhyQ9ghNVAX
dPt+dN86OsBEJJgFrCMi20R2nfI86gRrMNfrjpn5u1KQeiYHTp2gO6Sf+HVo4Jxm
hD8l4I52GReRQNkRLZ7HicU6ndIArlfPRZAmn4kKQobql1Tcw/gFxapAekPMYk0n
GISi61YXXIcET8f3qP7NVvo9QgV7fQ8mR5ifrKFc/N1DAQE0UykaKXsJzcGLSlES
ann7sMGJquuAdRLxhXJenWjIBaX729fupl3MyBGgQfuRm9IUetMvCVSfont1VJLP
yEP76YkZF6Th4DxOiuSgKw7Wa6Gm0xy/2PoPfQPC+boH2ivAP+FeS4SmUJUd6Nix
/6+Zp4dE0pg77ngwjBPxWTN9tBq7F3F6CfWEsjWrhiKkZ/9w39J6WOfePUxJTmqu
9BSie0z+G3mXgVKNseHZYq9XnLdJl29lEaVtRhHHupuiwoc0zBwT0FA1zGQSPBDv
noCIpVinownlqFVmUCWvy7SNbPxVW/3OAA5bBELaKPuHnItAHOz7dwqWyiOtjjOo
n/KK1rmad7vfctqKfs0Dfls+2NckAxwyh1H5txtdXOvKVLVhBQG9PxsU/OWZ2lCq
2Kk99uJio63r/ntiWBSQoonIDgV4JQO9bFkBM+SANCr7PvyiZlQxy93E71ErY6RU
2qT0DnHoIijS5LqXD92T/3CL9F1/KAGiDg0EImVyPGh+mvaGsG75Bwu1chAIG3HN
94kST8xUL5aDLOzLMTLBwieTF/t2PGBJc5FPdjij++QmAqpeuiQ3vJhQHOVdJeFS
fCcABuUmGrcHZoDL9lNPFs0IcAPmgpjGFrrE49YALtRxQEQy7SokE2MfE82bZEwi
0Ye9mkMlojZHffQmBzMHIg==
`protect END_PROTECTED
