`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYj2h+zIPQEe6prkFezHO10k5YcJ3twCewjmWar7PjCK/etszUPNhlHZaDZJzoYC
XHodrDfRd0WvMSBsDpF/OTYQ66iKf6CiwpkYPmxV+zXwPsKcKq8Bh40OcKUIUvGo
KZCJTKsyR0Fx1QRdnMvgiT4YE5Nd7vxEdADuQmerHwJydi9Njma96vAz/6mnn2La
F7s6R9EC8Pn7sn1caA5T/1TCBMJIvnc6+nDNa6OKx4yQ7XojXYy1khloZP4bZ5ep
LjmqNIp9URwxdS3NmV46PSDlXJYdTqIB//vyGYq0ieL5JPvBIalb78y2qUQVNTyG
l0bsXHfzKNvWHOxRAdpytC8+98x/7BypJyEkXjKwN63KhXEapi6xuq9W/uZQW4ad
b/UgpwYVYktLFBjjQd57C9LyGFU4eAJcH93b1Xl6BM4ENO9hFry2Tle8E65KlfT9
vPZYFnP/4vUJm8tvrix+ebyiEaF3gAjfp2XeI3vXHbI5bTkfvRDZkBlcvfzCW+dL
L0IOS4mzT25TrykHW1Lhbn1MP+9wTjx1WCth9NJUP5dMwmJBhJi3ByVoB4TlqCso
as5PTrbHgybEsziCyBV+5eOi5lQ7iUcbI8ANy2mP3aeuoqqZrkO4aBKqbfBogoc8
pj4uyyCyh3083b3EsqUW0z50lwKsAr46GG8mbHZNknzInf3svqGL4lmadj7URAok
pcRYttWishgOt7qathPGA/OqUNAAWcyyYyDKJTuV5Bqqe2HPHVz3LFhWItJxfeTx
POiz9CjGVquuqJLVVV+HLmcF8iHrvMRIz1HYecH+O9ZbcfN/A/g4AkW/S0MAXEZW
J74UMBCNlPXcskoaK0nDAQx+EEx/zSB9pm5tHWayCXZsx5rAuWuAjp4S9W+PtQvU
CPcqkzp47Avjx1qjYar5dm/l607pjlUnpx5yIKkgNj6t9rLCWb/swfSumCUzVgyV
wBUHjuO3P+6eISLeSFU5MwP0Ydc9s9Wy01USmWHok+c=
`protect END_PROTECTED
