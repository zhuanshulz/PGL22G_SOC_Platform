`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IGf6JgP6JPlB4BIX5ZzRnwaOFM3obhrv9/B1EzsgBMoZuJtyliobECNYiGm1BAqe
2toILPuSSUXrNhGX7J1ckiEW4wh33MYMfkcWh9tjbVOFHUii1ULN3WYc1gzKFKFu
ivaqswT/sx5i4A2BZE9JM3LAxTOijryHhh2wKlfKg30p4atgQz3EUCsgkSKVYD90
+BUznLYE6vhQKxp373+SDd6JCKyrEAV+r0/7SisRzsTEwh/Xrwn+5PNet6d6Q4ZC
4m3h7g+EBhI66iN1CEZDFdrQGqJO9SN0dxqewsUmi0U5jcWePQMLpkumFeISFLSz
VCwoOxtTIkhfttxMpX7/PMR5jBl/TkBxfznTMWL5nPo=
`protect END_PROTECTED
