`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssmJDBIFwNaH6s60tshlx4LL8ORQdXdHwsspod6Tajlyt4tDby1BPLtUjYhkdxuq
LsHsJ6ZD/JoPWcX6kVFoV2UDwRnWByNkiLmMUa9ZZ4yopNWeUtlBts+riNaWjpKs
So9zQCHmlDWeKPA0MUXeLFSEswh4mxGybeKFn94bT4sBOflukpVKgn0cn5Hv/cdV
6UUkzVZZdthLvQfD0Tgg17SAoKiZp3aPu59WS0l9Mv/yBv4vrKbxLIPYfYvuOLse
NH4IsNedJIefhGxOSJP0kHCqtbz6xCfUiwK1KflMi5GkumERXq5oOsGkw71nI007
YXka+qetVUufX/N00cpTofmShdXQuUG4wtF1gLsRtWEtXkoLXWbrFj4OUB5kgiMQ
BLeQ0E693AzwG9c/p0vTGhRMa15LdpmCcwlxTPaW2eJfFd+9s7g7EYqkbu0sEzju
jOYvx2e9n8J1EArRIHdG4FgvN4Gl/vni54oXmC7ZquhfLLEQnCDViRavJ4LXry59
Q7f4O/v2adDhl0exVQeVVg==
`protect END_PROTECTED
