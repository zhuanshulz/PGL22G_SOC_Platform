`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmAH6hwjq+y1q0KDar3GPl+EyHle0aIpQx6zZNePmHpUlvVOBnQz3AOBSUrS7YH7
VCdf/gF+geW7Iw8lbHR8Bbt0Hgk1lXQDPIHtnkpz+R0UekEZwvx4ygauUJnu7O9s
1fdNfKZihXERtAdiDT6iXYmitBWYKTr4/vjSwUGtuzeRmS4izQxq9BMWMo0AE7/4
TkvpOyhRhbVUCAUxLqr32UnV5pd/NgsTvnAEA9HFXWTjF98Y0xHiTfbeejHhwumQ
OUbwwPefzBToJcPlcSRu5ctl4cJ4xeSxE8H1eebkgBiMKBgDrck1AKwtMKJgqZR1
2kmKn4pb8hLTPo+Yhb6+QkaNop1kuMrVEkA4vNATkTSqiSnWzKpf/BhOtQnBsWSv
hivJsWMVrLSK/8sc7xpkTVSFD3kzM369UoinR29vKNlasnmTki3TJzFAWOeLdq39
sV1/kyTGHu6khmbspHIa0E903ukRXaBjLjxiu7Ls5joDaXBJYCBrvVL3X+QoNJ/r
H/W0w5qpi123lqulbH7B591qbdz++KHspNHBw73ra27M6pKgv8gQ26pYGjQumOks
eMMkRmBKnTJWoRCOgBxfXrjc8bHTjLw0feDwgZKGwbim5DT0gTvzAZaQbOAESBwM
lQxg3sSMf+forNTLgOE32BTeBDuZlF1dUP5VpCqZ51sIMF0KmZwE08VIgxUaznwG
XAZCmkbPc6r9NhVn5oK+rzr2hBh4YZ3pdZt5/9iIww0DjfijGwLtNQB5cbqk3QzN
BMYJNekShBSTavhiM9+b99PIRThGQNRKz6rOwE5LcCDqg96MYZXCMdG/Ig1HZqpj
xdKXC2Wc1tuA6yFxZoFzFKe8ziFksTs/A/gGAcuyTtJNgZYSqQ8lAJfxuV+Qi5ZC
TOdSmuWBASHzSkSkzoNibUAlw/MwLggcljG9PM6xfzuIFXRS6GweFGcwpNof0IS5
BDoyvArJIxs2NdiXY8xxiXJL8d987X7ZLwTLtS8Q75vh+o5JK+R7/w48a7yKTWXV
2lSO7+EcA8cbqtVos5PJSmJ7EMxMGKTU+ALvc2R4tY1NaU0n+JZulf5yezgz2sKs
7drFIokVFMyGSMEXxAu7WXiyRbUwa90vCnlda8c07mPkXLZeP0zwWjd2mp7OBMlD
dFJLKWLLD0JvVq+LqsUqtGOgnA5o6wppCQumSqQbFAL04LWn067Cgvc9hdPer6CC
pFmQ0HTr1k2uWOn02WkY4o+Fjo7FB+88S/bskuhLDLi9BvnxmfFY03VL5LcxbFBB
3dIoWqxJLogWPfRBqN4TXqk1YPGrUC9NmMPBOl1ThYWntJDHuYZI5oo/Mp8m+JEh
m4c8D45GBHjMrsiBrImxuKl7lf1MH0fClNoatiUFsCcKFrzcJXirmUI7gNDJ70m9
66cSiiAJHl3UJIXp6BHJMOUR0qLM9sbaiXOO+TED5GFpbpBt/i7a+i6wMIk7fFVV
eYgoloSFO5QZuX2A7NLcc2M+bfuM+bsTgfbTW8FpwpCsUKj/akOL88WpBszE+7ld
qvkzdAyr8NUCjOMd1dBbh9jaOPMJxLRkjmFqClCqWbXOsxytGtilqdL5LHfcUSY2
ED1/ZAeqtKqxlbZPdLvFTLB47BuqGv0pF4rHZA2nMtJX1DZ4MME9ZohiHwh7OEc2
ZsBfcFnbSItdolGKdewrd8fue/yxI92iXF0A5vpUPXO/cxPgWvecS6Xzqvl1lgep
U3AkHcHJorukYHdF+D47pQolQgLyDO+85mk0y6o90h77a+IXELyokOg2gTuq3wHc
85EwXI10w3aYG7kaNMmZl+36VES7TfxHAKbB2vYU/kACncYrJAMH6YgEim0XD3Bu
5kcggugrfqY3A90RyRyOSUBtkYAb4XwPHWQPIv0ZSUgGRbhgKf7nHv8+yG4v6D4Q
OMxoR9HCCam17q2lQQP+OrY+n2LWz9ifovBGdXC84nO0aePVAWrTBGHNgW9fQWbh
zEHOj/lp44Flie6BOC8+WDfgm5VcUe23NdsMBecr5ouMWwokkG/Mc4VJmY/dG9gz
C61nd+c8ab7KyLHuuFBEAkjsQ6mDbyHBbn5qbCVDw86vqbIYZbXCxkSn048GiTdf
hkc/17HtR+TLtttmDCbBOyqnbgkDTky6Klb7b2avUl2KVZByhKAKkHfF1WZ+5QJl
xU2Wm7MDaPFkzBdBr+XaP71WLU9/hdcK+CwAtCRvgkqQvbH86UBizF8+rxD0NKaU
yLiEuHfVBry79nlGtGZybllu7c/F7fqYFVDgF4WAZlVx9W5NXrBZrVZoWnr/fCBq
Iw2U058Yuutuifejf2lkavqlC9pf/S9zPt4WyjqEo+cBxU1SetIH1ESCLc5oyB2J
dw0JrjA3o2MqqlGxFJKrUoJyM+rdNa5Uc7odbAyo0pmb8ld4qV0/D+jdRZSlVtIS
jgYDgBpV8vfYtbF3fbvaz0rDnSLChAawKwkUSt/HnKnPF5y00kyER7K/HPusXmiC
HFRe046+gjAVD6t2yFr531g00CNSABcZ86IgC2KhXWvof1EzCdmFsnbO+DaQX5WO
YfzWFK1v8Cfl1ZIe/yhCu/fDRTQgdsAkVaTl3EGOa6xekPfF6h6FNeMLRKOFZ3Wm
5iDGsQ+y4X+oqpHfsHmCHEcyhq85P3ZKvVw6l6b3MHt5H64cc1KyMIlhaWplVDEl
h3b46D1GoeINKERF978Su73frwwbkFcM2xLu+TuHUHK/tEGeT2OVSNK9IXyUwQEg
AnXIPSoVSBqDxzWIe4pQKfktpJNHf1d/o20+heERWvPBdSOjvfvmcEfcR6Upa7wM
BTcdEt8M0r05QHrCPYHTTmBjc0M5RW0wBO0rizC/8tYxYInUEdy9q888cR72uI7Y
7QL4LhHEnhxOqzp2q9w6BC06Y1b4l043c0QOdS2DZ55vRvJ2k10m7i7TTJOWZijY
TCwlMJD4hAjc8OuGoVjF/anCDLiASo+qDlaWVu8iRIOnxfKgPneQSyqrQkXDGe2l
kcJoCcuWpQXZVcaMBQE0rdaGJZIYWx/CbmUCeCptJKHq3SheqzM2etIWdd75JJ54
pyIw4Y08SUtIcrey5xIZLL1M3m/rlHgmdsr6bzQ8WQTY8FEK6+H+Tp3flyGXqk47
fbA2O3G1UqAVZXH5jrDi2LVs/1aNwvaFqaGBc0bZarXlGFSUdZzsGDxDP8hXtjve
ZyUfrXtQEQIKqhK7enWmuKNwqQuJlzUA7q2CLsr09+lBo3V2IPimUnZL5jieIBJy
5TGRbSX1Qs7D9OrUyZ3XqAqhk8ooqEB0wrK7wznHt2/YKcUc/8DTyeKiC7gyOy1h
Cm1rhy4EMTKqhUbp12HvOMFPrKsUq1XPSoP0vPQpZUUKDJgxidSvyI4nsnYYgJdT
h+U0P1MnJdGXnSirDCnZwd1YPMMt0mL6ugPOFoK5PF6odBRrk9CFVq27kgphOCav
FXh47sY6o10KZVD28tw+n8fs+fWWD83kXQeR7lSTBgq5lbHrudT/jcmCGMAOWTw+
EwbejjctGfXVIEcpOlFUD4e+zhtCVQ5XMl1+eZ4x9NXzdxerM9B/TGl8CAlmVcHU
MVpsGAgK/XYvcn65NAFqIL8V97CEAOgIWip7kVAw/LyAATOIBYAbLZ5jZcX7dTPt
yJwrEmvE6cKROb5IuaAwq33et+mdKFYU9tu0d0PzobPkbvLGonT8x+jdJch53iUP
+lOpo3/hF56eCfnv6JieJ9u2RORg0ZLhRSy9RnIuuu5n3j6s/ImxtlAsI3gWh4dN
LDmbQnTq8YUm5mgSrwdY+hBDPtR+HcSMk83NZSQlMl8T+w1KeAYT8fP9Z7vmL9R3
BeOZkatwMDa+FiBMbgeKghpEM+Q0sw0szboyVn0n4r9t10C39kJl21rtR8sCyCOv
VRTEj3LrdUS0hRv38F64fOJFTC5+FiB0IrhhgnMgL5foVV15qeuQ7cRk7s9FvYVU
mnu6D2mjtKPlAZkBOoeu6rtPwYmRLTCZ3aMIIJ5ZCO4aOP0334BVqM0NC8yYQAfm
olAneZczd+Ku6atF9dX3QZygsgxOrwYnHdNSJHXlBDqlkwau76DXnq0cCSVeTYND
6Dun4Hxo+IODcW40ugMJIpeps7Up7Qh3KVdLZNkDjlLIjyYD1UKYFJbMv+NnNFQF
5cVQPvnBNufH44uu03Sqphm0ofYBhJQGAEoIho/oT0uQVFW2Ndq47L3ly8dEtE4n
oDluZFQgfBiBVFtsZGQacjYTYqG/u/KZz+PSktv+73Qq3HGIcuqi468E7K32R20z
DsY6K0ZaxxyNZizXF4n8GmrL5jb46+zCTXvLPemuN8ZBlasz37/3XweZG1WD9fKl
Y7motVOUINsBdr1QALsDSzrCa/vWvB+551PjUBYJol1fPa5aTM0wOSXRe8VHJaLg
qgrwmte0eVVRElWAIY20G60493ecHoIpSYdqLQlT1PQirmXOoeWVkpPE+FjNmVWq
7yYEaUriS5uzh+MU4NsBhvc00+S4Jqhud0A8R1PJRFVG07YWLdRfd0pHqGllC8GY
Jn9Z6YS56DMEifGpsc0TzfhIgVS93kIMpNdubXaSfccm46tHeX+3onr3bm/hnUZ7
gDYO3eTkDnwGxlaTYmKZ30Yp8n1/k7dZmKHao78wc272dWBPVFfYGFbLnb4zgNaK
2L0YX5MOkmsvB6uJjafigz5SK9igq5+QoD4qVLTGEGMI3WeCm2vioNd4rEu+0UQz
LQ0+pWkOnP+bkKx4Ke5DKjsosPALZu+X9EJu5juFQnsarrRhPax8DL3czsvFu5Mr
hFm8GABE9caUbdNdQY94zS8WBvuU+ZWcGVZlf8SvSLW8kDGdNMx48jRNEdGoL9H/
SmMhJVKbqjufba8ercUVHi/IteZByDtGDBoEfuhTOs0P6Ia+ZE3OV/pS4534OphT
kf+Z7xemc50o1cIzQOlbehRc9bIwqD4rS5jXHHy8zncTk07JYHP2TKUGo78n0Y1V
1uxoasJv/mwQIXW67CWyQ9FhzFrG4GCpLB2YiRYQ/empsO/ucf13SG6PAezzfqLh
cA/4zlc8qzu47q0zM0SmaxPVhY4eYXVCDrNfBypI94E77RQWVwMADuicOJ/xl2hI
AnxBN3js67clhccQBUNkoR7+CPQJV95NOkcsttZkXztYDPGHLE63fJ0aAKOwy6pN
uMyNnlVaMc55oQkYLI80ZxzPx+IwT9d2j920YlrfVVjwa5ucgh4Bjr9Az+OpQCRC
lMzh6rV0z5Jer4N/Mkspb45cuKkx0lyMSRJD5Fap1U36HnviUipIq4IOe/ii3FSB
FqbCbiMklVm8fm9a96lfZ0n+kuOpM5ntlgRmq5I0by4Kf9HEx+prbJoMi86cfrCw
+aDSsqeD0IafnT80TDLiS/QS4EnIsLw+LPnIK8djEYiiwn51QYQ/bTbpUxjdYkC8
IEh/QHANgBu/wiVkrH5KF0ggiNfBoKuVwIynfZmyuUoBm6e4dfQJDbhegUJr1pW2
f9/5rEXJSD0V+XGv7tFK0q1kIy+kbUeM7LQGTdSw2f2cIKxOAeES137e4DR4+oO3
ryOkknTLHW53VMMNay398+mO2ynI8XAgIOVY9yCKZsAUHQRtmrzJkk04f/CB6tv3
Uc8V1sHHMYMBhELeMs7l3Ohk2d0aeI8zjRylOh3VZBzLBIalpZvZGUqwOwCjb9pD
kljk9SrpSO5mQEmJ1NGFCSNo1UAnBurj7e6CP3F4o+YxlzX26U+YyferZKuuniXZ
Ef8gr2WhKI3OdW3HlMYj3cXRfB+5oQc/5p4dX3+pl6U2kbzuc4G5wWVxRtFdkwbC
QOhzvLXjAg/9DMhM9Dm6r2kuWnzzqLs4OK0QalrcKWaesfvt4EzY4Xf6m8BZcg2A
6dsjA8gT4fXZ5tpABzK4JSlhH5SWZ68XYICwE4h/p6vjkH8F8wSq056Fz6oIGwbI
Udpmt4SlZyCFWCI/zWw2+Ox82SyTFQPVDAF5pogExxUlRKp50oo8g4nfRpGHZJHI
h8wXy63u+d1J6v5Q8lbPriO3z7jQvbFp6qvEyrVnLGqZ9LwfHVtovqOUhL5ov16o
yePpQCrZPY/JH9MLivXFW5F8Ahp9bPjJaMHHVJkAJzYkocfJ/74hFgOdqVBkIOlP
Y0q3oHFRhmq1p7sKYAZmGnawA30ii6d1AbVfX5wTIR8rmRgA/t+s/OG0js/keYBo
zvs6hUoiWV+8R1S0KQq7OIjv0kLZsplqM+gs15CV001vZHAhfqOEkNlVs1VKdQse
9ACoJZWFdQ+5iN0DlPB0abWHSQoaGcKssvCnPxOpL16+Q389vYJr+S8cY5mJ5rlL
Q3LlI/RyM/LQCsd2gChLRHRcthbwf9JqNFzmJMjhDAoXWFfm77w5pNLOg75WRQHs
rxBfq5VBI3cf8ogrOz+1ZVpvJt50goJ/j49gYlYIOn4XslqwUC70OmVhELebgvhp
RdHcPUIX/1ZFPbZrrVQLh2Z1QOavPIlgORwyCJUqq3TXfyDHplHG0j45pfNFBN5F
8QasF7iDGkFl2qaNj6zE1VkGNRAmBjdWua26SxQiiicBCAIYaknJ1KfhdgIsc9On
9oqUBo9FUsaLhCwcOtc8kErIthgue9WClWwteVq3u6+MXK09jINcDs3H8Pj9g6kr
m1mRhYk1Y6N14BYt9rvjh7WR+Ux5BODQ+enCrtHGUj6Pq8EeBkLR1fxS6SPzABZl
yGXDHfNGufwQs/F1shD1rAN0ghUY2/SFZXf32BHioXpB6bTN5jwjgg+g40e/Ht6u
k6JyUIh24oMBot2u5tPur1bTczoX/HPOfrV4R8jT8c9Vzdu0VSv+eOpeqjCoN7LU
eibzpDXU9ShoAQNA3A98nTiyEJIP1H2thQYYgoMrsLl3QQdUSbtfeX3Q7Up1oG2K
FNnWxXslF9ndbAHexqXLD6Nl+e0Hbrym9HoMzGKzJZTfm8dtsjEaHukzMd/G0yQW
mP0T7NgOxAb67kn1DgJUvHBMsqqs7LhujPMTeCcwcAkylw4e62W460DXcKGOkf8o
4WdjNxkKIRUJov8VuovzE0qCdqGMqJxcMEJ+qJ3koB2EcuuPqmZFKP05TRH4Ys7c
ZVvN8BkTEpl5gt6TQTmn1Ef5hsYVLFCsgphoC9R/WJGK/nfzM5JwdPSBaapubMec
UnzY9zUL6YIVkCyu4NPjPQ2n0NCo8ghnYw/mT081gxenr+XkhDWWrMfaNDoSXoSZ
bQcs7qG+46HgnlWKG+t2YbX77Tl7XYjG9PS2S/O0IB/7utjIU5pNvFONHGAAzeF/
WWjxD6OMPaIGCAW82DLjhOnH03GIlR5Y8OGgjvIFn+SY6CehBu7JiLwo01W+9Ga/
sSKCLuf523xl4MoF0etoEUtM599PZnUhqa2HexbQyoxo5eYzf5hyttqp9eb9HnYf
eQbiWpQ+HE83HeYy6YR3uOtDTJaIUqXkDECNqOKX1vcfQWZAEzYFmu3spIiRrl1n
eY7TAiL59XeG8bZH+5aPK/4OyNhKlYMi472+KirlwaLwPo0mtEz3MIaY7KMGPqBc
Lr6hhZ3uoIM5bdB/e34EglV19FB73+07Qzw6sk/NLWG1ycQwE1EyyDSHuy2ws0h6
gkXQ3u4BcoVMLCginQZXlVUyvzgh7hl5VmaEDHrCThez9Hsj9L4LdG5osmlynb6y
EUHkM+Iqvi/8mXAcD7faoFamQsR3oa3S3P/GPfG+LBXQcTkoiJqx2G0qaBd8BXlt
3+nkixKIPPf/XWnorTpnCPfTWp3QVuWp6kIT7wIP1axw3+wf+u2pgaqnhei11Bjt
+eP9KH516BH12fx/JD6UqdKcyeTsNMydbNeZ6RLYc0H8f3F1u5L23BnPFJ4f391R
SAuvtdYLcuBrpSu4fyNL0yg05qTjwCCJ6W9BprNLBbo3DeUCTwou5gmTRrRXOO04
rQ9P7jkjUjCZ9DI8m3wC6vdnHaMqrb/RT6BBI70De582W7mn1kqlVsXYouST0hB+
6N/qsbjB8MJL1RXvQfCLjFjxphcBqjTfuVcgOvCevztVjdBoE3Oa6QvgT9r2iO8f
k+CX/HZncmsTZAJxl4kxwWDi4mYNJp9jC+IH4g9LRXA6dbS5KMLKS2jaFEiWDtRm
QS4tAsvVkYUds2KbYtK2X4TB0Hta4WB5spOWZ4356Kdyx7qVncBiCoO7yUSNbbww
tTaoPqogrPIxTY+ZQ9T7iaRH+5k3oSh7M5V7MUQZ99AL3H7H6/yE6Slz7CtqDH30
JLaA0KesYy5KuG+dviCaPG8YieYVR/L77ogGhCIeUIibqwRvcD3wHipSZxkdS4Jw
EWA9NApGezvepaUiCDcX+f3JKOOU9nwSi5DfaE7SsELhokZsDgh92U0GfLDQgRV3
hUgqJkBP4vAPddvBP9BuL7aK12RVbtelVUcpriinynbclkcnFKswg/Qk6XRIy+c9
unsZ6uGjVvRiG2+fNVf2wrZP4HyzlPtY6N1k29LIY7aTNfttGqfmw2jsdZkEUaDU
AmWbPDc7frjy+GdsnCIYwhZjTcZ3L8pJTGRAdiLc/ojDbdnjFnSbmpdho9udjm5U
6p60HVWSy4s0surJ+PrukDZDSiTtk8JlcVqobj3up1ErdkJnZFRIlBdqDQ1WWOE+
qnWqabQJzqAEGbZa1y6VggP0ZDIm4rmYeRpUfUja2LQOQOBBIk3dpaGEyedqYQ40
Hs0QlFcCpxkfPUK+rc4can9ehbYeSMUA1dtEOiAQMs4y2mbK4Lna3XyP6In04/5Q
86PkBGv2usEOYaGxJOpWod7EiGYHUsgE0FDLH5+S+FJT4acmNcTfPEYlT8bbcnI/
c8BktIuTJPikNHDsz3FtWBd7xMi9fPdp2T89tdjXXBjZRLsZasmehuvvsGEnyBq7
dDm15rRTTsoy/0E4GmBhoVP8bKP0u2HaXCQ9ewiQTNuS4vAXxwKXpfz3LPXRptbK
r1rLBmgAjJHz6sgQQs7JGfjisGBSlRBqnbxy9P29vxgOPHE/NXwI42UsBWurnRP+
Y+Fpik1Voez5zMe2LGAkfQKMk8BY46M+oN9LjMSxpD113Mj7yD+iJ/W2iz+P9Vez
mW0au2mivQtusKI/5UEREjMV+izA0jjb6YY3uIQeQ/6OvsACzQ3V6pGx9/0Xh4VU
jMl8rPkoqr0eOm1IHGIlwK1w3wZD1l294etAXudiut9jaMLBIkKpZovCLndVgAsG
d2gesXff/FyNiGV6GR0yH29wyHoJYFgcashAVHBlpPi3yXd5kp1CL2ucAUohaCET
aQGEtwKOJiwBrteJMYyEGtd7/K1UQ4+wgOCdpOkxdBOH00ieMrN7IPTr+S/1Uu60
joRJB95RrbjhTHl4qc9zNzijRGSAdTIbLJ4crYg4LU697x/pU2ouVYbgbAhoTOkl
KSAIjMIDAV8ZTqCQbCFJ58UcAncFFXabxtEo1FtS94JI+r1ikfETuqt22mr5IaFQ
QFXNqCGLh5V3nO3FM4XiadLpMwXeRB2MWg2atDM+VXQCjrgqpvYTctnLLTYGtdHi
0Popap3LaEvxedmPeiKM78rBvwuPMv3MDncKzfOEMZqdrjSgJ8+jcYDrAdR7FH+J
86LcAkj/fosD7MDODVG6vkBmXqCRijLibRhuAKvjLPKAiiIrlhlPw08NDceUPMHR
FNhlk8NlGcU1VdxNkEie3DXCJ9RBJXN3AbaIOGYjASFEmxByeGdR2hhz95DXGxmI
nrZ3NmQLKB+j/hkrdgq3iVGnuVCwXcoYGVuH1N9ZFRaEbAxsOVVHbJf3f4RiCLch
nzk6ZD+ZYm/skSwGmtRUdGTzoLPZ4scevSvUJqZB6VTigV+jSDeMPMXM51YNjIsJ
kjWHMtQnfnlbiQoCmnL5Cd2jrTDGferfPo7IMYAZTYs85vP28Dk6t1aUzactth4s
r2pTbzl699pwpF4eQLjkDA8E1pjY4fynoCu45kU7zzByiWxm1iRwagwHyS6RdeeA
CdcOj1MUi899DpORW//jw0Kr6QUDHKqUK2lDcKsEp8m+6G59wOKxbW2fehIJs1AB
GZGnKj45zc4QmbRKEcFROab85J8ZewoLFdOOIskJ8x+C2YoauO1tZZJjQ/B9RtuL
gGARYbj/4bo7utoU0zIMK4KS/gXtVb7RdUXC6FN4XdX4G66heRkIQAxi4HX6KFAo
YRMkVZPr6MQ76I+/dErdDq1tBKwR1FMBf5AugoTFmYlL6FuIY0Gqv7ScdCB2lbpc
ChoeG0wFnUf5zbdHUZIDY/XM2sZbSJDp284fc6+NGbxtPOaK3DzUPeWlcru3pbIW
/Gh0FN4LRWB6glExNeVV5UoSHH3NzXUm8OB1A0JdF7Tu5NktRdrQQSPgmq7m/KC+
7hdXRNL0Gu9SO6cFALyBtfsb84rh+4VVAEkgwnfVZ4dOCfUHfRjXt+sp+iKw67F1
gIUIgHFsNvigKHVrstCEsydFkP3akpZu48x+tp0mbzyeyt72Ll2tIL7rMPmXUc+P
EUbqTgJg3aIWtVvvhG8/rlZEetOSpgWaN33tlGc3p4z96q+doDG1Sl5eMA/4Ej3z
5zjJ0EDgb3tX9s2DrY0iNlWE3ZEEJZrUpNCOvbeM4UArACf8WWPSs9004GMlE9+t
xeigsTBPJjbHti+lg/25jVR85R8CEYCEA6roPFDEw4010Pz5VhdlSpwuQqIMv+Qv
dp6PY5xorp5pf7hcp0DN8zJzfF7FZS3xI5y9xgJhOgkiaU1EuqVzRA3ou2cmHCg5
JtyCAPd0TBNqnS/fYYY9NgmAjzPRYwB610W05xjgyIyb75hQTJpSoYW4J8bP2Qvn
fBbeemgZrGkr/LHPvxNmYsaJsiRUaL8Mh08vvGsOwY+S2I+buVEhJ7w989bbtpaP
q4zDwAJK/Mz0m7SAIPei6rjsqPngGMsofr81T3zqx5iJ8ArsrUP6F5eVoO7VvxhM
K/zqGfTOHcnk9mD+10je2sU9F2Na6BnP5hKuvVISa/8Db9Jn1AV5AxzYU2yEnomp
4bOKUTKJxMgcQmsLliA8i/KhH0BlKdNa4yxlNC+394s3+ExbNiih+mT0yYXo3XBC
oEymLQ3UUVJDOiEzb1Yp3iI6AHOrMS7Pav/P2pHx1bZPqN2AwsNW5XuSLETrmUJA
sXG4pG8qBUqjxs8f46XwRfGdJR20mMPREaGA6KhPwqToox9mbV+SKHiMt5Fe0YxY
0B8MzzCz8SH/9UHarorBb2Z9otAcCNkoFSgUSAPPup7Em/WEoHaKIBmHomEAhQ4D
DnrKpZ3JymmTiP3oXv0f/xRmmRrNbBPJXXmVIQ6Sq+Jiv/YP5aQHu22svUBW4s15
ym/gvlGkjw0UFiXVxsC7/uY1qG3MPfRW62TcNzUgQUIA8xeTBiB12LJmixWHQBT3
NcFUanzwpD8EMsMwiVAXDfP8NILYHfimht+dcIGhimWA1I33H1w+nTk0vBOqYp74
i+HfUth0QaJYE9XYvn9AGglMmn1wzFs+EyROK6WUnSqoJ0uS0x9aZvLuGDYQeHmA
f7pGrp11SPNKnxRPf5DFAqNN2T9JqJslHsu5lBoCLLVsigz4wutxQasCufb5t0gj
gvISDw13o9xig35y1Jkt4HnhE3V84aIeXcgEnVMPO8KzaaGJ27LMkn+ykCiz3tNZ
LOfTbJ4uNWMAil2JJZ3GGhj5gw2betwm5Pf6nacybKwdcw4rgTNAG9yLsR1HtRrL
EWLXUP2OlFUM75SbzukiiNlVrW/laOAAqSXl+nmogNKuAeDsYEZ75n/LQg+nAWIn
A+bNQOPEcrAx6giabbwMjDtZhCByFFuolyG92Gh/ETjrJf5Du29BqodZqcjsEzX9
d1reppqDOJuTvLTCWSfwCzwJu8T9VfOydyByNZdYYdcMtaWMLU1uMJQGUnkEsd20
VbOq1/UQvLCnyZjclEgBe87oGYKkjlxp35X/Bt6NBgHoc8uGKKh2Dxov3h6OkWyQ
UVK3i1omHJXreHBuM11WVqNc+1UibC0BoCCp/khgxpKcK7b5409XT1Kpf+w57aHM
AmYJ1I9JcfbTRSCj1iWSsqrE86ypgOax+clt9dTpHqzFpfvpyQDd1SRaM/rKfxna
fOLZYVK8v/Ismv2iQYm0sdj4wdSeaIsvhL25vS6+RCT9piTnexQN/w9eKqMpvhvW
0Vy/4bDOAlHBe0XDKP89wOvm8BkUpb2JgEnidSd1KjXiKYLamDAgOL1kYRa3b/u9
W81oFoMGQDXvBBBXevPsqsLfO6nFVlnQw3/nFdHN8ZnLDyGY2+jVKp4wI5ivv4vI
817Uh7Hj3ecNJaOLqYydFaqymX73WROg3vu1AHfpF47IflMmo6v8PTQRc8FddP2R
dKwzhy/fbNmsgn1voXDzKJ+oypeiP2Imbjw3Map1ByOskgokjasTOMfgFx5TR7To
MlKH0pjFTyU6R9o94NRCbgIQil+NYuCDGNwo2JSfE8Ue4ZJyQZH1JBojtDeJuysk
qiZAMJlVFML5mixRKeYoENgs2kPp6muieiCAe6m77x4IICxGuHxOqAp7o0St2fU0
BsGvTWxefbIM0j7U63BLMECLOned/MPDzRpGCPWK+x32ALhu+GHefDo6Qq44qTSz
fKmJ0GyGWtxNlJHQjuYG99J6FKzJMK+Pv2rcwZ/c62GKWG/futJchESy2eZtv4cu
LANuNOMfDew1pMWy38jJ4ccljrS+LIR3Ep+Eo8zESOxLn0nobfXg3I68Y7c/PXSe
NXoUZ8AVGy9GyGY2DzKhGxZ8rI1aO1erTa75vajBfiHwmcu0G3Q87nWFv9ZBLx9l
UxY5d96pPMZ+wikyiqtk22Z2xdKVouuGPIGCK8QNHuDBOn054RM8VF6wNQHi4ssp
eW5L+CrPL0/uQmiNR/gKyAomlr2HmvD7NZBE8TeaV8VAN7gxousbV4y6g5yAthN1
POef1IAOahtTVRwqiD/2/BcK7we+rgJBH8PLLgUkq2w0k1dU4wGoO0ImFPerH8c5
D2ESMHvalMmZ/hodnF+98dwxaeEWJAzIjevUzevPN/oj97mHnw3OnthF+4Ufy3Sm
wwMbpkk0KJqoFSDchGpmtLd8kCQfRfs4ZTq5Kd1jCtevar4QwWyRiPMXtIerhDhZ
9yxH3EeEHRRpUJzuhrH7USIe/g3BT5VJO7ARVufJ8LT682+uePxgRVNdHSqQHd4w
iPkm1jHy9Dv3zgzOI5ucdU/h1wmUN4wtFM0i+/zf8Lk1chRMUJ/ksDQDGBfwdEnl
DkXmUCHFfY58PrEQyOsQmd4wI3N9Dmdv5FtY1RFIWwTGTNcHOg/6ZWcpaWpFD+9W
ibPMlBmCgCTSuF3KKD+6sqS8WK4qPWiV0yCcWCOPyifs7XT+LIUiZGF0r5vXD7t8
moKH+/lXuuMybb4nC2RCToJVDqIHPOqUJMbQRr8IYxI6OLXNsDmzJM1i5bmZvLXE
srzr64fwOvHoNwihqkfcrpOSmFxEaQQwnxtYXlr/M+OwNmABSRJHcbCf8ySrDFmN
E3xS+J7cgXiUGjzB/fzTBQM30dLVTqAa9BWFe4cwdHxUdOAVARv/zpwAX6eHBPKK
9fCIvsFDvS++yE1rp7opbnORSGyyGR1opTrNCbFotL4yDJ8zCjsgF42oD2HDD0j6
t0jHkJGN2aILL01AgVXg4j0wJ5vlWEiCyZHBnzfPqJzDN3INGjuZHZn3B9CJNdae
7ewDh/8pBvbjda3JY9wbCVpTCw9PKVLzAawMvjfPMa5yvyS7KWYMSwWTnBQWqMR4
C12nPFQ7Ds+gk255nR48PKKwbAJW6APsgJbz5b2RuPom7iM4SFXgfrIdJ/pEzqX2
2spG1yU88nxBDH3TiynC+ic5VF/TqkdLuE6VBswdjf9IGrae5Dq8mJvCaQX73DyR
WFMkFwjMFPM4jqKuX9xDwjKHO5rC4RUe0aWcTk5tf+S+Nmm48kQoUgd3OM0T9/Ux
4edHXt/CFvUanFriPf66lM+vTeRaIo8EJQROiO74+7JK02g1Iq1qrERZCmecAExs
yg8EJPEin0KWt/FtS1sN9ZI7I3GYNoBBfml+Pte4f7qO4ywU9Qs13lv2+8rP1W2N
pw2SJHe7SQoqw60wWTmJJZOo26628F/HezYPlwwsLs4sO21+jbIhHgSNsh50rA2P
wsTSXorc/fyuGOV2EBAmT0bgQl5UL6NprSPa3LoOkYe5sgNhzN7lm5s1KHx7CbCh
dssDaH86eq06BXGLn9MkZMMRIJ21b4Q7/KCLoVmPrEU7ZlWcFkatkIhokILHXawf
OhvwNssxyrx+qsl8JGVyNPziJczHSvR4LlicgWLm4R8Z3lMHbCZ/f+2PacnwEuMd
QcAr3ylFT8SPgSdkfH+YuqAbzzK9w8mQOSdWj0ZIjJYkNhAF9p0CvVlozcPCiuZB
VpTOmK6BAThVTHhqFx6HXVYJdQ2wiC3NV90Tp/P8G4LUEIt1D8zDB1iAQsZeKjx3
axjjMSB12Qkm88QVUXf77G6igQOZD+HAe6NytcPPekewdIqPQDJF8nTobMNn4MT1
EmnX9QWmCCD6tjEN5BPGrGBVyioNImFlergPmN585aXGOUZsJGOrXPN3dB4vJ+5P
rPxOApGPR1rcOxjBSr7Z++ouDxUNDOBwOdKQe56FTT+SodJCt+pFdw+jxetESJ7g
3v02FjzJaLXQls3MmyNvZ969SqIzFqulSWUTgKBQP7UXAyQBbXr1lCKnIqLqvO2M
5nM17ohjmipDCYklCYBm9Q5TKfSKfS66TPWEKtykk6VDSYnAvnoXV2buXU4ZHQ4p
5LugQghrgsXhP6Ft2pSvGOYvSHHm5zeOMRLlBwuRu+vv15tDVpJO1vudf1HlDfGQ
4BFNu95O99vYljE0EU6L+SGV49BVGJc2pDCbsg3O/guYgcZ5C2glhALI0OQ3sZgk
tDvikYQ+sJA+StuzEqo9LZvIUkJpL/BsagPxghOYdDbqD+/5M5mW5gdKFquaG5xn
0F4GjmFFo2vN/2n0K95vDNW6mmm9MVEDW24xvIWcZm8H/BeoUUpcApb0mB6wC1uE
x6Ks8Dq7l5DNmT+Oqc/jwkYED/oHY7KnKLnHEhA+uoK+Q1Vzh4OZ/rpe+HASFu2l
UGLnCX1q69pIkrEYAbdM3+4LlPVc4ve9cajznXbRDi8nUxRi2ZDamN9R/YFHfnYS
tn9kw9WZx60NM8DKZMWoj4atGK9BgypF39gmLOLfv3qTbOqV8zO55KL6u9az26oN
kLStnFcGuYcpotffFVE4QaGYWFa+CEzuO1AEkYwOxtU7lXM5fHcxpQRF9+VpAfR0
H4BUtE0DAClxvTad9iK+B9fIkOKV52PBHMnZktw0OwDXmT3Cx+OQWZVkF9jzQXX6
03rMrK4i4N4iBSWikRAJB7JagrUCN/4H+I6Wj8rMscBv4xLR7uYY5qSqiekqqknQ
IRU+j0Fbcq9EaDIFHL1x+aZoWj2CApwYkd7bdQSwsD6TMUCmzAcsWrjnKrtHLA3W
kla1WF/5h/Z6pFzGy3CnMcHq66yqjzMhffasLqmZmyjmfG08DIQdtdied5tUNjKu
LfJcjei4Gdix8bKVLFO1iTgR+2X35AEf7Ugx25fSO4Rp1kweqElidKmYj746lB/6
fOcX7OGXiB+u7TMnO2vkMK/AMzTEhSvbuid5D+6qEKTWzVcqmtWBlEZt5FzAuYTj
vsED1dcWPE/8TS2OmuW8KODceEuMGg6XIVtOy/TQn1srhrMhrQeejaiVpj/lwFAT
xRWeDf1r90GHZu2WvY9NKXpCnnzyFbLPABXz7dh13rcziNGhfihy3EY1KNSktB6h
sB6zXEqp7vi1OTVtWFRRmSR3q4oTmZEjveGRJakW+sFVEIdig8PggzxbS2Ec30iE
Llv5WBS4sKRQtR9VkJQiS5fF3kdZYf7YiuaZXDfoCA5oQujogC3CqC/GbWwWHgi3
lJfdQFI7SZqNRERGSUJKXsWpDObb5wjhwCpn4FFiuFLyw5OJtsSxqWqo4OglG4/b
YWXKmcRTyFljtYFjDlurVxBju/1PYqj+OeIFrxXzo+0CKO+eTGTmbF56OUplAp6X
3ic9Ho7rpFWMPEMahlhT/QaX/091I6b7KGBtKWPMVROYh+NfHDdK+A3H6SqGqDJt
2BUknt9y1Z9MgZ6M5mHdcBxr2qmFACg5mPdkXJawwCCLo0cKppcIrzIpEsmjGe48
Dvc1aXpwBQ2HpSFe5Rji9gvIANCyEt0j5tiBy+MDq6I+jxo695GoR7wWO6M5bLNi
`protect END_PROTECTED
