`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8R1ccUsz1jILUzz/1MuDmxeXx14IzVCzN4DLfrcB9zrTm/LMSD+NWIyO176ncTk
zKtl2RWmVUwSK0HIOBzUPdypPzAjiB9NeIaa4x+x8RFDRFzft4RHS4V/8bIsArjj
AAac2COwvVbh3kQN8smRbWeQ2fyVwutWe8xsES1NCAalv78Tha3A6dXNIMcdgfGw
SJVPMVKhN9kMX67uVqiqq9H1rbA342nv9SYf1TLe7fDjqvd+w/ad/Nkh68QniorC
DsB69xv76RtD1F6S9IC+VhO8H0ELDavG7lRzsW7LnOnOtpdivZB8rHd5Cxlu09Ja
MzBYNDPqmAb7i8awpARF4q2ZupDbGgx6jGYkLR5ikcqkmN6qnkZlmlgca+4hAOCZ
2tjwcUExBfgw0BR1wfUAE4Ya1TLLjFviteo9f12qQR3WUexUAN+fFuiKYuAb0alx
y3jMP1IqpHZ/lEnMtXrNPSgWwEemIudGGWbd9EfgwMsAtBbhtMZa40Wvmjux63E6
8+KwFyfarTEmDzs2/TJEVg==
`protect END_PROTECTED
