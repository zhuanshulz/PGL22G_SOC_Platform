`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9jtLsy1XLfPt+kdj9q5BFenCfskuACA+zTiLhO7bGFYQTKeeAOXHRICiWe7m2Tk
0xWjhf/iUDGN4PmD1aLbcEzVY4+ebiGvYJpksKu2bbWLMKorCjBHxehzOxNVD7t3
s03O2i9QpZEuOF1WXCBcMIs+UBdWvuarfybhYh4adtnbmsMxCMYv7soAZ2PQhqh/
mpElZevl2puCcobujm60fr2K9pbQs9h/J+qT4rFfotdI/eiRF+VA89AUTucV7ty1
u9+cw7fWpVpN9b+fXqF9YM8Dtm3nGvMlGIVgjzHK67qBAo4s4A5zKNG109d/v1u7
KRyKmCuv3R2zubNiCSq6WFDJEqzya99pXHJe6SYMRN1CjDxqUZ+dn9DXEdYGxg2Y
eXxBgVJmwL2LYG8ucSDwkhWWaYwn0CDrKVh1DPHvPH4DWXh1IFVpypdGM5zKEFs5
E2AEiI9F3jz6Zx1HAmKpDoqwnM5XsbuNfrE735lSc6FqDjUlZzwWn9UvCDFc4VxZ
NtdRZKOhtx+n+JcDiYK5lk8+RQzuitLsaDMTE3qSbDuhK7fQ/wAWzqdYXl/dXeoN
n5XP3UOgfdXgpY+POD52PYYuwtM47ixE1hGqWQjclQ5x7cZSl7qIQA27wa5kULdK
ys2kC1r+Fky45i5RyNVocL5U3quBXVW+ILS4g6l7UzX8LzexcQT5CU42A7ZqqPi3
i2RMF97V/YKlHggehUenHpZ9JlYlPK90Jm6DfLPXrKWbsMExLc1dciNuoxraEX1f
ueUheqcxZq6fBS9J82qvn0ouw01TMASwwVZy0crvJHbdDYz8vdL/AYUXGPwL9Y1f
FmRh+GE8F5QIiAjD4uED/S1y9uZOPIQPMQnRHghoWmF6CSBb2VqC+o+/lleqLfjz
ngFd79CUYO+cX6ETV+WwkLeHNRsHOBd72Z55J1/3GIU=
`protect END_PROTECTED
