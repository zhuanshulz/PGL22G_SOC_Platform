`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AoPl1eqWJS/q1yChMtTsWBBt7ZH45bN4syBtDQY2Kb0inF3rZUXdyhEK74hRpZd/
OeP/wTtzJCtQX2f0abH3t/B9lhQTuK/iPqVkYmKrXmQRUx18F+7GPVTz9eE7kNM6
S0C4lGo1QeFRtzTjNeFHLl4QuBifjsaPQWm+73Q9WMm9t75SQvF5h+0rIgR1iI26
Hg5R0r7hbnR6S01JSfics32K3WD9z/SyltFBA6VzpjiNW6S+frYlkf9RmkpNqUeG
28hwj7a28xMz37nn7+LRUPheaIUDJZ7u/XP1xiHc0CRLQJS4wQgBAivm9YExGfFy
kAO3gClwg70U944tFTNtKyf56V6drYOoBm7D3hRHLmUuNIDpTPdh6WKb8pfz4JoP
9qHNy9+cp/1iBzDlhlX2FM+PZK4m4zQEjCwYe3ziCqj5fvOepuqnctX/CbSNfAAJ
EGwBCB0lQqf4VavRG2pxqTBsGlWfC/I/a6UokLz6s6Y0vUfpzWn4eJY00aKYyLgb
FD39nLwy/P9RGLmwRVd5b5UmSiS4xNjyu2iALNyQEZOgJiH6lTkBc7aluR1GHzWX
iyXJCpebhSgOCSywR/0zQcYOwPjzP5YsVneOnfvDPTMFcVsmKbvhqBeF53VbLxKq
da2Fqfepkh0pIq9s8OuFYTdohUgduVbRj2PeSeQqHGT1iUjgNhmsQ5R+ssEIu26c
5y8UJx967u1N2ysOE+3+atfaJqsyevqNSbRNzGCiWuhjQdj5sMmeDCAVgImCw4qg
sSlowXDc+ybTrLc1gjrfWfnyVqjJwVOA9LtPrBc+Gtn4l5Nj7a4LdcJMaGF3c8pI
XVSM67Bgv11jgi3UPLTTpOqqXcZS5WT776RoB3bcW6f7paQMf/4jkwZKMzYGRfhq
RgQ4FMltr02WPC+7z35jQJZGszL0IHdANmumhWAClpd9GMHbyPbCgK69Q/Vn7X28
SGbVw9LRe1tKDCOs8QtEUnlkulshOboADKCMv19NkgqgNF7ZMi2kam1O/9aYqeEe
LkxWNEglFNmU7YXXD0QyHsjIEf/tjEzVfqd0dsfOIg2qvSUAcAT31qs9+/lwfsCP
wUwxfDotkIE5iApgshc2sA+SAihA9bKz43nB4ZiviABPGingNuJUuE5yShZ7x6RM
8MxV3THo5fJQzBKHTX3UwMw2fImpdrkjfS0Rm5uSDoR3CNYr64Y4DQtHJFpZVbJs
UPTbUwSJL0Lwg03kAfiiSdZSwnv/PIuaY9VTScdODCF5g3xBbAozF6tY4GZ8laU1
In1zQrm8WVLjcFJrSW2yUecArdwUPG1gWd2N48Iv/NufdojaFoT3g1Qg5Svy+YOP
rOwJG0S+jFXVRSDyBP5zL1IMpUVX0hAPCY7I03A2vb9Mem1lPToRzZqpEIQtYLzr
rMGEjcRt2BU6aPD7StJFc60Tcp2vMIWrkIOqTSJNFi4XWMQFJiK6x+bdayGt1qcx
+muKy2I/KprURJylcZyBEfpiFwaBO6ezBcptMJ/PL/B+ViLqpepGaU3FWsvN+aOB
2G9dRPkbLwoQ+JBNdzUW7Y3o7dc/Gca+YQyg+qRftPILn6UG3X3qd+9dLp72q2Ny
`protect END_PROTECTED
