`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNQ8AdQ+d7QMdAHuc18hJbooxu8kKBxH5wLfQmJlsUwCZYyDeWLAdstIyGeylkJt
WOlqOWF7ZG/o7DCBznI57HOeY4xXxH/ee2PTri5LS2edfcd1qQOy8ZKG9Mvs4/rA
FftO47Oq1FdlFejTsnCsUYcXTKE9qsvofk5fWa8ms4U42iTOWrIrEDNtoSPKHLyz
JU6byQGGJKK6DHIvSgun4nhUT2FGWwiatLlp++HJ7DA378ndQo7dT8olEMsx6dZp
E+CbeIh5rIqOn1BpSQDHHTwQ9LdiXm8eRnR5A8Ufhkpqz2/p2U07m0YFy8hj+xdw
Vj2o5DXZPMvnewfUFvaHKGYjS9RJkSUCJwC/A3oxPyGP0CaYF3wiXTC0xvyVepk2
OzfTrI/D/GrXetjsnFtK8tivLyWPpg0RHc/SsD6k/sNdO1fUViSUDTWg6ttNCEwI
dbH6tMvE/sf3Kh/2INslqPSqQX6n1Qr0ll51C2rxaAD5uLjfBi22LoDjvQuFNmwQ
i2q0jiEuYE8sQMPdaeov14f/mIs81oMY2axVKImDCI7Lv7xX1F9/kTZqiHx1KgXB
y/pd5EO1mH7DQALHrhV8d4Bb8aAT+VvMPUcfFYcCW32uDD8tqjv4LrDt5XfqrODX
TVXHUlxbnP0f/gexXAV7RfF7QgQ4zQsvoWjG5FR5mNr/qERgB1fjik0tJEDnljr3
6jHO/t5wa9G3K8UMSVe/nw==
`protect END_PROTECTED
