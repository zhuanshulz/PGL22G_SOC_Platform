`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lyh+T0UZCPGd4vu22qlvUbt5tlfJuW06+G2wUThmqYU9t5ymBmIVU+HI1ao21exY
4Y30N9h4Ny5ploDxUVj9aXWB9fD9iT9XulFxbfFKM3b74HTevLn+axaqfgDiPJtE
f+qs/X7JPkGSLmZHEI9pZFGb6qi82q+teygfNxIrzfAJO6XmaNDmcscaNXY95Vg9
n3TlFMG5cFFxbNzHGLFQq+aXaORKyQ3y/QPvF26bcVR5fQeNOWaCiuyXFA/2K8NQ
CVi8m4W3S3Fx+cpiwPiCwA==
`protect END_PROTECTED
