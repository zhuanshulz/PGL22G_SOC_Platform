`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DwpjZV+7gBpzTcwIz/aihqvy8OM7U68/cWP7jgdJCWcC/d3CI7AbBr/A3Xgs2JcF
P+v3oEP2TWhQfOjDexbCLuikgb3soQXZw4DF/LSBbXdawqtGYx3VzkPJBTtEAjoN
TjscpT0AHu+qxF1ujxTtYLUKwZFcNyEo02vcSdrHLtGP9VaQuqoYC9vtaJZ+ih2p
fWZj+EKsbMRW7lA+MUGcg61uYbu51wwugRVmQTT90DmFIYq47I95zYw9kguP9K3C
d+MaQafv1h69n/kkoVDAs0qcidYJlIDhVAygErN/CV4qBxaKk59cRBIk/fjMeUFK
12xkirHp8cj83T4fqJ+L/nHWztHe1qsTogpLp8PGenql2E3uCOMsNpw7THpq6eWH
epWMEGatNUkIIAKVfSZ4d+eKfTk6jL/vzqEDjQ+3JagbBfOcuW0W3ZWvvat8uJds
fTivE6hxw49A83L0zWrk7mW0cqOTwra625PUSW/vwau5ZnFa+bTq4wzfns1/3zvD
jZDhXrC01R/CTrxvsDUJew==
`protect END_PROTECTED
