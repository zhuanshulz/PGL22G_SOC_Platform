`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tbiU5u7/KA8rLIrF373nPubEOzI77EWdpUxY5BeqRVK2OSN5gSMxch6V6Hgy7FA
ziMAm81cDL4PC7JiU1uYoqrTcOUgBSAsY2LDTMZfKJPKuOOX7q4Jy8RILIncHBwT
uLZ/VQOnaCkrftVY67MJ0HcVYU9daiFwPScNwByWr1IcpC/qm204RDcUDZu9LPBw
EIwa39kI1kjq70lWFiGy1YxZtduUety1laWGE5qwOXjVrOuQWn1YOoU/pUtb9cal
//xrCCb0nFObJiRU8OzfxEv805W8mSuE+VEp+ETraB3j/TBWVkRpwz9R/2uIKxd/
MIuSTxn1gNwpFG5c9AZE8JZEVIXBNOr3RFJKCjjef5gHZfjO3ak8z+zkVz34Smqm
PbsOmaTdB1bWtwF4xckhbdCKDdMCbBwIujdpTTi+L72NAk72kDNb20lHqbd/qQRO
VaBKKTrWP9/pmYcCZifDQ32bLnrHqeZA3/EDB0LX2jnkk9NqYMysB2xF6q0mu7k4
omYniA43sQxF3x4aEqHlh4d3pmdgfDEo14dhVTQHyyit09YCv19/0TuS4qFDh4Ju
6h4MEg+qXTi+/v4k/5oIfzqfUwd1r0SkfEbCKACNCpPiH9zeNsuHx3ozF7jVWxQL
/i6jbHwU9sCArkkb8SFj05oxAyrVDT5+KYeZNTOJTdabyo89+YOxlkanSqKufPDl
vLN34vFW7UO5qAur+mtetp04Z5rux4UwId5kdgrvyXzR+glsUVLlTIRmjK6cHcpf
MMnXTuvRWGy39J2lfoNFZtMKCvwj6hpzMYD2Y5jHhJAmVwcOv+XbJmyN6kfZSa5F
9icBiwD2G+OfKxKMVWp/PzhByXwOya7PTKAENqsu922drjND66WNPpRT90kYTshg
z4F5vgkOj7MKEiMXbYhD+oh7PVmOe/M4xjixz7O0F9kyGV8DJTliJtkgD9eRWZmY
IcGJyhObUDxOiKLU2T/3Aymc7ckRpGx5lKmTtju8bte1dHJdye46F2z37bDxsfjc
`protect END_PROTECTED
