`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/7y0qQFebP6kUJ/d+0IJbYKZ6Ijbd0amSkqgg6RBFTa9ca/A/7GpBty48cSK9dt
dk/FxjAuDQvk36OLsWYOvTAw9ghhuB5DmbpezEt24VQMlvNHuZ7R4qNn0CTyzFlb
g1BZQZbMPnYWOC1qoNDZ5uTzDJz0fYZ/9ZCVdYhvrTVR7ZEzSI1BDFmrwuwuJj+W
gSEI8EnM4Xp2AGAUsf1kwkdRNWoGmvzapeoGPtoCV/8ouGeZ+B7N4hW89haIr9iO
mPvK8iP72YWE3HKvjs2YLJotdStyHLGQB2ary9SPoP/c5Wb1U/0pvRkZlEGHGbYx
OGAXh1JZoJeY0oaXPt1g1pgjYIi/nIv1aaYCDCvMXjg8Lk0K/fAxpCYYdFngRk7z
6e37aQ/eiftd4o3g9d9qe3Jt4Ajs7/paxHohlIL6nqnJrC2tPq3Q2UnCYJSA0aVR
aSehiXSv7rcVHIZO8zMcfx4g1XFMDevkd2RPJ86v9Ly0Z5LQcDObSgc7bvjTmurV
li90uNgeqJvy2gXHEU+Vvad13JD4PGqMZlqYk+RxccY53m6q1WgXquwQOEgEaMoX
bFzVxyZWEbNyfoAaBDWa/dqCoUaZtUIy6sE7//QvgYSGv+1Joa9Sid9h8Dw4jzWB
uffHlEP4WTxw8JVx7o9MvvSOs6BMEqgASrtq+NmX1xnrPvPlmmSUQ0R783+c230O
sh6GR9VRGK3TrMGY5a/8UkzM093yfCp/HUYeGfZ99vmQov0r44dCNCgMBTylvxF9
NLlMEWpdclodKcOUunHRl2a8VCPuzxMP40Fwk5gINxytWP03ZPl8ICUuUtmPfm3y
hJ1QELD/3oSlfaOqsX7Z0GBA2AVG321Yd58oehajVbCY++rqLcBWnzYimMgDVRmV
0ab/F8oZnqfAlvg/A0H8IAVHMVvfp6bjUjXs39geaUa1yGIyHC2h3mpsC9yt8qDb
xzHZx8Typ8NIMTZokvs3VolzBUkl5E4xsMgRCEh+oh7+fAwms2SQZfyBy7osQGFO
K8kB7H1sHRKa0UjueHEgrrSscQJq/tOCIosM15xFVs3MoFWV1bEY7MULsCjKzOZt
68G1Y+bRqpFcrzsYIzUlqczW9L/is8J9cy58ZHHJNoyk8AW1rI8fGAHgJwSj2/3p
0MBLQUYRqoLWbvlVugiBDzfZqiGOTa7xzzhbxjCUbHyXde5m6JgkLBQHVEkpl+nj
MhvBbPoFfYQyHcuyXE3pFMduMDMwEmNAcaKaUcdgNMjyu4ffBa9HP5lcdf14+yZy
e/fUnJHG+HvLMPtWTOpsasipLz3LZXN7g4GNoPLN+ntsZfE+nTeqkbEhAZgOk99I
b7ykRrQOs+i3esAaszL3R4bRtMMQ+iEPQdS14laSTbe/d6Ur3dEW8EFJiiMTxsSu
ccKQvSp48Wv9OLlBNwGIQ3xrnmrNrdX1AZM/h7v3rja0V0GxBa5mgLsLGIeqp4oZ
nCOM9c1sHs6wWgPG+6KJs610Gw6IuPZt+VNYG4H9ZjU0rgzAjajQjDlc7kw/qmh6
20ZhVYxuyY4x+o4NN+7MMlPT0aPP6j1rrQbmm0C/fScTFTzVzJCLDxvf3ayBMr5s
rTkyZMv9mZX4R9UlAFZZ0rohR0WBn2DZz0o6936jjl5BBRytWIOcD9H6aqRHwjmy
wq0gtbZoStX/ugSrrco0L6GlP4YAeg3OcmuJVLtOkoQWD6QenxzCoaZm9PFz2fdc
XqtGIxVoB5D87Xa6nLRa/4xW7D5vI0g+tUdWGR92B+vftNy526O/kTXId0dYhzU7
4/neD+/NSVJ+epDrE1rnodJkOid/3e4c9NxJBr3lMNQus35urEmIpClk33RVoz0W
SEmwJmIjmkK+uKUEaE1ryqpvhpZ7BzZvnBkfGseALuyIUIjb36WzwrcA/EUJDgtR
s8Sfrc9bYWImNFDgu/Uyl1zfuxgs0HhCA47MSp5vaKjoAialhfCx++MjlFjIIfcP
tYRnN6JMP3y+JiWQQ8Uwt15OrOXWQI80cEUQHTmaI2WX30wU/69Lk2C7kuaWx08A
pQKs8KKq/ala/jQmEAnEMQ6GzZXWmQCISG8inKpB7DE/mCLEKXYx9/5ojmgvGFHa
VPwCgPzANnM+ux11CC1j8JEMvJ8d9sMf9EeXpPOjJUCuCHkrRDpkruD4GACZyHcE
m6jNLg0qjCkx9AEmT57cBed6XACW61n1M5xRpCVnMILo9QWE9UO7rHV9o1Vkb+aw
OHyvnojtzPCHnzs63T9zoTAPdEPvrZy5asfZYjeIjfRAUB0b3igGS2tMk2WgAdv4
jir96Xj8KiMgtNFzMuQdblS6WNWkXeKudz6Q4walwby0omCS9YZLMeQx0szgVNO7
kAZPbzUX3hj5ngx5Ktj8/1tSrxz7BxlK0F6ME0vnmgWP0rpJkkGsATyH0gLxt0g5
A40Ko35WnjCgfWjvUt2XGpYuvqkit4OrcLnuKHjrsWfsr9P+XrPJZt43Kvnyd9A0
5ViRSiOzdn4+rWOHe/Hc8kUiV75njDYtEvQHp/76cPrSOZ4KbImOJ74eRrKxbXtO
ZUSv2+TsrkQVjGYMn6Vf2wOU16OjX4H1Rs3m6XuRGITHABYDIHcbVTBVbMYfhHYV
M7ooJ4Afz916BJlLVfUCT8lC0XM4umHCyvP5aSlsHAn8ST4w5gsDt1JRiwfHDTgw
UCuFkb4wP3CHokd4g2N6qZsWpYNVvdhMvxcE8EhQEasA1BOvFGRIaXH1zT/+7L+Q
AhwAQwIoZGCo4kZhHmNv3T6JJWJrZ87jGdvDHMMgoiEpqBSM39oy9R7QLnXuSY+S
3sfrQww0fg3I/z19DsHvDmgU5RJKxb2tleoGGf6g/Uthkot2hiRJ/YaiaAemos+V
/BeUjLZDxhORSo+3SqIrQ6f+v+jccz6D199PVa1Gp3Ovyb0/QgGMxC8otlse0lUa
9VLkdt55R6pY6vtAoDe13bPhM4D3wMIXW9p/7vMgX4XuhtjiJk/Lum34Y6+d3N93
66G/t+03A9G+wmlyHceAf+K1A/iCyaLKWCwLEHmwY2d+Z253KqIUpawfulfuBHWJ
5ytB2kimwz9Kj0tLW0C30bWaNJaOquk1lhPOi7bzBZiAQYtjNkzmbscM3SLIaFAU
16V281SVXvy6NUdjOZLyK+ymSbUC7kzauHYJQkWq+S8F8SkVj9dNbimiNZz4Q3Rh
JrhaJDCbbAueE7vjd+vaYIUQbnhQM7Ln4WXjVm1cBy8Wkn/5QeMNOD/lArWvF6bf
vt4dAZA7i0eqDdrA1bWNbjL/VMs89dUmYzTvGr0ACB7a3CMDP/il0RWsnBYPR/mD
pyAvjpguem7OLZ+0Suv7VNMr3hCvcIug+GvpOWyfek9Xn8CmSQykuCFBiNODvwRT
/8T8ixYH+f+QIeLWOIe0TXVml5kpszQQlsPl3y8OwXYOdcVEXkTYavussK5e2sMC
MtIWd0rIfGqqFjAHl5oIctCvWo9LElQzIPp/rtOOVvbh6lwi8LyR6xFVeapyYj+n
202oAl2xftYnWRim+y7J7F8BCNEjHaQDJh74GnC6pkCM2pV7IiyDCqINGyiEJ1U0
NOPl8Tm72QLqW+2RBWrnodv4JiIXw5bLtsSXNUkIlj9A811uWCanqLuNumPPwK0W
UTLwB4nLneAQRj1tFmVnk/05tjVDHAitgPPJRXygZ4GJHK3OD1b5uyTSb+z+xNaZ
jZyx7B+UnRRyv3d/LeuRC5TP/KEEJlbVcM1GYN0DN6yWj5WvR1xt6qhlbREKzTS6
MUL8nOw5cqQ/r7JOF7gFf0BfHtwSkY1PbLa0BgwiV++AQTR3K9oPI4zhAROjqZLH
gGrRlQJQV/HXIBHz8AfLjLR45PDC1fVKRPsgNlIMlB4Q5fD/dvy2OuPJlbweE/5W
mJym4uUU6w8iYjff2cK4BUNZJfXMbbqnGf5Bm1BDn5uIRRvxzYCklmk7yMHz+FBQ
7hEPngeVmc4tKkn2z2aup1Ci29aBxAFqna5us87JDgLJqjMiYpQ32dyuDpLuc2ey
ef6+qoeW/UwElcL3Rz+LCrsUgkCye84DzxuZr+Yoay86MsFUc+ScvDqoDv1U7JFV
ZJV4MJ03Qoyd8CbH9wWgLv4VfghQ/p6jW9VJ9yNyzcw0Zfow4SK7iAg9PHdtzf3C
FkSpBB8Diyl+EtO7G+AFnwtIjIDAWMk23fIebeea8jzeAWIly+NLYoX9aVAMqQGB
KJV4pgOOqMEsgSnG21JqYUh0iF0H0PZ2j6xjsthy4HxfTkgHt1p3JFivBKTGqdYy
4qnayvWuaCfvPTbp6Spd8jxo1HAnZMlarAUML1KqVkhqJ9KxJoF8+riJRntygOiQ
Sor2bJvzI08cSNXRkG5Kb+qqNxnRzQ1IvxkgB+pdsBWeOkjel0YbU8XG0yoUArUM
xzNJc0NxM7FJQqb10N/SWu/y2FX8CRtz6vZ2j2M845VXI8kHsO6jA5pRJGk5RU6Z
174FPY5Gn9MGTcDAI/HqDM+SE3+BNK9Xr5293I5ovqaX9u2GWOqThWNNWjGHvN8l
kx77pbQil52TACGDqOFGCQV/cie/oJaO6s04KfhJmrLvM0j+EJAmch2SWVbeoJdZ
gajkPXCZG3QpXiu3Xp7Eb37jooGDorWeopkfmNJQ3Cg+5pCu91WvHBt3U8e7Xrqv
G6PLV//AzNS7F+oYsMjSgNbYpzm7UUFiZ6Vh+E7q1m8PwJuVjSsrUbw23kJ1vVSR
lp+EE5ZjX+6VSiv4iVc3UEI1hkeZ7AM/CQrDjqt12VxVvFRNjld+8aM+7jh46+g0
MI2SAa+VWXlZ+4AK4OGmQO2PiOd6JlHTKYeJoEkpML99sGSvuOGu9zv2uwkf4u6j
RDacGSBU6V9mpLvdI3ffv4ILqoSG/jQgeDJ02dtEvp7ka6iVlZ25MoGAuXqfENrJ
ftVkSQHydshqQHgc3JlXU3vOTveaX49FOcb2cQy0tKF27hXc9lxDbfWVS2zTngO5
ct8tDvOe7WRN36QFvn8Mi9z1zP5lY5qAlrHfKXagOfusiPNd1aAyZkppEV/zMWA3
0GT5LDnwoEMQxLlsFzxqjrd+GrdKoZnOZLySD52FYBi3LhD9CVTBg1qQd4iQTCsk
jndIOHTcA19uBXi8BNHT/FGmM0NfzdaqagG/uedJy60gP21ZxhCbZVPmwhRw75K/
ciZaOKQQkiGFQEuwfJoalT1NZ94J6Zdbhmrmwy+cg+IIhOZNjtFoGsGuIpyfwvnI
Jhlg3rH+nLXdP5Cn0TCIdy5SmmZ7kxHJaywGL3PubQBn8pZQJtt2ZFn/JQn/svq/
PyANdKo4yHjQvU94olz3B3E4rsR9SQlJ1haJmxKwLjQAGOXwrd4kbmM7kF/K9XGB
Q+svybicF3SlQvOoFTBtFsZg/ibo2bLxlBkBov4aPwf+hBIqraaoQMQOTMxdw4gy
X21b+RFf4PFmt4UL68J06KMFeCx5tmKBOCnm25cV8ARA1EAqj3H1xgxRDoaP74wD
c1cywUTWkbs7ItqtazlW56fzTEhUeHBSToTGw0YA+MSvpvcGo+S51d7yKpGUKOWN
GLLhtc3QCqfajzRsj0QtbomD2+UbYsxhqgorgnmy58+nG/RkT3oSRutjVZxKZEWM
dMkymFXFLHSKaUnswgw7OGLOwcRmcaJDbAPygDU5nTYzjvCk4v7f81s0Eh2zVZO8
Y8h5fOh2OjlMkpVzFCkontALF2WR5OZklNgDVutn8Li5PWMjwfdZZqLswJNTkduc
l7NADMiDQ2cnW3YE7HWrppNpsF0Jlh3gCmYL4R3zB/mNbfkFQFckY4PwhlFs9CkA
zHTZY25jenxq4fHAs6cfdO7jnp+MYw1ayES/mw7/fUD+tfSXryM7Fc7nLLxhkGUL
MRwSsAgHdqjcbK/0W8rIpVTZg10o9SbWBFtWV6Nbs1mgbfUOXd5CS9xQkb4lkHCB
f7C8I9mXXOTzude9IZzJzQ6tj3o2RVJ+4OG/S0wb1pldfF0f/TXz0b5dU4/ltHFk
YukogroDd3iV/Iy/6ovVdTbMo62bHdCiRGEXl92dqyfkK34o5fqAje+h401icPQX
351icxuIfPlR7BbXlu5/FSVXhFg4HqM4h2hpjP9TcAMVn1TLdaTCEgge35yMA5lE
zyA85MVW2/lS8bFEAY6rBkCql4rXj+8qTL/ocwumRJxpknLQBYliNU1hYaN4SkLV
8rku+3OsSpb3eNsAfKiMDrhoVb29ywgyPzTzvynSdeDpIoNrKoJTbJisSduQIc6W
OxaYzDbYNVlFUO2la080OP0sfviinqJuq9Zs1HF48y5DWzLy/bftmk8ZurZkIB0C
Uf50+7V63ENW1GHVDeNfFQ/JthV1ymk++Z3zfK78DwA5BPZ73SU8em2VazQaxZIc
ykTh4V18EJG2kGanCRB1BclIWsxZvu5qkdgwk37z3yEYkWU7tzASCz/9T4HytvP3
Noj9ZFVsNWibERMp+In3YCR3pGEZZIoNSaAW6SXBlM7Sn5HP20220a3TVDeQ7iec
rZZywP5kxGnSl0/lVhPRhx04BMPRzafvM4APegbXIayU7kBaAlfq/lOq8+eUU8Cj
hNji3j5aDN694jW1rrFQNR36DsGJGsYgpd8tDO9BmMaMAwBRcj2BLY7cGN4ISqoS
yyKVyKNYqCe23b/kPN7hYxyBs1m3dvnGxFmstax0sn2W5YmRXwKfJRIR9YfdhKjJ
q98hgBJGGIlMMtl6GvUvrTXVndCf2p2tq5qcED/IUNjHo/8OYWbv7K7yeF4chh08
5d1VGKLqIXU4kpq1ncbyNgkfC51x0epNi8siSNc+JZDZtd5iF8A4sZY78lZiGxuF
mLUThWDO128c6vaQwoBbIJfbtWgZujzHsAIKqOtda+GsN8/VFY7hjmgQm31ycvte
Ya1xKHlSXq84jTxUIXyaYrLoBytlAOZw19qmw4/Hdnhdix58HbROjW70FgRTabqf
b1O2viN+bJiBFj5hUtxhDR+adXR4AzeTNbL9brjhbHBWwdLsD0MgQjftdl1y9thZ
0WtpBzMcQz3DCAImezLi3thXPIlWF5qcgV/J6HjVe4trkRYRAP10qiCynnttc/2Y
w4JJJu8Sg4YetXnyN+dkRq4V1nq79tviPD56KO4z5DJSgSNpzoOt3lAbPXAmLSRD
ARkSXAtXhGjSvC2w+0cNaZlBDwCSGVJX9CnRMXvVcNWXGf7lAnq2ZCLdQieL3iJ1
7QKT+SXxqQ2SIWa9t846DjAruUg+qVPnij6MEmA7V0Dj7yYJ3DQvvPruFa3hI9Au
2ocRjQW72JsGbo6TlNvyvrvDx7jqbepRVNmISLol7YeOY/DQHeiDcWHvuGaxGsPG
AXMQq2OOwdjbxGWx/zdj/MNSwLlgPUDhDVjbrkqmdHzVOJWIG1Ov+mvOSzTYp1Py
pq1py77tPjgfGtyQh1qsMUILWIidBE9/hHrChYaVaoEVFVSgu4RrXYRZ5FcxJh5J
mtKKfhIJALHSUusSUsa4sjk53groJxW5H+Sdi143L0mLJmLQCYzO2cWO1yXFFN+u
ndpCvu/WaGv50so/3Kip2CTcL1IvJOtJdLjk9INBwxCgSLJNX/zT+0t707B8Dhdy
2yizI7hF/3gxeD8epuIYDA3ye2GjQtVbhz37QuwthYS4Uyk/5vcz/oyo9GGaxVtT
zeiiogUSAljK9NQlEaO9m67ZUXW/cqN3EUH2Ig3alkBYFu+GXhlQz0I6m4ewhgF9
ygVhNQXaTxRBKJDin1PRfPFzRERp8ncaTImByDvo2XrReY87zuFXlx0pgddrBRsi
yub5/Tceh204x0Wj4r5leGhfM3yK/t3dHhnifTBXXl0v94TTuZ/JTUf6l+jyMSQX
MzczAhmV3DPglXtApVAzhrDFB0/l23YjpsqeSc0vravY6x68y5XQFlUoTfFilSnH
FCcSC+666yLVoaWWBIOp9L8ONW0qh94iHd18ZNCLy1Fe0nd1pWOzLXhPsa2bNT8R
SjRjp6GJnCg0dWrm2fsJ551oVX1k1aJippGRSelFBhKpD4BS9GvSlW+czdW1mNKj
ivkBqC2f9LCIksSwHtT91bhZYJNN3RGzkEheq7lgC388rVv9Mgtksmh5jz+IEhOP
0EimiwJUnfQNyK2KqtzKxyjY+cv6YJPrTTOX78vGJhFH5meNP6g7w8Nhq0YU7/cw
pqo4UwJrGnC7z9awngYsDxiMhi4Cq+JNh9GaWcf/u38S1D3VwArIQxTu+BmG/Kqh
ZYr2Tc8PJxTBJiBZat9J26xc9ApbnLkRjxmVMZ6QiaxMbWMxO7Z+EsjH/uG1zf/k
p2aVTnO4bbb7MMH/6bf670K2wpARVKo5XS/V8FU0Nyt93NI8pBCsv2v5rA6gQ2o9
Uyk4+F7TP4yBJH/x9zFFfeLF8yV00BF4PC2ptoetuFeTinyG5/xQMqOYo5h01jH4
Vbt7a9vYj5yu/kZG+y4C5BaF2zEiXPmKiUnkSa/fU5Or7Qd4eKvfkr5o6CIN2lrq
jyjH0Hm1TcWF2ioXcHT6zQM+lRK4OuMGER1Cx2FQ0MClTqiNf0Slgez385KKRtG6
7aX43w6YbOfppUo1LLTFIiSnHbYRvlXrodgxafZyUsl379u4lwINNG4bjh1igkgh
WZ3ZOodcyrjSB4O3zzko/G1NjjvF/5ZPFduQLfgqL6jBZ6xiTpolb43vmmdmxJWh
S7aw6VhyVzIT+Lk0z6D0YFUQG0ch2eDJz/dKTz2ymXri05VSpyuMWcbCZh5V9ZCG
ukKK5EgniJzObwlUy6RJgtiyNqnKzAPKg5PrCBUBrVqb/UD9Q9P3WbiJKy89Gzh6
fQCKxG/bmTkH/vejWSKCd0p80VbJskk4IiuMHuMDy5GZGQSErfPsICjZIgrcCqaG
6SKz7NPpdDs06z0yB5yZPCRbWNHRdpp1w7wF500OyOru99oOm2mz2bgdxL8AQrpG
U/QSjN9lgpY0Am6uDDlCI1VFrnnvMr1whErnpPImcthHd/hKTeNLMlKbt1QG+XPq
foHG3kWj/7aoS4EKPlOXSlqbVMLEYtxe8LWvLmMmwGw1nDV+olpzNvkpgyGB0+jm
RiyIEI0/myVhQZhyVGYYRD7ATDjlKIx2e4H1Ys4BLqPmXS1849qX+JEgWOLzoy9k
4K0pptfitjo0HHBPrxKRhob5bHJSR08oSkqlBmk+hjuvI8G9NVgY3yxqtI3fIN60
ENSTWKMTHJuG2eZO24gyKIDVx3wdcWT56eFb0SbpjVoAShM20xzX6dBcOzKzhQD4
2ve8J+QMMjk8RdDrevA9TekTpvFZv3A7tB8LMW2qoB21jfJfcwVKNdSXg3El4iP6
UU53FsGXwg+1yJPjD6030aZNDEC1bicOAs1Us7o6jHOQAuvo1VhRiIhyB1EKHPbN
dR76+g6TtxPH+WOpVp4QdcDvrfv9tiB6YaztMV2HXdfe8arMNSziF4gkA+3ROwk5
/CWz4hVXVx3JOGKFTNAwAxFWmNjxEQeIxo0gUYZxxc1gOLHpkCgCMbYvuULj0AXN
J/y9Tjhhklrpvod5xThvlh7Y9S/b96+5UnECs2c9K6su7nwvkUjXpwcdsYjYKG3A
8LDkDJ3VnXxmujMmXo1gSZH3IMxHLs7O3W+FmrBjKHD7m7wv5TK48FNxdsGrErt9
CaQJlgdWru6t2Edq2AxdMOIGT57c9a+o0Q2IN3cQ3B87KXWVjNkc9+tXnZZCzIa9
ksrcpfMgvoN7Vrjv0IDqfVue5kFiY2dQueminQVyMhQnPyO3fBch4v4SukRuPSv8
yiUm0J4IQ95X9astt+0avClSZJQ6Yyxe4wpfVAodvMRGl0H0/IPyMn8Q/1Ew+qtv
f0LzeUikTMPVyyD3n0DwIxfhH/kScRgIUXDBMXvw2I0jGQkm7DOkGYskeUcaC3F/
nfUO1CRXDcIR4br8dx58vsiDihf/g6aSwWurEclHKPTwRZ9tpwnZQcWOW+uyUi+A
zo5gZ3oix6DhvOajpO2cz/RoEnXAf63NHmDYv2ngyD6LLrjnHYVRcaTOrNq+JnTU
dc2fVNEta7eSEYWMaVXK7K6G0wfWd/cImz/uAoGEyH+Qt7N9BRp657PEaLR6f9Bs
pfI1CS8B4nDaBiBLNPKTMDR9Fc9O69GPi1M7368TAfTo3Qvx61WLXCwCCBwVbEVA
UXWTT/ffYUWip/JzrECSKz8Gg1Lef0MJKJPokcn0l85rAnGEq14Y0YKssNcPWc++
6BXHjhGoP4BWPGV7XAciqaKLA6K1CD9XgZJGzG80DavAp7lGkI2WgUxtkJwdjs+D
KPqYWsUrQBelsYuTCiKIA+wqkX8Y9qpC3lXe1+PaVUl7BwZBkKQMQ9XjHzFEBsGA
DFzwpTNakQniYkIQHD6msW4FTedk1qQDJuEWKMATz0CrekQypBH7Q1K83vDl1Fo+
uW96hAG146bTO6/VyucGLQ+mo+tASOQgv4QVo2g6IKj0jG5tO82ZM4s0uU2uq3rY
YV/AY8uLDFhWqkMvxxZk5kzYhcmRRaPOUHbZlyEe8ef8WfnnioLJIDm5Kn2P4/6V
bW4tMvJ6wqAC6z5AOyfby/9DtqPRn4y9vk17lPwmmwiWbpW1JIzKfyTXXlUfO/MN
u/m1FFZlz8a5i9/SHl0V91cfkWWSffoEwEeXxiUnJxmZ3ngWAEKqIb+o0UbtL07C
UosI++wcLXc6UBNZk3+1CHmVvAKtfrvHo5bDCUQQLUTOaZuPPCoxWyPQMMkbBKwT
WzBHxvoMdwa9wasvqj6Tb1xhZJLkp9xvP2Do2Dr0GLbf5Nuc1vzkYz2sGqp/BS4t
MR/hI9GDlOrJJ85LtfWNlaEc8V1+2NTqxWSBpnQvS1ZsCNxEICFptiyi+9AarLZT
TkZnnyvWrNqZIx7VkAeKwITTAgnbQSCg7P1mL4s82twuM3mnrWxTsstPlercaDAy
erFhfZasUJqG9IUYRCZDlW907dTC/X4N90RMfApf7+i3yIJm8//dWVsTDVQJ1dQl
JrENArcsIbRGTF8eaCJYoNb/wJZhttoLoH+V2dU4PDfncytsPebLMzmZauHD5qEi
Ob26N2178/G0VcItZLZs23OsyVTdBxt563R+l4zzgn7PJDamGY8gHorWxcLJYpir
EFMvag7dJ1KbKJyZjs5xtY05/VGgFODhGcxfk5B3icomTN4OuenceHTC1F3umDg+
IRRZt3XBUG08aW8nXqiIkmL1iKGy44r6fapNj7bf+R7JkukEFhpb+jH5zQUeFRZz
g1L4uyE3gpdxRMJj/5AF1/8DxSj4lZVjEMpwhwz4aP/WO4d+SbOSjCKbCpEYmQSJ
Qe7QhnIwCDgCEIEDUc1fSXoFIsyiAHUUO/mV1Sia3GG2E/xRC5bdF/cQzmy2ysVe
PMwgfIFA1FAQj7T7iRvRZxEdMLNkGuu0Eb2bDzLuTdsWnXX1t6NbflhMpuaWU+fD
WyHU/CT75jLF2nFw1mNgQeHQiC8cBeEXq+FHV13AfMylna1Ft/6/jObiDujrhFVo
vVgCpYJJtrFwjxfzECd10ewosLc1Gjo65e/yIE4+ITnEGsRnGXy4P49s9gVbt/z7
8RGRI3uYAwj18wux5dmBisqdMlRa+1h4YTTb6029PBk3AIeNfuS+gQtxcOyxP3OD
///pMt5hqg95q1lETRyCedd7HwBA2CvpX9a+lYuLLkxnIifT3P+9LQ8WHpjcdMJC
snaNTr//FMC9U9BgqE4Wh9BhRueXwqArLrGwxa8xbAfzA7Qq33iCnqPOXQ3rpSFB
ju/ArCBkdP/nopDUveLWWY3wjNN050CDYJFTAhluQCJPvx3ehlgAp17o0b+iAVVK
ldBOKQ2H+qKpqNXt834AXHfE7BGG+8Xuo0ZFhq+9mXH0A7CKFu0zEwQ7nB7bsAqH
C1ILJKysvDv+yvfaFuHK0hjtUEWWR4z/58bQnsWCaca9GTXvlhwwxn4VDEiIk8IJ
6i3S6OwIkwXWWNkPvnwixQVvU9et4GHltVKi922Gycq9wP0uYzOVC/uarTpSrUZT
Ln6z3C6Hw4hyqqEYsIfj0ZlWQmK5+KPh4hVY+kZi1Dea+UUphlNp6lZP49WJ8w4O
SM9jN3lYODySLcibrcvaymXj4KU9RF37drS31cyY+m7w2FHdQJgTC3LPSjrPodc1
aZd0k69U91O85vBsE5h0YoV90kKiMbPek5lPi1YoM0qsuY7hlsDUtTXM8/3Q3QR2
9op8FlKxubESJHdedc6vs8v1ErBdc4qZ0zFYDcdhq0MHAanxW5F6nHq0WkVbwCAn
lPzHcjsvzBA6pHzpRpWzbsmWNMXqA579Nt/HqOX2MW0coAFuKSzxPynqnkRR8rAa
kB/VzEauYmW+JCqhQ6brXdHXBEw5MvHdYXlcUBITfucPMgj/4TDmcOhyqWJ8s/2B
ctvbRlhjspaD41dBuVDTG2Ix2ErKyt/4aZCjAfipTDI8UoERiYQNoHeNIjBqKKbY
15Ti0dqfnbmfGtbHtLtKT/SlKn7kShkpU217CFhip4mZqi7OeCkwHJ/5/UQUwHTe
oz/B+GU2GHhtEK0v9ShTY4HuAceobu0gSPMbRT/ybrZGcMZ+kGqJj2q2ud8srcgA
Gvl4np20yw4ao/il411LFQgJ27Br3jrr4oOgFyf6TX+YwsUbsdcj5QPAqLovhm8P
xr7jUuC3oo1SH8Nm7GZT3MOUHpE7xmgL6KYQF9Y9BFR4YpAHFZUyUe0K5Q3ZAfxJ
ztASjmKmdUmMREosKxck690FkPIMUTmM1ooSBCmvtRSE9RkH+aW6QSO670ujCEFC
/aLMQDLPy9b/wqLpwRrVWJ9wlPPRmJX0nbwgWTr1u4N1/9bifGn5MQaGX8ZFfv+N
682kP4iJVn7B+DotmhURoMvrt9B5F+IqTZp65/i1DMDPNvmYbjNzUo0dP0XYzICX
178RbZFiGvmaVZE1dLswHTaq6E79CBl+6lhPaRIU1hE0DpOM1jP684IWiAJ3iFN2
2o1D9wjdEUjXzlB0cZHhEkOtThZsQrw/2PjOSl/xjPaIvJlB8/pNxv5bSdsGeE/8
rxNyXFfoAuLrK43wFIcbWDVmpknVy4JJBOzBp+6l/+sHyLHNhbwru7M6Qc4khT/G
CbDrqmCpoCEWi4Yu9eU0ADMNaZ9D8NCGk2dJ96i9ElsOv6S+B6OQxzIdYuZhJkMJ
Tw1f1TVAZ+/NYh3O07+kXVO+2f3kmzS/18H8zE8yGZfKi8nncazp4WwRidFLOVC8
4IrQ9O/AgNvfcN9nI/1Sak3KzzbLNceE5DjKBivDuHWP2AmE9ggmjITzU0Bfd8jo
jSfipI0I9nVo9NcqYYlXV14I8PiF307+IkVnI4SOCU29B+0znxsiqmxkOkfFN0en
uhECg/BUFD90an13Z2Tt7EP7FhP9QsgiyoCiHh+uq0ELzNB7rSoHgEBqXlyJnqWb
o2ujFP3Ue8feW4JXUi/Mpo5yEgzMyJLqa3ie9k24znLp81evLw/aFkV1kY9tATHF
qin5I7yAWpcj6B9DR6F92EYiwng1VE8hNyiPRQKInpLNVjnParRSBKyddE7JTXj5
/fJoIlwm3/oBW0pv91EcRP4l0/TYk4v/9j5iVb9IItB7uT9w1ujhGCTanMdkfVFW
mcoOdNUI0oz3XJZ2rNyvsYWvz2L0XcVLZy+iwd6D1r1tRJraZ93n3MYvI8Jc/f8u
Y1fw4Z8GqNrUQRbkrQI2dczyZ5sEGZbAP88cYmDqn65InrrKQsKzyoPe6EhTRowL
P9H1wpzhvA01HOvmiTR/u9qzI/darhB7zYGPCXZTpkAJUIM8rVc5eo+fL+GzrJGC
aivbPeOvb2Xn8sFMrsPLYxc52kQPifPk9rnvQPvnH36NfEgiA/0fBY4xr5LjT53R
A3JJMbGsqp3PFup5v9SWUlNUAef8vGD3H1Ui9FvjDs1yZeO9wsi/nS9fesWNJXO3
Fa8y3Kqbv7g3MtYkV4yPeoYu2MKj6uygnyppAtMIFPNOtYrpbouEtYortQSzLY1R
bOkrbqRG8iADvKhrmB5rmZDEn8zqIr39LP3ikXCJNQdT4fiRIPCVoDDgAznjxRGn
5KIa0dUMo3Uv5ugU9Ihq082ojSNgZMBOu5gI58MT2qu81M6pjN1Yo1XpgcR25YZa
Wog+sG62Y47H853H8mdaCrqkfTsLVEi5klAykQk2EhNv8NgU3hP4KR3dBPMLh1jL
fIaUsa2kAiWNMhQizcUKLS+odOnG3yGdJ+qc9+GU1vgCN4puXl25iMQFXOgL2MLA
WXacRCqKNquxL33v+lIYsLBkR7LQunr9SZYOgV5P5s0jtNxXu/NpX9Di9fXp829a
kjnbtQhGgTgbJuapPPEW0jgTA7N4IJP388GkQ2sQ1a3ukAx9IsKw3hbCn+OHHbik
QBm2mkF8RjkbRijbpedJhBlkW5+ViMTG7sA4l8ScKYr46GwjOMjgiWwN6Re5mfb0
DkkT1laQ6I6PtcRh9ipVOYvjh1yK0Ylp+AjlI0MVdSBuvlICcgYevkzWNOeIbodw
vhUGJ5KUuDdXcgqmub78Z8A7pfUXBevDjk433+kCvRjVVscq1fP6FLvebLg9LhxE
XWx4bx3rv6Ty3q1Ru/iiJPApxM2hnmMKSp+U/JpN/f0AEtzjf17CU+3JRHlYWCwm
uGEliIFUI51yT3NNvQQdYWZv3gy3fZosKd9wwpXYDwyGrjN66Pd7Zus83QsPkhYG
8gwN674O3bgd+hy+tJS2zcowLIZsPI0x+/snW9NpG0333j07Jx7tMjiS/IHY99Lb
5Xhz0/YZbfpZdiBhWGbVaz2tOJF5HNDDvKNlATiU21TFC8Jis5Uy01qWQoOOH4Th
BlwTbh2P4x1QIbznCMmdcvv4jkHR+JReYtVyc16KlWJ1A4TbTI15q1BpDJsE1vSt
GHJM0NlIf7g9BDttmjFMLW3NxH584caBdXyI7bAUu+dtWA9MoD3GHWPEMl5DgBIp
GXME49vZCNsCClCdquaQ9aCyhkPdRMgIvHbZQhDUk6DPnrP60TcZaoXdMxuDnN45
6HcwcITk9bcxjZay61uOw3/izpXJrNlxJ0t1RigTv5KghGIuGMPFyA/++sGK47o0
IHvX1tlWVVpW/GwWYLEOkIe05CWBRseAj0SXG+AN7y1kbpH86TcsneODLWWOJCHt
Umft59fa+rarsGYH/Xt8/c95iKo71Ww5H7hI3tMuiciiuHaMuXZPZ9eM1wsfnq3B
1xCZNJarrfIHfVc1ZbEEJ2ocQkwL8shS0HUm7ydMJvFzWIPn5tlb3z50EVQLUhHU
c5gI3khdCE0FxVRYEdTqEAUVSx7kWTFvaE71nKOmQfA5jzWA5lMrVuzTRzD0UMga
YBG2MEdviKWmWISJ6akD2o4hdkHs8mtoWa+D9qaX21sd9pP8wiBA+TUcstaUHfhO
ghwAuba5RtrjwDGdNQ50QVLHnzPaOrZ4ZZcUwvE+918ey+UYk/qxIRazPS7nCIpy
4zmjtL8Kf61wWd7IMP1maBQOW1XsjaQhaJrIgyd3e+pu/Hk1UUGvFYS/03ukXHtH
dM7ptWsAPQx/RD7R4LqswjqOkBdA90rbVyZ/tBtE1MfD0vhoNpLxiq3yHLjvjvrJ
yoWAyW7kb41kzJpOgcVa1GYfkIIyI82gJfNLXBGI3zUWG+rQz36tCzqKIYgEuqI3
PyfWzcyKEnmi6av4WfaAGdAe793ZH4G1i2e23+8qf/SPiMi/GizA7DAvY5ri+/SR
7LCmSZLRZBkfMmxZm0rn7KlIOfFZQ+3hgRN/tTc5KMLp0Anvsp8SBOGUS0D4PWOy
jPMelUO1wYCI82lR3yVx0zDC0ocHOzdoRKRVrz5MbQSBcTdy4/bLszaDjZm+XPlN
PYU36ysJAIvVDE+wBzMb2JrWEpFRqSMcLXZ+OR3XhLYAkYGjOM2kaf0mAGVI51LZ
88+6/AIoiSCjFVspxkSSzH9fbPUWME6TuwN2w7Do1vjtHGQtnAVRmRMB+OMRB7u2
6PJjxSXkHBFVcBSLM5Bbf/5ebl91U9+NoEOngwCP4OFYRSF9GPzHVzfv7xKW4oQN
JQAFZVslb934Y5sU21S/QFtX7AHXWU6gvuIFFL3vaOLUEn2UnClS5HKDL2wYCL3V
HKsm9o8kQrjCC1vhs0Acxh5H3L2BTVSLPqx14vJL2whqQ4yPnZqexXr9efuTC6wI
LYc+w5pGDhmPTHalj5E8/cYinuduszNsAfWQV7nHcMCGJJxsc58D4FU0n6ygTuLv
Ns7uzoSgRKgEcz3UsSXa74rfviNKWGlXXVx8I3/Zhakr50/de+UnZT47yC71Sogv
WLSV6o7/dbO+tQGZ6Rru6lwQtZwAQw03Elsw7f04344dILr4+CJwxZ2El2XKy1jN
s0WNnaRZC4zb+Les/vy4GNWM/xP+9ywGzw+pcwwKhUomOT0/tWnmERhDyOv3Mito
Sw/9AwWhXksSz1tBP5DhuSDDgTNQsfS0SzIkL71OTiatFmA9dGuikXeIXvuDFdoR
M3R0wm2o6aRqcRG/qxEnaaN71NnH+vIxAmJH7+p/VqFhoS9yYoNe2bRpYvkYW2qZ
OvXvZS/EfQffxNLut6yVTce5s5Dpxdn1ImE4x8jWf4M3xWRIXyQ478Kypmn1+Lku
muUFAVaxEzvRWsn/VsCTWYtSIQ8hkAoY3eg7QlVIhesDRzfDhkp1KDCF69ddRC3H
TU3/zKrZY6ZUff7zOlEGnmKzSK9BYdb1rFh4GehFalvTNu051FdZc4hof64myIRO
IgIPwcd0bncKnCstpy81v1VW1nFFklxlDQBKRHj6cBr3QoqLIarC7gDtuATJDaXY
3ZrAe4dEWWxwSNVLqLkj/PZ09Kq+8kFy8Te0FJrPPlVD1E1Gtq8GcL1rDvXxggtc
o04umsLH3ogSw7Jf8me0Nli2AeoeOhm7WftJdxRNb+yTs9FWoXcjKMLYSPDxDEGN
XgEHV+nzJS13TxYYWs2pe5Tw6PGe8tUsyNnWXif5HfcSLopHlILeR2AolXT/Oube
oLkAJupOg2vII3fXA702r35uHniQzWTrA3ZpKTuu2Nb9SdjWYnEjM0C3/cFZmxvD
AY7Q5ywdgo8Hjs/VjSQ0Oiw/JEDh97VXQ6EJjUEGcsYTxOwuXb/B7XHI6Xvepl5G
k5aG9+O0VAIDKMQ/oRCdAliL5xoL+gR0iFBGm+CmmTgJG7Gex+5Jv/n8BPJISPDi
94EdTrOs6+SJrRbTK0eLSiy7OtSnYMfm2NwnXeDIajEq1QuPkp2gqqLY0iFx52Ln
e3K7DlK0cl1bem/mLZcT7adkepFwWGJaeGKIVPB8lu4+kjf3Eg2WdlabTONXZzJL
YGvd1ftlZD5VgJB/uwBdCToSuiCPp7s3rd1EEK83NvIbSbJTRVY7aDTSAh9GYMaJ
dsUA11g/4LgBejCTTY5m3IaezYN87yjkcxWTNMt6lSDIxbvFLQ6wJnUWMqKT/UZn
XvkJ39/Wuog8NxGItUY/BpGo5BYJrwTL7p1SH04g1HWesfjagAVaNbVp9/5ioKDL
m6zCxhMRSvbAuLVsphY3oBOXMkR3VaaGWVuQxaIcd/CTEn490bA4QYBEADzG8Jb9
87X7u0/mbfa580uZ/8UZhTYjePr7wg3rz+pOuUkVseJjHu94ScFwqGDV311t/opE
A8n263xKCqSA7qEccFtQ3FhbhDgFow2BPWfbc7yXoWERZoK0p+DPtSro+1D5j7Zp
eptaxCh5haKh1WDasSdJPuU0zoIefMXLmmSz+2mBANvfPRrt3OuQ5f9QVMLT1EVe
qw1DuTLv5rMQZjKHeTMEzW4d+14w7Erl7+XyrlFPH2/fJ0+1kydRcAz/3cerz/pr
ny2QKhj06Nzu7qof+DhpsPhZlP3D75r5AfUZJYwtGQPRyXh7ZEUdakmaKOV3bfVF
jqpRP9zdxgItDIs2eDFWd0EcVh9C/dzmUZ/NZAsizmg0epSwQAmEwZF8ni4/uVH1
Atk3EoQ+n9YWUYQKWRzvn+B8TypIVWl8uKmT42kx33ISFCXD4oOLxgR/9E4x9Psu
cmBV4u1h3m05UGczuL3uXE60CFf8EYHlq26P4CvHCeNZ6aDWW8w5Dg2UITZMDrg0
l8bb0z3OKFqatDxxZABIzaYlJiPO3QS69snXj8+9GIK14//qLxm4+aN5+GxC0Pe1
IMigHfEMozskTJpD24++U/un57lvfVfYT5L+XfirntP/ESX3241v5iwWPj2N/B13
wPxCDC9y+oy16AjoIFTdqzW/05weo3oN2mh3FRQ2nV/7RRX0diY567sW0JwumKna
JV1nmHve24ExbtFED8+mRi9tPP6aD5oSLUdkAYjTJaG+UhnNZIONyBqcaOt5ypnq
rEnl119bgJdNWHtQ9yJEtVob2+Olb8CVFFHfwKEa3PEvVmpT7UXlMKQQfPVZ+waj
BcO9YbwvIKacoLGou94acBCd4B4ipVuxwEaR6gdlDmxwO8V9+F34wAJOpHWKShw+
CwZD1SJ2mzQtaMZyAXfdaikaCYVtc8fY/GPnzNLf8ObP5B4wHqYeeldlrQeLI4jF
+astAk2RMuu0+LMYjtT8BaLYDSREk9beF64Vp2IJk3tfNyZeKfOimdbcAHWNbrTi
HOjSfVdEFbItruXG1BO0+BN1Ev2hi8XL4luyLl2zYwygRAa3mi3sTtk1DXzMpVAY
emiYXzng81s3cpc+NmFen5BscQzTqXWT4UoIGqNdt3rA18kkdph6YVCoNe0gPG06
XYnIQumrmn/J5rxH1SWeMbONGX1wrWsTduQdPcrWqi/HkqLB4BGP5csW5TiLSLhH
Rc7PiZ9s6K9a3knBn8hMn1hyKOJArj5sczrUMsLeIstd7UrzUuNFM+zZMtdUkeTf
l6b+q4JPnvWKYIp3U2l2DN0/Pgek5+sY1/OXi9OmqyMaCpGcvu0Muf853v/sd1PZ
dAfcm3MdgF89ViDSE4X3YLrOG2NGinGZruMEX3GuyQqXxjxBmHw/h7TGzLW+06FC
oosEKtdwgQONhF3greAezfBiV/Urea3p0qbl6i09B8lqKbdw4nBixeFsWhl+CJ5F
dZT4CvkMTakMgWwb7AvELelmJpH/PpzOPEBFzEY3Jfy1En0kj3Pc7ghYXuQeQ5eL
GNOjns6SzLcQDnkid3sGCElgb8HgWJfZvXhNRJ7iTPutfdSAmx6pi6LBrcH9gjCF
rXmqelqEpDDuRWk/6CbTZXMamPzJyJtmF4Pti6PequDZ1AWQZHnwBcqWbuvnZWNd
xIqYNFMO7u8dSHYzkHl0CISd56u13tbE3nnFV7jCkt73kzq7HdJfnFrb65vpWZHY
E12Lk3mWUo0j0LoFMeXD1hPNqGLUbVnSfJ4r56bh2bAXl1PbBCgUKv1i9I1LZdp7
7F+liQWeBrygqyqXRGIPiFBfHaROC1pGnL/CtMRkybZ5kKp9qOFLygtM4DoQTvNx
kKcF7dZwg6gdQjJgt4SP64gAkr/9RDfVpDhupeNmxeLjz12yTH4e+vCsG2YIl90y
1738zSR0a8/8fx4YaNlQ58F7P88q1tWbLqXZ6jxsmraqKfGuq1g0lYIX1IY/MOgf
sQMOSUFBHFOZcztLKE7SvUTOdTikyU7i31T2eezt7o6Q+gsHPAZIm8JA5ckXy1BW
V6jL0ZXJ08dzM7ySFh5XJ8cjzHATXWF+r9jn68PfquxtDgFwYtqOm6oWl+UptzLf
4wKnGihOTB8B2a9uDL6Lr3T9nxIkGLTnbbSs6IcdXSuANNSIRZu7sfcgbvR7oY+X
0F+c0BPAHgesv7CkGEE77vOUM/nWsSpJ1PbNwRUuso3f3unSFCyQESdWWHjQ71zm
UuCWoLZeDLU3vhdlfMCAg+CQBEIc27JwhiFrsgyfeWzq31GooB2FGdgbgXFGfZof
Kp7dGhK1ims5x2rTI6XB5LIY//ZKtY8MXzWk6MJmISG/vpAqjeNIxh5CZQsg+iQp
UuCEEe1z/yUcG6i/2n3kbBwIZ3bOwqk6mvi4Pwj/NdHJV7foJtMTh5C77B5mUOnp
tEl/dJG9GU/aAAREH2N7j6i55FUN7OYLR7e645NTOAdteURwM1ntZ0k0SSsrVPNt
ogfBfeOTYs2ydeImG8BF7bbrFdcJF2q5WzbtNYs16Ly5U4ivLLiAbJW8sYpDa0J2
KlOnqfTeBPmosz9pyi7HSJ7/MwgtNvXrOvuhDhxO3OmU8FSjYgLs5npghqNySPKP
oc0Mw2MkB5fLdtavgyKnGtQ4PRhj9upIyG9edIKlvLtwdNvzRgtjqTro58VmIxST
SV+K5FH9yiNP6NLrSbJBcFcuHjJSspd8a+G5yMZKN9qG+9+2uRGpiGtslpymo+nn
W/nqW0o05JUKk90yUiRhvheM+KpZ3c4++MGcS8L635JLN/igbefw1F4tG44WwaOJ
jlGiBR+vJ/suyGRxVLgU/IVcyQS/bI69eFXHtv+XPzeuIc6mOHKecjjTqagjf5BJ
zFzkNZ8Mknqn4JmWjHZpykVd8x2zBa/IE4Q7CwcKd40Pvh/x/Xlm06nvuOUlob44
aOsmSoBwNPQmeHLbWYHFwYkGU4+2aZVckw1/jyVWQ3tKgAB7oVk8lIDQddONItx2
rXghG17KwZxrTnmBNLIyuxBAzqi2W2VzYTg8IhbRqE9D+w79WxpR8MWQLZJfcx79
3/sfWlMeX0imoszRUcqK6Ax/D6NpQPfHvO+2ZHpfqhvmML9VtZyDA+JQqgra1ThE
P9An8Ak11m1ARyqx/RGLSBfa82QQnHL3qOOX1ioM77nQCpDEPrgYxv2pLgOYFJkS
UcBszNCocm1N/4obfzmSmXWcsPjVUMlegykx3drjIN957ERGqqBVAUxgXg5+C0uy
J5oEZWummNzeaLqmLNWNlXsdNROhVLzvSlK/6PlBuksPziaiK4e1T1s4dwsSKZrR
FftTS/PP0rq0TWj+PqjFcFvA2hNZ+qPPtEcVVNI7/iZwz42BktvL7GwNyP5Nv4Ow
Ab6SNpkrC8jmCrTRYJd85S5/3hRqnxrh9mJOIN0OYjcO3seWyNZQurIjzT/+yy8Z
16zn9q44qZ57mKBJay6Eo0994GAgvyO5yBE+mSRFSJ+VwVGAqOjqyFisF0FtsOqL
mvp9RFaQqKqQkc4ieq9CdEDbKPgx7X19euwdfa71xoDbwApVmMU0839G+993VCYT
2TSD9rtJZVRlO9pAcaqMS9SiqQIsk1bkJX03KMamf8rbSj2RQ68nq7Q8bXYK7BG6
ICardx5CYOs4fkaXqVlUTWlfBgbJC89JeVFv4gjHE6HLYHT7TBEKoMYj3iABpndm
Sh8OP/KoJ5btDZ04Iec5Mq5gonnVtCU8Sqh+PCFhmuKh++pFepUp+PCoPNg2f1ox
QwyrVh3Xv7wVwoxLILZ0Bf9f4sXII1zE571TXL3lHDwmternEQAK4LinU4Htl70Q
5sQWffvJk56lpP08R0Q5eBgICzuEjU8R/YSHlWO6hLWcYKHh7lcSlxncK+KNTPy3
JlHHFKet2xbl5mma4j8NCBKIU6idogcWfN4rDqKLAiMRFtdQw168uf5c3PmFXHvn
Y+ED485hbxlmxobbQO2J2t2fbYzMhvrs4T6hF7XXSNTa51pPr6zYUikCLJtNsXqq
7J3AtK4vThh71PivQ4DeDvOoRdesG+WnVZCP9LG30O1wYKp4iH7nab/IceJqupeY
CPw/TtThsD+yxDbyt9vpClZsl3iK3gKBNq0MrPYwdghc5ITsdeUvueP5eYq04W0l
yqum8qLha8fHuRoXS0y2i5jri2MpLgmGsru1ZQLxXWC6miUnOzWlh8Ej5Ylgo8zZ
phk4ncg0C/lrAM9nM7yjSPO6SuCG+aQX5nKIPJCszktWWFllJ17ez4cqfje05qxf
uk3DsMz7ctBPI0JxY0RzIBXmDkUyEldV3GWbvKX9bU/HIjeUTnAGiCE9jhQD7E+2
FCiQUtjr8bC3Qo3EBMN+7wDaA+9hl6O/tLhR2yy+y8wPVmo7mTsjkDnAAb3vwZnb
DJbL1eNMGGtx7MiC2oZw5c5vcnhgsF4OoH/5PWmrcNzs9/tdSKlEk1TpTSkwO+Nc
laP4U0lBx/3xRi6WWtYADPIuHBjkshrwFjR78GWmK1ObfSLJG4PA3vhj3UMR6KS3
viDbLdfXncSZL+cwEa7H24nsGx7zLgp4HJN4rcaVwJ2xc3Dp2fRDpgsklEpKxOMh
g1uUeH9iUA5XJj1SqCTKMMD7vpWnt857VciTcXx2VFvxzvdWSsYCjN4AezxQrgxU
52SQyRI5akcWSWgUNJN93ugIJvyvXDF2AVzuPZr9nnD3dYgO+1GfEkjm8fZKw0F8
cVC5pCCiU1L6Fqyf1yC2jMt9R/zvcT3vvERD57pTJzNTLbLnH6vRnvLlx1iD+eIZ
SgBS43TgrngOznkaGJMx8vQQhK5i4s8e01YTbelVOGHV16/B4cXO2Xfv8lOLoVrv
+x9R++UfSQR2jj+jG3gOrJu1kgf9WsrHAYxQwfGJDWHPPC3y1WNzuQxkqVEGJyVt
3LpgKGJDlzUPU/VkVmL1WybyDKiSGoF5ZYm4DjQejz/pD1oQbBJmeXtpqLNUAtea
tOu2V2wb1CAZmJ5G5LlTikv0GTgQunOKZvuF05i8LeEMnTN9p5Z6eiRxFUuB3LRj
ZgWYv5CCwvXSww83PdAdDZOkGZ1eTLaOUVysgnRB4MFncgshHaS6NK5jNsBqMAtK
w+AnZk56CeXmAGGjTXDLfzV4Ls/1vsnPkVsY7M9clSFp4FBJruP5QqpDyEUQ7Hfk
UO2gZyt6HAptTq/rMngg2//avwSCSeIwcjaDy9HATkyvDsMT349iaG2MgAoUP3JK
LO1SkVlB41XqmooB9yi6ZQhqxWhUYWFs7x0edaDIAOtUrS0JLZ7z27cVDS8fXUuQ
2waxEYp/ffWmIq1V6WlvT8Uh8r/tA/4Gz6hxx6mhJBzpy2+H+LPiLzTDS8wXKw/j
SgJbmvuwWcMGH9DB3wUxOyg1y/WxJiJu7KD+gjTERhPBplTTn2/zC3ElG0w/GhQS
sYIi0ozprbYR2A2Yv834g6xiTNQ7ThVankryxWoxk5mSwG7taaM9chj0sW1wlVvq
eyqUIhJ/X7ONSbriRK526H04vz7shYq9HJkbjn4IeIQfOx6Zvz/boZ7/2X/JvQ66
TDBriZX8uPKQtrAOIdS+hCNSi+G9nyDbuJsqFMLnaSxZ3nq3Sqdnb0F75pUO2jVJ
4DkJCPIkU7cItaXuk30UpE4+s5QDs3DhG34GTedqJpx6YOB6zYpDB7v2MEea2sXA
KvvfD7qcbEzTcQZsQ/ZZGtoLpK0GaPctr1Je2YrVQOBPp8do7yPDSSNgBFiGypF0
9csPacYi+SigpVJEzTw+c+kcbfjpyqwsmCvyR6Ln/+gc6txQhiwdZm9SPwWh7imR
mVkvnYJVRYdxHQqErVHuf5DVcqICOAvi9JTbKJ8udEVvJy+qld129Cn/kgAecN5f
TcDYjbaSmq8lgsSq0d+tp/InYGza9I371YkvaBU57nkQZgLYKUwIJie0sX/V1wAy
nCBwUsKoHENTUYJeUsjKEPt6qJo8SP8oOZ4avXw1xdYaTOBCOpykxND7gQkJVB57
2yw2l6uyFr/h+04fKAWRRdaBlCEeMEdcYus7SEwGnACKOwzy05wReq/q4g2NxkVI
CM/3tq2dkUOVbZazB2hqIiDoovG/NX6+LnV87iAYoiK3FI/hiN+SGtYCzpvOH6M+
F850HRmdt0V/Z3vA1gNNofzMA7kh7cluovjRr/HPzDlwJZ0+H9fb2Q/N+BJV9jEM
A+f76qm1Wj0qJVLjjbtX0DMgpadSJ9RUDysWSB1mywoTGyQmUBsPJM90fmO3RQqF
+K3lUdtLAXztNp8KdNrzW3JuWKRIVKx0qeRS/+rc8tAa3sTIN+NtsKQDsLbzQw8F
DzdlSmpMZ1UP4xGffGMYZOyLagRTkb+l7cSq26aQEzOFFvNNjsDN6GH+kqOsBcYI
j4pnqz46joG+gptqXues+rB6MG02jEskZO2B4ecaUHOupMadanhW5LgAPSTCVmX3
sc3RqM1uI2n5uuCJP2pYH6vD/Vowj7QWvZxVwuXBMSfFZoiTKa7lrp1O7ntooWYb
/PDLOrydpX4/68BJp6Xv9ghpmqEBP1uTWZZccgIP3JsVhKCDzpbUxf2wKtQXRMLG
KsXPOU3NATm85/milB/7CFpxUFF2uRHdq7RDTUI6730Q7woQQqY6m7STORPRX3kC
uRo/uWPr8+RfMlP2xJGOnLVob8NJvj3NvvYOxl4eU8yH1rIzglzCgayBY26g7dW1
6E8Wlmzda06eQwyrhGK9nhUAeVaGTno1jEw4CXNiTI5zoaGj4I4GKJUvu18F1nCT
b9yOutRouqaTyPvibu79J1lPTKIerl6adoS7zWtM8xgvwwuME7j/ATiylQEsmD9Q
1jP1Q5jYP0McLqSbG2JhhZ5va0uGpApX/1doef4l1NgL/PjnebNB6Lzj09S4cBGC
klkhbDduiFDoe534jw9kFyR6n8t43uRK4rze1qG2jBs3SVj4bbhyK33ykLEsq868
QrpQ2JVoMf58uBglHG2NFkEA/LJ8+wXAbiFHronm3MltilNTfg4VBND6JYEvovWA
PIeM8Y1RJY04SiJaOVoAgZp8PX1N60emhZsB65LcA1LHJKb5Cog/QOLGLZoYUZbB
xJRKe11xFwzlK+AG1jezQrz/PuOZICAbKFOKpvr76LmU+BX+LS3aFTyqdRBIQmR1
FhuyWfDMb4Jh+iYBIZ5//uLHHrylXZPAnPc/r8DGNZLB2nzC8evSvflNI5pYauZH
KxNWfuZem3S+ptgUQc4DIiN0EiXU1IXf1qnlFxgun+1/EIAY9Mw1PWUDBcpBUjQQ
9bHqFH5dffLnVRsghgDxx9VcnwkKxl7R/JRLHalPe3oEq43nyFJ3O9MT/sdKDUFH
f1lktCCSkgSP4BZmHhO3hfhJ6bri8TKaTuKF5UCp9iHXwqunHiCjX5/PQNNzT1XV
VnNvR1QFjvyYfz2Cuv0Ib8Ai5CJz9QtioqJtJTLmwtuFJANhtRnmUz8g5PYRgYzH
dlUtnwWYGA3NB9Pqk7aFZhp+hmCZ2E7kO5vWBRaDFbyhmv8NBoHK7FPkgqwzV+T6
NtwQkcn9d5Z0tWTuVE8lo/oYsEcsutQMDYOhG+M5Rri9vHQGKbpXcnxxGCOQAYdg
rtP2TCjYx9te3HlOjEZRf8RK9SdnkbOHRDKe0W8w/oIoUCWanGaeWuD8CtF/xAKw
5FsvJSSxkRyvuy09mcQ8q3PKHBL+4C30dqmyAT7xfNVCMrLrkZ90ydKEwC2h6E9J
pbTSaCYIR9hmBzZHOVTOU92ZEQu4RwPwcS7Tp/8P20XN97z/+fFeCnDp7X3iRraN
rXJQ6k1qDIP9SMTjlKW9EwnLhROSzavX+8iKf/gkkPNjlirUixX936Xygvy0bsp7
lXDEn/QSjCbsnN4RqZ9XRaqRK4sQwdCIvkTmaJM7EtRtBcKTPdCeTxL2iY2xMmYZ
F91xCvE9/WUtdCU+CTh2D1qMiTk25hrhSw4wuDS1k5FLK7k395e7KckmByse9DJo
wiwKc1uHhLt/uZd0LLFgxnK0ugFgwlhkIx66tw12bJMDAiUYnk3DLWAOSc+ZS++D
6povkrotzBMqt6pK7eTQELd5+ULcqAB7fkLU0UpE4yvVeIXTBfhL2tAjTcaGuBo8
Ovzur72IrG5kukcPjUd3L3JOIcUJ9p4AnZf4qc/e7xQD7KDvGzJdJ5Oi/B/q1WzR
rrtvpfS5zIwqnKu9+Dsd/UHjikoNOhsnDjFmGMk/aEWpiGqrpTCeZzJ2qQiZP5zO
VMpeNH03P3A0H461UiKCGn85a1yA5bzz8debu/9F5CSnWXtnATpbcBRoR+FABAys
puRJjFCZjuRo6eao4vCty3lyDQpBP9RpBrd5UDUtyj9I/r/ghhg1+uLLhvX5rzt7
h9RLh+6m3FK36nYgNPDbCIPbg+RZyKyYNmem5a0yg9WyvITGMZ3rr4yUfE7FqlX6
IxeGlmWXQ6UmPlTUOR3UKgwi9UXYN0Gq0QLmjYXlcNIPBcCUfT6PkvHnDvtEs4zM
ri5v+LYiPuzmgVXeo3iSk03UPWI8KqlJuja0b8tQl9uVhv8ME35/1cvHkOgNUzXm
ra+DqW1OVISf/NFgnuakhQA77+3estYvDtymb60SWx+8h9kue/cN0ApUs51w//Q3
70RvdhBO2y43YLr5sG2RpEISIbZ9PAEF+JhJSQYNrIUmC6J0J2rsxRgafiV9YTRx
e2QFZQHux1OvZ+FqS2BTjZYxGc7njfQ++Oo7SX//C4o+Qv4oZwqzjv8SKJoazHTz
RnTccWHlV8/gEaNbuUePxaH8JetdPkvRBGfXTIlwRZNaQNBjyai9T56Q+vPLcUPC
GsZMHIX/Svn4cm/wOxbbeyZTV1HtFXFoPQrYivOeyQipRw5K/54UN2IOMcRh8n3V
95A4oPdjwXdFEGUqwjF75VZyAkPrd2QZvZiykoKI7e+8FtkbGrPvq2Ho7qQgaJTS
iQRcCxc7ztU/7BHrUX44VQVKk3bEgc7AsfHp9OrO7L+5TKDklmFhnRdL1P9P8+05
kpPC7foBfOMjWSC9dIz4B8jsUB70haYMJBKJop4P3FcX14le5BaDfrFcrq41CAV7
UaeCqF3OOCMJp91WiD4SEAo281dCc+8b/ITuDSkhYOE0jJhVSNIV4xA7TR3bdCEm
gtg6n2+rrUgJVwJTNVV12PLrcq9ZIZlfgxf9Fy7fg4BUwh1RZS72D7BIJv7eKHRP
hSQQl2eXLKJUjgY+KDbA/r7pE3HorWL5dR6dMS3yULs7/qGksNdG0HeOY+NJpgGc
TozbT1QSEAjCcGVpwMY9udgb/BeTvVvYnNnUlnWYgxjnQY/D8KgSrGpiMVoZzCb5
Vwhsr/Er+zrkrPB2KC8A320gIKJjWs6678hq/b7yJkV3UlCUmpQAPobb3ebEAFZK
OSSdQJ+yuingNkVBBIRnEazQ9T4g/8Z4oUtmNUqrsnvpcc/gbV/HeDcR/xxzw/o/
27Q22JLpvnAJMArN4fZ9KRRU7+UsZNCca4MQluuaq/H6RyvX8KqhAs2OdiaUZhJL
priqBRjy0oG1a2JwN2bhe1XgB1fi9CZt9t+zTDLsAzEM8JA6qimClXv3eBTUGBq9
EO7xNmqFUHbJ5DlM/WhnphILXaguY9m1QThORcRuWPPeHEmZc192PHe19PaeQ1Nw
85VI6Sj3mZdSfcLsWZlyUm3uVw0SfhGtHFWU2Se6kpW0Ber9/XPmis0yzuO0o08Y
USlJGJm+42RDMmU577aLRLWXRDK2r5rhUgBBFL8rzmRKmXQFyeKddwFkiZgm41/3
todOUjdR+CagEJ5LfuJDPUfGoWaG75MDr+TOY11tkdb/5j7DH2BcHV6cD694Jqw+
7aE9vXZWNknba0K1KuUj+5xcdMiGzyj+oe9/gkt+5WJ6V7rk8xWiGAaV/sAFfYcd
0DybGW/Qdw6QhaBOoq/5EqDG5TtA9W60kKz6SJ9jKu8sAE2mnuolJcpvim7GHEB4
22VWZ63UwUgRmSlX7KBsWjbyL/M92gdcK4F01/CQSEiR1n1xZeb/xzqD+tmEYeRp
Elkx/lGyQ1jVEr0InIFFXSOZCpENHu9P8PSnueU0nYRpzAurYkyrCNcIV5dhr2yG
4CTLLYpmk5/xbJIwD9fuh/bYVdg4f0+yM55Ejzyyada8sngpMVrHgJEXg8qAJ/1u
VKhbXkNE6XEXBvqbJh8Ob2FGofeHfnQhFedNHRHmQaZoRzsE+H9PxjyXpjUgHlmT
1z737E/WpkjYbaYEzkloAvdvxY0m7c3hsZG22MT1ROam9Q20PMDN9NCMwAwNv2jI
KkAyW03GGB6iTwPUfIZNp0JWficteUi1qboCzsLudvNKAEORflO9F7zalyB1iaQc
9v2CPjcQC2vLZEZFNZecF02CdYDvsPGoIEMz5w/qjumOSy8XD/svv0eoU0/R1LGn
tvkz7vg2IW8EcLIX7E3icYYgJiO5aBx4xa3i7lzloFlHN+dy9Q2lQ2FB751KMU1S
4grh0iHAwmF93e9Rjy0QYQcUGaTvMLBTJbdRIykbcBBnsbhV0KEwPwyCOMaxi+jq
NexkMkzE3rSJReSDA0BQgVpgatg5JW9OBfJjGNXqBgNs2Op4gjpSeaS/BhIW843A
L5FwKEhdNlN8t7xN7r176i2Ch+gb5ExQM+0RfZas+w+ZAbzEfLM3U4u5h+LvIvcD
XIiAYmVNrRl7nYrBGTUd1MI6PP4Z9jtPHmJBToaU9m2rYz8Qk9dr5ahkt7Rd8QUi
2nWUpymH+WwbjLGBB9nZ6/U+VoDQxRbUWKWyD4ZoX1kIFamE3XY7E8rszFLUm8Rk
g1YU2QN94rprx0g5A1MD8iONy+WJS5HZ3xVzEoEq5ZftqioOHCdV/Kh6SGOUni0d
Yrn2L580gZ2Xqb1VTGycaThYBQzmaKqFwVzlyIAvZXmn565zRTH0IDVKozYIxEil
S2wz3h0YURCE1HQxAUQYAWD9w7u1cFwFgFQcXnSo9hF3uoTA+sKmdLx+l8bnNsyb
ZocFveBU+FKXNo3BOwUukCnyFgRdGscYWPv0lBOptlFJa5L+w50EuSrRJUDCIC+h
kroHoD+qNyFJxbi9pIAMhqry/ILw6miRO6+rAlM3ZyS5IKH4DOLpYbYB1BODDML8
Xi7/psVU+8FX38p5EO78k1aghzbShXLwOziwH2CvlokY88+PBQnYpYQdCVIZepav
hCFbuYcdm3hA48+Y6/WwgtIpqDe1mZs7SsnHDct+Vwp9E3HPlFY92ATH0P60nK2m
/WvEOFYHMzroMZzDKi1myyQUSdXJMqiiO69XBB5a9T7arf06ZepUMntmZcLtIdcr
rLCx9os4WuqP/8Q4/1Aknqbnoh9+V4+M5MUAb6QzbZBii8/zC6CRJBBkMEPO5/kU
Uh23gFFuPUEWW+brPMgICozm1RVKRwylnJbr07DeZauYBG+2snXc69x8MortJ+0S
jxMQ3r7XJ25UyNp2rraFV0jT9BoTZAUzUyX2BvAF2YV2pYtEfUOov7HGevLIt8CI
C5RugyMnG6VBsE8aVYoUQH2bZ029uDfpVgnVUrdOrpi02TLVcmEjzTuoLvTERT3Z
epjtJf9J7v+9a0kg0dqXIU9K82tdc0dNA2gMxW3xFrZzyjpFgaU4hbl2Y4BRAGjg
ksieqGLHSnuzuNZ10I4C9HtlnFrR4iNT3xEeMP6wttgI53WmFLLSR6VabF+JZCpl
SN4JBvN9+HQC/NQG+Tmt1Xup82QqaMAYMzpgvh0cjMrg1Xp2inoXrn6no/4UAwpW
Xdk3vQehv+1BoO3FTeZr09HWfn9GFt+bZnDHQmDdEXp3ax5dnfhbzzSUoZ4btE8+
o94twXkPu2ThVetyr06OsuiOquN7HptHSAJedexa40135dy/XtQ8Uvkap1+wGBjc
WoPcnhxPNQbCk9XyBGGQ1T1X68prF0xiKtRDGD1aro8CZuY3HN0k65h2DiW7I5OE
oydItRem6rf+YZI5+794AnjEGpK7iKWmuL2ZJ8jliFxnOFGrq89eJj2KRciQhGoo
kc9FZrYkysrYyCQheh4rIhy7xPng3SRMHYCt81n0+UpYbgKNNFECcoeBfvjPSR9J
cCEnQp46RoNWIw1Ai5d38V6SimBSEsKIKZZUdvjovydkLQQ/by26L54XDOrpKjXZ
57UCAERBRicxyENJRR/EVu1pYnW2Nw0gECNHCY+9jOiHjxJYhzlOhPhajXIuRUX6
f3xR3V9x8apwgWqfudx1y6GXgLTQtEzHbHmo7ynRBJ2/Dq+JpXZznvv+oG+49x+Z
BteyOm7lIl23zsxpG0bX0PAUDHpfIB5IcMWBz3WXTkF6ll1uTS8VruNAI6KCKgNH
XGKpIG7IzfZuRyxgQn7WqOZoOYX6ywPkGU/MqzCVYoSc/rKDherYnVf3DMgh/XnO
Fy4zbskRVuRhBnI98KnfgyCWozjH9q/tJntfQr4vSX4k8YMFEHSx+HeawSPIdJoR
WQuhKHtGwpsq5TEoLVOZ7cwGXarVrLiH2K0iFOAqVlXPFSGfAsDITT5Gv3Cy8Mpf
eVWEvLoOYlif4PU0epU1yu6VAX+tMs5UOCgYWa4dPqSs+6PJdA7+/FYSMHM8HP88
lheeXQofCIJ4Spo0wsuZSplLMtcjG/yV0JKqt4whvpHVxtDYxdsfAKoB+OLYwiMD
OOarLlrd8at4iIgNiKcudueRY3Wr3rz2H/TjTsASEFHlNrGUMRg8IFtc0jr0h7qf
llOpOJtqCb2vKbeoSG7EF9xW4SlP1SR7Yf0a8ZAU1FSO6+62RE5Zhc0R8+yCBZhU
mVcfWXdc/PS5I3B+HJhDiobK1NZiILKiLQ/7GGW0ieijgZRwf54quiO4JkVEZUgR
oE/QT8+1j1ucTtXFW40e5GbXwSOIN1QAI86c4Q3DEkZSZ0oSazbnwfGGYvU+FGOv
H46PXILfjypCEiPA/Y30ITVyVSu1+XFcQQuc7cYwBdNMVScNC4cDonhPFghHdTIM
YtO/FgGsersEr4fcNXV0lvh4vtSWiIZ9HeaSD6KG3RAhXVtJjG9ieIBIB0cm73L6
1aCDC0zXXWO1EMSBbyQaruucUD6ZslzRDH/adJDs477OPo1Ftv+oYtbeQUstrOIR
dwftmyUIW+gH7BTKAJyAnTUhMyZ002v9TNT1dt59iFbgLbjGt2ZGxldGEMZvN6tJ
nc0og7c30JQpJKPAQ8h6rZHH5kX6pMkhmCswjwc0oMN5unuOFA/fqeQt+GmeEfwK
GeXVGxBgk6vqxhHUoEt5bHEEG4P2drAgaGYUpCPymfZzyLukblQY7MZVQ84gm4gV
crPHPu+W+IcopNSPSTr5T0qZjVcQ0kXx/Hd4rKQTh2yibTb6KUeFO89WaUxm485Z
VDISkvAlAFTvJkXdInhGyBJF8hHwmdp9nAH+nXpvg4Om8xPru1O2ZH4shvTWyjj+
dyEeYnUEfQgfOPutXDLNpcWO8QCUF4O3/vFi+wUNnjnEoLMztlVvbUUcCSu0DGi2
YaKqQWlLfaE8ElDdOgHpU7pb39D3B3ZI5/L7+ODx1YtUrB+yzVY0JPWq9Eu/p8Rr
48n1Tw+YncOaWdnhRTift8r0hzjeVWdQLp1U1iVJ5BR5F/VsK2mlZp7JrU4VvNEn
No8f6syZOpgvRbmIuX/FVH3o3663BQIRwEhL3CVjG4MHWRMOqrWrRFjoL56zB01a
t8G6edxuRcmgPojGi6yLZwi60gW2UPQfQdyM+jBBktJeevovwHTRdjI7+xHmhxmI
Vb353vv4hVdgMTFpgVyBrJhCPkNPWsAzNNzsOFC9NFEzee20FBbrC5W0wtbRTgUb
sn/yDP6D1rqSNo4XURSqE8sfJmvdfAeIrLRVg3hT+TRGyXZ3kJOfLDLDS1010gD9
LnoeKwem+EHamALynU3iC1sYmcfboPWZYeXacRD+V24WimRdLNTwEUWodE9YywFC
lhJHbAlCt6NXawq0+GP1MnZKEsZ1sKCwzdtFcvRhI49cJyy8QinK2Jjosf0+wECr
8sw2e5GQIbzE9siZUo5B+Vhu0P5Bv3J+WSu3n9bUI7f/FrdHR9lYAfvh0YzItRJl
Vy7IXkURKWx6IKN5czazo40DSd8EpfL0CwtJUzoZK26zNusAFKyesdkvVy3N+Sxv
jXDaH2nBDS1YQMKoRuf7AHdU7EkiioyZ8SxkzSyRKRdxy3H5Sp824RAYLlYJlj0r
A/vHcIWGkP+sMBQxH0OWW2mtU/PYQgJHcdNE+DSpY1zLuvJx2OvUXtWABNz+hTP0
agPwtyLMwdq8E6tEE+9K94eLx7OFNIi5dYMbfxJ38MDctFfKapUrpdjNxuBPPIUa
/W5miGw73u9gzlya9hJtxmfh82gqBzP5zCjUyKGZsQ5re1Uu7Iv/NhYxLhA//Dr3
oo2UiXNOdSv67juBcL5eXEWIosjSxTD7+vnShjhpPj/bNubrqA4s26CQgBKe8aOn
MAgGP36sSFvf9rRLfBp4laAJOoXDI8xtkYr8UbXXjkmnwV3fRlfOEAk3mklgj8iB
Y1sJRQ2hCZJTflapMzWKVMlJ01ox1T7Jy+WYcisAvi7eWcvaasc/F/SXTgZXBafE
HCprMuNEe/vSBP21Nq/IgdlWR6iOh1bLvxaswp5dBVW41BOirXBEQun+KQ6aCxXj
GkBXVKwYJBgGn6Gx5JklyqTFn/P1KgtxgHzU+LtwXLSPQ3zu6/53L5ARIvIlrDOS
7X9UvGthL0XCSi71A+Vv8mOb9nmhGXgUR1NinDa3rUxUnF0zh+n4wHnt6HH4pwwV
Wq6fN68Fzez97z9azunG93TP64Aq0J68iERt8InYKLArXLQjgW0xTvtOz48A90z7
yMWE2wMWK/O4r6V084SY3yeBWY9+2HAmzMDkOaBifIqR9DH/8C+a1SsYnqrN9DiT
C0Ti/NPOCCOFdw5R6FIbAxjGdAllZGTDmN0Fv/UMsT/YO14x1Zg21joYKM+LEjtH
2UaKD6KG3Iuhyc9wpnG8lNi5DZOXepoybGNuJOYt5LnuPrVWL04rCB9twCOR3dYa
YN5/DTnmQA1ZXbSRZUCR758ZyrOApIReUpLwAqmvf6pBKpVehSis3iWFZEtk0id8
+HCF56n/AkmQIwEjaAfNRyq1QZgDuzHY+UFJ4fTDejYwC4LkbLgjEX2RMFKsdIu8
itqkKZg8FiSVOIjpjwPWh1DDWXeR4nR9ZjRHWfB8670FS2thBJyQyf6mxxUMAeUp
jRIjgQkZ8J+CaSwTKhpkb0T9FvoPZoEgN8nfjWGVWhp7gAi/qxi+cKDytpc94clV
RYsjE7rzurM8tZcku3JlYTVOfn/Mu/lvQxzbv/owZ8qZWJvCdE7p6B14gmIYO+h/
gcKWzNjpcX36ePrxKd89zaSLzwxRz829nJ4NsTz/vbCbdpcEll2gpzfoOVCa1G0R
fYTRij4vLu/k9tvz29bZ3EiI9T2MarcfqKysSgHP35ubMhxPXu5WBI2bwhszCyBQ
xN54JbQS8l8GB6+eBhiwZGdXMCnPCFS30wazOabbdSvbBUsp3SiVvHzKTMaepjng
7s8V0emknvCgtPNx6rjaaYOcQWE1RrMXM2uXPdgsFbJCwO/EK8PBQlmUNzmA4mC2
msA0jHRUYXw9ZWE+jXHldI+aWTHIHsUEQxLPuLj7Jg5evBzO1SZv4z8B1y1TIMK2
l21ArexKMfroUPExYRAycJ+ENGyjkjq5Ibfz3b796AS7crbZw0DnvplF6/NXo8pQ
g9Cf94LpjIa7/tUqctXVvTrPgpWT9nrT1oduB28tAGc05U+NVz9AdRAVsrjXeQvE
6ybpGEbiaFCy+FRmRebC0Strl5//ivWgEElfaWEhPjcqUMTbZMI8gUtRXJSnAnwp
iMNMO4pPG0mDU678ZkzWwwDisBC0MZ9e9JeLzCz5HgDM4D6p/7oQsWbiWS7lggKq
bW+uaqesUS7mf4v8z68s6vD+/p61GS9LvzEWuhYFbZyXkj8p6CkzAx0u+6r8PFZh
ds5S9/z5SHcUP0HlMlWhZWtYXrkee+oNKckGhQ/vsTCTQuVFALFk5TSpn4cdzZAf
9TZlRO8akGkvFwF+GukLZjIBdIWmA9H8XLljvqcEeRJz73McZ8Vq9ARam+cwvRyE
4USyV3ITzZrBWo/bU1/SAD0ROtaSmBsxPkAU2nCr+UdJCxCH25UuudVkXMkNJLzQ
fZ6oafnyX7rWrG36SMwMMtVkQYhOfP8zFI/PQvzWArc4YsaaSkkg6EcmxZnFsqVo
et0g1UolduvcAvQIn6Uw8VA2AsNzz4K/l4gVDb2TOLI+N8n2lcOUtQxFfrEHFIrJ
PNVonZ5V6awnC2jMtzR37zZPMQGoW7M2/4bVQ9dSX/0oVzEdg669IYxv3BqtUye5
0s7Y9p9iciKRsHXQBmtxtwfQEAbbb/KJTwahqj8T7kJABLVz8eqSjbHKseiqcjwb
/GIjgwPvML3sUBWakdDy9pytEEXGcmIiqBras1Bky7C8bPD6YuRCsr/iaIVwLIvV
L7LGjVIbbu9PVxeC6H1hjoaM8EPHfvOBQ5hzPTDjyXA/8E9PahB1cx4AV5tCOgxT
64anehh81H82UjofUMekvLBbRQmrUd9D8ZAOqLtIIhT7KGqGkSaBFjK61UvBbRxs
O0eMEhd56pmFr6pD8rJrzmB59lXiAYCnotoVcZtDAXHdzxUR97C8F5lQyRfIx6M2
Z4C+738DT6oPZeNPTldg1xVHbrmU8Bvx90rmcZP3LQbOxzkbd1HeHnI/TPUDcFvT
huusTN4mxG28ZfxTY5ybpz6CLR97VqP8AOqfJBi6M+NE3zf9dRh8hk2keNabGM9k
BRV9HGJixWO5PgTLgmsMLZmqqnFXxF+/kLSZezRqwOdF3mFePgtaNwmp5aUcpQjL
MP0Cfar3haboppq2RPB22MJFz+aYqkFj5vV2r9pkiMYrygfkoGCpppWAwVCWW6JR
1beCSivlktt5gkgXzpHE/RxF3BRDjTR3tCCrLrdI9liAUV6cTikZRTPIJENi6b/8
t6v8fUAITGZ4t15H/GTwQ4rSIoT+voI528B8yfLXJifudURBSD1u7qNhd8A6KlZE
h9eBR/hQmPuYyI0nLMVy7RmOSn/3LvRZDIl/8Ilfufw4EkcBJM/VJ/fmwqU95CDi
T+eHxnQm1OIZEPl4MCVzrti5Z4CJRu+HByYcBdF1pxKBhoyFs+T/e6R50uvahMKk
frUiA8o3WUTOlMaqRCGmBqi27oFV/kjmJFEmSPW3rqvBPwwt+51lsc61VgNU9VZT
zwxATqrz7oYgD9fsV64XXCG5FHkVSjKH/DzMezrXuOudtrZPoHnjVPsGnCQ15V0S
rMKf08P/kkLapsnGKmytBKHSiRAyyITFGWSsg9fjcStYXS0+VG+JX2SO0y0ONjKf
vFz4702hvxHYqOzZ/73iwanEhmAk195rUJYhN356DddyQEewq2jtm0fQZxgIchz1
E/LNgavz0Hg0oG49qxssvP1h/BlRjpMu3IJqqAnpPH0MnbPwsYqIZle6qqCZByXI
JPKpRNKu6lbEkJFz8APJPZy4X+SSWyss4B/+s6RdXLCx/uY3uBIWOiAtJKoRJRhT
Ehz1D8v+dytX2Hp869spqhOcTEMZt5OGVo1KYUjTI1qJ4x9xtwTegkN2J/+My4Pl
cl21s669bOAjunO5uoD5PkZu7KBzQ6ZZchtSgvcdm+0DicP2sBsxI7mHjUjCrEf0
L9gFxIQQhFtIbN9a/PgEKQlmcNuxQUqbGLpOc7rtAlyXe+VHLYxW6Smu9t8Y+xe1
wSL6Y26a4Th1if38yzTqZAQjkwl6bqBEzoGmeqkndSgsEyVWBC7idE16BlQcFHZJ
np6Pe6nS0e/koZbTabXwdir1f1Go/sYR71uhVDESyC3CsDe8nroVnXeaCJe9RD5Y
C72DulETeXbjRHNNoQaLlrqBaAgTbSdBdmUph9BCaL29S9/7f4aBKAf+Pg/oI7Tb
jArofHuesT1WONyEK0dwdRbIv3F3pdDOgbLxMNOZ66o/JjaBsqou8eeaypv059i6
FQo2DAz96lpeyibM18WrAF9w/P/S8+4t8lL2I/4R4AUzYB8JsoRMSvZVWtVE7XDv
y1faHBbc0yOmdZA3FQovuNnl4zABH5vQety8Sudshb+bw3zui058PgN4JbWlioyJ
jZ33PVC+KTdbVOfVut0AwhD7qqz3JX691sr/U25MQZC1whUGnROWnTMG+lhID7ES
D36/4t+UCpgdG4goOnjAzwF9muGRRCpbjeAN2G9E7Cyi4FEEPeDaXZFLWav5WMsC
Yxj13VYtz/OpJLntilgF4kO4YSIf+dn/Qgxg9rCjnlJubOo8wjXex1tv1orolegy
tlarN1IwPhtrVg55tdjyJ//CGBYy9vvkND5GGjgBN/JdyqXEqEARdce2f+9M5yz1
bsiWnenv2wGiOmvvySOH0BljaGBHANGEOZV1RMISq3rM2tWKVD8fDxuPyeaT7zu9
dQLwtzo4zEwQT+5MpM7DdgjUR6X0bOXZtZp9m7AsW+Jkiasac7n/xjRf27AvdEzd
TALPJNs2JTr1OeqUyWQJ9LTleXBdk6Nr3di1tD6ndamVr2HrRRG3NIlH0S+DkU46
jqSu0kVgdzAyQHYZB1T3J5QVlvzEZqRLN+G+EkqX2FsYxZVhExTHZs+jZ1e+CTOG
MjCjikm/BBNHXBo1D5TLr2g7oLa2K304/5U7DlWrtgE0F1nKs3/GddO4u6pvQrML
VOKiBH/skNVX3R4QydLr+99k4KFx3JA0Zqsk4BSwp6zIpsdg3qaUmidV8yU9b2ze
uEe5SgtUQlUsFY5UZfXmMGvu+opfyUwUc+BAaepSoMqYvgdsl2mfd/xMvMwP6OSh
aXjnLxEz7q9S8Mx0X7wZ1BLT07S2aqLhj/5shImy2DMlAlIuigqqRzSW80lk0thg
nhU7/Wr4IT7xMrPTA/e0E34ptuEEHtguzNLG6dgwQvQVXDFmN5QBRCh/4XNoeLeQ
raYx1fr/2zv4/aRYkeSqy9sIB/yYNoxPRX9Z7mgw+drsrXYOJDa+LgIUheypsRQk
4PdBWUrNhPDEpiTy/xEGc56De3gMUoZxjDbd5qinPjqr/ZV0Y1CIqbfQJH1l3n4m
1RFhvLN2h5H6JWh8Hr3isUlsZq3qWOBnoOg6fxa3JEE64nYaLTXmVEkTqEiPpx4S
xCfpTvuXu4UVjLmUqLWUktV7ptS5rshaOhpUcNxG2j7o9Dy6udeieXgzzRUodnVO
FD+AaU055NiRudE/BVyB4SVipVv+7XOzS9PamoUI1wXRw3+Hip+ZG2CtwqPP5oru
cQp40wP2cndTm/K7wU+HYmlGovJHvXUGrtq94fmJi7CNcWRvFIwAknJHoox0K4uO
MlE3Ut0K6Wo0H3gCVpl5019s08ksWeBDizoJjVs/kXf25p4qFVbnHDOHfQkpCmL9
6MDGxBx4T9qlfBZussnRp9pBb7B9Q1w1zVPDoolDNRmN/myyv6YNKCIGG8FoDrM5
8vfwy89GdOJvOmnXjY4ccklxHKarKDsTgc4lrRPNlnR8gt8nihuZHHIn29op9/t2
KS6UoZWABoHAMU8fpdd1riyg23a9xNQPHptke/5Yz4V+nvYaB/FRrL8lt0gNXwCh
sW0sYiz9PWkO4qS4Bu1wdyDzO9rI0cnYuzsy7yqb1nzfM/6BSUG5+vwNv8T3YJF9
6AySjaAHR2BBIf+18tYU2Ao/eZiel+x5CBBS8bTS6bBQQMf/AaAJdNklVQcTvOHf
zW4Mm+iYt2v92Gnsu8499pcPXdAJRVwyAk44QgPzhtsBZ2k+yNeSY5N+17AZeIGH
m0144rD0ga1Bov1EN3IM+78VRqUoC+tmA34O0loyghzaihgo+CvE3ibCqE0g0OY7
RMyvH7emZwElUv4cs7+B5IUUmYgbMe6KgKA0U4V+BG/oJJAvDFNx3I1n4kP0Ji+D
MRBwxJLTBvoHRBg2pYsc+gTzKQjpQAKK1+DndSNfq/1/uqXFaEGg8OWMOdbK0A5s
XXkj9wq5Pxh+k4l38jZcqvESXchXWQaI4425G4gEl8E2Ajxiw7daFSSeBvBD44iX
/dkIOHDXfnK49U1+jc5SFiWv+j1h13OOrw0ZNQoKPbSkvQY60v1w0LW7pe+hIGzr
tRtxllE7hoy2pdRrm6d4Inpmgib0ChoYlYOSdBIRYt8TS9nfcpTtm+24JvGGoWxc
apg3WEgeqa5AhWUEIaIn9XZ5ksK82CVlz9mI5EJWD3D2Tbtlwfc8PrJDiujrjBJ8
yJop8oDXR6iKugDqn6qEIKpWb9OZ3Lr32o/hvWN4CmoULjyIK/g7IDjpD3OR8ZRx
DbstlDZ0yjWN93dpiLwecI8rQpGJhEWw2hpoTJWicNBDtPegk0qBNbe7oWNO5HNc
NMZ/XwC12t/g+fn0j+GvDqJV3Jm4BD89RCwTHCozZ4abwUZrnOTRkGOSUxnWl/WS
ntiO3o3T7xAGCXJwz8hZ9ZDmbH9CyaBoIadOfY/yFUM2ZJJMeK6rnRree0iBC6YE
HGf/ehGVM6rRsNbQ2BOTOWiAaBVRAlGhG66rxjLqScUTMyKfWmQezefwoNvu7OJw
PmSfuXG+q4c4DnUtmI2egCCLaGIgzZRgqCrM12jgc4Yz7ARQ/GRuwEPiNb4QoqXq
k0vT8TwymEVrmpjEF0t3ymyj7ky7KpzJLV0oNhtNHkx3HfK6NVCSlLzB6FWn84ap
l2/4WSMHhqZj9ut6zzO+BduXnQ4nclBgNfXRejJAJvUGg/al9fo/obJ7Vpqi50Cn
kPFxzYAsjeTtQ+tiqIqmUWsCNvqrjQkoNIt0QL20Ux1+WUBePz/ntHF6EY4UxXur
z30WSV4eUfaQuYXmcBurScHfpKiCthWBTOn54ZotuWaPQ7cLvYkqp0gUzKzAqcxl
nbvrSgxg6PmkJs0VJXIqju4N2WqT5ni9Zjt8vjpbdrJYRCxStkCMbPlKlmy2jrU6
pnvsrwkD8krFZWR/VmRQWCeAgYoDMsxWCMxk4GGZ5HnR1+Jz6Rjd/LZAgAOY2ml+
E4XPuhGIJUif9Tn2n/9Xk2EVOexTuTTOnnM4HDY2CH4eJhxVucyyutZnYTimI31S
STXKJiQaDPTXxnnCOqvG7Xzb5OA/L4TZ/E//cqc0cJJgNpIpCXL7kNggJNPfW9nP
lJxoDhY7gtGV+FZlhkSn7LjL6/fqcpXT67UYAR6wN2P44hs5IR3FXHBXxN3Vszwu
synzD74/josEGndfdmO9vsLAPiqT4At5xxwKQL0MEF9MHmfJh/oML9QeMLrTBe3E
agsP8lPhCSAZgVol55q1Lb+0AzrTESoY2nltLUp1LdNpMHrq0Cmtg+GX8jr5D/Sc
I9KxOY7SlB8vTeOjRfZMvwPXlFgrkqqlphBjNYMtEbVjzrYIYrWjsLes8feCxpp5
8fpvVwBnWugbH0COeCLmp83yE1vNgVHRpEcVT/Dz6/MP5hcxoW0WyR2FZWMu2vkS
OrZjzLcG+c4dfxavdwY0gmD++ToMmKL5XycC6BQExLmrxox6RFpwa7d+b57HLFyR
6mGH1Ptrmey2KhbEIFdM/vMlT1S165VkQzd27/Z/UUDVfRjuvtwuL6NqMDGct/4H
1kldgfEV3AxNbPiK67g4a4Lf5LEuQkxPDXs/jL6u2hRvD0JvBLI+Hj1Mm/gxlfyq
0MNB1Ifdwb5Oukh7u0jBAh5I8wq9rg94ZbDn8kr6a26snZF4+2U6x7kLpT2Lpwc5
lxrJE/sZrbmoyKwvpZw0VB2NAukxFaXvU0IAbKjnKpfCtCdUxbm+FJAYlZlwKTXp
vlOWNwXU9E5FKWHdXbstEyLUxHcVttZX2k5pEwKiNo8UjH92CcyCbdv823vjRw5A
6BemKBRrzxW55uoRJRxQVTFAfbtEHgBpaYwxOsMI34lUWB88o4crw03MgL0sRGCC
doARU53ciWbwRjmmTDlGuQfXt1gqwdazsOcVvpmfsalYBdDzbqgrWwz/Ww+oemqr
AmeWy8ENBRJ4Vefmq2g7GVWb2vPBCWcreMFtkfGEm3SoAXrJSuQukE9MPAE7YY0Y
NGA3TInX79kfAuABcve4lE4YQ+rSRZKmd5jemDJ6v+kI86zscU0pIiZZ8lnKsBhW
Bu99SMENBzQgZxpIyJmqMxut/0EarsBnT4VzbbIDvGntaKJKTs0g3HvY1vjUSYDR
Y6/HO5HR0JnVAxHlbTBiOlb9cQx7R2vcWspKInwoFf9q8CycF/g9cYpsvk21wQOY
A3Wut7UgrS19tC0yXxOdaiTcn18TuVXsoLqCLEh3Ygjs4Cc/GeX11uN/Yg3P6P7W
0EdNSrO5gN8GOFKBb3ahDbBHl7+olehH7c5VGu4L1F0BIV2VvgYNwfcoEDpcVta0
kD+IMH54Bl/rs9GAXzH7D4V1epK7GwmJwxc0/79iNQ00P2T77XHNvvwJuE16sOM1
hPjMd+J34MZF002GbZAMWZgzEE5KMqLi9EQbKCzfegrSO8v5KiR1/Z1IALEhU+Ly
SwlLoh7PF1q91bVowJPs7Z804R0nnoQ/gz2HN9gzi3EWaOZWQUYF4KoV3cy83YoL
AGCma6xmPqH4A0XMA1AX7bSkWPCKJX06pI5ZvP3H1JyNgZEnGsiUXK6xeRowzYTZ
bYPEvMsHYl59ybA7MeqJBVOgH13N9OiF9RWp72+3mvrqCsj7VOingPjC8E3H7QvN
Ktoj1IOyK2sX4DffPW1t0wrOYqCZncG1DJExfh0XKrycyW/eDWcx34+qRtjgyjLb
612CGySe5RLdWcC/N+Wsc6zcFz1UicU6GriyBj7Yrj0zQkInuhIktFW885vI9OLs
zE3k5a4FskjT4twTP2UztW0I/asgsd2ttHwbEbRjagEl7fsMAkf1DLksmfHWf5qI
xVZQGdk6Nj0ony9hCvf4JieNZO7+3Uj1aAIGNiGJvgQs50tF3O/nADLKu7GlQhvb
+QByiws2c9hZOmHw6XNcaAXR6UGoxMVze/yDoWrbOCekXcWVDfSgomOgFZ8r53V9
vrH2etyrz8hMAFOph318rvyWDpGQvxgUO8V6QRruM0eLrFrp7xuhQBOvffx6IRZE
A0rfmUZ9D+4ZmR/3UDE+7RoKEivQRzmRE+l7eLqyagXusSHc1r87UW9F3NtZHcdy
71lnV9Cl5vUQjwtSo5CA3cim+dafR+qNKp1gwofV9ouljvkoKFtcJa5TsVCdWH1h
GrN4duVCwET48kPmChmsDGA/Nwbkk1ndEJ5CTooX0fbRagjvi52EzCCQYUH4pK0z
AVkr1E0p0IzT21L9WpqheqDtrcEbfar8Ijihyqu26beB4Yu7cbMdjaH2jRZ3nCcu
VMLT7bVwT3rE5h3VlQpqvo0mYl1P0G6GBpb1lIJ9M8MxgjMQGaRt6LJ6Gn2naHEv
hg5cIAMpdZAUqY+nwMhlUFUjfBcFuHfLkqMtz8aiZcGNzhUK+iEqrmd3la/nGsE1
w9YyTYUUuoe7QIuHWgffRC8BMIscSDrYOCbhOJp0ub7gcQf8GnGNPbFXxLpmeu+E
0IkuSVe8/zgIKQyrepH+4nljgir78gwEMcA/Tz4QkDLY9VM1QMhpBEXnY4E9MVPc
6Ev2DJDSLVbMx/7/LqzRgoIS2uJeRgbUt/zUe7rKqZhosekcwLonrHwfSGVBpgwC
7eb3N6HgM2SGE/ATxlFoti1BC70dpmpcqWdmxKmgZc1tMViHEIIUR9Haa6rf2Rlc
JVFtdF79YcR+bBmGB/zeishFi7ykZV6/7Qxe5h2Jq7FmLdX6y+k4J3OEg07rIeJB
dPXh/kEIotsl/v3Fq/gQnmLzffTteS63iP8KLBJYt+aQ8i9/A0bQNe1lezkhzORM
xYHLziFeT1+u0h5TLy7NcwQGiZwJxHTA69lQhYS4SAFrcDUnM8z5kvI0d/RV/qP1
MP78b3S0PHqS8vPEOiOAlGsiYg3DDgh35UBBMQBhrhhbtj2sk4L6cESAJr6ZhzTN
tH91RKEGSQDNL1F9AoRQLy1ZSpbigRVFOLYAnqZR5bZ9xgWXT3vR8HgbcxJFLJwM
HgpIwN/vEgjZJbQ2oRN4rY4iidhQVxYpKG+OkzCLZIs+xH1mV1iDl+X5B0DP27nn
0IV5LC3U0uaEYBovQPENMARY2lr6o7GkkLilKZn3ByIdaCLCmN6vn6tnaRtXZKJq
Lnil2DCrF/fvOZ7K/pyx6xW2w2o5D+kJwL5TKE2/9VOaxpLvgu2bY0r8HYIMvGfC
CBejPomgAPwGrFJn2WhSLwiVMvfALevFB+mLcpl5iW7LTTrNYuHheLsZF0LeHIo7
X0/WKOtoyvsOLVUt9jwnyvLaYxyjUfB2xQCV29hk5NCQjcMNH/Ul8XR+JtOW8hLW
6Rs/roM6PDiomeJcWkCRbttcfOLrOmg3FPoHrxhgJIiUquAvdTJvQaR9kglNw3xf
wK5e4OLH2Kz70K2s0R4iYXUJ+VZnnsvabYrimShMTV5Tdhl2md3gK2Vo4z/oq90D
Oe8VRHjcsaP3S9beAz98nlu+D51VTbdKgWIMm3K7wT6bwjcAhRAhjVBaWW5t+ByX
UnLbgHVjxU7Z78zbGfoDe8dLIcQvG/8s2rbeD3ez4CChyDX6tS1T+rvr3+2x7hxx
swxaPGzSxJmkbHWNi+5gkO06R3w+toyOtKJIjnsxVuV2E/G0c5HunVDjJJ3iCPyg
lz5Cq8l15ctiWRZ9Cv8J3qdAH7iIs/AzHowGIAiSfhkRarQu0cJLrGaM5o8tj6TK
+RO9RVpzktE+ZbodpSjRoNgDa/fdL2yd4Jkl56Zz24BzoyFcArVj72anApTWHVAx
o5zctYMM2vCTZjS4xzj4LNEDvRo4V5NeTzASQtIcfTFfu0r5P7bVPngHPBEUBAA8
8roEK/YOg3TYvzEHA2MNuGmNXgO23BbPjjDLk4SAYtbNXD4OWXBXqHL80pmvO7uo
OB5k2dr0QylDmVsuhOS8BuzRb/vxdTrTLJsh66XwwLfuT3tQ3kimR6k8gSHt4ceZ
qXIcm1JrRkrK04s4aFmc/mkl0Kz/pOJuGxjKm1LV4xTnZJbGaoOzbN/nao2ST+l6
jp1txCu5hRkAl7vqhnYoCgqNQZ+fAfeuA6jGOmwpDNVjHX5caRvq29ljYyLN/WSH
XF3zrYQZNCR4JLrUT8HwvgJo3qWMiq99Zg5tyghv9TN/V1VJLWN2x8jdyK/2qjBs
gh/gZKd+wdaEWyaUSnrMgQBMDkkjyKWmkfVWWx07cgFvA684DAz2KqU7m6dTHJ8j
whZSfL5JaFfObznUlA5UYX4+gCmHKurr4CIJaSbQm6XIwyMgJJwga/CGGy8lJifS
EsbVuN1QhjDf5Yrf2PJfKVrmuZyTH8/7PZ1myC/m4s4byTxjQHZ5oHyyRSvq486o
rdubd12WllVZHOoDJGHyL2IZ7UyUaeOF5l8L3XdgQSc/31DsgTYykcNVu/70J2tw
BxQsLQbeV4gz625SrGHCvNzlDP4qJdxXB2G8FQ/d1Gxk/d9WDPgnBWJ4KTGbL2TT
cMOWMHrJq/OLYH8Np2z0xmB7xYh0ue7aRnDgoEPQZxwehVWG35TdUblXF7ys7Jul
MmAqnJvxavji5Fg2o3rCRbZtmPQ6DrkVUoIbHjBr+t6NA0gKEiYWALvjga/BQSoH
qGQZhQFIVC3gOwvlHsVkHGYUWUGDZQOvTq2QP0Q7VKmH+stfsO9YuPOBtYqhwAfF
eXCVu3GCmzUjv4JmBuuaqEF9n9x+BVlLAOs9JMWqXaJc3fhbigj+yZ6w59A9UqqQ
ZYwykcWMyrmLBNJnY97y4fMf3/sJV1CcRoUMfsM7iIJ7uwfk9KwZ1OtsEij1P7B/
Zl9rCAY+Gcfn6VMTLL6bsEetbIW1X8NZ+mXEdHQOZGIVO8sQda11vgTEz2X1W19A
lDo3OYRNnMH8Z8d7gq7Ix2Nx3DxQIVXNksOSmzAulP2Ffw2OvZUCRin/ZEujPrdC
LO87O/vKkiaM2VUk0fxMoetW5Qn8I+lHBpqUV8y+X2lGu2LfhmOKYjE8a2DP2CHT
U4kOTVHS/MsYje9R47BDWtE0uKohr0A/pK83fZJO8FKla8KGLT9ZP0ctjDUffHYH
vnwn7QLowjY68ZPEwWsDRxorbjpENaGZacnte6mk9QotG6xpQE7/6kYyRTpjC2Fe
MNeCG/Mlufdj9WcF4joWd5MZgwkaoxdDK4B/+OkafaF/tNOkWBFyGa9fNCmb5q5Q
q0MA6JoA3bFeH6R+Etxb7hvS/PY437fejEG58maMVVbonI3Gz8jAItz2uSFXc4w+
GloNy1xsosTzkhF+6oBklz4S/jLgPCxaVAx5Bd/u6maYLhSB+5dDaN6LtZkcNJJD
zMsnR6bEIlwZEChuiuPcJlbAlF2cRcJBvZ6rBO9XeOVmGbh7wifxCBiTyKUjSO3d
OT0uevwiWNaOj/HQ/UkyJ/LhpyTW3oaeJaw9oXJmc6wyfb4gvpDtieSVQ0giaGUt
zAf6a1Qo38KPwq+Z7dl+i76Lg+SV7JbqW9mcm66Th8ZGBUsN3zl/nuw4Ylu5g54k
Gbf2uY3UucxRl+UEytZ+pQ7SC/X3krRVWe/cV54z8mlIcdptYinuyw0vlp59ltUD
DqwUhsQWXDjSgP+ZRqIUFAZrZd5RVEDmQmPXvLE7yHzr2+Jgamh08WXenEEfogeS
K+ZWR07K0VXx4z1iFbsfOgcyCcpbDTODlSJfoPQXFJhEnCjC9yySieIj4qbIm4pG
hE/rpMVmtbyYiRwxDYeuxR3niXMRZR8+qV1RbiYm+itrHs0Oi6yKZWXqgYK2lmdL
2Y4nH+Q5tUn+2+BI6Yhxu63NCURnJUZ/udC2OrQmRjAPsqjxIKWgpdXIuKWTJNL7
3IcdTFhPPaB06Qo8o+ZpHnDvyZVNWYbb+jWV09pdfim8DEI2EMUo/kHv4NQKYEO5
ZHG5hVP/WQjZcz1Y8TjkI1TTK3wFk4hCXZ6cDSZUnCliLZOqcoCWiI4p14aw3DPs
OWMC83YiJD6jniU4ou18KNrMITtep/o5LhNJazUDHai1Wiy5M91t8Y37YP7MDOiv
40mogb8MQE2thcMWy+6hJ+TJZ4V6uf/sc+C1ftrMNSbO0F/D7txazvY9PRHIu4P3
CdN1uYn4hND599qVVM/Q1jj1Tjnrt3CeO7+4ZX//efs0A4VH9HTvtSorrDL9bVq2
UdLFKGCEdYCNCdgBPJuWnt6/wyd3WxNSwq9hejDqIJohmQjJfHEzqf592bFWOUq7
r1I2itaXyipZKcUxorNFdb7F5rvDjBebgTMjCIuiTRIrl+Tw185gpF3aj1z+Ai3O
KztMNtEkASsHHRA4eOnTZ23g4WESNE1F3hpgid1HR0WTwSpsl5Oa4dI5clFCjoPp
sPfHy7UO0worxo6YXNglSJqRWAj+pB/vEG+mnls3IqoTP7ksI+reIK1TbHfPcT1H
BHz5cYM5qpNC+jiVVIPQlr9R3mJ4ceByHrga7JlPful5DeTr5RI9/5AsJdMkd+Y9
OO3JZU9YNSZhfBjB9AEBz+yXOUZVkwyqM/RgI8r8t0Uctj50T3xPdqaFhwPAXGtS
w9NW0R0u9LTvlsqxHNMS80v54sd/I8MONhpPhwSu+/KEhYK4DPBOT/n8AM9Cc/Jl
XWo8kBWlqlP0pmi1rwU3hvXSp51Uf6wQ/VW3JYlFVr8o4reg8WJ3MEiKSLKWYeR2
mNXTdcaHv2GcDlbgMIviUh2YfPp82PD+MR0L4gsR8FJqMbfb1mlmpoFAcUSvvMXY
Rh30XN0CDDRH8g37344xe2Xk9u1SwOcTc2yfcjQ6PLZ/VYbNQcv4svIMmxAPB7GW
7+snZB2F/YpJt2ztgaVU6Owx3kBEgiP+7W1vcoI+7cLdZtSicq0RPysbLV9dg9kj
M5TcrluKzM0pKrh6VfwizoYHqZysaUk9Qo/r1wA9lkVCESwyYrqApizoMdgsv1Xw
gMteRrKGJ+IFRie2pxjf+eH58ROTGOv/2GXm1kOzZcK3KZ2rVHBfwxrUBWuXcQn5
cyN7mu1HK+DBK/LMdfXV9cNRTKiXdWWHbpa4l7hkljsTn8dD+g55YBboI6JF/wdV
++EgJgmGnogvT+7MxNlSD1xO+Wu+EdtTi4IFHjBHfoVD0hfkEKDqaOgvIGTENTQY
+PqKDh29BAwfLD3e5aYyRW7fAI8m9A5pTdd2Kjx5tYQDLZNuQGUiCMEgccLGaOUb
lwfC9uYl/igwEil430iq0xpxUBuhM5qVxDq2J7ifS1hdgdjBQHkWyeto8FQ+5wFL
/RKcbErmXp94T2Tuu8WZMNyO2E0pL9eQPUVse45yj5DDYy0Fqje7OfGZZSsaiFqr
cx0FKoz/ODrVUvpku+k+JgVzzbnMvREdBkUbPKfDsvdsCxCsDwqrGJ/sHD5L/MP+
I5ZBptr/qu/cdGOCYoSZpGKPVsuzKGtaAI+7ejl4mNki/7uMmmWIU/9ceJOkcZ2D
XZ4UDA4YFQZ4q5wf8D8eaWV8+CKRLxgDVSvDm5m2AFkcrPT5enm2JB5X6Y6WOpeo
olvelahYxOOAjlb3uSzXEPI53gAyPHhWjxUSuOxv4bRF9X13W5OJ41bO/1OiULcz
z3C1eZhKBt+vFP+uOC+MwtRjLBun+LFoyv/AN2LMBj+gs9ht35UmvCvYshgTfDQU
J3TtezLyLQq7mkhERmh3Q3SSuKswR681i1f2OmmtwyhvLgEKLxm3rshRlD8UgLF7
YR/Y1ytC5k+/9/e1Q+cVmxzyrGREon9T9YJpz8VA0hNcAqvdTj9EcwC6FMg0I+K2
fZDVHdUDVQ5VuOGjIVR0mLqCyTKvvwR0waIynl6Z6j38MPmTl/iMuyjqCYNb/glo
w0WLfRfVSg8tj6a9G2YnyaXTsl2MLtXuUVVAyaK5vKuP7EhcicYEHLYOqZDAloY4
wwmYeVoqHO03HvGl3LcU7xQFvjiubDy4a7zzZ3KpFkkyRXMrlty6FWEbqL1czN9G
u8dvIYt+TI2I5lG5Z7xqx2KJq/hoq7Ergot3XzM0JflPBv0DrVNFkDckph32foje
WNagnWbbRQ/zf8VF7GAzZJD1nsGkKEnzvBt3OBvLSM6hQEqW7PyTc2S90IKnsMJf
EdkArTVcqMZbjFZ+Rwgb9AWjjLPUpDnc4PzU1PWv949N0tzesEFKoN6aJmoez7GZ
syrCyVUsaZMGoZKF8s84BFZ+iAbfxMseTI0hhnv3kC4i+dIl3JpAxGnqM0U5ROVP
YY1gFi/9uNSEFAXnAV12he2GPZviiFvZe3LhNvmfuUjCqWMj7fWQGvzzonXI9Hj/
XLz8kP8E6NnroE0AFM1SL75tenKOMc8bzxkoZ9h683gJuhIxlYq2mj75ycjTHOqG
oq24Q6N3aWzcoBHQ3myJHN8kC13nLbzP/BQJQnjy++XQYxYrxrt5Beg74EcfT3ha
s0zlU/wPArr4nNnLsDriMsY6ie3/lJOX/fE9rLgy9134GCu5JppTGKmJjEyvLPog
UNiYxep9hPMCqvLK0Y632DpQXYzq6D0cStiWhG2UvfxC6oFUOxMltYl+Umh7ZmIh
f9HVLCGEaLFXonKSxjTmpM1saTcl7znbZpzUwUznC1XhBRVeeH1Vxzz697972Qe3
pbwdC8YTKqEjOVk64nF4WsH0rsbBkNq/OmOpSJl7N4wzFKC1XdBnFLHDJsIMU1uJ
8IMPkWsvAZhcxenX0oyjPsPZNwdaxRyemUmnYznNmuQ8VjdBZikJUW11mBiGp1xy
/Qu93JgHCUG9bDOb1qXqweiEhKG7o8ucoiwwhk+MwuwAerGDJm6eYk61tkkuypCz
WyaJbs/xiw/kPYor9fohTwWW+3K3tTOhb0f4F20zHTQRURGu3hDR0dwFSH9m9f+b
ht/+vVpqYUOh76ERV2OL4W7X/iXcAjhfgxfWY4x8dHnzmilUmqxHhcxQ+6vnPPM5
pfoFucgz1rlxEVqUe1mlQcgOyCXNyaXB5bAX2y4uPnSamr2pSenGaT8+4HoG+wIx
XTwc+OI1vDKRpiwgb2zuVYqEjQgFiignQFYggtWxpfngq0jjWjp4e09MlPeoLdLm
G2K6NcDrFvXOuHouk9sQd6Lm2hzior8NngsD+1UHjJYVbE1pqVed0u3Kn/okvy9i
7oz/t0hjb+dBfSf/AeFD45jE0CsFlWUXNR9/egQWi2HXuN4NdVhQwOQv+xj1Zdv9
wc1RWF8mlHmupSg9/vDHQWhtUSWROdjQRoSLFz5odc6VtKD79LFkD5xSEfUnGnFX
JhyfKYr3ObhTCNq8DwcI7CvuN3mfdIB78F9HvYPnqn1iygoZDegSgcnK6EArdKBG
0i0m2jO/91G2Vu32fkN+LcHftS88xUkxIYC5YcX3p+V8mAHryV6ORAMFPtRgE2zM
b4TaxZ7evPkKjVOas6zXrbxubuEpxjPm5cR2EOjlVx5iuhNPwmr9S0JPFkAxuDBm
8NE25HzLobRhr+2ZMkHw+vr3U5D3g+TX7wGxPe2g/tHODsJul6WAEotYLwkYjyDg
nj3FUGg50qe1LUr8amDqEk4O9M13KrvOFe/tSDyYZSHbr/UXqWoQEDap+k5djbPO
uQJ/PzEZkAobJ4PjJ2/nP4MitAi0QBNSf98UFDlaKor+O2coYYFpLLYWPOkwOlXn
XtWSLsm7+XSaA+w476GrmbXHWUwYSjc5ZmhxAQzv/vA3jK0c5FzvEXfO7+BlTvIo
ovh8OxJhJDZP4RW+w6yW//bTm3V2LUouugQ9KdvBv4e/x6bEsEJICMbuiHDfawpw
DuMUycx8L0e7xzqgOKv4mP38Wc7yhEwPrr8GCqJQYiW4CQMwrbHdLZrnRTqQMDWG
ECNFsW5Hbokdu/Pe09+S0DP/TXkQuQRn5wkzHTXuBRmAhMScraLrhrIwpORhT4QE
CRWWjO3ZwGlVeD3F0qU7Pr1aYEXvhWuHFY9rM5dIzWd1TIfneiyptxvet2W+jM+b
Cttid1Lfbm7ArJxPs2hn9QLL/WS9G3QfsNECGgcdZmFKGosrw4Ka0ijYfsvDlLeH
uxBu5cay5P4E1GWSDVnE4TAo68w2yqWIhB1JLNdcQLsEo7SXxnk/yx3BiVkZ4wKL
00Jq+sMhCmhpDuEqWUMBFoY2RPzKhrP3IHNz7AW0wwgm4y45cL2jIBsYXxwyxL4Q
77YybtReOHrduyyneyB7m0JFJ+8hnmvqRgDrc3/ySnElk1iHigJ+yKbmyuvrI16P
G3PYCidm1gKNZoEXaIWcGTtwNBE/wGhEM3FYLy1qeLIm5ITKwjpFOjFRQc6ADJV4
sVJD7v/gM3S8KRROTO1zy37qT7tuMakqmOJdaSl4t60Bso1fLg/EuwzX2+pTalVV
8qAoQ+cdpid7k4I4HJaTfSYvgbAWwM5TA5eMeDzrMxjiEti4qztPvN0XYV/VGj5a
3SpvzX/NhYsgvQlnusrCKiN8HuZUY2N/4XmdNhW1whnHtgR86ZY/UyJDx1BEHQ/s
lb5MrECD8RR4VINmJ6wY57cKBWbrKoTMZhO/4VcQ3pTmcwSJh6EfFr8jw/mLLgyS
Qt3m2JMPX/QIsre/N8esr9XbGtM+GifaJob0ooSFri+xYbnFPliPjCliz3bTl4MS
CoNcbKzhyGYHgMMH0+WOf7grccQKcBnMsart8gKdvdp3X6y4IXl1+1FccRlNbN0X
gAhPsdxfuLeCiDF55LS/a7bjyjgi9REtM8+vGUn1t1VfFbcTR+k3XeGclAnG8cPa
P0OMS1RoyEOghTAIcJyYPuQoluZsMYFbDF5T71HLcVVfZposJUg19bsgPSTfUH+d
tzQ+1mTBbzZJTrBC4i/xhg32IF5vWSBmtkOZNlFps+nAe4NbeDB2Hxl3Pp9zvlMj
2cSxDdJb2nMeDosr6hTPDQfe7nRnHme/mu7750+5oLnPceJ8Th5RyHKxjRpuHsRJ
87xr9hrsdDfCQmDiNKrsU9/r1vCQ/txGGhdrzGrq1OFAYBuqiaUTU4s1KXS/oxuO
rb9q3v+qasCV/mIYGS7ApkPFpVEfZdnK/m1xFys4jbzu3x1iroKQlJx4d9JAyxyQ
epZ4aYadNFtKZnOG7EfntFarbNknme/QbcHNFow7nojwHGWt85+k9Ho0p6MBKz+l
XHnElFp3aJg3Y69uL/d/fx/klesapwjEaMiXz8JGwlMBkuDZ87fetVVLTqmuqkzy
GwC2o+Nvspju3Dzv3XmYpMSQDZKraEF19XXoN0oY3KWR3xrgDNVj0gs7sUA1jKna
Gn3bfca39+KmDMIbVrW/f9isgiuM76ByJSS1PpTVk+sfuZ+hB5COwwjrTjECayjL
O2IDCDjsKVsSLZC3smTPx141Ts62r02lOzGeoXOvmbaayaDFJOb7B1KGv2OZ5BcY
IW3fgTKbSjpK2OI2gbLuF+8xHpOal+CO2JGwzMWB7mG0DDBl6l8KwqTSrsP1G3Em
nrIFmZBW20YuN9AtFBXVZzv+Vap9I9kFMeSxGqhGsRJvJER2K6mTte1TejXNEkpg
iV01ClPyvECec/M3cDhjvMTOMMbMLhEkpWkkr+19sKmC3+Y2KtN7GkDhKvhQA9dM
eEV3d9qMhrjXfViP1HWESieVqF7sShi93DvlUHSxKzHIyPBmLrDA/rZXgMycHVgq
aIZk5+NeDu+fDcH+frYkfjiFrHkUBDm9PzJwicDQDopIptt4llG1N7z5L2gzW/Vb
IVxbEAfpPVSXn0lCfVECzFB34lFshVTzJl4mcYC2oLhC+4h/K9ymU8ddHKDiDgKG
M2MUBMQ1X+8juU2mdZ52sv7h2BtBIQfj598pFsnMlf/zfYu+htvEKnHlr1RtvSSq
rO+PnsE2hdOeDjj3HO5aL2A+j5ZSkUeeYVU1OP+ONX6kgURUSF4/WkfZ5jM1qn6F
xyLFC4kHUhlVerpuIGHDnrO0Xbjl0RTRWk5lfncSiI7pkj9PZxJyVK0eofdpAQY+
EYVrirdSeaBP0Ph1YnlAKqFhp9sZYtG/QEN39PJhJyNOStjAU3jCLixsrbKmqvVj
9nexTj4iJUv/Mlow4ztHGH+3dTDaIfP2Bj9PKszleASZKkXdYvELsikT56TauHSq
qnVYb0mm4LMzfI9s+qBLfchcHmH8akl9YMtrE8heZocb7yhpSn+9WeUQdz1NQWKl
wEKYPgxL6gStboThEHry+146z+L3bUONoLdCkRZtCrggXSbuJe+JkiNDGhAFYbUh
Hoh42XD1RMNZgOiWceBVgzJX+fOA3Qo+6WkzDjJqzQedDrDmOowtgR8RESvrzzDg
qXwLYr+YEal9NjBprGf7HtowI2KcDb4maKGYm1yR0XKpaTP1Q1SY8KbZjJsus+sp
KJl43C9FOuTvat+0AqWA/Zcbm+VPAFZSruFTvUyF/8qzW6ChqajwWHWiGUxEdQKo
MTorfL9UTjlT8xgKGileSqc5Nk1YbVQ+YIazkslCT3MfLAFQH7lJgOJtn2hUtP+r
awpSe3tdmLx7NixOwM82YKa4OK2225QNSd5aplyUMUIUTdvwycDq5UAH3bgsEM3k
FGBBh+3mUIa8AUdqGnp9uVGuOrBXAZnL0jWYH/LVIQAToughaOm5cf9IAyjTGuFG
b3VgdQqgMN3nebtADivKOtIDR68XNJ5RoR54QWLFblETBqF0iMj4WQtAmBmZJTGq
IT8D98re36+M3m9fWwdhyKDZ0XtoCnuezfYQX4l2eVM/MSxGXF7gJJ5DXItl1qde
AGwa9eHSVnxILx5ERQ67Or31EX+0lMCtU2K/D1zm/fA+cI19+Wsbhi7YDYTpCuJt
XALGsiwhUooQ/SOxmzrjdJXKgpPrYNlgQ2TTQ4NrhTxH/0//02dVXiLF4fvEzab3
8toB4azOtV/WZ472udVJHXUv9hiuq4Xag5lNoDBVHPTcrRWARYdPAnzPJiDh+GXJ
nPr88zbveBu0eVv7h+bSsabe6kaQJe4Zh/U4NvJMMO+XGQ/FNdHh5OiZ8QmLTK68
XtUAZLbETW07+jb5lj5l3oXmMqdLthVnrVJH4w8qghTAYSRlZMizYRi4FFrOeKN9
2KgolfbLmAviKNOrOkOJLul5In1WNv5EtlKokVA38dDi5F0/JwUiVEz1zyKdqUM5
XQy/erKIzhCV5JqYUB606GPWJNV7ym/U5p5n9uZrPticgVKLQQJJmNmvCnrne3SG
OlsAAUyNrlHEaaa1QEOWelIxA6P5lF2JRTCH77ld3EgXMNwL2NFwG1l11DSgn/Tv
fX5pXT2ODI7lkDDaLxiPvVwsmkDvZbCtc+Xcxh8Laje1pShBu728lSmzG7iJhpo6
yp/Vq4z8h5rbo6ddJjfmaA1g3q+09+F1nYv0x4EJM5MMAmV0Rr/5VrA497Ncavxh
5+XgeQS7ZivzXeU5Ol2RHHD8NMnGWm9kHv1WNoXdlLF2bTq5JvDHFU6gBEeXWN8O
UQfMm77+9IHlJRRWcVwVcmdRWoHu75xcLFKoT4REA3jEkqQVpkNNspSBrS1XkjDQ
nYrTJrazXre9fERKvkVN9idAdteEmz/q0BHK2XwAgah73qs6OFAf/MPGzwvmvOqd
1v5zljjXD5NMixtbTCoDnP0AGlr1Wo5arsyMg3BBLJLTwkijL2vRXfsZDMqnUYor
ihRK5dg+mK9zlOqykeRFEmsS6Og/cyDoQvEPDnlE3pCVV9aAqFiJzOSPNTNBzp8n
q78SAqHtTU1nVwSL8+7TpocXChWOKmM09asDUKH2Jk0r2s+/BC5fbHSYmfi369T5
LYpk9PdCippjugruiT6ANyLPK54XjIq7wo/vywLMu4ZKkm8mr0XfnwSzUEN96FaQ
r3J6ymHXVb22YkjEYvqg35+lsrYjK+ZFiPuU4g+JdO7Z7E2SXQC2p/tVW2wcWsVa
xvEgZBhMfoFXgkBuYvyRrS3kmy2/leUxrocVdePDSy48k1N/IPii3YHfDG4qyFjO
5Z0SOVMKjtPNzkJsIZPun0V/N9/oRPMR2XuJnW7Bzq3ItTQLtWEv4xX4AQvTporq
9Woor1o+m0o3GyZdQazUrI+mdkOq3eHW87GBZgBWg8Kliax9i7MzX2f5tMGr1BRJ
E5Tgh22/fyrQxL2TV+AgnqUksM1GETsPPo8XEBRHmDgtNUJhY86+fZwGauePV7v/
uX0GlKbkRuedUWXlr0+ZQktfuwV2xKrsKBZVMP+93w1dXoqIrMZS6gDrl2jlXhRC
EV+5UugaIXAibvrKTx8DF6EhH/YqFUR2pDnBKchNC5GduNssyLB3bYGtKJVPOi4G
V3wKxTqJgmNBulsYzzNUv8UESrPEiQlQqVnwcSnttNxiYrjoBaedJF7F1daLZXSM
0FS8IB38cS4DN8XLPUO70ch4SK0BqCDYxmtWCqEqIty781mu1XUToJpkpNacfQHA
r2Fg8otinsuLhfPpc+wx6itrvvuxGJb7eczkpv147y5lfuGHYMxqwUQPPgHUY4cJ
sPyVbd3CSA05MtHUEs/aJcXcG/Tj7SWjrYnQmTZPzgsQROZJXmW62+uzZ4+nh7j2
r2qcS79SQiuvqqQ2rPllqahBPwdjmvqYtcR4MPvTh7r6uW/JthpgIj5z2Z9VErhZ
Xtvic1K3Nqwa0qxbvMAt4xYPvEEM9b+7+u63IH5hOn4Adhz7C1afVMeAG8SCDwi4
ZVWHS8stNjGDwnFQIxhjzKO9GdaJvIPTmIGnnHo26vVvheTQgJq2SIPCQGL48ejz
NOwoeLCs8sRo1p69vHfnmfc4+N6IExIRUlu/Gae0LYF6bNvDXfMRWPNuo6fdX521
u0DpVrtCCMvG7pztaOCS6zi2bKTAY++25MEGUMK/rOuQbMK4dqzgM1hYtUkK4YiE
MxH0hnei/cc2wucfP7WMl4c63/ozMWvsRJbZzto6aam2A+BuyIq/CleBiadVOJo2
hTj+ySRbgxggO+hyGHXvwmquNkL1CP+elULs9WBM99HkZ8bx+zekcXzqN0yY/PiC
91Jhq+yx4mgBA4udc4sAoB59jKxzToLsPN99CBGhFNkW7pY2rwa2MWyUKEphDcx1
NikGH1gM8mFUdhFG8YOQJjecqvgtyrIlixZVTp2I0KdrXEYK0YTecFxylYv1ONAs
Rek4rDoMHA23VeJLJwuvrdHDwfDnYNY7KirQTLV3kE78KKrgyoPeBaHra/KzQMUR
fXTUO7wVubmN+qTlZKziKL146pFvzSFCp/gZmVdIjFLQse8in+sKxzYs6eKsZsqh
96AzL87sbtYPKMlqpAvZwcPTZX5bSD8/e2JUShke5+VgzdAYyy/w7YUr3yHGfxXE
DVQfGG0U4PVEVXnR89dtzI6oacWJeKtYGkfhDr6SKv+GWBLe9Z60O8vVLYataz83
J2yuxyZDxeqStq0SNAu6usuaeA9C5LBwGjbPoCQKVMofAh7FQaaujXVBfc17ZDnD
LUdLaE8Wz85aQ+ES7RjMoGVzqw0m/QRUuIjac4X5zi5XT3XfIweNhHVeRxLPm8gq
jmJUCRhkxPtRjug0uZLe7n3NA5dRI1gFDOJ3R/4DsPDDRNxKflPwcNRMvLrj4jjX
KxG4F8LOpjXJPZOuj0aDln+tDlKcCwnfdBD6BAa4MYo+tvr4EYmCSA5FAMglxoOL
18Bx4NZzbG8NQp2fD9w3Mn5bYea9MgGqldQIRyvS0ofUrvV4bjEwFAzOU5GvdN6q
8gOVMiFYE5uKLxY/q6Np4M1R//Ibe2SAmatpU1MZrFqNvDELmnISXwyjP6w+8UlC
/EyKA1FtKtDNFPMCe/YGpZMK7D1TZZCTDQt1L3fZm8kgDjZpiid7HOQ/Bex/y8c/
ma6vCsN/lMDGgrYT3UO4IBgcfA7QTnkt2bpdjnP+wlN/BZvG5vp6ehjzeGbRVYTI
Z4K3AJltgDDErDor8fGW2OXBPxuaXiHO8QJmE5G9yaGln6gRqI+B1LDmKOixpuQj
UahqcAREcAaUMgEELEj0OcG6dLgAyCMeOsBtsgXsv9U77Fi8wFC13Zq/PA4pMnTg
7vbjJJRg3TRHL720wPYve4eowiU3FCs0SGmed7T8QtfwGJGnIGPVDR0R4baudgs5
UQuFyilDXp+5cuBKYKxCJyvDqbscxOtyQkq7M5leN6gSOnTisuGYDt63pB36WYBa
PNbcV6tME9JN158sue5vrlKa+VUSRZWg3xJhQK5qh9NNKQKlhyHcOdP7FBR0doe1
oGVbo/QaImDgM3p0pP3HsfEXVMvyU40Z/fGBAP+ic1RxvqhLQjqf04hUhQwO65r1
Td0AqFdWGoCvBmx8xzOWBlR4m6RTp/pldp0dUW/syvv/pypt4CHk+ndOky13WQMf
fxrbh8+8xO/Kp8ut4pDXDdDYg+HrU991ICf3AtdJA412KlrHz6Zo7KzZBZZVXiZR
FWuNizh+LyGpcpKikneK2Y678NLAPbIklIHH8chj8meQvdsO98JRqf2wUGmp1qfi
93lVMpyLpFH1tszuCUQwXtmunR+8gR2Yd+0ks5G2lLmbcpeOBUHp7kCSxkbQXo1l
LKUxEIdXU2WR90RDx/Xx6MQ5iYUG2OwtYjB3IC/p/kL6m1sJ2e/cQqQCXEnq9wOC
bJPQdUo576DZHT8nGPBdhT65JqmGuvBYbSMxZTclxVIsN26zP6+jiq2VhzSfl87O
XQi5aEnW0v6LxsY99md46IaADLEUeHO7ume8Y1rWMjW11elMyxFar8+Qjj5J+aCq
bjw0ZDdZIPMRx7HKM0ranRvd8EKQshIyuAicOds65nyMkUBdskID+2gaTDS2Fv22
sH/ZuSKORRz5ZFFskUxKlsOfDG5ilXsSD3VJ70NBcsbQXAYsbS0s8JoL6ZB29Fkt
cS0827Pg/aE3YUvA0CGnL4JeAjoOwsRh+FbGs8Qh655AFIMuuiCG63VSIOR2KhiS
UaiTjK96aifISa1rGPsrtHcuZI6PTju88Txa1+cJLPZu7ql44CzBmt0qMbOir+Pt
10tQQsOq9CzwRTr4yD52M225fN4XXIEMUJps/Li2iOh11Li8q/Y8UBUK1xaAL0rE
6I+/o/Ed+/Ac3fTobkFpLejPL1ZrRuT1EFYCpnOb0DdUDzmqJUM9Ec1l6E3MJ2f+
En1gnS1v15lIHdrwHW6n3sZH8+KaLrNzXA373zpqEDhp+luDXsKzGfRinUMIQCfF
svz8TsGo6GHBX/++q/CMtM7cpGiIH3g3Hw7bzCSdVJrk9l2UjYzqn8fWVSfQoe8X
PM2LtM+dPuuyFEfSTCLR4omFNcwDmfYEyp8g8iYyg+amDfXRN/lRfizPn1qp6wuV
betwNGmmkNNC+337zvbhP1z3XnqEHp9MFNRgJcN0g32rR1/mL2oDoK2a2wbc7KQ9
PumEcPLStJdv07BJOY0AheQNRxrp5UBmNg3so4pHxvHx9B9d+f+2FC44v4rJgoES
+0GH1qvPZUvOsGlIoPSpUJswQVr/2Mk0So4Fkx2mWH1bcDIhgy4UuztAl8jp5IwD
+LxhMZBmcqJ4eBKUybQjjJ8K9mEpw1PsdemsMAlcu/3s9d2Wc86QHi7GzHrtMXDg
xTfsdrd+zHLcluXS7FOqwqGAN+AULeVSJf6iQj8ca9Y72VcdVEgQk4C4X+U6iw5H
x1uGNgau+y888+j2Mtd+C2KuSWoisYZEAIEARNAijXPfEQ/51PStRDuAzze4x2dM
hE1Xd1tWNRDzwjOexm362rh+b4m2yTD9C3D7t6/YTHc0NACXM19JtJxnxqBbrhYY
KGq5BvPFt/SzNE3+DjYpgyzEYg/tWm3f3F5ClcKSze3/Hbpy3UZnN8DwWxptwh1V
r9cwBk2Mfh8o055bF0byP1DnlANMCF3f+ynoyWYcAIUp3L0nn8a5HX7DKMrS1GY/
w3/XcC7rctsYUsNmyVvSUlY3GNXLk9jTeWkMe8/Ae4OZmN6+d/UeaGX8O7Er2QWf
mnWxd4satzyAY18AVE5Q+ftblaTR2TJXoS6epEUdZN/+/5sAWQs6VTki4VZ3sg3J
ukUuS3I67oQCJq3rjEpmneeo4EwCx+93B9XjNs4/DBTgqADiPDckHsNYxdLE1plE
8r9rXgoROtc/RkWBGCX2vRyV9LDYlSzkRK8Sfd+zUYrDg8SDPK3euQV+kZnbiIN9
KEWrrFaFL8NSLxSgmk+YU+f/L4O2dvWE6OfX5fou6jEo1BZGBhqLcUnUBDDgzdHU
wZ7lPPzH0GC8NLBIJ+/l9BgyMhJxFNLSh3DBc28snR1GmYZ/8gLsQI1f1ZfraN/L
f9D2clDTuI5HCjUzh9Rz2Xa2PVv7RUOAMfZS+fa88RY7S/ojLuN/QlwnR5c7xmnX
5sNovKzB/G6rk3pEc+YFZo3v4A3QafaDr7le8fz10DuL/ixKfHAkVI0cp3DxXXmv
jExR4v/Cb82j29EPm0b/AFu82dK7XOuHfByEfMVk9W0/oDviUWfm5Bp9+SyZSlXL
/u7n5zq5Z+DDOT+nIAUku3iamDLNJiL8anWnGyXpDr+10y2Iy9yc3EqyiAYWpsva
H+7pxTuuZQS3WlhF1Vi8sHc8V02ow32Y0WX3YLrGKP95i6GrUwHKgYRH2hdRy25n
U0lR0UmB4H+QznFnBzToUBwGtGHOp7ITHgtZ+0iIiOk37Nxch//02Iy+t2LoUrKm
XpHTTVoAVfMZCER22QtFghdWHIuwjBG8OjSJvzvX383NP0H601n5yo8IyKe7Rlc4
gFpb7sFwIu2JFuH5J9rk5PJRbq3et6eXps11CA+wDpdE9f+0Sn4s7sNzagZ23N62
owtjr12BrvXMc/RWD7LMDKemH1Tors1gpMJTpaS9gegsvmzT+NDXnZmJQnSsWvPw
V7bABm+A6LhyK8gymB63AMdtKup0kWOFO8AclusXlagJxJZ9Eq33ktgNVvnMI7gz
fTPS88oxKW6ZZrJ1jQKDx1udeYY1MGnjv9XmqtdMF17n+gsBelBQctDTJEemVCQ+
cb4zeAsv81Zlw8a0cMBuzU6xp8CTL5uUaML1E7ITUe33znT4QS7emXKLRGDuIliY
8b7yd3shJJ8Q/lq+TumrwVZ1phBNtWen6pGlv4k9meAgxCs2jAdB8M1JU8ERDsuj
I76/Aw3ek8+KDALx5fhRMblgdABNjW7NjLxVhSpNhvOokWVUwCXmJiCIbIP0h+Ma
D6A05EJXnka4MXvteDtAYpwLw13VoJ6gpPJwFedr9HvWYHKLFLxgciSCMyIdZxkW
YmIntN9+zzV1/3fJ0XZC0QdaM0Dz1KwATwB9dKMaeIXZW/h3Hx5JvdAgPOptsqjn
2FTLO6tzdMoQ6xvUPcnJTFXloSe55WzXxzh0G16kapIYjuiyVSr2qnuM1FmtBQ/a
MU4kOtsVBBnb6y6JWEwCK9TNZl2CfMQ/pBvgu1eIkc7kMQ4/H1Mj5uhLNrVFjhLy
WeK0MqqKOxX/OZ10xBYF/RpRVnZFLVPuCO8eZLpO160s3uEkT9LA6W8VXJ7rSvXV
4OHl1c+DSKeXgVvRfv93/d1/wz8iWc0IO/yMp568Cj+0KaqiMgINdmvUDvaZiu5d
TmgLjKWSehcK2HLeRHeKjkU3MKgjoI7UeJ35qgE7Hc5JJ3KEI7tzbPX+xpkZ+7b2
wD/tFfjBaMVo6DQwOvjXZymyZZI6Ia6Qzm8xbnnTTGyrLCa7VBjX3cdTA30/9WO6
cqQxan179NL66JGsCBH5Ttdo2DYCJbkj+e2OOvb92h1kz99majchgNXtDJWZjMtK
4+ci10SPiHAXcD/60Qx87lmnr3AsJE39Tl5D3BgTXPNJq1tk622esMywJQ6m44YS
FQvxbI41U/WYmMz4GM3tyLmh2I0Z1UgF61HzcizgT0s+kogCBTKy9edgNhYvu9DL
xknJ5fyrL4D6T0tHmZIjQUK65tPUeRgfLV6/QEFA2x8XYLz0TghALfCmKhcEYrn+
RQwXd2kqoApgd5m2Mbf7PdCWAnR71tQn4xRW/v0w1E7tAcam2d4CKL0SL37CJflH
L+ei9js/uQ4YCLZCD6Qf+WPqtELbu9gTP+Ki++WugB1UK/5lbUZfyiCaf305Xy2s
RsJAs2qsEatTf/8L4MyGdOJYvaw5CTjOHnT3vgd1/MODemRd59vuCX4YbJnVCTck
34MhZLdDKnB16xFTfy6Zh4bET2jZSWaAs/ADXcADTmgWO07cOJHVEwKkBQY5Ek0M
BcCRcJKJEJ0IpCkmCNZez+iBI4QjCrLMeD1pNOsqAczCfKeXgt9scgmIEz+SEKGu
UzC80PLWFcGGRMunhuEgyonhhHser9fmUiNJPdf3nqxB5510H4XS6KJUXWTLJcOT
qleBPrAIvgbeaymgp8LS/E65ceA3E5wCUlrCvea/orwxNQ+wfvmo5q4gi+th7w1D
ZBRSRY10J2HaXQpoWe0Y20oJAiiKZpj/WheP650x5T8Epc79RDUjO3519U6XuYok
RMRiWB7Fvw6gG2E+KeNkAk25cIVO9634nr2fMr5oDS6/DvCuCBcEkIyAXEM5QDJf
kquNdPF95gQiDpL1tCKkG0cIsg6qbRXQTvOdsuybPPAQV1RMvkwjyQG5hR1Yb22g
Xm1UIGIUtzN7/hTOehY7MHmrgl44lOs7qP5YjhsTuAw/aa3LKHN92RVVtT3l8FXf
N9pvymH/FxJkcvPF1PPUPv4mTZPn0imeTiFUhgPKf+GqBShWnwdaCps6hq/fJMmm
g8A/or/pO+dDfv3Dl3Txz7Wr3j/DlRTEWmgzV5YVylvPSlZGff6CA8vJpe9kF04Z
kqCPJvimWTzrkdgBTz3F0/91hL0qR1Q3NjEaXVCI0Co/UwvT6Rm3qCt5Scq97Uc1
FpZlIoBhgzzFSstPMMAb+Zo6EHlzLMVwpwAsJFJOjV8x4M6AxzCOBjmSHzoMFVum
gUXRQ7ifgEPNz27HxUpphyjR79TKQEhI36Q1tff8SshnPQGwktD0RvNDh44F8gUu
NUqEgsPEpeqpy69zZqHSgYmdlDtStPmObYxudexin2swhaWBHRXp/AkjTRJ7Cqy9
GUyJ4Ru3VQbWz2HJjPY3Z53oaRv/R6CG0FKqsscvU88bgB9VJXX3o5ft2oSqbZax
e+ML27jsNA35JSwYhhaMFGbtAmEQOpy9E8OJagh//1Nf9ynI1aK4g0JdDzE+GDzc
EdBQCjJAkBElwGUOUMsg+kCoujGE9BryvdAD9P6ZV/QQWYmpMZt143q3T5YF8xb1
ljOqy7vzpp1Eu4f73S/YoqviJT+AZVqzBRT7EvSD/HYyVkFzsxIJpLu6si9t7Tw4
NhJlmuTmTH7yffqMrN2HOgqK2S//00pYOrmE2INnpdURpzc8bZJbneSNOfw1qag2
ewBa6ikwmJ+oxNcull7aPgehEAHOeHU8gsjJLjgmwTpgpetd8Lo2R/vs+5S3PM0t
u5sr4vT4FTZbKtNsB7FcCFuU+h07en6nDpt0tmHnfDtXmA+lICcKVYxs+B+zS+0k
e5BiaPQkCWRvNHaCTRqFeCAicL9SER2DntHmMkBiM6exZFVWrEZL9wyPb7K3GAGv
Odw/2mhyesLprT4vmqqkWAeVRxiCkK1yZKNUpxUIOpmKfRlgcPTn+hVgKGvN01o/
sJXEMj2TTxNbdsGu2mg3ju7tDJ8xIsdhYbC7TMYrr5m5fqXFgp0rP6KdOPRFVteN
WvTRMFa/hw1CjNfdC+SdIiz0eO71ZDbFD5oWmVbZJ/SoBPZBg7fW7jD4iyV8PWaB
FfibDL2g/9nGLjl2aEDt9UnDJZ7nkmbuL4LxLQV19HTmdmlkFiT+CmQq9b4nAnZb
Aq/aVMgDE56M18SK6HJsz4WbqC0a5YyFoOUSNDMNjHpz6qLSmTHo/KQj6Z8SpFOG
evB+DZdoWwCc2MVHWd/yyVi22baFB/omiMUASAv+BZm6x8VRX8ViL+HvQqNuT1Pl
7it4N1v7UZZEq5FK+rdYYxofiyf4m6vUQmVYi9YoK1yH2PHGlnXq7cFcNzmTR9Hc
YTm+dxqCQLulf6Rh846//erCGdTY/zIlO/QuhH+gRKzpjATchXMrPa+7BGUDuQGk
1J3B+kF1+EyOofkFjIHazWWo51vVSPTXTNr67W6kLIfgvWAe/UhJJGb9SmGbUNXs
q9ZaJcHjoiYQkyKvDRSADvJUdEpCtpT5YgurnIAK0KHuvkQVoDx10YZXAe/EMocA
osxVx5YYaJQzfXB75HuHDlPm6x5Q7s+f94T3UCNhq1Cik0b8JdnzJVm+uFqeZXZr
CVJz/GN9mjU8CVT7XKpgerepfv6BXFihRP2HreRgLvD6PULZlWnLUyN1/SzcwgfV
2cqUo0hYLEpF7zfeJ9tMeMeqvJh5Oxe8ijBOhSQGUs+0YvP3wVfH6rYAmptDdBxv
g8J7VQRKvGihq+g1jyRa3F3MmAEOUjtsgdXElF7TBl4L4Y3PW/Otf8sFazU3oMZ0
/TTCzb35gn24WYvmF1G2PAfHAUH0Zl2wa3+rETxLnmNdhPlS1bJZ+eBrnS0h/H9Z
Q9k5LGr2FkK//nbcm0+xPDQfKv5PfEGTd+Ex0SYFyGzOxCyxc/fX1yyc7oBhk9Uf
r8M3mxdx3NyhvAmI98aStmKUzp/95frmWAGz4dgetA7snVbcXEUHbJE0fGEEgyBI
xrQZSmsEAjHdBWS/HsgkABwKeOb9F2VzwtdXKVcaZx8s7Epcqfo7u6+SYwTM2IBj
oWqeE96Po+65ghkSyM0cKWZehdlo4SrXH2zkk0F3sXtYPCxUmiEG0T7W/qnywoJb
c9vp9r4yrk6BnoIT4TdDtgVM5qYYUGApXGhtJPrKtlAn6hXDdpj3pxEO3SdPmh8F
b6eaq2Xe+qAk/HydtjlWdprqChfhnHa5e6K7MqoPZPl6sRtl1r3yaor65rLvNGWx
YZuq1qUrxxh3MQXYvujXGsK3+/XfyMyZxaacb0wCnaQvsvXwCuOeawIInWpickul
BONXOoDMzzlg3n+lEDG9ImxpLGz0QVyLUPP+ITW+tzDril72ueKzn3bGPMU4AH3u
jqQCPdez7+r3JbJg2z0/6UgYglImOH1emjqhor0+m6PYfavdbv6QQY1WGjkr+30v
+zNfmfpqlsCJNDkFMiW6AcaRDFuexrKwL+dYpIYd/j+LqeTeElj2qj5WGSI0bNrr
tDIPrg7Vo4fVTktsZZNgxRVZjAjO13K7orTE1PeJ/5PQUeJF9EoSIpZ5KZDeeo5Y
aSPWa8K2RHVtQUhvHwPO8A+lAFkUodt5x2fQUrMxg8TyH3fUMTCNQfpnkD/3yt1T
gHVA+pB69M4u6KaWhBLyaAFjDujqCnhmdvDlMgNqoGGp5O4s1sFvJr36DwwrC9/t
7FdSYzlZjG5PJSZBYn145GtHw+UaRdiF/bGUUPKii/PxnmDLaTsjVNkFJegFG5pG
fnd/upDIv/V2Zeo81eUstTKUGEL9Gs/lZHhv0CrCO/rl54AETMYzbNELIqabbrQZ
wv9LJGsQtRCpOqcFcvlJlHvFwV2oDTBFex804GYQUjvct7twDJ5vjIyOIox/nbQ5
ZzewEH7tlZY0DuzFSyS6oaQJQPza01wwT0h4VUFVDllpOyqEwknDXdEu55HEpKHs
1eUN/uGYW9wC9NCRumCXIt/g2b8/09q0mGrWQ7IuuQOtuMhwEAFwkudPFvUC/nhU
pNqm7ldGVf5KulvTpdhnelwjMlwrcdgNwZFOIg+z2BS7PdkbjQI3n3tjYRtcViLX
w/mGDfGf1mAzY/On32mXFumWpNF/omJWTOJl4da+QlYOyfuDy/GJoYghMN1uI75v
VvjekyZdtaMjWQyHC+Oe1QXL3mKPVWOTWiRA/Ha8kPONoUr++Nma42Njo38b7LJK
iDvW8vZLuYTceqCcRr4TjQmz85sIsZqopCreWH5UokMESVTDaXtFOQfyFGOkYZli
NPu+wUKwcwnmdw07R0/UWhf6WAO0MYBJLFTIGlX57IYTRTGXig9m781qkyQNTW7+
RLtiTmu9rxdfl7ikWQ99WCxjT2OUhQ87FpfYfhp8sBXVo9vYvJ1LFEh1wutMZA2H
VUUoa3Qsq0k0i7dyIj5ls3xUBpMh/S9jk5Gc2EF45YN8WLY2m7IoEARFsTyIKExT
jhYYdG2WNPIQ9bODpwWgDIM2TasABnuXeFnGAx3gP4JSjE+m5PtD32dzPWoEQRLz
5eApysXITikv9/uS1HQefvBFVTPQMyhEGI+8Pb6uKJ8AeDccvJwfoGjJsA1fsF+P
7RJ1fNeyOVAmzz/+dSpJbzI/V8p5WAOlnC74y9Ut1G+ovbzHC4xtVzcbP3jQYpJj
qA48b7wAPSCcmK3xfIq2hA0ZhDCq7Xa0/9RMx3VqNPtjSDkfDTowdNviZFVnMa/d
sZs/5gHtyn2znKi5BmN8B100NiigU7xJbjF64kcouz94WDgs2VNyLraTeSC6ier+
XSlvHzJDxX/qolNkZSDcbfYVfCwWC+ZCbbDQx0Mi8uN7S4XmkD/lrG2Sq4L9PkPE
gYUtssDke3aZ36DSsAsoJH5UVWJqSaafCoLP+0rgT4rnqazFwndtEnwUMd/IWRZU
k395taAni+UohJoXqPkOOEXNvgPjOFSyJrAfyeacCZ18VlUNyIZ7/81dbLLMTAD7
pMPf7HOEyTuBlCEWm5xLbLxG3ehuVMRqCuqmi2Tkv+fFIAh/QE+z9FzeWXM4l31g
DQBO1yieJayGubJIIiV87S+THC5RbJ8vCRZlnTLKaFZA3UvutmthpLc+2tMzIXey
Ai6O0+NmYF6PqkfXtMsntf+HtmN23iLVk82T/CCmkNIQ6XNqDme2yZ9Kbc2No1r/
qIkBGHuV8M7XcmlctpiFucmwVQQF+Nsgfnly9YSX3BgLr3VSO4SW2d2e8OOowiIa
l7uvY0ROWoIS+XtAqaOUJHXrZ1nQsIZzjWDsHp25BK2IHREtPfAE74yaJsP12VjI
JEyoI3eMflhW6eOlKa1M/5BmuUiudd/MrF4gKEgOZ12wqo9vXeu6MzhtIy9Lqwhn
kRyWY3eYVdeqoWnCLePX2mz+wI3ed6SgUt/HxCvvMlJ5cO5vB1sLQ9ZHKQ/ybZ9L
9O11Vf3z7c8A78vMYEpiZY0t10uZiXhO/RPZ58AXzpkWxNVyw3YkOgmRkzio4gzt
Q44sHonhT/y4QmGQMqJal2CH988TKGwsaSKM72jtoiVOIpr+mAYS0+gUt2ftUSNz
Cu7VR3+B8bJo1rZ8Iai6RG7gT7Wz8xS9xgv4Do2S9oFeA7gowCb0cDWX6wCd23d8
VBs9IyUgMzw4rxFZK6WHlfH/X2CvpvpF+H5r+L9kCSoiCCNP6BTxO2B8iRFLBXng
vqYXFQn4vhzHBUYIwkmmQbJyf+WBr/7bIHZKcsEZ0CMxaQgSzZNtcbQ8TAXaYqpz
mugRJ1qQJutqxq9yno6MfYJzERcfYovAhdqkF+K5AOc+qkGaqkwws557vPbiYroJ
Ct7b3rd3uY986ilWuF1RxV/SP3UWN/uKhTaZR+IjD5MzJad3YvSutoiL3tn0+nrI
r9BA/SB8lnzuheKCJYuO8kBAnfUNRkfH3sF1Fa/c2lXdjif9h0tmyrgDm67Bp9UQ
dhJ7GvIV2iiVDf/zNlAbDVjnBHPnaAf5KS+Fez7Ixlwvpz2RjTOmk5mv+TqMzmnq
3CWt+u/gMQPVhffstf3NlfBdYwAnzGluB9Dfde/92rAgDpK9rWWbUk++RJid2bvj
j1ntJkFnNvI1MRwP0Z1bTZLcZarccTbAUdSNDDvom5OFqV5w4PErGuMe3SVoaOE2
235Td43TSL14ZVkskHzXqgpcSm9Ps9dpKx33/c0w8Df7Ho5MlpPXTL8+LVybsIwk
XXGTIdW17GokWk93ocBfoCFDUAw2sA2FEAOoQeYau0vreFlR/kVkLFSEySjg/WVJ
MZ65lUGfWcch4H2vihVUBrYVvBoDA+IpOh81XH/3f/nmUC2e7IxVOT0elC+fUcs9
G1CjxrmRDNbDFhcArLUMKeEaiSBZQ3+a6rBBB3dEouLmU1dH2gTbkwUB6scNo/1s
gj+mdonFrmABbWTzXKyAR/7cCy4uothgZMmGsQ7ThUB0nBpaeSc6DqMRGT3rTLkx
lBmcmrerkUceTa9Zj4Yq01x2RJu/cnw1+iHeWDcbWkcwo/VXYnt1MSecyV/h45Kv
DNgvVjpZ4LlQZn38eUZZpCKHYLZJTF8P552NXdRuqigHQTOFf6LKPlLqXQQWo/ls
UuQB6PrfhyS5cpYMK2Z8inn2qIZJgi/vc35MRhnkRSEB9TSAP29vPbhEhys0gscf
DP5oHD2uXBQgYb1hZBgYht/wdxHQg+AaTQbWpbE+D7Y7KBy4MMfaime1Y0AuPEIR
HorW+2A7/06i3K2KVI/RWe2OChkYjIJg0Ge/E/Q2YvHXi/Tzc+UZEBdIUWLB/krL
MNXs2xqI1hL2NSQ0bye/etaG7dEbuqj0PgALi7l2cbIH1R8S9kIlRYS8NA5HPFkL
/0415FjXcVIjt4T2pdFXub0c2kSL1k4FLi7BsgaG3klCE5cfLlrsbED4+gmZAw5W
avyoniWzU8OR/d5sUKuHJQ4nbf8+zR4uCILzYlfQECh5396ey3mR5gPKw9tT92+p
lHfhfDV257te1eaJzl7uKWMWSdTJOJY6XkYY3kxdXQ7DTBjRBDYHOUMoXijKh6Gq
s6lp68zseuOHKWfIomDoLzyvAojrwrogoRlUC8osId1gQD7hQ2F56aTMsmCJ0DWM
1iBPztAB9pCur6lESd+EYJIib0dJekwTU1EHSIXVqKWcynj+ufgIoZUvtNsrP5vj
5G/UVLN+AojY74kjNXjpXD+rBO1ATuUSHgOOKHMj9ZltqOKYkzpyvJhho7xylkxb
7kZGCyR3QFwYFkAmVQDEpSKiTPh/rSDDEbNMG4NDJ2vlt2DadtDk+wIaDbrs2Gp5
dYbkmTxTH0h5qq1ZyDLOSRgaFiU0hBOpCTbE9bmbA5Ks0fwxEYEUXp8TvG+1aEwe
psxZ3Y/0P+SZ4mRdBXMuXp9i6sIdVII86AzW05xnZJuJUAQgI9jCYVqPQKslwywn
ylTCk29hLR0Mn2tEX+18CMORrczSukxjsgGzv6ofXLVvxShxouMIsAyTxPOoNTJv
su1yk6HQhKrzwz6tEfhVIjcnlG9ooIx8gCXXCR5FEmJPv7BTCdlQddvCg8Si70IE
9LAZYDHjU40+9dMMjmJMkvYau220e+E+aDpzE4qoU1Ur4cihPv3o6JhOaylFuRrT
NN8Ef6KG/KIoXH9TU9zVRpISXX+OsfBfU18jI6URTIUzgM2vDlY3+vet4u/Ozqdm
Eob+x9Ubh1baxUmfmzJ8bBw6zAHleKf/CS96iwTJd95pEDkMa633Z1sEzSGzTiYa
VqjcWmp9WWpZxmF9PekUy1ufEwuJXnSIQXXon0FUPfWwb7QpZIf3WpssCImixFHm
xlYq5R9+Rww3BrdaEXMp/fpuQMMzd3E8mrjxTn3bRtYi2vY+o5nZnJ8ltJtbwTWc
v6etZZnNt7cdBe4sRHU+qq7rM9JaBFi7Bxixafr7G5Sf0xiZ3RWg8G8BcK/0mQpe
aksSRuOmiT4roUb5QSwGjb1AHSndUJ9P775/N2poGpTDcPNskzARIfbl8sz860K8
dbudKEHqDxr/vkTzKV+tRltfxKZFDSGpTqPEwYmtUWZh84xzNwuQBzBhNF+tze7e
si4hHDMulMC75TovqcWoICBgjiwrnG5JT4gvAgbYg9hHujqSVbBuqLktquXIL7lq
Xqp8Dcut96QZ53aMnsrRjIesNcHRSLSmZyrRtai8J/d/LdxFWPxUpF73aYUPC5xV
DcBpOf+iGYG40rmfmkKYyJxjlVguBOHFSEXg6GUtAVkY8ph+kdGv2fozQ8vnDIym
r+eFvXW44lSV9Om+/v1jy9p/ulkywXwUKEzsFr948msjP32gkJw5Vef/MH0dBXXe
nHxbT6QJfGg6so3bAcCwfDWf+k8/IxBGHbFuJo31foh5K+sMqhSZF6qwz1L04tkF
satzo/oFAdkrXlfsIRjRa8SEd2Ml9X9lbStHnYtRWgiikQ/bWbT3FCMBEqc6OlYj
t7XCTWMtJOQh1/IyuAcWetzDexmO+Ju2GgZh1/yxixA66exa0lLD3n+aW8g28UYQ
e119XJsIjhaJ/MHl7gOwdmeJOA04kmbVx6Kbww+ux6LPK7HkGu0aInVYlzAfX35A
DDAGl0bvadgWhPfVdWoQLOu7WVM99NathrGCtNVWTmbWW0gU3AUsRD9g/DtOfCNj
DBqq0YUVEugP42VhWOPs9bPbq3heJcJterhxGbJlbi/bCRF1o9d7ZIjaIM6m00WY
UgsrWfrFnO1yK0hkElo7ZbULQF/3BHTOE2WI15h79woQtkYpTLVDIrIr5e3ORgtZ
rHmXdTVgTxOUVcGNuSDMXSpn4RrtyFdjt8gl/DdPSe1S7Ja/i2k9ahO8KKWohqrv
UdvpKilIhuLPRHv/HZnwArhv5FqxzR24zkjzLGWnyV65EBdClLrKJLGShFv93ZSR
UYatHD8bn9uY8gH8CSvtV1qLo4a5vKqeWlDu5HWnP6YjNViuIfjP2JJvqYiUrOZL
wc0KitIGjB1/2sIoIjbL4cbT/VvW0rP5J/QT0BSmenenwdHdHEDK2WO522CrgBG0
+Vyai/UsuexBftIqa6WP5Ut/IhT1GFyPqyKMQws2beVzB+5EqdtPpV7y3uWUWTLy
NZskrf+dCcoT5p940w8Bj1q65g1d23HxZl/u+MyFmmQklpQvGT5hSf2zg74F8GJ6
SrxJrtX1757dr9zM7hVk2IAW75kKoh1m21LriRJzVvgsvVO40v4JR8ZjREHAjKBr
tQY0OC1X1lQvIi1JvjZhroNwjOajXuZuuFN32iL2p8pqOu9ruOIeCiCFSxpw0yzj
wCqDWj7D0oYPauh3+sbqXsrtd/AQsoMahca4NYLV/dPX7D4N49CpEeWhigvSmueC
p+r/mqL5z5vYfnSH4Jg5PGNTcULoIYeOglsC3CVaRh5PzgRoFC1dDOl32/jN7Fd2
j9sIWhSCNVghqBKTQFhOO0k9ZRTkr1gwo4PffGiQYT4FeE4+grefaEf+EbkTwAFK
e8CzvKbja0Mojio3GNpTJxZ/a/EYAH7iu11sTKuEH+3OtXytVI2kQoVx5OBKL4RG
+PWl5cKTykuFf8p8bxbi/iiiyhxlUboQYzcYtwbWr+nWBvbCkewfamZAo30J+iuC
gqc29vkcT11VOvsBC/9EbCpfS9aKlxprcLg9ScTjongR7YTUAM2STj/+WHrqqaeN
DDIuBPD5NS9BI7akpETEmw16b++LcqxflaBAJAzYBMIshgZaI/jnwhTRZKhaOXZi
o9CejtEYkwnD3G48G4f9aqU7c5AeJ9epBad/6xIDIH+OVwjtUYnYHWaHtCVNcmYt
Uc6KM7BH60s+je8R5FiclHdfaxBAmOBvfJ/jP/T/zqV5gJp4BrpiZ1wYqqmnhJae
Kbyv1KHNLKh83Pruza/cvY2OBsuhytegNIrHkZTQjWs/AZB6w2x4AKoujwCyHSW3
9BYEYEssWcYWNz7wGnQ/i5hHIZrIDfiwYdDUPJhLWp8sNl6bTcsZj/OD4PErB1o2
sEw67wbzqeZ8ra6T9W6isY0WBY7A+tsNWEoPQs5crF6yIcQwJISl13/B40qGANPD
Nd42U6y8q2GlQPp/0F3SPPTiuLqhm/23PVnpkeYsqwUYrK1Fz8FwQoTlx57e2nOQ
YkbinQmf1SCIK/h35pnhtRYdifDgWLsra+heG/RV3r2UY4OWUYR/uSsJISgvst0e
aKyU4sLdixyK1n5kMV0mmW1aGZWk4KVIuR+uipZ+OJeeo75KUK32pFy+96Dcjbs2
bnS18xPTewm32iUbZd8aRMi8wkVx5Gil2uiKlHFMnbs43+5MJiZeaj/+eFLPkOYT
NLgnDAp04nNYv1IcnP5KLp3ELFIQN++KhnjHnhzHJmWndZO8zYNBo53+bq/c8Odu
P86d4Mo14NHGB7kCqLFum/ETdq789+t9XhKulE8mOpxRdwo8EBcANDBCzcsGIIAB
hJGlKCn7nKD+6qMCJ6kk5i9/rRKIiAoxpIHE1ckg1M9wlLrYC15MANz/u4k1ocY2
bMlyN0NvWWIPcd8FNouIqx1IYf56fj71zJwlMIZgYUN4YuqHYbVYVrpmGN45OwLf
raQiVAfyk1MGqeC+kACW4/0MVNR2BJXqHoHXeV59VOP5sld/wOOXJKwtnupOBNCB
BO49TKqi7RHp0LiOhvO0N7OdqPFG2GffahJmzApY315Mhg1I7ltm/0mdwmHm2QUU
uf0AKZ5N4MnopEuT36fCj8tu25oUL2pW2zOcBFgOi3891y3H/Ko/rXcaGSFK01Bg
Fcz7DHeYOTkVCa0yioJLxHUnFg9pauhV53TXc9saT1qM22CC+SX/xuiB9Etx0DrC
LTLtqaHlSSHRN1lJFrSGcxs3L+dFwrWpPaAYWnpXZE0DpwKt1Q3LSdYsGrYkzJEF
Yc6q2YKdAVlBgIOGclshqLeaNCMVcz1cmRjcqYIpzDgumT7L4bvWFAT978hU4IdH
0iOg4cqxYk07m+5EfiEaj8eOlCOfkXbU8Rer498JQDw4U5oEAkE5/XmlLsTjZO5w
2K+fe/Jn2i9cqMrdaOc0Dpcf4OjsLTIjJkVqJaD5TTIC3aELfsbL7k3jWA/AwYTn
v9W+Pu7T6+jEdlbZcftBkbBHgUyz6WgBFFAdHXExj1iFilXIyYTH/AhbMbSlBwwE
aiNruXRI3MciAgKDeK505z4IMGLtvr+97tsNZRFE1afmkKJDSh6qo6ttiyB1vClM
lvRHhii91BttIIGpcd73sgNMb50A408uw7Wt6U6H17JB3lfGxx2Px42+kzPSWPCU
eN+dbPsinPTPzmMWBhN95dwWq9uVrXVyx4y6TmaaAepwNVpdCcn7LBtn0uwhuNpJ
k2JJ9Xcf15KGxZzXAGXO1TWH5cjAVeaF0HVO2y3n9PESKHC0m2W8ud9MnVuY+jPL
SEEvAzdoIRzLrnO2vGJp/vsNwKZPNB/88qRb1+3qWx5VIuJVTmz/PHcjIkTJoqJZ
NAjKUxUK1G/GE3FpCg7N3UeicIyAqLzCI3TgjZBpOWYOzwe3BPEm3E8loSwlSOOB
3GQXAGMFvw03mcvinYS3BNMzGKhHkSSCc9MnPyNxjt9WHwbtLNqNOvdt2+m1osvC
PJRN47iEmFKM41CAxFe81Pimtx0VRGld0Z935rmMAbVA1zRix36HrFPCpxeURIxh
oqjnDFKVDs6EEAeXg4sZk8+B1d0koiqxUpKSzSLVxmeTYR2cJoFplklBiUl8UiuZ
sHcEHHJoU1gOlq2FAiIMs4mfDftaCWRGMvqz1JPjZafbx0W47TK0OJ+RlUlKUVpr
TbYbOGdHCxDbkJNZuwZBmB+CVbquYpZ41Q9ln61jT0g+o+PQeY6AZb5/0aZsXILX
gcN2KORabfuDg1L88gP16eekXBdfpLk44Xf6FD1cOm7Nd28LuRNOxhZq3FVhdYUC
kd9Xx+lNFoFA/d8Eeh5Mw8IXzv0zesqwA+mf5mG3tpAo691T4JPyjgtGAlzx8Ej6
eedkKoliLFvFVAzTE7Eot3EurDmgusnd/caUYk6+BewU2cqVE1gLg4CxmBS+rg4Z
QKB0AE/GmgNfUfxuPSZcy4LCjdnYLUOcBlD9jhFrr3noGsWKUdV+X2/RCaywoKOY
hLCXgFNfqV4bKYur3k5WAFV483KNzxR0k5ft6AE4efFHlzPIjd7edePTD2KwE+T0
LiUey7zGlRWrrtfJWiimU5fgAyt1dG7X7whrLOtefzivEhzmflXFHZ8I+9tzjtso
4NBy7topsCCjD7TWFt68RSsMCUxeWaU7cf/4xXWdPN4axF8gBDapbIPQ4wu2kcRZ
xZfbq/GDSkHqQM0KbUb0oUGaOtClvQNq+Xd+V5V4Q7trH7hImO9NA1LlSUbPSN4B
p9t+vLhWKaQd6bmkGxEmGKMcIeHhfDAksXn27XIHYQjMzOJ3kKCzT+LDxPdSVz41
wcqfuJofJPuMoJatDp2OItSqjFDIjh4COz7UV3sr25ef6qksg9JaxsYe/rMnV5LB
rg9xt5Ed+U7tafH07r0U37WupqqCbiehEEIUwBji94/u4TN8Qa3/ZXC4tksh3yf6
iAQnGBukiyFR7qjhi8xIOKisX32FvX6Hy649Gg3RnKpd1LtPV4IjtJeCxhcKG/hD
VgfV9/aE76po2OXVC7/t1zzp+ruTlft3u+FGvnvWDb5j0eiGyo77lU/dLG+UoHEN
Lub+37kPEQ5yBKHGgJGU6OYdCh7KGTLJdTVAU0SKL9cQ1XAfCYarpd+/iv8zrFwz
t1KvJz/YWDIS/IqNstkEZBfVy8DtVpJABgutIH8zDTGQ67yJ9TbzCyMcAPJi0eJO
plPGj9Ou4HRs8evFS1OR+IQwAZU6WlkUcKgge/LM4BJ0gEZrUmafVBxC86BFuE6l
mPqvHj4j+bU9SZ1GmXJjalgOJD1OUIGmQg5SM8PvJE/MWD0ic2iL4cShxMslXs73
ejMtKeO9e/HlILMYMVQjXnhp6liimnNfI1JZQrQKM9O7rGi8aDfpEff6dalboG2N
wYduWqtVSBXBjneT4akt2wUPP9y4YI7315acrh165dJ1Ery3+v0wFHyelAysL2Ku
teJkzmQXHMdF8HlniJ10udNwtrDQFdncuqHOl9+5WYZ+44I5LemyaEXHchjm8x89
Cb3s9VA83DKAVl6AsxH3vXUrhqx2KBftGhCb6i4ROMaQTdH62e/BBkMTzqKrNhNe
mtWsK5m6nyhXYrN6D3Z4HUBs+AaW8f3TQk1hIKmbNlQIVvr1+cbJBK06BQ3V5JRr
5hUqhYWW+EeJ0QNseYqR+zrPpvxKrNyK3+psh+hNDDN4P9TPzEdKx5QxlUF1X3zu
TBFKPhTZ0RkPVsVp+WlAMmtsDTaw+7AbmHExQ5wpQoQHU8DuF7eYKiCepTcTONMl
za4m+G5shKL1mbC9eiH9XcdRfbbH+tYdIW6l+KzKYbt77wE6DVJOrB7PBZ7M0BWw
HDsAXwHyLJT74U9fPsTQYWqWLk6YTm2SVkg2dDmp3p+e4kSLJ8A6xBnqN1BsDq4p
gc08NpvS2RHLPWGLRuq1TNBt/fL+BhOH2MFSoRfj5ymLSRgT/PxskHgDVnHcVGBn
sU6yjDuvk28tQ4pFyLOpeGugd5nWnIb1q2dIwjutkfLIvlUhOH1HAa9E/4fE+g7+
RuS6L7OoZA1ELkE5pEBMgqYJWWyT8G9ARRKc6t/wegVg6wweNxJrwRpfkXu2V654
uU/1Do6sFs9RGqcowauWso6p3C9jUsKDX04KL+496YOMB0cmjy392cU62pHPH+sP
9qEBGS/p3+HxjLbGdR6i1/LkBEw0bhhWuYYpl2Qov/lHKFNJyqrxbwpptNkc6g5O
XNguJyNb9c2JK9CT42tooR6adzbOq7Squ0ObOxdg9I/DwJK2pwTsnFay/+y2kTWp
E6QdB4aDXHDUfkZpArMdg2STIJKeyL0V57yHwIXDhcPtagMEcUWjkdnNdZnzi8lB
md7XIbzRR9NQ9E1lNnvTxoGui972HD4OFvTT7/Gd7yry4feeimgvI55XuGi1EOPK
CWyDbhH7Y6qHCqRdVWPvaX4NIG7CntxEpSYKiDZHhppIROSt6iEVBRnkT6PRd6Sx
Pk2ucmH4DHElmcpnPIcFL8fLnV6oMJhezygLlmzHsRW1RFXp5ncKKrkgzRwWLplW
L0hCICBzseLx2bYOgNKt73Jd7N/yMkmrdXzj2jiH1Bu5G0+m78zXtxwKVbnAGF6+
tkACCRUTOylKpRNjnRb3JTearpoYGREnJjQzzvo2JBAVvNutA8JReZV8mpOMf/YB
PCqDUErQxbtO4uWOGUPDXv+/5a/+/EOxtSP0fCmC7tAnDrlYNTN7/RwUR2Qh4hk9
rKEIwaJUT9hLf+NjjY/7u4pcAOQmFm7lwESYL3PNqlJvbqhDTXYZr6hyOIJBKOco
JXTunz3ATCoPW7YNMnN0DELiNXk+8Pv4QWssJ8US74BDdJiYJ2J5exBvziF9bapP
5LJfeUw+F5Z+yVYOf+/We/AHxDXbwRysWP06gd/eXGry99doPk1rJWiSBNuMpWVx
MX3UmPUIorVLFKTBjWWHOktxDtV4G7k8z/Z+luZRxRBUBS4STLrSyAv8X4KEiOaG
pF0c1kS6AnxMEUniHT6xfj1QIbW/qlenAVMAh9wMYTZYPKv14hmeQgA3Q26DYfQp
FRFNqxhrqlIGWnLW/PX+WTCmGzAS9sKfCVKawsvUyLCoEF56z4u/A/z00SFtfeE/
3lRXXje5N0XTlGslElnXNNzMGkikwPLhphCRTgHsE0mCmM5o9sAyL1UnnGNjUcG7
8HAzbbL1aJVzts4s2JEYLCTuJSDPxxP54MdfjRQBZhbbWIwT7Gd3ksRgO06Io13X
fX8mhVVXYZeRXt4sIRoDEeonMoEnJXGOwWzNCrIWado7I0ylbiubdpkKk1EHGVnM
8rWMwrLOtJgmtbQomQxOsZQbOi1cE34sIpOHejBpKwaNaiB5dl7QaIMURoMZFgOi
gS69Xh1u7K2IJX1IRHF7zYbLqk+JIV5n5/Bl1Z624r9Pl0DT0qKc1rgRsVOO1oRs
d59zTXsDfdRCbx+WzeX8UkDF6nZaCZfviDGMql/J4aTCmC9Cy3us1XJJ7h044eUG
P/LfmLwSugxulqxVu0IWprouss+pcNtex1QpVAoEO57RgosLWk1P2C0/kebGvJ1j
D3ht44fe0dKeRZpxYDXIXfTK/gls9Ko46GknzupWS9ehshq8n1QJtz0TTC1mcpSB
8BiphLDBdUqAMDxEe2590R8pwzb5kucqy6ag2MAipdggk2ZsObsug2XyG99FNq+R
WMpIVe7r6XxM5QVfcF4yu2Mtq6SGU++eNMf52M5Qem6lPGc2ZK+f29phweo1cRYM
/fMunEe5NZmJ+RL4UTi/Q4tWri5BlypXMXJDnK601f7HvgTV2mUDCkS4Mnp5rslh
TeKvlnDBb7wvwFLg2kZHnNnuaALp4Q9ptOGOGijeZC9qQkhvPyHvXXcv8GA/drGF
8q9ds16YuA8TLRi6CxOwfLLefDvaVTxFGJXd2KVQt1Seqf6TsHfS4siXaOnCIWu5
0gOwBDeGO1lgzdwQbMo1ljmRB++oPKepGlNBIW3U4CSWVjKX2zgPOJlpW+nh9Mt9
DqFOTgbKrjJEpjm70OoABCqhyc2J2JiV+FV0P6RZoWHVDsyBRyb3FLzCGI5d8G3Y
0sxutQXeP46Mom7LagP1rqusyS6oUNVKxj8ID1lGYlhaaZKrKGeyyq+bEDG+OaZe
Ih/YIHVor2NVqNW8+9YpfHnFj0OBa+r8eQhKHYd61/7vMA5cS53Nth+/bpuMQKxL
nVEQhYiMPXXeys0p+VogefXu5ChPbm1zHdWjc13OxLWj6FtvBnkQvnmYwN5hXNtn
RytnnXHMtM9TZGiRHexmZdfQbxnSdCMy/bZW7pX84ZcbJzhP9yQF/+GledK4lDRZ
9lH1LHsVw3kGpXBupDEgtNCamEzb+tS4UpMWLIUUpwFyMUOA9HdTRphVR0jFSYZ0
MdfsVh/McTSxWuVpdXcW9+6m+aKT57rtz2ApisXL0e8JSqknOS/paSQokWJbyh27
s/Xgk3DJHCngJFcPZcPXssTnQBT+DpUcDrHOQArtdvbH2S7yU6wVaWGN0Ad0g8/R
CU2XzOQ/U6bEVl5CtT4XNUCrb38HJxFlyNOnXMhCqa4ZzYm72EvXO1/tMw3SQl4N
YuZASsaBUXgLAgX0pL54XEl4PdBNUkhd4WwWrgQuB0R7SAMZvML7KXtFcWDJabeF
Udxn3FMRZTkJwTHM26JpHtdDD+Vu+2Joq00iV+n0sFe/Azqli0IihGYBOWk1Lx93
mliz2abS0kP0anSVqZTEaegVsF2s47mul/NPLteWmOrHzgoMwOcoC9uDin34YfvJ
bvJgPxbANdRD1Vl31OIs5xrg1+K36wr0zftHvVdqRKOrsdh6DI8w+xbhLINAPAhv
Z7IIMX8mOr2cZZ9CCQNhmgymFEZSeLw1xoAVsRT55TTh65nHWKoXRRSLx+XLibJy
ejD8k14QytKN/dRzx9sSCsnBrNzuoP95lqwfr10hz0OOHTO6Kh1qDXmmILEfHk2L
AwZisGei9ylkgAiOdVzm2FSINy6ZH6zfnlLXCkoRaig/GTYjT9iXTc0roIFjghyt
8Zu+OixZWl6vA6VrVE/bs7Las7q9VhBmRkwxD7W5gRkwWf9G4yOtqc2MW1aYf34+
4uIPhb+K5JYeuFO/ggfocYQ5lRTm71uRuvRrK2CEqPmVXdH3u8wdJeGUSJJwWDHA
BafPkETRDeF0BVVxkXYYeAxyNf5o9BfGg41aaEM/BNJq0mA8CKFFOWH73Aw0ohjz
xKLN4VCcj2bfzWwc5jF3cRKePEnb+OyiC75z9HBHWH8Nh1xkb21Dy55/UwccyaCG
ycTUKjkjW880gfjeiF+bdxyWlA/lFurSjK1+Jxps2I8sxSB+kst74lqXxsXKDDce
Cs68YEhkbpbu3zsPitadprr7dytdtgi4AxcjgssCrHq8tma2Ys/7s91CLAABIehh
mr55Q1qtdhwW/coDP1NRB8l9p7Hr7hsXXEcZTNj3YaH9wvlx3qkcH7KWku0Ksy5j
c6fuB18heLer/x86LQ+MVEEO2Se4f+dJzPyBh+T7zQ8Kc8FFXlEwS6cSGaS1pnAZ
mlYIM+Sf2eedhDuTcRzlAMyOKExAqN1CPc9wCAuzj4riBi0lxlvNxgdB/lymmKZi
ur3AFLfO9EtwfGut1yL2/UQ0IgtX39eSyuMVd/ULwrwWbW6O1qwM8of9LA8B226D
V9Qjxv+3Ohp2Ky22P7AxIYCuNoxBNTg6dYMoVmlG6EwHs7HS88+4BMhrY9urQjCj
bsKEz9ZYQVy6WTj20FSL/RuwN8tuLx1OCHhCmf1rCi8w2VI9dF84dbWbQtRPotKM
2B9qKBInUq+Qk7RTKOjpxqnSEQP7q3/zAYhNDqvem7ATYQaTisIE+jwMxT2MO9JF
7EbP2wq25UU6gLRhxJ+KbsVuyIil27VH35v6zd0dGu/eHAdFmI1pRhytQSOm1sk2
GUKZGHzEDQ7i31r82ASYQ1b5YfjTbwmcm1PETqVM7miZlrkpq4oPnW/TSSxHimSF
vFZg+WCBJ1BeE7VBkUVs1YEguMHwWhB0otjvSZqwpkIl7c/1rP4J2XnfLGt4wxbt
xZbwhFHa4ug3mQ1K+g0PelLqt+X3zJs6hd5zTgD8Hj4xfJogS5efI7R8zjUJsngd
d1a5VjXxbpT71YPY7oc4TFu22pVSOabcgaTc7nKcqlVvGyEEjoki5ZqPMrxBjtV2
4FMjLLCbNySzm3I5KT9qOYF7GZe8rAS+QZLjPRCaS+c34cefWZ1a9IUF4xBa/3TX
HhiTXz1J3I43vP5htkd8dvtZt8Uf1y7IB9dwxbqOVNRH5f3t1mbOLb7nsHvg6uau
CnXEOVxkqp5AGl8XwpZBxcXT3K0R/cGOH3Eml1qy9mW4Gu0R9poQKBl6eo34y15o
432/01QLltmocpjwE5USVYYhlbhCRiXtO88jktinMFsWUE61VIIgbqsf7v40oC2K
SUd30tReNu+Cnuacue8Ta/byFSgG8BwwVm2LjImFTO9wBy6YedQI7ky3y/oQJYWt
3ExtVf/mFefnoRqakL/KHMgj7kh2u23zmJ0UiujueeNxauWQkhSc3R95ZuFr8VyC
m7JGlQpDH6OHhUSClXu3v2cf8nJlGnkjP3zT8gfY+2J086pYt4ldpmVBYzinpaO+
HiBPbTUtVnSxfwvq6TqUtFxL8FleQvGmQCAgGNZ1jT1LxleBYbgTXLXADjaYDMJT
kRVqi4gjVgRibEnKYm1wvmH3HdJfvjMAQ6ZXeVAYyvkqgjOv+dsbA94wJyQZ2jdw
Q0FC/M+VGe2KfzYVFnpfajvwvWU4ppOYHE0TR/oTyhinzf/Mw51xgHXwzoty6gNe
R/3wePAVCri9HFziLesv8sn8Q+N/GTpgIyi7ikpXJbxf4euYj4fUk6GYmBc/j2iB
GJsFwLCNdeHLXk2cyxFZy7W07vjd6KzhVwRABhQtbtHyFLZ6YAEq9sM97pQx+VoW
gNRB2LcyZ0zxXVvtBLO9lDCPoLVt2dLZDXYFxSjQtcHjaZ594KJ6q88woUzXrLdc
AU3YutwvzOny/Sa1Gu1EeeNOZoazr4w0wFzgB3LHOgxcDqmVKZuzyB8R9sNAGhZU
nLoil5VHXU9eoZGPto6mEksKW80MJOY1HwwvwYpQoUyD6HirAEKYNWyD/yhsPf3D
Drr1S/xTuktnN3QEoTQqeeMmk/i68Lh+wf0nu5q9mbX7AQSI6yoVpUad9J4YoUbe
j7k7DFDadndUulxpfShj7cxPXbeNx0wIGPLBzvupNEwNP2EHf5PNFdxSyHysibBv
lzMQEpARQFVjS3zZtL3mcBlXs+U2m+YAiVBXFADlIdHHgpg8Opjo7XE88qEY9x2V
b3intKXvHBzw1XYrlsE315QAzbDy7Hm0cPty7D4kNTp7oD6snDeB5IkfyGoUyI9v
fSUbMUJN1vPwFLrSvPjpaUseSY5R6YlhoAC9Fq6pWP7fiw0LyE7cka2754F0xF2P
T888GSP2y/XPmbuLiLQY026w2uvfvAD7GBkRPuTKz7UPGcydMHPfn3jafuPm8O6T
EHerr/JzRUyygDRXkTQMBgOJ7QlY2PLoeehD9G5ebS5vxhQV2vf0eMQyyDfXr6P5
vYqu9HwSxqlpWXpsUnliEBPOsRJ03X9FAFBTCMVoARPkY15/rQugBQY32LIEAvhe
WZ2uma7UngAuWJXvN++r99c/+s0jF+f5tKtqfV1XkNYvRHIhrCdC/CpclPx380vA
Wcid8jDyTId7ddcrGnM6os3q1O7SEjc4SEH6M+HUd+hsdgknUue2bTriEpx7aQYF
8hMEFpWqka7E6SOAOLObgbcBVg54Kus01roaRTBdAmv4TGGwPGL89JvvuooDHwQn
KmUykFti2xKGdgwcqhOY8W06Ytdi8kEGXbO+1vXjV+9dNX92wXQObFdX8HVZlpHK
4Ro0QbPZ4k/wxmsXz1JS7AN0Iy+vfpt8UE9sUGGWYlHFi8Sgz58b9xkKynjpDk8l
W75GVuzDJIQRAeM7wERGK0Onk0lLsw0s1+Pxlh8D0rKY2x2zYipg6DOeJWnFGaPJ
1nTN9/5VH5XlbmkpzfJxlFmL/rkIrPAjl/Bou2ynb8+PpfoAwNSxaep1nJs4rzd4
FHCJFHPE7owlvz2ZHktgWNjmMrOS0IR6xKSOmyOde9x1pCGW80ZkeG/iXZz8iW4D
41HQGVWcnQKaJ2ZwsMvhdpafyGbAtBpmPCOr3cZy2bhMEVCkcf2FHDsuiSblf67Y
rjH5WmgGpXsT0yp7J4uUbbJME11QHzvfxEyCqiaAWM4oPvnFatgRHt3Lx3S5ofJl
7Zob9VNAHGxoyqHZlOptQ9MjTqYMlyBPpaU4Rm6ooeeHyYOuRMIFtTEejM6vk0oj
exoz6OFHCG20zlmsTBgykDSgr6z9YN5JPBgyUzADg2cfA06FvqhVC3B4z+er81B+
Z3gIkIvJVSD3yZEjs/2lYB42bIIvIVMK2KCyigowT3J0YlEsgzrgP6dBTJ38Ldl0
7S8596RMWCaS+Aw0N5/L7Jok5Hha9EoaH59uXZymK5hNjyROavfCtT7P42Vx7eBy
t01kaS1tyiU5AW70mvxSFuZ2fmfaI8IoqxT58KUbWsDEtsK94j8cJbFF/Mm8/aRR
9vIm0Y6v3VCDNtCUxTLQ6I/Bd10Oou8GiWfybSjL2KbV3UFlukSX522oIS5/Fhaz
Js2OiQCc4xC15gA3+6duI0VDAOJFFXTEp3z2euZu9MR/PMNcyvhJkd0qY8HKo0wW
queU9vMyfwMcilzZmjFU+DGEgOMcCRuMfcdTz0QJmXLSNEWOgDqzHYQIQz2Ys3IM
qnJx0+qdqg2UyTV4KuOrkIO6gYO+priLMF/4N0URX7HxusDojk2TDMjRgLeEAwJV
9PDAKXihJWnekaMFpqmiO31zoTOnxlXRbkeWuPsGZvbwfMQ/HvjZ5crPi6CAjyUf
d8kp9HbKSmWuNgHZZFkPOxHrer9yua+0HWeiDIH3ZGMJQpi3lBLTL4HNJPpU42Z2
1LU4k0UIr2KBZQmK66HArOsFcLyPGfIwGwIYhQQk1LhTA0Z7JO9Qes0Yofd4GYDQ
XTdO/ofwmBawT0bV2GbwH3NqQr0tHHjfoB2729RC1YZUR/r8C6c0S/Ut39a6sarD
pxaSgc75fS1M/k91Phm4j5TnJ7p3Oeo5zUctftBK4PLJWKymbRcepNRhfdYNlX5a
0eM+L7UqmbeMV1SKqRoOyCGmgacAwXAcVTwtIIi0145vczUW3FXWm5plpY17tR43
Rbkvjzg1Mo13y9scL+x6+uCb9xgw/F72OLPKwPQFKLmJ0dUCPmzooCPs6CQqxzcj
9xLqCs8aB4cvXqcHE1LoSIQ6Qq7EEjva3cDEDjVUzkoBoatZkXyMs5xgYRWAAenw
pP4h4IsWNIEQ4NJyDoe+mDoKc3U6P16M+dO6yeMmrN/ESET7RCnchi+BdhcHwiG8
3k7N3R0aX6XWUKEwJV72wDtA5J2eXDqJvWOY3K2O+YO+iCSdC9L0oh4aeLmI3+vX
sDS+F+1kq3JdLBqXeWjMGaEgbVBdg9GyPMscJKTSzHbt1bqzKiVzFRyJWXHOOTr/
IgpJq286gBffvOZ6apoLjIKCYk6KIn4LzaZtbjz+OzuTMhePs3bBOnMVblLsVDjB
fpNeZciJe4Eh9gQE3VB/mG0bzjRSTRXn1wvvMU3lR0nJxUHe0YV93+JdhoGunkah
wjMUDQOHhXmKlmzx7q4ni/+ypKWFlAveSwUwDv2G8fkWxpxJnniWnQcEAYvWwtou
hILNMJtSlKYI2UdgmJhz0IFOh26HBeAEe0af3TQKe3dxNLZijFTss5V7uThHGmGr
wYXqk1gPaG51qqsmBZ5tvdxxpKDJ6J7tFAhReMiJOSHNBpXHwIpxLII2AS8jpf8a
uonqH2cGdDm8i0nmEPN2jU6P7VRkukvVaNw0pIIf/g0DzCEAFhxrrw9Tr9J5AoPT
0vco+CbHwbjentdTm/ncwmUjY51oZf5Y8aLBqF7JUDZMGeNTOG1zYxSS2rv2+U4G
+dxvSWPN9A8dMcElp7BjSi29MEvtG/qWR/GlDlfWT2brQ3VhYpmuVt5Pvjxnhc6X
U2bHncLf9IEcUutNrmnP3eIcnYgBp5C7Ih+jm74qY2z6s4bzqiA9mjDjI+pqKthY
belqmE+72kIIJDmcwzWQmQHUWobXO1SMPRX0qjrV9QD6/4KT43jYn9Phq+dEQaJq
jrO4CGUWBPu1E03BCLuBkNjQV6oHnIO7uNh9ufkH40KNuA6E5CEX9u/QE4u+EMge
JlFR+PVO1cy+ghUC+C4HMSW2+Zvc0Jo7L6moIaflTAj8LqNR0zGE+gy4mHuNGfqd
2XuTWVWHcvn2PP3Ok1kWwl+7Pk4emDNBpukJH9RCrPHdE1yFAGL5EISjcnZxU/vJ
skCu7ZkCsWmG4nDwOpiiGeZ9eN8dOx07wbyH6kaH1/h/RGw4BlgfQLOLZuWPH7R9
AR7YapsVk6WZ7OIIIa4I+8kFWyMFJK8/83J4JMljtyNWOSLRzL/tLFBY0B6FoQl0
LwUtEnHp+t384c+MkBUbKjAr4GmWDPjD6rS96SKh/llrWYlBV9/1yL07yngwuN+K
aeKKDvDXAOAq5R/TMgL0jYR8uT+bN631eguqJKWzWZQN3GxqF19RRK/eYmvpBuQ4
b8h9rgnU3XGEavx8nxCj+l0ihL/6fGvjAUW5FmlJYWdjj6BsZ3df74yuAlbQP0a+
xCaK8XNdQL1VNjj3J12NuzxfZo47DhPS5gelIahzTwv9GXCSJeIsmCx1EaIODS76
+X469E12z2SzLHdv+Rvgjw9FW37J65/97Km5d1mVAU28hq3XuYDYFg6B7NwtkJGn
xhmJzIary+ptk1oZx8DGhcdVE/HLg/c1O1Q5iG2SDDtSKmNq0tK4EpzjeGy6Wrti
oNAOHoi8W+9YTZh6gLBz29OT8tUtXopdW2MwqdHpQX0a7Eki1GlWFJIITgaFmG7r
blZrRi6xPoYDQsK1NbDGagsLjHmwjko8N9CVPS5/yAOzywCGLejeqzsLaGPhgMvJ
K2Vq23oHCnFrnDiOFV/EJAcrImIXD+eFkplnGg4oHcLjWqhhDMLxpj0GxraAbElj
Af4rQ72EnZCXCRNicDZsMJbn/tSORFptiWe89o38Q5XSwQhHMuM4LQMYhY9KW3JY
4oEOFE2PilFSimZyeHrc7UcsrR/4y5L2AYIXRc/j4yR9K3H4nL1rccuRHNzIqXNA
7L4RjPVtG9I2JBRVfQvf0t3pY5hDN1tPrwFBUsbyjE/VmiuYXImEb9aW/3QzZTwT
v7T08OlNhpLlKj3Wj1iArMfaKjf/p3MsXu0/Y2z2vDSFgFWp1wH6skAgjSjgsFgs
kLB3MX+NsnO3vTuDpXoCTV0dTEB4Ska66tm30ZMKXJkD6Gzp5eXFkhIQRDihPxfi
yAbC+ZTX/EuQ1l7/F1gL//ZWtJmXrHY4rhDMgigBSOMmfvOPva7FTqSz/UZY+PEh
sK9M8XTkxrunWnxO8cMiWhjIZUvSq9wzuR+U3YBKtjeC1u1JE7o32KuvBHYI++XQ
l40mE5O3RtqvlloxtRsT82tXjXHIyZeSIMZ+bMx8D4Y7nTZhiWTQVyI9bKUk/TU5
8sFzpVPR+bj8fYi6yhaFRnUk3QZbiBC4aLQZZMsNSVZ+8ecWt8QRSeYltvgd+qwo
VE+D7LfJdJZfMLO67A8TleWeVUd4lYYbriyDyRDWWo8pHP9pvdF0ilORSXkf+DzK
CXixua+KgBURNYh32TA5ofKmOY+fwpqlyEzBZnDWlNh0q0F8udH5WiOd3HvpY2x1
5Qkk/0tXDqMRokVDNUGfRGDBB7HKrSrgxUbXCZcTKCMeDOgfd2hejT+a1Fmeiw7e
srtAepqY3ZRYPk4c0UtftCMLC5NUqXJcVjOWzvh8JF/vWZRarfkHij1OT97oxgZw
MaMsRVxBpUC2euOV1HIQrYsJ1/PkIWEfyGz+bjNRUIAfwwLl0oLLANnD28f7giHw
iYYzVpKEJcX5adANUaGUtjR5sbO1hsLHNu6m18a+2TdNnEQehg7IISTOtbnNxpaQ
dYn1MKNjMCFU1zG0p2g5iQPw+t3SIJj2ZGFUkA3JAyWQk0VEg0PWd6wAvVuslI8Y
ISJjMhVknq9S3j9WOtDupJpGUYxf0PS4Pa88qvF9lw9keNelvQsNYbzLGCv+eAvJ
muq9ykzIZ6bITzaGrALvZD40Rv5vU6mWAkrX6QVR751CLdH1o89A6kXYL/HOTlY8
ZiCjedyCzsfuVFz50tBvrqYE5676xonDLHXB/0V9sr4RA43H/i4PAMF9JPC4ov+q
foOQfLOaQDhAGQGsu6JBxPZsgMwfi1PUlddf7aa4udgpd+LXGOY1miwNNnM3hvvG
iPpAAKUJi3Mm7utpBGib1bNp8eWMzmt6iH+6k7Vb9itiJvrQIBzVZpLMkOGw0exW
rNA2A6gvw7zc+L/CnfJFhaKNoxc5Sla85fJLfQHQWumZzAr2GekcfHxuhi2SPAJU
Hlo77//YDnxaZR6hi5JPCiJFj3mhwU5HfWvMHTaRt0EwA2NTlGR6KVWJMLeYB5BP
WVrMJ3pKNbcPYCeq3jWSf4aU/loVrkoCIztLxK18Sq5fQLFPmMx2CB8vh7PRvG7g
hpAn3WOJcmsyZL/tTv+rnadgvhUY3+Qdo42EnB9pWsKvSjUODea6TgvKShh8YpYN
yiLhslTa1Sjaej5AbT8msjZa92KabGdPrwIVONXkh0yBXRqgYDgbpzgScK19HpaP
31sbkT/7YGrDOINkW+gaX6DR1BbhgagCH/1VIqtUSrTHrX2rZ+KmxN+MmiWqVv4C
LINDgRisxCdFywfn1hOQOsjj6YQ3q3zSbrWkGykuEsYIpaD9LUS3wi/dNEgDFynv
kalCHxxUwgyAUea9kMbXDexNpmJoX1mDxn1Wxfw1XIowxPFszoO/yLnss2FstBqD
nyfjmvuh41gvWX+OO5dVbqkXOlfmRQU1BQLsJpYyS3JQlo6e5iCupWV6DxEvqw+V
n3rqIoA/45aVNNRhC3uFRBdPJGmPmPDhuYyr7py18zB3y9bDYEh6N2Oa8MjN7iJo
VtLF6xF5CA/yepnmOAExksDOPfR9fQ3aTeX18Mp/irLMghcGWh1+uABGhQWTYjHu
cDuGGtEpvFQXbFxKcCNVn9BVeviDGb9e6tqhSYXUZX2qpW7FYcV8wKJGMXHFvlbj
5LzsMU14fmxX+2YBgWwlgJouP75u2cMgTyd1cRneVFpgIFZ+3jcb3Z11nDBGEG0w
MOkFaIEh+UQHiLYVGDyCTGDd7tnVZGsAfTbwhYjO4E18NthEjTPA42vJmSlDSmvh
EzzaSZfurl1PflIpAuczZO/7dxXEF1NT+M37SwLyPVbb1rbVXMxIWENKvN7wxXay
oj5eyxOlOJ8V9Evqxsl7buJXSYFPM61thR0cksCabHHQbfyblBxP9szyPbtQMuY+
c4BI/LAvKDHAUaJleTBWnqN4IeIUaKv15NuAMVmu22a/WxkivSjRVx7HzVwGd8Im
BOCo5EzDoPghK0gvzsqMtimGzZu+di/3gJK7exoaCC1rxGfR+L22TBpMFtk8FRtl
oqc0HgUBTYiOhbTO19D9KMq49fgjRbNLGOEgsjQP7ZGxWYy+8Q6biQzWvY93xqey
HQ363eqeG21VONue2t+qd1eEh7H0G1j9OiDJW2rPYvXHNeqadUHrkofPm2o2nzBz
Ae2KShtZSifPvkwWLG1FhM6OD1uIoD79ZsGtFfeznRe43N0z2C7w0/a/L49IxPS+
0Caj4MNjxX16MHTvIsh+a4PCJPRuaXV34VhGf7edXNJiLHT8umvyfyHg8YGv9u/b
J13xA2RNNzF78ykzsFuCgv1Q77g2QxX2GfG018cdAQ875+wHX6aDionUlN1eNFfR
z+x0haHbFW9ABtylwimnL22VbLnNFmcaq+7oUFCadeJsxxLJI4EiQqHeVuk4tDKf
zQuYsFbLAAUFyOXHgX8re1/vr7u+4nCaFLVV6k0kXzPNL0OY0TuLb8DTnc1saMsw
SczgnlGvEyOaRRF+ktRsq4Rv9fARiBnL/+MtxiIVwGlEN+chLFwJaTEjXT9J5TmG
RdtuOJggZRPLzrhYwGIZwhNQSVrRThaxQPRmkT/4AtS6C/D05xZl9430ROHkjwy6
Q7tgcWck4+bIXSJplhRemGvPpGgiVxgw9TNt7uhVE3IOw7IKYqDsuIp2HR773wTK
ZMrWoV4uEHHf6Y+w8qVQ0ixXqDecNf9jfjT3hUsyScGI6FYKnfKheBPeWMgAEuUb
/+w/JrscEl4YygYbkly5kSgb1vJjcXNBdJg+zDQftaibZV3hmMnbU50DSWFxBAiF
ILHGB01xR5Dw/MF+cLLrKWa0U+ge9JYYYy+/msBxfR1otcDqAy57gBfbSxhduaMr
Oj3IUIfnROqZwRsQt1ZuYK5pH6g0BtfQ8Juq/8n3OVlZG4tx+rEnN4jiH1dP4tYj
pmBPay/WaPV7Zum+9D22nbj+yeFMsR2UMA/darlAcXuUvI0eXN/PEo/1bWSWJbIO
V5YFFGnDtM4u++rPUm1dc6ZFvqu2m3uyIulx81KXowK+YqLI9DQ9xu6h2j92Vpt6
iFTANIr2j4MTeIBhQ1bwaWz/RrbrHAzrH6ai2yLDb/JKYQHDSeAkQtZ8pGsiS3SA
LF+aBLelyLHTfJE39qaILZzmHbJYPk0IKBlc9WLGwTlDQhCPtcb127KDZ38iG0Bx
/J+ksu/hARtqaUCBJl7EVfazb0ddp7z4M3kLKlUz+SQfD7RlmbGffutesMu5gLot
MJbNCS88e00DvRwWoyFjfZuy466ZOldJMFsrzERCtLmpieJsKBiI89DAEpCZfAkl
gGqkoTANuceg9VOBJOn0sGEPctKyMpbDwjb7IFhcNgjLf0vmZwIOe07Yiq8itQ8W
T8RwjSlYwxEVT6vBXea8WO5zKMYsrMy4l6a3u1J0vMcq+rZnOMOuEEx84HjANViz
JS6o9XPtth+V7e+recWeAfedmcqMB1R7ScMHiISNohb9boe1cPSLx4QQp4vMmIwR
sTzIp8Hpmol9J6YrzvD2sFGjYabpciGA6y014jn7ZDloTyk92DNMVrEXBUVjmqWO
M0ZY1zZXY6H4NH1cynxrGTZNC6dAn+NGn69kUFh/rX8fkyXdOdJ5pck9C2zxUIU+
DvCpEQoDr9uzESwBqIk9IbL8bnYqsc3gc4n78O0VjB56vtz1K592AE7C2qwWv3F+
5V8ofJRGz0YtHIiQOdIsR7Vnmh6wdmHl/BlenAL9VuJBVMdpxqtGk5pke90pm0wO
iWnH0JGE4qYyxw8H56gQFmEq6SSf47Y5ndJFZTXGVXXnnrlzEymXFKX/ZPrEgsLU
yYNJgP+Q+8xnbr3+XWwLE3dUrJBaZXkuNHXoJ2EwEetDTrPjCxvF1xPYXSOfzOcn
lps79xpQQLCOCdbygMI5wdGE6qO5MFHBmZq3oMAkDQp35RMAFhmyjho6tAUqDZHJ
G2KUR3GuuKaCb0Th+QH+l/gBMnQjzbwJcOTCjBb4mjwb1+sWMQ+eJNJh9aykrcm2
1YQqSafxdAjnbTSpBNv1PfBDe7rQQv9EVQXa87biJL5hovZGCL1h4MLGHYLXqg1E
/EjvrS16HNSitYSL6sNqenaeyAmAnBbshnvFcjQhMntvzsdwDoOmiMeKjJ5OG/oN
qu2JmmPdFO6H88JqfJ3LvV3y/o+KOtdxKsWweF7iZE1rBU0jXF5XtwOPKVFJv5A4
rUnygHXl96lhOw3m8yAoDoO9K+1iza3qf9q+W6QgK/hB6qox9F8dwjeQHI9l4lVp
JR93OYu7MTbO2fcWhzUleH4svgluwIF0hzN/TS08tukUiHwfxVwnK6zRptmd0ciF
BAZ6sdjzdA/AiCPF9c6ATblVWp+v5mcW1aTAIYUbmNr70vu51p75iEr6FsjxBfVw
csu1+CfZFstEcGg7TVMV5cssEEsy9IuEokLloIVUUc1tgh9mFnNvgGM/FRuqF5C8
AS6jMXQdI/yYsUl3lbuXY9yEWDC7rPCjaKlsNZPmc94SxmubdaUQGp2DcEPhaa/9
tpba3YrHh4akWCbAUIACa86BL14NV/B3pTXXn/JJwdyx/3Bu0fsfYLCJ2DelAi8D
UzTBsokHuy4BNVvrixoHxD0neR912kdX+w5bS1A2cYau+67OYEPb6QvuHxgdrLO8
hD/3kr2m1XnOybMdzQxwUYkTIdJs4qBoz9W0gGgCXc+bqpvxQix1zHVm4XnSWaYo
g25kLRO1W4zN3NzBZ75E51AvgkNw9rZAL/UCyipQ6eAJGVpNaMfiJxMOQlTmlIme
A+0zlnGPnr+Zp11CHy/Z9GZYP6i1gQxo9WdhLVNn15ykUzwROFhf/CzI3RYduPkm
b6zsOJJA7no0zj2R+vHdlx6473p93jjQu6VLmccZADLu2S4YLgq2B4m6BmubVJZt
cZtNQTaR8W8DcblBPGYQCrNnHcRlh5T/QihCdpdlJ5jVUUXvDuAEAKTvvqzraN2C
3K4EN///tMGXpR1BADqg+bydFbUEi0kaDH2lrcMlB4Jng30goPKtJqd310B7s2cE
rWEIO+p362Gcz+wKt4X17kYLBXb5lWCYjslXZK7WNZIIxx4hQf6BNWROPddjh6tW
Il175TuM8W9AEinUrJrofo58TVIRTXan9r28rEhBpOlbf8T9+MurNhB2AJkzPCc6
UQObw3nF2ms3Cw/LyoN62aj0dmtbsDzB2Ccz56l8h2EXgaWJEtFJS1ua8la3d4eJ
m1QxyerEQAAI3tHwH/M66Z4qTuRUu57bp8EdvlrTda4va94Y8o0cihhUlP5KqkO/
QvxhowSeygnKUiDTPiFw+ln7PcmgJ7VqezLzgbVMuUA6fEAQxSmxXH6WkCdGqiXT
0equU9uCIbkwZmVf/Gts1RMIwVCobEhhLZZN2iFe5fklCQ6O8FiD+v+vTq82e5is
tTzzxGOkEE6HBPolLZYWmbEmtpmHZQSWXvhdG1Ug1QGGVWsta4qqkTpvs/feoLa4
7yxvEqw+YVBQg8M8BPwMz97xE5UnSz7mN8GJUKlo7dw6CxKXKlZkp4vN2enDtnYN
wEtBqpyQGEwBFvL61QJTa7X72BarSx9Ph/bcp+1wOP+89SB92rWJRrrsdlzLEgua
NSP+1lfXWmItZP23i7+IN8KAYL5Sa5eoUedYECy6fpQcr55Wt8ap9VYEY8T08seq
/fM3ZBB23bEK97ADZr4/xdM1fVXLKy2I5SOC/uyjCfpKWs1zQi5lcmQ6ccBNIo0Q
GAi1hqAvmhBiTUFBMaWj7NC2K74gUuK9lCMALxh1XkaYnoTJBx1eJxJ4L3a4atsa
iUjxZQLnbJ1TZyzCBxanF+zrOKoL6FFY90uFvN0tLsP707DFZ/Y13Dn5SNqZICuH
Kg6sCe1rE/A75u1/X/TweyYe0BCCpqxTnskhDmOKIB20w70W/rixA0IchkGn7xij
4+EIFcspGW6fIqRrr1jiZynNgiAvkjX0NYJODneI2JgtXFd3M7JSoMmsSBis7i83
IjoX9l0ebKMT0ww5WDiYvCSF23F3N7eYDNn0x8Sr4UqL/FPkCiX65aHMo+pk2k4U
Ml9VGr8G4jGKRwLoclc0ABT/CAgN8KkzK4eOMhp3aR3ZJt/WeNDflhSE08McaANR
b479nXZEymTFZLv33xgii8pRsdPm6GNStFdBCEWwRs2O1IMTI4249nF7bLKXNeT+
5kwq9popL+0GLTI5fYp5CcISB4IHHSn9L5NgnHrxSJHu/aAmKcxGYAWdF2RHo7HF
PXfIr3B3u7GZC0ISiPIrfVaXiF3qIOeISPjHfRq1uwqNXQKXLHmEAykajfMCONBF
aIvumQbKAFHU307qpnZLe4Eg97bioH6nt6uAfbmWNxm8d21gj6lJeI6Oa/QvqNB0
Wmqjx8ikq0n5RGonVhzHHfSSYrk3g6/7yjx06uAjuvNCYit4szUtTfl49RF+8vXJ
Clusi8eo5DcxccmQzmfzGQudzo2bIuaOBSCRS4oYgBcZ/gD/pt8OFaKVY4RZVE/y
3McvP5SKd4UiT7j52Zqx2OXAeVSqeq9uauHj1DK7V8WIjbeEddyVTlB4tQx+sYYe
PTMl0Z/PMHU5lPx7FjHJ7sc2toYmeN8lEfC8GXktsZjiB/4jaK25dMPC4941O6gr
FZk8Qxe0g2lL8yQ66YvVttSSb5hEAVTYLf6zTrt0Q5Zg7KDZM6NX6vTHx+c/6yAO
pDoDsQWjILcvTJD/Is90pwlxKph71LQ6vVP0N3jZcHQhuVudVSVigFGjaWl6Jx8z
hSiNvw5ivzD6iti37inSYJevTxZHzvI0Ay4yZIMdvMpaIa9rDBx8/EZsxZ5mF6nj
DXoYw+4tH0YNu8bI7QdBrnJ3v85FaKLKB1iYNHZQslPsDtWTKV0a4e/vjhhGJQLj
lZAnK9aqRiYCVXOx+LETY2712CCfBTk+ISs48Wc9BrriXCOM7Fca45ayHf/NVP4i
Qc2L76c0N7gcf56hZPwjlH8Tfha4CQKs6BMHhcUEgCm+R8E7oa1N5AS/l6KIqG01
LwrQKCEzM5mCXqujRHZqsb/RZb9K8jshAwP8Spz5bCes9kdYAaDhT/roKXO8UM0k
a1nJKGXWvEeQIQROZB3iPVRHTI8OfAVZoiOgedVq6TclH+iyeiDn1qTSuUj+pSF5
TIOiS3r1zbvDdQFSvsjl2LwkmLi6fraL6Omr9hhEUkOekAI0Po4zFiQX7jxgvSPK
Go+2HaJxm5cngGeJHYG+m+cE6Pw6XVXfNxIGrrUuzaGDgz4H2SIgJeh8iQeNTtFe
W+SiTaQZTZGxrui1oJYxDg7S0uaPpOVA6uZUW53No7gMgEKcviZiLjKT7IOMORz7
ttkpmJiXmLp0SMZ74A92RGWcCUeqlKlacAg1MG+Or0tL8Xu07ZlZvUM7SC4kliQV
84V3YjVBrjjnZTyUKH5254jlt5/VTGS/k3QIfzLZ7j0NKO73MWJq6hW/rDoPiu0P
eRnJp6LAE2fkE/PoAR7pwed+lFz2ms1QSFkxcBkaqqlPr5hcde4WZwneKqkToZLN
/fZyVz8LLehjuuCB/PRP82tgRk7lJRqWUXqTHyj0nu8+DKvV3CKvrfHrmMn32rZb
SCW6JiGP8NHQBfBT0xQ3/pQbZ0/a4xau8IgWyf6mpehjzUPnwxVATo1PhqwXE/Bb
Fz/6AGINIsd/Gz/Xqaq2yZ49U7hnxPoyL1RnMYNbpfcBS5lgOctRDctCX8FsarZc
FEci3UkEpI7lNWTBBIG3TRzPbfvtUJCi/dAqoO68PxQ0u8jqgpjb8lYhtf24BNsd
qyou4grzGAx86rxIBMq034s23Ky85cBRvfaC42sqwiRnsju/xXDkbFhnirw0eyxY
aIQs02pWEiMAkMgechXB2JYhtRcN+ZjhbwH+QavUczvW8cz1iJ/Q4xqryj4XyWST
nl7Ew/8l7R8xWXzp9IqAMX7/vUwgBt0SGwsKiBv1ip2DYzra6MVGUBWYkAl2+LYe
F3TuFY7F25GZlxj4Q1nnYBwUVvQSBmXRS7qw3Sil2TKkz89LFVcAMGgL6CcEujSh
OZ60DkJCSYe9G5WRF/1A1ePYE05VGoTVwQUSQoYYF9KvDsRXNKaYtq0gVn6PvK+k
Ijq98sBIraM3rRg4vY/4w3s0XSD/6sMuqZ3Ww/nrGWZDpYoXPw3fm3j2c+mujQ55
WD6kVbdB5G5epcHt8zQObd4jSu41k1fQyBzwE2QnEudbaMQ10PY5ss5sHNTmb/pY
ywDPaxrTiaFa+rAYs/D6OnE4AXyEQRIljZFPQedm29+ImQr9/kCAIyXTcwS/ohW1
qZYO8pNqrKlEhpZ9YewgbMJ/43czk72dkM4UozEpKaP314uAH3sI+OSJC+t1pF81
TAOEku6meKF9LUoy682LoQjNdOXQIAEAwGSiksVp78T366P9GZdJzSqgDfO1HYcn
VSbrHDZu104f/gT3whE4ee/lEf9cCVB+t1WEig2mUScLv1CA4+qx93Hp6gBD2pmi
h1Zxf/fWLjPfJp+HPCHyQDexfsJ7dK5WuFsVQGj3yjmtH+QJN/V3c7OWqjgAREBT
KaJFST+13Lgr+QPOveOa1LmUJF+rDk3254fRn3jWSAbHleAkvepjc22XUBMmx74E
f1Du1tu/LW+I4SfhBBQw68XMj6Yoal6k4DVYVmWRmOCP0ONvxnt+FZiucsSJ4Yx1
DXJ174GOooo7eVsvAOI5t7WddnRVWU4nMd6DOzgZiyAED97xi08mh/Ea70oOjmnp
Coyl8BT78XOrBccYQTG37ooI17kw9ya46AK5gSh1jCz0zen8s5AGNQ/SintmPKBy
1hriGYwVWNuG7BhojQd5CVtEtkCgM3/Ux6We52f8+Ts4KaO72j2hktIAgoaxKVUv
DfHInHZmpLkWlQ0ZLreEAgmZcXm+xzFWkPCbzM5YaFNSnLMiWRvSqmC4Jvi33wEy
M/zSa7Y/XZCA8eRJmIG+VxEznEEU74QTpEqnj3jjujlb0QM5y/6DiJSBkXOWvr52
eiMAhKNJtMmX4ZAFMS9GZfdY3sPuGj9TJXUiMQRMvAGnABcbzuXJvxTmYrON7KlG
LL/9E8kU81Hq1k9tP+8QThxa40DERb7Et8Nwkn+CWM46I68XQ1SRE8/Uh0e0LknW
NyNR8BswIzGRsiuKD2YNA26Xk1x+Z0jnwsy16y+fbAFz1aCtP+c8OQOOWTiKqeQF
HXT1iyFJlIPpmHAvKvPcQ4BNQHcSoVzTZguvQdGmDKAneNZ8bg/A75q7cwLu/bdi
bU75sjSeEpwlntuK4Od0tR7T3G2KYYvwtmSUKO91syHh25kgaJHXH/pQODG5z/Ys
GeHwUcs2LLOGSCDzontrUPyCXNT/1N0BIgEf15rV9w0raXWMZ+YhESMKrTEo4qJZ
EvcfNR7nIgFqzsN2Fe4TD2bEGRZlIDYOMC5FKlVmsbNkEpNd0Mz3ZDagZWlPuvd5
tPDwBU6YYTpepAo04TNAoM043/SYIdKG5FriwJ4xpfVOIBLSvAy4/PdDXI0MdnsC
RFN3NC/rqOK8q/gEgiEy06kIpRe0Qt4x/k2L28vhVzmIATGQVQF4vHc0v5tD3voq
1yViV5ByVwHS/SPB5xjx/uZWTWNJcsdd8SxpPX626fE3TE3Cn9DOsgcTtm+xZ+by
l0ct0lwm7AASyqtJ78NQedfkv8PkjjvTtUXGTDMhiRKQ//Md75ox6UEg430CfpHd
zL5nbUwyMVI+wwvqtMsisj2qpSflv0abHkYfcadytlz29ur5PttieA7xTcCYHzB2
+r78fzs0PEnmfXRl4UCum1KXpZvAx0/COcjjyoxpav8TvIAx/m3UwhxW1pAizMRM
TdY+7BiPQ7dAV7bnyrLJB7R/6PRLuNoQl8CRivy3dzicmo7LVE+6sydN6aR8PRdN
GSwsZWWnviubpJi9vONQfIL98C05uGdd7xvNrqrwkymIFb3E4HEK3tTFfHAb4iIl
FiCa4SQb1Eycgew99HK7dcT3Mf8YalF0+lGBTr9qw1qHii53X/1U15oOORxz0IXd
cWI7OMUw4oHT/fw7vJi39rmBynKY+w5rqJrqT7h3+EFPHKG/E+AHKwEkJKVinDfR
RyB8iPcOcNuxxxO8IfaNaDTIEW7IZ+lJHGqe+OqXKlc3EXEll/oInoU8FhuywYtt
oQfNbd/CUnk+45vah1jGqCTD7yMaGfZJPgeUK4cLivl/IA3KeIky2BB4PQHW+sPQ
9ASn/oI2HehIlI2IkJfxrJlG0Ld2NrcDY2mmixcTHFRmUwkTd2wNMzufty4tzMdc
OtCRFZEkl76K238wyb6SS7RvSG47RhA0ivVoKFu23mIW5dU7KGyeAtOPbevzezOV
T9V5QSdcT3hVfZOTf9zB/hL4BRUgO/leuSfxmHDj2XqcW8TTHMfHavE1+RnRE55p
5eOlyiYU0aaoLQaFQ/Moe6oXFDnXZyWmSpfoPYHGXwOHEA9uzu6S1DlBSetyaMYi
mJWuWDVtI9Xo3RP3DnLD5k+mYECC0PCQk+dLzF77KJmql1chG8tiBnEKWEQ7QZeM
DS7Nro9iyQkUarf9po6D866mhqICksLhoLScss3yq1v0jRbG7M+HC4Cpl+Fzk7L9
EyRsXgnUIt08+/EDvoQA2gOmlpGGyydyZtScVp4LQBlKXQvUhsacE6XW9AeLyddK
ezXKB7ASkujvBea4zA3VDzbT1ZCePDkXTvetSYU80+hbLzURHTXROAoImpmu80xJ
00smm1GffqJ7z+YgZGAHcvMy08RAutnNCSxwyj/Gebu/B4B2uZM2qmtXt2U4GGM+
HkGlTdvmsWtvWquR1LmQjohpVpS3SdmPXqIwtXKHAoxD8Ar1+le9FmNlVfUO6CaY
ILRe6EoVlHrwe9WA8b24fPE4j6slz30XDZo+Pn8G65tmHboenSNYR/612ysc8nTA
2mccFS1e0M8ANXzMbvkLiwPDJnilJqqXeAPm9powLiEdtrmigEv+ZUaW4fdSABK6
/Ox9smuKs1R7FQN4ZwU0zXWibAfWMzOg+VKYtf49hVJ7YL5fstxRCEqHcUj0yZeX
bsQnFERPUrx5TgkxjRHeAMT+DNNrgzZgg81zmyKNOVXnQLbEvNN3/pBHVbBfw3rh
XwdGT2v2EKgjQZjEfR+8MJ4K50v3e6w3OxhE8ZXyEF1Gx0t3Wu+lJifI8AMLoZf4
s8JHzMOI6iMCUE9DWHTe9R8Ek2WDpZNRbzNc8x17qm3DQWPz3A+76sub2+DJZhiI
uuonNP9ylTMH5YVOzofOmXndLv0CzVf7jr0/BoWn8xTybF85ThBe7+rH15P/RcMH
1O/t/9EZuVg4hXr4FB4XIGl5beaDiGNijkTq7bd4st0B59C5NAL0RLab16WLnvP3
QweDIZOZkNKvGGIs0/F9AZaz6rv/GZgf3LknH3m+jCvjZ5qLVzsYWTqipT+VPCE1
GJAKf2HnNJNBoMSQeeug0qyJqqiWTW1kjDzH/d9qg99gHdPLMBiNfLUJzSMt9UEq
FYtd2e8VQYY4pQxqlBZsZPbqql17cF779V27IFIcBBKv6ZrPLjpECcKeKok8Llhz
giMF1rS6vt+e7pjSb3qxDK5Ma6bFzESggohtq8FqHE6KsUYYPfjzPbcn4A0jdGWH
igmeKWDaVPRR0o6f+YcAkxgoRwJGDj6JTL5WJQ9dVLeMLiM0fgk25/3MBoFjtoYh
BdGMVbQhGVsYwVJ4X25Y08nnXlN02W/hCloUgTtSxmzjPRYMFyRtgsW4ZOH6/JON
nLTknXgSz+oCSlfmNqPV/X+RgsHhYzyfM62N7JO8LCep+RoLqyfv1LhVXxBV/PBJ
KDK3Czfb8BEQWkO/sw6SyacStMd1r/DKpKulDvafhPNgr/kDtWQg3kDbMyAOk+4K
HD//IOenawPR24whnBqyhqgeal6HxoV9chd0s2+HQIC/zp4XU5NAwVhoAV/40uZb
OWG62WecHfFqAiAz9f1Y0DtPJRWSdfNiIIy8Izk2ZYjvxsXUOo8nvs09GaubrsYf
io+3bGCDHOQbCkjKEmdovD1nwVwBbESJpQrj7dGs2Z8w5H0poZ5jdwnugb1Iw5XW
aLHM7xwOe9jYmzkPQZFy2xKXBIjzIhF/pY0PrjZP3jmPYUQad9xib9SpGS+DXraU
ikA3eOyyy3ACtqOhAkbnzieCTW8hFM9UL5NaeRAErDBUbOTZHOUJpvR7mw8PZcJs
aaxpNogCWqLEgdAmSq7ww9ExSeCYM+GIIYjaTybwFyxcR6iTCuQ8ZziJEGXtlTat
HRQadQJgdnQuTLBUJgp93w7N/ZbS0Ym9J6Rrpxx7v14k4CZ/DGMwV1prmfm+GRqE
Iqq/XyGO2CLPW2NnzUd/VXcp91Frj1XuTBnRhvlrqTqpdI+aQnjD8DHOsM9/slKr
6Yu2yae5ulwLS/bR1CRP5w6+rprbNJLim8YJVdkSiRIUr+1xTG7yTDsYKc0/XUXk
TW+uH4EN1O4Quu7yOQuScAP7EqN0qIgLKuGF+fPg7xe3f4H3oznVvO1tF3EUDCWu
PRFjA/jeduOH9UFG1OdfIO+8e7WmVFAmnBoc1JHoDFKdGe6CQ+N9nFI9eIdBaLjr
ohN0b8sc7Ru/ZUekuvZWhncE52X0blQ0q7i2dWoSYhCYc7/Qy9p/Fm5lahiGFL9H
lShTZavuLLaAbA5cEU8azvfq89Hbc4DCYuX6sZFShM2cligJEe1oRC4ib8aFah1H
kZ7GcN3dvN9SYkqbYXzGSvV0YUIRYpwqHHBVSpRNxoV+JE8QsNTNe8cW7hKgTj2s
n7FaayUJfE7iJOmjC4grbOHaiIvHrJBVnnwumWNQyVdcNfFOZUz/dXOxT7PnJl9f
XtzSV9/jha/mqDAcie9IJ/YqY1j6zt2lRDs0MBBSZmZYzTZX8gzbvtIx8e0jqdNv
qCzLpSj1enPbwnz3JN/M9+2DXLovEEHIwR1EwlS9DFy0hyRYjTfdjlTOa6wRcFKl
URHfIsb+HtkwVD+ioQKGv7b8ArTXgDDr4T5jnCaYtnNPTI5lY56dC82ysk+6lIzg
9AR9Pd8kA/f/aZZcOeqpL3V5/rAIAGI1Q2XQ86h9lkxKP0apqYEvPqA7lYD8l2ze
RFZHLFo+C5Vscd7DqM+t/Vh1OJIyV63Q2xgoBQdOt8HUmHjS0cDVdIvZqOEMfRP0
QY4sNjdrb9jQgapZANS1e9OlApozM2wH/8hD3lXnilCgHhVMS5eOh4YfMFk9G0at
/tel2VLZvIcefvC2bBxBOshbUUEJlTX33O4/n6FNuqUHPVK37yiO5vtX1q2z6ELD
ouJPrCyXYDg7NeBTO+w3JIP6MXUOBvXnfN6TuIP+BW4xo98uARLjcj0lrdcl7O7z
mNzUwhUMgh4BywTQNBR8aBS4eginAF1GGUGYEwmO3Utgnu2sA7vTnrq1+oBuN4uL
GAekrkg1HUpYPOU7dQNmptwk3gKiwjaLFqco8wAbjFtzb5Z4FyNiqMyVzfL2SfpK
Zm/0kI4YbafryJOEcrB5lQ+mpYUKv38WAQYbxKevqiq5fwDKxPKpjGVCSrx4K/pm
+z7+MrWJKqoBcbLTySa83B4mpVQeG5VdVAUplA1IE43l+t5lKg2BMA5+fIykEZmZ
Z7JCfCHSncDNxrZHtpXazNo6oqXsgr+B189LNnXE13vYIhh2TdLaioI7CGJ2PyTI
HTazXS9Ftzvg17gR+I4u5EJvF3q4ORxqy+2fbryzl//ybEZrK4DWBEPj02tVtrrI
TuAAxPfe78W7jpKFvaAXl1803/iETOCy+H6H2YlM1pSh0uXmNbSTHl74MEDyiavY
VahPFKRQIB2nhBt2Z2YdaEu+ZQMAaLq9LnJn+f1U7YI8n4wTHTGeH+QnQJaiG1W+
NFwGxwhC0AhbKYB2rWjlf/IXreCMCMCm2fi208dbrWdhvrQdA4zkI07L3TVcVAAG
Kdf2nOAtXpay1G4zNS/Zu7bqJ6M0N8BrJidiPu0u6NqQXq3HsrJ6pDvI6NY7+Skn
eBRIfTMn4mK9PV3W544S2IwodDugKkdkd6cQuBM6Pk3WDPpJdg+wsK+22+Nzq4sy
932bv433othZqXVcFXLd9be4wGSkhyTF19YES/DLro+qVgV9x/hS0xUKuF0brfqh
2jt2LOdfoQQV3/J0ZNqJvXF9bLy/JC8Arcel+FmIrO1LkwkFx1Kjt2/Ljk8b5a6J
Y5KDRIJQ8lRSGhD6Cxah5e5xG23MNCEwoNZTNllqFwWy/r4eoEwdCu/AOziJrUMO
nBCUplimFe28WOGnV2KRWuOHDAzGC+d8sVVjm/wMGnRJhzoGj5PBNUaDgcBQGgGt
jGSBPCP/e6DR7Csm6iNf/3pE7s1Ld593O7bXxTgHqXqLprE3LUW+kAjAFI1V+l0j
PGDzVXhVPLwiEQ+Mjn2qVwCwT3CY/SrUTErR7skWBg2nrNV8QUF0bUAMRuIlLlOH
JwwzTqrx/LJITcVGJ5pvJsnGBGuGQ7dGjrJMM33GQ4+IIQgf/NC8ppVKunkLKlbn
jvCO/QV/gvftsbQzWSHLoN025DZn6HKUmAEng2eGfSsfFKIUXuWDq4PSo/r5lFuf
En724Z8LRrLLsePWRWK23eUPWY3QZPP9oeTLhl1cNlwsF8xyJhbwhU7+rBe1wr2e
fFCbD7X0xzIRGvrDiSsSvREIUKrNiUH0nliX91G5m/gZnZAX4xQ/PQnZus8zI8e3
6ApJXibe3+Lv9q7onIoWcp7HgtoTI4ZJNJcUpIo1G7D9AN2atdYiX9lVA9oZpHzn
nA7RVv02WDw/jUyy/Ous9mzFHCgvQJAXkQS6OUXlAwJUTjFu9UBL7C7zPKlIg7cH
5ChfbcJfWW65mbCFyhP4k7uHx5U2SGS7mzbPFE30NZ5/kHop11LYcsqfEzx2Hspj
c7h7gmhnmrFb+L7+hUwNW9Z4lvz5bDAccPQfOdEDdG08B/295Z4iOY6LEXiUVkoC
4HZQCUgP7eqI7KrZE3wyCb6qsWbKz3UDoi8kBn9AD5/mZFeZ6NiZo5atWGdurPn1
JupinWsk4EVbs5A7P6pJYZIcoto+APupJ1ubuJZLPJZ3wHzpZhwN50hO9W+c11TC
2JXZVOOHy5uvVVHWDRLsL8I/V0zl/Upmf4ha1yuO3SWNYmGcMGUfTAwqko45zGmv
tX6C/p4WMo68XRWbAm2qibucDf3CgNPsKX0z4sXylFnIRuk5A0PURw4qNss3i36F
N5tBTNSm63112YCsykzndy46cpJOAuWyTdfZoEHmcD4Ux2tzJH2txmdfgeQcb0lg
eVfpB6NqO5qwouIUZhaLGTSyHY0UE11Yum4KeBMww/gvP5Rv2of8DnpBvT2xftni
3DZeYmdxtppm5OyRnGNYjoURsu3jtYkklV96pbtjkWkUKJkQV16c2KHawR+VBj84
r3TU2wIkbjLHkZOYemtXCe5veOW/TluRTAqGiUGTd+Ig1H/TcmeJ6YvUAVgnPDEB
j/ewyvytI4kasmz73jR5JprJt0tZ6gfdTJX/loSdw7PGBrrjUdRbAHL3rHzz9TPg
c9OVMvDuCVbOTyTRxHeY5CUTslbIUJ0UMkqRj3GXeM+ZUC8RlCvg1iq5ZuxKd966
7JngJEQrTJ5vuTm3vpFz3LtC973kbuiVb8qRxTJCxf5oLwCKo8GHfjd6u0oAqJKb
F7OyFO0HMaSubLnHc0BAeZEd0cwLl7+xwZbmw5wJzZa9CxQ8KIPSEwI8FBjwmDNE
b13fkjuJJhl5qU/ykgjbISjU8x8Cm0uFRUuh1ghnER+OaEavc9JnICYObHkB73Jg
zujP0xCOGQ9oSPoR7g6L5K9jZtXb942i1PYc5qW49NHoJUY5rtriRJXkzC+EXAXc
YlQvSzEuz0F82tP6TSrqFY/D8Qkww54L8CB0cbsbRXjop1jdUkZNvoWrR7A3Bmp2
5DQUyHxDdEZjpXFf8bepjwmjs/NNbjml41K7B5qHNmT+kuOmc2UWyaRKOMBlVp9m
GYS1/LUL931wz/Ryh6aX1fHBHtRTJPobQ1d4Eu/3/wDXJPGfxJSkp4dtjhV1ytgB
aRmr0waYTd2wbJ7jDhLnRxPMPuX9OTJv7YQRlHWs7gcYXzCW/bWSwVvqtoVAF8ol
Qv458hJCSzj0BQ9fhmCQczwyaMh7v3zBU/3mqZiRChPggIqq0NFQrg34ASG09yUs
1PHeh9bTTBTnXEySaOsMjDdtznW/0DO5QNsKZLSdQILV0zu4H8dtK5ZNPc3r3Ox1
52bK6zgs5YvFskJamwx5HsfIxRTPyEZJHZhzeJFCcLCRZ9S6xL2RTjnyAlCIkea8
gm9Wz+CKxZJtks++c+kTOfJpZQm5grn7seQK4K4Y8SwkKx31eWBpoeYKsCUzS9KN
R01i5znuvAP9xGSRN1DUY9vjTAgfesceBWr9IQ4zLzK2FqaYAs91Sf8rUcBayq74
BYx1nsGnxplPX5GyndxUkEWaPgJfIOva8ROQfxOkqGNvQ11eBreh8mLjRRuJ/oZl
k45Qd4QgQWTcoJzf0XuVUAWH/BjdxwZsqB5PUA+tbyJ7PNYExdjI817cXf1u2HtB
tq0pxEsNbYdfgC6TPw9XFge5hKUAzHCRdmuQEWnB+I/MgvK/x7liAtLIhnYV9Wki
E/tvD1Ag587H+zvcYCfRLjTJeU1gcoIpB5+1fJ9W9cHgFkVdJEggqnNuJIYQjEPX
mam8q5XtVIDIIa4SOxnLb0idXWi3stKv6+I9HQBuG/LNWuqurr9uG8QxOG2wsqpL
ODwCLHzCw/KcIMSkz52dhacgJdfZtM9YuBOb3X/2il/f/EuynDp3Oa/6VTF0Cyyv
YIa20Ms/puLQQZWy6ymE2gRiuXUivmjIrG4BZ34yan4BTmrcSL1T0LVp+3iZMw81
PELeFeiK2k3tZkrXKliFMq5bqGrjFMjiO/56rHeFewaBprrs2S1k1ImieCPptdgQ
s2KY/oh1brh+r4Xqn/hRH3aWNfvKnUDBq6laggIwZiLGW2YRxO04mnvg+2nFQOgz
CKeE1Ju8ycee8Yyuu3kQ4VvHtufsfy7Qy8m7Api7cVcDWAIikfayfoUSX+u+Wzoa
cD2ytUcq4W6E7dIY7d8yMlfQgm48qu+X+dsQrtd7q7ukATeuasCKYNBt65GopiVz
AI6p9nLaAX3UjSfQWM9luUwmTgJoAqE6d6l4Ei5znEbB6NeyxriftzxXhiNwSxkr
/irayAxGX8Llmo1AM0RZNlfFKqnYgO0jVku3vNealGHT5LJd0c9E2fMoCMPOdwK5
uC58C6Lt53f3vPG/AGTCLVphQpRX+nqtcj4puRUzE3SzBT/dtLy8Np1IOo5clbLG
ckzxNU+07o8X6HXzqxKoT6LO7k+aawhIdwmLCGQGJ5hqluaj8YOsOy9YYhZ3m90k
UFYXB/6pfTP8yEXvnsBdY760nzme2aZEG3NTEXWxASgxtZugPgsKkHjBisYtynGw
D7GBRyu1il2XgivjVlhKgMn/flHlzK84kZF5Fk5Ifi5lLYKqL2gDwM3TeCQu2sfT
fFEolVemqs85XDzSr9nnR+IVEca6Z9bX9VYUrdp8McC5p+6k8rNwn54/R2YMq/2+
hWdqeU8rDFIy60hMPWdEoLQAHpqXTw88RLw5dfUNy1DVIQZxvUgQ449yQ0Gt8vf+
qv44Cfqqdww4uvnRAIYl7eFVfIiDlozZGhVELkN00qn48bg+JncZ84tVJnz9VXx8
gQqHnMBBlaCK0KJ2Wag7s45JAeqK5jgRHVXAH0brP22z76TRop13deQPyLKUSSN0
ymEN3dc5lM9V/oaU5qawVA8aZ8hgJ+waWR9iHI9+rU+tgG1LeMAhTU1dV8aJwcel
YTyfdWtg2Cy6Du23jXsoDiMBa9iFZRjqjjNsmhCfnKC4aQN0LxXoKn1JwDv/nDog
WJvV11qB+ocAwi3V+jvmpzI5k21Jc6gyGGfq+LH1TYaD8BtjxEN2zUcZaZmLawES
KclhPZl8kivWpnkY4fR2YBeqg3S1jQpGN+QLPaWR+QGrS0FuEhgdIc6fMGrGnnKz
Q3OTFXY8Cm4n5WIQYxj8rqXxlIeZTzxU38GrFv3gh+/quJYMJvXWxo7M2vtM55ko
xBxMWjqrfHwHtf0bszdx0F5S7QflqpOSYURKY515pmSBUfbkAGnn+TKRzd5nM6f7
5VEHWUsCexDF10wTjEEyT8hnFtVFSLhafp59IsH1U/+LTjpV+76MGCNaLVJ+mbe7
+zBsTnAr4bYRhbli33CDC6rrzyWwkEtK4d36E0LuuCiqM3hn2ZJPypL8FQSvVwjI
oNBUqe1TC9YZD4jjRPH7iyaSHZ9KZ5EluRxNSX1xgBqFtjDwx958aEWxfiHwlY/O
0w/5FNaO8hG1okv71UtqPPYn+5wwYl2DUFZ4GT2wws1bTU0BMffqEUZXFFnrHqxT
Dqc9Dxgz9/kOqWNegHiY5zgEkzQAHV04vwBEfBk2nzIOT1keVegmXgz/BriOgfFl
5pvtdGXKWnLgpFSg2rMRgruZr1P6A9I3Gm0F1S+3MrZR7Ip7VR582LrJ4XMOWOJo
yf7n23z+R5KmgvTD3jkLviq9xfFadvOxYr7ZVJUTzUADOykbe4r4ikEpzNHsHHTJ
5KJA7mzAWj0H4mSm6ZAftfMHdVDWzUkcrU3xSi8OrACV/kMpxfSVfQDuj7ns04OJ
slxGopjShd32XgiYavzeVS/XztxSlZ2qU8Rkyjpudn2qBRXaq+/RSDn+dCdHt4yr
ir8Azly3cj7urGvFpgUYyTYWxgVdAoTmM4I94d3tVxAf8qv7k3td9D90T7DAkJTF
aRQn3XQD4NbIVkGo0m6teFHUtrsdCbmt4+pUdg1sBjO51sCIBHf5Ew5MCNNosWPI
oT11LwIuqnt4zHj9Ty5kaNxlEPouHL9+kpidYw3HNhBDj5E3IwsbTLnehDs5bMx3
GRVHSuhgypbWNFn3cpln1qKMTyKUw3zNBAMiir87ua9aDSCMpHdYJ7eRm2cR48C0
ZAxNK8BgTjUCmlrs86lTk6e3aWStvMdeDMNEr2VaXp0IHRAVXgS9qZJUswcChC9c
hY39ZEjYEQmSWIE+x/uscjaaww5CaI0RCBuPq/d+nVsyR7lKy2VFSNLZqAtdSsTD
aBquhWbS7qYer7Wj3WaciaEScZvTVU7/5MYRDlLW+tgXKXqrFiGoW6WV5sl7cPEV
8PexviVjDfz180kRJ68FeOKpWFvpOQxGIdOpglTMSjf90tnKhUXKBzh/uT3d23Gg
9A63e9X7tEHJmbqQnJvOo7aVgKcmGUqGkzyIGdpNge1KlSlMzt1pty4YKex8F9zo
gV/Dar11qVQTumyI5sc5gelXbEKIdvjms1v/qVt5eFOd6mdCnb8Q2qLYR5pdyTLl
0epj3ppVe+zAEMSwdCHPa9MOEKAHYXh+7wfPtwzZuxUtfa6LiKUjBrTBpkoaD6W9
sASMnrms8MURr3JK/Jqqck1TscQYQ0X3X/Eamo6PypKf7AKBpUMaPORzfZ+VnHaE
OTIMBP0ejfOxm35y7qMy6RYdggCbRaquq21640oodY5HdT2BFQoRZtdMgHdsxAh/
Kv8s+H/xBJe2kO1VVjjCEd5Xt3f6gFmxTzVREiRUy/6dE3MRuA68R9phUCS4YN0+
v/toQ26n2j8+MRdCX1jYrMqumFjxDALZfcXk2iXQjn2mDpcuq40KQocOkx7pmqor
9IN4Lz07B0CKAyv8QuJgR11K7QBbUVT0zSCRjX1pIGhMEVGNLuIIHLEscp3oVRu5
8EBieM6mmNnTM63UVBoBdSqUT5r9BkK2HYlOUvR7A7yAlj8YMk5h0uxwv3nYdzR6
YximE690MRXJStLnpjGX8YPHt1jhAA0nuQ6ZkaoR2z0LXGJmmknKV9UXmGtB8Nmi
E1kEXNQckcdHCnxNMU+BdGaCZobnvaOXMMPPLyJZzjgeJqrKqWU3xxDeC6A72IMB
T2AkpVspMnIprbHc5cD1RmzC7iBFKxwynZnys5Lq7rcMjrA1vPrmm4tb5i1ASljl
xWUTQcuoGMGOE/VYbOxIUMg1vS9zHWlyBxgLPN2hxXmhX+SA2CXaNPzuIqZd87+W
NiQY5KZonZ+ilb6DubNtNkkxpUXGZorVQ5oWOh4UU8RZjj1q1b6Y9Y8VnV/HaObJ
Xfeh9xWvJtu2IOFzpjodfW+OJ2Uh7EjfwW3gA3oVYUEQzbj/HnZTvbx90dHSrCBm
PLPqM5nGDu9ZAbBPVpUDJVUwijV7vnpL8k9lJtDlFUoUTs5ANjGvexLELK5++TaU
qp3AN13WIhlpG2oQrjAKKKrWYiHqL1KjFUznznivW2S3OmXfdGgwqElolAOECl9p
0FPiKjOKq6DYJlfq5RROe/s0zhQVxmUeh/9xEnBm2tzVyP95BY7+tpV+zJ3xDlY2
0rL8U+OZqqLGvvyH7e48v1/Whsjr3k1Itg9yYmbuQl/LZ3xsAVMgEVFU83A1SOfB
NCSEQVNo77RJgQv2K2ij4vF5q+sn5zsLfgvv4/4yTIClBmkIsD3P7XpeUwrV/qFm
JG4dbXX09nQ7bMbYbXGAX0+neqRPc8ghTuZRUy6+rAbl1nV4OgCkn74NX6xvSpQ8
EdqkGj82lthMl/oVVImFWwdhyyYXIqldg222oGYvn0g5+99v4jIqgHGPHl/n8kXj
HImkYVhtrlY+JGKjz8HryNcwkmm0K/iLyuD9DjxVcxY7ogZJ9+zDFkesWgemjLFR
FbikVYoW9FsCu8ECTuc17Dva+waY7ZnO55EHhmFseZhEacAZ2ECDsVVedYjCfDpa
XEBjesc3b9EBPEPBwRrQCVGWnzauSVHvivaoJOl7SoPufXiSRZPpoELY9PegiLva
5AlhNS0VIIFxK43dNMSEQzf0yfEIMRVhy+TE6Cc3dXgIDLXt1oXD1LPXxZHWVX3c
zcjj1ZzOX5s7Vj+2oHRtzEFh0WOB8fOwpRJGDjvTXPcTbW0pI/gd0P8B+/hd/kMT
8pfnVh3gLhgkFDodtONR+OIZhAP+jIhS+mrZVkq2jcHbShLMM7n9HPlLeUOAXvcf
xEiVDEPC0qM6MnUBZi/i6Pl8ndfMkDCWxmMxPcu0dchNSaHFRGYOb0BT2G1mFfWR
L4SWFmlfMWEGUXLeM+Y4RJ8+g3bn97VASS+ZdNnaIuO3J8o0cSMogruROX4vi1G/
42ic0i5ChnrKTVHL0GhZuWE5M4K09Ya/94g4H1eGtPvjhVZcb3nzug2r7qYCxRnl
UoEwHJxW4+F6nco/Uul5sq5MwgH2PclZ9HmXW8KivqoKHhA+dqr0xAXNIyKqRig1
9ONx2SmA+9LjgLmlpUt1qgmTczGOyvC+hYzM0ryZT8GQAAAuqE8muBnU+er61W3P
FDXN399omhyZE1c5joOjEdLZknEDaOdih1pBtam35dPqhon6gxm151Fb5nahdF25
UBvnPHtUkTaxQb/QIsrxknxZSVwtdyHwevK1VJDjF3pgNoKv7JgmthsnzewHjM+P
JyKKLmMHNn47H89d+AXBDSyEm230siVTWGJ6m3VLfM0emqREggHQetgUd8NLQgct
Phxz+VFuKsPjzCnJebC15fvmmuByjcxH2SswZ8fK9BpH1Zoz9R74SpLveSzpaq/6
WJoUwXUv/efIC0sK7g9EfFdnb8ZuNx1Ovf9hKYVpyeIrPzWWMgdkQR1qK0g6ClFD
gdnyq3OoWqL1E8itb4LquC+9tpq7+CIDIIIkza8fclZXJRxfudmNcRiaepCD/Vln
oxM6TCsHY3rXGS3MoTaGuuw94X1yYPCudIudSj9kbt4ykcMr6RXs9REQNN0SqM1a
F9riytKJxUvQJfcB4ulIR+27/CIq9vqJOynpaP9IllBaJ+ZhscxuRS6+UDGr081e
HwXOU3U0UgW/V2MSCpqlhMQBgNeoPiJmTCPp+hfsWyN+icEmnLweOUoKLhwV9I9s
oD/4RQ3k2EtPyONJQbXCTngvMcutnDnGt32sdIHzLhhdd28+hGvKSdQkPnYuF+iz
/4a6qP7/8QvPa+HZzDOAPDyH4E4s5lSYacokTx6T6P3ijV13QuuxbuuZq+0pQmjf
FQdMKtkcMplH1p2OYtxUHe5I7EGUiRxYATCkrDTEWCnTDXV2R5SEkTzupU7FJH42
aGM56Hk1BYWrxaQYc9TyRjqKptwRZ+NjRI/wDUiATN+YTGQOkOfZYsX+JW6ZYDOS
Dt0Un+79QTmXdQSgdlEcxvuXbFtp5QtVUxjtnZnI3N51bUnDzQj8lwITWGB82mHU
6tEewvwocrhrhf7r73v/BICfWTEW4UaTyBPVeytobz/mJSHoZHOp8Yuph1j7ugfX
5IHpWIdiR/z5zIZDtWCajY5WtkdPsooa0//tnS0MSx9amOnJqE90mmnvr961csCk
36rJwTSQWWfjdShuT1PEGHdIAmn3Z9weQ5tg6NAgMCag11/CapkGRQxC6fOa8iCK
Qhcshfo2eAYnFH76unW2C/FGDqqxcH9Y+cITaF7IDEWiwXAM0JEEKZvjmySYDLMD
MV+Jq1hf8IdzJIpFRkoI41mMeV+UHL8QVOZAGSJ0UIIGLwdfCkjrkiOJgSnBfw69
nRXuVpZC2m//Wm4dilDm/9zshZw/68bCbjAeOz9eIm2SpqOsXHD1GxRX9FKlEUSm
RHw1iDKlXYWZ58sl7aJ+z52NfOxJJ5SkPViH0zW0DUJp+h1KaZuG4L2+peDTFuiV
F5cN1VPQ+2jZDLNl67MsBw8d2bUeuixvYbWksYSvsSfWITnySApXWKXegNf0sghy
jSjzOalde2myJHoPaJeNcaQVlo35BvJ8RNM1JHMap+ogcCCrUakFN8MU5Ws8/J5v
dYXYowqGBGtyacgFzPFKvfmZhJ+yl2GeV356gec6LYPcKi9d7KwE+VkX4fFL3V25
9oQbThpGxtnHAaOrIeQX8x71/eu0lLHFqm8IyF/QCfw2acbvZfQ17rirIijKSJTv
qLUywYUGM8c8sBmT1d7RfzzgYMglcr2cDpa6VFepWJgW36KwKUefZGsYsE6YIX4V
kL5issCglXCYFWVSMzScRog6QnnNP1y4beX/N0JD4EydrWFM3Lj1QyaNaVuP6dcb
+TbEEIK3RUJ8gQHifXfaNQioriS++dhAcSnRuzK2VrSlhz+IkMi3B+BqiwHGC+4p
fN/qJYikIsRVTpg3aZ21LVmLG+pPO9BijQuVx3q0aulJ3NYbkNrA8qjrHGtwR/J6
NQoibPPvm18PNWlBRlUtKaU98lOoBPle7h8CQazzCMNodiRspSB15qZnQpOYDBjT
LtBo2qwVj8wP9ZJ5oQr85wlVuGb7+fOGZaqFXwQKVBMaFN8DqK2qtIs920UVVvcr
sy3HHs1YcNzwwfsKC++7YbXLWWkmMy9/Ap0JQNbkUCSl7lRPlO+nEQZqITmqHG3I
mCSmoGC9THsv33PIME13DvwccpzS1QOwSmvXp5IUtmFGJgEq5Qw9aDgPZnj7mIdG
8/b7eUiHkMFT88lEI7FqgYpD1q4i3PFBpXc7gGxcSRtUpZm+1G6G6NMSHd2U5Lrl
GapeotMw/eDo7k+8zFK4QcCTOL1z6ypuby8ERdeXwmlYauMlQ6RGu8SPlhIyIL4a
dbNYjUrdvKoTPeyuvaxKMPoErCNo2m55dr7ngr6ud9APN+IKdJeaPjJY0bjIjb0F
8PIJsKa6cFJvB3LLYmdUWxp8pBb0vimfKgERX29nJVU7bogORdU7gDT+awKfdUo/
KfCKZJ7cXDjHzpCQqqbxbWYB5Oe5DyMhELVUo4tsVM1kkr5Quf7rvsMNjweY94ge
pPoawldmnwGxkJ1KfDr4vNuAGDCkKXOUt80vqDf1Tk8dXoioSlCD0zmX577tdl3j
1YHmuMwi2dbVa6rhGDXspvNkNI5KPrqdfTWChtBIvHJIryWinszHKWwPK765/jQB
75ndVUhIDAWCqajwGFXDy2DUv/8u4bwxj9uyomuY3mNT2gaXXZ/makVkS9ucSE1i
X748R7QF82XOwiOjmNT3ujvdtriNzmPmKn8e+EyMGnSH5KvuwvjAxd+Vzy45tqGB
11gVJdbFO8RsMimcaDeUzWgjV6wcxQ+IVZnr5Bj/RK7W1Zv4K8brgeNXv/DoU9uv
Ml/4hwxNAx5/aYg2y7Gjsh/CMtP7qhSjtbYPAjL4jbMgT5W5zjLMRWA+vy+qzz1S
7CvMmmR3rGNDHgw8+KBwJPHwA2ajWXR4Rxl5VwyFeUOu6dDx1hvi5P+DnR7ibtcX
cKpdCfFJ0+FQX2aq0YzZZsKB17nRttzy5ly6c0s6XNvp0Pw0fu83RPqmRnTlkFRe
20qvZwHQIBCaL5f6IlFq4ECIr7tONd6pfgJlcB1HMpBMEc/T3qERr47kXDSMM0fq
ynqusXe+kAno2uupXWOpdMRbpNtmZyp+l23I6XfVQyOHhsXRCzis/Wc0CDt4qN1s
yrg2oOX9zYeyXn2rnnK9MHLfXbDH1TA+XD5QQMHC0nOdjGcDTTAMFTIAeFXLecM0
KEe60XNqWuf7JUbre19soUwQH5HfIzyGermaj7ftsqM1cpeJfL3FgHeJ0dTKrNOO
SsOhwQ//Nrb4cHzCEemt2GKf0qHXn8J27L2GenYnhJea3M3yy/LRXnKEP1CFHdzV
lYVsHna7Jg5gdmwtKRGh/De5MtOSTtexvondo4pP5x4TwQQ/o9lLB8ZglBn00IMY
AxCzQpunPI7OXUDs64PyirDYomPRO1PeRCvkEEPlQnKTtjTuSURz4Dvf7wVORGJn
e814KZ70e3LAuRa7pX+RvbZR0Mk4keT0HzvYJMQO3n3T8ph4ZTuCI/5J7O5pTitF
8174rHSfX3Ja0twBRqg/wa463T0rHTqN4S3aNraHP2ENGwUeAFAJRc/4gr6+9gmM
UpPaTTTHZTaLNzgJjzKFQEzXdggOJlHSqMSGiR7xukPrE2HE717CN3cvJ9cnt/fl
TvC40ueY52mbXkTz1rtVs46lKTZMmMiDk/79cxgzCjkraQX+iurzKVoOj/DXlo2Q
GTW2y4coO8NWoH4W3GZMJGS9VsQAPzRjRBv00il4mHkpv47aVbzD63idBlgfD7UT
dR0vf6l3heHPnufijKi2HMsQVh1DwZTNLO56za4FMP4uTcKVhnmiFLGV5VeTTWlZ
lI0QfP2W1egGnTpnCI5S4cGgk17Fas/VVkYtuoO9b5q7RlZ2ONoKvXcnBKacleCV
ppqLMdj0lFvzF/vMEKOZST4usn3TJXjFIhJsxhS2NYGuSEUtFM20IzHLGIpRcURd
30oartXI570VuORSScYNKmXxbKUyMEDenN23MOGHkC7g1ZyvMx5bCHXthDrtFOI3
Xg3c6izEv7QeJVrGLPUXcyfJ5vueC6ll8I/DYAlVHkVLObOHahSXTrkJky/eMdQ/
sVCc6IMX9Jjgj7Nq7Cd1u0UdP3HDmW4K2Hi4bWCa0TgLhFLdBL5Hg+jjejJ0d8VG
NDb94kF+SxUQHPQV/iIXfX3R9W0ea3aJlPwXYcjUE9Pi+yatqH45gbX+38b4s6Ru
TUKnnQ3VeXCGuesksP64n1nDFhDLN7WlVLKZj1hnjNXe/lA4HTulpoOmuB1XFwL3
Wj8EYK/76+ha5tHnaY3Jf++F4eOIEScFWfZ4ae2c5iiYrBKmVy+avrn9NBpqVL/h
DXq+BzcYDrgFPUwPXZnWgtgONdrOuMsLTiHt9yZPZou93pJ0GpzvI27z/Yyolvxl
xdDY1ieCSKHs5Vy7M/2ywoCvZMl0XiO8zZoSWDjgRjNVYDT59NRZmmuNJ+/VnWux
yiQQJPXmJy8wsss9clRdWjWYAD5zxOkDhhAqf8hCdB/D4kBQ+YFX6X1aR4UGHwTB
8XgLZSno57E+2JEVzreaELLVGJAOXs3iGsqYT3ShkgUOn2jcTv7LCt52cj3EwY0h
Vwts39eFcZQDohxiWghHTk5C4bA/x+eTBNwY+frTyWB6Us+EBCYp34c3TGQ2J8WA
ykxY13Fuu451XIAW0k4GQsvBsO8H6A/iNAswSVQCwVBS623e/pQgDj+wihV6F2jP
viPBYbx7SsymO80uvgNxlIEzQQ9rLbLl/ENdLeduk7/F+Jn43WR6ep9lPB03VIKd
3YR4ExZI1zXW4Fl2CAoB6TJlT6oy4ZtlIQC2Ca44NQ0BGldYQ+MFiMKXPHBCyQoV
EtY+yvv6tmaWVF+Baq7MKkMFwWJIdvoipp8kd2zexAO728OOeiGVC/O27WHk7cB0
kO200O1cxxXo0AUSoWpzph/Xn1JsmY9ibhdQRAvi+8UmJ4J4MXaEtOXfnB/7AxXH
aQ0Fy3Wm7sQKvciqaCE2LqYGlbkXAjnGgM8YH+A76LqByV4oDVFlIlhznbjs9Qk/
nrdjvgMAa/LvKWWITb5tgHshLzcZZe9zvfjA2VJ71O4wV8aTxrKwN7VanROTTS/6
H7yRw3fvO+hL4Geju44gOZW0DJ9Ysd4LK1ked0k7hS+xL1elhguLag5l5fpHsgkh
uYmjBcskL5LWN069oxWHjNGBZ1CsK355jQXffmO4LLWpFjvEEvdJk7Ppmar/mIKD
P57RsaQwCuKOJu3W3jXyKvYqnhJyX4ZNs09H7cPc6/iYxcsaluLfYxJdkRVz23E8
pULtPiVdJeOPC53eLIhCuEhbzzslahszhAlXiEVkPNVjLc7pJ4fjhH3yEUZWIUrh
bHzKSinBbAsAkcKRCfCkJweuWKEmKzPcNowh36S13o8hMhrAIYt0mwovS8KcUYg0
p6mwNr5FqyJeEigfUgSpR+2DQKv8adyRxefk3sUCAxbuHMHJPd2WeAnZ17GneLZM
9gya0iRDfyXG7qcgW78snbW3ldFJZXScb+ck+p3lV5xHDAIXg7MpXFfKaYdhXnLo
HqkUZCyLcAQSvIw7tljNoYLaCwn/PQFd/ilYVwar+LdsCiVPoW4uiY9Xzx1kTS4f
mx7mSZMUPva77U965PIgIMBeKpjDsiilsQgO+fZm2Z6HLpv/s9WuRF8xckp4cqXc
t5+hR9u8pVSvz8TKuxRv3F9R3ozsag2QG2VYKY1DFSxRA5o/o1wWWcZCAvBqbAHT
XJadpWDeqJZNDzioa5IEhYLjcvTXjzyLHuNfq8A34zUMEZZID/yb9lZOebpdFRCb
WT9c1IkOp7wNpQR/kjBY76YAKQuwmZLHs7tMSPkhRl/eg4ci5qYbwL+/bKiThOzq
UCuIVZuopNR958DxJFpQKdbH+9l/YtqzPlLRPUJ9unjnzAvsp+fSPCJ2fWYnbPde
WFL2JlP45HVEau9aX5OfVsP1C26AKTdNd+oYwtDGqTacUM0LD66E7yz6L9sP1TFI
S3Us/EIngXEWtCEMb+U6XM+wwF4fawE2eoJmE69OS9MIJNxk9O3RPlFvnMWsBdr1
4L9JjuKC3iqiE2qnKRy6TIW1GOshYviJsB3DB/2gpVrWseMgcjzUXvHENakhy+z5
rnNO0jKOHuU4/jESv2VPX1K2ig0C1k3yGhSD3FBLy7v2dINaaIUGzh2F7Gxp/BOQ
eINWHUaRFlELySxTKKP2hyh9M3p0a7YIpFdEDh03lMVJzjH5aOLKE9PHBcz/TWR8
s/eVwu5me8/xGXcj5wmlDcuJqcNjw97A8NzpEVZ8GQuI31yTWKZrn8FfE4m5KDQp
rK0b+ja6uguspf6Nn8Ivv0troA9IzCr1X5ruvDD5sB3PE4tx9p52ZlXzPIuRrVXm
oQsO5Ddcu16R1CFtHBWqpACnOAVcF6i1s0G2kvoO6Q/4LvYhIz++F2zggvUmS+3K
xntRJrZSri2EJ3lG7gmCiiQCH6rv+RRkVx0vnXFp8YCkxqJqLBw+lD54JJWzSTR2
743yaWiMlhQq7aruPy7uUNpTW/iqheO3MKjiRQWPQL3+IDjdyXRs5llXCBfoWIum
Hw4WG/8rwYWPPIWNlfnhZIDBLi3S/6rMybvlQ2qlgwcSy7UwAKcv2tVHbaty82Aj
4MmjkkmLlW8LjI6nWZ1LmI8Ir/cG2qEizHAjIHlbpq6lYIzs8LrN5d59AcH4FyIs
h+pL8DwD9pKjdyD8MUUvFvUrYA04TlD2Uooc9ilF7Fe/0kXMVQYcBugPO+3pk6Gb
slHVVUv1jo3PK8ybC+MtHQ+HFvwzvDn1eS3hH9gvM5QWhYc3bdbTQiHFqcYX/zKE
wbeRjcUYhsJY4XKftGpt23B4fmG9ko5yy3xMx3gVcJ4JqjF+j8qAZz4W5CZe5NsR
Cz5xRpj7rTg90rgveFDU8Yl7NCQVKCYxqES5GT4cpVTO82KKrR07Y+qAZYYfhj4z
3jEmjz3YlQ4f/gmePAzEM29o+LWJrEMn29y2+Hgw592zAo5UYJa+dX9CeXjB21DO
RJppFc15+IuL4J7fbq1w92eL5KObDJn0uAwTOPxsi197M/LanJydlkkrDmQEeKT5
rsS3yxjGITmVXx/f8O3oGOGmQOQ5p/TJ0pUR3CgGR9YP8kN0dIZwTFSxF5wrY+0W
l7PrykICO1K6MkDs4z1YNB9QSh1KNncy++tiwaquod30KLDnPe7NHALwg6XQAe8R
N6rVmCJ2OTLXeoqc4klXe7hNuapIKlZ4BlZoYGz9CGh879tJQvriV9AqbrhadLPv
YTPnnWRu7iSW0mCvsoF53gAA1dT3Ry1O8k8y7/yJqF5ReTS/xB6q/dJ4K9PdkT7F
zgG6ZsKevv7vAZ8tCErL9Q2iT7R7QIs1Q9V4OfJ+lLiKP7jXgqlcIBJ/FQCPEb5u
WEZVp2L7S+Wdq7Q9+rydkhj7RnhyR2Iqyc5F6BGET6uQ8kKbQjYFBSVaMH53Jf8M
DLQAbW1IhlY0gruRzS4LKzkkT2NDqaOP4MC+IVtubx/Bh0xDlOTbP8rdi5lo0B/L
Wy2lrmTWFck6em5K8j5QqndX/O3Kn0wNEmW53abFJmWcQva1uU57x2zs6y3sMpD7
o5HIoiXcupoDDHZ2WtAa/QkEBPyWYYOf5HsrJY6MGbpIUiHdrU3pxQGMZ8smfTTq
IoITTG9QIhXga1+E8dHdB39ejib9iWyl4WUYF4C9kRpvcBNym/+2H7WTWKDXxTdl
zJh1YaxrA/Jk81tOonkgqTOzhzbBKv+Kvv0co1xvNfgyROj9AShLYugvCMzVYCtD
SUqRZUbsbK5qBOrZnVgNYY2oTa4ElwFzo4d/a6b+XKtk0f4YMoA+9wvmamEgbsEi
VVdaMzdi3OKgwGtlvXk14ntmlWD4u0R/OSbLKF+II30FG0XTRC+U2hUyNEbR8AVc
Bi/5AYmmIGXbfSd3PVq2hmKnlWRaXOYAPV8lZUIgt0Ir5zO/iEPgkclILO1Xl50c
vC3oXIMKd/NYe9GOumBZgFp6KySN2dJ1OK9M/cUsVxeVi7K9NvmQz8jU5vqGr70q
nVRLTD00wLBtirWmF4KrI9Jbe5OKazSTpQM0BtbPWA6T3MzWCpURlf3AoPJ/TebM
CLe1YErBXIlnqEvUSmpt5wJxEINc5sIPDPV0jFTNSnIQjjZvKmiJDEDXkpIUVmxp
05jrBdaLMv9L6EiheTI0R38cCudZsaOfShgzCKiUcRWpSJe/3Ccq7mYH1EnAsP2V
WAJqkD/JPtI2+lQYH3fqaISGgOxhGFUpsWTl7FsAEp/ayzZq2XVzi/PWxIjzhgkC
scMHSx9GoEIMpvgS9jf3mQfzKgtBbwohvqqFmRkToJrZ7aYo3Mp/yNaPFhBx9Fn7
kMebj8NeeDJssIMupL65Sb7v1w6aKi4OpAvVqsw29BbGNEisPH81QLgKO84WkqfN
BUQDsGV4uzyU76hQ4ac33cs0S99LIfnilTf7px5a5TOW9mBmfjrDTLgCMIgchjbR
1z84PNC1inYExoNu9JgKdXtmdSV4+JQLAECwi42PeVAiX+wF6/CZby5Lu6xuWUh0
VU7h30ujDYMUq+JUSZaKJp/ppRMx49dus38X9t2ZZKgl2l0Hb4Swo/7+OP/YFagb
oamo48q3Ehz6DzFfOVJqmC2JsxhmbjT2hl4mPg8DlIAQzU5H8l9ihBedkTul5nat
1cKwIuEkqf+JPu56Yt0pot8fDEtDhJuM3CxudX97vgsw6+mFK/7tpNwRl2ojKFRH
8D6Td/YCEJxfOKA2H8z8hQTG/C5vzMrq18Cgdy2vAj+YF1GCP0NIRnoLE5CHhBJ3
NC7Ey0es3LLWLYFf0iJxZ5KkaBVSi6DjnpjygiCvpOQd+vHVQJCl8MoxB1VUKupT
fRN/OBoejk0htbr3EVx5NJQyCrtnZkvs+VGK+QZLTuEUi5s8NqjdcRzEpesN35kw
aMqTKBEoBYuK3Nh90oNTZ16l0SHFtekRG3TcpAS+fJIdhms7QZiHpGNBVKPX8Bvp
Fw2oBYsZ/E4HlElefoRCSeb6m7mn7jwBDT4LTfza1601g+K50mNwAdeeS3exdAHq
IyJ8QPN7AqKZsBPgZZghLq81QSs8kX5Hf4G9/66Q0jdvSJTmpnkNMdBT5AwDo7O9
q14n3D+hrUJ2GbGcuTQbW+hpr8qZ/jn4H5IittSx+YoWJwN3i1gJsTqmnjNDmO6S
yZFEm4gHKmeXX9SYslYIsZROhUrS7SAex6SjEnexFSewkmuOVM0+eMD1oxvswjBv
uykYm7NsV2p7jegDJW0Vfn8isV+fW8oYxCFUv9sRWXwOjTUSU/oTXGL1Zj67SGU7
ToyiHvTD5v9tZ1puKuU3BBCUm5bkwW4QcwDvq6/LdFeCLuI4qVJ5WviJvrPQbkgE
75rBTVXes74u5FbQ77jQGOsaw9xuarODiG4UIZHlirMIDo21Qbdez1kJTxj90lvG
SeG3mCKRQQ0mUEo5qNsvjWj6oLwL/CEaOLuqANDCuQfrxrl1tl5zGOzgiOxVcvpf
hPj4aPCubq+n9E53exJ6lACOPyacmvcsTP/Or2cRDTB9feuIhkaFXbkcwz3Qp2DM
HebyggY51ZnvcWU55cB/0Wl8IKKOS486mrTGGRMbiYXcXHcbJIg+aVFTLl1UDi2R
q+AN62va9fx7dkCtpAgTIL/o1qNG4Vjxv9XbIab3buUrb/i8J//NBcp/phaxfnv9
irc5InjJx9P2UeKkPGw5CBHtvKM5b47J3lKeOIUg0DQGWgWOAfuyS4d0ieln5Pgc
WtcLuVzDCtIdEwMmC97thYf9XY/ABsFzZSzBytva9LyKHNqs85mh77msZWw7f4tw
n9MYvf3ql8m9Lv/GA88sKFHSTKtEmhH1rQEsxn6iugPLY/QQgjEBx0rTTdUV7a9H
PIiPGnQWGQRDNvT2dRnB3mM/II6xorJLoSscdnPAxlocRaON38+t26kw+2QDjyK5
x4exRIxsA/WO7sMVtR9hUsIcZY4/3svIO3XKq5eYgq9JZw6tfWBlul8Y4HSPGzy/
sLDUM8KBhHx2SH0gSqmFnHq/0+jTkm77Hd36n3HCgBayMWQuMZbfhOSrPBQkYcXD
D2S0El/pvXhPbR2jQoi00ceUxskC9rlYiJmZLmDIVFYrz2E7NaxPzEZR/sPjFzgl
JthS5PLqAELOQF5I3LHQR2OWboQppBLjE1UM9I9Xhc0nUWUFZmh4HSevN8OrIAFL
1HIcUWACQfoWNwbvvbTDre1TTJ1sOFYU/aGljo+wzhfH6EPGnKaoIGXrWaNbUmAh
WNlpcb9U0ENzdmTUIzKLHwcP7Csm5r77pew/Da8TB4WbKcrjGz6D6l1IF5HzEZug
cCDJhkUO/qtqveE3cO7I4qy4F+TQ5r/I1wkWLEZu/a4vn7QcsKvncddvVVh0iA2X
2fChUt7zUW74jbFHoypAwpwtGXLXDRokdqS+vJffv2B4IvEQp3PcYse0bFyiQFs3
+xkkZX99iZdzFew+7wNrsHUaOFpC0yQarem8C/rHOLcvDK/WjOWujE/RFKHQnGfQ
5cu1OS4NrbB49NuOE3rLTeVw042dFyq+YwQmlMpJ5xnZCoQucGvPCbOTbQCaS7kO
8wTW18E7yJA592T8O4znDjB2J5G23M8TjMmMuw13ngmrqFF3GXZINAvO51WuDX5E
WGdkN3TlYmY8LCR0Fm4dXhMBW0IjBva8K6pnfHZuIWsGUuFTzH577yKDRwMg2XtL
s6Q/3xMWtVdPO7hWwjSSGBnrbJxHG8Z5fj42VIjwU4mqwykTtmAzVZzgYFImzJwP
VjlZqBGERKvz9Q8+3ChIlKOS6NHGxwQumzBffgovsWbfeKqQ+x/Qhm4fHNC2mxXp
mDuMMzd6SSNkq19xRCYmRvyu0dy9ra+cLJZGk7LiKCHeUNVtq57JmaWkz5c47/iG
ZRcwzJdj1GJAhaQ6FmlYBkmybojh2/sWfYtfPHrDIKNM4ksCM2QgwX0Ba6tb64J8
cdoLKPYQ+IQ5Oq8KWybNQ3S6gLw3MkgJ0+3gW07ugZg7/zgc8aYOfpxSQrH/9LQc
OEAYHETxeGSFMbHlcnxIShoowVn2GPuM5mQ4KBVXTOxfOgdWoClzzDyA/9arxP3E
ASkXExAxWT8z5jWQ3gMlSmE0FjghAXqgynl6g0ZPww8TTy2Uz5w8UaA2sp1oe6Lf
KOvtVVRntMWH04uBp4XYvwiA8Sfzf+DLIwBI9KG6Tca0+0yYDXdcs1t4HjbRMpgV
otw5mgsYT3mxTROJBvt+oGnCFAXT1v2FlTzU12FVQEfeS5MFDmZbL2HdwWm+Z8YC
9w18D4NNYw0u5S6Ooz+CMOI6Kix2SdhRTtXio66zaQQgYDD3h9laCKTrqpMD8hO/
x3gDkg3mTZGhjUFFgcFF21/kAr1+9W6co5sSBsTlDf5bwCzqZap94sO7Bl5ZVjVO
MgLo+030jS1jQrZ7l08cBtXAVZEhckpaMURfX4tYe068DlzUBn1uD+LPNtTUfAkt
N3skX9cIjE0QivVoh1E2xb16F4XRJ1tfJh+CSjF4aioz0EZefMld3ySH8CsTUvGQ
fkmPNhRRYy+Kbgx4eOiqqjL0XsPkBpAZFv6DCpd4uWvI9a5q79prfIVVCPzBYiTm
Y5LC65E41MUO4wWDD0kf+ogrMU6+YV1tcI+Ji3pDOwAMyYkrVyYiGaLFdCIp+5jj
3zBi/i4Yli767zl+WyPaxXiPf6vaB6faeyDuOsOWsPOpYAIHyUuHZ+XIpiLjH+Js
5f5q85x8sMIhrFqGCB4xZQXB1WORhf0IpmJ96FSgnZAJYlNZ4vn3qDq9ni7aYAUu
UGxU+l41sY+IxUdaSM3wwbtN/ifbJW3lrwTir1i7aDvWRJ0fij5RNpBv19l6GXJq
N1GEnzmACTyYPOnSPtueppfW5fpy2x+VKETczdBfb7Xr6HOIxTQVmqhfhxSktEGg
dFABI274GGKdcj6sNgpgC3nl0h2OMJoxbpoMDr/EeIVCXboxipxPIxjfy32Yv3rE
azd6rhnP4XkEI6+oJFzK5oByk7SP2B4JJriCPg1SYZJoxzSK+jIp7jBU487xWPG/
ABBd9vXzfOBMbk/g7BGbQqXDBCAOuDm4L96zScvo1PvmhDdaRohp5Z3A++fgbfjE
yRHWjvoQVRdKDULq7EPwe6HH8WFD4LHjtlryNyaqvTN+lCmOCfzWWtWU+8/YYmB8
8MOqWzKLEbAifUJlsuwqaRlazB74qFKIqnREFrvqgdAbGddJlSGtc4tKgyTfpz59
BD8ojrgiuSxgjM9FQHre7KGeSx1tM+dZMG9lnVxHZtbbtj4lHFVO9tclkUFNbI7i
Lssofr2lXhDBDISf9zoMV1QIM6WRzYRU7tRyFm/KgS6pX8Imamzv+GByTWAPZJGj
ZVFZbsghA1Yj9OTCREMcw8oVgjmtVlTkFwu0VJFxewsxAC2qiflIBoZkweevfYA6
uGySoFK1exv8aYriBXCUsYIYjWx+F56pcaAaznnqseprB3mMTIXsyqCmv9tWMkR+
GEr/6uVojDNPzBx895pn3caeQFTJcGBokO6JyQn09DsnGDi8ef/x4N2nnpvAzxdD
6fcDvFtTKS8+hzbXuJ/2ymydGE8Zv/mLYS9yoJbzEg7qbzn2BB+DYBYOjbiGPsc8
z6uKWr4ZhwDLQFfBGGUXaz9+LNcCaDTugQGl/5bU4rguoFw4zm0g9vQjzciXEO/k
JCq9WNi1APFNBTMv/Ti/QIRDvMOe1GnMliaSENiZj3B8XGPg/XjW+f/eYqNi60T3
n6lRjLIQnPrz4hGq5f4zIXqKN70D/yDjJUdd3EtCYBKVPjMNRxbVUqgqJeRYOEI9
SK8VLwpxHPHSM4TVHg3MTz/wDqFBn9Nn57bzZJBfUK4LOOyT3nQcli0dGVEsZaaN
VqAoZWynZBZhm3voZ+gDqYTPb2svV3imRI3QMgMm8aZyXi/U74Ko29q8b4U4QjNL
Sc6NhYUq9UAM2cxQNQ73OkkdPxucH1iJKoI34gQ7rvHYqfHKp4XJRdzLYgljue9s
Fz3QpwC5nr8F1Zs7IP08oGjWycjb54vCnIM12JzHw4BrRgETZLyOi+PJaljGlxB1
LBbF2iws4mHQL5e1nvGC2Skb3AGpkSlimrhAk1hsdJ5/SFngmbxNPwdntHosAHk4
TNMPz1SGUyk7+3Unvy1JjHIbdS2HzJSbI6Ivd23JloJl17Rj6uTwnwS/c7B3CsP+
pjhLcjilp+htqJrt1Mwm+McccWE/v15/qWmOn4EQSm+gbdLx3iyVu7gfoMuJiEuU
PeQBOd7oxKCDhbo5s4OR87DPwqvDi4O1wron5EnltQdskV+7lthEAYQR+V5H11Ev
mkWNLUmGXcVV9nqz7K9XoeLFsl5/vcbPSgWyTyluKJ+Ukk7RdWiJ9H758W7vWONC
p6ydKGf7UQdwXkpM+bSDNbsMmTpgLeajDrEqzU3PrkR4iN8ndeuFuTRy7sG5b3ZH
J2XiMaKy2a9vXu9ST1uSW9s+toWDI0uWdEMWMAZN8SObNN+HEC1OUGbynpn8mWs9
HYWw8uQrSdoVphBnbP4P9XwEMHFTQYsLJ5QUk8I0lW6TX4pPXkBmdZWju1OI3FUl
Y+AZNTZpsyU/RjdCnM3auCxw2ZglKnSghED+qGubeGVBpdh9xDgQ/thmY8vyiUrk
aY75BiFaBM7TEDOr4p6LytOm83xUoFa0zLKYeAu5+584639yyjE2VvArQy3wnrs4
9YOipo41Zad3SFqwIv3BRbCxXPnewCb/BQND2h0Dm3zjzL8BCFgEhP6+5Fx1eckk
NYnrWzghl5v9qzO6B4vFL6GOowq+benUQkBk7JD4TxmUiKqrs/G5Lc3/hqLNemgT
4Y8DaUMJX08vwg0h6qSqwlgTAlQrP9zZy9/4c4v6jhXE8bVxTtBiRLXiKBebaVIp
1pMtoy+ClpBwrMt4WEYSqoo7YX+RFUAauT85jJewsc+OS+NC2lJS67E2deetxRvy
GL4eP6U6JeXyMU/DfqcTQ/660i23D/bi6YpluVna+8YRZYPYg6zy04jEnFCscM0+
eN1AtVzANj5nPyM89zWs1BPw/gMdyDehG7uxerqjte6HgvSG2YKoArqh1H4xBh18
kD93Sm90nB1Cxudml+GkJyl8CwmQTafdBnX9vAP1gtzcOEmjjIIIG6S+UEJhQNg7
7V8ShdTMadj1U4qIo0ZDaXeuyZsNm7yzGmTwSlaBptmWQ5dAoUo2mH7/Lc6yCJnY
iMWYwo2F+Ty6nBiufDiRje+9Hlk0eDEl9SkAlRJyZmelvilz74d07CctBUuQlA2u
Nd3PSqgMrTsDjwsr8diYylFol3Gfpv1I9X36N/zmdsOqLmKikydJuyOezLKTeZw0
EL+bfi1dTSX3SDWh8FkxjczgOGpPL6p3FKAhb7EZtR60zKiIyD9VqvlutntdLuRt
KA8AbxIj/tcPQhsXFB6jJ0gTmnXmMtETae+cj5YtXFepu/tqc24tGC4NC4tbROPS
es35a06m6v2/7zNjXhckrfmB3YJxzJzw/Hprt8cft1DHp9nFv/t+VZpuwWf7w/Gr
jP43+2hrjv7VbnSXPqZfbdRzCx6NredzHSICe9ed1lgXDIb1/slmIYbkd6iX8Alw
vovlb+PF4n67ayjV4yqCJUor74VV5bNmAicz+wU+E7rXpWNlrTIKWmChnzAwVFiO
OCrSSBOPPIVX4nfmgOdw86umpxXdZfQQKabHFjNDc6SscaZIryCG9Pf9fhoEO9XP
FpgWsogP+kOx+4y9jedtwT+4n9lsoIWGItyWyuQOXtj1SffHQCr4XP3APEAo+fKT
4uup+3pq5iqKC5ipy5H5RD3xrlE3Q9ldWl/90pDR1xAot+mHF3Y8R3qQBn+y9yd3
yoOIPRt2inijgZJsi3JKvn5SXhrFaGFlj6isT7f8HzBDrUEBtuNMzivICYm689Q3
SuQSmN2HSBplxwwm6M7idWRk1ytOiLG6in3H3BDN0OL9vCJMe91iAaXga2rPBCCo
BMFmcIbKsRlepRuxme1m6kL8GkZLL+dkJsu2Mv7Iv3WTZa4cxtoTygoc6CxmbDqC
D3kcu912vVtVPkBU03HRfQEIMSXDPdZ4SxHcaIpLt1OSJQba7i29doGJSavjcwUf
j+xX8zvitlhZMX4SEn9a8l0D2x8+8GWES1MMe5Vigu295YALJnGHeDF+F7MgNhfX
JcsIVTJN58TXA0il+nGxTACV4rlRepmuR3aUmBkgrVcCvvZh+ZaU1YGY6q6waHOP
J24BwnsumTi7vwl4HESBOQNqQKTMm7Ff46R4ZQF/1xOjq7J6c4drC/c48cx7V3sG
i3dj6mBs7aqcxT56QNoIPB/kKbnQAFIEIJx/9P2/bRND/M0pb1TVB9J++IIuFXAb
SUWAstUw2fxErIXzA7CVFPCrs5CW5WNQkN8BQ0KeJl8y8vbz1dc4d5WOVOMDDxAh
U4qUkP1VsVy8U8YSkYOLegpW40N4Lf2WPNpP6vyD5WG0mYq2+TFHZcKcfuOt5eyL
51TVE4vAcrqciOGdL2D+PlHHSXbELYPz7JKZbJ3/PIGV2Xxfxu4wWq5HpI/Rhppl
q7vaPISZ2nqjoM0l29VWy9sKZP8Vx5vOEU4KJSLMRabgz4GtEyRh9xvMXzOPAlQ+
Z4nQUT++klrQ1W+S/97Njy6n5TQMe1JZCXyc7gkbUHfr7AOL5ppYnmRN601rvY5a
SzhmmHTGXe9dgwiYSf/dvoq1JI54pN1y9YmONtMf/SPaWZeYT46z1NHe8P6i/jvY
g2S8U/joBWbhptkkrjH72fWu1E9haKYsmSgXEyQKbFme7AUqcsFHa4WwmFdki3Ci
XmuEPyS3V1ntg83foPojAqUsQs/GY0CrBryHjYYMP+FHfVupyWiNkg9DkTJYdD12
v4Dv3thVvwblTXaJehmPFD5QzFyeAe1wpGNQ0GgvxJTW8nS5WYMtpuptEGEID2TS
UsDzJvtnXfxEqxWfcBEirEjefExEQkUnmM13VuTt2oBubJ+uR9rNMcekpiwyUV26
TtfVTTPixY2bvjv6ZlS8cqo4LIvnGH6gAjYgTFBOKg2kQVEyl80wSXzFTkX+Hqe9
7xbqvvxqD2XBWKHESOI0BZHoALIju1s45mcp4ZE63XDNvcqaEH8oxGxwYlp3jrOO
sS2JSoK9mGz7+3ieKfCZPz1JopzvuJEHITJ1WbPAqDIc8W7hWXjufkwjgtQgWhgj
JFMK4c5O+AmowmT7qFn1lRLRT9U/eB50AiaMT4F0ioJ8pLNOyAkssOcgAUDTv2bV
0kVA+xmKZ1oa0ukC4kR8u2M4RyYlYP3eB/6sAonjGUjVZzz/xnSsdO92Wkq0btz+
h0zol41/q0bUFS6BgUk+HDHIX9QmZ5qL3xL5OF76QZcyuqKV3B3euXt1+hyzL6Ev
zCYGfnC/RvEzi6OOHlRu9DGISHP72GGzn1jNTTZpV5Sh9bgEk4NiEBWJpKxZMulR
KGpJ6cgCO+RbgEdHHQ8KyDaa/Zmt4u7UC2WZr66CySBGJRGJxBtATwUp3yJaIZzD
8PBs4GwXevilkEfetyZfnpGd6d/gq36876LTcUimFyamWl8iRElNBpRbaE3Rq4X5
/6HXoZRuwyI7egtqetfhePvz7m3G6M7lXAnzZOdlxYla17G7Sl/g/2dHGioXxqj6
jPZq99byf0VKFIIEeIIkheWq1pBhEK4FlBF4NdaHYls/lubtK0mZ9L2PSPTkNkhr
Nenl2k1J12napZ5tG/dhJt4f5R1cLGKcD9jXx/KpOEjqwYmqwZbmZFOXIocG+mN1
mgOMxakepJmXt6Mb+QVqllSjwoJqwcOs0rO1wiOCrw5qSRWGIGyY/ADXnF6SF/Zd
g1KvBykuAazPVmqVBc/i1ez6edOk/Ir8CDmVQi31L2jvJ7vJ70rIbxcG2l1T7/C4
9e4RQOUMB/AbG4dp5K902qdENh0wQ9n3t7rEo9N/DC+cJQjudkMUlGiqVVYHSo7+
URs7ziyiZ8seRCSOapDc+qUivhcOJKEGIcuyG6dgv5ri46auYPapjWJgrafmIuq8
npoKqg6+dSoMVR8/ezrETpsuxzOXvg7e2ycCMqOqgbJLSaeQjFJqStKwN45Bgwvc
0obK/4nlIE4eE+X2zsHtlXM5AMy0/Kzb3fcy6bvSII58NB9wiIhI/BfXICCwSUBX
Owd8NksHq6iUtz23wNQPeJwO3MfEqTqfzz2jwflG30gs4pMOepyDp9nAP6jBlZqV
dSobCPdNvuw4RHQVulih4/v5bqgR+GSifd8N/V9qr21odBZYndbZHd+fmCW+pbgX
WYXH0Fdwu9e2aRya/lwK4mMwIlZFcXHeemzH5wG6Ee1U9L6qOZmYRDs89amXXodw
V9CRus2qvNF4tGN8uCeIt/zzMK9vUC098H3e7ZV75X606w7/OO+39LBZz+xgZo+A
fXhq2UhxfWOMyOljeCLcAGQZoa80LWtYzY2B8N18sEKXS9DeJaWLu1Ksmws2cuh+
CeegiL/Imse/OKKaSy1CnNLBkLsB1SnPu97Qsw0piMznQT+5vkAtXnDy87MjQgxo
wOpLEmgvTxRlUbbn7kj5/3qxyNFzZ9sxJvLht/rwIlDdWw+LR8Q3vdKL4g3LPEy7
/BWw09N9pYpcHAlcPz3soyT+5vcatqKh3MoK49YyDnR4R8IVqJOO2EmQ2dE99RRJ
fuj+rPfgvLD2xUc4OumBi2U5W40VfkSQXm1+f0KaA2wyMRlZw+o3HyOm6Nqp9yFN
lp+MtYMzEi8Vnnzrgao175Ufe5SrZUItjUWenRQfQc+wVBIerWa6j6lh07/dG9R+
7EsJSEj8iTkZtqsn5RjHtuXdJ46wXftfLVYBuXqF1c3BYDsNFmBxosoiTuTexC6f
0Z8RDhApwt+Mx25mcSRejDteuAKVsgaOnq7LjTwQrvhWgmycAP09F80Bc8+S1tzZ
h9IV6M/aym2eO7NLsHS64NZI8z6aoJZG0YZRMm4BYkH6CSGKIvWDPb5omnmvOtMq
WYY1kjx4E/HBXhOuD2izvDoVvd1+0JHrysG4ESavYM1ArT2zVULzbR5uXkj3bzbJ
rZBwgizteDiaRrO7JdGHne4KqXF5hNmBme4G8jv2a9bA4IiKfN71BIX8tLj19h2U
VB72i9md2kQU8n9A3lCSySKEvSvWK7kBFaoUiOGNRrRASPYv872cdZldEHWuFNZB
a7xHAtCkekUcPt1JpVmB58685jTedBudeJWzkKnoy6+ooNJ+81KQ/uoBZ9ZoOgAF
wAd9n0rFSUpIr34evfhtcZeGw0IOuwuZHym3reUF5PZoDmnBD9aeDWeu1Qk9v7GB
GTjlMgDUY9lerBDdD/5QyBvPmcoH3xeV88z569oVGDeteSc+f8GtJO0T3gjSESoM
8b/kChfQMIhytX5qiaarDnASfUWp7ngzcYboC0cBpMWBgdgEmeX2sMR999Ju0Hbo
o7XmT3zvfb88O27CcJBnWR1FFgUVC1oOXl1p3SAp2i78P+P1tHr/0YnavFLDR0go
vTsZZ4q1KdF1r+QT494Wlra3aYu+cEmB9hIeLXGnyaAsx5JjpEyl0D79ROhgpz1+
YkK5qw1GBi9iyb94gZvVEbNlBn4tBoodMJtA5yN1FhvlxsoAK3CV4YTyjp7pvMVA
ylw5TTp8jos7bWc+OIa1AzpJ/iKVUdDawt9E5BRwo2+cePTuopf89oPf/pT1/lyv
w2CMLZqP3MKYbgwOMZDWzVUOZjTOZRS0UZu5ADjjacGwId2gvg8sT3ULdygz+lyC
tYvRkIYRn/l1Akyr1cMElsZzewu4UGUUKYTZt/TM4PRWQ3g8qnNEOf5DV4PZBHjC
8Z0M/sZEmjH5uvdcp6vDxHaMXZi8OzdwzSa3Jo28gd1B9/7qdUa+vhaCsiClmhiu
j2cJ5WgdpndIrT8SLG8Sg0AnMzLNT0EzPTtHxyirbp0/eS9ruDI8kqfX+SYiw0SK
hFKP51I0xXeH6QFf8mOBFyuXyINyay5vbdujTINDixB4N5BrC6A6FHGuaSX+TRuc
Afs+ze/Oak1WDZFt4wH9a3GQ1MC2Iqmn5tPAn7x6QzDI1xaxbzwinmJUslHJuy8E
UcG2k11Od39MOxCiqiASw8UulsvTWULS/dwIpBn+q6YSTszMpEzZdp/WhY50GkLO
QXZYf1/6M3AAQQ0cBRKhx3xODDjaUrC8K7aQNvHIcX+jCrU9tIwSNKYCBlS5OU0L
akdYrs0MYb7t6+3DMm//PlYaEV/P8axjatbtSEfCc/CiOdahylRaEVkmK8y7NU0Y
umZRuzOsl26EC7xsWJI9b60M3PZthBjKY5x3buminFPwPkHHeL3U2+a65HiSQ4Tl
xB6IpXQAAPNBbW8dtbALoarQNrw8QAnH0Bmenh57EKejXxANTnRGVS9x69qa+45M
0yhPFxYL4v6MB7ON4Vswx4eSZngH6JQ1JiREMz4fVQlepLp4T+sH7bTL+llGcJA1
nUg1zLnwvaljtUBI9eRWXoWW5ppSVdzZW4kqzKT3TU+M58GOK0/kJbOWBZm7OUFw
rqKYRx83oZtBNS3NlW5YXCP6TVvCBAZIIwJuTtAoKDCxlmIv/QmTcstEYrBAZHGe
c+1uRpFTtdY4v0MGHWF4lPjvjyOChhDaN76EreX/u6GqpjdjgXv5EwoiQxvqdqH6
UvHjNEBoL4F/+7HcMS+3ARUSH+1fiZg9pa1Rb8BYk7WvGRooVOGKwjXCB/0jqizo
o/5ksL5G4K/vSTjXZCP6ECa3Y9wKwuO/+MzV8GfEBugV0l+ABnXZeBs5cxKqEnE1
ZGRiiUuHZdnE+YO8dyjfRU4R2hJNsyr/3Afo8ZIg1LLANj+3Md1gbdW3PjRqKBRj
UxgMtOcbr/56JCN7lOnS64bjyZyDJFdg88F8CtYGt3NE4+Bi6sIHVc6BLgU/oFEg
nbluLLZMCRnIL96QRFQ1Ep7eT+AdCgvO4GmybG0UXAAvUnNQKgS0RlrVIyGshvuS
7b/FEIk50DEIzF11O7rTE7HxmWKvCw4OhO9J4sN6Wivf+t++8xE0OdTHsrhfnyEZ
liorq7RbFigNHhZBpoKNEQmUe+bUH2DZACgHG0i5Z1Y/hgp7IKTlSoKYQIgc9gyk
jWx3Fysxs3YO+oSFD+ZCtGZIZ1+JeZHG8fyBnYyY+6hvM9OoTXbf3i1oeQforJdC
wpogm8fHNJuhoSQHOT6HgAHVFMF2NUcria7WfGestDyTgPUWtTurZZn8JLL7ePQ3
QYjQu1ULfd1nu6hZs7bQ0t1bMy9Fhwnky4nxSQcYNXmQ6xbf1T10n5A+cz5zJYRA
kb2WF31OX6neU6q1FXUty4MgpJQ/zHlcNPNEAf5sEYQwcbelme8RoffamgQQQeim
Bq5HiU8WqqkyI4Xrce9MNFWv+nFJfctw6AefcGBBEbRVtyo4bNPDc+CoqJzx5Kyo
F7JhFsCVUi73fSA/NpDQOjDmZOxtuiJxvwM/1BAtBN4nqMPB5pESxpXmsPeH/jx2
gCcasV1WAyIghwhLIDg9383QraNiIf03d5heXT0rnMdgAxISRlnS8aTHKGEx5NGU
3g8/sMS5txdL5O/EcobVrSv3Cf+m6xsPsv6fSiG/Nw7ctuBBC0ak8cHpxqTcXhBg
xTUi5jGjTp6HIPqojrl8su79bFKbJ7e+5qzmhoQJCQ3cXQy6Cq3skfO7lnJtGzlf
rIl+snRd5Q0i6uioITpc3p3RSTHsRl1aF7iMz8fz/pHrt+WTv5rarUjDm1IrNglp
ArmAhooogGcwGhtRneHt/PRnbLm+wwa7IywRZVJqewLOsgYr4EHiBvY6RQZ8X1kb
GAPCC04PPKOSUmUlEAkiQ/QLLg6vCMNkAinAYKAWDsZl928ZrBt1kP8KWkqFZuUS
kdyZgAcyDWf6DCQ34u2YhmhirYtZrDVINmjB/oI5bV6uQnJhnV/NuuDAKRdBMxcL
l9Xq/cUGOTvYMhle+A1Q00Qcr3v6stA3Q+nPrd5kXMFZRu1fk4D0Y5xJ3SWC+Dc4
VQPW1Wmsxp5afN/J2mPhWZbAoH1FGurXhNkbnJ4ySRl3qEwp1fIfNi6+E6nQoxjH
OiZcAjjGU45vIO3fxFd//p4Jly33KXSS4Wk1XIL//W3eR4j/Cc986Fk4nMqk7dbe
RsA7ESAiSV2nAiPfa5SG97gwsczBT97H0FYoTn3/M4e9NWxi68HAsYi1r6m7IceH
YrN1QyhNL3eMALMbM6In7ApGB9fYwGYLsEpP3L68sx8AYtuqdb/i31hIpdJyXyp/
Aa4x3NQ1JqyGGuJ8NpP2WlZk3x+uD7o1KxlA041cCXaZsHG1nE2hStx+tTEKfrQ9
16eEFoxch7NAivrPT4JSAdjQcRO/yVoM6dD73txAVPfHzlGp38i3OZ4fO0u0sI1P
4Aj9CBQ2OI3GthLQb6Pc5IAfYUqtgEl16fQg+fAakTIqsMtfp694cplnrvwd7UCe
dPymdIKg4SoqFoPKIB1Cv3h4jSkQ3ycDXcsbNywA72blaosblKlK7UoKU1sk9NqW
rn2EEOSeJXkChk8NHp7oG/Sj+bMHkuaoC6AVNpevEYWOpE+3QFgJ5FxZdfEEG/DC
zCH3pDqHcyw2S/VPrgoQ8YUiT92z+QQLMgUakJjvVMT94g6GEp54w5yjbQkeY8vK
7rmhNo79gpfiFyNoiJl9VmoCrLF7YosnBcgih2vBH7p++hootVy6pLQ0zVOrn3nv
USpm5h00YYDZv0alvOb7maAWv43R8mI61w/p9Uz/+R+m8cGvdJd/JJKKd7lXp3Ed
OgWI6RglwAiuxUZ6RET0cRMURV1x8qzzsdfVqPAsW4zJ4TL++zRnDcYGdpDrTReo
AAecEN3nA97ycgPW2c38OLtuPxKQ7FRBnhb5AhXD0kIkbz/jKWM3WZxsg1wYu1gc
aeh1yY6n+MGikc6Wuux3ORpTDaDsvClNBZAfAQHcCgCXOxqCktiTLYfzusm/2TNU
uQ4UZfqsAcEkb2VUqWHBhmWNnViKTOTslnGSH22eaut9w/h+wz5cIFtGc6VXg3g8
RUgwNykQVj26kvdn6F5YcO3Xd8+L+dcS6cR3WMtFAOIckzGcn7hjWkZMGRKQx7x0
a7oaX65BQExOxgGN9Hok/oHxvoRqVZz9nvt9P6lh5VkevJ5Ms61heEC2/aN0JhGz
1i1tHpt2POuFcBAB4anED2js/p/vFwsKDjCMVmWGXJZz4ThTtWK/nFY+2xeKSVe1
25umIKgU0QNMuQZyBAFvaQXz2eW+M8tOipGzbwhaDjoQwbDX7zkHUI8IGuA8FpU2
KpDIGSsA3YFCTeUzjCZJTfDvEsdrTxBxYU2ZqnHdSFb9mof4bzY3zHUtFCwNoBfH
61hQOVKTex07wLjLEEcYvsOa0MPZz/8+Mcn4XGELyZzofOv2dE3xKGhAHmH17Ipu
nuV7pXsov/femJyolrp/WWur3xU02NXf3Ryq9gcqQwWECXpttMRDtMr2byf9XdSo
90IQ2PUc3eUKA9C5w6jHhab/PXnnKtNpteSPjYCQwYunqPN6E/rnWWZE8eaK+6VM
vlQ3WlFixHJ7dLXTNCANXiwhxOGBQWAgvHf8WXL9WsYZzNjsKzbaIfWZpqrNtPLo
TfGiI0gEMtb0Bm/7M7zDWZ4ULBNeX8m4gT2jjFzGM57Ud6jfLGCSg2tyy2TxPPrm
i48sZMXpwmBKHKtt/nyYReON13K5RVRZern9FMpSWGz0BItkgvYqpyP2C0NOUmda
To+sNSUh+a+xrj8a5Zp49/Qpy5bpHEcGxZ5X++Y6jpFNelOOdNYlhM1adquDl0+v
oCMVdC1rjaRIkxqFVtV6H7dVd+KQsoosTgY67/NwQoIfDLMCI0j/pCHas/Zr4xMK
d4dJUmIc7JPNhxuuDzK4kyJypi/Xsj4KzBtZQO/KyiEY2ajNDHB6zi8AwoMgeF6Q
iKL1xP7IVNc7mIHM40xJv48u562X5WwN8AF+JvpInApdIR0A4DETrcuOMHrIgYWi
oQ9MMYV9tOc5txOClC8Kaql24EHTeLa1ybnbOTuizu5QfDb709PC3oYrG7zfTMWm
PAaZOn8CcxGFDPcNW1B0HPJvuuacjtYYf3irqzBWEBfUxUKHe1age/TEtNpHwnSn
bieKsZwSlsvno8q3G00fXWDIMT2mzpu1ug5RSQtKHkBAsNuYgvVu9dP9HXqnmZj4
Ugnz5/bqVD1yD7zT12kb/A6hJR6LECAYm6WPeon5gaDV4+TyCjTbt688WhnTGirq
Ka+Dgw6WCnJ+ZcYSBsvsckLpYZUoy41z0utmDu5ExjVUsGaNQLCGmRORXNcuohxO
DRvMEYKxpvL5R9sqtBmVPHKTcioKr1qFGBwTQ3iw1gcBpexLa4z0DbvXCyBJ0fIm
DOVIzEvFhOebq9ykCxlaRFPL20OXztHm2Y8dv3x9es3MshAuN9DNhdZGkydpPdHT
zxJrNsZfWBb5vYdA4Y/02VCJVzrkY4YEtzv7z+EVQSOIpGb7D7SIt4EeJfasfo2g
BPoHFestDOs/oYHEhRLba9aC2qYF0RabnLWiD+hLaoy9uSjWx5XlXTbjdP3cGpMY
ErXvzFDw96jiaxLNEqbKNo6WmTu4ROvuXw1mbe63PyOXXuzupCFf6+oFQRzI2HA8
jrbGZ0bIi6mQeOE+4tSaZKv7/DVPCnJFUmbYsTKKN9nM2WrFfbRj+wPbMJFVYyBR
kIwWJxyLK0ftJ36zYEtCdNmH+E2CrDXP4Bsu2wHTbTU7Q9suspv3oNQLOj3NPDlv
7q13rjHo/+3zzBbYS/BmuuLBEjERfMsv/Tn1foACSxMfkuh1jhoeE73dSyZP5IJ3
RVwTyduhWW14Ih6KIXlX2+eZ6/6ch/LpE2FqBHSQvoKCjy91yOQ+RKRrLiwr6Pkt
+kZyFXLrlv6bFyiOBYBwcGuOyX1siHFrji3a/8xR4YkDUoBonaaCjXGYwpD4yOPA
0Yr2tIxFCWSA3AVizGMxy8rdfrlat94pshwos2gltwvU8Pv5PeTBsnpIunxFBEqs
vQlZCbSRCfW0lZ47dadN43n6VxzKsLPma7v45CDIB2F9bKBXm8JLuOZGva6DMMqh
Ok1aiGxNPWSH08qHBrmflGk+TUe5sLkZzeDT3AXt10iOGGGXwczNYj7Prea11O80
0rGOCUloWhJ16r21wZ3MlHdAWZWo8zU5NUkGQJFv8WE2kGfaSTSSTRw6gBHplebi
3aqztLjCOafFfsCBEd/ewbBPC0FPq/Iirol1bPNWshnuDnVFzlkGNqn+KHUjBNxq
H49R+pM1ce5wfKqtm6aV5bAPI94T21zps1r5KfCPfQLNBDbc63VKeUImoDnsOePH
3vNwhedC3hIBJQSjtSrCpK+TL7oRSwucrPubnprz6CutUHImLErkU8Ijoum2x3Qt
aWowpir6QdX8Sq0GlPxlb0+jf2iPRDCgw1U7FzjhMs8jLfZdXa6PHE8DnyKR5a88
HKXNHE+8mTiS6vQaNu+KUcy+HYTChS4kZhvAoeR1zS4ZIs1INEbEHNMtJny5cJcB
oNRJr4YM2j7rAYXzPkIm96diyuurbLGam7tjgBjZFhZ7Ql2tz5HGhwXSzN7FPJtA
uoOASRW1ngeOX1ab+UUfclJ1PNerturX0p4aNrAuhoZGbvTYx1k2vzKA/RO80kfv
eH1ASz+Dp3NGMwZjOeq+Gl6ZHJJGl8IT/ucT1oQLms2vLqyIrdRG+Il3hZEkHj2k
JhwCmZgwdJjOa8XLsE2NPisL1BJHS+f8kuzKEVaJtclv/sON9WbhMrfqmf0iT4s2
jTAXGUVs6IylLPufJx2wLpGacemnBjksZtAFhcl2j5devZz/DKmY6zb1ZyXutLKK
7qK48ilK5N8kN5pG+ihSX55TYyL/DXrbLhDmMHQKjwZWdGLbFHmrxkdhkLwRcYMb
gdymzqRuWnX9yfLpC/Mp9e33iREmfcj1t9yXYuF6IXKtk2e3iB8KP0S+2DeoEt6e
sWYJXWjH9DNVC6nR4OfNqhoEmto1queo+TJUuOJg1r1Ix6wUangjYY1xsF0cZDVg
lFpZYHS5p45iyimxWRvCKj4STu50WVIbt8ExgR3YcLMHYl5nVTPOFvycBKzgnOS7
S7J2EtuRXcGCcWh5Mg0b3pJI3pzTiMyfUpjIRRz+aNa7rjeHmAceEg7gxa+mpeUZ
6z7Oxe0a/OvyhW1G18ehQ9GF0uuJRvADUDyHelaNTmnnZN4j1qdWvsnh53IzZPe2
cHtKo/e1wqdQZMC8COmQyUJCq3eaRTDzQX+piKz+pn49mB+IQOb3aZmA1R373rhD
2bgN5hlY8tiyIu0DOV5TeiftUNCP0/YFPFb/IA7CGANNvTuj1T/vm5RQQzZ5UDMN
q57F+NxHuNRI0OhEkTZrfXiWeplIVknigHGPBYJMIM+faGaLcbpTwb6r28ossYQ2
JIrGqRH2Cg1126gb/Ya/mEf2q98DrEMEe7ZMCYNlSAN9HqRAOKJx9tdgeUXb7enx
mGs3sPIoAo1VBpSirp63AGI7seHaT9HjB7jXWBoDrP1NSE6IBib+sHBYUIB5lQeA
BBWKWCHjBjYwwAzRaurOwgKjmc+p7GU18id+bgzXuNJqOYOdqpRzo4QhZh9emoRx
um2E6t31uDwuYGkG+QlOydYpZgjL+9tR2yyPT2g693DUd6LPxZvwX3/RPKauoTa4
ChWuNWdyb3VmGpUJL7FIXIJ01j0x7lXTYV5ODzfN4PaY8hXiOSYDuK7ZcH8Vf3xL
QT2YaXq+YIflN/ek+Twmt439ekuD1ToyZGsWfk3OX6IvBJko40WRNrpCDpFfN8R8
sHI6VTSyZUbD9CwnyErJ9Wa3Ho36XiBTOF2R0tjNr5fpna54oNmAP3UAGUT6klM6
VAnVGN6stMdUIwsEhNKnjMT0tU8TEEaEjqF8/Yk1V37ux1Cuo/VBRoT+MSXp/kNv
q00+Ufrj7de5aREEkaqqZT/+HwnAe4CGQ7gmjx3pnZpHttmgF01t3FSWFY2MJLg6
qQjS2CzWG2a3b7JxG9r9C0cpZUkcJLT5itiT6pDLVx8c3a7R+Gjl5Gz/TwjY+22n
c3WxScOo60qWy8dCkCGTVbF2S+xdozbjsExRNRm4ggOofH36XHINnVRZF0En3gt5
2fpATdgXipD2BtCpeHO5MNUdmR7cmj4qJ5VYQ9p98CPoXvEXtXu6E7tr9wvlOcu5
K7bLXF4YjgNTKYU8L2M2h6wFyh9W7x9ysuhcAXGHQVIRDhoF19PzguutXSK7WSBz
nvu1fjgjClNATbeWX0XVm5ligNWpi+xpUIcmCqBehY1c4X0MkJyzPIZ2j9eoJ7nN
mPGdh+iBbaR7uYBde72qeQcI390QqpQ69o2ZzlLbRUO36NJYTTYp8L2AVQHL6Z3U
Y7/RkUcWJEFGDbOniNHPGOihdGhSD8zveiqJCoxRQT1Zc6CMGwOEBaURSe+J8p9P
mZ8i8W9MWC7iAQA5jpmGJxQ3INQQwaglIAxFml5ssQ/OhpNAVT4iik7AWykFvYks
D58iYoxfzYGZCi/MqPBMnGT9ZL7vVOPKL9Qb421+hGgb3e9HL7sfOCGinvj0+w+4
Q1kFm5Q6G2I0FNU97EXNxWQ3HMUGWwlC4kxLVFjAIro2KuZ1WqQmYWFujso31PCu
c5nlRawFIZo2Este8bScWQefcGICxRLVrPsUkg8VfE8rOQtYUCD9P3QDmZAxvza+
ACVtbFJ0kuZZttxoX5ziYSPkEQ7zvapbrHkHG+yE8+f2ynfrkzebkGot+dM0fxNG
3mBXYled6j6mh1m7BTzexSsMthnxnz9bK6A75UDsxYs8yw1AD8eXJvZ+knOhPyrg
hV9ie4nEhVd9RgaQuRjVrPyiHNP0UhxCjuMTttwCOWcC62tePSPpY4FcHS8Tw2el
ug6bJVhNgLJlNwvqfecufio/VjOZoc+tf9NArH7CUF7aBTNNFP5zvRMfPCBWE+E+
BOCuaGMRaY99fGxjl5LX/CHg0HSPz24Mm92KcuVMu1Y91OuWpPiYlGm+0noAO3ne
QfptCPImYFd4Ek/EhejNDm/KiJn0b+nlujda9cZRIRNhLtr0f0+oiJlkwHM6EHh9
uH4gfTrVB75yWOvnumNydqo5cjdNo5k8/4/VrOdPSRSZNvNmN8w2DvYKnWFdI3pi
qzJHoQO44/XibpO3/sQTXU8LidAv0P/6Y1H0iaNqvcd9b/X7KFqT/MDaU42hmUXC
RgTu8bipSxDTMpr0Qir7zX61Og5V6qcAyhnvTHkw/ItxoQwB1zh+RzCprIiWSrd7
FFiwyXRiTXCmvbz8ixskDE9oAREYPNR/VGPIIWgYOK85SYPs98ZnZkpTCXWS9LzU
Ho+ReoB4QjB05SBduI+53t7vSad7ZMNyE+i7Ad7ai2DSTjM/OTjM+PfnQjM31jxd
jGHHEWwEbb+eUqhQ4QnzGFV5/TkOZacmdjyueJUOCYAzK42qoIWFqA2p95nTh8RJ
SJjLG9FYAHQdP/4hyLd8ZX1ZCQI7/XPNxVdLPI9XmqfkFtFp/OjBojcFoHOoOuH1
aiYUWeFW0uyhS6VTShMjty56Fr7PDSU3vD/nFi66s+FTi703R8FiPnmm/e6BcI5v
yUzvdKLs3Oj+yNMGGPx+zJ3hN13nwPFKc5Dx7NEZvBBnHe/2jMsVDgsil+tJKcux
whKtfBs82wgGKr3LescPqu1JWfEIxc5ISBDey/rhd1oHun1oeO85CsW2tcxur4zL
pWTcj17F2UcPkfGH8egq0cN0aXq0aTn49e2uYqKQ779DmYTk0cpRQvxmUeGmfKQr
l3TtkX+tIb8QB6oQmc3trjyONsmmlYZ6oqz+TsddMRExstWp804snKP4B+INM1+p
PpMmFJvRMowTaTpPEIE2+gKIru7EnJzWzsQggrOvoA8RAyZQDgXj/dZZkSVYVCt6
yx6M4BKWNFggF9X2dPd/KLhVXfayiZtfyW030NJMnFqnHf81wjRZTNMbT8//GMfy
1zuUyrU3kNYFrXFrP8dbWCuLaGlsn+kaSQ/prtCcwEfRKSHxxcam4c3Jr0pnV8Wt
IIkcouqLEAlGtAZk+6MLKR3r4u/kzpQwyVNlYelywWSphmr+TzkOS3g1jFG2Sz8B
G9pZYuZktJpOTYG39sCEcEOX4TYek0ZV8R4Ltqi2jKFK9mVnGMwJYOv+AysWu2qd
KuZSEMqR19eiwd43rtC68v3RCB7EVy4aKL5Z6okbXyHnZOthJ+yvQsaeTAIETFMx
xACjY2Sle++CRmFqqz9s3OZE3XJX42avidzn3l/3UwMU3k7oTXh4Pj5RAooJ9O/S
mP4gcWzqrBzueOW4wvcYIkt7aeq+T6HU+UtnTMmpXJW90VnXpiJU8UAqappvu9Eh
iT2SBJQxhZtOU/M0QZvowB+3W26WyPUJ2nrizrpR+NhivYQ+eQ3RpVCCHduRtWP8
0Ed39bUMDubWdIIl7uXfJyv449Doh11AbeHbnPUavaffCorp18QNKOm35WKA0cOf
XfgfLzWiANVmV9GRN7Eajlx/ffm045ohJLKbJ+f7la7fymj0AMtPJ+PrYo5qRDgk
x6eICGcmFUd//untJdpXFJgsJ58EwweKP5BDc0Jw4NXUQn44r+f0I3GGLNXSquYL
KtHc+AeRtLzDXVnZk3ZMVb6Kl+ezJc1XKlq5aYYRN2gAhDu1Zq0CmKA6Y/rnbka/
dsPeL/MhyYx7IzudiA9Q2Z+fj45Lsilr4Atce+klXFJofCcb/sDQtScY9XSsWwRy
NI8Cla0uEsuY9A49DuRU01LGQuLx3D/deCFbhC4HILJ4hTKRRHs0DL2ZFOb8QKin
ZQ2mc/FID+PIrT2zFncGFyEF2CY78gpqoXzf4RGvlTzwNnKFpS8bWjBhO45poQ8E
8XTSVPo8UqeGOb22YR+W2mxTh3BdsZ4bGKvcag0ePGJL83BSmabVwDyjpsqJaQKQ
OGok0PqQA3d/qj98bnh4sq0km7eKbNdxQ8v45gm/5bU0t8zVNtnBaA5+GJRC27Px
KrA7Lpesy0nueBO1yjlCTSD86l1YJ9BGBk5TGEAvY/4+ATeha2nhbCCgSiHfhDDr
0YQtZLpYlJScmFcq7hMxDQlGhfztPHUeHv+cvN+HLsUNFzerzkfFMuQnOV6Fyomm
nd4Yaw01nHQvpABoWXxwJj3/Sm6b2XRJjvK7eJdCeDubI+WzRz9U67M4V0djx6BB
B/pUGlHnml7quxjrpMn9mAaevtJhA/pR80BhbSsUDHLUTnfzM161X9JD5/Cwov/P
CBBk+fnRrBTNcfVQDd0/rEAf67KzTkrsKjqny2RO08YuT01IJp4myqy++Bn5Ti+4
IfJx61avBcfJVSNQvc7nyJ17xaZgOUxbcx3tezF5ngvzyOH5PKKFCy/at/vU1lru
8WKZhV3KN2XrZA4acXoxO75qS9KTHfg2wZoOK7hXqfZ3/yI/rjvEyACx2cRrKtw+
HkaVJ9TpG1zcYvdZnV3C8BntuFcuDnsdkm/lPeDV4pv+FZyvvfFizs1Z/OJ2VPlx
1kCyhWn0hrhqVxS2QO1sllEcmPbqYIDxtVU9H7QbArA7WGTThP1HJbyH2LfH4QA5
Zx+1/qZOxmubyhwBCeXmOWIIKFc0A6S28Vc0zITNWktGyKbdLrnOkk3J2GJuw+/D
UFH3f+z3AQO6KP4+tym8cE+HSNRZiUf9ge6r68xQQHF1/FJ2r/yXRX8MRlt1q23q
lBqNcU6jOVMbyGKKJH33SrhNBS/NESDybr8eCeC7N8tfSEgGXj81IC0OokB0DNgn
CyfyGDNz+tMtDB+5/AEWskI1Y9aCV7M2FFQWZhPrnTTZil25lSORFwgR0Q3hs4K6
SK+Lu40pFd2irNjWGYQq/a4AJRL9Rx+nhXm082VbLR9gyDBS3sYgF9bm0JMRdEMk
599/SrJfZj9oq+czz6/KnME+lo3LaEAa7t3wCtunowVUq7HkMix3aM29C7toTLfL
iu8tosKNXd5zN8w4uKqbMWcjCsWzQZcJc4ov2QML965+yHHyD7I0EUxYfKTPLQ76
ceTgYlRFJYf+VT0SM2x86sG0nPeckvUdkWodIGZydR7hZcBEGHnedKvGO6xI/CFm
YEpp5Pf8xWcUDKr8yZ+7M53EM4jQgutH8rpG6fZhGMjiWUtwgDh7t8RPNmiQjR/n
3XG7t6XVJoMuvOGg7Fu/km6lANXPg8LdfA3wJaYf0At1NlqWyO7Wu/oBIwgJKHEN
gTiMIiuejHRVGtWRfX4TafjXoDuD0SNMW2w1g/XHzJCHfvFvBbTIiUESQ8UyiSKU
k/2E7ftW4WfVndoHnSmYHQMth1yqwhVMOIH5WHdqNm8KqK70KNyBtDycmHsbCvwo
NMCMX9s+tKQuSgKK+Xzj2Dt5hBahozvx1i3s0nKTSMuWXxVaWlKUpMLngPslBc39
36cBhhkoERDcuGlacFIFsk0JVK3knUB0GEDRrlstZeQ9i7z4ZULuYPFP787vFRjw
PjozLZ1uyyO4cfUBkBkRT/EAj6jaxmw7bgh9jg35OezCA7KvrYAbm9RAHdSIAhCz
cn03zdVZA4tGdynHM6GJVjWsO8yv6J7M6LLeb1k9mzx1wVWYpGuqCQACW2JuMsmj
SmIRgjzuwx7DYWhrG6wIDK0D4VXzTqiwWdM7fP4Q4lw79/X4UEaOpWD1aVOzi+NU
G4tihKvNssGp/zUliIVkUp7QTgH4RKwiVk5Yprqbfyu3G8/xns/LwSfgI8J9XbWy
MSQVfshOIYCdHDlGf28AgkrG9DgPY9ctBnGAQLiTcoP5SAMbb3a5q6LDJHQ9jPwp
vshpETJ+w/RNEeCyEc3IrLArEVt7jDrHqp+ndFm8DLs3cOBX+GqYSDnTCufNAkBD
+EFSSIe3ErbGLzALgQ2dwiNYYQE4wGlBUnwyikSjxdghVNL1XPv9ELWRubuMiO+z
bmZOniHMycuPedPJM9GL8YGbdFjs144ejHSq0p0q/EXUTlSb9FYNT1B5i1uhIr05
4lYOQcRD7Vgi+AUyTcYCTAn/i+chA/jUj3zU4VsRq2qWVFbrjWvAd1VMO2bH/hXS
tQnG1Js3Tj8Eki3P4qER42aMNOSGuUBPdkf1SEZIigMy6PHPwDy3EQ+9afc2vc8b
2Pmwk3yscMaiEuH76Yv130PN/NgTbGDkqs6jwPWKPsVfeXHammmwjm3b0kdxxMel
J58pwY+eOt0kgF8NpR5TEn45fPU78q2W7f+wwgGe9naqmBdhCYlXnW5z+0AtI29Z
BJxo4OHCUjUx2aXU1GBn3aqOKrBgcvFSntHi0HzdK/WOv1L60UDgu7BMHCIF5w7Z
pddMHeQ0FCzHg/w+E1yPns0t+r0nTzaKIy5JPYR+vV3SSvVPNLjvtSJ2jM5d28xj
X/wD4ZW80vvnLUCa2HgA/7RkgeCYML6fhWQr4wNT3Gd1TtHyukUlpJip5VlwbChl
NZlDsH9LQVxuWbuYAjtL8f3hTGc/u/kB9fDeYCHtfbnQITnayHrnb82mwXuv+S+v
mO2mBqEspDY83eYgJ9quQ14hr8eb7IcBZbh4NlGxKLcBXb1PWpofLv0hYNrEGmy2
OsnQd9on4+gYkLpb0tUJXUOgVvbkyzHMAle3QM7qm66MiKNWxhpsGtGtU/wHmofp
AZ9zlH0+uZuQjJkqAI8KlyGZwfh6uSLRcsfRCKRyFDLuMJoR9uf2qJFTUXk4QN5a
0gp44t3FlaOOzbvxrI6ZOgXkvpBxn9vsketM8D3DUjndUwk28ifysQ0UQ/VZKC40
5B3Lxsm+Yg8jHB1zDamseK7QZyuDPiyR9oScI7S0ij4XEdWALQSW36x/dk4u7lj9
3uLd8GVyhjzqDANWU0zec0tIUO7H2VImSI0LIP9iFFrAI2eZPMsWDSW+jFH43W0a
3WRKNXLLww0yRHiiXh6inT4+FRe3nYRK5tJpFhfITGGXuPipYW5nckeE5nQj3sM+
D/RWp9DzeUwRlsTkLcooMGa8glc7ineFGiARwF1N8aKbKij2Dds77Wc3LM8JRdDS
gU4PP5lmWVglKOUi7LjJWpXAqBXG13E7XiKJoACiovmg5nt0bH34hx+85FGrCciy
1MVyXAIyIte1GAliEVn7Jrr/2siHVziJyChMhUK4FSwQwLTHhCm6FGYKE0A/QJ4W
u3/dim837BOweOjWLxdvcW7CsnX2GTQPwjyHTTy3xlP9I2V1StCHtcg3N9M5hHMS
Ehg6ephWCwRfttV3ntXmDjOgMkHzAubLNNBxZQhvfkdSNkdv+JtEdP9DkneyiJep
S+FhuiCYGYVObd1V22397tFbln+cRf7t1XEzPJo7kw7Rl4ndzy5Y2SNhPfE7Ozz+
benoa1QKnHLBK4i0r81Lz17zcs4ezmgq+cGjllsC2lJ7sU5EEFTr+kQCcdYNlzzV
UgLeOVKeTxu1S2VlzGPGKbH/0uPoeMApv9qH2vdKhNtppiQwWoTou7c0f+iJHuL6
Lfn2DODHvwdNFkToonGDbXz7mo/B8xvHriyAgVQ8FWggalnScxYlufzctH/aurw+
HFE/z/22w4G4fg+QzfK0TbPD3WIhlvw3qYpcW9xCEz+OJUbLOAVrX/PWIrePBtpq
Fg+md+fRvsAw4DAHTYEpYz79Q5ibvz3O871mfDqJUR3tzxu6F+W+ve5IWD/PW3z8
tpHbtz8TuG2XMb3I5hoG5GAv3F2uyMnqzRDiN8t9wQPTAAAqWVYQHV7e/QOh3/ER
HBqmhyaZoHZzamNDyMdes8p3roVfzjP3LDpIHAMgABmpPHYlcAUDH0XL+nr3nqFQ
UOOzGclZZ6HXCx/KPnnUXeOdgE7D5y7KrL4YLdo9PgvQZUvHBjwbjUaJy2FFU3pe
/oizXCFKa+BJX06HpyjqwxgNViemGYnv6ezl2hAfDiF7Pg9/FunXqOwGQpqW4KYY
itz0l3BW6QghimS13SVVdhNRXUkamUR99da1fXdhxRHux3a3BeEAADrMs+/qYPrz
hE5CVg8nYCuvk70mE/fgz2thd5WGcnR+txhtXNc16g0xRgBJ4gWxHYfDuxjdJ96O
CphlEAjfvHoePnr2ng5AgFjrQSSnTsjB0lCyL+RnZtDFNmJE/qO+0SYvSlygMmQb
kwbmWT93fZ7D6OmNbdJJSQWQOE6WUl4iSDJVbOy9omb6SrOSLMxx2ynExAku+GSp
y8oAqvF+BcaWI8JbBsljbbxofQ+gK6qOHoOXM0EV//KslG6LIS5yHm1Mi2cxu7SH
p8T3AlmTPNABt3Y4Mc7B98N19QUakP8f2bhmFgxzYO3LmyUgpdZCPmEbQVWKuqHw
MNCMxj69ClEq9u2qHHb5A2dLRx7ztNX6stSpgH4VIVX6sX2gJetPXHPYETt4RVPb
hHhYs99an2h+ZRsnq2XL9j36dxOQBT33AQHIt6Vw0MRVIELX2i0dcMH4oVn4U65C
a7VHgIL00pAAlWzgig/FePV+A0I6zDPRQGx8hHLc3m7IyESNkcNwxODPARhs/rXp
v81trXK+WYVgYISMZpdEfoHG/3HhYquty9J39kEICQcnM8SkjxjilanGPVACpWSf
A+5IzMqNCyh6IKtryUWSP9bP1NaKmQtuKF0ObcuBkXojwTGlLAJ797nEU5P/Hin+
uJg15Pd7fQc7ZZX3mDmsB+IUrtt/BsRv75dct5rD6K+Wnw1WQ7+kLi9EAgUAdS7L
SS5+OcYYR1uyw4EEJmDGijhdmakK5ugMXHnJ60b+5i1Trv3spM1WFIeZ+/7IUyfx
4MFSVnsVsZnggo6fglXmAS1wZr9SGkcrJUMWw5k848WhaMQ8iK3ZpQ+tMd02EDja
ds5D/V3A1im26zOLsCf6mZ56ZHldSkVPGYQDNIiaqTOI2nCdf1dQKyr4auI1Obhm
Ztt5mq7EKUk/WPsHWCs0sygQYK0o0CvzFUqY9GIfAiCBa0a603n6LxKgS8g4PgDh
oOSacn612mXHAkfkreWfLvJBxtZpEmZNYkJu2dweWYQuoZDF0NQcuAQDEcKMa68v
V8CVCywTslFODolON2Nl5avsy7JKig3CdBqnf6CG4rOsAsbbXWlG0ZwMb/iXH5oT
nUjDcDPYeTyezpUv1yJWTizRkJwr3RJxNrGgX0CY/7SI7Bq5+9l2WBje2ai3PUSb
/tm1to8OkJfJW6isLZFvIltuHcLxGEWR7PBnVH0DBYk4kTk/D5hxzg6c82WqeugR
XkpK3D7zh/TleXrXrj/e4Z7UeT3l+MnhPFLNbx0nRlFsQaTC345tqWmUY7HeTfH9
Pd9zEsljN2W/xDh/GD5bboJLTKCrcFgMUOld/I1X2LoI7EC9zsZDrVYpx4CRgfd7
K3f9ONbF7EGVgWmDotEb2da3KwEPUlPpuUYxkRCfVLa5/2flkz1Te0/mLpve70az
TYRjemRBjg+q9J3n5iZTEVzsGEJBYnpNsfFsTVUWCKkXW7MlMjQBoJ0PXgCZYB79
MywSangtC4TXsotUKD2+8g2WhBQbSVhMB8UGNmZJkPaULFVA8sgje/iKvwH3dgal
YAS44UcmTDl1timEq8R/xxL33KY0Xwh7EtAD0mhpmFfctLYvsGdjWHGpF1e+Xti1
pFeQqjj2rJsnBi5MHpbCpRJtKWWgN1NJ5ttEEp3slieg9ugAcm7Tl1JB0R8IFIuT
bbHfeA2M7VHpoGk771UsHT3X47lbSFbExoOAFT6IvLhcG+I98gToiIZZF7i5lQm+
yozYuKttpIIEMDAiBtzdAzuTmnmU2Sda1wSPQelPMUXxxA5lKH0fsaHl4rSKDlaL
9tC1AiETiurz/t2DglDHBJzbkarPdprP7trwMuyC5V3ARbapPkccHLp1NDalnWOY
oR3HAxCh1qfUQVm8oquJh2yHVT2An4VjKPjP25BkhiJklvrcAYZTY0pj9VvNVd4u
6gIwcgV+I1g7x8M29bPA9f6jEDjN2hJWZ6vySvDXullhvMz/Fr4/4eDWHT6T6J+U
zUFNv2JQr3yi51ciwYEmR31JI11kPRQ6FSPfWGZPW82qy0kLqRwfM141MQ7kIVwL
DQVICgNpqPN6e/ldTC/mZkBJoGhSP7JByHJYcUV96e0jSgnmgzY/wVUL5GfkDIVv
rYKgdgQLk1AAmCqiZGoCkaRobuS/vxXf54XsYONSmPY6sexKnV8OdwY1RDzkV085
E0edTg93DjtC6KTN9CmO5IF1nxhPm/q9hym7la9ZNquH2Lm9Wj6xHWndi7tKw+dN
5N7umaVgcPKSHMPWOKyvXMQytSZzAF+SM7eyMQozaBI86twf2ikSmoWyZT37FmVz
HdSQO7FNW6bvbczx+lTwduEbI/aCteE/mQHFHux9nVraT8bY4FPZKggHrQLmhxJ0
f4w93Pn1y9vuasNGYg2Ta4ekE69HVz4LHVIC0yObBSVjUe4vZ5imsm3c6Vbs6I7e
MlZCwwTZyWSAQ7Fsuo1AAVuBtrUgqweWNv06qe9FiPyh/3Hb3ehiZqj4ed7DpOlN
17OEbi79YULFTzovtVEbIJXUqrs9dV/y5IbU6qs8Q3S/64LDppla0UXKkLLQ/jbl
xCsPVUuMZ32x4q43A7aoBZN8PV0qLYkoZ5gzDPprgdKxYffwvRHygd8th3jwE27C
ISUXL7F6E/Powd341iLIEkuzMYP6imtWbWoCLu11lqMUHMJIhRRFqyNePsu+ycyz
Qgimr4YFXWUwxByoO8jvzSccm2lcHec2zew05grE7PBw8H6anSilvlMON4mjQSiw
PA8qXBZK02pZi8eBL3FGzvuz83I5+dMheuFuUi/OBWijiMo8s15buY4BtpN29suo
xSm+6MFB3jyGr/n3salhqL7WwNsWhhnTzTMLW0tzdCm+q/mC9EG3YH8F639foqVR
dhGB712+xC9JT/aY8I5+ylRji7XkM58OA/ROp9ohL9wb+FLFcwp9TmJKU/0+lGUw
EDvx9S6dq6YOjqZe3BORZGrYgIFewHGhQ9UswCY8lP44Kkb31b/5DevE2ALJb0Ez
oWNqqIlMPJi5nZcBBRDlXaBZgmvrlChfTR3MwwXumB3np6P+wW3TAmINZdrTxAsS
rCg75HmrPhjb90dewH9tkr+tt86GaH7g4WKjJeE/BgtqtgqzrgxrzSFCT9flavss
my545h2GgTAqg2r+3LXaeQuIfgXHNQVP4XKIVxeoWTRwu1NGYFecTR/pcx3ZjFAJ
vurIwvf/8hGvP/sGbv/mBjr/mINNJlaQMrw0TAskxMXx5fB0JOSJKBfZnfJJRdAS
/D8B7Ig5zxjSSQ7GJbxFI6KL0W+Pg5s+5ojM3f3i8j7r76coAsdDIQBPmgH+Cbl8
2SVegGINon9ErMXL9AxstIJ3KHyNJWjYJiXlfNz3DdIvBR01VoEetAboK2dlhTlt
uJjN1IfBtcyAhcXfNETZw9f4o0HUl2hKX65aSvOEs7JOTiJGdJcQoSZ/0Ib1zCBg
C38fCZezzrJ6Nn/Nam81snecFjXOk4f/kmsWJrAuYcoQOpm0KgQrP8YhJ0e4z9ef
0meRDxRY9m8rq3bRbWmxvxt/gP43+SpYou+ZDZoPq2GSYGG6iUlpdBG+nCRL3E4R
z4sKX1aQ1uxpIHKj/VIfCBLuR/XwdRCspLv6wS5pUUrgk4jf1F+c5N+EWBcWkCUI
+G/EmpXCsqNxJVtkkviE8LsPHylsrbsiqbD92DDh7qOXrIsPA2r5byvLVciYR4aT
jLMN/lpGOhSDilNr4Wr4EE/9B9BRB2A3d93jgwbdtalJz5VQbj9lCt7wfle84/by
hsYrrv6LLYBUl2w7rcopfXQCy58W1NtqiNxODMHEJ6JuQgQKiIhHNEKN8RRV/srx
iQoPQ4vW7PFpd7PS00fl9/nP5uS1hMahHOIfXmbTAlG+tVYLY8Zq8wovnEbATnmT
+sVgwaBBbP40lIo4tYbFPAFC5MYBCN8LTVnbomoPC+1p4hpvHHEdaVrfk3fTzh0h
TrzlK8gVeYCvmg/s3eSA4XaUpldxlnKfEjA6Pr/U+kGAkkHvEfD0ZjWzSaX6+SUB
j01+DFicY+LfX1OfpbC2+hBjBVrSEp3Yf+MuTnH1nKQ2AW6CEWE9PFxr3lSUxrI8
apgk/xPz8J0SOol7yAj/qOt7kN81H13bIeZVs+U1675vD4hofUJYMsz8GIx3slr/
bF/7+SE5ayDp8s+sH5wKVhJQh8HfblmoG/ocbx8tFhtshRKN8r59Ne0d8Slf2F9M
kfSjKAEX8UNZg2dCu3qtAaIC/Ha9/JLcoo2wNaVRbx12rofnffJVslqhYyPir+q7
Jwwh3s/S51DMKd2adeO+piF0ISlFVIDRF1liUJ+i+rGwXwBmfL57Iwg/1uJKBi4N
1PvJtjW16L1VReX7taDTTtV4iV/kWlby8Z3fppZo5T2G1Ok1PDJ1n3kBRFZ+TK10
uF86OwmimNQHDyrX8aGeHcIvhdBizTPbZ5KO2tYqeJM6WjZ+i5uyC79e4CergwCa
Llpl7gtB0oLKK0VXOvPz72XO5j1FuCfay7tRg2zN7bg1sJaRi/o/sduSh1AkdZYZ
YgtY14ReXx+8GDr+ArHYk1OJwz2WIgKJxtZb659uNI4iuZ6T11G0eI5DhKn9Stt+
aSSVPS8AxqCsD7bcI5ZStqVeYiCNRGY87nOHzAHwCtqpVPavk3lLl2N0aC8ysb2T
O4y7G5u33ix2/L3eoJUjB1idbf0focMZyjHj8camkT/zYePOoJasdpOCXv0fFWuW
9zKFaC9mKn3eiqYFoIqnF5ySySOijFWMJ7O+RlJdkaQtr99+hkfpJule3svMFxWc
v8ntNOFTF6DGdTAf7glQwPeZFEXWuPve9sPOFZQ4GlWlJtUoWTVbw9PaAae5bpWT
DyoCANq1rZMGxn6l81NnxheRvJ/6OxGZFIuoT1QNVV/lWvmR3/hPU9bZn4MK7/Ti
DFH5eQ4JmyjJS4Q78YOEnXrMVDccxbZmxMZW0kyHurwUIcO0QYo0PvIi9AvVr0P0
Z1wIz9TcWR2aqFMC+oqtDc2ox2QGNqeLj3w5pTrr70ygIMFD9Jb9ohVfz1usX8dx
Nq5RcTuYNs+wOP07QzlEj9wjrlnpGpv5bInsIVUs1wHzzDSZFtZrIpJkMAoV8MwK
iZ+weWSRv+u5oN08Ugbm9pKMgDFYAZVvv4U5Ib6eIbBfbV8K6OTte89CfFHLemNU
XvEAt9RH/S/PkZ/v9MjxxcgwMhLzedHc6g5diEJk/gyj5YMoek3pZ9uhxzadf+aT
J4psnB+jPegq0spi1PllfCramqtFYH26tF6Hrk1NpW5hzYhtKugfrLrBvdc0b1ox
4vhB7WBE6e0BoI9QLCDV4HDaVY1nlQMI8lZ0hh73dlmcmqNOELNgRZoQMFLfFQHb
ZWfkn/Z3awh2Njx9TPw3ORvTmaCAs5nQAi0xFxsb/xoqhBftBnenVKGuMVlKiBKY
XtN6RwlAAl+ycbMi6YS7OEEBU8At92ZbIKdSABh6jCVET5SbzdeCXF+Hqdd3B6s6
ws72bjSeBPi6HNTgJ8lHgFJJ7dFzpdEMG2o8dZpwbzKVroeozdqJeebGZP2FAPzt
ghDpAV0KnSSXzKuI4BbNDVpeTp6as255adWeE7PIYkMydgGYsro0cDCIySoxyAR2
6RYFTKeje2R4OCnnIUwx6xM5vZ5AuWOzH+T73XuuFLjBeIrvTnMSMrEJcoph/gju
GIAtR7WOIAF3JGTrS/0qH6nAfRmOErYLQr03itHErrjN627AlEMH7yRdCbOVxlz0
k6YRAxgzT0Nc88I96Gu/nb3UuFVVUyiBLK1LOe4AeuKR8xzAYic3ZEhkVIofnCln
yscMCNBKnMKKQsJnz37Gc6m15ZP75owZ1k363T09RZgjnPH3zSuvLKg+pRFL5lmy
g05LD93ghzlhjyiWGuFpbZgLa4fUe3zbvAQGmTyEDKYQs03aRLalP87BtML0tl+z
iNqC85ANwywE+LVzU5WInbiHVholw2QLFzfLyEX7T9fbOFjPVdvDteZ6SP/m2I0u
5iabMYreAl9lG+AFbEM3JQqFErRGqbm1pdcOWAUzc767bHBcNufgOPFNS72UzahB
SSGN8suxdoLQHuSo+ta8oS05p3LYbG9joERVmtgBsyod6G6BdFNuxnu+x1ztYhFN
enPj3kr+H67LcjXIl8BQkchTT8QLdiy7EqbFg8sm+yScAvotApb0ZyOYfxTGpFci
zohqMjmTdRcmHTorjvLf/aXhjck6aqnn8i/QOv8YOER+zY8VVjI9d9Sf1FomRQ51
o5k+HgjmySBn1em3RyMIe1521oNLscZ/qX/Do1oj2an56iThRLywl4ZyehSV5uKr
mkR7ArKPCS4Ar/Dg9CDUvFGnB1zsfhLFZoBmhGQJt0zhsVb/wsxTBW0vo69LUnBA
EO2joklOzOQzym+wAz9L2Rd/3yN0Sgm4q5KSOdm/gKwx79Fo6uX1a/HQj+Jb+pCe
+muTzAuEp9z6ArDe6i+jJ2Q79OFEGjh072A9ea0RdPyWkAO0u4c6Ljwyfk1AqXiA
HN19xF8ylgo4SAawPn8yYphQWic0uGqT3Sonl97yK3TRdRU8/UdOaKCEJvNKJ048
BuHcxBViRtb65dEs1qvOZkZAVMTjpiOVIzPCl95KfL+v7FGUxvUoFBdJefMmfbMw
5DWf39t5Wdj7bkXyTK9LOewsJrMS1VwkqIzoLrZvlVFY1EBB7N6EJUng5/7zy3rI
DYqdI+H02qqyAMR9qGtGVRY8BHeNy5hBT0nL7e6i1dPXuRPVVYaTpOoaCTGjFR/X
xxWKel19Grwr5vypPRwQsjjTdwQ0bb5rqDyk5L3uSBjxklbeXpWEiGVCcgYFO5Ys
wV1rHyyfFjak1mb7pvcU8R3FuHWj6UlBqIyDZs/75E0j53pTVA9Isj5P78YoEB8Z
WdJoCe6vqGWOTHvwshS8an/c6cqvyWimqREt7CnpJh+asm1Wbl2H5KzH/IZaoa8h
HfmDe80oW5SK9IaOuw0sKyUCyl2UrXRQQ+jaNBPfW7Wxvte/k7m5Oy3NpSJ/TgUT
1ev+92m3PLFeFqEBdgmLunqKHYsuHsFMBqhcOyKmvnknbK9EAELgyBz3oZV0Dj0F
aicb0RokZinBe38gmAoF2iv+y+YZAKQ71IbZkeYGLyLiZAFQD1rs0PIT+e8/fTbE
2mInGEL2uhgHW09jDp8QrFciS2yeLDRrgROQRxM/27FULIKUQsn4pn69oGYV3frT
0Jk3GDHU3cZgRGi6saTnRp/VAbgfgvTwLS2DoWm6sjsqHuTnYkVNHvv1HdbqI6eB
zs2kP/Nko+yDshdAoJq1o0hrf54BvBbrbJtZkUixBoLCwJo2Mdva4mMUkoJfD5bu
+0eKX+kBZ/pPJZahYHlaZG31qvDNtVh5ojIg6xdmTRTTtLLqD3eLHl9VInff4j+Y
Y8n6cdlQQVQ8mweTsuvNEqk2qyTTm/vFUWdF/XlAJTSI2RStWTR0ViQFETJL55No
QcCpdKrjouP09HFI78t0425PnwCG4x525+lZIbzROcK0eI4WioY707RfIdInIPKL
8UrUoqMfaCEpXaLzxLHab2jXKMdX5WZ6E8FWcXfafl0t0JL/m0qKaC7i3QP93g+8
fjVKhSZnzfreV6Skh2ugeeUWvSh783ikJXwBGRdt3iPnx+5imHlxH41b2LJiEM/D
Mz9WpPMPYuGYexEm9rZervVk8OTi4pkjuMaGG0WggP/UMcqjlimVCpbW0SD6CzGm
Ey+wV46MIKGvskihzlWqVAq7IEzJky9enFiJ+GUdVQhDkDeE7tIVkVLMYyOtmghD
7OLzkcVj08BVSyeJxscILzqfZ0qVr4wEMRM/6vevLa57LJm5PZWp4h/oi6nF+NQv
Yk2wC+DPWooBMQGq7A8OV/5WNPBrx9jwot/0UQTKf6lm6dnUEPrLVp8celY9Smzw
HjLsVbCJAxDPVad6t9ytJVBxvbgnBLmdGQ2hgMl9KOYY/NwkX86lgwevi/HGALGo
Y0QJ11K5mS+AKaKGrsmXGJof0NalPAPLJdCiHyvF4DOlXycmP4QT5OvM6snGvpSe
eNkUl8c4XNBhPy5wUdFEiFNJRczR1Fq3LbjdHBQNLQEQUkUkfGx/TSXL66qcsqRt
TyYnxdyzeOe7nWqFUwKGfsaOlj4scXhS5dOGv7Gt/jQanzB8y+AndxyEEww6J+CC
bS39upRJ4seXo4vjagEsAxUjyhDzMssQMW/vg+wWfMBhJe0+U1MICT+G5Sx/mGrC
cXGVpLWJ5ObCo3XwRw54QsV2r6pm+ciF/+K+J6nx5RmslL0lz55VZQE1Drqd1Xy+
Um/iHLxvlKiPXCR2KqsVjwey+pQxSirSzDnz/c+PvOR6sRzEthXsZ+4a11UL33Id
k3vtyi/oKPVzz4nZfJfdquyxZHsM/6gJMWHvMC7ffhFkzIHD7+r0AQE3vHkQfXZo
ABPQVSRuKAaYM4SqI+ELpuI+/2MoPJsA40g7o3XS87k4DcQuxKGAbWpNzlOdAK7E
KElzPZdOjk37kBZYc5gSA+QopCZdpXQ9C+kD9ZzQGrjCwW7IGNtWvbGF3JDXFpiZ
bKrVb2YvkjEAORZgZp3dxrjtBRJHlpou92GpnigaNLtz2VllOtgr/9C5NZs2Qf2f
xFyPjH8n8b/r+U1uigvFrEcSMYscPQiEGn8BqqDT4r8GQprzx27KoRlOJqs0FPWm
QS3iPPYYz1ZW9ep59tk2f3SBdy+VgJP8TqYl0fNjIusITtCPE+a9P8IPDAhvUqJi
4IHPFWrwUR3pbRibgOHYHFx3XcVmD77BEkLKspbjja9sJ1czzABUfEKQR3Hl/Tpi
emhrB7h1XgYjOaVXdd05edtReYTUqZ06WWUvKakRhB51287wimHy5JGYQgdk3vXG
HKywhAXdrEhMOhMLiAJDj1VMf2Pqdp2xxnzkz3M3mjCodNdpD6G63/Ovch/Xthk6
yRfvVtjkrUP/P6W4mn1sn7DJ7yf6l2tNG2RBYvqIdtH9OF3VYC2JpXjpoqqQyDuo
4mE6DxfOBhjxedBeKuVMfi5seXl6RaZlELhFR2Hjer3RaT5EBwcbymAFBaHYxWVo
WByILHIBqAIQvWM/UvwRRWD8A5P7nInT8/w3bw2oTG2Mj+HWv/k4ml/oQQEXdOgx
4WmJr9+mce2C8ZccCkDL39Xy7Tdl+xsEpdakMYyb5kDNqMJ9MpvKfP1nUPmpPRqx
MMPajrms3iq7oC7P0DBj78eEluGd6LcOkoxO+Kwi9bGpKgaYy1PHWeuuJwbsvebc
VZtM8pNnwDsr/SY+ZqDINAXbLMZ8s/wk0lwgKL7itq5op5IsNywST2qP/iEBhMCl
NKiI+RxqBR6g3+VPcu6GetuiYWwZlwDUe1/O0dg2YuxflaoPwSeYrSwadwViyaoj
g4Cb5qKRL3OIi8TENtmt5Ygbkq/GoICgBk72FIfxoCDbDRquzOi6XlNWJvc752a/
DZtsN2PX2UYu+XLe1mDbkk8XveFHagYceOc7OihJpxOR9h6vQNSPFmTtQvPq0DLe
url2cfmhDf8yXqE7kYAWPZ6A2PGtU9Dt54evCsy+eF6F54NwS2Qad6o4skn1yMk1
ud7Q2AwtmVApvojqJDrbWpddw+5zFHrr1YurNGSKtRncnqpblYoYiCId9PuJn3EN
J1WXtybbXIpvQlyZ7jbP7zTWqnwqewl5a9uKQ4UKa5VQAjHk6itHk355CerTvUCm
GkHR6yi4kT/mK8H8Rb1kmOy83HWDn2/JdzUUkf0DuG0ok4vJMl//aRbyrMxJrFmj
hDaaY1jcABMUJVZxKwqE/nVWRCu2f0hDmwT/gregqsOm3hJMpwNbKefBvp+CRT/B
q9U6bpbvZq9zztCoRJT3FdFBGmPxCVAy/xIXTIfLVizLlWY0A4yH9Z007GA2Af3N
B2F9x14HwNVpNzDtal3H9wy/uz8OEQilVwnz1gEJ5I70ppIBlPOtuQ0bw29LW4Rp
k9cSvg3V2cSiVs1brzCu+vFi/zbgL8p4uLom6VilWvyX0yCLE7QNl1G4oJUQ3MVq
Zls6Zi0PCBkwjQ2DevFSrFycRekG2dofaNgrzvorA958xMHWzABHymOkoyESdUr3
+sWCgI0y1UGLPUrlNKV5awihvvKxJVuRiefXizP9QJfJ1yhOTtvOukvAo6M4aT/l
KE9+SCv5VdBH2VEEbsQDk2MBAXi6HBnEAc8ZXfTomd8y6HZvqaGXGEo4Ni/HgFp1
7wOX/7R+TwlpL0gnE8kl3UojDAZ/94jcvsLiih+2Q1qms3A/7M+2jqFRWjEPjIsN
dbswxuRqqi2gpG+569doIKC4usJxywLz89U65fmUVJ0lut0yRh91lWObiIPqGfXQ
IB7dzZ9sEu2aPmdTDdjYn8RWAMVABuvb0fDs3MdbeQ6LVnn/Ep9LORoE447ne/nv
K7waHUj6Aug8Qiqihw3V68P4xo4gWnOPHg1tOJEzLjwX56qNWvVtVoWspOvD2VgM
gGFhGAVZpk4jpzEHU9MfAn+REzWJfDYlMKTdfqa0B0PD5TUz51vEBVtfZe24lEJc
kF5WiBMagojIH4izVj7iDks/wPliSVgeVbaWbtGXKShcUurE2ALYpNMyHR9pz5NN
f9Cvt2KYm0kxRGpFzyMI49kWYehPtU4HY7TqHTBylLNf1tHoDwP9+cjdvjlYTLsV
4jjXbWEMeDk9ASOuEHpR/XqTnvrYqyw6mt/tA0oCujLuqiJ+jF12hiZCWKQ8Dd1t
WTrN0XR4PHeHKoYsnDTfTDyVosSaerk9GddRJkUeYcieh5JBFQu67AVrH2Ffz2F1
igivlli00yEBHd0ASt94DiGkF7gAsZpBsLel6zOeNpFriH9gCiym5N+FXqdVzn8c
LK9JuFYFSoq8tkLZrvI73JKL3zRZQ9wbEoMbYriJlC2SCtzF1qkvEgFzVX65RIWe
JzCM6a+YyI/5kPBY1OF0vJjYGrm6YbJZyOITyBVmCX+KzlURPcl7R+Lyq5VkB0yV
Nss+6wtHoYT9aJ9XiLm7ANgcRbfw365ouLfhapyuRgea+RyfHDj5pOv55R9TXMbg
xvmHSLh8f5xzULml4zeJb5PpvUKwUy/SjBoBCr7iYmYcC5RrHUmTgVX3qp+3/5ux
w6xL2Vzs8w5GU/S+40vi2lhXvg8YEeRWJxf+fR6IEUnnVTaAO7L1CvFs4FE7z0Do
MX7T+EGC6hEShQzbHK07JD7rJCUj0qZVpuizN0U3oQXnR59oFFmgbrgvsNDSQ+ED
G9xN1Jq69Oxtc5b371HAJGJ8fkkoncpAAW6tna0L9TRV+A9cZYNL4ihCkf6KbZ7c
LgJN2nu8VNpC+sGZwkLbnz1J4OBr9m0JTML2VeFZVR2xvNJYdBMnWRPPSaKATd/D
7QBBADwYuLnn6Jn8b7N2Bca+dtgU7tDPCAY0pS24LPKjKI+njaTENBZNYBvsTC9E
UhNE2jNIPrTcMB4SQDlOjeKvlUJ9rvpyBMXkkJoZB3Pl42rmGn22Euxm+EZofQf1
YYvTsRykiNMFJLarZYNbjXPwQB4QIenS9LYnYIYrVLkE9QFoUwkl++AeB66O5B2E
DUQXNVoSQAMfgo3jF/cRDRRKSnSOEyyFAv5Gr5UW5Z2z+Eb21m4gsftUAMcYctRu
jCyftTttRYidCLVTtD0holjW4ARe0SsuhxY9KrhdxIWvjRc4F/CrBiSVHdxDlVfZ
pPFja/OzDlsTn+jw600ASMyrwVq/GtRrGNf2JfBWam7INWbsX1M+Xd+7cAwChD8Q
35Pbzr198p9XbVu0C1s5IIS7s7W0yfnPhNyhp4bLnGE+8Wy0RV9X/6pAjBzryhVn
+gDqleM7CxrMTvWSSdC/SnzPRIh6a45nQ9KjqLOtlVMRbzqgEJsBaZeb0nROo5SP
gQaCHzFjsQIhu8WqHFe/s00PT9qFhgD1XcSwiOi/ubpMGPgaZ4q1FI7ciQ0qBNKJ
YQ8J89vuLko9Ox8wFgwbu6xtbanHJMmEvQqLMaAl6OHMoza5WPk6zGUwTlWC5iEo
IrGwo6hWBc9C9jpfCg4pdy/P6P1bsjBAqDo6jtxg+TmwYSF/ITItKRo9adJClp+3
iHwfYFXbBWqGfJGdoQVM++fSqjzPILOrDv1RJODBT8gVedQdYK9RkXzus+iHY71P
OZgUg5livfx6/CGsQVUmMKVrg1wl4scS1G16FvQ387iguPZRgjc2mIz51OmEFNVC
qNvzoEUR9mmmP267yBTF87aOvW1XBsxMobNDG2SGdhBILWexGh8W94hZbN5Zj8be
4uUrScGkWx31TzKgELSk4UEND6o5UzecwDWPXRTQSjUysif+YwBa7tmTU4O1KLw6
9ZrHIpyrHielG2/Ap8kRYI09iw6I15wTwpMt+D2JFLaaYUvtiHgLFGo1OFOVHwIw
F5X+5Ns/IQClZA+zjKH4fl80Y9cpYVk0p1pkV7hWcbmurNeMHZmzj3bUOfRKWkSo
xvaK7rhwhE1BvJnZqUAzOaygTovydP8MvzUA0rr8YYpD3+tiZHlRS8cqkOkl5+XY
ywgdYv1wAdqTI1BZ1a0kog8ofl5Pls22zJfJZyRSWFtXkSmJ1GdrFO14zFGLyois
1fR/IiQ7fqBMODS2RCEVBjD0cz1+10SZkAtd+IiGJfLCLkqW0MqFVxtsvZk31pMx
iWQ/GF/58CT02YBkXi6VpioZso0huy7o+OgsGU3x17iW+iJb6/umJhOUIdTtENYP
zB9pz05J5WeOmY/18eeiQiNEh6+gLIqlJE343bhJnkTbVpRzYkxzpo0LJH3QWXLh
BcwNEqG5/tLYyYawtgIPjshMS9LNQQEqVMJbvg4aTIlbmjm9xdgwq0xAMAO5yNW9
s5Da/hkF64bzw3eV/42mMG6JpzAvc45Ed4wmD6/aK0C9BB6ghu5Xwfac2vrStlqq
znkiTvd58p+bHtmOc2S51dQyH+1ltqtHWvtdjPFSxnTcbs08k1i4c+K1zfsExfGs
oSUKfMhV6kTFVtrOp2vjT0z2Z1N5ToPW2dJrllJpWXq61yIEWw20FgcOYOwAKvQq
rxrFhbWCZ49tnLR3pV17w1t78ip0pjDcE/ojyjznBF292AF6DlQ/x4Z5ZT8tcirr
RfY4JNUTxXmb/rj8al/epvguJrj0jBapd2jKYHIq3WrP0CnuOooy0ZqS4worYsxC
Pmx6UrZkiW5Obje822ZUmPG/fV00JSuf+UQ6bp9Z4GUxlnHgq1Q4R/dLqnSxelTE
YsOL1HCqVKV9T6JSotzjCXKLvobK6rCKCGP8zEAVxoWOjDijaWq2l5DDlWRLxTaM
nRdldLLATAkmq1P7JkGcJEzQMTzwq7KYEkisHqtiaQe5m1g/3N0LToD2nievLcoo
1VwNO9otgr3tZ1iH5xwjg8LNG4fT3l9/msujtbB7689SZwXwB8cK+G+nLvMg5Dp5
TzcVUeTJx4OpE9lJT0VEmL3klhjVyQ5zR+LL3HZb3s8iiCcBgFKh5aVaU3jljGr/
+NmIIpyRQKpjloTei7jzSOBG9PrXHNFa9RMlwlXIkUTylLWRwh0pGLwE7Ho6Wt2Q
ZI4F7dBK+0ECx9zfOHojmnLQ+9HF6vP3GeNFWQ/4VYhZRbemBffLeGvdbITOO15M
HD6uU0Mz0eemhSWdhz5ZezeDVob68oljt0kQ+Xf4pSQ8nKcbZM6UbXGE79WQv15T
zJpwwHJtdkkiynV/MMPhUso1fLJOkTMjoQfu5VjcKbXrngtMRS2F8sPmCDx3Krr5
FguO4t3MmCE+S55M+BiQSd1DbJEO1sYg1IbZyN5pWr7DT9tobkw/KAG7U5IANyyo
a08/j1t0GNSCA1tfzvCbVOCDc1NzmOgjxUhJwpvrF+6C0e8IISJvj4D9Q5uyY14W
KmivwqEHQ7V2IRmObz85YRnJbQb5RNHZz+Nfy4Wv7+cFAAwuCrer44hPO5W8TCW/
JsCdrg9wGKjNG5+homgAQxtMWScHHqtYxfPQ3Jo/KHtc5P6F8/1wmn07egtG5jgJ
+8G5ua+9VIe6beJYmMSGrBcv0f6cDArX9lF2nCrXyfyfXZqZlyrYBMIGEROUCGzr
ZfLTI4H5XbnAUbqyhEGSkLRJpOlxnPSPyi53T9LtJt4PiFlBm4XVrlK62bsuEWja
PhnI2IC8HTvfV1dli94aILQGP9wEucxtm60OYpM3+bRtrq/6i4YXHeUGnhf/wcWm
tCWxkngKtvBYjrr9H1DpaJcK73WuB3FIjcEOmnzt/1la5LJpNJp4+Jk6L+bg7WMc
l6sycVcUiK1EeuoumTu2Kg6KUxhmOATv20I1SS7iS+acH5kmYJa62sanxiFR/6gW
rYsgHggCLXR0TZtuP1kxRJGTTr+gE4z88Qza5lp44DfWbiBg889PPJW5iz2iHY9m
7eTAxCyQZdXlTc/ThX8UcsKHsp56FbCIPYRNqv2vfvsQv/+DOREi1iW1a90tJz7z
f7RWZYBAowIXXyBoEw0iSOOlKhsk3gdcqbp8ZGQ27BzZ1zi/OTCyeXdCuIEjh4qD
t9RGbjHtLwyXkLRYD2KioPuJcR+QyqzoFShP3mEJrc2lu8HFbsNDC69BmROSZ3Ol
Mv+1oXXHm0oKD968gdZAZvpblyC815ceTiVxFVzTfyvkASVExUxTzg1twi6exOpv
JpuDKUZGXvTSscF09NkLiQ/Xb0913FrgWhSesMqKbD+jCknIBJdoz7mg2DNgE+TG
FwZqewMoLMD8MOxM0IBWEi9rHNyTmZWb0t13cR0ONcfk+BYrfSlsUTneTDi5Y9Vr
qGacnt256UkcwNIiaNf8sf/yn8U9Y0Z8qWjfejwADrObDb0fpqAXgcDOSroSlTJE
6BOTFheVZWTJxtkqWjs0o0XgI2G4ef5PSnh3jPY8FvsiY1jQPbRd55W2tYgmzAmo
Le8ewSJl6TQIi5JhDsjgOEaQ+OLfxTd/+QvQvjEoobuyK2WqJEmMK+meU/A2O5Q9
n3ndLrIq/m2enqoUEkPwmmRtv239MQnynVQ0EkewGARZFj7vxwYtCjpPXabRMUTc
cz+FmPYmPFcvEWc+O1I0OzfLlzRQY+H6mXmuKBPGcIONH6tbVm71liAOlFkE0prd
QbfvIYX5i83v2KoRU8UgTbtIxehuhESoL6uP110BCix+6tqBKUQpaSYQzL9XM8st
tBHMH1YyuYVRSghmk/Y1JiWCbrL5jroue02J3D1+7vGLfLp2j6GB0HEgZmSJLm4R
DWUKaXRdDiQh1kBVcMCD676ErjOxxHgAG3E4aL9iCJ1POF21oUi1PLZMUOvAnQXp
ue7z3XD4Y7Y3jUyTiejSA5RZmtjhQdzdj1GgSj8IPsSBMfBAf3yRxO/uWcHSxhV5
OrGQX/BKThdWnTzGnQ7F/iWPOtc/N6LVBbO+aHXAUlvunmIWljdFc/+uqsMOhbpb
2AyB+LfX/xmYDCcjWz6RttVHlonQkT+XDzRvO4F0aoUyr5+ZJYFBsP/53dquGOiW
4ZS/FQPmyAaRXAo6KdQl9vk8mnqguUN1a+BOOogzsDSURwpG6oyVSu6+XIiQAL8N
3gvw9QImVhZfPn+z+lzNBDsZTEsrC0qIiEgSlFM36CJoKoNLR6oyAXb+u+JXECoY
tdxiZ4j/6IqHQsNysBCknqg/l3Z74SnKRwIZXiuQAdTCR6G41O7vZSwuOB2kFfrq
uVRtBfVZPf0psytKGKYM7Y78yDBzZw9zWYuqjRkwqJLRkhOJFRLkFQnwqVlobhe6
PmAnpgQxRwCfHlhWXJ0d0C9sgEdltVlyvJLgYsCgCh4f6C6TiOxy/+XJ6kKjvxi5
kt5GMQr93pHGMn8Mebe7BZq0+lQLUCPvCiZh9shPZ1EDQ0IZdb8ZxewZ2olE7LQ3
LaqbcoNa43QEaMLLP1Gfn5mkPy8P1Z8KJvBErY+lbJM7eme0Id9AdQZi3FSycEP2
b21yqlDoAEy3h2cvupQWWVY9pLP01HJyRrYN2oHQfHTdctKtKcEpsza/VZwcu2Lv
siNJIlFFCCDGH/3BSOnPp2gw2BsQBI6FLYlsmpIdyumo3Kbyf8IKlgPwrNHNo1vh
2TtfxRnlRy5sl9wqjTAIWF7rvr1Bs82eF18m6LZbNABAWo0J6pHhfMP+Fzv0QCrh
chTnHHJB+fzLP9ogUk0uTUNgxfTqNXEJ2lUpYNy9njWmuCKgpr39VdkFc9BByyaK
1hrRcTHqmp+ejZdcikd0Dc8rbYMn1TskVPBEzu2QzMM4D7WaMUKwR7v88fVnRvV7
o+4FzWk91Aw16nh9dJe9u/DgLcrc0GOWBe8+fiicSTPmK4M63uJ6gNDz29H6NK4B
CeM8dvrP/k4SL+hP1waSTbtkbnAfrM2EASa7f6yOFWd3mWfIbarvjGIdFr69L3Hx
O3lWrLTKznei48X7JsrkIbNhCxUdr9y/i0jSSYsg1nts1R21Bek2gNcbcY0I9+S2
uOmTSay0h9DlNV50JaLjMDGY6JXzHtPebfAshGzbeOZvdmSnvdYKRjlNUodM1nMh
v+2l/fF2PlOP5+EKQly2u54cn7llO/fBlKkNa1iWIxq9JZwBFt2+xhFgb3iAK26b
Lnrg6DNrnr8VmLnSIuwhN9N0Z6S1d8ZiVBW/12SpPHnJHVcLvo5Omp8yAbGToVuG
+FLtV+FI75YxgkmiQjEdlLvOe9+/UBXorW8D98UT2Q4rjef7WtjmZhu/oq9CDmXI
wH0wxwdLxi5sptdWmRQvAqRfgV8twYFT3IluH6GsmdcJhwTCmezfKEriwOuNHX5y
ceBfKA3S3ULHieItP/UyLTQ5OYlMYVNF3p43RUsHsX2gpxKpfZM3kB4wbA1O3gE0
Bv0QnCDWNX6v63EdYawbx7ZPzDjJbe5SHWFKPtYPZqGZ/jOhv6GyEI1Lcwj8F/jv
ykpy4w+NueriAfmCt/yK44CKuybAiQSarL4NyPO3asHKGYi5RDeEvQo6NtJZp+1g
dmPZMxET3WbuOq0EKsvSH0YEUYqHERLaCpQE5kq6iBcgDedqNJ7tSbtbFJ6YrRAv
C24ktiwGIppAQCVNmK1M1Y0ayXkXQ2gWPhZvbG8n6WTFE5B6PQEurbA6bdFXZzTB
hgEXg1pyqbXSGywQuKqllGaD7tJFuAMRGegwo/YI9l1i7L3DQ07PseQBDQNf29CT
jRv5fwpddj4pOlikH/C78XA8fT+jMXBn63lT5stnbNhWFAVL6R9j74TyxgZ39akk
OnMclRmJILQc5R8cYwH7bQDBeLGcaO1y4PaR5SngdVsHXxag8wxRaj+YUrTWf4GE
dOwx8u5n3COotasvbmNalQUS0UputBlhIZ9T/Uy3coCV2buZ6H6tGo3n64PS7ilO
7cOvjJARTTJ/0T+xhcTUz37a6MSk9KjAmOqaHf2wAWFqkhfjcyxTZD+QowSevmAx
hWt1qpD2WcZaySKoN7Uxkz8j+K7vIfiKTIkPu/m1KuD8wT8y/SYrcC3mHdM4giic
lEyRpu7DZ2OdbAKycDqugFayFvPsQIohLQDN1+YF6JISJ+wVP7H/Ky8+Y/szqtwM
o0EZUSmOr5/WcwYfLo9r2tYiaSJ+kNTLJbvnsupUcz+Lr7pea9KMrjrJdiPQGw0B
Lg64Zy1RfiHxg+muNH/tM6lJsqvTlWFKeEIZGYw/6PBLEWZwgsHYejXdNY4bjjkC
HlVayRH36QAsUsXG3K7tkDynXvhYv5pmiQBNzP7pMG9Zb3Ar0kfzj/h9NKn14PDJ
q5oWukFUFojbcovFpeqFXqBhHn81l+aEa87YRyuaCqzAUZR5xADf41k7y8KA4HXw
GRcK8vVYZdF9P/LfI25bFvskIC0IhiNSmTzk7jO2RxDG7UNmVD+Z3KsmHcIntN01
xMlt2kfhzsvnXxXOdLg4zMUOdqaH+HgRd0zo0bOGhiZUTVwttyh+i6rxWVXK2rff
f/dAgxeaan7s0m9MO4z1J3BNHKcnl0igby4ILMmSuT7kOTjL7W4TNW+kOqc6KN3b
7ZMqpQpmu1mEgy5nP1a6dvhbTSOO/p9uKMvcH6TVzAB7WSI58YD1ZFjFwXbiaI/h
1RrUtP6eCeXfEfGaftvcLnEQGY8Y0pyKzpS0oWB3X9MNw3V3liC6xY7iCtpyR1AP
jrqXnzariMauUxU18ruiQJkL88ODv9kaxyITda9ZJsFvTD6PmzhfXhMJoQH58TA5
FK9dN8Ei6G6Ck0xQ8wjoeUNtNTG1tIMg0h9XfPv09uGsONePQ9FypCOwYzJS7cPg
HX5Rf9REyCaKNDh4s8U1uSJZwAr88Gp/J+6LDajV1aQn6m1Jf2LxlhUohX8OjBdz
mg4Vo/qY39q/voVh4edmJ6IOFXSNxrft/TNTodNR7ZcFXlq64DshvJLwOTx2G7LD
XUcsSodj58Vh8+jhOEv69DvEpdHbte1g+1NEBSGFVqHaFHmeYaJKiKrRTdsziHXq
It99pE1KaGNGlFkbDZOvsxF8zZMogsGvhe/CKccZhPvODq1Cd1DlaUv8jwAlHWuT
ZLkLvLqq6uSeKrPJroYVZzvvBnwLWYrSZQXd8MA2NpM51Qp9ZoHLg7J6XdnHCTnN
ZmAVKlsViKMxdHgkFCN+yYEYAN7WNKCqJx4UTIih3/pjOOpGX3GuQto4TeGNUX+U
6hnRiIyqDGbcvPpl1y/YeHlUYutmxQ0jNX+yF0qz57MIa6T6LT2G5SP/rWofPVsD
kzolULkF/okZeBrJ7Z6bWRXEYHyRlB0d7mPIN8Lf4zcz6AR6QbQ43+eodnKj147Q
Od7RtjGpam5y508efSm8Zz2AEIjJS//GDPvYoqfzeSsGrQsXr13Jb3Quv6Q8SKxf
YrbmDBEl0Mxf2n3s7luSIZQgsd7j/hpIVwJ0Ai7+U3eX9PkqM5tiIB4Dza4ad+6r
8ToVIqJoAzngwBANcB6u3SMVaM6Jg6aCbwYQDWzWC/sfPONGshgRRFOMckuqjfPJ
610d2QX2lR2DIRhunR089G/l+eC9HNpxgDVx1umgcsAsoGr+v6Zrh2iq85oU8WQf
QXgsL/kMDR5Y4OEZF/UnNxafIsTB2Mn3kqFsDIFQr18F5C3NeBfpuvWKBLrwGNFD
uujeEvicNL0WZs3xsp/A8NErPeYQux6Ooxc5qjw77XeyZ73F3vIR3a+UAbM5J0gu
KQY2w/SQfDt0rbk/f9K3vlRZKzn2z3W1L4Nc9zbcXOG0rhOzvLBVLjzLhyoGt0Sa
D+Z2zpF5kTgPuK4CW6Td63wz1zpeNWZAJdkxPL8HOqdnu2LMDlud6SLxZo2ugaZu
e+hwZxTk93oXXe9QFzUoYu7r+HNkHOVIUOIftU2PUuaoiiivnCZV0VaEvj+zmmQC
+imzs/wcQ5eL2yOHFNk5Y2C5hrjOiO/cXSfT2eW0u80atzF/QizcUeN6GUxbfyjV
hPD95PKgrzuTXdcazozq3PNXPYEXw0m1kUmAy9qklGbthgZY7iAKrbmd2RDN3uZB
aCCwtWSQ65YbCYhbyQvsR9oN8wPR2BI5vszolLmUQggt3bR/iMJk6NjfAFZDgqSS
dnVNx+IRMNoHPNE+NGvmfVLr0N2vopR8ZAZ9Q1MlIJs14B4nFrK5Klyo8wt457QY
idDjqkwL+imrlibJ6GkW9f3hb1TaPNjwYWq0VwW7F3o/ZZiQd03dhq2BRjRmaU9J
g4r/TN6TCpG91OgkDko0JXO0yhiVWSANyeMCi23kHtCPhYW9boiukbMGze/s/98d
hoYxvvADd4or90LhImSFgb9jg872IlGJHwt0O1jjbBcZYZNRJkdA5pS3c12diPIV
GFHpphuYOf4zYNXOQQ5W28uVWbfMdTAwiFBbOEG7Hfzgt00//iyB0Hz3pLeuEHMH
/UaYL76bVML6YTeRnGsG/xVDoGpQlM/Ycg7HIf5p81V8vaRG9aZeyNQE5xWs1BvP
taXGEQ9IEIZW9Edl4LH8JR8BzVLt+A9nQEAOs/rXbss3tWDHLlfc8X6QAvNoJgLx
m1KtLvJ2dbe4CJxoNV7UWETTQLk1Ddw8jqBsoOS/rL7ehH/S92VnvLU7E12pwPP9
yLlD3Srlm0HU75rUYDGCPi5p+qISmLBd+5eRTGlXgXv/yPrcE8AxClAzNjl/H7xI
2Sxe68VODbtBiIEKvA9sOX8x+PG3/96NxMwcfNQcxKadaw5noajOqSY55K66uR2o
BG8c5oeo3lAko4z6AU5Vn6BTdltWHMPKq2luYceP50p14WAb2IaMxCxjFqEm3iF5
eVIQm9KNoxetlByGCbAvU4JacLllmk7rRCa6ZaXn7aAK3nrSU6fGIAdijc0VVf3Z
RsKZkloZLNs4BHZYMw/9ks2SOZAsN95jlAiYw4ikjaxyKBtXDvNEVKrgmGkDNKD7
pTzgr3V4V7K7hZv5V6R36tTiAY7lIdmBtU55lQk8zHXLwFBd95Z5aKLiNHRqY+Th
luAsV/rbSg8jpzhb+6jzxS0TRyFRgU8Ch6LqwrdpKrTn/XyNXxxY/qd79NghI0Ew
z5bbiA91n4Jf3xUT49HQEOQvi4/wNnxaORB3bkpSePUQHxo0weC6aaU8L/Vob41w
CtnMu1TpZMllXan2NOmfhJ4Yvtzz6zZzEheMJMeHTDRuv3w2LAuVlV2/wD/oVigW
Tn8Lnb7wMs/nsSUaZ+et+XuoSWosQW66XFoaTrkEBrzgiPACwZMLnWW5DuRc74b0
nhrskkCCMr46eI5hcdR06woggMmj7Dxp0TInuz14bRNpjoMazV41IMZWgi9HJY/l
o+/SqmzN5Htc08dMKPdl38nOoRBX1SEjYK42fRTER4ACCHhYhNtCfxm49N6Qtjuh
i/TgTCV4U/eJTEciYuOcC/Po6yNqMwJFm+HOxy/pYE2iQgQKim2QjGKS4bEB2tqq
FqTFKZx77Z01wg2OImIpONDqaDmKZZfQX8YRx5D/sT/CLz582wlCp0XxaH9mRRzL
Uu2UJRe5OQQ639P9Ng6BVYXeOqbjtmBKsHFXvNaoRlPKKHbMFvWsizZi9wTCNzpx
qkNjooqaRSHeCmpwbfwqY4b84YuekEB9ZxpmE+JUq22v6ZQrPzWRO6eeX0y3SLTT
hk0rglzjQd+8tXcAk5cjYTfJCg8ngF4Cnx0B/PPZmZ99+07mPKXczdGr+3wa+F9S
droF4oF0jBqNQJK8fUYw5AXT2CwW3Yx5o3sV1I7lDI4JzXDhkuZyBAiIJaUItCo9
JUpa+QH3l7YmuWnSJAfhMe/u35/t8VcSfWz2JqSegzcrFEFuZsvhUFFbkBSarS+c
4YTjkGAskhREHVEZWTVqMEd6uCoexIkIT5sO6et5ueIrXKTBRuENlU5MYMX8Dhmp
2sICcOlpsZfGN9VTNZnfYYQWW0pyMF4QgbD0OuPJRnpDy0Lahu19o093538EgeDu
aTrfqNScl5JlSApk5lH1Tfe5V/GtiJ30JOkCoRubOVAWHknlicL6y8TolkDGPGaw
+MZYcHsgspcCw1o12Z+KyVl7hY2GixZVpzKD+dQ1lg91YbZ781R8K7k5B/4tTB8V
h/Usi/imrEImAttZ8BpHeLbS6eS8ExZB5o1576/vUx/iH8MEuM+mFbPP57FlvG2q
YHG1VKlQ0mn7YjspOxnlWC5rziGbIZ0kkMXQogPLtVz1Ixhx7JMkePBBoBL8evq8
VwSO9Am2StMg30nKLsP02007LH+5tqtf8Y0kZ6o16HpTpnvZHZXemyaoV6enWLI/
MTmeUY71qZ+FddPDYQptFUyqoYwj8oJvOz1l8SpR7+GfMAsq2+R95d5MtVFHpfv5
/yM0GaqfjZCSOrdj/SKGnp5DUr/JSWVBefdNfNaNBY+8u65Jt44/k9jslS4TM0TE
lQ280DaKp5Vs+3oKzYXoMbFYW2nRz8U+CAf2eBVjdT4IOb/C5YgakPiQdnttH5kT
3au+jUH2XWrEPhaTnKh+NZdm+nXpmww4+nBsIpfvpCcvnYuzwNOcxD1/Uj3Tdqcl
Si/DlFGcSrPGNJKHiTM6oRdU3rqVmRcsmN7+LEEGslw1OJAMblSI4MHT/5i10QpY
WU/LwoFoSXe9A54uuxvmbMY5s2bNqjJeUnjN92F0uq+CClc86TnISMkfeLcKWVlq
jdQ0YtW5bD4NoMSvPbIUqslneyf4D5qwi9QHOPe0FqeMTXqbXQ2NX6I6gA2DV9Jc
sO2M9yPvVB8SfW1f4u3Aolabmp3QgliZu/ODAdIlUKPIRngDmRmwOVH3OCkNSYOg
BIl7TKLs+0PLQ2vy7oTHPxBFcrvFgrbC94UQrhmYKKWhhEb6TPSJ7ONwC6tO9KML
aX0JwdyEnlPKvLC1ozVTr3vYvB1CL+ZGtzbxfpVXX6JpN6aPXAURkcaWJYu3oV0I
bgTp9JuzWxOzpx+lPzdqIZppri8p5yFSWfv04ZdutAIRFo5nxYtnGg0z0klFLI4t
XITcOsMdwuC6di4dwpE9F2EXFHwwwgv+r4JakaNp8IwYp2Lb8+7buwwNuFQ5DJ5W
hOpSLpsT9NelthfnV3ojbPlWa5C5D/RUNIkAoNOwN3xtX0EUKfMRA++sUIFVuBjG
xjhZsGb5pRbGpyLAjJqTxYInCRDHvQZFrFjIbanNaMGTiE48uSVJ0FIAf3F0xVWt
/En5K56FfdbjC7FNyu8faLAeCTcNZcHViph8FXMQS/8ZUHUgUacTEqAS9JR11ZlY
Hy7i+HxjoKtcjK+b+X/lALv95Pgfez7KvF8gO4q5Ir13dJ8Ud/tpz/dSL7jxmPkB
Xitesj63MGJlPl3yKSfuRikdqMyskhUhZDd15tLs/lYCKn+KQviLiVIRDVT1faou
bIHdhOOe6h997CxK+Di1Xkfq2NR8ryhOMw66HDquPJ7arcpbfAIVOcgLgVXapqAX
EQBiVeLx0+bhR2pEN9OodJWYC2MrH1/aLw3K3e12k78j17JNcG5A74vGm2w3Vfkj
igg5s3d9k4IFh1PPzK5fuH+uuJgw1cLKJxLNaCvcxyV1G92dAg2eTEuNXxF6DooI
1jbcHTDnnqg8CNvUZbpfXGTKfSeeLTj6m9GS8fqqTQlP+lI7LcFawACbmhvm+soe
Q0zA9dL6nkzyICDd3BjfVIYn1Rkr8qvQiyllG/8QgJVToG6u75EBYdfubqb4E5P6
Q7xkUL29Uczv6cwkFJKXYsCY7nyOF4Z9QsJ7II82T8rIVe2vwlQ/E8pQwbTiQh8T
JAHknPahIcKKvd1etJY1GOcDA1ZVue+TlKoy9IUnFJN4b/Wt8r2SuqAO52V4EUag
AcE4Mi4shS9pfLBaK3fjbjIC4u7/6HPZRXLmCuUoFwRGffC0t6DfV/ats60cW/1z
Sj4MeRR2ixxIhiXgppE0uLAL/uiJqZu3F/sc8c7nt19uThJB15dOGJsu/FawT7uE
dbPPJmUB1+oRVBZd7bc6A6vJ9VhcarJbeEXiAspIcsbZDNp8Qfxwl2pEAZb5BcAZ
XlEcnvDuVRMQPJX9nij0F/RUt/5pngC9g2OM+II/abl68eCSzgiZELarUizb/7g2
wE1s+p8QthTIzDwCnU/l/No7lunzfCaGLqc404RzUcf5+m4gaDmb9OsRY0rupZ8N
iOVEFzYBmNLluZU2y7qt0O6kFPTQlwnCsk4JvQArzq8rYEx96cdVzhTC43Z3N8k2
Dk5hKHNTWx9NdG0d8doI8xEovd2iL2e6l3NPZfHMFav0UciRUywz9mkhdPWfBSZ0
8nXz15NvirENASEEP5IXvRxEifVfL/PtqNPJ3P+Sy6fut8+C1ng2IWKXexVbN+nw
qKhJr5EGOk3DfvMz/MtNqmf5+i0MKqlPsZJhZWOhe37LRDC0+/6BXVDE7E8Q2hAl
7/77FIJ/X8b+2qdwAPzK8YKLMI6XJ/ROb62hkR2tw74beqz/Bk1quzDmAtHI1Y+d
3SqR5rTF4V1L9jt08i3s7X/0O2xp6rXJBPqRqiSKTKrGIiaZFW7vZEBV2PzJu9Co
F6CljwvfMHi6NxtEFm5W2N9sfB5ZaQL2JCeq/1EGRl3jvdUKwUwhkYnwSOnOdZEG
B19ZFtXao7kR3sZa8St91qaIsQ6jmk+nkHaISFIa4O+6orppn7n14CEb/YuEK2sG
lk9X9x4XVQfGgKsO67jC9DXC8//iIiNnYnFQYdCSffhHLejI0PG/EBUmHQUL4ggG
touJnw90XINBW/zkipiTwct5WfR0tbH6ZsAHrqt238LXo+27KcWbQ7ygFSfO6wJx
NmVEd4nPCTbIHjyhDRp0Rpr3dYPo7K34YyFlR7k/8QuaOW/WmrmMjnKnSmCUgM97
AzSzZ983YuNGqZGIr4ZyPsin+fFO3TAvp8NGxGSVRMyuNvhg2sp1ktPpWDLv21yZ
8+9aViWUXjeK74faCdb1tG6JUy2X/SIS3/I71X99VpAOioNbQBaAgSmfk/dF1reb
6hxz3YBM6tHEWnSwx5LvDpQIWpJH4YzvRiXu9WQ0xG8oQ6/qw5r7PCy7sLahbYyF
yZx872TAl9Ui7Iz2mODcIacbPTgulvKO5GzjsVcnDVPvvaKViZ3IlqSjh6VAuqHI
dIELuGjuBr51H9h6R47ByLz+WFKnPZ+ImtAhjz/Ts2OUziAmT4eAwqDW8z6wP6CE
LPxrqXbEKlP/gZaUmhEoevRvCu0uVcvh78EkGugOVuGaz7UdVJOlblunn4HtbIBS
YAqqi+AltvHKI5gvpS0WSxIlMHh8xliMuwH/Zf654A2b02pgmCc39sTHJJmf2Fji
vnc8+ut1SydYlM8CLCpXElLwNO0dCboUFCSRlQREqiKiFIHo/rWQHlA1aktYrAAN
OnxdaRI46rSNFQv1elmjlOxkqT3lJ0EPu7e9U+hdw2t3/SlGouUUfSOFn1qB31kx
5Dg+XT/lrDknl7rGSyr428hgQxKnTW8EZJfx3P9ErkHsCi3C98Tl1wm+IJBsieNC
8awWKhms3S6OWMu7mU9L1EcDIZ5y5urQDzs455Wl0lYTwGfX6Rlrw/jCCfw7VOah
LTfZmD6e8TnOVknAXd1eOHQL74DrrUidGwSUpSh6c71XHZLVPEw2XuTUnhmjp2cn
P54GU65oXbML3U7TmIAwKoBUFAFlWrdZXwqaUHO5jZS2GpcjXV38svNzMp4rFwWu
e90CwI+hleJoB3+Wp+xXX6M+LCYiK5feAPOnLi4MRMxXEeXItpB7G2O7jxs0Nngh
39uDgI2JNtOOiEeDs2s85GiETB+BPayCyEtmEBB6VKwMx0MDzmxrFy5I2RwmRnlY
12v3q22A6upMBBkHj0V6xt6v9Z+9yhUB6DVzwIHj6gMEGf9LThUahmew+QRYWTAK
QUn3ztzKyv9n7l4gWdLYvRxEFNW8OiXEYOlss/DhAkU8k1Cw/xzGF593khIMrEy0
n2lLMo+amj8txzjufuaqTJrrPr/RDh57j94gnnXxOkl6NHLAyZ7W8FTa0s0hXklA
sTdY4F5RmBZCir2XxzdXjKrVkI+SWVVfTB6oONhTJkXoZ9tY65BOQ3ftjt5i2MDo
fSWttAvgZ+IDnQvbZCFjkbNaq21Une+ZG+kUqJcTYI+9yJh9UPi4mXg1e50e3gap
4eFl7RL80t6qpgrezDweLxxa1JZgDHxNWbEWyqVblbBa2E9+uOJKI3PfLaW2HtLd
aqZyynG9chxGpZfd/N7r1cKmTrEIcLo38ewpjGMDQNx4hx2mhAEN5HKcyHk6fQyC
ZD2N608jLT2N1Uz/fCQVtmCNkW7c2HakzHP1u59vLKWrw0D5GxOfvNmURkkv0ad+
BvE768dKtqKj6tzP6dH0SMSUbVBRYhzAwGU+ILvTreg46rba1wzfe8V/mQucmxIE
02DCnzfvpk+m5sGkV7Kc5D/pGEsE29/PfSQTFv8X15BgC3cQlKLt8AjxQcrUI1kL
A1vHMZMueaRkZa5P+MYBlLJWf5nyYvRYlLFZW0XHcvK4pr31JXveBlHlOJZi/clF
ILGLNbr/L1MglM0OELvydEQLdZFt6ZqGpqpBYHpkDobrKAbTyTBh5A7uXswreYwK
RXKe5OU+GqqdEX0ajDfDVvlGSwJKDjuSBxQR+8WOi1IpfPt8xZj1Il5RS5t+vgJj
OC9xEPv6CZLM+M6DhAhi8D+8uxtxO+xnxg1HsnbNSYxV64Aa2NNnynMdQncStbyp
UropHa78bhyAo40/LkB0WQSjhZOrUj28SVXgVNezhsYbibp6G/2i7p6qVJfDncHW
zwKSJBC/cqdG57rlaMP/mJ1rGD6Ri3BRgIojwxzvUAM08T3X6MUkkwsYMlcC62kc
bM2+dOEps5qt8lB/6Fd4WJTZ7UQpUh7KmfXhYg0AiaYXwZ1V+dqT9G/jMK9gZI/g
WG1xXcFrijw7FPncynGfVdmTx8sP6lgKly+zBbZBRUH58rtL3E5RdRDID5SAHdZZ
N2xJwpJaxXLvgXKYkX3rxtHLBPms1FKqH/HRnjjX4z6ObM95bbXxUYs8xr+CJWze
F/hlM1yEMgEBBXr+mrVnKNvXScXUqPROLGr0SMkvUsKJOKCb2rSl3R0F3LtsMhqh
jW89eH0bS9A0lPyv93A7Q70yRkurbDdzkOLyCb8cayE0CZa1+ub2/XIcgnB2o2YV
/WjohXDvQFNYnbyI1nA6mjp3QwXmkg4jMrarapFdla/5Ldwi1+H7u0TU40jxVnQT
Cfqic+ZJcXdYPDzMdGaJIihakkDJOqe9jHPgfVHVmgQxmqb02OaCV2a6ysZhmzr2
hCBgWgebzMVPqOVU79aCEPTc/HsyWr+GZy2UL13LGgMpcnT8QP7tQAFx31XRfmEI
MrygsyKQGaXPKSSW5AdnB9BH6loLxoFwTRwbThn+WiAwXnwVfYqUrDIzUHJYIo65
fJXIs3/ti50bQB3mjaEGTFW3C92g3cLG/vCwDAgRHUrH+1qqlWxrWtRgvQLBs0Ve
pnnsiT2H589OC5YPu2VAW1G2NoBhQCRNWGTMhO/U0cwUVSHMU1Qxv6Grd7yB5bnL
ZWmP1DGtdppCZH0Qn4NoDUnQ+CvDDCLU+7V1gfm/fY8Nk/KSdo+vMwcGxghjzFmW
9uIsAOUPBoxvb0D9MLXJ4WM+5CSN3uMBHpWx0vS0lIfhOxI9x8KFTjAY3B5ASgPx
z4fkxF0XPh5lbKkBLc5c4zobIgFZebQmi6pCrtE9+QbinxjZqi53jo+WAoGbMt8t
eBs331XZlL5nFFuQ4dxobc0k9u1mK6kUliF+LXBZJqGCX1o/Xuor003U3k5UpqgX
QU+3oBQoqT6Beuzkbi795rO3+yaccrnaWbULLOYRBFbVc1deczu5Q5D6L/b70QUJ
DyWtaFm52MuJVYx76u4TEe1hHkffdHIi1PeaeZIWNwqitTg3CWEYUGWiSIx9olZ0
7vqZkOZ6MeJ95VTeDNlVHutkvpbnjIbrPVrCSGfBEdsK2GZnXy9zB33Onl8Kersb
sLe/YGaCLn2R6vJDqqKxsD3l5xibIJPcKg2yWG4bPK6Rh/Dkk2LOVp1FP4PGoBL5
2LtI4W2lJ0ClSZr+TI9RDTTcuYh2VCvvUJ/zgDAEi06+dewqeIJdLzUnUb0CJ/7I
HGKWU4tX/XdMg6243epaL3geEX51NG05M77qtj8VwvbChHvpi6ufM/9l3gokMTpG
gCKk08DUnuHmGoK2tGx2F2i8eS/h5fq/kO6Og1D39pRpEh166jWKt450xb3+4B00
cLevg+bS6sAVs8g/igVB5q8xsTUzs9sjkXUMsTuaIx3Y0fXcHrlXryVAuZcGLeDw
/DGKF7Az5FD0Nc5WAfRMeAEJvqpUWnuHaYlsBCICwO65VLIY7D0dTgRIKbot0XvZ
GBc5AUIBteC2vptNRrKourXsGfP1VSUuqb2WkzPWFpA1XMOPtkEZd8buxrmjw3yG
ZFzY6g1XKQzBKw4XE2Je1yskJtPUadIk07Pctvk2wDvblU/73hDk1X7v3RtkB9C3
R90engqI9GQr5usjx6mEP7N4ogIXnEzY5hY3yvrJ4E24x00Knhh6vdnVAD9FWu5X
Za4sBAIsP5WM5sY6UmXYWeQw2dMuJ/jCfeW5asGsCelkEmP+S+xlm5UkaJb5te9P
sYrgyA2Pz0vCNmDI05l3obQVTpWASzTjvxbZpJ+amA2TFYaeYYvwgeZNa0OYLcwU
Zt06Bkgn2WpdX5OhWClGqF+bR9mne1hcqmvBM2q5ixfajt2icwPVthTxPqyFMCFc
QoUmliYYk9RsWzwJCsYlWWdDCdn2ctNMbqlF+Rj2xise1fNnQAiJ5aDJKE5GV3Lh
vt28vdtNu2IVikduyMhInQcK0n8vLrP4ZJ5apgy6K1cb1a0AI0A/HIrpxEBBLVEL
ml9vw9ELflOlFU6Cqia7SaO6hnJ6t0FGh35+k3Um9gj7IFoGYOtUZ3DCkRMNTG1w
jHT2sCPxRoAFx9NAx/PIZ+WsatIXNmDQkCCXyORjxbM8fsCZIMpUw15a03Dz2swf
9g9e91YsXGUyMxEsJkwuMNY83LfQ/4PI4rxNqeor+OcMn8FdGZD8FpjwObzoh4UA
PtHjYwyzr+tYlTPLIhyOQ5+VcP3rG730PKO62JAV8cnC5u/INjJoXn9GpgHsf7Ml
DkXu+YNTx2b9FbzNfYi8B5FDa7MacATwyzszuJD9lveY27w7OxGGrqfdIZ1vWblO
04WncigSiF5NZBrQU143GdH6xjpzCjzar/IBrnHHLpKpHcCcsT+OOPiikI8MUfOg
+qcUwLMRQXgjkX7/SROvEHEnFa8ikqGQXNcV0xzp64/CbiMy1nL8+9X1GKg2LxkS
sUN6fkPOIzAxgaa/LvOp5AmonA/s/vuvnvZ/1vIgQTJ5zUOvKlwx7G4Onc+Xp3cp
AOfn5qS91sgiU0IeNgsFGor3vayIPGD/Wtj+gIJfTTSImS3mT/ehSHKqI5Pib7h3
NCLghPeR4wWdq2sPefkTJSq1EDOvRjJtyDPcwgcty94l6uFRxOPBAWb46RfFUd1C
xHJ9xdprxTgsPFpopNS4zsTsUO6OBiur/91Mlcyi3vFY8tECy3XVhWuKWGZ7F8KE
qZpt8RQcgtYXpBGTw4pPyiZ4AJDZPRU2M3SyhIj7LK7ieyQktgieGAyRlIuC9/4X
Ej9p65NwmU+TXo8PkRruiGAd3G5wfrX/GmSuunXO7vi38Ra68EcyuP9KPkaG9fct
hrWHbIThIYe0NZfk/7wzPz5vocvqzVyjIjicgCEJUB8eteNDNiBEcXzAW1VqpvGC
XhNXmJ0QOD4Olx5YQJAqOD9AlLb5+HAl5ZHJhHvdcULlu9y26eiwS44ULral9c5E
pX+OK6pHi+1sYc/nRSmlkIvxwSNQyXs7mAFiMNnZ7hklbSgG/xiVQqbCI+Jd3XpW
tm5q3QSwYbin9gOF0eDRP43NPWjM90iYejn03R2qLtp7XH8xP1fvzi6HNWPOMT/h
3dBoTmSN+5Br/xuXEObv8stAd3fy5K1oIU8NkrbijHPFR/dCMt8ue818sNYayB2w
ZwL/iEZw5SIUCKzpc7NpYeM1vqJziJqyEmmkQmernZApdKEtIsUMbyRa9KzIW1Uu
6ynVi35d3rTCrFMkMx885bY0QZuLtpywBmeqM1AAZgoFHpTlbar9+PRAi8N6Id5j
lUEHxp5jxb/3ZF88gv1xkNv6x93anojkDOCwAN7j7+iOn/TcWa9nN1JOONfsWKmm
LggW8Tre7Lonq9N3W1HdDfBAEagx0NxH9OWgq1Eh+BYtP3BBNT9XxNvb1JYB3Pvo
izkpCAoscOdx+otUpCS6V5DlwTrxsKXwb+ooIYJiiIjYa+vaNeJDAzG1rJqB1ndy
3Vc+9j8zfdktFv2oLNopsQ/lvfqtCOUYkxf6PKWhAV+PPYv3/z1Rf1BcKFx8O0P9
3TUs4pu87OOFhQTy+qboaGKPM6JY0SVDstfCY+P00BgzbevGOl7L7T7eXMkV0Ecb
a8ccASO3yiIpW60lGawpDCYhL0TDT/MTMElfvsCrXTcWDKDrLt76mYNek5BJIjLN
2Cah5aENOjOvvCpMtHZXHFSpwahHKNu+H8hRjIDY5Wn7se0urDyvrCr7Q+GyaPHi
6GduG0VImOmpZLaHvi9Sz7WEVgDNJX/k3dLDDE5AxetZcNmFTU8gyJoLA+3DZYVw
fz+oC0fL9gYc1smJSMRJ1v7kS8q3viAsuEN6A02mBSZHp69lmUNGeAC30/syDJ58
qk48RSsc0EnM5+CRg2UqnFjiziS6452nLmw2kD4kMBMYDzjoukKhafIu+I3jok8C
Hhk33kQ2JgrqveOQpYqVHy3JgBmrkIljGssOUyQpylnfFUMP3KjCP05haWBJwYOV
opxNhwBhXoZLsqcix5bGCXOzsifQ/MoK7AP1LAzZpbfBrLYEPNeLViINDYAAIsHC
nlMK5lZ6v7AaTW2WppiBK+jWimCsw7woKghovN9Jc5zw+Pyekd22RC+jEc8Re2Z8
m3vMUvdNxKvyD4Cw7vhmPi1Vpd7xTslZV+xs5h4H0p1DrVh1LgtCY3nxMt+izUfz
sdfqoBP6UnCMsCockiOM7rEghWHoYzl31Le1dfyR7IJ8hOhdX18ImBe9i9PDVZjo
roKvEBul9Os5K5bs6Vl/vQQA/pnpUMzv096dQCvxSw4REgllT7BgEsbmCvPXovRM
IQruycAEatZhgOL9D3L57he599yizJxIRFZS3JhyAeeSPVBhxHawd4n5aswVVkTe
CSIoNxUa+HnivMEPIr5p08DJcuN/JmjP4ciiXWoAXPZ4th9744cNxJIXlIXmkhJ6
fSeA1+xCwe5jPz9hwBhkDIS2Y/ONxz9eto8QEEYWtcRadJx4tmdapK0Ne8dX4enX
RbUtQ760lEXy5KC5slK0ar3DUVHAP2tQjiQwAYGHk1mNhTh97Nu9uw/viwk25Xst
ASJkKb0tgCFhSCxn7FNvl4cICZvGzW/ttypvCWAC1UgAIsRWZOjg2jk/s3khbCR9
LGPl3SBBfuvt3P001QtKlfRggJC9F6K/zyychzqU41/gKq0DNC30G6nxC4n8Ddif
8kAaBh8X70Ux3YCPWL+O8WYXBh+D4vOarh2ckDpNdSHe2JkqaHwCfVkjn39kAudq
ljgFX+DYoTpDce/tWxZAsdK5Qc8FUJMPHAdfsEDLNiwTHjo5o3Vz4l3NGtbVa5r5
zTamg2N9wGQg0TyhOAjXSMsYcs7K/d1W2Uqo0zffUI1rVuvsca8xBXCynv+y94Pm
bqemoVMD5HsX3AR6NcDWqPE4oeGAfpn9sjBnt4Bxf7pPq6ZDPVfvKTZvJNOdlked
/eluKdgeV1eOYy3MdVHx5Qz1aKo+zhFjeViG+g3ycQHUv+wTQRI7umSSKgEQJNmv
bXXyUmr29HLpDXRu0ZnkaSKWF7jOnWoMIN+U6TLcWx4D0PHWeGCye6Xz5u9oXdNP
5zXeR8VIIsi9YbqE1YxZ282btwvI3INKKCNUXzSpfAL/2kb6mD4wo23E48V4F1CH
roNs5MOcpw6wo9FL9hMzAQTZBtsWRZQING7lErFKsfOoy+rurScsJpWBmWLhX9cQ
YJNHqBAihcWIGeU9F+h3XKxdTThsOhUsGOqpyhszk4C05DpMIGffAuRfql16OHJN
DiUpk88eIznUQvHg5TNU7tasLoS6la3emdOYhUo/Yw0jJlrFeAT5kkfp8J0DCmB2
+H+t1emyvnZXxjDkvwdt/F8/GHLCkV5vgora9O2+PK7FiMimoPie2DRrnUQE1rG1
FMQ/h1gr/35YrQwvgtzckMF7MOTqbiU//+vJb409sRTAQ52fN9EinDndNWcO5OUx
tl1SfewF1TDLISn0ucIAyM6XSKQ+b5FaeNA+on8TVmGkgIueMwYy1FSnD3RELXTU
IzPrw6tUTNA7XA2QCMls3pjrGGSJexQartP+1WXkNtFnJYP+gTRE4/qMq/LHliEL
yvyXwEKo/dxFpRpxKflcGNFDUmIndC7v8jSJPNCX4KOSz2P0qtfi+wxBCTrJpoY/
+q/ncCIdERfDJXQwF4nIge/nxMDtJWtP9srJBvw9888kDwdXPSUgdOhyFhdDuEW6
p6XmYa1Li306bLBwzeiTs5SMr//bsgf6lVv3KTmj2S1j5cFdKAwIwMRDE6dGa6JE
GwazuQpRokD62FjEOw/2cNDW6pQ2MVR50x/clDxmZWOU1P2Zf5XdiZNW8ADouAJd
C1DKe+ZlqcU5XTc8bbvjRyMnIHhb7deaT973RXd+KNBwkrgZ0jRmCadb1j4CzoWz
VWgWH2NPxs8jMant+PK68lZtyWhsKD6cowtpzleFgYkVCEW/pLkl1XB50cTPw7Iv
+cGR47b2YaYddu3+DqWgARgdLNJCJGMMrkG5HFYrAvb7xVk/HEyn5xdb7kMei92X
Lxy+EdaH3byUeIE6Yd1gEaQ/q5czmAxK03CsTwHdKJ7OHd/bTxS9zu1VVHtT5dBU
ia1JBeAvpQLDLejBE1W4A8xE4gLlOq+L7gdOqul0jusNGN8FeTnnM0tgxCtw+Fd1
+KsMLwjiNNm/uSiIfYh7dDnIYN5rSodGfslLmNh9WTtLD2IRVp7eAL5bFNHvsZlU
FV8dVVefmf/MlQdYKMuhYB2aPFKUvbmI4KLkKHM49ao4VdpyckEDgO5p8Rpec/MS
BIGRJLWrWQ+0PSX3/eYVFnj+lMaZ4azZkn0CgcGtvz+bGBBzkwOcYr8kVQbB6Dzi
yO0JhePsB92NOliSB4Vw67LFp7HWFkbAPUpzYiWWIvFZ8IiWuG5+QeiurVe++mdy
tuKFd8hRUcjKPie0rw4RBBt6+nEjySKNJhQS7HRPWJ/8NsET6rB+V5V5B7LL3IQo
+j0hgGl/joWh7nK0yYjimvOTodBcOzLICJqM/EOXZ6WuTOoXUQQXn/zsexFFQlFX
PXsa7iDdqWDFV0xL84XvwYSMfd+cgwaEfLxCLl/LoMa1HXbvGYEJF2SH2CHLJdVi
s6Stxr+vbUiR6G/swbKxcnxClyB1+y9UNTQOtAbubIqNJ9HHXdOWch+S/Ov9LGmm
NZpJ7EXpR3k4FI6oTqIIcBkSK0/YDC26bstPNFwY9LpVxtqZoJrgz5EVpyANQKI9
JcSJLqv4O0Dq3OkTNXDn5ew1meQLnLDjf4pU+CnK7yl5H/R/yC4jIsAV/Rp8dhFG
VOTtRFsTzldq5IhgLHt20u2VUN8jm0FJ/nzUjYKBbmFOdQlP80APNiY/+qd2j+Ll
Txe8kdc9/m8NJ0n0g81KNIITnO6iP06ve/BE96EKw8iQTvDLImpOUwq+XdEpQiBs
XH2XI4n6Oz8nq7cTN8doXVIXN7ro6pFPg29S4ENqzPxYpqO+gemEhpJylX8YM1DQ
gQwF3k4A5eLsDfofZb2qE7bxiKVQ4IXDPuSR5aBSNfyTuGHLmbbRF+kkfWrecSTp
CLoWY0U9aCQQ36ls1gySHZnKmbhElgbV2rvftuZSEMqxKvB1WE2YsFnziJPSwn2b
pmjUUEaz174D5pjjL4OYOxQtlA0yACl2shGsL3NzwcV+XfDnKzLd5GjOt45WYOC+
9zyHuw3uIduvLoQ/J2m+RD0k2QI3vp4wPchgc5ymKx3/Rjn8iv3Bnhr7kX8OgttG
l35kr2KVLn9ftfXr7H799jq7orMlxUgr5LwbOSr1258EN60a5cTY+xmq6kwgreUP
oXHfF4w1CDQy6j1IxKTvrxLhL+U8jh+3VzwcOI1BRQZnSZPRIloI+fF/A+IrB6Fu
TsaTP0RzlYdpHdasLFbZiYkQ1j0evGa+qfTBHbOyRZvR2sVvHyiPingJOdO92l+p
46vkF08AymUg7jJ569EmjwC2GqEMp0sKLYgmWTjVBxitRFdiCmEh4H/ijbeaLUOb
0LOH4YkBYG1PBhL6XHrL2/wqMiNa8QLQuDoKPSVa1g5v5Wr5zenUnpnT+i9JbdfY
9/K48bDY5+erD3LVu87MZavG/K9b9Hnargd/06wFdRHT1w8E2ep/JW503PeAXNkb
AGU+VSaU5HqdqXxCb/lqM/RoxGQIr3hrIElxIEigN+ZPtLP3Hujmn0QYfhvFZu+B
h1NPWBbSp4ikv4NOJmZYKaJUPYYlPDd25JjBRTFSh0fLrOUbHwgRc4AiFdUFFgt+
V85a5YWGpwFhbox+zbyfHbEcTVlOkfL9LptIg/4liXFDXrA8E0wzgWLK6xXyoumL
PQvUDAt31EVAU1ZzWnJOGnc7qRR80LEkyH5K4Yzbl/rCKR1dHM08QoS+A6CNTUpW
D56u3B6OYer08zbu29DDDNGjt3KPA/KGvYmAc9XM5RknwCZXdyKfVr9oLdfXxgfq
aXVGF9PXBvAaK4llH+4qBZ3jmp2e4n1jN/HAkfwjP9NwDFVb65JBSPpIqtMQ8CvG
TymLO3M++DZuQLdvRCjjuuubJJfU/bjouFdpTlaij79xTBMQQw24ODfiLvpOGC/F
UGGkJG27mD8hRvs0oOTXUyWA3acUQkV7AZ4aNX8ugawM5NqGV7+PoxKdansST7Fw
X8Zv6CMrhemTG0uvaQ1JgtsBcq/fhIohbhUfuzGPj2FfsMDahu9f7AFk79EtGap/
Z0rbdruc/r600bVZKDhQBm5ZD/Yt5wN4GviZTeLZVZAj09ZDQFp0KoE/eyi0qd98
VOeHdA0poUEVyzrHsl2wO43pQj5VXJIzabgy/RVXfdM6WqZnTIbubEt6E47GjXdx
6pBnUCl1+jm0gOylpHxmcPckC3itL+mLvOgxzLYa6SJ4ZscYYdMoXnB8vZ7vDvTi
D5fcoKM1NPVxrHCcBtVyjWYfB+JHP8jgQKHAK57omqMt30hQifTFOmmmHTkzcY9X
r1/jDJDBK6bZjE+WkXnKU7Parl8GTd6Fn0VCG5ycjvgAbIrtc8eeW8kJkXJtepRT
5m0eyEKTxEuCnRfW2Xi6n+qYEvuE4Nkym8pTgW5bA6Rsx9p9PD/z6tAWMtJsR/eg
KR7InosIrS8szwjL9UJNEHteefADlLWLHuUXUYnbtO8btLEB5UmVO5Nyu7wUHnkp
rDSxBlWcAb9NDtW7s7hUwnXMYVphCP/bIzSuvsO2ArQm/UhEE9H5cpZLVrzaVLWD
+gEkUvbxxPJbze8AUQS0lOgi4Nb7EJiW1GN7cXPBxD/+fl8MxWpWUtijZhchjDXY
HpQPM2fr4Uta/TSNzk+KohQQoWoH2FXcepJYyY6kxSJoGApVVrOEf4X8MW+hK6hp
t7z9jhljtjA1eB2pUzVLdu2fZR66DXRRC9tRF9CmE03L/VLmtIpfM+E4VxdFFjq9
R8sSFdagpBSfiQUXO9yFTP8NNzEGRKoa7heWkQElEOjlhR+VNql8jkQ48gGqDqzP
rUIMSkrBhiyTvSrM+05EV4kTdY2T7zjEIPIYXJt6PXx7l3MQWQaFHz5d4iXbU2lg
YWWoM6eXX3UnpiceGFkwfjzj06FzC8sKYMw4AsiGyM5WXKrWUbveFGkxmGOMakr+
AFax1IAy5DW18Q6gW8/VFb+LjYROsEg0DjHfqnbu4dfR/eX32Gky5WX3UDp2g9Ul
agoAZ5SkBmFZZpSkipxdY9myiWuMbcgCxY768wwHOZuuTjfOWDmufe6iBPfog1GV
L7FbNpE+AGbt7/maWHXl2J1WsaNCPD4iereaI+ymyb0Ro8MJN9S40U5WXgM3kZUb
8DcdT6zrnwffJY1EbpCZZfw0gJ+wpKff0xrc94LmUXidA7q2bazeE5QM09VvVtm5
4Fv4B2j7fFBYnBKMkAgB8+V7BldbiwAUI5T0VYcgTk+hISwQCSMK3CbNhUH8sMZ1
u1XhEA+Pp7HS9paeVq3W7v325j/+1LM79ygUZvX1afX78sxhnTJlNG7LQT5IrRcZ
BX8OScrFQF/nzoyHEybd1CYO+kwRVaBq+KU88laaUSNbFPfM2J93ZKCjdQbHqDJq
On7piCoA9twr2mndPm0gGamKuY0lTN9paN94LXUEGqkqiELFxHiC+OX4Oyf2EjLz
mDiuhstnlsZoaGMzWBiKTRVM1vOqF6+pi1pPo3LuC2qVaO/Hk9/ZZyhX549mn6Vw
VFxf/EzE+vDiziTlF7hERmUuwG7POVnw5peh8juNnf3BNc8ku241mxxJru3sDRNd
Et98D+T0q59Ktw/mFs0Qb78bmzMLezaGE2NPp2U6nOZE6F8EQRklely+lyAyPIet
egUtaQsbgi546HXjuE9qftuZo8cqjCeeY6IVjaQUCYiFzEAv302hNuIms8JDaGJD
MfFxSLHeK1IznHpxL1fApOFygY2jTIcJTZ4bkwkcPuxqCLmioeUMbMVSBFmVbmly
k+U8zBCvN5rmkRx/UQSscnkmn7jy14fDboieJ4lxCtRUGWv45wQhMohPh5/jr0uh
6yHpT2x0syjWDGmb2MVKJJFL98ZgyIXVBoKepm1rConu1/VzcflsDnzoEKtsBOdG
OS/cXTwRsTL+Wtk+G7WlKvdRT7Bh0mCJPEVrslAVHSRkUHWQGAPJg9XFIY0t6S6/
r98cRdYYgQpKvBIMO26diCU7VJ4IhhI3eLdxetIScc1uR+3zhNiTKrPD3p5F7vp7
rM30W6jBtmdbzfdEOtcl5OBC/ksTeTTiK6tN1Z1dw0UPylI+wWIpICHY5nR3Wztm
aMAeIIO2OdcR0eg4hHf8JQEY1i7eMT/s0bzhjcKBK4HJBsndaxbomO+cUvO7HvRL
S0tgRjlg7ZuiTM+J5hpQ/vS7/LsacLCdycF9DauNAlov0k6B5jLlduD+kN1J/Bfj
nDoBjABYkznVyNYzsMDBXYxjVIvBS27R3JuWQHuYwnfqkVcD0qFA6B5vl4sadEGq
/OOcwSwLS0MOKv2byp1H/DvXk+kKBVHTtMJ0JaupA04c3ZO5t6uuaqUZ+SolkPub
NUMhr4VJ9SdCrYsBKZvufQL3aD5yXEfG0Jk2GOOIYtmGlGB57T9vEyS+ih3+cp1k
G5Q6oL9iNioOJLr57mKYyLJZYxcRTBBjzhCCdaIPg5DCOkbnPBHbIQwfPyLckYV3
1rPhj6GW68WVMgSsrwUeDcHXTQZm8PbWlocO0DEJJdO1n7HwiyGpmIMOFXpsIjTN
fe/OYOZGTmBjA+CnnZPJx9LRaap/DbvsSQDKa/RccpSdtxDt0oqjUKUkekX6onn3
8byL7ns8K8d1ePsoBktMdAWUULZ/1iho4RF9Juoi5V8ATLIJ+1IPe2xnhgVonYqT
OcinlKjUP9RGoYPgFGEQsUsPQOl3XL0L1l7YlwdYnJFpiX/g1oDFuEp1Mrd4HL9W
VeloPs79MFC6vgV1iLKagmNTaeW4JYBq+AQC2FyFjN5RL9RwyonaUge5NE2STbzK
tmCmFYZ0Fiie8+vzfGV9sDPusLgvUBEWZBjO+eGYBc3uXZzNcoCirRo3wWZ1I/GR
REGGyLrOwt/IhOyjFhyQglTn1Ys+WnZ7+FWZA4fVNjqwQ0HNzQLWP7imvW+w69yD
tvfMDQcMWSHrzqmrvpXsRcGbOR6aR6/pamIejUHYyhrw64vcSbui1aCGgub1d4FE
3hVNTo3CljaOOJPipTrYFSd6TGEV+kreZYVEt+gLDOjUxuROgxqFikuYQoXWUFpo
uH3gwPCwRH2aVuekYXQ6RuLHiogygcAgg14DpAZdl6w4LTgflNlp1ucQbnPOzFi+
qK8jxa0Kv++A6C7tEwT6UcMAJCgPxG3etDzcXKR3ETKHE7kPtbkn65yqkV9sKlSr
ENM7FUvUwIWautm1/VY2C7KrwzWDUk2RiUnkGeEWiAu/dbmOXRu/l1e53R9zmLTb
AIUS1h+ULxdzVhmstOxLFES89izWg27oqDv1M1rsQXBkmR4t8bAyjMtt9LqB9+27
/0sccb8Q0w7dXRmv/k+CH+AuJYP7HoqC2Bf7TU4A3gJ/HbBvDvs5EtTOcPmwQjvd
YCNUTRkFXV5amYSXqMgKcAN72GZoG/nSTf3unmxMCpHfWItarlW0W6OS+ghPNwh4
2bYtmqf2XuuBiNtp+8t4qcE4N693oW8db65aJRdCC9qgCCPKwlOa68XLP3md/VVk
33wGqqKF0nrUdNYmEjW3m9bcNb4BNP4bxAPiYSAVrOx1iN6aA4NqLMHFGYsDDUSb
7JhVCzBPs9NYIaL2YEQtIzN5H2fZ5ZQCW1W0mtNa9s60injDZCTF75xujH/LJxRO
JcwYpk6KJyN1O9fytr71Dz6r/380LZw0N1vuknmu9x/TiHeAKc2Rv4O9uqMtzEmu
UbSdxAloN+KJpMfV7YQMfay0KOtvl/5kRDUcdAxd3U6AFNOD9maIuKLVpZk3QWh4
1Hdn7hCaQHtDEFtZ0E6bnBNK7gZTOtCQKDg3URGncn/I1aarK2h45Kk6t+FUKhmo
8GcYpECGMJK+a6HMffAreK7XHWSkzcbzPa7encqipyzRU5P5cPA8iFi3CKFfGIC9
1zq7GJRg0BC6lsj4eNe1FxqMga9ByfgmBhGnN0m+nLfjWbXevIbLPoeKQpR+TL/y
/fNCUskIN0Ot1cIPIa0SbOsSxwluZIYIVg7aaUdJub4kObyCki0zMWsTbIIk+jLR
zWBqCjyqdvwv7sXmIIL5AlI9STOlb2vOM3wbQ1y783gHOC9hPaer1A5visBj3xYk
ApyECDUO/tLFZ90p0kO7FTBVsQ5QdX3DHgXppr4xsutQ6ZIXNyhH5w6IGWTLTQt9
A6iN7MaGBOj3+WimHnQw7j3D+HiZB5M5eHqpnrWvV6JH27v+FrjP7fP+DIJ+cjwj
TCkdlJ9ezgi3iMYb553CugwBL0lhA/Czlte1XprKsvDqc9Ep0o/2CtW5cYU+9Z4k
aB03pCZlIeP1Bc6LKCMDR1bZZ3BFo/aL/KY/Gd/E9Y8W3fB96YBagOXo4xos/57N
ICraMHNoFYGJsRl4f4jGywXcwWrirZ6oIqCfrLu7OQX4LfFniaoyPYbGnBO0qm+J
IUN1EPDxZQs5c0jieMglyhWz0p2WF5OM834ZWiSwOfjjArgDJzjPimaUaTCe3DWG
DRPqQwZ1PfqYvfCtJ9+Eb8dOUqQcOBKd8gB6hFed27Pl1BPBAqBI6WTbsPLmBSoP
Nt0k9oyu85ogQMP78v/ILvXYDG5k8XrruuZGp2+GmcPheJUfA/xC4OT1wDv8g3BL
YugF7B66nXCTSd0Ym5J0bdcfmUtfAi5aieGBHGQHVo4DqUmZz4QFjJesRKj8wIt2
YcICgscXTgf9LGkxhpuKSSh0IFy9zB/pvTWrLsm0mveRFGQBfOgXM/8OCPEiQk3i
9hVftogbsdVemRhyUiu+QWy03y+owPlRHljxAv9wtcJ6XtZmXyR25yQnKkQQPXli
LjnGmb41NRZURJcvlTi4gQwjXFY7R2awP37tag5ou0QSgEXDVtmPz8n9Y5AYYDUg
QAofQYUW4csIB1XCks5ceyNeaVmIPiH8AruOaVSXyJMI2o2gn+xXEb06NHVteZmD
o4uPOWqYT22m0BvZaLy2qHRCmGkbvpzuI3MBXBtI7C5TSz2VQdz70HnshUVTaIiE
b/xOEYnfrUwNm9A+QvGr/ekbSUW92HIST9C17+bUrvHU1NtHqdLGxwE1nAsqSUnl
20AFPXClBXA1ux3AmDnn+SDIZ7IMAD5xaq6Oz0Cl+lmiS5ifM8kR3dx/YCgT6wwu
FQKMjMEkH6MxKe0Z1sXH2EQi9PgiME/af/ciSvQ3SYydwyIhqHBaVBAX7blPCXNQ
8KH3749F+Jjus3obezzspGHzu67xWujnfYyi8Zmze6bcAzDeZGrrTLBg5yYbVPRc
HqNn8eUApnaX+T7PabyKoSv7kFcu1iz9f6A4ac8xQN9EtPHnZWRe7cHUQTVlY/K2
OSpRXFZNARgJuUQvnUGQS2+Ljvkfk6pMWoi0XannGC1/sppulqU77874zb1XQ00p
GBrC3vQ+pnrEd64xUHJBHiOD96FmuQJkHwGIRkfSO5LtvqS7F37c+vhUxG1YyJ9I
bATkWGVe9OI+2j8+u36tvawGEYKUCCt1oHagnJXgAf46d/Rc8qPooEI0tpqqsbEi
1ZVCd01oSpFIaz/QJQH+dd1DvR2mh9mGRT+6F19DMWkSpGY6m78yPeVASRBpMILR
s1isj3QDKfg5Ur6YnvDW+G5v3dMc/xNOwiEL0zoGBFLBPtp+OL0nJtt4P7hSpRc5
ZDRgksSfPyTsfQEM4N4N+jkBEKlQHrP3BalV0Xa5dhg6gZx31J/4odQKJ8LkJr4l
Vn/+ZnWHiJwJeo5RKxJ4t30cn/RY6SnQH9Im/7qXDr3kJNi66RFS14bWcsMYZRba
2rX1o+9UG8mi9cN8UMcWUPnp5RClFodeYOYRKg2DRJux7B7APoqVA8xuJoJgjx7i
LrvIwQAFw3scs1V3zH+V2DIS1bhIR+Bw4HUWbg1wt0gPFtfu9EEVQ3CZXf79SWhF
0YKGzyj/b59rf+C7S/qxbwAhAXeP/qnRcnVMXrDl8u/YLdZugaIMOAtq/JfBxzVm
tZFmJCEqEHnl52cCTj5N0A1Ku1HT6f6ZPWU3r0dBi3qP4zyzz3tgLVqKMSCe4/c3
ARd6x/Jm2ZBG2aPxC9v/luKh8/MmuXGwgQ2daVCZcgyf66wqqS9h5rVm7Drsz/pb
P6cnbPGCbHNtNIvADBBBgS+4inbzF2OxzulN0s5iOqzjqF/eJPezWpkr+/dKcviR
sSTkjSw1MfF5AGe8jpn/ysMhkimwUgR4SgapAvXFGd+/paXeJ8jGkVRVCogonH3G
b07BVOQSpgg1WTePnqcZQe+IyY6+sw02LCb4yAH2tRdkO9/VjAkiEE+yBmTbPI3D
OumL9eAkoVlZRi9fb/QaYVGikFm09kJnWWVOYf3F07gYlguyIhWrziTfX5ap1uOo
LwdMriywwmk/fYXwKBpFVRrsJl1fkGxctvmx1ZQ41rHUeoFMIJI+nFPes1JK/kjn
c4+PCbxkCQ1EsaS45kDxg7aoi7NNi7dCPoyCeLPLLPLYse6NsiGPBrT5x17W9je/
4odzQXef72lsx2Xb9Uk58B1d3SmMFLvxUQ14Up7LFobv49bJK7VxSWtWZQ+FHOyY
rmxFULyj5lm0lzBxyXhy8yPXe0PsaDA2HZ8pNJXQGuEx+Nkqvu9EBJDND+iakbn9
28VjpylfNZFlNV/CFnfWYrvSrW6tBWqoeFjMdrFRy6sL/NspBqmS6uSPf+Sps/29
RJ0Vit1Qrs9dEoukKnHCPU80B7esYiSw2rwChjFUhtstOyTHB6JTYLtY7NKljtQD
Pq1PguC0+5ShjfJUHlkdVyvAVe2ZM6R2HSQZlwL7ZADId8AryKioiIhj58lWFS3K
q7lYSgS3WUL2oFQ6I3vC9iqLeEa3pauAUdLJXLOn0iPacYk2XoNh7+xboTSMr323
LW2uwUw20YkbKpEjKJFdVRoUs7+yByWBF4m4KBIjvChcoKrteAOZPmZCDlQkbn73
mo6UHdj2ZFPRMXDtDJlFmfRwLW3tLNuQUaSfkAOYq8CrB8veDW6QhBY1wVG4PWsF
vl6immbVXajtSOjiF3sEZ8n7Wx3k7FJc0/FwCOKX5VhXACUPOJl33gxBRMmRWYqN
T1Qq3Ab3h5DUT2hR0jmPvaVR5VDIyWqF5v8PpLAtJd6uqa655H1q+jCCOpgGerHF
dInZXk270/9DWJuLrQYzr7MmoXG7nvQJ2h2QeokpRtMcEe0T2+V5HVIbzQHcpJdw
aasN4xCmC+j2P7FyeX2UdE8i5wIlNCaFew6wDRieqe7lmP7hF3pNB1D2z+vQkf84
IMgf4G6Z1eREm23Z6gh02/GMwMiosKYflX1lkq+cZB/clpoP83cLZg2coXU9qgPT
ZqFCaTtYBSPzwGQ6BqhEXg0QvFR+VrncgW7IdriL0Cgu3EgdyajWF2KVpV6s6ku7
QTrAIMwZ1RQtuYqGbVk6iBYifg9OvZuQI4GPJH7UsBje+jAvvOhcSIi99KnX5YqD
Z8sYa7T3EtR+tlUO2VpXqwE2DrkTDG89PB2TFePfs1ysSTe9OOzOZ+bYbiNCc0F/
detM03aiaT6tVw4rkdEGFleNarlnuW3EiTCmgYd5xYcZsRowSbjudDg/4hZkW3yT
y4YZSqwqhqYPppdPuwMT/v7kRutSyIRMmykaNxuVNyY3NfLnqgRAgnp/tE7uOTX8
CyOxJ5yKxcOQJUazTggvy2jalZFW4EhbluRqsXN0rC9c23j4lWpBnVLMAulGJo9V
p7rwgBJtLTopGn1tCsp1nAcDLoTpn3NinjRevVLqlqwVya9COk3k5TzqiM8ST57N
cOMWFNNPPWxq8pbGimiYkFgU+QpznRJNHqyGdvP503qtKzrXMj9N9NzoRVkaIuzr
Q8D3B/SwOdJxGfcdRrtPmzP00MMgdOx6fRQE2GriuK8h1qv0+RypKV3tJa3j7jmQ
nnELVVA3QJKJ2KZWDqyeBrsfdC3ldi8lZaXse9w9J5bXmRCcfRH4ZYb/B5uxnQ6J
BGvLI+TopJgvEWV9tRavyK7eNJQo8xTUo17voyY4qNX8X6Uj/mfZ/moDih2Fs6T0
QqUq7rh9XQwWcC++fBbX28uJyZodgvlGlgA/6lvIrCtiHqo050Sw5v4WtV+u9yMn
q2nAl3GkFXiCXw54DQUosGEPMQPcr+Qh0LK1dutsf69FKekA8l9+ey7980vB9UWF
K/eYm+SjjcrPDPi6FDsASAycz5gH5JNOVo3Edko5LLYLUT+86Nt5Jnrkfc/uOwP1
p6glWMmk0fenbXJtaxEjUBFEkiv9z9iUmc55VvTiIdJ2vrJYRe0ueI7EmSk8uHGW
PgcJi+2ooFiGki+IMeO5Fe8pp5wyeOTSwzjawyuDfe2zPRwzSqNlYHWhxPOECXsP
MLS6MwXjUqcQmaT9TQh5+OEIhkDLqHnoE8wiUooFuwDQ82y4dNiN+4PPfZfXM0Lw
KC4muIwLlL4X7+X5RCoTrawjrCDUY9xvVYqg2XHx3wfEmeIyNlX3eAXOv841wOrZ
5aZSKFFoHtyKFLo6uG6pE59/aeieYbhN+5LkKkn0h5QsAEoNaqrXGwOQ3jjZWi7H
aMWRjVl5woUZrTweSlEBoz9wqJfT2Nq9eoY2E3Lzcd8rL52zIuashUyi02IQbYkf
4mAqzjFdU4+AJZLq0GDv7/tdD1Ma3NzXJ3+by3IX8jcxeLfgyivAT4WxA+J9cWpJ
XCGThRI4dsAU7LRAR1c6o5Sokyj3E6e+EXzoTN7bYrywri7ngex80ncUWF4Fo3kW
e8+90m4d9XXSBmATVA1kgtCbCKox5VK0Vq0nv9PGIBac1hZGdvdb5kLhbdMXMTCQ
kb97pzrD8MLEQfq0a88hVbHDJfHg73ZctklXNLYMMRP5mbLucDyb19Sps3QhDdnX
rnKj/ZkGKuH46jg1oMiCsODssygTqb136oK9TPGzhharUeaoWam9dUcomCq5cfZR
yeYdaXT89DvcHVPLlEHLFbAjkp66ZVVpdNc+sWNZF1wBVoI6Fac1NUK0HFyEaWVT
98mNYUY+7KZu1Zga+mC7pfnmwzePvLo6W4tEhCqImh9HImLH0mU7LTNBwsCraf1M
gLFPOHf1UBFJd3cJFtjcnBB7wwBCWiz6dsgpuWtYdgXLTO8E22B5mxTBnpn/wyuP
PR+hwVv2DlOZNTfsBH0ioRdTVfOEIuk82P5XwKY30krwLAPZlMTywC6nXhNr91qD
Xgle2ITIN4w/Fd/8Fe/IcLm8blyPsUh4V7GbI9MGv6vpeZZJgZM21XJEn1MfcEGZ
XgUSUYOcli7OuNIyePO0N3+x2kezpETwXyG+RJdIZek8bwr/6w9AKxVfDVTR2HTY
/IehPCzzZTUElbk2+KGmyb92sLeoi0m+Z8bbSkr9LY/CicAj2tlCsquZNE0NVkcz
m4Vw0mbPQq3cgEn9avMyeOBLN0uJGdWdwHKldDRSY1aXaH7Y/3Q2O2ddU4rMFble
SG6soTYnpBULh5HTljQZCrkzsuz2VpsaaqFgtt7iW+YZ+reoH330OxZUAmkpxUTC
aYDEftkyedQvodfXWg7o2EiGsW8K6ilSYx/62FUxyGTfIBhpYqOOUZZ9BlN6rcs2
gNYueZcswxDBmdZJ5w6IEl2/KGlYZG/gagXNoj9I3z2nH6tGzXNf465PuumQVeu3
Boqkix88OxO2JLsuTWWwkLUqI4bgT1JDErgtSXXpfIOaoH1DJilmUr0cTMrV2ehG
VGnxRMRNwU9VKwcBclWMc+DptiDkvms4/WnO/IM+OpHccdHnfJaCANBXTHWKQmHo
skg+YdzT7fL2eRN1akpu3OHp+yzO7LuxPXM4IPWgwpHbkOhGECjxE6RIh6PGjEpQ
RQkBT13gJkyOmp9iq0PiJn51IDR6w+Jlp+Ud8JFpNjvRv5/e/mhEE+CY+GoR4gl1
UL6PWSX511KZ0myNm78spMsIDudTJSSbbLOdi+V3JnV+zNirH8zazBJ90T6j+83c
1WU0mh/nWsNWU3AnvBfXp1phyBYNwRCTHTlzSdtEcJbZ5qhSO3DeuE066i+yGdWw
tnj1ZliCnmAMZeBaK5YUk0yOb+xiqKtXQl46VbmgM+XjM/XIPDAfAlKMOrKIZPIB
T1RqQswO4tBoem8rvJ/wHuykk4TdQhk+0I/Op6GZ/CLggZlQTkrmPGj3CM7NnUhu
Z16MbOvOJOq1ARpHpEtasYeQTGUNN5ZSPuRhcZZFYFmuo0GEWZVZPovOW6jTLLGP
KL8cMoWef6x2EkmrBtVJYxAxYc0QMZMIe30lS1xL5JkZ/Mh3b++pv+x1OoiN1i2g
8ZBt+OZU/5yx8djgPocUIk0ZTMEpCPlbdTz/qMCs+WgnIRw2D6zGPnHmi3QWgr/n
+Hk4tUp3Ly8mL9J6kW3TyMFTaiDlHH7l2u+8tR0UngmYxSm7QOnluwKn7J/nevHD
lZyPuRgcd4qjg3qrU2988DIIq9OPBja05r5LuiXekw2VdiMgKbPHfTQB5GlD146+
YEN0z8rDqVceBgrrLHJ+qHTL0HpT95u1EOCSVHQnuPeJuSi0IAxXR2S70LVO7yBi
VF0AbM5qkXCz7xDEW/yX+tH7yaDlm/hpsO5R/YJDkI3xnc2Fqxqf6a9HYGJFVrtV
yVH43CbIlP1BOpXXrCf/I21W8DLCj6QzUn4tC15Xy+0NT/V3fAyqmiRag0Kx4Ht2
ET7AEhdMyUbah9vp2oY9GHdS+z80lX8DckyghHn1G9niNoKN5yGppznmYwYsxXKU
PA7QfSWmKiAlheogI8AO8yR4wKFFeWODdmwoF0Z9lrZ7belkK0tKCViM4wg+wvk7
w7cYWsI5iTWnVQQv5TzusN4+LBTdbtUmuRBBAElBKtYF7zrsqf+G7wt7cUwJoDIK
DZBGQAMqWZ0v9XiqdUaD5idDXwhxv4Mv4tJ73wwGW5RC80mnVHvjqQAMgwTaGsni
FqZPSU9gPzcVecL1H/cDA0jcr11IW5s+P2P4UUO55eTY5f7mJY6qGwNHdVon4RDt
SdkUFHq5sdnz4GT/5+jx2uBVRTfgTs7CEk63igYSDHxu79k578zZRxk2bCvtC0nv
rTxrHRjXut9fXgQVNnu6jd2Jga7RTkswWKGWkbrXIMxXgE65Q3fwGX1h5rAdUBYo
5Q3SdMlEzM1yoJBJNr1PCJc6uvIdkh1nf7UzCCXM2QPzSXs70BjUmmdKzE/la3py
FgJXID+lIp8N1RCmdDI9ywy8nEx5vWeY50FOtaBtlfnjBVKqS8TwUO7s+GBG36gi
DrQS5kE5a1HDp8rge8OeMmZTMOCE34l7GHkJoRlmSOGAauZeUm7jBhsrZafODXt+
qGoLF+pU6/HUjPBSc/XqUeq+DZg9PBCVhtFQ0LtWFJGCBnUGZS6f+JfD0PyKowE+
Ut/y9KNhQfbGbsKJ/9hG5LUGMq2IzG9KyESMSTVkXOdK28T4BtRNQLyU9AW3IDs3
DCjL3UZOVFBq/ouCK0l4LCKTgMMkWVoqtj3otroEOJ/noIb/yYR4Oi6nqGbjbZfM
ddyxmmYZHODlayEL/4tfPAu/fiy/321Mf7SvwzdHpu1pRkgQXKStOb5DTAXwYNIf
1+jUwZ4BfH4aHa8oNc/8UKTuefTiBgGV7Wgu6znWhDpF+/bwms9NGaeHGOkbrHDG
PWAWw62Wy3imTc+L6vqvTnirsNS1CpFJBBRoRqjy1UPj5MAIfxurGLRG2sGA0nk+
F96cGFs+ofM9Af8aNgx4cZ5lPe2KyfdMLw+t7nGumV4XqCs6Um+bX9cur7n+pU0y
1dmxdr2OynJswkXJuPvMNHlSADBgWZy5+fezNIgkab87hj9Aj8oOtWoZTo8MRe3h
95WZcuSjAY9gpRLlP8RIVuTjfoFKQM6wTgG31Gwhwk3JJ9/nFQtXTsaoRuqvo16V
WhBHyXLBfrFv7OQglQ8vqCxMNoj9HSsni0+ZREVWYoxrDryRYJjc6iT1OPNwiYKw
Q1pB6yh8YqOWLLSUmLcMC2CLfTeUMOZ3SticAYmLwLcOzxau1SRrwN5zZXnCQpUh
pghZQD/mDbR40h3WLVKwd//2CVvIz2aSD1C9pY1FqzNtO7jDGmkyWkA16BTyAq5P
Ar3omylnRBYslDT9IyWCt6tNvs/Ua6YirhjTjbfdXdUKlV9wWUHuNZQFSL+Z4T4i
UQfWT7pXZiGjh0I0tBtULwgJC78IbxM+uWJbbC7fLkPy6j7OktxRcI6N+BmPJe0q
KTiZ2AuDxpixDcA0wIQUrqG9NazikU4O+aB/BOzFIqsR3pR7QEGjKkf4pP17kC0G
zQRT8dSxn8G7rd8I4IPm3RRF8V+QpOESwWcgrByd9WWXy4QYnrlbeRBab1cmnfjX
Y6kEwAg4tCW6WxicnqGkrm9MScTD2ToLj2rF4JKo9QRGaT2QUsN1SNM/NY+oceMv
NMwhwc6VA6mYJp6u3tpTmCkJwr05sGB7LnypMcbejwg7k5j0jOdho5yiJi499nUx
2huBKjA8F4LicM9CQEqrcnEYxe0+ssQuGAC4A/cF/JChRZu45BQ5EEI4fu21Hjs4
HGQWpwJ+VwL404vQQ2u9Xw+b7q2OZwsX5yreHDT1Mqd8Y/VpZNbNCo2n0lkA+6SW
QK0w9dp4sA6EmLRHJ5d9JNWjDxa2iFH/E5gfaDPc7mvNLjzUXu3p0g+3GTh/kOD0
Hw2QVFsdvN8PzVlWG89kaZDuFSK3DkoIbSoUPYiV2vC0UgonWQcWGXw7IEzNk7XZ
fGfthK+dyQl5OIWSKIj178B0bm+EJg2kQ1ko+KZb4/yQoMYM6yHhR6yoCxeiFuI9
s5SvVXFA9VVGNnRK/belXiTVgMGHaZFcSlS+DFI2DZMaWBAjDmJzruGLE1m0CD5K
Cp89pW+pGCMGOapCSD8rnDsNtvz4ZIxyFJPRZG/6/BY15+Eb8kyutvDjpG+OgM6J
7RagU+uy4lx9fdzaUCTtW1+L8cmBd/+PfEyDmWG+LyYlqCw1QNGh5NmKH3gLc6nb
O9G0cRG/1K5WeHzsYUyHOIuOhI2FKk4Jegtfz4w9m7VgYPe8giJDjCMXbdiVvv8n
GpWRJD4a8PiV/23W0TulezH6ibiHBlmm9LwAxGOAbOZd3j2KyHVlLDmlUT8hMEbW
p6eJs9y3bppNeoovd2WcCRg0X4VwNcKye7T7BbyXhGFCDVBE2yusbOy3b86j4yHX
OxYRAYkKSW26x6ch9+ZVmK4flGDjyeFXj2OI+kxl5iWEoMtVezOuRS9zXJKD+2ZG
KcLFwMdoYMSb0zvGlQKmurWmXSsC2uaoZyncB3krJ5CQfghEWTy/l+SeCAEPVcAa
uyuweh1z3m/g66TCWakYljBY7FEYJAxo6b1sLnYVd0sWhYyfS2RLjR7wM+UHLFjJ
5CRCEbD7Yz8ocQVx1A4pLXk2f2tHKf62lssQ2V9CUvrHuo6AWAtJg7Ptzj7Em/Hr
rFFMdiw6TZAlww2rge/qXP/VKMQygjLvMXLd/PXptmsvrMxsc2Czp6gRNhYP6d9L
5jmo1qkq0X3Rzjt2qVOVAXQmUi0sewLl/v32RpGxiOOabtAbBE7CGZHaq+ESdVUC
XdPAeievLIjLxzEQG2TwkhV1aaPTPse3jCVK9pV9bUPLK2j9BAPJZDnTzyo7boGX
T6PQ0IhFlJMcFO9/bEMPwlYfjlc3woFrl78P0iuFzxkb86n+0QryJEMWGnfGzjR7
SJ1AJ1nVnpDCOO4Gk7Z3Sh5XdbjVSAj4bQRulfWMahH+cHyzW40DHFUB6vXXljlK
ZiiM5Fns/WDqy1JT3Ilw7O0c3uTt/m6FmXuJhqnULZKlajY0RUqHhR6JlDdYCjZf
J4H+aRnSlOVoey1L1axI6wDnga3gb2sFKonYMVm8tzVXFsDEq/5vEBZBoJAww905
S33nS3aBdeoNaV8xN8cjSQLhE8QWwOASI536/QlDoQ/E1kXbcsPmFWPlMFk9hW+G
CwmUM4LH+CwloecVN0g5kkBw4yPurH1VFAfEUMtVJdddHq0RDfkIy+VHjecO7ts4
7mR4axuRUlBR7n59Jh/G2yBCpad6Ul40nyR8+gHM5dcfovoPKnzdLc+fH02owSLe
D1BYkByT6tuRrWVfoMU0KVPyQEU9UhNDje37uoEbA/7hNiKWf1tF+ccg+KKFoRZU
gffF/Es6wjF+tQB7GrQuH5qMuOaPScXD7rT9oTmIhgP1WEhoYSqJN11P7bJ3oU6O
x4EcO46WBRYbN2SAQb+vaHmZ5DVipMycMmdp9OPD7pEit22VXfvSemotzd/HijcW
FRb8XDun4tz7cb7EhnuPzsi16CiYrE/Xqtvgo9eEW4CGY7MWBmDSq1sncqcuXQC/
7/wWNR8+YXXXTfpfWOS6RjG9X1Gdt/J0oV/W75H/wYwUW+U8ySywhkhUzbQecEPw
3m/blsg39nHl4pNVftw5zCACAdbDz7WzEvU/6K1cVddTbVxAFoIwV7riyYq2eGlj
r1JQ4qOblJ3L5J8R0eZGfYzHGXezFF0T6OabsRnCNBJr+d3q5t2rI2HvdcvlSFyM
9w6QxOzy5DiBKIHGtxX8aQekqfCGujL/Mdg3EVlN3qG5cMPx1lZqD6sfA0sHsWZb
dL4wo6aq89ZcOaR2NAwh1dF0F+iaug6XLXoEXSc15NEbzo1hAW55txa+YZexStBa
fzNcNygVcsRJH9c61zyra/1v8uXl4hZ7cMReJLVrUpGZhQ2TOJXJHH3F6L9/12Xo
nLwe3R9QbsrmN+j+n57Fq/U4lHgP+so1KMCzITE4E7Wh7oydQIahy/u/KIDlIWax
AYY2+57gu+OUFlkLry2GAodN6ntqf761UzYdFBPlcGItdpM8egmnCSCD+BXq/Vop
43dg9U5vaqD9ABXlK81ki+oiqo2ruY6qURiMoX6+njp7cgLVYvZrWkmVW8y6uE4D
jCsdGatj1HacS3WBnIQpQCLO+JdHYzPBNeD8LWRk1+HnV1QPezMlHBiGr/i9DRVt
Bh/AY+Hwq2sxSivlnrRei9yo8yHs976Kr+Ta0S0UaiXAbesIBXBuyfVDRBifmDAL
OHd2ipi2TZg9pAWlMAEPUrSGycli/3B++6rBiPXeYfa58idFHCzhh7tsLarWdzF9
w4iEu7iGVcAocj7FgwJMVsgf+oR0F6RH9NtD3+mvF570Gq7ZdASPhGiRYOVFvEr6
AgdqJEkQhrJGlEKRDYj8T/9n1pfmFFGzFY9hrzsSIXNfcg5NVIvwi0EQeaK80Why
3dRtV5RPxWh1LRuE2D3NDFyE2IZdGnXv15iHYrJXZkPqGL0c/bhbvMgk43BsvvkM
NDD0liG84hhfvRLPMDfuUKi5gralKXa2ZSZJ41Orfq5n+n4Cgmk+OUCq1zG9P4H0
1ZUbeGDOabjDkCoScHRbiIOGisGMSz/E72gbSXC8hkJ20vvN3aik6zKHsWP5snSP
StGqINiugmvlrUSgAlX5iHWXHpzd+XNgSVVFA+vZaa7l9Puu/k2DnTTozu0R4dbD
KgBFZXNi8wLKYmaPgLkmGWaJ3xKGx9pr/VeYVa2r2uiJgaFvo2lfshUwdzQKA5a7
hHW7LGBdOFFsa9VyszaTg1IK3p7h7oQFdY3wvFT2V10qM6EmW7Q358s98N5pEhTc
UM9rdnf76Z/qp4vflUBWUS6nsNW9rjrjJ+SzKOzkpKBrb2NmLXH5T0K1VkUV1fcv
32dfMqm60lHCGH3i2lmIrmjh5YT/gTqYE2WMwcztNmxwe17YA9NG8JY0IN5AgQjV
wOCYqlWhgJB55YGKJhyFGbAbBpJj3NNeqDMg/IvaGQpG1Nl4Q2CluascHYT3ulVd
Pu7Rce9q9Oa6jlP2ekJVt5iJdrxOTFdE5oTbiZtYPnhxTJPGQT4y+RNTS2lOTAEk
98YVeJSlugVfuYjUUODU5sBZj6jGsY7jeSPelI0nzfEm93KBwyPN6W13UzBkApZT
1yDk53GoD4dxSC4K5ECq02KN4aP8a3A2/+nOSCyYXz+hTAm12C0Rp1DhgLYQyxAB
ohddNYAHTTdnOkq+xnn1qf4EjyIAWLKwo8FrqRtH1Ep9rnChjYIG601zvNC9iLrV
egBUH5MrURcWW/pE8fOAMBCOGyYCb5QjF3BLJyxgJiuOdwopsyMUdQuEwqf2h0cS
JcpYm//Z80QL83hVYUvyZPEYxzIQX24kRzw2PjNjK0MhmBF9vVIioD1TIy35hogw
Bkw+wrHSfw9UMG8PGUpufqceK4j+ZfXaw/N0pT+0m2nRBuru17mLFFXfEsLaNkC7
cd4SmGl80jsn9lmRHoMk8ckpctQXvcPjLj0gqurNyVC7z48WUj6JkJKD/4ZfzswZ
sOpfIbwA1kAV81YlT3Cf03nBUo7XgyuesDvMYbjpxgtzidQs48r/801NvUwNcWNa
IccoQaRsYp45TYw0mrmiNlAoe0gitRkNbVKf6AMeyaN9AGmf/mZghfmv7w5oPHXO
i2l/JUprILX9YxnIndwsnPeKY6g6KoSLlAGpTpHk02/baNoW3G5yityV80mtnrlz
MnNjNjx/cQzAqIWzwmTOGTi8suOJbXbxSWOYSIiXqHSy7RMHjsFfhi8hR4S8O/Wd
XeGg9KyjGVckH4zPZoIXSLSgonONMy2WdG6IEfV1Hq+e64OJBa15nFUjg8gR+j+n
ZBBR3wo1oa/TZpGkoAFM3wr5rUIum05zd5R+MxlcqZ0liRPjex2sC3xkQc5vw60/
6sxX/rWxb+hmcUoV7xGiGwOagw0let81BNwrQzqlVmU3sFl7hLoNt8b2E1RjeD4i
TGr69iQkHif+R2ddENIDd5Xy9QMnI9q24qjD2xKZjpvi2sHRtOjOIE4nefPcVred
GoieMwFTxWXxVOANw2ghYSg/f6tGNVaZQHfAB+rbVjT5YaUpTC1QBSye7WurJ3gH
Y4Lm0CCJ9dkvZ15V/IY5ByGgtgEiCcTfZ274ENNTTEH90PzdokkuNzAQVyV1gNvo
cE3ibsCAtRfLghrwER1r86e+kdVCH7opI0yBl09DwpyMWIMsqMINNfPYjZSobda5
hVjiktMgbJL8B9r2xSTKH83zToroWQb4XqYBXvAkJmmHKoJ31TpddFisE46ZwQ5r
rNRUdPjne0w+5YCYaH8cXJXqG1PG5Km9+rQ5PJDKfm8xKGYQMtvU9lKgIBTm75L6
lKBhvp9IDtTuN7miJh7IRJaP1MyYlpLcY0bUVP5aCgCGdPUMLZtLSGYWHXr1rOIt
2nCzOqNQ+JekDEBNk14Ry7iAjMADlbpDtb1gR2PbEDdHfsma1ffBXAL7DyMwWLRB
W0sIFHBts3OY60nzh/EpI2ww1I8fMu20cVMcMwsQIFtseRTYyl2bbAe1xeNu+KI0
6M9NayFYuxkz5T4vZSVTpLVSZEa9z/0Uaktz6TNWIyjDpLrHP02ZoF7xC0vGeFlc
nPKqIPvZTZEu36jiEvJnzogkOIV+QiPN+M8mofqp2tSWtKmcbS8cBIqajBzF8TCO
ud2FdOjhGO3FAdk+gGYg93BOxQtdgfCchBNsaj8hFI/suRDtfjPNuP/z5HMPhgD+
jCaAWUpF1T198gvLYU9G0/4f4x4QFN6Xv2kT/334S3yIfK5X3/hatZr+5nNBDnBl
WxfNB5w/N/nTXqqMjfdG46ocXnImPpRgRI4RNEp0DqY9p+Rsqg6PUDvEyVtEG2gS
XegGAxnXpVNsBkqvWEY3thRJeNRf9EmPistf4WZo2znUVh7/Jhvxyh9rARm+Zl2J
cqenGWZlwKN2dgu3VEaS0DBoQSW+X+ewjXWjvpM3WyzUndlElqGMtcnyn7mhqnRq
sjXIiH+lLj8tINuamHbaJRKp/QZ+ZdY6vOjvwu31eLrG1JWGihqDoe+051rSio0Y
ULNNjyFMC7Y1JC/F5JPptnvE3xQo8Pz02ni4/tAJdpIM3k2DhuAnzu0H5Wsi/kLM
drH0K/KuQXXY67xLWpTMrAGAFaYECSv877qjL+f9t1q04Sv+zq4+eC2g/3c1eQQW
adT4gIKB3ohm+MVdCeD5DzU8Gm+c4lOberm7MpuBZGpYC2/BOiWa5kRgx+MvUaUt
mOKpbsVPianPMhZkr89Y8MlVMO/n6nCxLdliAJEA5aWFuuh3iNq5Gr2tlXQ9VSjS
4fk8eZ4c+wrupL5tYrfgN2DgjYOeGEeJa0NNP3ghXxPF9Ftt+TVryxSLZLoOJD3f
TFCOob8nywcxSe+3NNxiFKmjzh849mvQEZT5Q0G5HYVW2Dz9b6MqaDM6OYbTBmln
EiNGqFOoTQRvjNH4v/QocaXYmW4H7eeqLpx32f+D3sF5GCYqOGJhjVG/0sMdpyOF
PE25mkiChiPl2PTVMEDhDJKc/ItCh/oiLaamV5UnP4xzwU5Cptr4Eu+zYleZDRxf
yDtQ5agknTNp+SHFu/RlfYzhxaMxYe/IQDYuB6u9qClTdAOnW92WEba27/20MG7j
+KCWRqUjFdvWT1ld/TRUBD4tSgum13epvYEUxYOmKUoqhhXRrCWcFd5SzoxlwDYp
9OIAglrkX0XxE51vpRtwO72EXvI2vcR4TQlgoIBvtRjrFZ9YdTLWx46n18JsRoXg
Oaa7x6dc1sYUhusUUGgL11lUKJgU7qcjOx64/gORboNhqR03D0cix3AQMqKaedDx
Ama9PMJt7S+Ew2VkzKetIZoHF86dVMtwZR4DI6i5RIZDpPA4geDlI7AcuxsOTXjG
RKmBXQsH4WCc2x4yUjJ5sVHQAy6bUXrcbgoXjoQfP4Gjx4e09jZKBeEvy5hEGs+6
Kri40aq1imQoLyfuMxqn8D8C3D3IvK0nM5v/7UsZo/rxiPR0/0t4bAy9rPBjdzP2
Z3yFdRvbYC3+xFLiKue0L8R0/+c66XiUdMpukjK0OhRI+VIt4TggzwHI/AHT1at2
2lbIWNuznz6bznCWU69uy3D33HSDzfQRUInhvXG6nnky57i0NG4ekdFUsYAdM9j5
i4+nc2LJROaQZt5LKUtLjIMchbUG2SGlkdiKi68mWoUbg9pvfXTE0gtf45cLKZwi
qkAr1TOEsTMQpt1baRmPWacfzipWHXsK8JJBLn92ZqvRmPjjIyM/89wwmiZoY120
PUCtFfcdnmCvW+yyYnDlXmuhV8txFsRadg3j52pbdkbhekgYvGY7soq9xIEU+S5F
wCowHZ+b8UoTKA0lQD1U8fI7Clg0BIq4a7s2E1lzNerTCsdZDqndK2k23t7yUr8W
+h3UbqOZmXXBcA6VOQBuIYOhLcgPWaF/W9hxpxrdS907OZw13TEK/nKakFmJ17OB
sYjH1TdvaoFfvBd348TjXIIftWZwq/EE+YuDV5pfPbvPKqRjP3LPvJX2BaLtyV/9
3HmWsoDQauQO3RpUqorXyyscpJWt58BnEDZAopSLPPRYEHpghK5QfJa3Y/s0smOd
AGZ4hS2oVaVHOnAm/JMyS12ZxfasMhRwWWDZKlKeuSpfEC2DfKqeZi8uJbkjBJM7
g/MTjtUHzRH1RiO6i5IzVLf3JICWw/+yrGMjFMVaYbh7VziMYnX2wp13VTkAkc+e
iPmD16sr7gY5bciT4JYb13tWPXCdOsogEMkVQK0iYmwRtpGqGz9xjv2YQQc2hcDC
MCpMFypyZ4NjFe8VYI35R2KMjBA3x/vfoXyJKFrrMnNRQlrS4qka/6O9imm33nYP
3pUBtm2SzHMo4f8xVNN+Dsd7RnJloWdUEAiDCSwnpCqs/FRsY154L2Ug5mUSoo4x
eNKuVwKFoECjMBccdBU8jwOHcS8zXfhrAmKxJj7pZq/266t+Un/p8TMsoce1MRgS
7OuH3GypXl02m9frjC1GWI7fVHAfGQlKRj53MI2qralDWdplWusFTxkHQgxiUp8s
lGw5AxuzBBfP5UXtJdYUiNeSV1/CnRVPrG7DB+/AQ4fqCBgmb4Nv1X2YteH0D+xn
IAi0LNlxbTYSskhUXp9pbGOELXLtEJ6K+vrLO08Y7LJZmuhdubP2zyrFw1F/zrq8
dPysXt18eO6Z4H8jU4Szma63zGzwrnb9MlkWocAam7Pi4FHT7Z50naugXEziIIXe
HSTTvwAStEy93BV2WYA2BpoB/dg2wq7IztlS6yoOu9ATEsnBPnSIwaehKbKBWfYo
IZdVN8+agmjc4FsfS52tWZ7rGXo7X9TWH2A1Ho1wyjPTOZUAblpIjCRY0sCA+qqJ
glFcJf/gj7gumEtZxQ0BacUEmATHLer2nqaBf0wr6KhZZp17KZtdVTOcwFvNr13D
TVMvj2rFsZ3Ez36dzhjMIluMkvhLmfRcBoPOw9c6zLQbvdfeHtAxcnSyKeS29Jwb
re441wxvH8t0G0XEktKKEG45JaYx0iGuIo8PZaii9nsvQPn031p/ij7zgRMn3m2J
/rpZ66lOVvC65E0ZlXH4qCWPOdPXHTdNoNyESQya4SbVvIkFNA4vq+45RdLHxI1o
5gw55FuGq+DckUrqmCFJnmYURM/4EEiiLjpwhMxHViWutiPN+3aDSmu+efZB3Jvn
l4PkN3XqdugrqaK/YUanrJl9InBWvkXd1QLOj5c9imfhF0nepRDZPeXEdzgHbqMY
EqDWdtloEOvOFLgWH+PKcVCIns+np75LydO+2n3/j1tqEThxlVhjbqFZcX79EPSU
/4TNiHLeC8IP3s0KARflz1YRgGnNSF46jgdH8SJA/i3pwUpfXRLp4d2dJEN1GBkP
4bb+TMkuIwXBBjt0zZOXpLDyyYkpUUFTA/1yBbDY51ECpz0UoQ1TZmZ/wCT0md6Y
N2laxHRiAEKQ3ehKe4hm6n2YjymzvaF4Myiq5PTxsjGe68dFINmWNDzgGIHn1bzv
g4S3EYRM930oADrtVXKr5qcaABZvE8XtrKJj2Z+wglHuNR6OjFItkPMFZ89w274q
RO+CNv9ZT8H2+psJog5yFdS4oFzaX03BP4e6UC+2oEgOezJnWMB/5AxOQFX36NuM
g6Th9SCVaQdRPRL9mfzjbkcReoAVfgTuwtdkeAgcpDN2NPeGoZFT6cJK5a9E7q5q
QHPy1ec+YKqok9O74TklT1nXeoJG7+uGnSHdJr5zG1zLdIGv4Jkc8Accz61NMgjs
S6Sxcf2GBL8zI+DsVj93tSUu6TW3y7WDdu0o8BtEp9o9C8vcuwAce0TeRFnRpz4/
C1J5FxbSrVYX36GD28VD+4CT1YrBvsLrQ3CqIsi+k3kS5ObDUoj3kn78+VSTpPdv
q7sXAcsF6yR48jOC/JX8cUd2P1kdIVJ/G5QsqM9mIFERwefmYk+6jLjOv5TXbnap
n6AqnOdmCxptprqIDiL5HUBDkieHWN2Zm8nVmmUdLug05S65PbeozOrDW8WMX1do
hhAgz1HQ7Kqm0Ha3QQSB774Vtgs5W6kBqNiJ3L1ecAWf3c7tBpBrC5o4ktbp02Bt
RJmgXsQjk47ejU74zSPb52ZeiVh//Qz2hcEccxWGLJ7Mdt0NmsAS/KXAAzMvXZrr
Xpz/OyKvAIURej2OUlT3TCXUkHohFOmNXZfloM6kGG4EQT5tvyToW1H+R8n2mKut
GWBeIOgP5m4eLljDfaaaSEj0HW1Wi8co9EshEarc6pYB1U9Cmi5vM364TYf1XoVK
GShevTx5t8ZqagmYIoJjRKs3JYUG24vDaAiY5C03uOEg/CFdQ6ra1mVpbGF+oRcM
+tablVQTDmgfigdRoV/eKmLRGjRmZbvJ/Ac9hs4mezUmxkZiDWQsfP+4N+J/Q9b2
tyQCVim4xYwJmaTF6Jte6RHZGYFpoIsWrYoVtMpQNmOMn6BJDKzVMdiAhLJhU9lQ
DSKYwBTNjGrAOvFuXK45aeTLfKU68tTmvWpnhZO2FkJCFUQOOQhj7B9illO+RrSw
obJj0xI5hFHFJuNUG0/l0i8KZ7MbY3gQFoxXNuG4DMnHypDOk1P+DE4bpWt/xv4q
/J4fpyWWcUgdlO5vMqx9RR7hYnhr15CRNtJt6doDxNC/sbsRGyPf788GbZPoWLo8
41cgg7nC42kS9Dl8GXjBTbV4tf+3eJp+c8+fDCMhGpTE4mkAeoe7VVh7YmGPvJvI
7iPzOwHOoy/zeltYjSK18fXf+yp4Sp0/s8H+xarpHXuPgUs0ZrYcFl8Mb3Tagp6A
Jt+JkyyaGE7EP4rzKWjapHuAlUna0SpekUpwEPV4Eg6W56ObZ3E3aJEFsYfvTCNE
OOCiIpMXIua82KI8+GEh89tbvApn9sblvkHRTPUqo+ELn7ehkAXX0mH4Iv7+mdJQ
gO+K6BNx/Ckot3hQWBHjiYEDVmCt1bAIWUOH5DNUdXdNV59oVZKVPPhnkncDyXnB
bCykvuGECzvzXPLgs3kAaLiyowYJXMdJnrGCbL4nUxI0FwOZACmwAUCdRnK+13iv
nw6iM06Y8tsDnzxa2rPYtNR8dxiNHF+QyDkKFTeIElJaovHaOCpYYJXtDyg3hY6D
8+6GJIsteyB43M8dGt2dwEWGm++Oi1msPHcGhd6wqlrAcfpl1pCkAXSLxzrg7fQ5
TvWM77fqgFWJt9U66a2UG1tu72n0l5Tnsn+PN4PcMDKI67F9GC/rvr/BGIwTDnd3
vN7LoNfFKvR1+R2DZlYaYKE6R+2/YTSvdGa4O77PN3XQxztYtzgxxD3krVjyMfjQ
0TjgPWWCpzoA6uNyoce5rlN8jb/sMGl7kdmxpnDOUTyKz+ojBFC3njqoNfqLgNGm
4iFSYQjxqP3wlJ6nLo0yz+xmlUpAKjMc0TqR4J28ajh1tpGwFgsFau9XxWjLtvsw
4PKMHCBk7BcqE2pMuDlRVItH41g8c3Ye9DYR0CC6qH/SvZYw55oVAeXUf32KWpGr
9+rNuu4/j6lH2ejCb7QHLDE9QGO4YZ5Djk+/M/L+SYJ3aj5XXsWUnYkShH2tNiaH
OjMw7eTqRInReRykJpdu9+YYh0Lb07BtRJLRDzge74ol2LUlKTVHtXRq8kTxzdiE
+/JY4it4bkEzFaJXN8pXMSppPZ0SSeTAFUKD/2+asv/mMErhTwz/bQcjX4qdNxzE
WXPhdq8ytIcS71xi043vth9ckuPXE2My3LPc+8QFRjHNvtm1WFjPWyDGDM9CBKbA
SBOnVd6sXHoaS5ChjQGRFZ8G8OJgUdbaf4VQG9C3xWacOd8ZB8yV9O5UD+0eNt50
R2Zfwu8j1QB3cgF1KyUV+OlJdJMzNpKplk5tnGLh9aVGhec1mF41kqdvLO8a4xGS
CX0mKmueV2rKX8g5CeA9ovDyAVTW0K8CjzmxAdqwcxGqNGDzKzQDOZxg8YSjBp2D
5loVRvaO8+AVzwuzosz001dmzcCOVAzFvWFpjytpUPRfRZQ10u92PGYynqYQVuew
LhzLVTZqFb6oFP7/6N4cji00PKrbnv0enLHAHJX2j6GuUNWpdu/nyB536FUoxO+Q
Rv+ei5+hvaygmO9fCwxhJLG1S++L+CP+C0uQLHkgSSEBe9DwNLdFoRuCWk32TokM
Mv4+6o1XczUcTh62ll2wG4avQ5EkIPDnhxr/YlIpNueYJlTBGEa/R5M+hiQwJTFo
1QIH1kUdwQv6ohiqdm8PZE/tXPkOO+f4P/3MiWWdr1zY7GabGS4shfjxWa5xuaO3
9vQuLIz43LWFInvVxxcs37LBVo21ry6qEkZesZIb+nRP4vy5fgpvaDz+27iTBmpR
ZPTkur8eQHlX88A3l0NtcPNwD5urHXLZjPXkIkUYgwavJbZVtkZ3yn6w02Rwi+Pg
D+y+gdFHC0j0Mp09V1ZTfnl9LafrzACbwR9Aet9JcWMK7/qrra7FTk9p2dTWc1W+
KuEXRCKum0eHbm7vLL/kvBnj2hkHCL3jbDmneC/6rMItDiBMgI+4S18xMaKAAn/O
QQ/B9v/r/x3zHyuKraSqMka492e6nxvgBdo+ZMqWv0sfnoyiCnvKwzZd6pYC3Lvx
ufu0AorcgyMtcR9b97iaJ8zD1arz2wVnp2duSkgQuUJb/dCKtZK89LBGlpqLW61J
Uv7d4+wYPvSfvRYD44s66vhJRgOdsdGt2T45ADkMwTdrMhoVFAAimdMGNorOgXQH
StIU1wSBTqPL4M3DGUARfupFtFrGOcd+LRSAgzZR3ENDp0xc3IkkHWk9szQtMBUK
tNSqXa6wvS/Z+RsohkVt+ahSZb+zQsAwrctUWYKfsNhz61hx1+1ktwHzSdbPUNp9
bsXt6M2nt7Y24bTvQMDJfpC8L28o0YNSvRqyfDEwYzk/Ytye8RttbY4Nvu5WgZKP
nvd9g7ZyAc/yDeYWdte0LWV6d/SI8wgN4SUCdIPX4Padm7r81Y0DlftR2zfnXqib
Bcxf1gNQ7VxnFDOqbNgt33krit/IwY1r5AmhXi+Q4vXEm2/iN47H/W1R8rn20kxj
/3JdkvWJovMUxsZQEkGsJnyIkd6X15J5cs8dfVP/SPtBWASYS+FnKa/yuReJWuHx
nO9uNZf8fpzMIzvHq7wYIY458bSnFMXnqCP+29VBJ4WUUEZmpvXvWpGacpKolUjG
V+txSFQidonHw/yD5AwZiFkWGrprv/HVMx6kjxY+E68JLQl7Yt89mUrCQQhP3sLL
bR6ewZBfqDHZsU0fZRc4jhynCN8sSKdqi+en8waZkL7QFKrDcD4qXcXM/sQUJdEg
c2eC/JKar+mGCb2kyAu1RtiktCMxWXv6AHwiXyAZlkoiBZ7zjhquftVlxlP7fpPm
rUuDXaPpPfWdvsMYx3ruMhdT8B3N7PUA6j2EIluJNA+uxsh9hbcqr2LEKUqP2xb4
wovZoisFPA90n/VhtfuhfuqIWnSTSryCUCAKqoPh4qmKgskQ/Za1cWBOd+SN7enC
DhIvY9tSW5qhEZzkJYphHHuqci4ARt38rCemKEO0k3j3oGg60UkOxSYzVdLAQeiB
qchXeLwn4fweu7oQOrkDmwIa2ERiXflNLuIwQZdwGg5F//u7Eh3Bpk9b748Axqo9
Bj9hdJQsXinHcKBOJfDY+EsfYfAGd1dIWeDbpp7GogcQ3KHHCyFxuagMiueME5Su
M9dbYoQX0OGS2VAQBCgyNl4+yhJdnoECoArrRtehOtdj0HwzBq5O5KY2a19UdFt4
RS6zVdAQsIpJ4xnNCKGYSWF974Gc/hEyvX/X45Wik79bfHMSpUASLmEiUM3Xda5/
vmq3q3n806ALOmGlrlvYBXtciOnYSH2WUnKoezdWNgTDTOOTEpFQmZU140SapycI
KxICY4Pn4YGpwpTZatj/sP6yO5iBh6EMbZkcomtTQOrjKcPYm5zDuatCZXxftfg9
aH+2gXGSkoD9iG+GySTo9numGD/Y+xBiuj8qBTRFTw0Y1lv02hE1GCzEE5o8vKht
yqW8c2vy/3BmG4loLOgE7fbVth3rxfml7VdWLDEK+43/0u9VkhBSiYhMjkbr8r+n
HqLV3WGVsni0Q7OwV3fAqdnkqwZOJpr3Gwpr9U1DqUlXtBszjagEfB4m7S004C0U
cKi8a3ASSKEhQ6Xn1p5MvcOlbY7wN53iLCo5zJH16pjyQacojJJYkkvdamSWLsYs
wWNcGYhLJnNkjqnvkLsiHC1Y3nVOkBY+4HDEEckAmIuYztCJeKoUUA0/F9LhgiVn
88jGH6sTd17MbZdPrxq9ZuM73+SrlxxptVso9W/pugWBQGFA+RervwRROiqrYIkA
KJQgNF4QQ5M87VuVahSpkms0Rkj3BhKg7cXKkOx4S3zl9Ew4EtcBfaGhpFreviW9
qVGMujblSkyf1jC4Tuxaa2aw+CV/3Scx3VMC7Fc9EDEqWoYYpuUytkn5uVQ+q7Rb
RNMjD4Oo3w3UtrQ3EalsQfIax3C/GqsF3w0PNMBdC49L/ijKrAW/lPpkHKmkMAnM
eNhq8wHqSrxOPY+uKuEQ1+RRi3fbxywCByb1NqzKtBLzEqovuXFDLT28S9NnFxhP
jEWppWVctm3qIF6Vzopjqlwh/S2GtHc1UQIc1TfDFsdvoPrPNEamOOoFgugMAhtc
ZJi6Qu/aJfPdQGU+3wbsi8yE2c+E9/7B7f3tcTsUnn6HzzfHI4/EMnuzW+U9oZmW
mwSfPBYXRUCFBaUK8N1A35ttsXPOW8wtFsUVE4jF5pOxFYacE/YpldcuMB5g3vIQ
b8WGQxkjqlk4pW50nV/XTjs8ekJsehAFaTegYmCjn2ohI2xqxLj/ncLwmAGOkRpG
DrCM+5rz3uDPn3MmI4JLjmsigTNLlWdzX2dm0kzQhZb3WI4itbpJgUNhRayIiBS7
jEbEKTCUCbHZyZF2jo9yNi+l4Sb9MwJmNmxDHmsMvlO8kG9fzdy0ZokT/kxPfGWc
k06ArVs3DHbd1NDKKT4AGkUi7y6qAnZ2mK6wXe9ueU/eMcEVGzJpnVH38OPwYj3b
uJH6AmP4ixNh7wUJysQczwDql4oGCQJNNAx8/lkk0fGqT5loTMV5WTZ+v7J06VRg
xXHJw0rJk4XNL+DshYAR160k1qHii56QpPX1lOpEx5vq3LG6LrNg7R1hgR5yAcsZ
2NvZ2P5x9j/RSgVhnU7ZRo+htWnAMoNmXHV/WnYBwoUJcPJofdFBjy0mCjW5GEH9
DuX6AI5G4PAzoKXvxoiG80Yi5jFTg+orBWKn/uX2wBC/ksNu7sBIxnxwb3xo2O9h
LrlOc5Qe5piDSDKQqn0d/NlfU24uPkIPu4tHeeqYH8lv3sPCX0tgTR2W3UCdfmOY
MVfLhbTJZ0b73Y5r97p21BIfaYR3i4NQVhHaKHD6+qRP1UbFE0gMyzMpNEdUnFmt
a6QmGb18kV/zt9soqU0eVEKv09teHZGk4ADO3kUosLCNcV7jfJ8QqsW/SifjYG6V
FmxtbLIkRiplji/iwb2JL9FChUQWP448368hXO7sanGpQHLgccsNm+yiQpq1Wz2n
ORMSxN4Mp67pLEu51rJedQr7qf2uBSab+mRH90yY5YbeSyXmp9VvQAI1TgOsr4RF
fnwWPsyWDPX4ZB/bz/DcUs6NPtPrAI5uBY/C9G5P4maVenEPDnaFmdtPzxqrCJAS
9ZcFDqXQ+Ck9SntLB4wPf2i/CMyytG5X0gzFkKrA0FswzoE47Ifghpp4nd7/GXEY
aPsdp9r474aFV0wPKVknQyQiVQ7VZ0Ks78oxejhwuwiDkxUPRk2rtW1DTbCfHL0M
il2H/IVlPiRCcr9lCJlwPCp1Bs75GvLFxLIi9Uf+94ilkvS5eO/aLPNvpje+KWlT
xcjs05hHXYIKbT8UDiI5a0+Nai4ABdqoZrKxAoVBT87kUi90qh2bOyxGaKTxkKgT
mIJe9upBVH+6kl57LfpQTeFCtnQrAYOTYg9cftkLWeISkBSCuO4Cjim3GoMxCiz3
PrXbq8hJfi4OIptP1aIRvhMpQN7dT+gUCztXMAxOlt2ALXVm5qO7Q2ZUFbDHGVs4
XjvDPXU3CElzhTxj1L+3c+stNXcwGQ/rB9p+WiMudFsL9YeL6DEKN3AqDjEXH+xd
Pp3bsYGFXre3vXgknZFFxp4VU2hqMIM73PCxf+HmCgVUZSdVcj4mAW6FnJ71Qsbs
Qs4E6vTvQtZ7FOcYics27pACo8zks+5ePGMa8ZUz5kBkyalDN/F1mAEoXRBu2a0Z
eBI7/VLptLNBTGjoYO3bcpizooUlNSx0LXLq+aSzLjdxu6uCVk9UBycijEWN+onS
LLwlm4saaMbsyEJeNZqkSTy44W1+e3SdkAZ4VZRAXEb7OjH2gdcVu67n03xDgnHz
6a4Q9sjI2klsCInjBt7di33zwMy7Qe5s7IkK4pmz9arV2Uj1GohhYUi1g4eZut5D
aYXgUwDdFkViB/cigXmv9pKGNbU4P2ognns7/dMBX/s8bZS9u778nQ6kSrtiCt6n
+/W8nNSiwqtuo9b1phO5PCv2TleeykWaYs86MIgk3e32bompo3n5AGeFXbIKEMhw
xIRY/7Kn7LFnXCcNXWh9YjmraoTbY8ZS7AjUks9esZ72wZiYO5aZQeK2fozHDgfO
HFWm2yRYvpQP976/9WQGFF9tvJ2FZviVK67tA086GbemaIplGfdg2s+YloPaqAq8
zHkDjFTeZnL1NBHTV29N7s8HmGulTQ2+Y0rHuZqZ2m/n9tzOHA0Xb5dokqa5IjiV
xnDwioH8gFssXltH2GPOGClrzPY6ioC+rTpVaz+K+KScNCVk2DAXWUqVjqdGsMJJ
f5KBUpSXk6hdUC1AP24qOXKvht+0Sa5a7pSZHUsmSSMOFnt26kfCB5GGNybrHDqo
ikvRvvxjyixPUq1eG25GdA3fOW9lTDCufD93fKCpR/Ydcle5X59sB0KtWcwEw5tS
EWKVLZkhgFmurxhcpcMtpJnTrUXwAcSGkGMxT8WltwQGFT+cm3D/qt+EiCG/32Tv
iY2RJAyiShe0Wsz6rC1B6jr5sLZKCnG33Fkfy3PXutaNwTEmiui7Lj+EuWD+5/oG
gYFnbv4HM/M2ngY7IMYgGnnWWi1QjWR7r0HAEFcSI6WbKXcmGad2psYz3xBrVetb
Lf5jc4T03aHO6BzSQl8NT4gXu4K1xUFOZffLmDcbGH6I0yPDyLwd25RU76LzKfZS
cPP67/QIwbBhLbsgydjTH1kIhcGkOlHyQSzVY8soxFjLhOEtrbOVFVAdqdTNsLPO
OtrQ81eZIMNdkHZJxBV86J65jqzR0Dreekn6DnAIPwNN1KVNeegGsgHh3DrgDp6K
+OwfWk6T9Ao805u3EqhXX9zadhdgz+IOSqzd22cS5taXzkFVYUFzD3Xc+KYHKgt3
f/REdEDTag22sNCZnHIx3U+eSRoNpwqktDn8CcVfbOc6LrMIb2WY9bR7AtvwqdO1
jkk2uphS8/cdwmo+5CSgC8J8G94JjdQ0vcnpC1HFeQaAutFB18dPnT3tKefuhefr
e9r/NBA7dJFY/0ugcXhZ94nCLi+nvYl3buLb8lurRcP9QVtuCeq2iVkKEbowAwdF
gS/ARn6CUihhY52gZnbTTArwf85HNoqP45x03/AQUsb3beJYR4qd3vtn5BB4U/Gp
WrizxqH+QbVEzpA7XmAC62l8pxOW403if/GQUenI9G0g1QA19FGgcOs92rTrB1PC
hFBoIO/z2JDddelXTDAZ1KtAgHLRbALhpPrLAiok3tgfRzphdBbHti3Q5bzibdnp
b1DDXwDJtdZkF4BwUkZtCW9FD0eevMRszg7tWyx9RG44+tgq1iMustNQhTWEFcX6
u0gWHboECROAT9eZ1kF4R0LzU47RQthdexY5RwRwIa+gWHjXRK4x8YXe+BtXs4wt
LFXdq+hYcjLpbC5rE5Y9pPRTaKr/aliEFVDgyUuSBhokEnQhXr4JY8ozvi7Mr663
lTxkUlenI/WD1DGHABEnrgwmhJQoYRF0w7DH1KWc7HSSQXy4yBODfHZMTcqHYr2c
2yRi+0Z8uKhxSOp57cRi0/TgJkSsR4Ig/eJ9D5fyPWKQnLf12sMEHIYlaTT3EfEx
guEGQ27d8I3FT1S/7h63nABeN1EAxhuLE3D8x2EVwrKKCapEVTJGelIOlbL7ufgm
PoIndPtT69OYIR6NbHJN3i868MJ1Ohk0PJNk2uaPJJd2dI4z3ejZFvE6wqi1d6rR
XNkYrefxWaEEF14utaPTKTuvVht+x1ErDND1F3dKsxqCZZtp7O4188qAmDwbzr0y
v8M8/HbKiOqhWeWz1jUHNyqMhI/aes7vxHc/gIfKdLM0n5LetgbkCD4OB8TemxyZ
q41qlIqulA0KNqKR4AskZJL7kFfOsHu2LTiX6Lct8GzDqYLJsB5H1qZ/Km9RFsX7
4I962rQ9qbhBeUbnYU6ngno2vwY9zNWDLVu6sS2vXNbZNnEk0pL0AgAI0bjf7uDJ
kxQVZp7tWSE6JL7Qh0WKGFj9qam0JiFcM8Y7vOllffLj/jtc0J9dwrakF94mvpaR
rXomgPvRy7nzcay4ksqLCzqYv+p1NDF+krNVasa0i7IUDkcANQJL1chlFKWj0hIp
AQrwaV91BEnCpwf4xUNCh6wT0uBGvN8QKLNdDK/SUWWR81eakZD/F11oEmsshKXo
ob1t/y+xR9OtLesoAMAI1ZfWv1gGuUjC+03VyklbPXJzxxuyCI+zpYl/IQ4+7Zw9
hfJDAafepxIrWHEr/YFFV310E4nBEdJqBWxIc5iHLqo0/Devx0cEGe179oT55zR2
86QC41PzQlw17l+ZgH/HOAIT/odG14ZpikJVFwghPA0lrsDSx4TohXlS1H+LXvXh
DAcLVHpXWJUPk2VUotnnoQAr3ILfmK8oEiLNLEDB+2TzOqtCJHzEVCIcU7dbHbFa
CzZPgysyij6nyFs0G/TcDGzczvthCt0mb3z50lC3lukhIluK78UmaKSqnXQDhYNF
7MAagLF2VTI+FPN7+SixFOk3Lhrg2qIrNSOji03GPrb6rTomdwRqSHkNcdziSYUM
8nxrQWsCfNyny/xABuH4C5A0T4KzGjNdwbYpiZ0tPfa/I4Q/B4mjSanfa3puihw7
7m97paB5xL2eCY65MmFeCPlR61Bq3hLikCLjU/nN5noKfXZYUZTV3k1ptlfXQsnl
XXOEPz3QLTc1OhquyeFTkNmQWamPgaC2Y/SSrjaYEIFWNZSEgJFpTZhF/2V3qzGt
pHyjXCAtwcZH4IfH/KJGleB3nsGdgcgPJQr5qXf1Gmwj9YA47LN8++kFHZTGQk4T
Af4f+L4ZpLgVXroEPWKURqBxZ+x1c2d/9NWJ9d1Y40hckEXoJlIee+dI4ojSqX0y
NK5ICEElFk8sN/DUP6SmzqvGJ/mj1sSaFaQLE59hsoySPfcU291PaxoVzs5sXRCn
VX5PffDPpNScTVELR3U7P/mRBHK3CfrJ4HckN07F5CByk3Mkt9TD/p/VJeq+7V8G
zJCx3N1Wc13FazYnjqEP6QWqBRIFmzCtlU51l4BlEiTka+u3fMUAjrn+3Mowesbj
GdNYSo/rO9u2hhgjNvhtb3dg+T2qhXNLECD29M5FO8JUwiw4FQpmF11F3uCj9d7P
W08VfSrvEmlFZdFX0MefEq92Ob4sNaXfInHQP10TDoZ2ABRm9aOvNn4yBeGGLfBw
3w4JEeLDm/W6sECs8lNcejPPrX/vmXcToA3F/Ex80IiduMe4bLpnuDVT9en/bVSW
/CDN0c7zQ/O2sulyCt9TNjQiZAqrUb0YY4Mon2eCynDNvRTtemLGWBdLnSv021fR
l/J/Vt0HY79itg/c9FZ/wRNilIIYzMvssekV+DpFeIRxu15cJEDBKZXNJnM5Fdeo
Jclpyx63dpM7ttQ7i17tL4i8sqdjlzIZiDhxIipgeGBUS7/YMVhsZwSqZBywPS2K
RDHQx6ZVVdKSi6L0zhHDTQ/i1JLzcrLfB4o02TdRS58HJua+sDaC1ow6vlcB5vLx
GJ9hZz2k+8b/dKJAcBK+FD1VUks7kCrMUURwTccXl4EmLTeDgI3Lw6SK5IQYxVW0
gEH330kvTM90beQyktUL9OPsA9zXy9plxQSRhLD2WMXpN4Z7keMXd2po77Qhov2k
5RxfkA4GYkRjr95CUhDhW+fN1Sh765Trggx9x9AK1MxTnSoi5Y9/4E+uLYvwx+fF
xjJ+vE2OnyAnnUsllyyzvU41QRozvwgilA8Yvz72giOynwxmbaVC6dZRNwKbCGhk
1zFcshTg3BEK5hz/hdhoTx/VlzqsvIGmVutLDSRNnYB5x5zth2968CRyzOA5XfmB
LtYdLQt3HEmf/TRyju02RGIGNQdCfilldbR57hGhmDIER8/4dfGLFB5Wh3a831a/
H0St2vmWd778QxNoBmI8gsEVy/s1g25deGtqrBUMPmoFCmHxG0ZShGAyyiidjydl
OJcr0SI/60GADPy4QZXhnX8AwoZ8blVt2KQDb/frYpO0z1J/1yzBfAc+pIMlsGpD
2AeARzRpQ8a70UkxhnDNQ9qrMINiDPkIfKU+DkVvBb1xZu7syG6R8rHP8D9bBiDo
SLGlwiMC4FBuMRLmE/P9E1mwetxyiChWQKS/rZQFYsrPLjLn35p2zxIkKqYej0B6
1O6sJhKVVKkS38k+nmm9t5nUVmBWtCnsUVw9CTrMHZgLRkZqEBzelrYepvHvRJss
rbCsbV7tTsDY9+beReH8i3HR7PYxYwAz40+d3ReXqvkDOPSSeucE5iSeDZXwRfkb
S8G+vppcCd/+oCNGtGLI6FvXAZq08/0c/vs0d5/X2f1x642W7ivHy8DSlJh/i5gP
TXoe/vA4//pdcOJT8hrl/9nPXUH+vnMbkmjowyY0wIgnokJFkXUPWAcKxoe7tk23
HFXHehnbR4A9p0jxMXTKS0dkOOmXdZ/vEV4mKZpbjyyXiz7s7ciC73K4IXhUBH+M
H5y8cqqm3FEklTN/ieHvf3oqjpYVbPcM4yqFJbCDsBiUsJSgESpdgetfPr/sGqsu
tUG7Aduf7+kFN/hwHUXIjjGcyM0RdsN2MMaSbG7mXvG+QIpOaHl1JgZum88j8sgL
P7KGHnEJ/aXvKUZfCVbr7LWcf+qxoVPMMvWTalNqbBDieKFEQ+dpAkWrrCU+4XG5
C9kZc1qUF661i8CZ9Yn4WTbcGemZ1AtNUzK3uKPlDs4gaWk8hoz3BLQkpZfj4NWA
6h0ZLit0OHvDu4VyIXcqIVX4BCF0/HdDS32ttESZ8UP4/dF/1rxBaWirSGaOZWUx
Z8jfbhwWha4xvYnZNMLKYHHUbWEMCtKNurCTOvCRkXZoiKEAqU9fUe43Zrt9KdIi
ituCMJ/HJ9/ZtN8GITSqXmGGDyilV+kqqPgz5SdxzMUHTa7GGdkyX6XeTvEfxxcv
oB448JAhi08bktOUe0o4oXZUQ0RkO40HFzw9B0iSRdvk14EQuBM6fz1g9sU8FekI
aruegtQQ0Nz96VryMP8j5OeyrFGLQC8XeTAiPZW4E93dfIt95G85VaIy8nUKnBuO
yOGB26qBWmjMMkQwWe/zai0zv1SqQ40bXPXIfV591s2XI4bZIN82T16zk1Q1bcO3
XQvTU/qILM/dIxuNEeruuAzavzrCGQjyYN1XIjXwrzymk9GKDkofzHHHimbJrUCC
um9zTe3RkBqX2HBTFIf5K2gRmH49AGFZjY74M+xRA/SqlswB2L7n0e4Sm20m5QA/
HIVDFAbF1aT3fl9nOfPbwa5GiRbah6rbrnXkXzoGB/OKMSLY9PfGQWYa9xbg63ll
cmHLK49kgVii9OsfbcLwzDt/wOvr8WiOBsGtY6v7YjNAF4FXre+/con7kQXoRVH6
Ziw7l9C5iu/zYMo+2cbP743thQGXjXGU1u2KxUdty9gldObWza/sO+zFEfy6WydB
KCrtqngRNSCJiFKojF1MO6Ts16vP9Uk8SKQWEBlRO5Xq4RNwjCB5afbN6/EOys/9
lrfe45JfJAanu2fbaxCdckMS8703xNqmxy+lGtuUVjNoWXyAenkfeHP7WA9kJ7gZ
5AHRVGSPzSzY/maL6uN05xCjfFdjX42/nqZD0J1cIX8dHnQ9vOratyDhqeF1eqxJ
cPO/haMXLkhjJtrAc6+BSnGQFzCFM6Izo4aixU07n3excssOHHSfke64yyJ8ab76
vQI+lrXJyooiZ0D66gARHY3FugjWccmKrVDfw+1QQVbgYMS/HfDhv7PrViAm3Nyg
C3UT4sZ4za6Ds5ozlFirO1lbeAMcVwKC+qzQCQsWFLLhg9ngcaYWpBlsXbUmfrMV
Yw4N6Y2AbxzrKkhcXkwwe32ifBD6zOO0Yih9LNYLLcYOrK7Rivf21ZzQMrE3kuUF
8ghfjnZg4/J51PS6PH4TZFQcCMIR2F1CB3/gCoIAWWWTSYVwlDHjsgA1UmIYUbGK
Az+oG+PqkZHg3soCy6wVHpwr9TAJ+EsiKntxSlSG0el+dR8vd/RYA/fqJ4blrCEk
ys7XDfnxYxzYru6sfKNnGmL7uQJ8Eqs1j+ajlbZ7RSs/DfkwsDz9GJzHrqwONsAF
dxkwTwxM7szSkHAXJT/dwGc28wsuaQOJ1b+66JtPZhv+TcsTFICXSIqHwKWOBco+
5P+P+OM3S+mrLcRmz17ZsWIqOcApVD9JZ06ulJYtOr048jgntRgVMGdK0ITz+cye
IAJMF5b6aD6t3SZI/xX+A/FawThvJRO/m8LrJnNvJQJFO1PVD7rsSmGRFdcUzZAf
vOadjHmJlOQ2g601n+KKyhIO25bkeb1aq3TY17IqiTRgDD/niI0C+2CyhdFVwO9e
N+/rj4q26E2UizuqJth9vBAPA7EwyI3YGaJGLGUJjWqS0duOXMj2+tnsr2oTItkZ
ERGTGnQwQytu68NeH+3VIk/bisZoEDvM7XS4muIXqI4qwA9lLX/dAzKs+CVEri2m
8w6cw/6wvk0LKFxNnqgkB+R0pbhxFzCWOhAL7qyA72qq45oMzvHqC7IHx4wJA/sS
oi4hdwjLMHZvFOHa/6O1eSsP7KTu7nGWFDdhCidOmej5VYpMQhnwRF/cyeqQmI8m
xNJD4oRTY25lgP6xjzfztuA07nPlWHKHle3KHHZolkDoQ28kqDqyFRjzoI/6bjZ6
wKIzmmEA+jyXXtCogZoWXUgv4cJbhFbp6cSQpq27gwFyKQRy7C5CrAW+YqVX4Axk
HzyrkQUS7Fw4MzLYPTlNYlp51Xg5nDsd9YwHU1Fo+6BgU6HxUTForHzr2/ECK2w/
cRQyQpc/NsNhUJlG3JRB+f+5N+iGHywTSg+gqtNu7GtWhii1ozL7XoRYc/TzZJZD
e1H8IBxvlNrXrizEKRNj68YlSipXVXI4tgDxR75lwrWT/cknL5MVp6FpsLoaau2W
/iOC2ELV6ypGQm5oBxO5t1VFzEGiG+z3uNdX9tTC6HVul/S9E4C922MHvtk+d2er
qdFOgm80sAalIjgcOHra63anjps3hpKhz3NHenOOlM6iADz2MEhaCShVwRwnCX0k
+FLPHA3x70OeGZkM156/5YKXoSpKnxnPDSMSBO9oio07qERYNiYuP88PtWdJG+0i
+BZf2rtIWU6Byuq2UyO93e4KcXl4U8aEqZQV4w/8TYeRPHgYQM5PAGUEbxUDv5fK
vn/3tHwET8qLTItz69JCoyqfGv8507rPMvV3/lYwNk4yYfUAZmhEuL008TK5FYyO
jyqICuDxl6GuRooKyF2WRdUdtqiuCfKc0BF+wSCTE3Xz8i1+ng+bcZLsoogbJxiJ
/Mnkj0u2GDbB36SD5RMmyaF4OILQPqxIHeEq4paoibYurlvAiGyGB5h2hebXKNtX
1V1W657BHcdQWqj9Eyb2kFw6E9zMyFf6hHq9neMUfIsTuy14ZV5fbYaJ2LClyuOj
PfdRbx1QhFgXA0GXXmew0NZf2lVfUg/O3Ro5aTCLlczkYIH1OYt2xFnqgyxuDAhb
9tBjOcncNC4CBD7LlYd3GGFxEpsZ8fHFP8iGxLS3ccnaAMiofI/JZyGmz9Hm4Cfk
DgM3zMaQvgsjKWdHeCtYjWr2up8fvBHPEli0E+u79uUuouo7EqSpBA/mOBOryEoe
VcNnRgvvg/4PqH55WMCItBjk44P9NgSaaGCDFVSyEDUQA+3ZhrlDINN23NvKh2NI
cvvskm5mJQcMN4nHivQxCd550rdBFyBEd+s5qCkH/DMN4N21JI13kbJ4TBmSeW/8
SH5TX/lyRsMib7L4jPGm1So7ADrFDBO3F0BO3UpF7aYgbx62c58K7cVQ9o3/OOVh
L+mDz9Qb2QxX8pAjBMDDu+RTuSXeaxNYhMMBBEiHlDfbzgWiAoPfSL+ugkAttGAT
sziLPOBS6t4EuyJyV097UvqjcTxm97l7ERr83eMXqvroSE59EWApaJ5q9/MqtwH6
Y5JB+MMWiKgaKxHNyFT1zPfiokibr78gmuv8VkjYq98oP2p8cyuilxVVkJ/vy8Tu
CeZzeyKDPncGQ/qEotvSrAOyuCL82X7DrCEa/6Udxq0v+WEC15gPhZpyO5hBI1rr
bhjTIKZ5CHer2xQriKOfO5ptTO6jFjgcEYTYKrgZghhQcdRQ5S/wMUTD5U2+mJEA
VbUTKbH0A6wiXUox90R8V3FCbAbQGN5vl5PJ0Jx7xzW+J1b3gffYx3XvcfDTiNX7
9DsWpOx3tyJAQmBELprYJGMOu+c+WdnTrnwrTY4oEhrxNpLoglwau++kJKRFrB8z
X3tKHwVcJ8mpaEzEYLbRdgwwwiFIqyZcAlpCy4m0oiG/WKvOZED3CDrcdBsQdLfa
rqBQAkZjuJ3opHESBASgddtFDis4So8Hhkys4ZUvmn8lCaaz94s+f15578akUu5D
C/r2RbvVDyOSL55MulYE49iiMhezy+LFqlzr33KkdmW4u0itLh5CCuqzyYyAcdja
QFd4Dej4rGKuJO9SsDEkeTGODTqsDT7/fcB62eJffpTEYEw+Tt/5pg6DeF3/tb5M
nekAb5ZLf0bCq1g2DEmmkKFRbk5FZ5NpoLGg0X/8THvbtO/W2RXDriMB8yjSDsku
MrY3VVmgjcv1DYPZeSqC7lf1UJMHdHG79kG20yvQJDa3PxEvt5WO0H6UGL+xVCH5
5CW2AtD3QmDQHCtrrszGn1AEH0tC7qi7bx4pLCxUvwZLXTJrU/tPzCEekMbMomBD
X7jHdS0srUMRbfPiXdesj/B5KFqBCGBiHmoB0qsNaOwO39KQX6245u5B3Vgb0/B8
QWHvc0JDAHQO6b0Gp+y3FoqRvISpI0QIHzmvK8aC8Azlq0PuUDGA6H8whr2jaTon
ji3VTqFX0WlVAmX8RYJ17WhAzyW+wdro6LkO6Rh+Ekah7GZVzn2a3tPbxYLP4xMi
u00e5iBu+ktp22z6ZGnGgHnJVCiMstSKPFjCXJ+ndhXuWeoiNVA5mpIshOpwRcv9
u2lb6MDdRnwiMYSGo9ugZ05M4R214niTs4BE2lIm8lbQDljgBeOqRZcIsmLkm5Ni
0kqG7YOXzt2C7CdA2rdR9xrY3PydgAwdKJnaeH/yTi5P1zLXyEZt5l2mhtt5RFq2
pCynBkcQ2G9FvgCKyehqfW5pm7wJq0oSZvjvBeknJtstyD4HMuWRW1seYYQ8BTG1
RX3hvNFaqM6txfbiLPnCekv8h20AKRzgZT2RHKafDp9JGe/VCZT0aOoOxsS141Hq
mbUMlHU6NCsH5kzncDiOkoJLeWlmP02hJVt2DFxATHbeKelg4kSp54OF0ilCqKq/
EZ4hFLU2PcDZvweoWm7ts4b5Hwlaz9SQq9CY00dv/eVMMVEvJnjjMbQdzhb1X87M
/7PQhx4Q5sv0DcYKtjisN0viw4A1rYBd6sXKqicaw7WtlqE3GrpmteSN9KB6VTjl
TaNBfgsjuyWRf0F0UqQXhmLabl8S06G2XX+DfVR032+6SaoKjawNnizwQV06aVqa
M+2wK/xxRp75CCqzE9XakGn8I155DzyyQjjYkP705cOAmy5r4o+aeWCYZRzURlVd
c3hTCH9V1KaN/4qJOI0imtmB1zo0PKlU3CZr0/RK/+Z+LK3/lzoAEnbZfISvmvok
cLyo6XYGfuHnbSZoVuXsWYZSdpSzvrO4YgmDeQa8Jaha6vcBATf7fEx+fFmDPxCK
ywe0RKDBgIceRwExqJ4NdW3SVEicujtLf34puKmy6qvodPmXY3qWp8NsqlyAksvD
1BMa6mwZEs4vBc2D4wk0AbdReHrjou3qlScSnmgRm0WH72mdKRABOm10an0VgU4c
tOjXbNOZDTuhh2rCQt2CpDHa7ry40GqNGuFfHMiDZlzxgrWjQKfjAqFrnSB+9Vd4
aBoaJ/4U8y6cAXXneUNu+Z3Wfn7BKyODlqPlQV2iZqJT6sNDIfxjMQgZ6899XVFm
Ya7J7eZJBOWWlUhaznUPrkYZ0/EVgCVEggpbYnnH3BccfSLc+6gapjyHsjFW3ySX
4f68bcVppNSwLn2CNh11A7yqpHThTOSfQbWoggScPuD4yUEEBr/xl8zRB9aK/NH2
bBMEmVM9lwvtV9h8ZchvODtBTMnKLcMr0YpFSNkUiWZj6bk5ce7GxnCps43TRAbz
Hd40SeG9EGXwjSwJCrNx7JazaGRVPQ93DcBexyNDNTefM2v16T8xW9k9ETbInFq3
NjHAxeoln4q1f8BFET3Z9PzqUjJRZLK4sEBtrDXeyuBirF3un6nws7LCN70U0M4D
S+jrXcXZedOC+kDhMUTNm1lvCHPb+15rJpguoR7k2rqZM/ZYFnK6D/vhzAkjHNkZ
9pALDXtZpNAULwgzoAuLqC6quM1Z2Ff4FKzuCwkRW4dFTyF/3kZzK3iCzZBZkuoz
gyb9x+XzkRK8+pH5sbCVUt8GDbadiTgMPrsoX6wFMUNG8qc8E8iENbtudJ8R9Z3M
a6MqTE4lHztisfXeKQqZ1RE/RfR6oiqxLkAnxMdfiwcQTqvasULHJ8eW1SgWaesl
p5D9Byw7YnX1aR75GmZTkyKx2+RCoG+rirZEvpVoQRNjXZYunW6X7HlnNhKuLGhR
eu4AjzqLRFUw9DLnTnrOfaPXG4Ep+xs2qdy6T4r3v+rhgqRwxG567d3qx1Z2RGnP
NKRi100rksOtreMSZ/yXBrKhWV+wMo65KuVXNkrE9jafGNqc/JK6ROozSAMYXOhS
RrjbE90qF17jyFJJZywFY4/4wdHOeEIJ0LfYcK+TYFwhYbO/hZcLKzDweKCW7lBz
dJ65v7X990LshpSS1zWg9C81gtoKgzdZgbjMfUC9kK7lKG+e8IlrTWfb7F+lWFOg
7++XbNU7v3gLMFAKILGeVqkJLDuS4IuclgmWA+jfw4AN/EeL4b+eIeRdXDnHIuy4
TSSuhI8PeCS396u+1anubJKAi651faF8AcEkvpkgbuF7PlR9J1E+b2wxqJWpZWoQ
mpBfWrewKVYpcm8ePSqKYMFpd3MCzs/uC9utvE/3Zn05TfJUTTjZVqhsvmOE/PM/
9mXPZk3rEfJEsVUCOWdNZW8/DM4SDV7LEZ+n8X/lTKXMpigN0jzhSm0Nm7PGaEmB
+YNHkqipHhC4O7iaT5sN0lP2givc1VEirDus6BgzUnP3jfiCFBQAkhffdPjNaWId
3OZ6W0PBSwyt7DwgmJnpxe0vK4BITzof0mI/yrH0evCLnIqXENYSNuIQ4Ctt66QH
pS6gLxIHHPgieisRb33ayQ5Fd9xihsL1IG9O5Fr15wxMylP0r7d+ZGIExp7/6Oe0
wcpz1u7sl7Ji8cHH5tA9PmtJxBxIz7O41YY/C7huY/A0cMEHebUCsuYzuAghRU50
QCgQ8ghHTCQbHPbrVC07/y5hFlNMPEwPZepaVDcpM0VZRp1HmYGJXnYd6aQyiRh/
dbBmKMnmy04FDzS6FeeqsNhMOTLWm2vF5rYOTFZmw/0og9YjBwt9rlvrhhY8qz2B
+F4A48ugQqnFAISRnTB8vk6XoyJrpffIk5+fP4IO5nEjDNzIkXZ0ifq28gnkDSu8
+Wx8zxNHj4iLfu/Hwj55xLm2it+9i6kiLxCt/0zo0Y/yW+UM1vs1C78L7FUNO5ZO
Kesp/SJ4RSaxvYfYBsQye8mraxWPhfdPaFO8zZOY+JUTfOOfQ3O5VX9XtiOewDN1
qypYPqSGmPmStHumxSplNOt7ASZLlsR3IsQBbsvoHqHfQrNe8e64H9IOlL03+2i1
LD9l4yT/NbihbIn1d+fIxymRmgfgQEp6bkySR0MQlCT59R57D9h9JrvRomhCJYQE
NyMGaJU2cqJvDBqRrp8AkHLZlsHdatX8gxD8f8WmSZjHPH/7wxartB3EkT3jc9fj
7TQR7B6q8J1xYbPnbsn6eVg4O8oCXb2pg+0ngWMF/nm1IqP2mFejbJL3DMaSgUWi
nyvrql8Uk+nW4+SwUzxMaEYX1RAWjuIQYRZ9XC262ZooJK1+5cTDJfEi3t3KSzoS
VrUF1E18cIkeHj05Ev58qKe4USCaFhE4JMHGm3iaJ0+OoDrbdefqFomMSU9bmQy+
mh9Jhbz/I7ve8y1HpGYO35+ZuUK1G0MfFF0GEjFfzQvAuOudv3mJb2GwrWObRnYw
nnWxGSCOeI84fcV1qQkowo4zsMRGaXGCB2Th3TOPF7fpf5nppDR9JNxgfydp+clz
msDpnXKLDqfl62EZF9qDT4/t+gzGJswwmE5+FMU+M0wZBKsfMVshN67XDaJd6F2Z
cT6Gu9zaa3+zpxuN4w0vl3V1Vgf0FR0y1S5uOXn6WU7ma/3Tc8icXP9vjeQber1x
ffG5XH1IVp+nB/XvagqA7uI8OLE1v7QJ1rt/BLis/ZlaxQ4yWByNNCtS6CH9dBdC
QPMq44TgnfQxpdC5MN5IIDUqfF05HWjcHIpsTxTDQYP3kD3dgcFMGFB15T6PgEt6
0zGHY+QfNT2fNHoDN8dqoV3aA9BkM/0Rsz/DxYPr+y7P7Sh7Bnv+7HvfcPj5yHL6
1LjbkskZsHBmhKah0iG8yAp1m5uiYdYi+oLyW6uOnxS7Zi9/kY6ZnZ/pyCNzJOiK
eDPRNWJl1jIlxTPE+kEzR14NYWbWSRSApDLlDWeYfaOHDBUWFDQQmFq+SxwycwDO
oYzEPorpROgqAsNg7oU9LMHT7jHK3NVTxQgt1qYss4PnZ4Zdr8m4b4c4sF12he3x
XBswcFkynKsfhRaMvupyQNOUS6y3vebBTiOvfHWyO81dxQxCFpso5Ljr/dCklD0V
sIwTjWMhqlwBNUj4hKDzqgCtiEsyVAezrNGBvU1dKltMa4F2HOObaitDiJnLNZzC
BSo8EmzDG84xzhTGyk4ZeOtZPdAEBiXOZsxeQ3z/T0POJ4Qxx2iuJxwyd/ZJg43o
tFE/neakt5Cy2uJckFQhGYqTgy8gvrr6G0KvqGVQyfog2zGc38nqTUpogHms8qDD
pPvhRHkATlqlL9EXpKkxh1Jyc8nIktBFKGLhVutWkGkcBpsQkRXKj8yA6FcF8nU9
GlD9xSjimDCexibAF8I99fP5rUP6Y4+mhuVk5ymn7UOdeBlcHkjZZI7zrsJUUEu2
lu/NWicecCahzs8pca0zUR0YaULQGQMuOMc0A0fCN+8g5AzXcChD1W5rSMBXQ16f
glgShwf9C6uYnG2KFLf6jaI8csB0C5cje47J5H/x0qd1vOsESpr4r4IRE3Z8QV+Q
vMlfcS1kyvGWm0nFQ92DxGuUF3iR5VP2HtWdyaBRoO5q0FFBMvjP+dmWpWI+YHQ0
9JzTVi/3lYOeKrf24NlrGBumLZLHPL/YjaN+kpvOxKNrCF81E5BG4tYTMWk+5Kob
uZdtdrONMd4WOfyTbeG0qVI+We8H/xpE6BJffVJ1KT2fnLjr8/7ahOYEaXAjiOvi
Y7EN7V5E8UJKP5/oTwQylVqnn8Tg1TrOKxytMLxdtavKLLvJkT7xfvtO2kYIYkuW
3rOUMWRkGrHyDpOPuxndD9wzstrGuMsCFWUgsMzSXqTKtsDb1d+1DoaS0mEskCqB
WxsOH7WMFnkq6m/FqoHy+ZRYGANKAypqrkV+C53AF/acgB9fmURCc1itj7pNnyaK
K+m+1AyD1LbkqwC8z2Zvj3NdJeZxebqgc8oEFFR3O21HSd4P6aLWtG/Q2CbIezhb
Xf+n5PgjrW4QX3hojmS1vBVTqb3tKPqzGVqr4FzSZ2IY7zAQq5UdEnIV+MweGgPc
EjZEIzfVddUAJBpYPXqnLx4A0PSyGKm/13TQrGC2wzavet/i5uNrz5zH2QGoNPCn
85txbuxRd9rWKVMIxRRQ93jKbiarfbojP2BreDTJyti2DnXZ7fNwZNg2CYEAVfxw
fyEB2Hw2T717fb4LsXxJ7WivNlWPV3SqisZz5bHvJLoHiBGWhUDIWTou7+4STaNo
RYzvcZz5CMxNQwVL+clCcfdeLRo7E7OEJ6ErhG5HpCljiaibhXS0EQd+RPzIdsgI
SAURUZIqJmDKpJFMDADiBKYrsmHR9N/MSWgWMFblvxVAmDv94RmI2fOWup7zQAw+
AlzBgKSmf6aJPC+Tee5TdP1zIDNU9Zp37VbsKo2M6tOQe184JjcAmr3g+4ZGFpW7
hJe+Hs2MJCnV1t8FWAp4ikN8vb/sDaxGwk8Y7yss6hzRwzjc6Vlqp1yBWgrOiXJU
6fau7BQECh5F/QQ/aiovu5nSoeG4opz7aVOn5p0g8dkN9f/wUI0eNZLB+umQ/+QB
OaVNgN0464HH1BRYInyVBGZ/c0He2w68rzl4PlAQFS7yRsNROCov0i+R4AsqpSmX
pTGhe/rTTkI+2V/+wMjF5ZYUlOkt7RTWMhRGo84MLhhx2h+J5P96BkHsndISBLyI
RaIiizUwX1+YLcowDlxJWCoK19XfR3/tYfo3Pdl2jgKD/iZRJ0lpBf2UqJPNwOvZ
Id4PqRvzmfM9UXGxr+hJNZrIvKsHEIKiQV0HjLh1WzCB9vjycFVrw7nl5mZd3vKO
s4VBgaRLsqgJFhAghS6zwQmR0BpXrvaYuj35/S8Gffa8un4nrIubhgmRfmtwxODb
rknvmj56iqOU2OZDw2lUewIsTvSm9h3dt2lbx96JqFU9wqgUnAB23QiY3qqoXyGj
SQqWM/GyJ/CJ1HFmKZjUy+gQ9irFOv/ELL8GDjNfLmjINpvuPKzKUfkuCKqEu4Us
G9vU3wZS4GoufpV2mKnkge2CLwkNVeB87I9jQJt5usIY2K8RDmozCJvL8oTMvCO1
WA8dRJUtYqlqh1TP3XXJFVIdGbE4oeQvAa4Sxdi9AQjRmOotmWaWqrvqaZTY8++3
Tcf3LiL7HRbP1LKpbgX1oKF4XIPiisXXTvXjgpq0D6iV6in4Dn7QtiCfKxyIb9Om
W/6VJp/3axm4Jp0ZeNXG5tOxw1E9qIKxsCP7PqgWnEoxiByLAx40bVNKlB9124JD
pX1VhzOUa/lhqmR6f4iTtE7fLgBG1LISW8kHvnhjv4itL0tJHd4JB/e2aIJopvZU
ECFZEqfELy3s9nSH+Nn0zCtzwDurVFmcVKPqt49F7yNLd6PBsOEmdJaxx0mgSbbA
79zibn+Q5rJLi5vFir1QdE4/jRzLUcKJ1g2anxBFC8+lmEO7UwSL3PZy2MriE6kN
vHy+KisOuZfHPnm+6Hd6T6FO0FpcttBSSq0oW9AI6aUG7hW3PD5zYnbo7qa1Fb88
wCp14/ktk9bXz4ytk1Ow86Ut3g6VrFeQlwdUwKLcIPGOeA3hD2rF91RQIu6xje4q
otYohwBUU78WDIsNv4jLKtdAWIFWqrNcZfd/Nfwa8wEYcBFAG+PH1STs9E7RI3lx
UDABF31YTIkcvOom4umzNa9f2XjkAVtl1MvA/UCgiSijZRgjeEhREQp5iT5g1ENb
xyKcmjZfNK9ynOK/sZvfI5n1aogZDmgE4BLYonC+BiRPzSaiG7gTKW0IxUtrtFZS
v5Inh+IQZNguC2JxeaFc6mWSlV2urhXR3WjlLg/HamTk0KSKf7iODilhZVARPb8i
BpVW35EPmlvtgM5HsRM9NuZ9I0y5HkcYymdinZXap7ABFlxfMk+w3mIg7Td51q2A
icRN9WSXoJp1JBzxfD+DPs0otZJQjjyfo7jSiYNU/FlyunKo+9J53f5tDdHmwtyI
NK0pjhfcpy3QoBitBFdaKIMqeUqvc5aO9yMo31cm9CB2KMt08vHUXpUBWLYo6nM7
gtTmU0YnUl1jt5sdk97TlxCoJgTHTGnHOTpEwg3cJuy+DcNQMUVy+n6K8mYsXS2k
HH926Zzzwj/BLpidYO2oOvi0LyQ2gFqb7qBnglOlEOR4IHH4Ji1N/Wr8172dyR21
dwwSBTkGA/BRwqEW5zzlv8+b6Tq4/BYEvtw1KstMfTzr1yK6e/81bN+2H7JrPj/j
f1PiiHqhhhCx0CoBurO1p6Qu0nMYh0n3LJWYXMtITgQxZSiIGQ/HDgiPFTPQ02TU
MrNJJfYNHxk2QjhNXUlqv0i6NXvOQLcchTLUcGwkiKuLs+gti7Rg64kXX3RmewNw
xmVQBYXrrOel/q76GcNAh4bTiku488evfifRepiS2twEucDP+Eo6NrE9nWqtmuQx
v0PmIt9DOvidto5oZ2/MNYCJvH1ZxyQ2FOr7Q8VRM8ji+9V9NxJsFUhcfQwcfGeX
ozF313FjfL5+/XycfxQJeNnjmX0TLNhIN9MDoKxG3axw0D/ZBT4AOmwmary1YSgg
bYZaZH7R7FdGwpDfHGFX8CGdabSOZQZYUphQMwyvBPqZ1sE0ay7ShbBIO7ySJbPb
w4Zn1tmhMT/6N2pnrVk4jkueXsiRSRJCOMlB/LDZpgMiwRv2f3I3rwigFjDi5GVV
Wth6NRwQSE93PnlyFHZ+Yz191esOeWWYGZrCoDBztZeuT3G+b3SWQ2OCMQoJhFIM
CT53otlnyuVjV8iRqHAV/q/caqniJfQpj5XSIzDHCRs8cQoAY8YR/ttt3M4+swRq
ywMP9SYg0RzWGx3sqWFzITHorEC2ZIMlNHLVm0eADS0i4+uydoV4/lADbhO3AOuW
LPKNKXbTfvoOlWpfAs4Nivw/XG0uCdWlXiiJRqdMtke/XTosDVNwLXcT5B1cGoKE
kuUII69qVucfJYCfi6AkSTlSrVdrkHLkiJ0DN5gmcvvHYPRnTS8vfHyjC5wVdQVZ
MsX07RPO7BH6cuoqhVxpxHVvbFI65YYYyU2CkGGws7a2AP04J6+Bq3kSu0HvFhSX
hw5DighwP+6zO+kvAn+f8J6fl/pQ5Qi87aaH+oY5uo9DNrlRBRjt92jjoVhD+gqH
SlY0Pqfn/vPps5yHVGALn8OvezKcC8b6MiToDknbESQGxv8ZV+8H9S6O8OYKiec4
IuenJya2LieiLG+RCfldz4P22L4S+NqpphF7YEHHYoGhVrOLAtDoZnn/PkxRhRHk
xL7e9GRhPlsgFa8xtQppv+DJywPt4M4+XIWSK8h7JSA6biqzoFRC6Kn8yDkHBwls
g/CJ255vBT1QFsltp7dXLsOfCoGYw6Fec5o6udqyrEU26kOqcVXRFFZY47UVEdFo
/5GqVxitaWzrk24fl38WsZ9AfTEt4BeOzjWn1qQe1ThaP3RxhGFcAdatqs6s/xix
oc1JBQM2qJDZCgMzCubsO40T4J6l+X8Zqi8AB4YLTCeCLu1xIC78vwkTAW61pKN1
U3UKVg7xZKhqagWSuYc3VcmNxNKoutGQVki0F0UN2DnMBrxwS2/rADP7LlOjPuVL
orcMjSdVTBdRS6BkvxPgE3vanyXfS+ufQuJGDn0dMYST0pr1+KH5s5lFwm9FCA4y
QpKetZYFXlHQZHNbPeFyMq0XqV1Wv4hB5684esbqo51gDTOvPmbW5NGhg8jDl6Go
KGSpvlzpsFt6Cw6sKoRFxZEK2v/dMHURVbK14EmYZmN8tSuYfZcUmf+AiqQD8IDG
dg3uBA+qyiaIv/5E79gzJTzy9MsgRHOk4OdmQstKHdFg0KzDGBkue8/mtwzqoaXM
KH4v1OhBUAro90V87XBsMvheKCDnQgR2jKPrMx77mAbYZqFFXcpdoYTnSwsAUV8I
0t7rnCwbccgQQuD7xwkPHZJj5w9RKnQPr5sBhZwFdJaSRI7uFev2veWnJKmVx4aj
EoKogTQufIrPlnwY/jTHENqV2DCFB79y+zuGBK/4Ijgz7z7dUFoOlt5SEsA+/Ytp
5oyrcRpdH/DjtZimcof9WIuLiAmVmqWYcqXx+Y4ETdfcyQLPgUhbs1WTvTxEcdjq
x/LM0FHVFfC9S+Y4PFafrjphyZRKGo8PcAWAiHUuUI463OIGHmv/e6Q4y0DqjqKM
y7xF904cT5IHJQaXLObQp/rgEdIvtnMIw8Cy7vzxyMI3nIYCsia/lYWf0u6hFWLr
hHjW68VPSAynSJDL5Vb0iCraWhL3xs5ZNeE7p6U2eCOoBmuJB826Vb6sFRnmz9Vd
h3OF4TjOKI+Y7UK82/aY/AFFfeWLzNFMzqtLhP3PHfUB2OsVp09FN3kKF04jKB/a
3zG/qqxZYzP6DYTRAdg0M83Ut/wGFJjclmitxfpOqrGRx7D2ts/lFjBW8imh12N7
8x/6RbwFZY/sekWHAHCnIE2PVAvalHLXnoKKn9nITXKTkseazi4JUgyBGFKgijQX
AplIEWQ8MgAWFci6zXlfB7NIRytv+13dewHPWs5UIQHjMdOEsIcwGF7Y/IHeMDFJ
V7dOfL1mIIa7XsJKzvuzRP4oZyHwGRJM9V1Devj7dSvzR3T4wBi2DpzE729U2fjh
GxdAX35bkbgpBiubY+IR5qw7O4WCFXurPl9bBZ09ZWLkSwCUipgrxM7VVGYOFuXn
9IMnW3kitrzu3bLnOYwhZ9W+kUBwJPnnf52mi88CE76f6u2sW7/kZLyjfTeATJZL
frLave7vdHKep/UxFRUVDSU5fPgqNfj9e7EXYAN5vgG7UbO6JmYI6NmWFDpo3LrQ
v1WHi8UIiBdegXgms1hcXv5iD/XRw5fk5vf2M40Xtv96lBT9LLo0F9xdS06GQiqJ
8BFbe90gqGkaIaSJ9JKPpDLJTjJV+dtx3EgFuptvD/4tZevei/URH7yqSOPqXST4
sCIF/Z1QH3TuRh7SLax5WOX2l4OcylrAfVKm5d816++/TcnxkkhDDr26RcxLF1jx
mc0NI4H+QWUA9AJxyfODf24+c2Qj9XvpclbXfEp8BF4/dg4gNIMXNNGIexRY+oXH
dF91jht7gsSSHRlzO58xebcbCFOAw7SYTIHvNykCHZOt71tDJVZGxKlfjYDPkZm2
OdypQXJ/HtKvFIhIRjReXSxz/ddT6ZVu4Bt/AZty2BRle7Nu2EuG9SOMZn9JvN+K
VgEk5r+jkO6NdVDT1ZEIdGH+z07H+5+jXKUPo2LIaF3k0MOPnaNpqTAaX2WFxs5q
1RcWvSI8BLZIMekmWRZaXXWmVAUZFhvlL0IX2C4IlHdn0vIQzS8AsluUpQLwMfJP
RwQ1kpQBD+TWQREfDChLkYPFTNK032PfoykwrDZsT1rnxiXyvLYY6l3SeOstAGJ6
wPhd4OFavnmsI/cazxgsjflLzpluvGaNmkV6euCK3Akk0/Evg30aeu9WM1C0ttGg
Oq8m8sj6hpX7WnKWAwR/Mw5vPtp8UCutGD+07FOJbTrBltneuKOxtjSpeM3tLXg/
9ykVY9t3QBaVU3wTi+iixnGx6wA+w2xx2PMuWub+4wqMMJtbea98/dl25JkHZk7I
RlFD7qaj7NpbMYJLsyVJPUaxSl22XwkE4J53oyG8Y5y/tgkNywYus2eSkwi3WOBt
Gk9NKTXjyrhDdVm1pu2DsSVoVTqThJICPFuWoGLXWmeslbkfCynws2IC1zJhX9h+
ZirltfZ1uqUgvugV/gFPr3zxEI5YxEuWwreSd0iKnE5air0BEZ2gsK+NR98UOo7L
3+oHWw+Az8P/H0Q6JlOnoiTLp8FtkdI5T6RRwXJn85P/URaMwW7Nv5iMjxH9vBLh
KJTDv1bHEa5l64FMosywQN5nmXtGg4UJd14k1847E8VQKM2Q0x4MjYtoYYFfmcoH
hLb2kcQLcq+kx4aB9rko5xC5LnYs22QJT2R3RweP77ksdCnVzIgTD0/00NRilbPo
5ZNnETY03OszqVI4F81y7vCGXrPPCw8bXCEu06D45iXUUB6QHsLTqS+DPV2neObd
/xpjp4ex+UrBVQjB4fEtH6CEybM+cgfgdwlYD0C+dsdO8xJNArQNox2m2h6DLIhx
7vs4ddqo64hLYQu2ZjCrwIwUXgZopBvscV0CdLSQRPEpeuREYFREOuSlfIULgksB
ndOcvLLfSb4i2qP27LJRHLCppWcTfsPnKHY8hvlH9tNAYzhh4QmDbryTamF532LI
C189V4LZzZOejqQ3yRHD5wWY5weO8VjZ/G4T4vVdZ6Q82OKi/Urs9ciRIBVjJ6Wr
x5Gi3JF9ijha4KP0o/6p3ORu4Qk00sQtvKqx8QrQ/bMBKVs16MTp6f04DRFwM/Pu
pLcS1lVoaahMUsTNs6ubDWxbb+F68UD+veCWBrOgp9jiRMdNqKALsirqX7wSRH3L
FmzrmNmUNFhYdh+8VePnF6NQQJji1AEYmuFYISqwvk5vIv0JQ9WbZSV2OnrAJ+tR
6QCh/j21rf/Da83zNCqiD5XEfKpRPE2skBwvEzQtrJpbrrcjTppmO8yTLVZ65L6E
R9OrmtbXWgzwa+FYPudTm5k+cCVwU6kmdLdOFqXMrBDPhvN9t4yXlzYos4ORQ6yT
rB0UNg9dNvnhQwMUMyqabaLA8RqhsNXisPdP2Bnsy8ft2y9HSMOk6H+66Fc/a8w7
upUloQBNFqQ/846P7pt0GyBy+4KfVjPwRaQEz1WfHy1GvrN7ERYkx0pjcQqEn4KI
GTXtlxOWin9UFq+RSYdWslIBky/Uh6AOgDtkQT97R7y/fu9Nv9wsHphlLimfiKdK
ir+oty/J3lBXMjR07MsF1JD8AY8lTz02xCdME9rQvFaLJI1wMDc7EWgbmUm14SpH
W7L5tImd9sz1AMsY81FZrpKH/C0kQP7Pt41lsIRq99ei79QUXGU28iu9omS4F6Ix
fLpcRbk9Lyy7bKaKKwjOL0ea78QlSMyTSigfrjJdUcNeNX0xetLZMSRJ5Rdxr20l
P1URfdOq+wpQrlR4WjGsoXpYugcLBFo3aD3HsJGeGdGQT6uVpTo2LUhp15crVLk5
C1dBVtF7JStrhEXvVbvVWpQxH4RQuziIRK9HlzvIB7NhnMtEmhqtevFriJiWG6kl
Je8C27fS2XfUwVasNHBS5IhfnHOIiex8zG4Lk9y8mBWD0l65DPVKFecNGTbXAewc
CSK84OaW95ryyJsBZWFaEPPVKs8yMjszQ2N5v/uqqSm05W7BTEIxFTPonKD0u75t
O5/K+HeHyJ3KKsC5VyT/CvzBIMvbe2wdbUpNi2JBXZus0Q/6Hfqlma3Gj6pela7G
R40ZZKBrjuxKxrCHo7du5T1n/yD/F09pv4lYQg+gMzFlDYK4qtWHkAlypzUZO0xB
3se93E4UyJBYYe+S2xbvnEhqwslEtV0wtJqiv6/Ko2bhmksbXiQ3BDec4wS/7XmZ
Mv8bAMGzYIl1UjEeoTUd/z/s7jK3ZW6B5fy8eFxj3MkGdJNPu3impgEUUDvGY/6L
618Cy21aSrnwP6/6BeKh+qvni/hirz++/4HYZtnEjZ8rZF8fBdjSnzN96SfdV8Z3
vDXT4s0Ih54iZJ2gq+iAfVmHu66GdcaKw83Rg7mbgtbETGsvqaxpuw1C0C3Ddd3g
JLoztppCHJ7TK+I3kr+Sp7uWONj0aviiHgl3Dn4C992Aq+cBPWK1HQ9PswdLjl1N
Y2H5seiDE2WmmtHfkjf/9zl2gCYJ33XTwZ7i3UvKvwyXUv8QcnwmFMP28K4Yu2rS
/bHyGwqyZWVnKe3zzRsS9wPTgvOIqWZbVIQdpy0YegRZnHiKUpIbay85prGTVybg
B65Xo7k5Z+2llwTNQSwvqQRhcHVhJV7u5RTZ1QEMq3q1+OL3Ytg94aZFOCaj9zMM
RSAJFem6xqNHm8hYYUbG5BCaAeL59E6OZ5Gff658dQF5ziCzUDoI62V+6u4CkoYC
cOJ41Ecx6Y8CH/l0iMMmK5OOxera4NdCxeArU3fJtR0ZtL0pe2xYEaGAH+9fsbNs
ZGB48KCf2JeMlmphtABzW5pinYah00N8iauPBiMXav4CYQwj/gpzu3ntoV1R0k81
0v/3sW7av2E7t2E9CCz7TCUUR5vIyld+Qtf6VzhVVyH3DeQCNMres/vwfEhNJZZh
TbCB/CvN0HvsK51xSFtmsdFQ3WhKfftQqGJbR7qRdvtG1pAk6bGBzqyq7QYRbqnp
Mh/iOUyjFZJ+nzPNzsqvQAaxuXO8+fVDpSBKQ20kKHhCyFTU3C21cbECP48sto3Z
Gg3gNwBEV592CZPYMufUFVQosen+ZthKpmIJ6/hnMSc8aQ6NubBIUZUaZjo0vC4D
QnTohH/AX9FJRBu0PiGKTzd8AEZWW2ZQCIy3I5yO85KgnY790n7PQx0afMZKHBDu
AIa4I/BMEYrkjAuPt6Krwu8uh6IENKPgadmGBwmB71ngoQaCP7qYg5iH46QD4RSx
VYyBl0ejP//R0RhVgQ/sPwVWedVO8pmI/V17OnXjxYdMkkMJF12HzEDmvllrPTbn
leQWTtB0yRr4ujalFmcIf5p2+jAOZ0V2epOLo5K1uqv6tB5XaEeKBR6nUQ3TJ8nt
MPSsLV1pz2KKzTD/H4clgAyHYmMbvqyFXOdl6BvRXWMoamTmwOEu/L9DGq0j5Svv
gcF/2dBYxcOHrqxqOM48WBLPoBFmnlojsC89zZV65X3Z5L5oleasKWxJK5bxUdtb
cpIh6TcLDHsDXX/aCtkCSAAy9q3Fc1ArIDirvSIGcpnTERbOc6PfLrKQLoqRTtni
2+QfD09XkGfpT2LB5EoCj93KjYkmwZc+M10EyD+Hq8bvgkKvjRfnVn7bewcEaNuC
XPWQIYZ4t4TI8dzvOlF4BJn8Hp9HtTePPfmZSx5AQO4QViv37fVw/Ho2t7Y6M24i
XF/dVn8h0gLnIRW2jt03DIIHQnJcnmX1AThHK9pLza0dnrGSrDRW95JaDBXDBIBf
h3L/gXM8lft9PvRy0sX/q+1NqcHoVRFfmFAXJ7LgyupovzaUspJKUNq9sovSHCgx
th/k6spn1y4U3RASkBgo4jPXTmLl4osZnqaeVxct7WEp4cEWeRUSGgIhi5ZFV0S9
/kt/XHJNersSf/J/qVYeMnx0U9haISsxZhuPYHHgmQsHuT/By52oiIhJC5fOWCpW
kjbPu8bEE62CNrHktBh0gyEyZnAbBJhgC1fIRYPx0mWBF44T7OXDMz8z7UkWY3tF
M5dJODDOa885CuMvUTOCZMMtkED/M0unoutm2/HbyV7G0rie57YA6C9DJWAqTKkY
j6buBI5RMkeU+XrFV+SqNknYHgjthMCYNnvPPJ+Bz4Q8sEQ4cSk8QTiM5Ty4T8kE
4Bydu51mWAgWbz5OtVg/jJtIg3OrDzDLdo6xDcUYSRMP0qPkgfAioqOvwO6HaiQS
D4j161ndfmNl2Gv0O3OmCdNNy+TbtOJ4dqe35lcyfI0DlxoteGCt6Bosb4+97sp6
LBIKlhXOE/6dDwjXyoHjuFVbE2Q6CQQgXore2xCa/SqIQuB6y6vhagUfyMS/2eW/
jLNzh9FDT/SHZGAyUk+d5lBeR2RRcEam77e9JxZigXb9GZRt5ZfoCzYAVpWHrZyX
TbyNkp6z/kduQvtx4QsxA033WAyjWkCATNG4d9O41N05Cs591aOEajANkVqReedO
RdgBJgAHrI1oTToJRa6ukHdq6/hZuQnJRU+lgta2y1gm9pJCQPwYCGwkNmcsEF6a
Ysh7v+XkEUV/JrscxQpi5FjQiqqLqP7+COHLR/H4iH4XOgBY2AFznZYu6r9RRtX4
4uZY/WxHWcWyelTqbl0eZasg8G8BLNy0pjNUkeH1hvmZ5atGGHEzuSIJOSQeuhAW
vq5rAUulPzbW2zcq8lEYSqbkvfoLZDEuoeIwTwPteP4KdBTMQgap16jztymEhkCs
gUibv914y+ZLqgVvRS0VQCXX2sQr/zbS23yDyWZLKMGBOtlvSY0YGu+VVRWfCJ57
IZBWtF7zQKhN7zQgybYT2bSpwijOCYtEWTwOvijmlDoMVzdMv8B4Tpa7mj0bjFs5
KBMW6CKW0E9FHCeQ0DlW+T064+rq+7386OimYNJdvdi1Z6CGVI9ENpjPwFnBPUg1
thnIr19D4uOK9n6MsVz59zsnT+9fWUIFdjdRkoMkXjsoDJFIP5VrTrllvBY9tlqv
oNJzEqmVuXsXQSeKbvTTC+ejLBSsULLIZ7LKnGhykSlAeJWz1Jc6m2x1VZDKu7OB
uPH/7mvL3Fx/2Jsm5Ucd8UZzK0LRPl30kljSkOuFPFEahWrRA1h3suBcM2xhPki5
LKbNd8S1i1Uc0hZZbuXriF+XvCkc77N4IozwHgwM0OVFRUzqEURtYHjVbxkxTeaD
BZ8zlauay72b0YIzvmI9gOgRagaNMJBvyVhP1TqzcAawOBJUpxYKA2p7a3c3aDaL
XC5LaSW8Q4QYZ+LDRmuSmCD8ki+qq7fI/OJLrUpJDeatzuiUDBNzxuAcbBNvg3Sr
8Mav1dK0tYhGoR5y7XMBkTzH3/sZaqxymEZ2OCfImJFOh28mV0NcJwgCMjMIqW0g
etUiYoSB/2Pr13fITKBbsYdxReQrkv2GgQak5+lRlku//JCXjI886c37oykISQeD
7h4aQMaTYVT1twxEtlGMYpEBaNhsekJU+q1DCka654u8E0W7fsHNl6opxHTkCUSG
l4pavi03VrGNnpNTXRviMz7XLPbUvqkNFg+XvWqtLITcAedPh++X521NH2RZZhZg
c4dqhw6OIaPQY3Qz5ULAn/3cMB2J6jScmKxU491navDQB5M/vJN0zFa5KGdahLOA
Ruh7bOS1Rp229+Zug0pp0I0/VXjIFwCIshHtBip49QsERkyd91QDfglfLSbTC8Lh
nNMfhTXDQIjwocpYTkSIJMv3lSoTxVRAS2KU+usDQ00KP5ZdwJJ656YgDheKiKnU
3ipQuK8OBF9cnXqR9zSNkJZZMb+Jw0S5s6wR/qIur8XBYmYIryv7Y+GJqWVLgwHv
5rIn1fn/I6Ab8hTkejPGUZNQcDq7brDYZPhLU0sS9Om5JgO8kgEwqP+IbTEbpVud
BZqyKTIBSM5DvOv9b5z2ZIsbujJbju1ZbendCYgLLVVq7mMYuWkNR+IX5rxNuj6y
mIjEjhWTOscxSZm7s0vF7MlX4eK8PJfOyUxrd9dxJrAU9D4AjlxthBtKG8YEpmYx
LtdwNnXb7MuqrOwLrjkk5XSM283nhFD+SAHfecGWBQL1dyl1ufNXvRsjheMkI75y
eBdLcfM917PSqHW6ghJsfvD+Zfggs7bSTjofSsh2uDmwVmqLK/+Q7L89nj5UfArx
oTPrx5unrQg1/xZzoA5rsbDm9Gbcd9uehNzMBLwVcSa2FMgcuHkL/guM2PpQ7Amv
OK95TpwLRs8AZmqQhJwMxsDqWdQZrbrvyvoAVHtiP3JtbQMnBJzxMRkSbi0rOJpv
VoxORvCaKNUf76BENzVmwCMLPe/Ob0Xi5sx2+WPR+jScr/4vqezelDVkgQDw42do
9V0z5MpCmwL7SdjiY3vJmql4oT2ieXr/FD/b+ouTfqoKo5hLNWZymxOgvPB06RGK
IRvZck0kizTHvywfsKXkgrIewyjA1wDalDiSQNuMhWcbbOLjw9wHocOi9GqeQT5T
u+G4q1r4pRTypq/+O915c6oxxazlWbyxHzR69nFVPno+coti5uf1TJBLhzurhvHK
QHvzc+7K+hT9JzTi/6X6zEzTNpLXsXLdKPQEXg3M9RwUn7LcbOb7orFdad9bnTSC
hOo3eLApLFU2Bk7IytHDNAEqjPaBMNspQ7GJTOy3ekxCVuAXjzdLq2bWX/XpnEeO
ihriZuJEL6+BSYTsC7Mvx+cML7cHdxTsHp/rWCaZioxZjIFkY/y4mDjc8YHmQ/lT
5vfoAF74BGyF/DBlfiKzlvUwDtDKxq0EKx1RrPvFhPhODC5T64WP2z/DCZIuy0Tx
mNfH34KYCjrjvOFZphYkL78serchT4q40fZ1kNBbWJtzncdrC+A/EsWIAAKTYFeB
XSaIjv7LA6M/eQ9df5W+lRmR7Hd4WpsfSscFmIM2nK2VvLYqRDE+qlHAqURfNYyg
RlqoQ8UFAcjeB5LvLnmve+LKyxOMSF28fboKj9L1Lq/hbdJHoZZy2bXJEaHA06jB
YFg+ciIe2P3SYh8CIlW5oxB5W7Y7H/0UzwS+aeV6y2JzG98bIlo0euCJXS5RKksZ
iUgcIHmtyXK+QLu0jvKsxi7yK/S3earZlavllSnyaj11uSJP9mNijA6kVqCDlHsu
+AvC8iGLHis/uRX2X5tCr81xkIz/mzep3ln5wlnCc4Xg5rTJtIMBaxnBAJw+bE/w
64q13pPhzwTKuTq85ttbsPUY3PJvY+sQX1/YPgz9q+GNyevskMr8bfCL4iNJ08/0
2i8NBrxLSVsyseT8z/LssWra0SwCR6J/+9HfDUmpVqdjpboRV31J5+2N5aHWbQd5
LhQfy5CBder3M1PFiY6ALOJSJJATJWrHPS8LHmG9Fo9CLvksORi2Q3nYOjo2qJh7
zzwqoJbtC93elFNj+PcYWtzprHfvqDLHpMxmgkcIS0nF5J6sduU0NQx6lZFyq0uC
bL6s52FkXxTIwKX8e7cv9qTFzX2rU/YjSI4QPtG7UMoFmSKuK4xALpAx9zNdFXZh
DvWecAZAHIaT4dM8R5qRJ0bGbiMT86BfHNBxwxFrr20t8po2uHdp6StlkYTZ2qRd
IMq0hGODHRCNEuo3gAsTAffa14dhItDAZbQ7DjYaDOMa/jyym3AlsRajbCx/KG+z
tcxW7lVWNyievoG2tgH9Hm+BXd7gKKo8J5Pz6lb3OYHkLVkyjpBDZ6YOXQ8MvgQG
RFngy1o1JFWQnXY9QQLmg4qR9T+KwfoBD9p4BK2y0qOTYzNuWQYqw0dXo3qBSqv4
Jx0AH/jMaXYU9ezEuIq1xXfeuXM5PRTBBUuURq3Nvr7kmhzn5KNo6dI9SPXvvM9u
udQeW/Tg/FViArL1PItDZIhaO7gRL0uXLhrYIbzqWHayalXZhCTFJgo19hElLZEZ
L7fw2SItmmaLYw9FZLSayf+FH9CPjQ///UyHMj6OOPWHnLFSJBkcO6Q713zQAkJa
21bGvfUMGhbfLBHNKrvWX6qmFDY3hkc6YpBPMTB+ere2gQ+NO+EmPFBn9T1jhgfQ
3cuM3xvZrCD+xRZqR4ZAXGxCNrcjnilgkaowlGcFITSMAsQBUjr0HZRWvI0bAp2b
Wei57/lTupXESQPQjm9VsHdDOG84FEISW8TgVKz66orA2RFNLRjghKSqLKKTxz2d
LfgxTAQhzp68A2SVyVlgV13aXT6QeJ2ZEH5RJMBKCZnUD9yu1S6f17p4G4z32C8y
0n/I5GvJtthE2dXaz0t9RDq74hXn+1lCnxUl6qwiR82vK2xj6MyRZheEpFXxDsIG
5ka8jjty9yB5SOR0AZSqUuGuatJBRe7fXjzw8drSWV2dosuEj9RNyDlTBotn4A78
XwMJA0E9eWgB12/zhKBSs0mGW0nxBC8JKp4FwiYyOe3OFP1xsybju/hCczstzXQZ
CGwMdCCcZCBMZQWbL5IwF+hT1Ifq9uNKa8JNyuGYtElC+7miDBhojzM2kJa8XEZq
BpCG3gGTUIC5OcW9GRUhzXql9Fq0Rytv+JUNVYNhTaVyOcd9jZj+N4TJvKa8uWna
VHl+AS5R8BkLTDD9dheiDZf5D9n07Qdr66MUVue7TzU27tT0mlaiTDhGLU+CRMnw
hHpUk5QdjtNdQS2i/+AiMrPEvcR5nvjj3GyR6MPobWp8lBEu7q/kt8eD3dWc1rSS
PjIei53Qb3ceuE360Kp1f0GS2OmKnDlQ29P92gYXOfB7MkmUnmx0NE/p8rsW6HG8
kVGP3I960ZlmlsMv9CVidJlTHbsbJf3VkZm0a3kfH9yZuwekOMB9oUR8xybmVJfh
tJHsj/Y/MuiUoLg9w7Y1KGNOqTr7jjlHfYzC5zSVikhHnZg5gfGufDtSKFY546tS
coAS7th0PACMA2fstkGrlJFifkcO6IOeHmm/BOVaZ3Aij0AvuPkNd0ZXoW5Tw9Tk
6HsmbPgjTTOEANIhXh89MjH2ZxQST4HxNRMFhc8HmQo6G/oLjni5YS4bIikZpzYa
K3vJ83na6xAiQnPn6sLpzqEVSzaULc8BsRMgElLUMppdqpEK1NftudFxkiZtu6RM
wAEY9U8qbE7FCfbmiuImkDoN9yXPmHi99sQhSJJSJqlDwP7eFgFaUvzNoZ7et0hX
khGVnsVg4ROLxi2SIOJO+yU0NpvbtDwe7Srbgz57lb9tSKx01ILNxSmN3m04ORJn
UmYb8/36Wkjhu3s98QIZUmOuQ6Ep9VRz3RswbZX9nNaH0iwei8bhMfFW0md4qevm
Phu0bD2BrdhTK+nIvvA53rnVIOY7Ufu9mFr2mCe8k5ACXp125HmvGdz1qnb4mxDC
O7ACwLMz59PSwhfjXglpNi4A/MLcEZj2mJly0dcaWdx+A1ZP4QLgysqd3+uhve46
TI61rKDreDU2UNQ3coGTZp4cvGu0Dr7BOKCmR14DSTthzGMx5wRg2KTiQMmwl1eR
94R7Cg9Xu5hy2HETHcwe8Ua9A81PiJs03ElCAE35xYqrEuS95usjUAUBB1yX6Ar2
V6Ho+tCVQa2KvrDP7OjMcho7x0TYW6q9tcO57Efr7/GBcWJG3ZWutMhHR08G4ytW
uRwwTdkPNNnFrrDos9c3KdAUL6Eh0OSJ6yKDAb36HvstLn3cAwMZqSKElKU1MJvi
CWDHxcXRi/FD5DSUIjAbeCv5etkEjJ26GI6vDxx/3VzRASIdHKSaf0qYcoITeAv6
O/kMe8Rbxiq6voXmlUOoEWVz/QrDZxS5RlLU150+AeJvQ3c8m7T/4Dz53hC8r/RF
c1wkOYAfUTegDZDst9H1Vs4jgX+CJfvBqZuXbSpVIH/YJCUhqWSvTUG+o7R95fq5
zM9lAfajP9HzJ1zsyaURTfSKT7oGzrybN9/WBWhcqVm2vEL3Fou7QRgj/2NwwmIA
AEMwY40xcOsT/vHrDe5YjQLJv78LtVSH1XH6X7mbaxWRF7AXeeJ8f1JQxKUuFW7N
kPwTO4sYp+jHiv7LBKK1yM6ncJyW7vNyDZFpCFwl3UCCABecRm/TJqlX5qXBAqSH
aTViSekVbVLcMPJNVkyoAwRO7/DCcaJr1idsWsSZ/e/yN4VKwhSDA6PFUNP6qu5A
g+lfJB9zqwhabfRxwvwdyaIGc15XCWPUXoVTAOSgubD8TC+YaktjUHLZZpwY/Kd/
giY0eC8NRg3JjnhWSJCTWZLtSr/ff/ADGyFNq8wCwsnIL6xDI28/uSOwxYuN87R/
CjgR2+lVXcluN/vlHnGHeT/Y2WiCSSXFP3d1YUIAJMdsJzHZ4sJWat6pU17vFdR4
w+dS4a0owDP1sQDBe0Gye6YJeZcKdYRR1fngtkHyulz9boCBws4lVNw8w0XzIQ2Q
fP+6TWfJ0VVIsR3ex2ay6Ghu1h1wz3AbAZUhFsA728ltl2dAr+JMvP3pgra+Rmx6
Dnuwa8wVFzcYxfAqiURNGLWhtX59xKq2iAsrXJvw5So79asRgxAgUEzJ+/3K8EJy
Q2iVAXfzTsEdiGSo2PO35sNVZzRtgk6HD+Rzkm+zsW2cl5JM5kB8LeyHO0cjtAnc
Uks2dnyp07UNKDm5nH0fN0SL/vJKqOHhtJa2byXRMwvrXUgjIMZqu+T0pEwXMoPK
gAMH4YlksNfPb87rrtWvHHiouNYwOlYKGuJJa97UW3UFR2vo4jy7OMz04CkbtMw7
86Gas2yQW6xp7PY4Oow4ycIgiBCOL6OqBv03OwiTcv4879nwF8VNFOpTFwDYNpmq
phOlD1xGz6J1mSRV6vps6z+k7ZvauufT8OwgG9+iFQN+MK9bDp9iwRiOQnCKi4D2
TwfKhSWjerR1jvD6CfB8Q7EW3bo4/dxYQLiKrSRKYdj0B/m5ihz0hev/An+LTqW1
NY8lIBNkAN9pPMF/YvrWdtSg3n8Js7OXr46jPL87Y6RffQ3KC3hTBRxCwR375Jds
QqqueYeg6UFaZ+jxuimiQWjLTbaJViLN6m9hI5v5b7fKSx0R7Lz67nazOVR9G0QB
NrZXsswhC+VOpIwMXKJneXzIKZ6YKeklA8/DOWiiCzIB9PXhdqx9n0PQ10Y0onnV
A73rX+r0rrz89IQjihTvVz2YnyfzyufkPqes3wwM6hlX7BLbIIBkAJn5hsYRpx5t
3hkIxpk66BI0KaG/Lsndrs1nCj/O4APnQl0GSDsVPvBaI00CMlX3lIQ/nbq4S7Qs
kM6uicZbtaiYGIGCveM2Qmi0JPzvG5b9Ykty53sB8rZeOkZ6o+Fw/wB7iE/WHZhf
PCl4XzI6edtXKrkhzvsgxwB1SzY9o5CD7WeVGoZdy1VNTcxMHpmPVbz6LQHSkxjV
RiNHTHi6EZDyHiW3SxJxh7n879PhA9GR1kdIKh9Mte7AuSRoRunk2kDg1f0a+aGP
TAyscEUAlKzIc3TV2rxqOUw1Qj7VkELB4WXJXCxGc/GzmhhqKM9Me1ZLRRMO7EOF
7hLvRgfbsCWzYmRrwIB0bfBiD88HJKfNkdCiFb/YFsHGzP3sLbRhxxk0LK2otkTb
k3wOxaoTd59fit+7RTBERQKdcmiyW18LjOhpjGclYqU28Nsn9GrNOneHsDJILYT6
vT8dvAvu0ln00mce3VLn7TR/HXcvIiSYxixB4n11L3xfeiBpX7HNH1lNT6dXSff8
L5U8EhnM9A2lokCS00SfBqUhJ15DyQdkpjg/Xet2IpWT8ecoBt3MDuaRxRXaY/3Q
XqaMdhxfg4Krs7iO/bs1oW3go8yOs51tl3VG//1SD5AEU4g4IC16dNmg4rNwP3+q
E9rcPXI0joeLRht/W/z1fXnzDX6tzuVzAtlPpNQhJxxe/s8be/OtMthXFtsJQwbq
reF9SPoYqSN73h3m7tjPT8ZrNafZYWmN/ziZc2CPy17rHE07D/jDVJLz9fAG1zqK
7tdSE9YduL6FrphWe3rbFrpu7on5ioXPWxDsNbpCMmyre+mV+5lL7VAikdh19SIQ
oeh0xlrYG0EvbJu2n8KbASe8+tqMZMvLDXdKWkWf5O/Nlymo9aRF0QPKEZDQmOWF
b+OM/AncpH7Tc4tsM4UzrtdzRGRAm3+B/eDq+2qwhIJfJjfXkYzFRbsgx3lQiBwR
JRQ0CiT1qAPulHbDQUAJQb4hYLXQ05A150Ye7KLVfCidN7nbR8QVtWriTyaErMgS
ZH8FHxArsRnjoFptP1QLfTN94JEc778//HsWIx+6SV5aXDh2AuUU/7P+X5ILqtuH
mKutJF/8p9utyqhpGJv6s6CTED3b5Pt45TUr0cfnQQmDixPzFSO3Pcy6VOR9f7QD
lbtD9lMnJIxX4iT16jV7zIDAt6PW96gwOp/p6783Jxb68VXm1N86uSPzQC4rfThW
kKrw+wFUGgi6KQT/X4L6OP5kKG3jXJNBR0kailx9hhBxxMYeaCUkfZgWIWQlZWG0
8EqsFKtdCIBWYR6I3KUXJutAuNGc81If+8xlp5RmnfhngAhsfkiHJ9tvln4Y8ftw
1pARYv5AnYUOyMGcA3HjvE9cy4XSDfeQar9m7z1ld++Lg+y5CZVuY3pVbOphNdUK
WuK6dbjyB7sy0xp+pxLrX5lrWYSgW09G9Ot6hzrAwOZ8ZjB/o7fndKlnzKKr28mZ
De9NsPix1lTcpqJSuoDidIHvNwhqckbBS6YnxDnmGqMSoV/CKk+pJfHCuELdgHJK
MCxlXRhNjd1fh4fEfL/nhJorUORDhHn6ljIOzQx5wTxOlnuHXLeZbsZiflWIqEnQ
jPylUo/ud62P+io1zv2YBbP5FiJKZ9CW5mNg89a25BTXNvBqHbo6iMCjobG7EB3g
eVddK9tCtv1yOT9DShdd2b4UMJKlLXv/PJSJjPH2LLh72ubIOPOcFTQ8xf+PnZbx
4UfM2vscg/a7LCUatgWNBXftuQ3ODiqOIszHILmpEjihqb2eQPe+6/wvH4gxdcuO
e7oMy1ZDAxE06ym2Yc4QRFtWagV9Ra/JsWCBlK3OT/MGFvrqzvSwzrfwx0uSs+H2
kYDkIcGoPmlUdQNf3dbubfJFfCroy+pRDymRgFNjafa6Me5MKUXqnmaKjW+6knwg
Nj9dmdJevKzwaZyl+lmKZczulRQEa/0P2ZQnGuX+QmpCE0m5vLYcAmafQW+Tc4fs
MbbYROC2eqNKpSEbdY0Hc1Hi3C+TeojTIOWd6rK2K1GInLP1yq5caS7XbJYVWK1F
3aN7jR+3YB4arO6cBzarpkllR5liH62ZrpTW+oJmk2NY8VmQPel/JNkiKzAklnBb
5vkQIVtXFHU941rEj7LF4c2LeMlbBb7qOdTWA9sVt5L8XVuSmJDxMqarnCmOMy6x
C/P8gcZp1QwGeniubTV1eKh9lph7+2edSEx7/yGOrHeA526xt5XNqmL9R2IleI9+
ZiKL1oerkMP1Z5me4gSMTZPXjvVwqojJXJyORUOqr2bTXvY4rH/qS4WdQ+u0yfG8
s2yOSN89l4+ke1gJILVzIXQ/k4zmt2J0x7UgkTJcpovxKVaUJQ7zUJ9IJYeIk6du
IQrC7o76vAULUck0LI/us6OFLR4mpph4HVfNC/Pz95UYkDcBAW/Qxl1ohOfToXWc
IxBJSAvQBL+ygOuUYyYRiw5xAndB2gylam+KpIqqkDC8OJ66Pr5j3m7xdWLXK+yp
ETiXAQa0b71T1QrDiJhuvj4keHLeNRXIWtUYvPJkSBYjKKNqPMZmLBtXrtPUzocs
kxmK6PTf1MYcsgIc8yzprWyAJmzh2NRcxdDPc5x/hhQAuCYgmHw5Bhg0uDFxEdaf
Eg1MGS1EfoNi65A8o+PArWVg4SvDJU8yxouo55eHKuSYtB6fKIrLtxyfiR0rW2ZE
VP6M2sA7/xmjvpqPeuHux0tcU1ihVfaqGoSP7LxSeHah2EFfpuOpNnk6uZ1tpwFq
dSXHguE/9j3hODE7r0VZzdhPtFmuTUkmrVTS68hfU1ruFgq3PYETpq0SM4EZOP8O
vmQzSBchvJrQIvS7ebd9sBegIdZ8zkNx6HcrfG2tKgrHGwHvR1T3muRffJnVaFq2
vSwjvR8Ym85CXreqDpakA3JsQ0mT1GAwxoI3MPjiTglp/7/yFhc6g5A5UiKENCTP
JOE/E5oiQOu5E04KSJtz3AXam1XSmAumVXxJK5KG/jzxSOWTIprPxMC+VF+PG2q5
MeD0UK6Se+VT4qtj7DHO22QCGfF5NfsiGVwtkdyj3D7r4wmvIivrkHWVsa39ffdZ
LHYqha0G1wHQCSjG0rmgmi2WHMh49nXVqPMn5NsR+BUWxdczOVJfi6Ml4ZgqOrPJ
rCWq4GbDB0Z9JYrUcL6lFTM4EtltD48KHSCdRLLz5mFmIKw879uAIx0FA4ECeRYt
nBZGdtLn/Thc2mq1MD3z7EI/M/eDyn0uXPwyHoGLEjbS09NVp/cQMacI0TnPg0dM
35NTQtSkaLrug3ePaKRZCogG5mADoPrQL/wOCuG5+iBj1I4jWi+Fake58ylo+UQP
fyrnVQNsFX2vho0qzHlpMpnUTatQLvZYhevTcc3oZIA1yBzvqNDGR3xy7K3rT6WB
Gv7IWdOmxWgbn4q/XWc+5GyQXJHjZJ3/v5Jk8KWSELRVPUskyU+yq50uJJQUgVVc
lcCdq8HHTYIYMXmN1OUTjqJ9vJ8FP/o/rOAH4wS7b6ZvJLm6daBwkWwLeHtJ9r+k
UGFKVS7U6aoxDcxhuaZOVsH7i7ITZaNT5949/5vnYIOQAvPb6sEvaxFd1lqG3bhe
tV8hWzBhHsR2Y/O5ksi7KOvKvElTi5ZolZ5zCfapt/abgGd9A2+CSvQyu0aMLb0Y
Fi3Z+SCtgw3NJ5q89O+2z1d+d/33aNgVR4Av1t0Pak5edHHp4XHunpPbEvSa3QK0
rMvSHoItGtkQIskexO4impw9TP96jxzVCTFynP7q+JEEJRMZsWELGGbEqN67AQzR
YWjNU+VpIPwaHq69W25kI3ykEE/qefDOuZ4EOLhRwqKsjuGRFD5ozefN4Ii8cAS7
qKhX77yP5YJ7EX0yYj+jkvHbt0u0korg7Fc64aVoK2Cl4e3f6CgsOvs4oy8huykC
fKIpT1OBV8+QVPoOcuf/aaL/v7jqJAkpJN4F6lHyemC1KZvXDkb7/TJwW/4fiJzE
W6S2XHwqX/X1W/x3sMuQP0W6OcKflkmdXYy2BbYxOCT2Qj7+VTef+izRgm95Ta60
ikOEnpupZBwdXRb3vluNTXiYlNuMdHi/h4d3K9S7g2ZY+Klee98F5Fx3+51gYdT1
Jk03e/OvoV0nK08nM6QkSCnJ8ol4+hLtoCjXGq0JT62R27fGiyFWWBkRbEIE2f36
SbZXoa4hyZFUuPnvfLzh5O6no8vrZ+SQuVvkEFH1GpleeLPUracAG9gJa/Il00of
gsUcjH8TEn1eN232X7bUh/4SkVefl9zvaxBfubhtxNmz5MfXthOIhmqEMcdQHbpJ
RFE79kNdp7mBTOHmhShYSqex4emr787xGIXODyG84FlN/7n/m4gFU2hQ4XYI/FbG
bOrt2UrYaIR1gjrI0vtJHCBKiQx1fBdwUk4KPCbRPj2lQ1YqYdi5bWDwmkY6oqI/
xnWp0Otf7SIWsO0c/M3uF/2NRBF9XQj62oS8Phdd8HI89OhCSNuIDJ6d7h8MZ+SJ
W1FdhAyvKh6oNjlHDXAfqV/P4UAinwMjsvafaaMr3llvduAZRwnQ6aGBG8MpqIah
RgUy+KGwxPT85oIOkOl+XM+qNjzkgU03Gmj6NwyrT5qn6mbYoTUWtUX8hw6gQGbb
rxMQPqEfYyo8lvdaA0VQrMVOhPLjF2I7aQiJRvVQSfDc/p6d5GL/Mi2yEuyWXVsK
ZdXslCeCiiiyEHjbbxhdtTi56KO/FmICbsHX42cn7o1SJKlldbL1iTrtkur7IqpT
X/xA7RJ0ht871cXARZRWbqcQXnBSEMG0hQAPmtDKKgMJIxB98m2UNq2yppd7zdtk
es6+ADHfvQI4+BVHDbGrwYG5Xd/K4q++okUfAElEL1tLEMVHqvdpwkqyMlhAtEC3
5dtY0MVMIgTRL3GjX23NvSjXccCub3EjXnDMI0XU5bENRDMhFuzijq3Qbg1fNalY
KTgsEw3BQ5h+l6cBSZqw0BTBsKaGe6iciJPqwPaNZGZV3+F1J0B0WXMNJhYQkVly
4Qaxkg5bykwLDPd0t9HGl+OeVN5CoGQPUFbnpXse6pAvkPDHqhPJb85DoG1Qz5WL
eIkvT5RcXftd8/5hpCL8e+Sk4DYcVTLZZs1jvHUFo0IV6IYCeM3es/mfiQK/nY4k
veZ8nXzIHBCt/1op0ya5lNBri7aruEz6XpproVz2PGK8y9sVV8jbpvWd5bvmltYk
oBEvz9mH9g7cameOEaFsxdFzLxF9cQtXy7fSFBWnUfSACMWWyuy4yoGhg0acfKGu
adVd54FBWxjf7CdFYFi2fIT2YmwxQTKTiGYcRLBMrzqn9iu70kzajw0bCimwVmEe
os2GKSGt1pl0zC9wEAciinYeJV1V3Mr7VbBtrTRhXGVua7+cHjL5q/8dQ8VfB0w9
3GCKFkqGYASOXiwGms7h8ZcJkEqmaiQKJW1pPcBDwNLVtMtpUwjbvEgxTgtDhCj2
rXz5VAm9Bc3LHKXGL3eUeIkccuKT7dmn6Um0T9nXMsKQhY8EUDNLvASNgowZNueb
MxmUVW/eqLiD7taxCqtxX3jO6rz//sPVI50P9OjnmK4Xo+gXwDxdd6+mozyBIXB+
6x9TZK2G+aWyA4KmS4gDaSgRaIjXRWNzFZIgkZxWsj2k1xXuTKDz8OviyUmSv3Kk
laMczfbaUSmITTCLGPTf4wVWBqJD0n062YKz6m1E5YS1RPp0KLEDxTXJK2ee53f4
0mC14oL7a7vihvtbOm5lzrxrA94gTlaEl749iCRmBcAwVvRtMxd+nvD/owHLArxB
dmsscAirjzxCFDEZ+mYrRxvvnVg8Dgch2pe0Oj44xwbUkHL0I4nVJ6JXRGnA5idY
C5UcKrjBJNFmuYs4lZgKmdgYFMe4el4Qhj7AJhpVUqubum07gzZold0pUsGM0Xbb
8H+UskV4zLTOaTf6aXyBrj2sNIBQPBa41slfUQ457v4g/0G5P2sxd9LE9UF9E+iA
ajqouDCI2Nd5QcpdkI4xxLL78AAGu9lDv+OwnQIxUOHKmi+Tig1eLJzj++1p0Spc
5pDHLhaGj+D3AhG8qROf6BOWwly78CszFGEWGvtdPtcqvu5RGrkIU2M2BsIMm/bp
38+xPQ6QDEC8CQ82RZAFOiUYwdRKgcKsw4WpQ5hM55LTQThZrgM11oKTSq0gYk6u
5VFaUzt91o5iG6m6A8ytN2AcHNXscyTi8wWTCYA+oWXufJfRPOxkeMOGqTCCIXJA
F6gEVmOKxFd+CQe+Svf7y95ACnKsNVRqbdi/mOLhOoll2qAxYOnpyXVDGVyOsEFd
UN3pdwNd7plr4MhxcNl2Qr1LlYw8eH8rzLyO+QxNHUbVwNIERoZlKn06geeNGiVf
8Bk+sS3eDgJTP9zYJGUjYsbPDmGI3FNRe+KB5oNTPI2DuS0wg0Elqt6ZeDYJZmIq
P4zhJsySgWoDxtnuEoPfE2H0ki2TwDFSwjNrpbQTAMmQ8I3qt3SjljYD6YTi4KWj
MJhYfvVJ1aQuAFApwtADLGTQfNWlgjd0nIRi0P63QHwIQYqabEsLRSax6x8BzSqL
Ia7WCA2A63oJ7S1cJHV/RktLEKkHAq2EXQ8Wt7nvVkAmP4F9iHXDgH5eJEleRI5M
OE7KMg6TNm6WpVsY+qbVmVQTblpdzcnD85ZoDwy3ev/sT47Jueyc0KP13lY8LhCU
e5fZc9Yi/C4CfNFC4xnXvHov25PAnyo4Li0xmkh5PXokQigQu+GTlzi8lLovWqVK
azXCZZRvbi8MsYh8A1sUw/wcDJBLCwREwVT3duREfOniByoxb2bh3Fnj0GosVQo+
ePcszt+BIoj3TdhzuGe9LbVHdcc27Gimfwt4C0ZjoWPbohMH42pPL7mio1jSijP+
vauDFzWuMSpW1m1GFwJ9NbVmVWLBeD/V0oZwPxDp8WaidDyVy8/tS1jrSDGpzOki
QzKNEEteJUml/C/qOEx69Qgjkw82H72Budg1yg9+pVmw+R2jGMjGNLVfOfwP/fwD
Kyg8He9Nnn01mqp34yAv6R7T0VgZhYeeZSK1iCSw69in0dQNGh4MaEvuLaK12Tvt
opH+FoSOrpDUv0iYT6aSsIrq8EteyJ5WFM6DtxtaGzKcYdjfVD/akynxoPRy8IMN
fG4DEbnkf4PCjxkGy6E4qAyEuhHI+wiyC/+itu/YNNXKshJwpGDmrCgAXYPfCW4n
4u07/9JijxQ/5w3Cm8N1jBJ3yWWDOOS0l0MrB7C7ej+lCymxc089skCMWf7vadSS
J4+CL0azinobM554FItrg0F0wWxplKakT80Y7ssFAYVTd867uGVnxOQT8deYqfNH
MiC4qPAew60Mam89C5rtGgXJXYU43uQhVDAQu9ZsTxPFWi5AVjZdYwQauloe6QSK
9l2916Xg+9A2LO8wUD7Tdx04y20Gh0nmKR99S3irjtmdUmVEWgRc7JpFqs/pASR0
9l0EIRsdMn3/PWp789vempbdUqRnfWjdvtSszv6drSdvsnqTECmf+QfolAxNEtyR
P4ADqemjX/ZsDHM/VIkXn78LFle3Osf7S3UKr7P3//5EuJ3Y+s75x5TpND5lM8yz
PxAah2v3OtSjvzQW2TWuR6K7J5HxivlqUY0+ijfTSF18ypI59u9ZCiRSO7y/+/KY
PZQFmhPqTAugdpzYj0uGENeTnpJoX5pYWhq3q5FI6dH4cPZtt5SjnLsjLLDLMQjf
ZA/eNS7KalNoHaUZWbcgI9ob0gS/dys/WVJ/pzuH+QwbOiOzZ++qLYtFfVbb0mY8
uKgy9uFu+mJT5jhj1YPFM8gEDdu95nfL/4HkxWzw1N6IayjHUhgm8Blc7L4BeUGp
j/EGfJIWap+1dzw1P+I6EXwCDtd45mPE0+BAhI6OS8D3pm8KPiCopRKtpW6Dqa4h
LdZ1onrVetn/P1sFSljZJs5pOUgTjRdgU2h74rrCTI/mixAXKiD80GdS0GDWerHT
bpqDqPcO42Sf6UzlV06bE9VVrRIkXfWggBwl9FTZ0wlweDHIJGw3J26skORgy2bc
7JCB6EK1ZV0/Qd4zXfQpmYLUURMrRKcFZrLeFL07QevEMdyaRwskiwLxtVdVeA1t
sQuOzfSrvFC1M0xervSgVD4PkiS1oesNwEsH6sv/MvYnt7xOqwDebYTxzGZ50rZP
bZypV/PXw9bPKXrI2uOLJafVnAyxznAXCXT7rtTY5wTtLW238Z9igOI1FQvCBlWG
3NlZX6+vOdn92nWdoak2x8e+e5WyvoRcKME/3UE9hEWO8SPkRlx0feRzd40F03Ed
2aMY4/bxzrc6Rcuv028bHnBgxO7vbcdC70oblngZLjZLgtpMp3n4+Y5ohQZALfhK
wDhTwBs0qZcLUfvgJYHn5APMtY8AQJkm8F8EejbNr2InUn056MeqlNM7ddzbPJkB
dU3AoYRdDKdY/hL0ZAgFXvQ2YLKHOChH80GLGlspT4GcsPf6rAY8OspdzCaYnwAp
Y13zXUT1qw/izG4Qeux3KElNi/nLy5TEMH3umwXZVGE2vXSICvr82g2rZw4U7aeH
T81x9HXk2IIDaV12DAOKQwIpjJsWIQ8hTG1KsjmMGOSqr1az/YFcakYKjcvdpf/i
4YeSTh0sYbSkYAdRGil+nwktZ23q28xTZvjptyPlx89TImGNxnYWrE+RWPCDI3cQ
iQi20789sRj7YepwfaXAWCsvsGKhVhXpBhmYO34cB8GpoIiBDdAnGijlYwm9z+kj
ZQl0uSrES/3+yAJEEkX15npvzABPucSAx752kxYgEGOWEFJbDrMByqcVEjntQyA8
tvPKku4w0lFo28lIVyHStINFlySbD8RhvvY1Bvx0pWrM6rEDl/pulUmNcoNphBEn
jzmZQqfh/OWeFXyBI23sfqkqeoq9rIBXLNA23rS19LqubSOMow9jK1XHp0J9BnpK
+akgL01gsP7zgMFh9S6jc1yNJiX0q7RmLtwatK1I3OeTxchmJH5tY0oNMttXMzbD
+pYGrnrjqpUYwr5GxtDnkaJxhgi+h2+LA9p5ED+ulV/Qrr0qfKlzQv264UY6/Hn3
fT6j5oynZVzwdbGJv5JdxoEgnZyfB0TBqii2M6pecRgd3y/lq05MwVEu9lI22BOq
/KajghJyiw5kRF4HBEWpsUzzKPysFr1LpU9+CHyGoS6O0iHpGEYrc9x0TsgW3HgD
q3l1al+jC5C+Oec2mMDwNsRjCD2v4vMtaTYqkTqPx4yGeYa1vYTjqHKydWCrS/l2
rkQhvB3HpwMxt3ZRU8vs6zke9ydnbgJxEkmQDc8h9zirEy4OtnmwkMn0h6R+tfPU
LRItb/05WHwpr+bkOyEF46ZkEraURDaZW5ZXqgsWdlCRVrELZdQ3nVBe1w9tOwYB
2aTjI2Fl8oa1G0Go6LRRlNurIBq8gLbLonxhFBMF8Uvat/zJ2KSuDq/Mh5jBMJeo
48RiSwMrQRZ/WZMf9MfvZ7c6rR1nXVNIKG0tIrQJYSWZIzoizZn+LQhSz8wp00nQ
orDsADCYMtAh4CTU/NluNGWw+IrjHRcpf28auRpl3lmARc/yHdooIXcEM5Tcj8LW
1smHvLjajTX10NwhXdDaTektjm/S9HTQnN13vn/NNS1tnw/4TThREaOAtFDpTKUM
jpgj+Cl4HPlQ+Su+5nnpcn5Knf9apzOnaC6OtrJ+k+UbFXK4AFIWih8iyiB7IsXc
7lUnO7ItMyIUWPj4v7YIx7xgavwf7gtNnBEPXCfeZ9WogsZdUNkKNK3F4OOrtLZa
nDqx7kSwW4yyyI91+PlgNpz9fKeKk9devXa4wJshJhMEzsf946yviYHPnsOxtqp2
vN+nAMyOOYPi0Ln4TCEW3tRFKKdR2Mb5lpEQeBWTX9EqNDsA0vXIUyjUd9S6VRJt
xqPQyzI5BKxVIVK9LQXKJkkD49bS8nsY3FUwHEwThlx0NVhUQ+UkyEqTvv6b0HYv
CWw69gxRyxKANhAECVNwh0FMgHsnf03Mea36nRqb1nugzsUoxGl05kY7CXYY8z3k
Hs+1XTLXd/Ma4jd9QZUDSkO4LJtd+ssLXYwkQ5LuxZbOiAUd0e3wJf0cjdL8pdUg
CKiTxzhjunQrJtxEAKSFULfSvosI/He3iuV5/LyL5UGnvxKToCOh8Bh/u72hqiQj
bVIIrbDRdwcM80ltfSxK55yCUKWB0nud88Z1EZ4cAMKVt963/5iL9nNh4iVT6qMZ
lKMnD3PJzmPMge07Dhmqd1py2ux1ZF+yBV28H/eaqWza+GXB5+d/iizk1N6cGlQO
hYXpOYpIeCc0toO/1IAT4bUWM7Akev9lgntl7GkOsGbPKuGIQx87usJj4QoM1IDf
6t0oPUNfFYUhkAkNQqTyrR5D+LiuMXpU2NIwuwf9BwCi2IyPeGQdSPoNzYqlCtyw
EQWPlqCfQrYKH3aYOw8CsydlMYqwKBY2sCUO76K0GWS21NlERI2SmnyrGRxMBudG
S4ZsCMhL7UpfjiuXM3ly8Sc5TEkBxVY+ua5MuaxMIjC0V5LG0buGh8EKzXRtcpVW
lJsc1XRh7tUv/VVHvcWtAPrDJ14cjEzr+67+ULP5BZ2p+gU/EbNwO/+bCwoEEvSW
cnm9+pubwlngRnCAlANGN87ve32qCMXiHP11DPpX/gs63IyJCgoa5neoqrwhvxey
p76ntRZJA8L38WyLKXaGRrNImFi2D31zINKbQotlkIUe9bVMz2+qBX5I+A5beV8O
Oe2sOsrjMaxZ02lP82cuf+j4o3ZS2VL/CMy5dgVdi+7N63hwl+JM9NC0Gd6asd7Y
CA+kwPCvsHt4zmXPDKdjgbC2FeltnXQTgm+/pmyMelmX5sK1dSI2Yk853iYActEe
ytJouyDMvYpkraNCqSjMIZdq3cpiXqhAKMV364BT19KrXJX0dMaJTy5a6ru1eyde
UoYgm3m87UtJ3MwtwlrVAED3Tfb8mFhDmeQqydUXNf8kI/m13VOmEERJzijiURiF
hfWQdpZil2NNNTlGc9zgbl6wlJCMbPXTXBpLL8HUZ4upFygpJQlqwhtl5/fG8OwP
GtUieSZ013mTHx5Ec+oWdlaqY4DWrhZ8rdxFs7rOALJqpraNyLnkHrbwia3OZWKT
8gmzyTXGYwdhCskjDMcILSjkC/IHH36OOQeyK9J/bArYAGU7nVaqs1D/IIlTDcK+
j04G7SlEPzcIbQJMBjX1wmUq173gpmvI5abCt8J6R/kG7fXfAiL5t0OmHSws2VmX
4EJt9OT8kgebzvxASWES12RkhD7L12TR1swPIU8UcE5rgljcVg/GV9sPt5pwQvnc
Go/w1Npb52tlbK1ofC7LT8Mf0q/PaWmKV68TVAOLZgRV0+wWv3auj2Sz2I/yvZdc
3lAub8133O4blUrMIlh3+nU6GdiKBr64hBlws4IqeuQ/qnx8HxclDb6kTs7xJohp
KCE22gkGnflqz4xzqxGThFuyuzbvO4kEPR9t8OAFIxoksQsLCRv4hbSwiEIIk7Z9
XHlf+daInZsG097aua4+izuvChGvW/r/+w5ooc7ramRMGEFy+nIQzyIgFhCG2sue
tMZLtwVPh0oqhfabcOPUqjyNydZlhs2lpFGKpVv779qoHUDoBpb/uuIK/mW8uO3W
ajwGhGUaf5iiuvDMfSh1TwwKUo70xeEmF4Jius04FkaMcb5UBlczsN2yVtkLM4st
4of0fW/zNGQsQ+7MsV9ogkp7AAgM30R0ORZsi4zpQuX4vkZ2NiXU1EzmFwizAdWx
uYDDjJXg4BpvWOy3noIMtVaEB5hqLKqqVvrPT3n3dmk2K99m3dzd+Wm6xOwKFFno
6rgAKpaUbdiOfNfK/Y1BJ6iZuLhjnTIGRXI8Nq/tc9OF7U3xX05c0Wa5pcv0BMlS
VlOUVr8chy4625QIg1ADfBz5eG5e/eT4BJ2UgowUYSNKPHxlY1W0CD11qi44KMjZ
obm5TrJMjuFia6v208H0u7K00lrdIdC0kzdUwuGeD/rt7Uiz1j5q1y2xzdhROVF/
WglvKzFQr0LFymFlLJmDJiTujRmfoCQ2uv6XMq5wBn5xCWGIFmdgnCD4Q/S06wL0
5UtdFXrJrTGESOY4K2gzx1j+xfX8cl5wmswROd6cYDTCSwceJLShaPUxmhhXtOB1
5ZeOgVNnIQEO3LZiNuODj3whBgTeiOXqsCkzSRtmNi5w0pKsENt/vo0AzUSBegrQ
NzvPmiEu/6ekE2/Ds/tR0SZdRi/XIF2AoonaqR4laKQyRTnmM9rQ819xT1SiCOql
WNsfkNxwABdFEtlWiROAD8cK2wYFbBvsXWzFRMA7LtfIaX/BOvl3sWavuyYVut9h
jSqgMIGjmSh3MKBwtsAGARExy/pgjU52yZy8olY1lXfK2y189dvnqlDbqL/tYkwY
DGvjZzPCDD/6aktnvIzCsQ+0gnej7WH02kBy40CbcsxvYj3EN3FzCinK/Nu3II1v
+skgh8nD1tMjvuLFovo3Il+3CWZgnq+vwLVpd2617IoGphVBPKJQq+jxCqNnphxt
YrSjXOfK0aGZA1uKeZV4zr26ZlV/I35Yg01mbKULDoUttyoFPQytC402tt+laQyW
sksSGEa3GU/G4VzGXMCFeqtoTgbpol/1LLX/85pG2A0tqfcZrZuJJsBC5k0IGuzc
OaEB+e1241UG/TrAEulzjgS1bLtj/uw72CcoajU1xUOExpgHiUJwwTs+o1Qw1/Wa
h148IgcUyawrK0TTlIe+xoqXWPE5iKJw/q9KjN+kMriMAFOYVS8QnihC/xAtjjJT
7fOfM7mEOvVfecMw4fJVNY5veHBHmbeEKRCMMTPCzV0gXJpslt2fdr3hFePtOqHp
vwmXW5Hcm34UkhKC4Hy3/be/BAlO83q55EnuWH8Y54PnZ9CYejftxO8iVpwlJ8Gd
RtxnswMd63+bai9qaMIjxuYspnd/BkdYb2eT/88kRjpsGJ/i2L7IOwqCf1OQczeh
wg1pH9yWXahlCdZBBkwRYNYxueMmAihfRdYHqXgvHqWqOUiCEIDMwGa9jjnhmePX
uQ0yEGFyKu/+4aPJKY8ifNcK77BZm8jmVF4HpGXyHFzO8dnny0p8HUbpLAtFq5vx
rgWdX+p1gJMBmAdYZc2woswzWT8PJM+SIx9S/y/52iS2rp37QJ+uT1na9twMzxqg
nYwu7yucR0BnIc0CCA/IxINvnjekWQochT8x8JSIPFHZLMlRE0ziqyzSd7jd7RwE
c0VY+pga8peSv3My0hSF5ON5DrU3DldBmzYqrFVmWjYnvF1QwqKUWXXxACmy1z8g
A4NG1ttE8QYwr4rett/mmg0fk/Bq7VtJ7Bgh1Il10WQAf+qtgunJz1QEoUMt6+3m
mcTpoZ7a4j37Yp2NN73YFdOu86V2HwofxRqcQ4k1yxG0f+0pCq4HQrnePcO2LAbN
yhWnTJfGixpYAnf8d7xdHU/Pl1IDx1GBo1qGmDeODrVYJxVUyPMIZbmbtcO6OHjF
a/vbRjaJKDxb0/x8aGazUIcHxSorzvf40Zh3bAL30K+K032NiRG00Vz4JT9mCgaG
5PeKxBySUVNe9lCY6+r0i0gloiK1614uCSazwE+Xf02LeOBkXksmOAjcVZQyL+UJ
qdv+Q26F+lvytArqONC4ceBDoYg1BZJ8P7jcUPWHGveXTh3gquNiGXqoTj8Ju7rd
o99/hs3az8QtfBrJivwtpegeDiJv3L/wZyoMX8njvMnivnQM0GSRYOpPyywap5cj
EQp1ZQ+vD6vHtO9xlLTLLssVGxfY3yhM/5LB/ZESnIrNJ04cuyzE0mpGdU/q47Ug
Wlp3F7pj7I5L8BTjUR+u/96IKzyyumBudlA7hY4weIDbht282OaSX0vLa/vLvLPD
mZ6NPqlwPUoqJQVOHRV7EfsNP/c4vHl9I1cQzEcdKzuKcWW1jXQm4qXxdmN0YJXA
jMoqt5mraAqyL+ZpvNlaxDET6JrVG+3QHmZLuzy8ZvfqOyRx2cDX7MBkTVI+wEgI
+im71gLlzNz2uzbcd8jqIk8aMglMIkrQUqm6x1VeFWQOgfu5HMXkVmuHCdijKsAM
3tAe0J2sFplldhaIk9NQv0L88i8SSMLviHhkYFWME+rK8w3PDXEbxUi2y4w6m/Fa
2YKwOs8EqOYKYn/4+ZEp8aDPafbWiaM8H07mSSIhQV36vQgWzL4oy7T5CKwLD2Yf
smSjdfPeWlGxHl0kXztS555wLRojM2x1x20/hICze/IaOBSxHmkYZwxwcCcPvzF3
dLahowiIPL7Ph3bzDzTeNZfc9GhSseyj+AAh5j2QaQNQ56vqGdY0GmUJTSaG7m1T
Nqh4Bm/tbrjmwxjvrxn5oWReaPBPwloqZyn5TmFKJ05h8Q7itoA1mqVZG5inHgWD
KCG+x3kxHe1h3lQBceOuprmF7C8yXCMIT12mXFT1ks0MdZAKjrJH+RyiQBOeBaiU
8zOkCq+mE4R6kT+q5FtQSt0dXVQK+fZJDOqCOKxYHa/dkZ56Sdx3YMeDfraX+nYI
DRNF27Oik3NSVL2/U8S7k+GCT3yr6EfDV8JHYrnO/wGoLUg2ve8e0L1VSNRH366y
/tCmlib8kMk6x/52T8xYC5kvFkkHIEW2TtztqUvZ4k9IGR6buf/E3t7gy+0lpMfi
b3fyjg8lKKjgHy2Hu9qvBuNGFfCXIEEYa/f/B6Gm43OuDy4OZT1RvkhN7rDDdR7S
q8Dvg7qRw7phZg9cgEHeXZGrgRgFc+IHaySy73O/Q1dydmZzovEmmNvVY8rUM23K
r4ibOcyjsXyfUUPlYD55ZIfmt96knJ0E33I2i6esJ5uqxqMk++JpOFWKU0m9EKVw
5L83tkQzJw03KSVlTKO7NtrxjqL3xHMko1X2er5ZA9lkvj/mreIE0qAY7yhF3Wlg
Yzl+iY1qVGOnLWpyzuNSTV3A2HGBQeRwoi2zhEgbBI5fodZvpmpEt0w+CPJyzUi7
lS87DV8iVCSco+xmE60bDTFSY7hjxRGMJwpwVZ2mrbvpVma1zRI8sy0Kosx7yPKI
N7aGvsfxFiqO96virY/VtZeWOootIQ713uf9DL0RRxqgPuqMJUcS7Ss+T9C1r/Sq
Bu+1cqzljVYY5MVB6RKswvCGPX6rHM5rulZORdY5DuYst7id5MQ+PRelx69U7Qfv
fhQanFe86xYuG3gAH2cewDMWAAqQo699juM6dUQi6Ej+3arrs2ARqtCE4sGl5Vpg
WzX2IZSpSW0o/T7I9RaggTQD3r0Gsc76GmyzhGz8klhtk6QC7gg/MxLRXHP64gYS
Po5r5+QJXdqUTEV030ecB5vboCMRfD56/Wd6CeawhqQJS6OesVS6kTdNfL2NFUA7
6jAVzSgics0BXrVLpaih6KNGlSvqKjk6RkAavMGW6P5W0kX7E4M+/eQAD9wEWD4r
j4wWV4wSPBOqI0BoWRZW+OuOR5xwpV/XRgSryl+4+RUM0ogZY/WYUeJPInGV6h0q
/KQh48lRQBGR7X0jFirLsyzTIv9GEpSX0SJekBp07uLA9f3vYgKO8TC9P+fur7x1
rDaRJbnXd/4ZbT5kHc1vkgM8o6mqvliAKWivSDCLeAdVfIx0wSm8tnlkyscV4CrF
eamtNsimGGGw0mgw0nYCVOd2cXwg9MTxEDGxrATRBtgyx/FOFSkCypiQykOUT14c
pAe/S7GKHGeZkLJXJCv+Kqc2wMDCS82ZMwYvjHoCoUhrso6u+YlCMI1LYvoKAzPe
y0PmcK98F5RljkLFpN6lmmDdok7xwJ6oRUTdkBiQoDWHj8N9++eouhCJnjRj1HkF
gOECpSDPR1pfCreTS2iS0XvaMwX+2N7fi9mqMKXiO2fy4vbtBfka8ieSRK/VzZuY
3o6pdqcxkWM/Ynb9/F+dTRSPeiS2yxl3GseSCaV5C+EP1JOq+euLAOPJ8kHxL8LQ
rRXbOzmTJTlARLh6pXwDct8GDJgCQR8BAqwlfu+f4vnX1al6+l6QizadI+22KxZK
XLRX+r3KQbP0ibQi2SaHtJxXh/fVx5UB3Z1ygvyDcsDfAlFBENjLPjJElvBQ7dD7
AjBodWFjJvM9skZTscStCkamSZjTR9eodmKv/SqTdCMXQm3TJB4vNfQkMIZ9EvZw
C0mYXNNyUb0rVApJXVBTya6ztM6+vIJCO0Rrj8YUXTNBIGxpPTDTmHgWwZnPn4XK
HpKF7y2DJDRhXapnBQd36YmhfJOPGAPoKKp03Jgm+WcTgz3OvrnzufYgA7r6ybPw
tyRFNwKMaxKgQZOu9fM1vHbMn/ovvHvEHTVnDb91AXqFhBmKv9zD/F5eECCPydA0
dLP+JAlFL4lpVCF06CmfT4EeRIfUkOg6tifnk9sgMDCCAfIag6xQL40W6KFHgkjC
tUB1MJADRzb8XkvlPjsUY5hT/YhapcpTrqBWy/0iYXdwv6MAgZtCLF3CNsKgYl72
OXZHtamp6E6AHswj2Kv4Dp7hAU2iYABGZxrFPUa6hMxYfjqBhB979pUL8t2c43dX
IxncvQ7FOKu3YC6hM91AobMkfFXsNKGxpntU4mUO4u+iD1cwjwlUDPHTKQOK6k4L
An5sfhLh+axLnGRC5vSBO2QLcpVHQennNHBDFJqbUQ36dlV7ipzVn0YvJXPQu/6m
0cs2YlEbCvterm1HqifWqscemzUuFPKL/lzgahCLS+m+ftaZrKv8kT0fpARZiH7e
Xt8X9rKLstNM6qKPgG62P8b9JjjjUcAfKLfDq2eu5pE7BGJZ5cOanlOl+ekB/6lh
LcIPEO36+22AuftQOm50pjrJ1fwkwJRnTgOYlayhht3GPRX6R5wKArd+smeogYdp
FukcYzNpXh3V7wI1Q4ud8fhMLqeOEFbE8hFG0wFO7KGum/Jhv2zY+/o+KIuSAkJS
5iPf1NIkvhx8bNe+Ll8fdCLkeR//wGbB/mNgUmD1zagvVLCWNxAzJW6HmXF9NtAH
Khkyf2T1FUv7PeH4uYYU1kvC5f/jI1aq+baV6XslvDZhuOZsM2I+MVn7qpnSIYPa
KJNovcUtgkfTgWwFiMgMrlx9sjwfMS+wJhf1o7JcN5a7vLxz2qNvbK9Ho8NFg1Lq
khZEnd3/YSj5LdqPy+X7MKpCQoKAcMeAqrC/bNq8OAQhOaGG81yFLXTFGwa823qe
bITlX5ydzHcda0od8KSGgqKxl7M1I7cAOxNhx1RV3xpnVW+05x0xElpv9pawLOyf
8CMX0NM1b138tlBge+HLvKSejffNSb1ZUawtfyLwwcRtJxWcpNDkSsC5wd5BcbT+
gSOL1pg1yEyl1VWMNE10Nc9RW1rUDVZbVGi8FCSubushh81AkKdJ3gU8+Nj5XgaR
EezeQIhKbyJT2AXQ05F5vCH926LFCbFxInXTZO5czJSFLhpWDAMQK9ONzZ2DRMDq
9ElVOX38lkW3YhiGivonwj1AdQ0ZZ1TP5mZAwdfTRbVDEOdYDc7j9b9MVwaWDPNH
ggMl7tBEC5ThzWc8W87Gl9EXy4btOj0ODQGH1NFUWPj0yufbHGZ2rnpr8SCgo2eB
LrLeAtP8Qt7lP675knGCLh0pxhRUvLHiW/eapIDD1E1Rcj6I69tAumdEIxQF8XDu
/O2CjvsTEJWzY7THYTbB/19aSfPQmSO9oXMf7IRZd2a8hKolNrJOqYSz1knFlES/
6Tr2Eih1F1hsjDSf5kb4vvQD7lv9KJ3jH4b2FfoewKadIUa7YT5JTzbpg/GxP0lB
wWpq6H9Pvfgp+6RYEVkHenrtpmxfKqHFMabNwRFoHr4fCHq/hKiA1dv2eBNb+GlD
8hrMEDx+PPj7ouNg0UYDf9Gn8IkN3BjY1Z47eUz1dFmkK0tmVBfKl5shB3Lz100E
nc+PfKIxD4pNF+sxWw2a5rRevQ5xB/gZmy1aa/2gNYAyV6Y34A+WEeDGbvTu0u1E
uju+uVoHrbL1TFWBZ9v7LMCn51ah0+SgynCY+klsE4/mqBIEerafK5ppQ5GvoeGE
x5zFlg/jV5PUZtROWgA9GTeLB2Nq225roacAq8AUkPnipNDhnUsby/6NDp+3pE5R
kcUDuTtsMotBPb/eM1NVJIOychYtjSuWEgWKJfLAB0tToQnQZrSBt6JORIyK3BMP
nkIL4R8N4XSQigzpnRvC8KppWAw2tCQXIpkjfL3spXSFlcpED2tVL0bkeEoM1BbL
g7k3gR53EiqybVxe8sCerkFOz2tg6jT2+F5yGSuKNFlCvshKkNmztK/8aa7xsD//
Oahv9IJMJfBoThYmJxCLJb4npp4vGT79tMXDci9GMM+Dom1GVNsDISHW0FnbD+3n
xpc5JzN80gyy1048PmI4OgAPeWXezSBxaNTv8vA2Vy5Rej/QpWR0/047k+hyTx/2
Dwn+ACxntavzOgxK1V/lp417x3NLAnoWdJt+Si83bRyUWu19Xlpy2BOSCLTsDwE2
3uZ+zgSCdJr746ZOaeP2y09fxnu4gEtwjsQ4AN4Rqj3J9Xp3sV34JL48gZUATlFO
scOz/irxu7bRqBULl9sLjLplZzYI1lbSwnrdLZdrjF0Dl6bBkSprmUFgIVS+0FeX
tm2/MNJ7vlAmY63T0d+vYs4iMkPL5qTCT15AaUypmPfKnqmYKq5J4RyXOQaIyGbd
ombBiINOmWMSd5E48E6lXOy+H/NTNVQ/ZtHi3wN2dmXsBuLEnSah7YTfNphS4bnU
7DhWuMa12KiPaeop+dZMDBHtyTcFrjGuCMI9gK9R95NhQnCi3CuL79qmNEHFVi6d
T8ItFmdq9en11Ugd5viVFqM5NGgPN4pQ/eIirLP+Gr5Zd8AomnyoJTAMXr07LcxN
Qa6FVhJL6U4nM7oV9NHhF+i2fe2UsHXoFthI1sMgqbMZ4vG4WhdlkI1p5vCZys9v
fUzJM819SdbY1sZRL1w2IpHKFpvXysa+Lt1HGA7arP3zjOsKvvLOzL8KYBqojAwf
TRtPkdih6Ql1GNvfkvgiCiLCHEiPxDKHTamyfIPNPsD6mSP2TqOt8ZEpY7tQo+0Q
jPFEbEgXAfwCbLZQkgEvlBoUfxwU+O3Iqc740XP14E1nbcn98hXszBsUzaAqiD/d
K1ZgMJYOioBA1f8pIf2f0dXiRKAM7oolsVTEK1d8P2hFAYt+Hm6dEbxf50/YyYDY
sVnOx+OA5b3Pd08K6NnPSdIOhy4Wz9JVXgfsMtQl9CNgiD7y5DyX9G/PW2hNuH1l
tfWUcCW3u5cq6eJGceweaEawSCfrMJgkUkNrYcwJ2ovXLzVeznzqRXQ9IJrfbNmz
/5cmgmz5WlCnBpy+4FmewWEEX09jTYkw3fe6BSlTQgu3pQ23Kb+xBZk9b4ihUWvT
EtfQ3lXbCHuwO5kdiryLaWohtwJkxredykr/EPvSkfuobg1WmRwMI5zsScmgbtd1
20mPwUPK29vibOJD7J5WNnFL894hvU3rpP83/AQZw5mAjLWySgs4hR2IWdn40fus
uVO0vzBm8wb+zIn5aVcTuUOMP8SOAs7q1uAxdgrM1MhCz/UWKE1rSpbBmFgd9TD4
orCSYs5YEFagmob8dZhcjlefPLwlI3V/33H3msGiZQ/6i/SGyjLepEAj8QJZ98zL
wDWXxbtiDdxnZWQGB7gUu37wNs4HrVFZbWEhl8KKT350c8gk2imt8nd28EgOIzhj
ZkWflsoVoER6pK7izHzWukukg5hVOgge0DUD8W3AQ+ziHUZCaDWUoNeqAnoi2UFR
l8pYeBrR8P2gYE1cQ2BBC0jKzra3D2ffEWNptKs7PsO2LHncd045O8/2jF6dszDV
nax2PgdEUp7uIrNRUabdyNannTgeZ69NOQmpTXCoq+pTl0+lyLHPe+4xtXmGnlog
7eN1czN2xquPa3jsubTTJEDdlcHj+eTwzxv2ZLoVGqFAZt0ryYnzZ+yWEhyZO4N+
WgaiwdhChXzvipwnku+5z2HMaFiYq8Y2u10nRZ5OFyP0vBFCdxzGRqoSZAeWwiqY
2EervxBWWq30iNRqFHS/SxwQHxge4VG6hGMADGtXxY3EUMtVSenClo3toiu4jojm
W6rqFOdSNJ8d9c57sANuQ2aDDxsMdgosXENOT19GDrGp4pKznE9Ni81dZHSrcmDH
u9o4XWB4vrIx2waKlBk1+ZgtQ2jbjnpvElfholjkkdrTW3NFwRmHwJNZh6Xwjw2G
KTNedxpL/SC8L/mA386du2VZ9psLas14byS1Vu1WF5V1CqNJN2HRjKTOCpwqfhgf
grIc5sMe3eqBNsQyM11f/670qwECScXela4wGSM9Mv1Mv95WkLjhjsE7hv7RjaRY
8PMrEiS5eSdtR5TefdmoHQASXcv1HI7DxFSOgQ1s9VigkaztcHKJcmHXIW0VOezw
YuNkDRhp69KdKH5WMInI+g96fzLY1KduOjHD/J5ecZUPd85aG0Pm/Sb0en6AtzwJ
TIJDNbe4IwR93CS5zQcprJRMqSJrBRak1eddIGw3IjoQBnEmwhGweHLYLaB84zD5
j+dWayhOQXpcrRbDQXg7FN+Qg8ZuLR+vejy+M9ij/+WCpC1gq28xbKv6wUWJEdNG
PgZ9A2Xo9Kiq7hqRGVDvRrWHemuxC4K3cOhFq1JQJh/kX9Cd2DHeWJOBukw7kJlp
5P6ZGDDNVFdIOaioLFtzVl/PdT8TVS5rNvBN2p6NHmyRQUBKmczOj/kjBilyx57t
TGdYXO4wta4h89J5PHFLrzb2LdlDJqc4Pdr/7nFJT5/x8UUTSzZarHM9jeUE0Ruo
MCjPakPyYCmNInf2rCcEMHIfDwi1v3F5HmC+4hp3bAEB6zbFFLstDbk4qih/5I49
m1oxRYQRIJhpx1l/Y8TRlWVxHNF/jzu2I+PjB8THgr5J48ezWzsmQAruooaMdc3C
rccshtPMyT+78oQ9v5bjqVEnlJl+lQ1t1bozB8Z0RHJ8qI6H0mUkDrbkZbRuRxp/
1gX3XE8yDjitGkFao9sHOWq+y5hYHBu8dTqju6Lrq+h6FjlNBL1Vr8lsC03R7YWA
zuDjM5G5JF/FbyUpNeOZApdg4bV0kmyfUhX4KtV38GtB8foE5Bhh35sk2IKlz5O6
E1dCWcaonqI5060bIlOi1ddc+fG4FzcLy3ptgtHzjWwAH6hamSwgb1fUh3s8EXxx
I53ms4ZMuUPuq7h7ET59AcWKzqcA+PpPNDutyIJt4s3eta1bMjQ2pE1V/DhXn//o
cnZ/MkDqWok2flFhYTc19AaqwQaFyCcStz5zh+ZUQAaIRQARIm2GI1TsMkRGJPES
pQdazAGI5Yy+/BbZ9oNHWvmiCBjUcB2YwJ4GmItH2m5JsEN9LllnORY6JRxY5RZs
TgBHtiwnL9x1Boiczrdt6pwqb0TQeYzpIB35erjqQZA6/rigxWhRf+n4b98CFy1J
GtW2zjwdTA/QBCeU54W6HmksipR+S6sWK7IFf+Lk/Rj2rTDT2UDS+4GSojUKQ9rH
Z5VZV8hfaj5KpRtE0xeU0InyG0/d+o2CiGMqsknGQe6cJwx88vRQ6noWc/nnkn+3
FBNY12BUEVdQyROvHp3PO1aM9q6b1ylzwIF+50iQ/3UtzpCccNqnl1xyA/qN+Euh
Z15LNVhwxW4vGm41BtVqLFzjhPmlngF3r1U4aYg3fCB5TqsigNUzOyhi+XKMHkUC
xmOsB+SHN7e/HsA+UuTvY1b7HDt4bsKZML6VFPbVHTN+UfBco8UHCtkb4tN6xmCT
Eu0PsXB6ARXBgA190usmu94DVattsuabkrvpRS4O83aHulY4qbY6zVOXtM2IczzY
CTaXQo0DWfYgUaaeGk8DR3ST9c2XnMgELjC3zIH7eAWtIKI2hTAcd5TRDrzz7K3n
l7CHrt/jr0+ALgvwrno91brmMsbTrDhXcNE7ifx85dSKiKel1QNQFBu4V2myM4AY
5+3/ZcVCfcexjyyXEdRQoCE1PfSIAKiRXgjNutQrZkzN9wXylJEkJf58qHAxOKIx
zWltNeCtH5gfa5xJ4KKQXpuJ8a7CcOrwukQY3VHBOlTqlzLkPQtoAxDiCYQz824y
n/H7JmR8f2a5NefX8a/BGsnrFgTRY0oJE9LVlSJJW/77WgiwET/zXs3NMlU2brBu
3aEjpuV9lIteKwsUW8HIKqbSQejVsCCXKbP6l2wPhYq/FFgmI1eCA4to2+H81LN5
qX3ByRbFtXP5rajef2//2fGkZsfb8T+qEzhCwB/N1cZ90mra7i8vsuXGH14Hftqi
mNjj6HMZJKNjejea6bEY8mzGrMAeU0dBtlZMV+OWkeEwylYR1hSm/WjnrbkvjUTL
vuM2D0G/PkJrEgltfpbFRYAQA8Jy3vKMyRDjIyn5us/leLz2iP/5WGH6hSs3/iGS
4uYdq55QdXBtCu5839FSRVZgLVu0SI5AClJ+BQ5Gk/vwHZfzN/XjKnhkSCuB/05B
nEsK5DSHOEtYBe9jJyjrA7pMiGKNBugYsFnCM7vjn/V3RZZhpb9zaS/0tIPwN04u
PbeTYDy5LKTideg+VE8U/BlY4rRYrDkGRLfdOPvno4AnJIU3eD1c/+opHv3kbHh7
1WAM8ypXW5urJXtFPPDOpOlp7RrwVtHbt3XansmsRYaeRrzQOH4yAZbsBTchYZ+H
UFWSlIGCk8F9i+RCgrGQPHzl+EsaEzPinTyYAWRj2hFZL6WtjBjX9TgOqtx/a817
uHgAcLomjpVmjwyWjTN9+r9Z8DFc/9sdleYq6dARmBYzoVWLg/85dG6sVUGZT/sK
9tWOsWraUw0yNNLrhtdDMUpgtdQcMz3vwTiJiKG28SP5DFBd0QEI3kw8bF7SE0vi
PWFwFsF7mxzvm68+S3fFD84JUTaIB7nXiRxjXk5v9Q1HSyx9OruUXZdP7VAAnq26
7ka7lBdFRWZCbFp78rwxY0WltV9JSM2M32wOKCjatFGq5X+6ARCrsiDOoIo7mKxD
8VAuL2+sjVuae0T1hRlRMwdvjqkZJb1Elb6E4tfw4TBcLrg1SBfVhdVu/0aYwbNl
JVVlprzlSo7LzoHccJ3V7J4lj9TX3Q+Z824kNjzEYEt1LsTnhpydn7s8WonaiB62
A1HD1yxEuIB5HLumrb+0wZ/gOg/a6/Hz3j7gaVD6nlx3U+aJ48pXCsd2U3kMFnPH
G+xjAHq/RYy/GEC8zprRfbvlSlTmqz/sCzxwu6NTnI57REH2tDEY5aRB8mcznUaz
eUSw/8eaccFqkctwV5jKZlnJOCBA2QgaQvbCSY6fR3267JNRuTLVGJJeXkq8Tqcn
Os5DScb1BVXHbVkQbXuwsAkYbZthp9oNUk/5766hhGj1nG8sDZNMtr9eAaneJi/v
F3VwkXHhobu4NExHHn13AkMznnM4oIiaP5UGojpXfQg7GBMyR5laabMax4DhfgPB
ObPLawE4Fu6NoUYLr0/RfgU55uucuWjzr2UsnxPLrX4TYk41CpvfX9anlrDHJB1m
df2EDdAvkbLu4ebxvtfzm3S1NsrAi/lasym4DhFz+XiFiGZPjRs8C/KnNPM0sKsA
I65EXAuIJka/OyO+WIu42QYJWohZRv3HKioMDlpdGErkCCGmbIMxNl0+bl+SQ8fK
5igvRixXXBAJyU4zu7VAJSc9Np8Dh3PpJyZ/5HGhC1EIEtuEYjPd7NWmMHy6hvrL
ORHIzcJk7meerX09eBIJlPEjLTPkh9qtBBJ+oZbgFR/QOPyrcYc7z0/gkT44qiw1
aD8FDHaNApuS7AwUBTcpZJl0AML208PkYXt/RuL3fbfJekO9fcnWW4CFvTjWgcbB
CJQh8vKJHDDJkpR+OrCPjuTR80Ye/OdfkgBmH4a8dIAfKE4gTSdLNiIUB5YoLBvA
AZuZbBOekXwtaWeyXEo6FBGbRIKN4gIMugfnh90OZ3BSWkoc4p56JNMvRaTPhBpD
a4V0sKyB6G6qoMd3nk7Zas3aFw6NoH9ql0RIqqaWRIB9AEHnC2IrAIz6nibOGIyR
HU9zRv26bnnqLatqZ/E+Wr3Y96UyLjP1euYel8uyMVEsqFenY+zLwR6Nc6h59LKl
4mtIBR+9IrU39n1hWcJVr3QGjH/Yk+2YKXK6cdZE0EqYShxSl5AiEZoi/h/oEmV3
2NjzWxIJ2nt53uTPqcTA7wXuhg6I18Ymcqhfwf3oJGBu+ypattegb6qIe4sQdnpF
onQ86cCRmMzaPsdpFxPbfBQ95GC78lT8j2XB4+aOPSNH12s6ivSteiP1aJUfgVbv
rIpjr2D0Gjkvdi2IuSjR6sM9VVv4Hg+PuVuwxHMZIl3PR2la4Ec6y8fFEhJuAXln
conqRiZNfbhtT71HIwzRPxJtsdc+cVI6VnNEtz5nVv/+g4kRhbP6phDna/ldWR4O
FN6gbFnFbgnxOLeZSEGvvQd/SZDGmNFHjLH3O4FZ/vwCu543jDRV8jd1IKKBOQiv
NVel3VEWespiBFPYPHYTgFlGYfxlecMf6Xj2f2RE9U5o1kXzt+qHub7eCopCBQAT
5nfeMsICdXCP97rbneGZzq8K5I51bTHg+7LxJ0iHvqNygHjMIUzbQwqK/CX94FGc
q4+lqoVwjV/DU5MpTD9YwGja7GfjdNTrGt6tfnVORcvydVUYF/9xTqFYwES7AZ6P
LonyTwst4swo3Fhf/3D1It9scmFTlhk6JAVp5FfXG2N+Wmt5zHyhSnlfvIlJtts9
PODBstigvq2Zcf1QGa0Y6P7qXBut17tyO8NxPtwx7I2QuRpa8HRwZjYqY+TUJBvL
QFR4wDbgR7W+UNcDb9b8lvOR2qE64FanRzExMIVUZ/0gGDZQoP2rQE61mPxgQY7A
+gAYju2LmYywpk/8XUJBBa0a+14naAeDQrPcR2TQpI2VwGwWVHLUDBbK+r/LD3gK
w3QajtPjbIsmCGObdPNa/e485cRBqbEqg1i1bR1d8SkU5dor2UilZIlifE21akHE
x+H9uLmIN7e979ckHjOAFE3xD56HAmPemxWl63IPF2DsktHfQQklXlKKF+FOle8Q
mduWlEZLNZPFs9xbxXNP1z68V9oyq29NuBtQD9EEkXi/noB2+3af4DAusjglT3be
z6ayuuhoB2isaxZLhVwNM6znGqqCrgiiyWuKNKpZOvqkrXvKhBzU7KR1ZOg91kiM
QUOorHCmXrt/AAI1TSojtl6GRE/e9zMRY9TPRp48BjoVUTPu9KcpaJ7CR80v1LE8
5gEM2o9/J5TXSxHKKqSJU58GaMiKpI71z2ukFqlOQ0PlTMMR35hVz6VIOHt7F94D
qnw3eahvTap3AXYhn7ICTfrmIErIzCJNUCyctApcK2A5Qr9d8rMKkMXqrxvk4ivv
EPtuVPpXUoSKG23IxW69zRVjeTqWPK7LFXWWV2vwEdmKvekWQfKsjiAmP61wDEDk
nidhcLugCREfsQe9+2pMIxlnxCHn1rTQnF+xgeGtAwUlJKvigAnW89GtEpH9KM1m
1D0UGGy4plMpmYRL/EircAUyWULnQns2nLsRle4X3Wr1d0fKuguoZOvRPm/rOz90
ejaOAYJIxMCkSXx+hGM1OhaU7mdVLl5GdVxQCtNHLWbh7klf/frn8AAB84uSttMM
jzC9QnBb0esVRLRNDyM7n6oSQ3JAJglXXmawN93OjRSA+IBGdNr/Fjll5c3jvWyl
OZbsz08J0YPg7bzRiOXZN7bEBJHn6XQi+dDPYM+aHlJ4MnHvPvAs+/8I73AtqWRJ
1sVzLashMiUCuO3NH2Jl2xJv6w/lO/ApKvL1HUpCY9wC6LXR4HnYBrTcBStzfA2b
E/y+sMoOJhQu1tI+vw0nU+pxQJERtyo0jGAnHUKWj2/FAIbhXkqLBhqEKLn+efp2
TMxvvT74z7PkrZUT71DLhedRxes6i1QUzO3baWgn+SpRcxiejUUPdSoi+b+87vFt
d/B6U4d+sKXeduHfbtVc/q6AnUP8iOw7JZgcnMKh/ZQnuSAsPluk78sN9VSqlDKO
nG+frkRIOeecAzfyT1aZrYqQOg//wRV9owlg94RgX/Zg+sgT7o1r8SBfiAwpvURm
B3ah1fRvbLlvH+IurX/l36VhFEjo3e/HBZSbFTZLDfL9MKVuOiZObr1Q07nEPveh
tvYREy9USN5F0USPTvqAElLnQh3mEpkxE7BT4KiIrzsAhDZnjQPxgXbs8rCYpsWT
sRVxdv15xfarB6AtqtTOEEbdoLyne5T+IhYwKO82Q7Uu5cvKhZGzcp//YT3uUm09
SGLAaE6RuNN/brFhJJN8V8NKSBUBXuXaS6nQlHKiKZ1KQPZU2QOJu73rFBuesHQd
/omtCeScxcjj3kOMjX7lhN5aBR2gb2W35b1OynCdZAUnNw8QkpZG0fdgVSCz33t2
NhR4b0txP00FogL0reV/FO2J5GqixYccqnqHhUJrk2nf1EQRlkA70PPUpi1AHm7o
CM6VqlDYGwDwC0N7lFVd50K18sy4jaFLiGCpvBMRnNO7H8dSQD0iy+sC2zgrH7Z2
OVhwkYD3PvBcYtcOBqjD8JJekovRJwEtXMx/E6hqBh/h9z49M7x5vIxHOy47KhVU
Cs6FTZ2HHrTwkUsPXs0IKdrp27xGC9wSj/abiKM338gVabqSyrUN1HhAkWOMHJHZ
ZUc+X5WzoJcu8G4zJ7aoPuUsdeh8jpOJP90Pgaxj2bL7bn4wlUywGXw4AF9PXNCI
rfBatdf+rOYz7vR8JRuZwOmvMvbjHlFOv4fiFoYZQq0Dpmw118NDahiQ1Sl7Fn4L
j/IlNVXLDLMUf8JdpoCVjy+FInwuucFouoeBlWnkcSJA+8Gy+mjDcwnkvMOzGA4j
BRPvnG/f5iFGo9gKz7pnGmR3XmxPoMVVS27UtMDj+1iCdh2J0m6E4X2o3A9yt/Fk
QseOFwNvu4yyyE1xvBTq6sdfqVZM82cy+51lbu3LgqalffEy7TDVnunLoGgl3LBH
aYOiJr9CfK/LRhX39bTx2USSJk+hMd6knRuzGM5m7NpulO5qHRqInCS4zbleewjp
AAcx4UgrRjoeiV6TZK98U78PKLTHJlZIZIT2E6rkGv9LkK9lNyw5bk6AY6t3nr22
78aBG4bZSkxLNeA2Y7QKvoVuvDF0pTqNQ4CMugj7MzH8W8xoJoHrZqX9Oa45JNcN
axuLTRnZuWROy+gyGDXL5LiN1kJ2p0qMjTuP20WlCH86xgzfSn3oR7IjeabQscvZ
gSiPEVun7gbADXcVTzNzccgJAH54KbquDA9197wCbIOsNqqRTQmuVTFtxLZ8AvmY
D429iFvZJ4LDC0sZoAzAItULv9EEzMsW0HQ95t4IjNKzo8Tqj4GuvEPtpVaIIDWR
FwZvsEplAZA3ypi2BkDyENmc8X67Rq03Qy3iwhbNdejGzbXUhSdIQIzKgoQu2rfp
V3phBDyA429ErGes3Dux4862R4yZ5Hk5e1zv50YUbDktD0c7urY9xEjyKNx4jKyZ
uxcvz4dJc5wBRQqbBIksTNi9ieRdDAkkSU65ZPec+Rt2JXuCS9byyehWR7h+vCzC
yUQC3dLwjP0/VbIfD5OduhHkkxfAq/ovQUBNNf3hBqTxOlrF6shLegZnELht332N
YvKk/gu0xUvI17MrhO0Lo+Se3aZrFkl8eTqVHDH0+Pl1Ro/RKkp1j9oUiNFR6g+J
zQTz1uFjWCHyk+M61E63DKiq00ZC0M5QXvPWA7ZreDQtL+cAEmg8g2g45t+k6qRJ
9Yg4o727NJjwgBQNMjIFne4xcyOl4gxfJjh+F7mQaDw6tuvyC+xgtJ4u/zC0F59G
kUiKQcqYDHHvw7ubuPX2jTNfzHTujST+CcPpimhNn7AU1fgAEMFYhPy+3+cLQplP
DgiqImyMFttOzyZmI9VkXV/215HP56EdF8StVZwJzcIHsMl+48HQ4kHanP/vBQrC
9wEXuPvpaIl4kYT7Dyb2Oz74JVwo7D8cF9WnUp9sSQ61ewt1PZiA0ngzlTlWDDJb
35elHQFR3CSmLM8Lv2KQBvaF3xOAI66+F0mnMyvC590u3mQ7IDcaG3nTu89QP1kW
kSP/trMJ19opv1Y4NmoQz9RLUc6mNPb6FqjAAE+vy6iPj4V3lOAf2L7fXIoNDA+a
OnEifCZ+sCB77LO6byO7nrSjL7S/RnaPLL9Fg4zoLnOOQP2U3vEJMO7OqRD4CKcq
ToHzUFI88QN0XMKLpjd0T73Mfhgs9owj7vUM6mYQ4/jO4nG0xR73FI7qvBkN9WAS
dPB9omvmkiNy+SwcxHrsKv/snjAbbh/AZe0vHohpbjpriD2WJOL9lauM4dUheCqo
DUUvvSrllaghEYOaqOiUVP0ueSO/8UglTakcFRoXlUky6DKDs7di3CiGVg8fO25F
hISZE0Uvq9t2dGssZLJB1BXgvSGDTBlN+kSoDkGWSadYcTedZVT12kxcEPdCju8d
F7YjZ6wwwEfLpq3t7+o0Ver+ry7rb+9zIYjLPRT72v9n281bXriFIHgvW0ZPB+6J
QdVRK/ERI2vQvLKY+oRwFBvTO9j6dzmSkZ+c6rK1yECfnAQQ29pGXfoH0Iv4QViF
kz8tsdXlKnALLR4GYQdxG1NbgQq6jM+fNpkco3q9N6ZqHBE9KvlwzJvTdIeFiFOi
yGaqV+8ijjhjDaldJ/0GdT1T835XcqIurBjI98lyraNNNhTKUKLPe4LJ+8ImTjA+
HtonAlpAer3eq29Eg9N6AwvMCrcgbYbZu6TSH8vc3v+JTwe9qN+D4YPPD7+5aMNP
dsDePPBwcabydMPx0c/PbsBsI9Pt94YH8+226f8wlMmFfWgbQwPxxvfcwvl1BwtO
o66xN7AWbUh7+vp0oXks/c9Ix+zjuWhFGZh+S9ddPTG95NzDLMWgf5dL3wfDoQxo
vfkLgw87AXUrtAWjjuXMMGtXz3daE/wML0R8k2YC7rrMQQ70GotMGA7fqE7Jt2Ex
6j9x3vgE7C5Tcx3k21pxsL9I9Xn+oTeSXkzYgKGCXYdYk9/Y8IaflFDwmofiosnU
fTx7iNcY+51Xdivh+J/OrpRpBPdda+gmF6q0QqyHOKNFpAQtpIy7iGXTruDEd6bz
aglmwfYXDh44bWEAQ8BUQZhqyM41TtfqJbbs0kbxNATnQBL7eyusdnl9AMrbAk4W
fqpGYH27Pq65zbfvrnBoD+lxzDdJgzdETexZtPLq9xcVbchZ89YD4thNIWdGl2Ff
qDK/4/0u0528Pnh7Qo2Oz+1SLN3dPXR4ZRjUY8GSRS/wUrxERIN+8qkaB+xVxEbC
YeQ9++VqyguS/95IxvjbSl83J9dBmMup5BBcTObZOZpx7TQyPdCAag2hokwUIl/1
d7O3vSuqGNaZVTxqikFE29RN+WXYV292UTpbhHh0kCjtOKJLIZQR2SHwgT9Vx/ML
ccc2jc00aC1cQrRtBeiKhdLMrrIH2hX9HSqhMIJIG29oAWb5P3iKoutuipcrjExv
Z+RnFcayAFSyo3w31Nf13NnvH58g9ajT/Bz3Bk8AvjGl69eZbM7I56S+F05ufWUS
3TizIDnA6xZjnTpB96G8f+tLdj6Uv0LbIrwQUzznhfenBIvDxqcPcdQj8mj2ZfJb
4IuOVHClbNDY/62tc70/xC6rhzoumwJAvCz0Drkcidtz5OyNFBsHROGsIUIDbG2Q
07gCFE65vkD+FI0hXQd2ln3cagXkqunbZND9Ta2TUykgRKmdryDmsOgwFHDt868d
z3qr/tm+oC2BQ/iuDc5A5tpPp5XMUm46WgBamS9DZtzSYsVAHf2WQG6j7mBqK+l7
dxAJdl3LGY/bH9CnAUElz0L3jomglf6/Z/EQq8bQ0qvSGAWbqQOMgjYS5TRfA4hA
NMFKXJ0CLoAD7OZBbhcrski6Leh0ykkjtHC0CaLWKWq9dfYnqfDvD7YrQkzhbtP5
B4b0tEtQToEQI1ErvUfhbv/go/IeWJZQ30UxXp1VKx2KIu4I6dI3wfKlwRnrEr9L
cw/r6548ksBxOhZWb+lmKxOUMd171za4oa/cGoywZNogUpV2hEDyWrLgf2wV0y4O
Hu9nDOJzrdq6OypLKmSCgtt9YcBK4ZROxHxjM5uoz97pnb8KYhKGILqyToYXyPS9
R2ej4ei0MGOJLxSNKEZICvhN4ut7f0cl+ShmrxCfAjvuk7zsGpjnQ3/p1UXcLNse
BF/m7d67rHrbLAtnGPly7CvccgfEBroYglYgH+fD200CJsSt/RWT7oAq2cKjLl0L
OJ4Zo4oFEshplisLII3WX0ZOHW4XpvSHvMMbgNjGT50WHr8fT6Y9KiOT41H+04ae
cpk3pSuI6O2DPjF6MdHaMGW0R9DjrFaQL5xMeKoZtaJ0OwdU4ouGndA7kZ1sTWcs
zZ9QLs+xi+WD0q5om5zvEn7XjlizHaQbMu9fetMfnVzZnu0haPt1tBPU3S865vu1
eQEtl4LS6oRQIsrFDg0ki5IIXg4G7P+zSrUnV3lPLz+0zweTRSRXItbKQJP5hSRc
65QuRATDE01mXMdJKUe4Zz0zL6fAyF6ugd9rYkjYGgLfC02pScWNWAi6AFbeyYgg
1ZcYTLlgW5ZUR9EniGFTZoYEe7SGPOT7PZUCrZ/ZXPvrR+BE08IW3iD3F3k6F7Dd
D0RvJgGuGNva1sJmm6Yi+PG2EV4fRu7H0Jj7n0MrzvrNEFeRXYBJWynFFmr8lMxh
Noeywc8XLV6CkC2D73+Di5ehaxRfYhSWWBgy/pld3PdHiYmVq2Y+/yq305j6uWx2
tLZ0QwM6DdsxH9V6VhyuS0518blkvOsDT8u2+n3eJfpScT92OKXGkM+6LJoJVmES
DY3nskcXWCgDeNDI0QMMSBv/cHUA/wJIRTvbHNXkoksxDKBueK/WnyJD+AxEpWlP
MY0HS0QfYmDPMdJCV0L6+BzrWKynn3gf+lX7uUFevA5S1FTnjYyI/AfKJB3rJL1/
ifCIeP5bYiK4tdKRiDwd2B+7Je/7vu9UMtGW/C0dJKa6dVly/JJpymKhv5hZtnu1
qVFWYT92ndbMdMn6oU6BMg+iFr0hpVK97OXEK0Eyx7WGlZm+DKze/upZdKRndb8D
7zqVTOmQnIsEYrkvvcfub6+h8g0QKOoC7TwWxHHQDrq31uxektvXuTCypw9qK2B1
JI96lVMEUy0UP3xjKhge9Od0qk8YzoJpGgBNZy4z81UwQx57ZJBcAq77Lepzujri
MF25/Oikwj+cTpa98VfCLL202Y4z3CbH4eL+dkMe1n+rIkkenrYpy/Fg+ac16Zkc
1CCMChu2VbItfnrCniPRIp8ACYdQXXegIXMdIYuH8is3oiPl13k2u2w2RXpJqtoJ
AMgL2HxwxVN6bL67zwD4XMZ38efTlL/HBdWjcZnp1c6RN5OO9fLEqDoESeciEIgT
EaDlIQOGrdDNLOudAQ5y1CWj2oV4jPpYOTdRc/j/QptfO/zMKjRPHSajLPUg8w3l
0FYFjKJAVTuiqT1LNwfQDNyngwv8szROvjeTRuHElPV+Im3cKy2Wi+Rk3NWXakFo
pdyN2tZ44n4HfUkJQzaq3PEMhE5jplCizTA5zsXaCBCpfogDxkKNALS18LJn6Wv5
Uuj+2dJfDQ8NKFEfBlQqC6q3egqAWD/CQObUVyobJAtKIa5eDcxxSy0suRfeHWlk
7LdStyI5bzHVrGhbb44q72vAa3ZgMxMeqZRDaBkW5r1eC/SMBY2Subjhzm9bEYA+
9btVVwbv37zI1tSHWsqdg/cpHEJssQj/x+THDevYFlypYQGs1X1TIBqPt+CRS/rW
0mgVtWxRx3bsoGBwjiGy+CujZ2DDURyVbCThs/zIMKhMeWs+HZwcBQMX0k+WkfRi
8Tp8gNRTJe1rmt/UDwIDjFWnhkpApryWotttjn9tJ+R/TG3N4srpTnu4DqZI3Vua
NLUmKbykz/84kgaxSZ3ylcktZ29VtuGA+Nh4IVxnXkRFnIGc53SaPUxD8dofI29/
fHbFEnXyo+3rHpfZdbNhJqCrrKptHvIezKoxITQEpKGwtWoLhBpB0eQ/RUNgWZKB
nfpvMSidIod+FTg0bsQNgz4PzlmY3VW7N/K8FGrK+7Noy6KWGbuIeCVfSShUUwyx
y2m1dXOWkCpHsPCi/vrevu4C+zqPNNnWmvuhOaFlp+DO+JxqAAOvAEM1RtwZW3Ps
lx0xYiFRuCOZyCGtX6OMWnMSGiY/OCI2VOhgftvHpNKmd9HDdoVDWYe/WV9dzg2M
gcAjAt0jpv9HxscFMJp83Tkx99l9o7qLnIz0z/F6QgpqNvG/JAT1Z54f1wi0hVl1
1c1fJXvCE2C/FMwC0D+zmQHZhpUSg6NytlmgF212jwI65sARcU87UtVWYGdYpV11
bwAZ8xmrzDgjabncLt4ZF/G2hdxS6Pw+XjV3uHjAGnJPB9j3ALsazk+nLTzQ50Po
yMJ0b08uIu6/D0zLtWz/6ZnEJYcVhsPirNgrTz6YjrctYsdwfHWHpDppqxe92QAq
Q4sb/nG92bHM0jbSGasBF2fmjMzZd3ri8Y/pHWRrfzErH49H6wpASQSU/yIE6GKy
+VX6HibbGMhpnq6GEDktPiKUCOjNl14Ns0E3uqFxY7p2UqUucGA2zpKhlidJG1LZ
D9y0tjUEf2wpv+QM4iB77pL9AdOJcsOvhX5dopCTK5n23pfg6yhuZ/H4/pwTlrQg
NSdHE8RVXyyCYbiClfg0Ecalx0gd8LU7IbLSKEZ2dj35My+FVl8jJcQqyzulAJJs
Va6C/LqvdsGpfu/3LpFpf1G4VSLeVaaSDnTH7eiciZPAI51aMpnEGbjwMa69BPsN
h04sqoJqZkKz8YFSpfIkT/8fVRtRwZzx/tFIUPrRhij7hLWuKtuXIYepvWNwSmqw
Pm513zGpiLbMyILnRZGnu/poduchwpr9CzyazOzBDc5KoCC3x1tMy+dadHi2eV0l
GNI/BUYDn5feU40iVxbMhLPgCT9mBwQmRyEYHPkoYPSzcyKyBb6C1ffia/P/ouJ3
IPWvVD5wuzNvf0M4QWUEWoF9tznzpbHZ1BDpAjExBXahaeajrqpVyWwDZwSWYZ2Y
K8GchAsPKcv9UrCwsWmbL+uPjU7QFqZqaz21VJctzduQEb+mTuLBD3Anrf3sW9IP
ewXTQVxg8xYBgZPHiuXal33EMVluNoIaJDiSQHvL+pRcza5oQiBvLKCaAj0yjYm7
fj7+4QPzBAvBQWsz/Q9vNKKKkq6yAGFeUVa4RzUUu9eJLaEN+cHSvk2b4PIB9Xp0
SSHePWRDWwgv7C/Mlv08ajevKDvoEJHL6H/EEt82Sm+wxu7BVLNiWiGqENxyciue
2M12kRSR32PpGDW6ymS7zZIzM6W1jUsPgxYzFzmeh4D+ch6P9x+/QItKvyZcuIwq
+Om+bP22/SuWKQJryUSfMLk+amxhJtqLvkN4oJnu80+ShG78jviSBi0s5RQcIARW
XmNtgIxBcWPMdg1HSll/an8QuHVfqRFFwaWMqtzcxFstkkgJg32WAqZEjrbdK2QJ
m/eTwTRBgnT0N6u0t3JpyPu12FDxYt0LCUR/iJ34JXQ19JFqi86fz0zle99eYxTU
YCAs8RKCi8E4VAv2R+Zg2fJUeohpa+49pcCUxglEA61xfJbuonrO+er582PYNPiV
uEu1wsVk1tdBw8TFLNWCLAKB7MW/MB1mXd1WHGbb9bN2Ln63hmy6EjVcKpoBvrVK
5jAlvCceP011Kx3Egjn3F05DLWKGh91Yim70xGjUVWFa3mrDIGXUCLE6lC5924KS
8iOqF22eHiApy0hcB3KuBA5t3m4LDUnRGfdyZF5kxQMAFiMJHu8Ua2SkGRSU0YNJ
8iNaY7neeJ2aEo7kP76coRSfVwyQg35ir2QcqM2C36E8UxtdNtQv0P/wF3lPe1If
SA/aKkMLJ9ftKpgSE0RU4aU3pV3GmwfjQHT2cZ2E39YYqemQjTKBRKTSuNSdMayo
ONg6x2i0/ZU/s7WMEAH+hHfBR4jWHjWMheH6O3KsshDW0tyaEO4bBMNII7JeV/HI
oQwav3MTG5T+FSOkMqpN778bfTpls9elwYITzwbtF6nvQZKeaT7RXc8QYLKMdRmj
Hh4SIx0C0q7Y39clYQm3qgqmWwWldaGO5Sk7dJ8R/laG+OlaADvceNg3BEmh6S4q
zi4XQDE3JiB2FA0mfLQH/ECYYPgQ3nowe+YOTpc8PvVkCAYDW1JhTq5kaIP4qIql
2P9THHrZx4qz9vRWJETC8vpRiP90MhxyOVaHt/BulMvaLtsZA4Q7c7u+yfHY5fSy
d5jw6cdP6sKXE0BjFSCWob2CzAltf2HeYGdoKmaJv6eTQyl8htvfubXUijohLB/W
53rAemnbN4Q4GQWwmgeGggLehRhwvHwTMXQv0B0hhjawIkMxapIsS7qK9L+reU6v
or+3aLnD47i+a5J38x42RSC2tT3xNudexa87Y1PqFa/mFq8kPSy6ybd0Vf66nCeb
qWdg1w1iWjlOxMx1FmUeAjz3yQnZZY8Scg1ufg4Q8JLxaOnST/Ly98QWC6+UHqxL
ztyZ8DhQPc2YK9Jf+/z0pJnflrP+XAojvyMD3v2dbAnlLQ5ENgVYCddhS/kuprDw
R+uucz59ZdKgn9/DEA8FdSKTAATKPFk5vlABU/YUCm1kiEP9ouW7Aor0bO4yCf5s
jpC6alwcDUPS4Xj45n94TReKa4mDVPxSByJgw5FNTOBffh7pbOrgLpTWngUUgyBl
9QFlixMjEs8OyPRwBUCStDGwEJRE8QFkMznkLPCaB7sDn4ipSb3OMLvdrX3OvvqN
0EN0NtFjU2FhTT86sPLkh7MLbqxRBpkcWgorWJCLjGPNYDxVJs3iLkLgJDVg8Ya+
p7UP361tc+Zx0ypQHS+0TL1vcZ6WRx+kpif0w0hyzuPVdGxrmfHwQVyvzB+H/uxU
VKf4r+DCHi4n6Lok6uu7dB9A0DQWVJa5pjDzHTmL/8KHqnwEiOgY5MjcXpph1dkK
OcqBNdlw3pPIlBgqNGHu0Ot8U6/wS1jOcIWxikl/X1jricqb/4byrdrC7JnpdIwW
mWGaclGMwl2RHk8iS7bPyeb4lwW3/WEXYV2/nmEdVukwtQxGWCqPTIt9OvPfnbs7
RtbMjCUzZrwUqVoAn3SQeV/23z9IB+6J0yIIsx4e+GvJMdF/mvESKPUiTpRCAbZ+
Q3ROAobzzmyFMXOb7bRy/HrsbQtnEVUh+mWkbHA34WKfiD/ovNbYVZt3yzKC1A3K
deKdAu9k0f4miVtDWD5ReVNj5nvBCSGMCpMbfXQ7+7WnxKAzKgWr6etCAyUM1pkr
5mpBvK8RnFfr9yHf7afQZ7rXCXQ+2O4iytAMf/TDckLYzgKg4i2ISPKW5ivwOLhE
70adx0Rnavm3bWersDWLBKag3AfgTWP1X18pWvrcDcp62Z/wFD7TjAZKCIspcFcR
XIifU41f5CqlItmp30D3K5IzbmZeHz73IsfuU4tOmlcuLK+kqHE01e+/Kf2vWG07
mW7qeWrO8YFWbJ7/Snjq2q4YOxFie83Ww3Ep5CnQhX/4+/WK1Skq7C+DpPGtMMFe
ovVr9eFiAEibvmKU9hZDdrml4Am1kRFWHwpy+f5NOpR/gMSOPPMohAv9V38LeWH8
yPOX0T2uwsSEfALEqtsnh0cP/i5WPOt8kFtMaLZHXYkGwGOkGHuVXbqAoexvsa7Y
bkEGq8WCyutHrq0iiZLZLiff3lRLkw0V+rnOkuEsGzYvulV/p0xZabcJ4WSymbnj
GLQutRDxDJCDqaXMNPZTnmGpWHzNC2jvvHOe/XUEajWvXPbzu5b/CdRkmignq2UG
J/9c33+nObmc0WpGKh7jZZK324r3NqIyrQrXInyqHeLfyGaNCxHWF5l5QdLVkiNY
A3eC9YPVMtTeNScxQ4pB729TvKFRjehy8DFmW3LxLji+S6EQjIscMYGtcur3PR6U
epRbP+RM+ILEdBiDA9bCBzThROcxyGtiMyOmwAINZ6KKHJXA3+EPcdXkMYrFT+k/
0ARD7n4CmDMnezoSXGsFbTYB+XSlh9rBp8Xs8LfT+LRxpIIZlnkSDdQkErp/yT3K
ixQxhZw3oXLA8whRx7xwEGPeX+FTOyGTx67u0IJTGJfONfQOj+Xr0W1ZmVm+8Zog
XnfL4Kd6cIRaO4ouOH7N5dnQ3ovXgm9b0ekKsio7xvDOo2388TqBEtM0pFCrG+8w
Mr3JMOkmDsTS5KwirCRIJ0iBTU8nERQ7LVlbQjHkuboOBlF9F6NY1csKZzChHjKg
/4Acp8LNqlY22ysU5jT/xvCbpnRBu2FrofIhJxwf7dzM5y3EW7iyICsJ+Q3+jbXM
xfcVZBphFGJkPpowpEQ6DMOz5qZSMSbY2lmc5QJ5Ru6+x8X1SItnOq9lPIaPOkjT
jfwshg9QMKjbXcQC3BDSA9AsTyEA3G9FY0Fn+at3cFaaMkgM6Ai93fxNjv97I9IW
/TSEBO/tOysDYhtuiHGYh0nnL54kF0i8XeCC1ArHQdMQwwZG3f2o9m7gRqStqUbC
guM0bSvezri1XALmDejilhC8JrzKdii53SjvpNfEM78KTRjkgLJTCJ2eBj0gAmlU
qL4Oo/zhr12xkdwsQzycYRVzwEmbMY8RZA74Cks9GRgiGSMTHO1rOL61ytDKZ9uj
ttWCVG+19EOJy5tuHmXNNSsJN2/BQtHCg+GncIDvm0L9O+CmOH8MGNOwHzy2IrQV
H+kC/UMav+yXf/csDfHTQp4HksC4wIHKOW4IDs0dIVQacq5ocCKoRIfiRZEXkZ9R
aKkANSkm4aPqVo70V97mOSwcV0J3Lyrk2DYU0KbDQWuVI9XVFrpYEIohZrscEl/u
snAbxq2Hp5jOOth2tpGTfmJVKRj4DOwPLKKjp2OyD8i31yuQL/tpmmY/3Ir3Vmsf
WACEnT0E6bw+FAIwxEjamakUsz2E46w4M17NHmJ7TxJmnzKnBuYmiy5dp0j+j+1C
vnyfyQIOKpL+WYCbyOovDN25ywDpJ1RLjulhfAYhNyLa08i2Mh9UBRMurQOve/fg
gwyQGqUMnuB+D+ybBq67frYBEl8jrlCZqvIn1+cwJzqLIcOhctopVkMkOZC0gTzI
MvzjiM5pZgGgcvocTQwrUFw9KmKQSNt8OK4wNM7TkkjfQZhd4vZMqszFRqDM9tEv
h3RosKdUM50j4sDWpXUevQ4wqDYB6DqxtxX3lJOn4ZLHp7SiJig7t/ujcmqXBur/
Ex5L47rXXM7Jbhk84l4hxlaXhfcHB33WLsg1DawZACpb/RVu7EG5qFoWPnwu6hzb
rLhYBXPQyxTOO0oMRjKe/NF62GEaQLXm3vYNIdnZR89SXtJ6xysyR0GU0RD4K02+
nRAAnbmfYfSIhzV4LRVjvEmvBIyxIEFXPwkfutnU46iAVl+MqpPxzaGY8+MEbKxT
CkK0V6AgbhfFonDgJaEbeqz5SZYRZBNF7i9Clr3kyie7Brxhdvc9r1RtreO9HS3g
sctdyw6gZ2iRnBVyHwHXqBejekAw4BQljDZqQZu6dMRWj9ggXDMLZnXP2B8Kz6XD
4ydqPE+4pdClLfmS97Jyni1FG+0gBbouSag8vPi521FPFAwx2I+dIXfQItnHYDii
DiT6gOMGAMQ5K7aQmz767R5yjQH7pSQ/cegVm5ydxk6vXqUFrRREyH8JzfXgw5cr
DGTsxvqaoBsS2aO+6XIcDlLmXpJvyYrDk2jAUEkztJDdijDxE7RXSL+kGajy8Qnv
Y8dPiUo+Ftg3DrPNVQAkjiHN9MgszIPfmIr3hPBfWW1N4daAOhKQjJU16GEGvhWv
obK7hfAopY8+w9PAWRXlFUN7NaRoDM16I2zpgcN+1T/SD0LbxlhdVjJlu6GK02I4
AikIRx2TauA0UUhKQCaGiOBkMxrS2J4Wh7CcWK+xNrjF74olezlIb4uw3mQ74BTE
T0fny4Wj37gLLFlBU9gisRNkSyXEqPu9UiLaZo+QxKIRh2s3cd16hxETSX1dxZyA
WOO9Bk4BdRlr5/Dt+FU9RAl8tGm+KLxEuUhtWA1Sfah+jNZTHu01/GvY7PjwGKWp
4ELiZlodz2N4N0UThHVRKXhoLlQ/Kxxc8C4OWH5onrfpiFJMXRd6ItiggNbd2eCk
LLVM0e56tyfYbOf+TbFIniaVDE1o/0EdlWrmtvVl+akAyDQCFJzi3yCinwO38flY
Kuj+aDiRNCR3tpXx5v/b+GZcQKTG3wFkIjR9K1QoqRrIZ85Fo3JevVJVF3Llncme
K0oIiWcBNybQyt0yf5iIbUwdBMdx+AMof7Ta8yg8B6KGndugEJ2lBA/T09N2hJva
a/DML6QBAdB1v27MbM9ADJZGNiXaapSSh81u0jDmhxgEk6w9orMpxW7hruO37UDA
1IeEmDiH9ZFKvjk9TuVutXqYYUy0+uymTDKtYaScQxer7nHNzB2im3beFBbt2MLu
W3LlH0wntmbTp+x/soX8hf1Vqe2sQLA7vEfFBcR7tR6MjKfWgQhEqAdSzPWl7Q7T
iLjOqTs5HZ516iMk4n6IlxX8rkvXpc7rFPRL3HOm4vY/24CywRoYFbfBctYGEU9V
MgdQEQS675CewemymSpTb+RUHiHkvZ7US9fQbmkNSTkS8QGeSB8TvD7D+m6Q8QBg
LC8QPOCELgiuP4iCNHb5WA9KJ6Uarxb7cPMSC07IPAivu/nWiTGGATi3gn2OnVeV
xxSEIQAyBwSPdGGdwLetlD+18LdF4eBtVoAzBMJY3/jhtaV4zAlB0uxqOLj3vrSX
ej/RSmVRsjBF5N7JHMgoX1W4rGQKISlJDXbi+Eg+1ywJY7GghibLWPm4k8Gm2qxO
VHtsJnM9/zuaDizFNUTY6C0+Khfi0Nl9jle30bIu5bq9/nA5Cjjbkn72/uBvxiz2
BQquWcXQc+1DNDt67t/TF6VebhxWedVzPdchA9NUGUphAQBdMQ7E5X49x/0uWRok
jmHUY0tUXE3Mc94RbldTPYhIQbuYOMCweJkxK6AkNUIw4dE42n3RhkWPdOJDRgYq
aFUspxeT7iE894wwKQkSX5hyskJQOVNsQZHFKAUmMA9HUW373heTlqJxgTmKTOmo
Jm17afT3MxmWZp8B/W6CDol/D59qUgMYtvtr0XP7Xnwpj4sv2XSnR0NCnvmybfaV
1WGLmlEQ9sZxTSJmghVxrUbiU/gv4ifSp7G9E4g5DccigUsge4Z6MOBD2mhh9p7y
d/uwUZhRO/pu2eRvX3qcK3VGY+4TBCppGv/Bbq3+cX96eWcCwt8VFABfsNMX/IPf
A2oMf2s5YptIHugttBb/8HGGmYDZ90mQecrf4WaD2xwI4LXNc/6k6JfX8byusuhF
S90bXcdu1pF8poNomUa1eEMmnH5nXGDd7iJMQ1g9r+e1776RqddAbZRpmySVRnUJ
NtfTOhV8bgwVdw0Vjwz0VVK4QAMqSCoirKN/kuTnw+xU+GHbswYy0iPk+qS/mQ/S
3MRYz91lg5RXMtHAuwQiwpC2GgvgHMiM3QAfylJZXGVzXRFL9VlyPL1+gzAMifU8
oq6TuM2O2M6/ZwQHpBYsSM/RdeYiFm904alFnpPg8gVpgqyERKQuXxbJMVenH9oP
oyORXw6OLe7CANkpBL8hsN9aRalAsIVdklUgoUKxSOH+uwtzxzNAzJTUa8JT2Phj
LRsUkorGg44aAsm7BC2rwQubmEc7Ts0Kkhyj64kJQyk1r6ZpJlo7P3xaRkTMVuPa
WS1sRUClkN41TUYPtu85O5VTG3ZsXH2BW7dSuRZlDTHJbCV5jucQPkJ1bEjSE6mL
4gQJ2LlQZWLDFmyt9x0nXBI5RuWeRj9SwFz0lWxfxKK8aATw6muUiJjGSc/OjJrG
lyvvwYUDQP09auqZk7M3e/b8Z022Jq4Tf95LH9YXHAXhD8u5YwmY32r1uFdpeVRl
MixoeX8MPc1HJu9c0olv051GvaimbCYhimIqfneJX2I0lVICduBXB+6nKjfqlL2u
8yf0FIHm0AgmTNuvbm+SvxJZG71sawbCKtEV/91zYCwZobxprnXqAnlTOMsTmpK3
wgvFkFgd8K8+4obm5p6bmnLB3x38Bt41U73pPutLSjxe5/NPAcJnzl7PklySm9Yx
b/3soTdPXP8MMOkGg5XUWbBrIkH5Sifr/nIhXSU8WHUpBA5YU92g3haDOnTKpk4Y
UQxjXT9zhDwkdAVwao7yo+eFLpFG3jmuUVXIuZXt8gekNHjBUBb7T4oICm/Rl+FP
qqfgxt6cuzz+4N2Bz0gspTqLwklA8LWXMpuy1bR39ecbBh5trM0rxr0O3ezYAfRZ
0aFIIjJG94SKnbctsQRqjW0vBQp7bolaRsyuyo8m7sLahZmIImQxy4lgR2WsqNay
/b9w0u5C3TM6LQgEInLZ5wEucVrfq3AYw7NoWpDVWE1v3VjB/bHdUDhlGUzslJXj
hAmGoPF9BBkKD2qG+mCg8wddV7G/ftO7Z/FD8d4/anvEQZUX1ShSw6TnDJUlgLTQ
yATS2xffuZ+IiZxq2CRZO3YsgwejB4GJdKfGBJIqGIkFqFC6HbIq+6RMjxK4TnMK
Tl0SZRyqFgLujZupAg1VPR7QtJyNmf9NvJaVxfBsqZJf6BcH4bPp2chqwDsQc7f3
eNnN8Mwx2OQWQlN29KaCYrJAnkx7MYZHuTh5fi9BDpzR+mVfG3hKvxnoQJw7ds3T
oPTQHEf5sSVUBNZOkOVsMA2qaYmkhpp23mcej3/U96xUNyERuuZz7hoDOn7UKWqs
byUPWYaRMpKuQgmVL6NvTfl6+tw0iHIjyLUCD/U166KB5Zx2Vu35HyFdyBC5B5OE
BlqvIXah5GbQyk2+pc7Lzj0uxrmq/LfyGa/zkCVcUAQRVLjFqUJpKJZaNqhkrePK
AQpAOorzym3pCmc2G+sV8V9Km+TFRye+NgggUQJkAHC/0xfPv1RCb4+HPVPR+167
vjVJBhp+cc9PI2V1wqK+jg/irEjWBfOXZmj7GRhytV8ZIEAjoIRji4TZ8r7sR1GB
JrnF4illSnclo1V6lQTEaOLD6aWOdJ9ZCt/nLWKwsG2A62MX1aP37gTCRyKgyaD8
SqlRZHqnTT4bOIQcIonW5hiHVggeRuOwHH5CV9uE2Vb70qo7ELfz5ITY6L+0XnYH
wlZvDGws0FrVLU1beDEm7pBgQ4b5pDcPghiTvTJdsRUBsEvZHAWYvNNTWwuqFKOw
xFl3CWVgjcymu3zIg/JhjvnpV5qfG2T+U5hYhQFCdRWXNC7SrpDdOssvTQHVMmEt
YRIBNap9S1WfLWyyotkX4sPI4VWzTppINSN1IZ6bTcxgu8+J9ul6F0JQjMwLhQpV
UHyKZEKWmpVk73X+oxK/pqJTS4iROKqTLc2Mft0wEG4hmUaq1e0oQ9ncj5hH1CCF
h5yYhd8wFyNDNxkKE1r/f5t+Bv6iEMoccWY2SAJRMA8juvVBh7vkxcl3w9hMi9Z/
ptJN8HvOLuoUpTJ4wgJVJ4jWwWqEdHGCXjoSjXVh80R0ddU5dGSl1OrXyFUBnqce
InwAG3yyqIuuoJr6ikqke3MJM8y/UGFEYtRuHaZSyVqnkLOPSpyzDHVdQBBPH9yK
UytOoJD23okLI5cMEPJRghtNP/v3JQJ4ujEkk+GfkZaqeolz4YWniNMq9/9RW3c8
yHyPcE1AIrehJUvXycpPLZlQUrXss/JO9Fnrd8ptV5FVKR4WidN3xML+GpGHKsiX
pPHsUS5jy35CmLwH4BqRsA1q6BBjdYdDnSbtdo/Vq0hVEKgcpJe1p9ecns4J5XXl
2wg2HuMTRCihWtC1XOTaqgiCpoabzJG2jJW62QhpKpijYUhMmygHWADSKygi6q9g
gDEvNJiV/jLRC9Rvifmzd3PebuZm1QkXzFrTv6R/6ZbnaN19X+yAw3Aif4lJlsXR
H6sXtLFJmqzpAAhLtUHd9Z6va1CxFLXzyrKBc6MB1cnEE1RADQXxsKpkpoqwm7T9
hFSZcKxYli/YoDWS4vllUCoJrKydQPYB5ZhU0OwgzoJ79u9/gSPkkavIl3ikqmdE
ZFE4de5yx1r7CY9fUmeNkgyHeqp01Q8B1uZeXt3NLLyy4FQFVnR3D2fpI3gkWvgG
LsgZp8rGotkIBFRi7lC6EdVygvMVTYmvcggldNGdiszn44nDxPdPI61F0y5/dBwR
kzq1XUns8/79DghXP9GYWZhjxR11oW2rnGwEKgUp4OChgR3J29enFB8iLjbPIiLy
JEm+1Kw0GzWMJOZ7pIY0sqJHzvWyxOWCjSjyduDsH/uM23xGFLO/HwSZ919QI/Gu
UR4QgnsAN9bzhugq9SV/uMdTby7FiRSxtF64O7ikpzd/ZI3+GoUEU5bhT0imDhB+
Iafoxt2BIpSF8hji6YyIlCmplz3AGAEv9jvJ8vMpnHtaWqE6VAlTuQsWTBI0Bfzt
lWJrHKY5to+BQFT4o5uu0qgwGeariulCCSi/px42MHS7qyOhBhRptkQojWThZjE2
BM2qzyFMdfXOGF73XmqTapxq6wqX16bOxH48xy7UpFQFTQedoZGrFWPVANr+yGtB
KIQm0McdiiBwdkVQ14auDtljR/gc43tTLvXJaBPz7V4/NxOPW27KqrhbaZMFOW/8
HoTe62Uy5yVdE6GyMyF1obB9jXexeoQnLoosmKgREfzwS9DUciXz9VjaQYJU48F/
u2knOg7IZQmq4vyUb6uLEuLH9Arrv1R/WNCfsWgdWvWfCMzIq4SW3zHLhhrXwCGt
8zT2znigrg5VPl+HOuAIM6n3/EknFw31lbtqTr1JQaL+5uxtxw+4gqbK74r5/m9P
M520ynQAwDXSoyQxB/NCr/+vO+UcjPKgY8taPTciRXOLX9cKTsauTOwo/hYjpDRz
RySZmfnbQqDF7xKbNw1pcXotj33LXdjLxvgixKL5Exots3/GxyOgtvjs0zKr3UCq
w24NvnlcbfuqR8kxnesTOPiz3NBAZQlSMUEvRMsI2tdVfvOnMfkxu1RvaU45dByQ
O4vZJVdTnmmvEqkd4V5DCZKHa539szhvHvotQw0cZuKyZRkOER5J3ArbGSEw7w10
pPszoKOcmUnpFOVUMHSpsfG8JCKGlsFfKYo8LPZuPNmeFh1V2rBlu5G7qN2vl90p
CJ+00hPo/aDy4lnrQ0aydPxcAIPQlFSFXF5HnQANllkKAjldnWH4Yp3+ofRA+OpA
g7eK+ohxNs7IAJf3TH0lnA6Q+ZAonmuaQzM6P6O1rzzxXJa4gd8ts20e1Sc8iXdm
PM3mtbGnOoP1sYyGyIHiCQbst1aE0U3D68SVABciscVUok/p8ZxeCvOF+2PeK/1c
wr0y8wip7MtuOaQqtjq+fsO/fe5F6Tx2THOOsk/r5OoGnyeuU7eyZUtFeHXKiLdY
0cKVFOVgDeDkm2RgOjOQ0GGpYCCzGWRd71K2TuhBgtu6VF5uqS+I5AXhTxhs6fqd
aU2nRxiWN4pSZohMveiLbhQfMtospegUBtuIYvtAo8sxrLvIfK/XiZp/AiMCtdem
GGbaecz3N/ShHptqD0B0u4tDunW36wLmLJGo1uzCfX5wZra0GXar41COOsg1x1Vo
QYzkrCIdOtKOCMABCmsBGdeOapUX954bvOrVCqy6xwJ4ljsCS272ibkLaj/55olP
35LRfAKpTW1vF5mbU5Z3EJtdjRT5kVi+xWYAVplW8uCg4uO5BqSjanExX9T+7Yvo
8IUM7c4zm5TgxK88EZlwGlcQ4HI4+TtGufcCttS8JRAHNRBPO2uW/oC2ZoI346h3
JZ/AtNACwSiq847ZFPS3ci1ghd+CR46GkUwTuTsSkLw6HYNiliiNl7fdvzLNljoc
jmsdhVBpQOg0tsRcVCodPGveogKj7R31xcJt2XW7hJrqXunB4YTi8s8zjnG89E1d
XVE10xT8PX9/l3GHa5lVgumDWLyeSV0H3DacFdOPAHcCE2GUsPWi1i9qN01s6+68
qIMC6GWQ+CAts4yxZyk8Ok7Rw2Tv60HHSR7COwIUeWHJFtqWyRYHv9pEd2uLSnLq
IJQ0MkoPr/ucWPknLi+WlX/R/mLgE5xpt7TWXGoH7neVsECbFZ9qcXImnvNWXGtK
F9zOxUuZRLBuAA8TJtSkklEA8XG+i2IsLbK5u1G7qJz1i7MEKrWJCAs/JOGDf5ol
jtU1N1fOxmzbdhkBDA7SxD4YAPQKV2GMZGoKVoKgv2UvIRFWZ5Fedp85SYmwRso1
UFlzi4eaAPghCxgbE8TnOTh8oKp+7VJewxSZLhb0+TjSaUkoxjC5f6tslrDrjfL2
gNOD1k7T+9+H6CWHrIx7ouAY+3DD2T71dIh6BnFVxypBwHg5xUz/7XJZl7iws8my
YQO9ONQ7rNP47fPZTwLBLgORAUyliLkHxuiTUK9O5a/oY5xCuZ94LkjkB2FmYIpM
VGWfbLNCu+gnHeXigubB8Y2V+d0emEA9P62b/6uYX1M1Q9b3xCyLCJaay1o3SpE6
bpwrNTpV9SWxDKaRhRV1HXXo4etBcb8eVMDcums5Dg5/Yci+KJw+9nnPgXXwe4yV
LP5CWtwbZL0JhTbKwIjiC++aBK4lpF9ILVo8fDl68ZkxAo7RoNYj3IC2KfCipgO3
mXIb78bI6KFRyqL82F73dnXP9hxJLiwhN0mli8L34Z7AI/i1fL41zq7/khpvVm7N
PGd2Lbfj4na8gStLBeCRe+9PSFPLtV5rinwVWzXcpYt5r+vOZwfK+MddgKQBR2Fq
eSpP1rlM+yNG3NIPPUKQ6KrgryiToIQ+0s+DWzYqCOVFeSqwYHMoHmX4dyjgwGI9
Iyf8uDLU9v5gzvwvMBGs9NWfbwRDm56ltgFPwGXNBj09vLUPzyp1idSxNCcB7MVj
u7+uM7SpqIq85IItAq7CMM4+qlEh2eW49ONDPC2C5MRfA+hJodxswaBcVkzR5fim
olrormhnDqWO9iNOjEr/n5qI7V8ZzznjLD5r1mnQiOl5Z9eFQ6lvbyrDBiHAu/YV
cY9Fq5Kcogf4iTJboO0/zkyve+VhYYhGQuoYDLWSOG7eCPKwdxJzRGxU4R9Q15AQ
7oTzq1KGmuIwE7Sqz2oyeIzITB3Mycpex68FETxhkzOowqVFI+eJg8Z7iTJrL+Mo
BWZVEExjCZsW63U5yea8lIyNDoMdO3Q00IJdTcwAnpauv6HMgbIN9BcBXdKTtVsT
snK1lsXOXDzaUkHOYw3VB+IXImy1jzz+9wDzKE+o5r/dIghHKWBUnvOUmvBmEeXM
+cP6raSBtHZLpugZVfPe+BJc29iSS9pDW7E/gGKS+o2SYQJInV39jOxuQvIM/iqQ
+7GI6d+X/B4vrE915mroQzSHehGzk4lN+IhyWCgVx0OVbp7euX9FnUqozAmbR9ta
tQG3tcy20UUfQguFbYJhNc4upRKPUdNdL5oimGUYzbxZxj2sp78DXlAuiQXovKZY
YaupcRQw7XLt9VPZRd4JJS9QRlDDscZaZVmWvWuV8JL4Jx15nUKboFkMo5GPGS4P
VbjECTJVdu9ED8+9MfXQPcgLWxl0QvzDmgK6sPc4f8/csToBws3IpQLcitplpqg5
S7jlfiQQei1yL9vlPmY+CEu+ENc72NQNZopHnWUDqmRxjVJrY98yHsuXFaYmxB36
Qu91JxTJWh6paRTovUtrO0ue9w4Nx38GoTlHYloKCKO0OTztHI1UioR7Jz1ed6U9
8bHHruBOCczC+7shL3pJMSjEtOUy+Q2PK/jLAtTLPy7Glqr/Axf/FiTge4GY8n5I
zn41FYbm496d8PJJYt6FFysZQa1xIKhZYeGtV2LZd7HiIVw+BJ/VxnFlggSYLzQH
k/M0+7swHZF5JmW8tpELjeyCteGA8gmjgizdLXB9V1D0pXrf4tEhVyio6Ts0CFCD
4GEn/RA1ySQjwRehlWVdZDce0L7Z41Xu+mbyrgcSMSrdzqFlV0+2PWr37iFgGpD+
MPAefQj1OQWN+yhvo0GEIsBaCjd9pkdzykx+HTWjyqKfEiVQFmQPKYBXx3jPpJuN
bnbl5behBRYTmuxi2P7Lk1e5EJUcNqxocsXzA+s93g59AsWLRpkrU97Bgyjvp+Ab
oKWLT1EHbXD6S7Mph7JmZhiTYEJvxiEE4q2mxQIAukGMb7dvL2Ltb8gUcF26yHx8
DniLlhxpqH+/eq/0GMi4jN1V0AOB1ZSzgm/2JQrYateYSSMnVkOzwGnHbwzImVr6
PrL1KU89oUTOlItVWgI5pAmjmADEFaF+YHWLGNN3e/TwUp6HPT4ZwPNPodC6Am5J
R9/+VElWHEUZ/R+2E5o81nKLuJPVET5JqF510foN+Wy/PuaP3o9NpV9M//m81kPl
GJJxz+XvY4zEuNzRx/b07NXPdCql5HhmgDHgG1fRISeIeiC2HjMwuZSaAXgXxl+v
DCFhIYDMXm+obypughoFT8i0XGPH+oNLn7VQs9bpLfjDeHH074UMenrljh1z7sR6
Htqn9IesEuie2spPed/4aVAHFHHgmKDw9J7DNdVl99bubt/YrefUENDOcGivrS0j
B6w+HcgLpod3b0QWvsf+GkOnILiKl4jl6mWgsTIIfCCzvkgQ7WKaMGZj3+kCfFFG
LnyfjYkvtE5Udx+Sls/0BRCp+kD9FqGMXqZs6lmn2dYruC8vEjXkwPqM+VuRvJin
/23W5zb8Bot4TXysoCo1gRy+SVJt+3oG8u0ERBiGXvDBc7GnnXGr/kpQtGk/Yajh
fXA1X19b+Wre0KUemZqou7HcA7tspjBitXh3boKCwqV2AAb6B6u2P0vdaiSxqybm
JmymeI8EFTjuBhf0AsAcayghfD+iNsg/pB77Su2am4+egmkrXPgc6h0E3NO3xE+S
O+LBCqHtMJ3W+35/taPtXdK05q3nqA/UzJEFhO6l0n7G7IFjydsI4t2O4kuQW+aR
1g0GZJig7wIgDSJ7PQSUdT4MIh0CSkgE5hEgGwnoUP7bLkcJlbkjfvLaeqjn7hiY
2QiU1r+UvXJfKBLi9v9Kv2HWgFNH08EWMzg2Vc9hlbz3awS6sNeH2ejHMwP9ymME
i3DgXqiA8w8OhX/ytrvAzuv0GM3rA+Fc1m1/OM8He3LO3yDJZkqa6XdUfjzBQ9cq
+F+MkSgWgcIqNQiH35mwpm6NFvLJPMViK82gu0bSMJl8szbHZES/ZRMf3PqHQXE3
Bb38DnGbOyYe0dXlHL+4ZgLvt3HGnTvRpesied+M6mmv70dTbWg18LUJsmDshpsC
+xsHkXEoAsdBs+dI95rPG3FvGzswTyJlFjccupHUBKv5xxL1NGTXaMNgSqhc73/I
raKAKL1DHxhR5Om44/R1APse8L2aog+OsQse9FoLGMJNXpej0E/YjbF1IugnCP9S
hMeVmefdc9OGpicyznCaDAabm8KKcoxFgvgi/jBdGYcRo1XO5m3F+Too6f2hHKZ6
Ggq1TsyuGtMd5N9S1Qzr47pUOy26HH0lLTzOhYA+72X/SUEob1NfojxhHxIhQ1Hz
utBCxmDVT6YXm/hQyBAnbEOya+qfN5DFpPJa3Q4r7EyvIQNDadbUnhkEln8kDvVl
NJk6PEg12+NcftlcwLVGFU63/1IGZZM/E6JQZvqIebijjwaqo+GU8JE9r1Lm47r5
SnzDO+GWnScvUKgCwMCX5MC8+Y07h+BMHp3GE8wuNTmi0odsgAME6xzubVcdZXCO
hHFrJsHj0gX+MiayaVxqZsQOGWJP0+ejaOnLtRNEkNQofWgUit0we1DFTI8KTaw5
7rP/wC5HeRjcpJpck5wJdMoPdCVlRaYTDH91Muh2iwvMCszYHNm6wJIoJRojbVjB
bWd3b/1hOwCxdm+EHxn6xq+IoLPzRABknErgP1PD+s3Sh2+bAHufDkyQG4tibGQI
A6kJxARAd1KujGGxZiAtDnN75Q2tYOsCOOdtwcN42Sy6YA0PjNRUalos20IRpGfi
TUAYSiycHKt2UySMYh6D3tTMxaaWn3VslPga9BupGfHZsnorMWHgXJEAzb/FdMiv
eypv6fFj2934399t29VhY8elbZZm5tIMSZlFPfDDcCUvM96Osybha9OMGYpqtI9W
+/bMuxM9wcw2bV3s/6r1XZBYluNFVfro4HVYDvZghSzJNMq5qUsyROIWNywB/CKU
OD1PAo6bB5CVRcju4ui4d3WMBCh3Rp1NS657NsPbiNS8ceqYfR4G10hhJDKbMNky
fOYPweGY7NZ5IwedleHHM2O48BWSgQjkncwBl8VXFf50DHLRFOxzJufwZOkhTJvd
eyOZoDtCzavBWW8ikLBJWgO3kk1mGzSWj4qXm5HTjx+y4Iy+HBwUVn9Ui7QaLxZp
rjCEH4T2FGX6O6oPlQaDXo9/8ObpeLzrW6JjufYTx14rdwYXa+8Xqn2cM0V+JeFA
+NBs+YNW/BgOGUiUICG1rrPOTnrbsVlmCh1BCozcwgN5FZ802DC7R7dnRd9F9lTu
0GcRm5ls+7Wxjsv1H+NuIxORBivdCivZ6nHdS22syaQcqsQnsMeM4k7Q1Ob75R6X
ahRZJ8kGMXa43mzHQIUbcsd+/Hfwg7alBjO/uh+l1z1tVp+32G3D7M4vp3UEGtDa
0IvvZ2S5ao8DhfS4nxWK/eAVJ4gVQcouH404wEB8SoJvtN4ZHcuo4P03jt6VuWFO
Qtum7P/k6Gvsm959J4ExEO5284dWcjLKBpNYvXE4FL0oZr38Bki9Cy3h069eg0YD
/p7yPekS8hRmpnAiJb0wn1v4BehEzyoyRsoYvmC2QKjJ8UpTAx0ci8IsVsZj1x48
S2h9rPMREd7UA56PU2a0o27Jv+YEi/mBcDKCMKI/4lCwe6nLY4zlnSn0t7IUxG/l
J92nJo/ifdzPaJzy3M4iHIsPwy4q/9gwVAkIe5lhFHWTgsNGpUNTnWfy2FdfuiAL
atTS0hCAaP1Ljwyr9Lt4HpaPFkIrJDvb5NX6aOvA5prAaNAacYenryPAjL+weAyn
NI3QevC2YCshvRT/E5EPC8UOVHhY3aIv4M1VBkFoy+4G4m9tcBX156j5sMiC5NdT
hxmwKqkaSrHJTKM8MLcdIc4DrDc3YK0udxN8oN4FJip8ptScEwXzLz+adauLGa+N
WKHUAf5jKdNEkEOvP1uHy49FcNSU7jtS0NE7WrduKRWus95XX0WYpcBF4BmqkUyA
DjObwvp4xBbJv/wG8/YBkyPsWQHb22zl4dhnBv61cc6EMmxuXZMKjT1QHY2aX3zp
7MBQGjEFoKL7buTHJrBA8ZIlfD19TFV4NQJob7cLY/GGRiPFPyZsZdv9802HSEpC
e33MEYGwZMhN8OvAti7lZiAIhdn0JeLp0+qxtektTACxuW+hyttlSkSu4t6TLdyP
l8n78Tg7jaIJnsb2TF9AXnmkGW2GRPm3E5i0ik5HbyqzYTkUwuPnUxEtldmPJVvw
AvGxHfoFnNZWuqOWIi/Lky9nu+nYOdT5R9+Hw3znLhAqxhuix+CVhHskexLkTo9v
mCqFZr5OeI9KDu+tblMinoD9/dobZgnT5cmLFigalkWVBVIYbMYZHEEnnd8wN0gg
H8vVxrV8SXK4sarko+bJmyemWNrBvKjRbQUTOwAJhvtzFwFf5q7d+G47SEmaZ+Lo
5znK3wt8MPLGmGUMkQx+XJ83UsHAnznjlX0xf7DJvOGqqcbRsMYvmSz0EDDjk3JS
6get9rjV0YuTatQxc7ejghHq+HFxMWPtcOGHdcVeiIdj9aQ4T7Io8/JuiKn27LyR
PtasIlejwl8CFK9Fn4BQRgmreEYSNQBnUUoWJ1w3UIEgGgIlryO1wDSDMZ0j2h3M
Q7APYigYq2K6KsQiemKHBqtBKO4UJBBk/G55tGwusQw9qA7y5WtdYpvx6et0ZTld
RgnM3zBmyKRasZGriVs2rCn6IO/NZ8RW0zrY2lm318huWXZaKnmWlu0LqjVwgIDq
/FRKHYRjDLIAa5YoG5xPKimiYuZgnW5LD666kBKS5wpfhIusaDnFAFqr3TOQEJQX
2vTPvBzkyLoLrI+XPd52R8sv/p4H/RkMc39GnH9+Zdx83/z+PjXNPD7wz4A6pXDd
cV7uBbvbyr7TF7RxSlI8Xrq6xI7CM3hiohfOGuN3+cDpP6M4/Y+f0XYE4Dyfn7zy
PZ/szmruiaan6X2Am3cMnxqL3ylnWdzfEvbobAuyAlyrbHVc+cI3WpMDA1N+EuP8
MBx5w1moFqSPrMD7EnOttucbTthfRSb/hBGmjCC5xNnKBx8AWPjZ+UHkKsYQcGwj
/zvaIBeWdd6IPfQ3OdsdZuPQPUXbNQmiNBmCnmu36r/OZyK9QuFXOw2ePYmxsDjP
Zav5Wj8er4qRl7rjTEoORsvctexMzvs3tNEJ8v5PYYUSpFTSWcNZMKS5wdxzXioI
AZJPK5Sxqz3F1XH7VjqNcWL8lpkNe9ryv2bcJV/7rhbbwZ/qERR82QA/njF/Z/UE
XswvPcwmep8Cfa9ohM/YB1zYwYqUjr744DUPtxdQRyRufC6tr/sR+rLoCAxc9N3s
xxhsLJ+1prdRQh/hXNS+GiptYCOEn482IzzTM79z0rfVJCrvSjLkf/OJp673t2mM
3GtHjae+wsDcxdb6TdvI4VZwauboZbDrK+GQ93T1O1jka8qHcxOIfxJiv0Fwn29U
oLbtSL91B5Sw/esO3jZy6ueIXj37jtzsqpcMefFH0G82VAsrLBz3r/gcsIeci5/f
nGpFJlfWrtZ++zKzh3iu2ydr30XL7S3z9FnoqVoGWiNT/izq2wrgaEuAs/eBq3kY
VOHSQRAPXpzkDLYi6/hibiFad+I/9+IXlj5b81d0/pSsyBXzkkl7wpbqj+p0I069
YF3tW76VaM3FA9Kyu+WACLidRlH510koDAjbdjIGwZWuiQsPsjTKqU64Hr04Niyk
TQYGMUoZX2G/eAHeKqn4kJhn9RXBB6ctXFet7sCcs3eydqSh0UJd9xH1P/kgd6+N
nyVtHBMmxkxIDlUnzHRZPZKF/x//okvLtbPjv3sLNeA0UuKkzv+cvo5IhB9ZzxHP
7Q+lNIoXyqTgECqQfjOggto92ES8s+I8nkifbRgoKPdj1Xnd5PUebFL2CPrhvK3X
zjU+TSA2Kpl/nje9DPVBNhk95aLP6w2c6CbEJcP8LVQqQkHrcg3/uscFoPSci8F5
bLoCorOYjN1CKuEmI8BzizHAFvJs/VBvZfuuX6QRhj0TnaMvQpaYM0rE+rMRxuro
CbuHkTCXqLNC/B2M2JqS3EC7Z08JwQ+sAu5wxss1v8byTflKMGqUs/AfmB4J4M+P
6RsAethyxjyGkn3hGZr3/NE89dHp443FT8PIu88bNre6pX2P0xR+VTj1kpl+JJeZ
vQCcTj/ptTQfsdHWM35MFu4v2YLzzdcQz9HCDrAke8Q9qTIjBaOCqFflxuafAU0q
fcZ7GhBHmNJXXqDISIKMfzpElAIX5uA4US1Z2+Il6duif0YWHAau9M8NyKCm9ixP
LIvfwIVCJ3U29nLVZJNUmuNUIQ75iOEQr78tMEuTxJTfVHBtOjef+AyZOuO/lbOR
iWCNbZ6rnOsHvRTgRAdnWZPeausBv7Lgl0nOi2k0s4uIfeQmnIY80HEkzGkPno+O
DH0ijUa693aOb7XoVY4OxJbT23l2UudIl8ieSyS6/GfNKYYwZdQ9bs8eI0Qx9ZnX
8d15GKFP31tDdbSizH/NkDus5guJyOuBu9Uf+V0OI2wjxHHfjyNo4bY4hLEcPwmV
4bDaVNjNdY4qZpz0AkWXif10fkV2poktdi7PUNq6yjUA0XR8IPyJbh+LrjvMbhNx
HmkirBVAsl9/a5M9V8qPaGjxizKspaQnhG2D6vPXnP72vUqjKwE7yXGDZUbwdhim
3+XH6U0UQ0dC3Oj9XrZfmo91EupseHNAuH384jZSmmzLFhlPn2kHHBfVLOp7k1Wn
9H7LksUet/u1cKQK1iGV9siG9+p2tMHsK9MEbQHrttLuwZr7eznreHr/nEuK+Pbo
x7ENShOQBX9VJngrPuPH1UpQh28p2dOizlZgFOxoVcZsFqONQ2+HHScGYW5NJrdk
L0+IeZQXuMwRtow/S99BUunblBVtB2jpWGV+F7nz5R2fWHp/wqeCdd+XDRjw3hHW
4WTUGBcwyNMr8PwEguzHxYO0W7rADXJIZ3DYVTtlbvYfqIMxPod59AeYq+B3dSX9
Z9fjFG7TnlCCr9/6uep87nXuacXFUqGk9FfGM7tMG25l3cN/gT7AZVsmC9YQSleP
d/LA6vy8IEqbNcCqzsst1pG0DywfDmsrbjSH8VJPOzmfElGfRhWuiUHw9jbtOUSx
H4Nk8ENIZ2sb4FmlElZQeXAV+VP/YnSYGPVRZJ0nVTahIr0RSRPapivBhDSNMcuN
5It34r8/LEsoLfLEUgb+CbrCQXezbZzL4drp8gUXmGlbQzH4K56YjhnxM8NCJxK/
ASYn8/f8+KFAaknUxebmKBBrzIUFYrkT8APBo5IXadfZn/CmaoT4aTS48DRKhNPB
OdWYU775+46n555WGU6INiUGcqDaAKpkia1QjIHh6JJrDs19XcTb5yH5gP7mNoQe
h/0ViCc8n1HdgQ7nQRj2aW6H5MBRI/4VWGslZGjSv3yDBIe/VvwvG7BE1piH7g1s
2GOX05w63ubopiySzPUVQJNURfhSAHDu6RwQiRLqMe/gyLyPL6APuocJYXQPfm4q
4Ah4TYE0qCrtQhoAKzXHf+XzsMZx0qzqhVVDd91rs1HnOFEg5olx9Pq9EG1qpn17
ESJcxf05hAhJfQwTduTugFuErs/kVyGD8Hm1/40bKJUtvDxzQ7w5lXI4LumdOpRL
p9GyUcOuswx0IDWKAnVa1EbXmo6yy4JDorniIo/O17J6WNpVEppW1D8MtlULP0q+
b/eEdFpbTltZyR5/3NGLU8YkgvFUTSK3Lvv2FyzM6pqNH+SIuZ1E2TFEQ0tKw+u4
jv6h3q/cnmtfqcsJ8US7i+GjXXGUuKJ7jKYnaUtubKID8vyEjlVGMWunOJoHX9uk
zABBIT4j1ziGayu5VZNqJ5OQoGnPYnBqTsoE2t6qloCv+PLEUUAcEEV50UECWdA1
rv+XFGnqS1WtPTQkSBAiVsAYYR9401xqufjWBphD7ov9IztWZLyPQQEWtzWAZ5gL
dufiLWK+OzKfXmI21xZpJSvpUCtfSBMGNS+WvJ4BKl2lxEeKjl3Uc+31SLd/smAE
PT8zN0D+rEL8TQCd41T01KdjeMHdHFQ60Er+WK+kTLq14vdQfIyI5oUKfI5XrBrE
zC8ATelFzPR8/Jd0NsCJhOs7gBiATNdxk/PJ9oEzruuVgqzSr/kl2xHwqMW5X27E
2tsbfh8OcpnaLGUbv3cx9v3ew1eaad+J+tF+dQI+IDLzUgoLJ11JLdLy+sS1Bn6l
nizsBSzH1ffRSCMDtYfMALg3dcwZ2lBTiBLiVoZUlP3wQJbkOtfo7YODm+5KSIZt
5zwhPt1tmAu0M0ZLJIhWe65Odoc3dUL9nSRokZNGknT0zxAhUY0HhD95VSAWKMMA
sTo7VdsG2PvRRfTUxqy4X6VOf+lpHWMuS8yS+ivMbphsvbg+QbWurhhN27doYtn6
cY9rELu6iea3qh+Shqwcqz4Qwv0hDkmHzr93GvcyZu6epkvNqbzCH7P+OzsMLcoy
YjLiL/9QUDcTxFzxxZI+xFo2XPzbmu2ujj94ElsjdW6BJEa4CO5uj+g/Jys6tJkK
1goGeB5VvO7kmkRbEyvaZCqfgDVAj+aCni7xrdwF/0GBEt6gjKQdKr0G2JwjiGU9
nJZkX7x9j6clJQeTrHHA53OXO0ww/U8c6xG1/1xo6GZnkMYY3tOpK51GFvJM0Bsl
EqC/Af8iRGewPA5RxVi1X+krR/WenCHs+T+e18+/ZVLqFkT59uPKZcyNZv+fUtbe
UpvHzsOYMQZsbu++NEMMpH0MNWwL7oIWTeMYTIIDdDYGckSLg01ssL2qo46SWNCM
DoRn2nAhYupvWiG1zPBMlEGoGB9zVsHI47TntymuIxWNAI4d+50ZZszjaWYALEqx
3ez2qzRmYD02dkvoZL+iye0m2L7nsRBGmfTeGvEWZt3o+icHcDK4kvMllj66KIgP
bhzERGSeGA0RXNhK+xtBgob3/Pj1F2qn5ToburFTyy7BCn1Lv856NMT3ozveiX7s
PAWLRVKqxUesxXlAc4tqc51L89mgiNCPDt/NWVX454ABYn2YGznDSxj0MQ3anVDy
fEOYIS3SnztjB5xvqCFOwwy/upyzCgEvcfnn2gsolhUW8Ys/I/OcfY29YfOurXNz
L9GImt4X2c/ZCyWRzanfccQQNZTnNAvxjlme0cBENff4oD4aKoNQnSw0s8lmLwKu
md3FuNFsyrLNiBW6Fc6I1FTUdajZmtY45WEoxRvTeH3mnn3LG/CJmu8stxqBBe7T
SE5pgYKkhKmn11O9hH+PKhSjPt6DJpc4AmEJj46HdL+JsbDWwaQD9joqTvVT29Fd
efbsn/b2Yc1WStVii1FMIKDDqqIPI3SDEDZx8IsDLkpVWuz223oFLU9++tgq3HIS
1ZZwBgXtrbwoSBRBBj+nTGexUPZ+VCkOxXLqXMXafOMq70Kr4uTlXrb8mC4It/xh
e7BFntNbj+RojMucHKyZ6zORO3tI2Db2z2UMAm0Hpe+dF99VTPUe3bScrQ3gi0u2
ioFQd1gcPggsrV+/++3y9MEcsDNF+safgCBvlPD9VsAHPeoo9AmUQS0WhgCWTaEZ
hFz0HGRe+ZtulzhW4qlqzaA+WjWBKYbNJszADyMMWcGc4qXkjZgUqbpXZ77Poj5i
epMndCEy+Vn+6rHuhR+v+i5hdV6GFXgeJnWNvkzpqSbnfeNTynhnLVEz2Lc4nh9H
14utH9NXIolLeclSDvKhy60tXC/QrYgYbK04pPqi9ojDXTVNwnB1EY4v3pvnIXaG
iA7q7izbw7dBXnaEamLXC6YC36ss3NEgNrTrc2s/iWzqIKRasLxrbL8LU64IYw7G
Q87uGybSK/e5Yu/k6xA2uEVtU/LoF8RQwrFNan2BvJDo3UAurBiaM/yhG6Hx6KKj
YaxyuYdLSZ3RXu3Mmbjwwt4PzM66jSUoghlNElR41tRXvaSKLNAZ1vJSWmARTF/i
3Wc9E9Pej07ri0ETUMc6AySuJQrJwXLHUG8GSrhewaADvZ46tGTa+pr4hs0ex9G4
xV5k2Nm8YkaCO4Nx1WtnQPnJvD9VFFFYDEORG8Bv2h6bZiL+Y0u7vAXsupViKgTa
J9Q5gWeznQ8AS/np1zYPX/pkVVHrn0o68nsnVKxnW5vEpgMwBvPqiuKd4QDUj2yP
G27IvsP+8qt0SZ6l3mcnvqMJyFuojmJkhF88IdAN/kM0ABXfxeX5/ziKxxMoJiIo
2mL7uOhTprRMiYyj0PPLD6IZGSRsMOyYn853UjvWI3/Yq7I09WfKy4gvTmwiWMeF
DeVUXxtQ6d1K5tflnu4kWq9ko2gkiqgZe695haIurOv3spmLyovSsGvSFA45k9u1
vjSnDkuuIXQtCxjXJyFyJoMh94aWCF6XhFdMTZ3IaY4SISUBLogYeGUCWeoSH8kH
wtT2FHQN3sIhLkRRRxVOKq/ezBiDerEvHPO7RsiPqO9Shmx2Il+WYZd5ml251R6X
0LgKNoXGfYebgsjTP5K6BO8b9+qR/Ii5xLhUA90LHbtqHPN7bjA4PNhzDyjljPFA
4ibQeM54m/prfFr+UTJoSoYBqvSU3kmBUswPPHxVITHE4frytbxir6lyO9vvQxVx
z8AVptUGqy0QTL8bUjfoitU9kTFub7FqJQKMEHiPI5H2Km6sV4SCK5J8xfvB7C0F
6TgbVFLnSd1WlMo+BHsed23/1VmcbOaghGw85AMB9giUHyNi1q1HjuS0EGCWtIte
pGDUQLWpLFMIfTOl86MRLbrXTK33qWWehOaRa58xz0j5nsDhtN+NQC6/j4rVRAnW
MYY6BgYBQ0JH9hMBKXkwv2OWU5QTuBtPVSVU6UIYmTAY9Zy0TA+lV9u0uUIENRTe
vSQUqqfmO/14fB1N1pHQagfYoGnax+gitgeOPnaYGxVZlWnlJilF3FH7Tvj3T4JD
Oo6K/dCbr3FmKt2zeWmk1RCm5w2WDvEXcEzuOG0eN52OlmpFF3dyM7xfAg5ns6xQ
BrBh+m6jRPyPamg2bPsJWhzpy9KHFoA5pRZ+FlKGDaggWWLjwrTTH/vOwilYGW1Y
IAsOcwjx1W6jSLCFdO9+f9wt69vlEIzlKSWtHVObUrL69tbDbAUEp2ksXgl9etVQ
Y7Y0AP910y5E9IPS7RNoMLvNpV/BqXerwZsktjH7iMWyEKVp3gazZbQJGSujJ62z
QNT+qIBAZnInNGsyDKlOK4F+D9AgA5+Z8Dq4qM1ZgdvBwq26pqiNhWBruKCJzmYP
FSITxDx6IAjbyhr2TwnbxY8OAKmPdeknI+cfh2hSokPIwbb9aPbFp7MGaE4znC93
Lk8+KkYz4KyDSsg7ZcLW+gQNzSLn9zpqkf3G3eQqdd4/2VV9o4vXLl5/QvDGpqaY
KaiCEymhoNe2hZiP+RlA0IYl4nz8CyK4F9iveyyTv2yXDNummfOHaIwPs5TG6N0d
Fb0Sm9Z5cfbFmnW0iXhLDs7gD9Ax4OQIQGPsgh7neDJqwXwLY2MlhnF/OxVRhbvg
aYHSeTGjasM33HLn6aW7YRGsZWnNHGz4LtTo5ZivhijTxwVvfa8QQAdeP0u34v6J
giolzOHrPiLsYSqzvr2RJJ3PccqUD86z7vJ0IXwM5JdaeJAJPAXeJLLjDi49KquG
85OaQ65YGDR8G+4w140V+9ZnTvr8ScA8AdYR8+5JY69bAFsKxyplg+7SVynvhCX8
kO+GHzeLqVd+VZlk57wqDi2DKhOrQSdsju9c6rY8pOsVMEA4ppT2yTs1c3vb7mdO
wZb/W2amzwAd3gHzv52dRDZZYt3QDnPvMUv4xXKuFi8BBEYPkPhS5zdRhGEvQZ/7
R4DizZSVw8of+ZjEiL3HzEV/LHzVhnwaQWOmexRIOsszjc97U7bme3Z38EIu6bAj
VtaD3act6pbRrvSbxJ2x8T6P5Q9uuYUcZ+ksnw+KeIwPSGkXLqMDxqHbib6RXHAK
uo1c+PpiJ8DRLsErZ+i89MdiYm2ahQY/Wx/FCON0d6WvAAuq0EDsaJTnbCHtgcz2
JiRP7zSg90+5IuoSk62Yxl49y7a+o/WIuEFjpzpqdWnYIBpDneGcc0TOM2BJeXOc
eIFd3Ql/NTfKDhgzKljyup5EzR1UiP3hCWB/EPd/41KjSB//aBUYsSMCqBwPuvdI
iDb7ZGzQcuVK1jApuutM6aIY6n9nNztUJuutLXTBg1zB4j+XQ4hBNWgduktmVZGy
vCPIbBA3S/zv6l4nWIqI8z2rOFpEhcGomqkGF+wE4JF9Yt+P5AwQPUDAXwDNGkRW
weQHzqpjDOLDbVvYv5b2Nd489yOkIZASQDXviqDyT9sYHi7fyWcrcdANW9000nhO
UZvze+lfRPTFnFmJSwHC4EmAIb/7iiOW7lAGknE9FJYmjmsJ5KnFk2wh5IBMSprE
gXuMS3r23jQgArGSLYi0vq4O4pPAYBQZqJF8Go2JMdNmC0a+61doBH6afMUqoHUu
8UR+XULWTv0Qfu5GbOTJCrrgVdKr9FgmINSfaVSqbGhvfYS8QAk+vo3yNnPmX5F6
dNw01H8P3u7RYwFUy8kfE4hnGuR0dA3bs5eaR+pevL7oM9AtZ5wCqIKKr3mqe6zr
HNaLE/lh+S9NUChr/0sRVOPgUOHIDkC/X0zNSXsx0FEtN8SrQigRNJonU1r5cBlK
yA8lSy5I8VEncI5fmZHMOIjL+Syrx+cZ3p3rdt77OJ0CEkfu96L0rqSBhsygRtuK
XkywIGCEs85A2qVqEVLMHRdwkQ0Kjgk0l64iL47ySL4p0sRR2xPY2BwLg4mhQw/7
z4SdUy/3u9psvAPWlGJD9JvqWtj+qqQ62rpdll/VBI5v2YdyNUvXoO9Puwd/PGGW
c4lujllbuPffde+CAALhPUg7Y5q+9WQT6T+kcbFMZxPUv2wkzAZvvZ+QqFhxge4p
PC/chWsbSc2SUa/T+uXwLEUTZqUIo9gbAwYBZ0AhTazGju3z0oG2Rv7/1jT/4Ynf
dWffdAy5qjsWi1VYD68eQ/0twQ42LKtHHBTFSieQDURLlx1rbUPdk6CBm1RduZzL
yPjAgWweig259VIPs9R47KA/wZQAnumPdzyw+koHsP3nxFVMAmF/u/OuOvurk3/2
xuIqxzT+4tiFrX8g+fbZL7USQD8xCUNb8JT91WAXh6GRVH4xzQ8qhOG2rWDByHgF
49+p9yyBJ6ceEGkptMLwIFkKqPMeZLII6sQN7ZAVIz0XhcNZbtbhhyCqJF438K3x
s8BLjsueA5fVl8x/BgcIK6DAruQnHfOJZvOvDRTsdmypIiGxqhTsHgjgLXbZApxT
1+8twFBmyaYAfU0sd0SYCZcgwBc86hb7ZD2XWgcbSCbWGjz2PddhbFJc3NZqA6OS
BaelmcZ/Il9NhQlKGJDsxVICxeEXim2jU72X9fl04n/d2z7p/MwPoYNagcf95qy1
VY52urZVDfXeInqhfx2pRiK34J7pD89NtvM53Z07VsxnGZa7nso08AGwoDhZQjQc
8NbtlcMl2yVCkmBcYmtc1QHbpK6wlxk2HuRz44Wzzo6eIN/LDaMyjVmRw5ifSAOw
Yz6OkLfOuQFyDa4fQauaaY1wznEZe+ivqqQe4ILEMc68XGF9fTcuPoy1F73LWcxJ
05kkxwRmZNcp7SCcGD2p8F8tOkYlfNz92JwVZjkdl/ZPK0SJLmNVPJJcLh8H8gH9
qA3g0qBc6bgKtO+NxU/l8QEG/Npd2MeVpNKOzAbc7EUfp+gy+wMqc9Zr9bSS96Wv
SDlCiVyBKt9UtFqQnJdHHQySya4XoAHxLAs9wJ97tAUHY4AWde2GxCvBlHRiprzR
eP9HAAjD3NHZ/MlRVJTxyHeF/3igllYJ2rGYyFvmzZkNDDLWyktb1WXWce15aBUV
Nm20gTvX0AnEKGJFmE8qtmAcrRSFz7RF8kTU2Ep8oYaLgVBqqq5LbX2MAQccoULG
+2Y30UPAZiRTjPohLQ+5OwtI7v4QxKG9dO9XbBTzAqPFYzT/o/i+Awcg0CbFse0c
affPpqZVUhmoLbgLP8FO5JsczaTiajM7BeavaUjrr062oEyyETKffm0f8hWSbIDL
vMIddmMZVimlTMv3S9LgKcIlJynzBknH/aY4+FhfodFV2lCpEQEJXmdjcQFinM9m
X97gKF+b0bVzeHdB2CokoddeC2msCjqs9QsWri/LV5kQntgKmDUIS/vaVn6JRXAn
Mab/8SdsynuFkO+5BvqoZdOEgO8tEmovRteuuL1SphF/SOBqFmk6346Xoy5NFUty
NCrjKdNyZPICjFgHv+bkXS8mOno7bcqMptOQtjIEaQWImhcGJ/QHh51mRttzi3O4
cfbBcoChPbQ1Xj0l0MAJG0gEYLYnfcgDTPTIyoZEVO4If6A0VJ7ft5ZkM2M1lexi
IMl8cko+1emNWMBpuOL7KDPQg7Yg9nD/noQvlsLCltsgDC10Zz1N9ZYwUER1CsxP
nSVWLszait2KiQKv6zmTjoIzhEHHqtk288s9mL4CXa1oru5EGqu4SXh151Z4IKVu
5iTRaZUmn+D3vmGEYlaf+qWl3wDG9l7vB9lH+6DbxZQf84ZMNxYMKWee/udd0ADw
rViPkUGCyVemnhR+q5L2TWDhxbMjzRx25T3bn2yhYvY8UKCZn6ThMMEa/AkKsbDM
V7lu8SwgB3UUTeyoWz5VCc8EoQUsaTegX46OC5B7nOsC4bPyhNsh4kC0yn8q0WL+
whM3Uzrtx9SKYTaSsXscK1+m5eGgDAYrQt6rSdxUQkE5LGDT75Hc8S2Vk3anqFcf
LPThXtuv5ho/oG5TP+PGJ3Z3ixmHTnk6Qvqd/aXeYimN1WtBxy+dfRMETZ8ArCuP
cypT6JpaYzin3MYFjODRBkow0Ev3U5VNfQ2z+JOEGnTmgaSuuvrpTuVFgMhosRlR
v38rBeIUKzcu5uqVRnUDBBRSnEk4bc9g74gWltIaqb5ymT6vUojv96LiIm8M4IKd
tZARiCVvzavmxkoTurKhKnVHxu+XG6boZxLIyxtsXMwP8VU/XQwPyHAfafyQHrEZ
QsMaNI3+XmahSP7Nb8bKSKn5b1Nn3QoQmmrxJaY0M6K2uu5GQk00koSt0LoV+oxe
6pujIpqoUC4y5xorBDdoI8VR0mI0xKabGGat7dDNobfrxUQ6OgMLWpLpF8oMlx46
1cwt5cpFk4sDCQfF4R8LvClQwetbG3v9FD3NgKS9/Hs9Prp8fK8cvAfoPKqQIkvi
LQ6V1mQWAiAS+WfwCpTP7w435wA9hxgDzoOOQl+GY3whuOjQELhqwYjcbDaCrb/7
NeuUkaCZvnUcqXDQytlF4m8kYICFwyGmPHrc9wik+pqhpbm6i1nhHcvGOIPuenvy
XUawMolr6oZUWIIBupyKKi5d8DYyPqBQ8IsGRaVaCuZ2BY1lI4S+War0FMni7p3V
opDvzuN/rwojL2PVqgZX1zA534iCURyg/M9J7wx9R1p2JjdztnKFwC8mXs37D9Pe
51zqbqulind4NBbO8vN0v6fQTPixjo8i/H2l4LXl/YBJ8vLpXFMX8CxYnfInkj/y
LbsYbLPfg8U29Xq6/ldbNkMCOfz2VW3n3HsyM+F+yOmoog2jJHeLgUw0APUbPFte
337MK1DZS4yHSxxQfc4kts978oYQ6biqkksDgPaQYJKt9P9RL2G8GQp1MFFX3Zuo
n1+EDXfL9FMfRdWmYriVpaMI5E0/rNboDqb8mAhbyVE8zG4KEi88jQvhV7YKfc4I
4I9+lyetkmAvpGi+qovIOlZePa3MUKIHMBPdm7zC5tdfyJSMGebk6b/jFl2ISiYs
ssJVdjfmHgSdNlAdaT8dn4O6/ZrwTDawN2Erv1Ts/9wmz0/b9K1kcIHt1zBolsvP
K8ysjFQ2GhtrCnEHU9jofwM5RyoxO/lBdRzI7GT3mLL+ss+1S+XwQXvbeiOB5oAo
i2Uag49UrZb3+Wozo7DqUtwNIdX1e/Yk7f/uqhrrpuo0pPmX5jrUsGQ1Vl07st93
oW9VKU5eWEc9lkwc5A2IAbG34ZbQV4ur4BErdeoCTp4zJl/y6xVoJDkU8FdkZnhs
D+Frx1+rWXBJJOoprA96aVW3940Zbz/HfVLtJpIIAlEBbPLAawduwTKqlBfz0PyG
3vQL/78+Jttk1u27ixt2sxm/PqkDUZ94erVNE9oBrp1h7d1AVun/Emy7yUEuprdk
VkKVG43lIbFHuVedTdUR3/01FGCCNVnyVYF9bgUI+ojFSGjbmzzBDyILFs1H57ep
MzAYOY4GXzVYffW0ZlubQZI8mE4TE4h2m8meveZ4n/K6oCSuw2xF1qVxyd00Nj6b
Fnz0wZcpxqsbAjei7yQqY+QQl+6cff7kzdxRkJ2d/mzwdkgT2czIyzsdKxabFZSy
nPIozvOjiTBz3NKx9KykxIlFpm3VlJPjePcN5UxSJZgYKZWGNhJsmYjmlX5SDkuT
WJ1LlJI13Bf0+MdrWruyE08kHReUHxZgyTTHZrRyUZOczSuBNaKucS7rPamt1s6s
WaFwEc6qHng9QwdcPGlNnsoHqtO5P0y7qCyP/9tMlv8bm6Nw+v8SrRLw++Np0Umr
h+8avWWXxa2F9O42PFZt9KlNi1PtCZlZHUEbwKR60ZlaYcgAdzAjQMyflNkyoHS2
8EIA4urC+SQmh9j9Sc+uVNlp/m4ka44+94Mx46SV+PF1M5jt3nw+6cFCokI8jqL9
u1CJsWjnjmm7kjpdpWa2C7dDEkC6bOgmnFbjVxcQfyD8mKK4dY3KvqyJu1acw1/E
GB7LtmfD6qyx4x4tsitymjn2S38ERBFDMVGo4/DV5zrxmWFLqWLU5LTniQfPPefn
7wLy27vD6IX5BqDacdBSYWk/8wzpivU2IY60zPccVvMRhqTm8T/0Ej9S8zTQKPAg
vrtVheXD6ehwdsK3m3+fnVzQrratxg1cb8Q8HhQTlEn04gP77d7BjYp1UxsGBjVY
zgak/Rvai1/FVG+y6oZbtVt3VoPoNQrlZTihB2XU/QkwzNmFqvuyeDQxy2vVztUF
wEOdxu+hwB0bdFsNFDx+1ggcNFzuozTU4Dc7D8EVWidN5MhAmrYrVZgKUWN9XSn5
H4Cfbc0Sp9vND4bu32EMpnhMJvd7dc1rSBs1eFM+0hGVM9fgmQFKtEkYWg8KACj4
VzAK3Bp7pwRvtFTRgrV3y0qd7zxRT4Y0GarpZ2we1McSvwD52TMYsTSAlI0rCdQr
3znCtKScr2CuKTeUwBWEaI+yJ0+9PETIVlPDJeloAKTwiX2vW8l0+QRzWZQb1eFz
0xEUeNIqYpbaDXzz7XK60lVoyQVjhtxw/powkkVaWgMq/2kW+RkIgUU3waNXwBFj
FWBaDVcGV2YUXzFN1+3mQEyu2FmnIYPXUbTqeyvLMwRFzwA/VMEUCU2hgEI+r+EU
8T8HxHcZuMYzl9x+Hjz6sogXGCDdrdYdUwLn4FW2yq7XhutB35Z5acqT6bSNWeJU
cEynMh994Rp0+gS64fgM5TdyfPseIqIhSCq6Yomb1xcHkKZRYF/FrMGLV3+7SSOn
YQFb51HCfY996nLYRRmdY4QWsUgAgeizumssaJ47zXgYYQtRpiQ+OvGOukYySrZf
DlPTI4hV+kGGYaBm+toTaIWuGCqQSxVgAYbeIqRU+NF9DijWV2tgSel7AfVlYZVG
tZk1g3fpKsgZr5j2BlA7QLK7POKJt+SUUBKcgDxG1t7+EBasVBQ6ySkqkEsUAKSr
XSWtUS4waSQ2yLf/g8biQfxwJLQHMMTxt53FdWJLrbgtzmPglrZ51ToqJV96jOd+
bLNsPh17eWpte3cwG0O50DekCcKQCrxTvGiucHoWrgH/VqgeZuHAJFCNP5yNWVvF
SAPo/nwPi85HT2rj0Qk3NkasRs2mNaiIXhd3fuMcyWOra7Nzzg8oS6UtX5yk3WbF
K91/0WYgtBiVYDdIZcl/03e8qXBWpx89KKIt3eEupHzjdKujk9ryXnB1WaliJgVJ
KsxpllWMiP2loyo9odYRlTjKThrZX+2ocDX95TTRRnOtye+FUNGbAenIKti89PPh
fN5Gf1KTh3rkKOGeiAV7RTCbRQu8eVfW7Jjyl23BPIUKKh3MJooaClBDI0uzHvdz
sguwkAYxZYBQtYo1+LV87acTpQwLaATik9amun4wmpsIgWbfyuic+lI3/4Ot52RR
SPAF9FTkgEZID/+ngnp1tiM1YoZBtUCo06qmg3dv/zzxfVb8a092bMBHQQoextfK
97UoW2DcKHNsFtcF+IL2fHSBTo1qtaIHqWlo4WIHyyYbEoFnMKR3ltEh8+7cHZ9p
gnisH+ZGaQCkyX2qiRxXxul2znvlusfxVHU+KeBdo+f/4KvLDJgqtjtAoMmon6f6
20fGOSRU9cQkcKTYMG9P6n2xppGaQoGO0NWZ1YQ1qfzs3A2FkzGvYdDEWLb7CyPj
/dZMc5ZMPV0ad7+nNsvErsyFcVzrGxK7IsYDp30s4CmAu4dZ10FnSpU9bvMqgJsL
4O9vI+mjAu+TTBvg1xS2aTfE75HQYJbp9Vwy+3pQUp8GiGsRN10NNPI35gcQNley
O0vC8Vm5rsWkPtnv2d7KYHqbo1JJcIWSh/rLhZm3wJfFbCzR1kGP2A+iQtauCR1U
p2wihahQfZmHcLTeIuuRytkCNy1dOLR8Vmz7vxhHNrcaEWA9UHHxhgf21OiJ71/k
rpIe2MiUbBdUMw6C8PuhJEnUCtiS61gCz4B31kc6qXFzOPGLbRE/QNbnV5afwNCo
67fCcO8DnqPJNeT5+cVKAhpPSoWzrOOm9/x2TCgdanjI0ITQBavvMaKX4rD4wpah
dobslC+nRBuR21EBv5OBKhMQ++j9MlxafsiFH/+eIhMuMO01VjdzxFFupswnsOtD
Qri8g6hQppzpWnHVpSxJFFoezF81jcuvgRyRRGxMOd+WLsDJca7qrem7hOHm7AHV
bSy9fTI/YhPz/zaBbxkJjfeC4g9eGHciYcFA5Gq2D5zcHTLkabjpuhCM+QHx+AOn
r65ThcBTXTnLcMf87TB2g1AX1TnWQmBaN3FltWlvGFT25ZN3OsIgCdqJwlT3o4Ge
1WLCRDTMqvYOTQtAu5GWX7KUqgJYjRxyF49yKG+x84vxXmFPlfpEQ1k4hLRPX9Nk
fRMoBpIw7olcXys4kpiiPnBBtS4uA/8qJhVNyRUUMrP3lQ80ejdAByGJtSt0n4vS
d0LXe31UHlWaK9vhmoo7+7RTbjSJi0U0iUcWtDli/c57vdLZr1XdL/rFqrWEgyO+
A/zG5GR6s5BlJEYwBrs+TIj0LKTDvn0Ge2z96HcHZvw1ezmrNbZURnCnevV0zqNL
fMTqblWO+AYlDvAoWH3czu73ZuOzXiidmnHLFL5uHl3UGdW2BOCSUAsSn0v5VWWq
K6M2rizrIcJ+0EdE6gRj8O6770fQTiXkC2EKvOtpGPfIS8N2Jz+oFEcfKR1upZpD
XaunkSr2T8iqytq49JFsbyE2MXYnzj5pgR2E1cBK+SQ6oTJUx3D0M6EA9+1oBMit
bc3+hotnfbd9kH39qitrhNURwtC9fQvMO0SNUhR47aZ1yZWeBrwqsDjXeKNNtFij
3DEj4RrpdychOb1rjDit7OEGEQ9pPN8hNHQ2vlM7AbVEalXD6vZcymaNFPgAmMyl
cPSYZcKoSHGctJ01mV9UspscsLZoy4Hrh/W7L+vaZksW2habGphQXmAvP3jXZGvA
oWXjkefq41pj9X9N80563DiOL/q9q09PNokdw2yolNomZR50SaR+58ty/j2PdYaK
jG37+Nge6mNhVzfV2rpb/NxknqwEEkk7ModPf4vB8Bjx6Ld4ylsGvFv44e27z6zZ
32IV35XKb6Llj87Kxh8/tImuH4FgPWplRh3LNJ38BXpivwo3J9eS9Ky2xO/OJ4qF
luIUpR8cf8B7Wvm1agZUcaBUG243k/W0SRZv8C+Gq1mUxzO2MvgXzES9lMpfioX+
NTsf7p6lTFDktVuA7Fa8EZ86PUSRCkktWCJzcFNIXdxKSyVKk2eV2Z9aflShJTGW
/ZByAzpM/n0Ti3POfcMDjyGZ/KxzQoTDOewstkX9Axl5NyTB1+2sBIN+9i1Hgrjg
o/u+dQvjOQWWpooQQ/OcRW5bFjYZK45fJ/ymKWcVjK1MSZh1D9rBItyC2qtFkRUD
Kbd3ma0uMAtXGWtUC+f+0iHG+DpFqlLC7IioCeLbxwAiDO17sIFtHtJz3sUgxnTX
WAYCr/f0Ypox21CGdM8zvTbJsHsk/SooHfbR6C35/o+DnA9HJNYZ5nznPSMUlAxj
msv1pZb+PBxcE0KHGemsQpPtRF81XzARqaBxvkpxzATNFjKwP7Fs/PM3tUj5asKd
/dasQp+3jLI5OA8Ht9uXHjTQQGaZaGHD1dbzhY0WQRieAEumZCmPCp+TWfmLnJy7
RqAfy2MgDcceMBGV+5HojlUOh1T6+ByG6KLno/hmRvrYIleo/CBB+kYI7ep24HrI
ztbquaoBAXH1ydBbUCIopmcUpv1sptA0GXo9nqb49ZhNCA6nG9X1ifybMspxmYTv
y8aiqvZvo9/BK79OJx8FE3cNZKFoMhj39qD6eiZBg7lYmYFIQkPzOzfSCtwaN7hl
REcsZsYeHdYU8bahk7tra73pUpX0Ha5nZmFInG3MQmAd0bQab/88dvKw/ILynMqC
Z5EI4PEutTtcpbf21qb8vj+XZMRcKQ7WGbGvy8X+wBQZWBfuGG69977YuJVMf1wB
3OwgIB+F9aIo7/KyEPF+PbvyE3Z+nGDKlnPHrGN9Rjyge4+rUXi2nASTuT6icEbV
iCVM+adWRWQ40FjJmXgv578RI5hNwzVyoEkVEDRLsGra7ag+Hs0gHyEkXTLoS4Uw
2EnaW16dn7esglOEKZs22yn30avB9su5BGsncNeBTybRpbCinSxEacQeVAj82zc2
8vMv2Lk13OzqfVPlxXq/XsJnOyPAiM68t/0MyIcT9V2cBlNJWotSQ+l67sZyx15d
Zyr6aFFxOHmPSN8H5hfMXEOHbhy8IHvQckd8MeUFCS2jMFSqCmlHqVJUNRX/knQv
Pgto6BajcgZeMkVTd1Ga5YjqDU817Mg/uwqG/5q+v17AI/ZpZEWW3eLiVHLP2lUM
XmX7GvedkcRBWHAI5F2r90rt/wC99aGUYk99WMB1Eu8Luq5fGHTRLTY8Q95ARMHZ
x0uTifX+9vFAZvzx4QcwLtibZdAfPC7tQ+M7epTE6zRlMpQux8cfAtqIm0A5aBH6
GbkpU+W3sSGQ/MSWjV1tXQAGdr83vbLraXFP4QUdNdnn6SN3/xYKWNNcDp1AHfv4
AQAPgRctV+e9nIyJbcxe0/ttBOdXuhEwy0QVPGMUgSPMfOGh8gqelglrmd4JNMV3
ErvtDlzrpRMq0i/VNF5Pv356Blq/Ig4+NIiE0woeklebmnogj4pWpY8arDzfclsD
ZK1wyymltcYy0Phrc22ao7bB8EXi6FOwEKa11sHuQ6z5W+YDXHZqPvbbF8EAwCWx
BNiC44oKD1bLF8Vo6bJcJ3/lqDrdk1YjOj5ENfe8jPWeUtR/wzhfx52T8WxDcn20
uER3auAX4eCom9EMQdHN2Rb0hFpjyT4M9XOvJqptbOsFBgOtxhQloR4zn0Svv0lu
+lRvT1DJObLhEQeS78cJkzpo47JPjhfZF1Un3mCzn/ye1gXijNTACewvUzLi8jNs
QprBZRKujElB4H4YKQ5gOsDlGffrIaKEcGXKZMzmw0b72xL1mD9inRNlWRjwhrPu
SIL9s+td1FtrFJf239otoYel35oxmrCcH0bfr30g5R9m1H5wK9ZTR5eTorkHu0nz
7XEorHcRDld1HkHxhP5VZw+KaNS1GJtB3smn35miQG0XH151WEesxoLycOu/U97I
OFIBTG+tf3pvxpLIzcmRVszj1H+nPY/3BVYbM8Bs8enjX8OJzOawimiMLjKZ9dqC
TKQ1l6NCqpgbBh8WXaGITX82FH6D07tSqGAzv/12IrNGhflaWD+Qnans6IeHMZDb
PA2fzdEKJUGuDSRCWXIC6fZVcQz7JGKQZWfZumiQhh6RUD04oV6gltk7eAwNls8z
nkAURsXANUmHoAasVlkjzgrsm5qzAGnJFeO/kEt8oxxcHa9ith3EAMorSn9CSggX
dxnElcL67zH+FASjl6Z0K9/pmzDe6vsJu0mDHzKg+iPNrZF6nhPnfegtyS0IaIG8
cnLuHZbJOJ+JqFxmsgYiuDjUkGi2b8Wu2zmtMxz91vrE+IJd60ITWWNO0WcPEitd
SJD3lop1ENyeXbAf2qsBgwyn6E0Rg/W9InrcbJAdNOqrTB0ma4RZ47IeCdEQvAvf
WQDSQKGzguilX7BzoJGzIE2wZ+CKpZKqXhe0PyNSbTRyYg5LqUvVgbSz2DROWIgS
1KF3fMjSPZ6EJM5iSrFmCMCfQEW9zZ+LuWeZDM8mMQTrzVRpfdZZv5hdwXHZjgO9
NE9PjYAB97I16ZPF4U4qYCT9Aji8yAdwb1ykw2CHW3YSGELccBOw6qhpGpvswxmz
5iTCrnDHDXuxl1EzrfBtlKSLkHK9N6qDN6Sd0tXPgDk6ybSc6nwv4ALqLpVBxw5c
cJPH3SNXBhsel676FRPNBwfxx28HzMtHoQSeV0Sg6r2pqxhZ49SxeST0TsV3GM3C
F0/30h45Dt756VnfMulMS1wfaU18shsWoK7AbYYLXamnwm0l2axgi4sWH3NBvBtF
udZrvFAy+Noyl38k6dq5MxVlviPAwt2gOkkcYVxn0gGeF4ZC/41fQTb5Wtn8eMNK
fWX0Ad475YPtU8jZ14U4DoJdHUKVhmX4vLH60YcLdYi/NQX7kJi5MVB2qGUBz3Xs
hil2HaeugPf3oe3RmRsmnO1v0Xb9cDpCYVjp1RQjrPWJVDcgx242fDHK7ssVOnP3
qD7TNJb0/TSUPdZW/d/XH44w8i9mRelFjTbH/taAtmKS6/TeiMaZB+U+Y8ab6705
OAvFdKdioRKXbmuIYO1xrI7ptlqb6TtxlMpdb88/GkoO80Dyq+S1owmUt13a7H6p
4Qeq27tJjsHmP0/jWrQb4l69Ix34YZ7zjHadBxLB2jvy8azQuAaj3Km0pU7+lplg
rghAYMm8UkjfoJpKw36T3u7EiicfKhQM69m1Vt5NxgP7aqdORYDzXYN47jjcwZKT
pNWQl9whWZe2CCJiH0ZqaosxdfiVB8UNquety9LudZ4KwRMxuOXy0zCT7HqtH4xu
+cbAc5APrM0l7uysYt7Ex5niaTcY7pidDzO3Iwqp/C7F6t9oCBbNYdrbQ3kDihr2
r4Hp+ek1nMw+m0dTScpKNBSTBRWKE1tPU/r7yHHfA+ffzRW5WOpD5xYqBdQXCN86
brCcmMO6SrAAzsQo95kjEoDavu9GLjG0t7AV8T5XMAKDu/dsURcQwuCIbD04Hvy4
eO0MJyWuowrgeCRL89QZiBivSaw4FcI7yhhscQhc9bHTLtyIQ9WLkrchBsvs3ZaP
0Bb53fARZdnXqkoFuMjIVhfFyWOj9HeY7UqCmTZgjAIFMVkF/OQkV6RKBEjm8huG
2SM1/a6iUJn3W+JNc/CR+LKmGbcNhkYl4oc4JcK/aNMvOZ72jUhDPRVUnMRdKEU4
dsAFMgJv7bHrDBvZ59PP3E2nxO3PJKzXSEF5QaOcnQ+tw0P6MzZjAXSs5SPJDFF8
aTOlSIXK3v3A+P9GifDdbQQQwH7leRimdhGx7tR2BSJCzJHMKXge9zG99wukTFvX
O/4gAPVvuWy5N2eVRLNaOa5CI0f/3V7XqIIGssisHI++wAL/jH40m+yjiZuUEMUA
ROR5qNuyEeXmZk3RhfQOHRaxFN2NbkoofTabFbnnRygFaWF9kpXHm2UchqILKhpb
L83O3GQQFC0vitLLTl+2J2M3eiCm7VtYyIA/ad6a+/p2QnAOnhrxTv93lmNLUG0j
wewd5z6/FJ9D51UBXTiU/CJ5rx9LiA98P0BZ7byvi1hgRf6PNSDFkGZRNPkVa+A2
9DUQEfofnpqKUjzFOFxsj/T58fBAqr+Q4LcsTawKq6nPXKteGN+GSbWLImJDdMvN
sdMIJ9lEdNTJlCMQTFG4ynfMEDv99jTAXeS21L0+XMqBjUWua1yE/NehRFz8eU3A
i2eoCBmipAbKfIltXJqdMx+Sw2l/gck7TDson8Tho3Fr52nCTf8OBOEp7Ydtp3/0
Hia0hh/vfcaWEIQcLK1oJ3jsBQNiT5d0rhrysLQr3yLfxYYVkhWYCjKaFa9rCOH7
fo/IFj2qLbCfswZDgSS4CvcUV05lo3QdHpHOhZrnT5DuX3Yier08e8jAGe0vgQmk
uP7lA+vn06/fHmEIfmUwk0N//TYasyHTQ36ridfR4SIrvVUvbuS55P7QaAMwtvf7
Ux+2pHC6exdg2XyqHTM0iNmLYS1FR+KWbg/T72i3426UmeSyxrg9+s45x1ULBcYQ
HyqnnTY+K+SymK0vYQY+LO0/fLuUJlIQXeqQr080V/NPr8nWXP5fztbCB6J2NvQu
a9sSunMMk+ID2af+PvE6HIxWmOms9nc4oG0zwGGxHsonjeknVnqvly2yDdN0T4UK
MyqTSGrBUIBmXkjkLnsiH/jl6Oz9/NhtFGjMhgfzf+gPIz2r1zcwDldezgmOHY8c
nK8XssHLzfwZPvYewJYDb5L7cccJJH4Fra18EqOrSMvhpJnINFrsd70IvQrrlw3P
UK32luQ0mf+CIvmbRPyFSuBgxLez/+rtnCQc7NKFApmnwV22RT8oADg6werlnHNe
iSZYn4Mf8N4Xiv9mmMczQc2Ng91fbYCOx0ftSshyK3i8JB0p8HYOIo5WDr1pws1E
B2H27pvoAow3kJGndv6DgaNNHuxZx1uIq5l+/Xxuwf97RMV+9Jw+sq2YeZlw/vhR
XwQe3Oiv4KJ2tCjLZR80MCETU2a//4vmUULv4ztC2eJev99UWE3vp9o2S38tzLOO
9OrY8A0h3hwXD//u5LWpEuhd06pQt7iLF7K8AwREjbUjC3ZmgP5b+oaXh1aqYWq0
jJD0FDOiikYBp6lnsXh5yYe+GOkLHEkJLkYCday4VPEHPmA/YPKeCY23v6e3fWbe
7uPCUQHrxngBYvgmfj6fxbV37J9b56bUZ0d28cpgsK9RtmrUDoJvXuXoXZA5D/u7
IfC3QFvKPn4VHXrnaed2yt/hV0LwVP6zQFOd152OvlOsVRaphHA9RZKnRBw1Ehoo
CaC2oCGGbkqqfMpbpLk/MLU8BBU9GgwU+x2LEKZvsydYql/BOdu6fgbPbWjBHIGa
bfPFf4Iw+GQYgyQF9OWW8yUNhQ2Kc8rs+JcnTae7zCRYhtoyi94XdQt40yjz0YCX
AJ7YSwvY2p/3lKYnMWE/2C7rKlYA47GKDFi3fstQSbXL/XXW41Vi7JdtwQ9MFX46
Cpi+pu3itTmaK84zkkYhmY7MzhHioWeKxRzhOCB4MwHn/uEEhdMxO05MwO1r5M+E
pMEH3mqSFETiVPoKKD6H19MxQmx0u4GxJcq4UBQylJtBdPJrrLGeW8PhjQ0mcB+c
HJ3smHiafLUUr33pDChI3BuIW5SBhyTrCXXKMvc56iQtfFzub4hp5GI+McTuEpMw
XOZW5ttGrufTWHQWmg7B3VrQsgIYvyMrnYdFpIEJZ8059UFQSroxdZJPALqyZBDR
Rzu1g+YglZK3eqOsvZmy3bneOPeTccAIjAdsyOwaHY+cO4jRPkoJt7e27ypE08Bk
k5FFwFwaAyrBqTI9YezhA+//nMMdcEMqxhkDDAVDE+2oXNEcE2q2q6eNR0MWS+WY
+sQRs2WOZG4FzWHqg5EbgMbDXBlulblws8YacvJQmLZYi8UtB0NM1FJ2FV8pmtDt
9YmE+PiuTs9NsalaqhlCfu8Njt8HLrsHQ9yyDwyBcMcmETxtRkf1ewQy9+PGQ7Hx
U/IVWGXPTFZCwS107kgWt7NpjF8NINpDh0QZtSFH/xzLMJKtzUs3uefakbv60TWR
oVFdvrWsZnZLwqHvhbN5ZxHZmqNEEkotxJYIzlXOQmP02pYW4aza2OdvqX1jnby2
xVIwSHk9ogKUjVCrVhgDnf3/z9xiD71PM8PUdPqEvRfnIiiIQz/tKd+Ih6nYhSZh
TSz80/iz2uKpIS0zbDL/ze8A+m6ZgDbCyeJyYx2e5TgRJntBiNuEEGHtaQCSBURb
tnT9Wod1tx0UcdUu4v4Sn0DLw9NLfweyWLEE1LDe8x+oYXR1szK9I7ulbPAsqdMf
9vS+pe2CwsXCH4ZpZmNPGZxb1pHnvNZxHjN3WaFcZdoyAkeqjCuWh8P4m2ob7zLU
i8xKw6zlVDn118pMeqm1rzjitnJxv/aG7zg0TqNFYIfUMDzrZERz4uwDVFSLSUIV
3appV2lvVvxcpQJ1q7bhUWqKNJXm3p4YsuoX6qPxq2IUECeZdNqfB5ORVGN+fm+n
EAG2aZIPhEhHAj0f0zCUByhDG16o8M0VQbJYYSPTg/BCZKY7gjKX4eFnyDWY4cAc
vBF71EVld+2+RuK+gL9kmzkgz/pEFfIf/AhRBg+ixk6kwg9a8K2EuuBSE3Wd10lJ
jueNVWKMGpzsVTtUCaDmmcMXbjH8UkxnIV6CiuG14+YGz6WRRpxFGI0K95bCUl9r
BaT9iSatEsp6k7QZO8fyct3XZ7AyF5kTfMpykco88Ew6oTHZ+8FoqOqu1iyHKf1x
XPXZ0ouUGNTUP2MDnrEI6jBq8qyPNStl/Fu0xob2yCHPq6QGKOPEe10EGyswhx3B
h045vu2Ig8JG4O0O57rTqIWEHz79BzS1Pnf/uesuHgAvS1kGyuLaljmFxWS+lomS
VEC9G0rdo6eqrYzW4gXPnxopvQ69hDjHIdcntP89ulqseUrhnnSdBKEMRFGqGULL
RCak4cYnJEFOJLjTcAB8gPyNMKROsCwFixavaLG7EQxWY2QpPpTK+Amep+s8gP9z
ILllASXNP0+5I/HCiK8hInajVilOPOAF6etnKF39JkKsCqTnf7TIobQz+aDaxAzS
lR9RTXpOBUqizvgJQzz5Zsbtl4E9G+1RJzaVcFSYumGG69PwPQmJWyAXh7+Zj8fg
b6dDexWeEcKmJblY6ktE3iYxcsSXq3Ar7ONflH/bcgxsDL7KX0jx70xXo/9v0sQM
pnvZbPwC6+B2+HN1vRjcJ0/GSR1J8MQ3zKz0OX2/aC8o07Y9/3r8aeyI0nr+pkLq
wbcsYIEgvd6yodHt3Xk7VBDHW3PxZhTRSXvuM01DUNy3+OuyDnlUfDpV/C5pLcgd
2YCv2YO6F17QWsbgcE2hMgTgun5Qi1AMpQqtw7cbTnjBuInt5iBtPj/m0DJ9485B
AwdH3RxbYkelfLnlu7Ns4xb6x1F+D6KqdkAkAB9foM1e6PpHcubxsP7S3c5cNOfg
rI1kHYq4oDH+ee5b3EsvMjAlBpHbkzlZxYexE/HU2LUq1butZfbshLFMDsE1X7CZ
/0TnVscv6rtQMvaMlFC3wxM1EL9Hd7Or7ourm/u6EuVmsD8Wo4igc+So7Jlagd/y
plj8lPYhwcS26jGrUE8sY8741kCTmAvBb10IiKgdOaAFAfDbirnnbt0jOxarJv75
YzseJmRu0DGSZQiEJvjNPqPfsi+O+niJkl63jvcDY1k59yQwPn/0oifMhsx49tXW
Q7e1Ra2CafZwQMfB4kHCRug/Jw5e+/ffUpZDoqiLUUmjemJVXwwk/nkUdHdxELI5
9gOvoyWkRnf76TRjzphG/qPvPPKuhfWGsWdkWqtwpI2JQV13BZxKpo9OUG64E3Yl
RGxKn12KQHKIiPSevY99SarjPQ9jZ4oT0CSB3ZdnW0tGEaD6LbQrOKgjtId4/aL1
BkCXS+T8SbGUXM5D65E336nBryXYnQBqL+76YpkQqbXN8kR/JrWEl3bIR1g+RneL
AQyl+PLQdTy2G/Kzx7Rk6T9Sx2ryTGscJ4kGSAZHH39gcmx1/86edTCCrG2igQvw
OvSqX9cjX3o6W+RdgAoyIki8D4/HY1xA7DJJBpDd97AAAj14rzVR9gLa3AqhFNPv
tsuxTT6ECNmFGgfFWDMa9HCj/TtRDtvz+/DMo0ea0G9H5VbXwL21OUFfqPxBVfnS
fUcmedYIJrR5U6Zk4wU3j1KBlVexsle6LAzd4XSm1c5JFQ1sFUMf/pGNeRdWDw4E
9XqLMv9scSDYXvmdsN9v8q/Jhhle5JqZQmz3w4n+KDLk9Qgf3sY1Z9HpzpZDRgpX
sd0yRBtzrMfybA8V3IEcQMy4D6zKVtfGWAwwm+C6r+U4GABWPbvoIKLi/sfBgdqA
gHrDDcDpemmSWbdOOw/nUF2e7DiEcKfnH5Mhj3e5na0O/4FGn0zLoXOODR1vZtKz
jWBJPK+7YoQiGqbYsMvADzRCOmhKJSB6tZTaE5P2wrdqaQGVbuUxmazNIRf0gohO
Ux1+lL+XTxcslSkDZ3B1B0cNad6szn6YXx8AhRyrUNX3hV6wcwEboXukAQ+p8HXp
GCt5r3kLxUrJ05tCkbzUD0aCMjB+eyM4IAiEmJFTdT2oGK3lE8nX8DKD2cmGBI9N
UAh/0jBdbELf2RwqII4mqabYx/BspWFMG0Z3FKLn0yDsyf6nt3mT+6M5kRfN5N/R
5A06PIoTEtbdVf7mJnNDC3VeEunPsZBKfcOSSzCYAFo3j0iWnIMD2kd88qs2fJoS
TMmk7NTfMbM7CjqDCthwQEZx9dTWZRqsXmS0CZtJ4hWlIoNQyIAdLI4u4hnK52km
aGGHQaaWMHsvN0HuKpR2v5DiC7WZ+SrJzDxSp0epPloTvw5dQO3OvAT7IYY9IVmi
MhLodfx0dDJTJak0GCqGI9dulH2cR+rM2/iqHyfqVOSGLe0bbRiiQubYOR9ev/C9
f9G2qyF+E3wdtwg79CCgLPjGWeML6jhHmEDGI9HeJI6O8Wr1DNCiXoIzF3l/kjox
ppz1GdzK4IaxYEtsrR9yx4SV+3lOxBP4FlchmCRAaT1fd3OXpapGWccRuIMy8K5C
H5Y41yXxaKB+viWkwJrAxcGYwotBN2eJE0nuumvMMh5zhGSw3wbtwFATgtwgy/rI
rb1OUhBJ+xOpz3NyzGus38t8reti8KRAPRwyl5fjuQ6siApnac1/FfGx8+DKxF9B
B8ZI3Imn5HskI4p5fwuU+4JxRi4OUCSnIOS8jMVVMFQsddL4x5dcSucq2EQ8CQgv
3580mWcMFjTdrJ1hV48v6D7thzELsNycHghA5a2blNj3Bur7jevLBdh2oreF5b4B
g826xVKv42vjFxCQnWvbLDak74jMbmvUL9EHlJKywaHzgQN1hk1yGaJ84B0O2h9X
9QADu4VAYBHHKn8rZDB4H2yhGIx/+623vfzbZdxAPgHUBTkTq7Z7EEEgRI2e6nv+
3Ghi1OYid7SpItnOtuI7WkvH0F++Fa3OstvIwLDDbHHpLOeF7+P7aXepgqMrbrvO
rOhl5tH0ZCjsTSSrLDNOhzAqoNNuav0hW4mSnjWh2to61en7x1bYiW40XY0oUvJL
wGnaJInYxoLrSrfywP+D/C9S4NS+CSJkavB7hbyViF1/1pnyVke1zVb6kj0+8Z/v
yPH7VXhFULbwalvu5PlaHvYR9FoY/HF8Wh0p/del+9x+n/rMdDTQaEejjCI0yrML
V9/LLe5cHqHpt0Ny55uY2jQlGL+Y+5ezvwDs9pkDeHokYxgIRdEdR383lOxhpIuB
vV2rO6osA8tWxI8G6r2Cha74Ox6jqqNy91GP7+JA/CM3Ne08BJ8v9gBaX6+9vvJs
dTiSB1xvmwlZaDljKUu1oY3cb39BHw40ZZJtVrMEgvntAIE/jxIul7YnEJzLI2/F
oqeENY77To/wsPkuD3DHGFOfZBghLbi8cX8QBpuHcYx96GCvL6Dx/ZH2CGmnBNb4
8IicxZCTRFrguP4e6coxWwFq9sKpzCW5hCWh48Md3RaZa48dWxr211nDagFjnCkY
oFpowQI7eKeIrEe0tvXIySXpS1eeP3kq+XBs9krlwWmfbAKvqSu+H0VdMiZnBWAx
A/uvuhD4vb490vsQZ6ooN2Bb4ZEvXRzeV5nmhDATiwKLtKfl71Td2Hnom8gj49++
LVfH869cM+xq0Xvcyt5G9I4qml2dkMMSr9J+C+XsjTrkO5U8grX+5//PJny8XYzQ
Mn168B1BEP8NfoqWe9oIpvKEKmlbbwkL2zqw+Fn2/WXqMQuOmJeuYuBO8+JfgzZC
Tb9eM8LMH9dm4FljCrCQvgXtkwX0mi3GSAWclU/W8Of8nPV/EYf2GOynwei6CPc9
Qp9ULPk1bB+0fuO9CMtmkLJLM/Fyne7ThRiOY6kSsF7h76kT4Bq65kc8RPcNucEE
xXMiA4LmBplpA9qEnSo58BZHPHxjM5fAor04Bp+O7Vk1I5TRHYFD6lZ9zXHC5XBG
lVFKlb1QtrlFhXmyqXXAhnCA+Bz5GWppo2xP+GprC2xjMOq+N/uUuKPSVxUh7bxy
hGrsl6/t9vAKrH3Ovu37/47GKz1XIZZ3yydNgnMdgfWLT175NXl7R4FcgOOSrox1
t4vLoMX2ObBelGtippH4UOFUPxAmzWQ3KaLDbhL1CE5f7UtoO+Kx+3Gu1Km3A52H
PDwkSMYI0Hdk3/01tANvsXwcT9Nq8PzyvVyDom1Q4QSKIdkKT6w/U7cEGmsDe93y
+5BguN7Qzn3/1AQgK9dt3c8DSbr5RwNiDeButfSiOGc0SxB5tEc0xcZA+J6mSGsw
nFuBYY9Bpn7xsvqd83ocj/YIQtgzItReoLUSWAjPW9DsCIJgUB4GT09cFOfRL/kg
n8LqN/dUVobdKUBXb2DdXSNN6R5utz1HJlhTbTN7Q7N9D+AxmNmgjD8DBjiyN36y
aMVgPBFpnPeZfd/7uSORjRwakcm/BF0kybIwgO58ZyKALczXh4hp+O7Uf605mHQK
5xPhh3pj/ruy4SDpMn3xv420vfa82mp7smHKN8UM0NDgH3Pal6e76baZH/uxYWkX
zH6sr+Wqo26Hft4TU7tiuq+/doryPw3Rgdqg5hLiXGsGFIKzJvO5g9tIpuIjnuXd
zQSx4n6eY11jbLOQFQwZxBiHktr4w3dGQ1138nv3qlPG4C8N44rUYjcU4QG4stlM
cJ5+ns6ThEngr1WGdD+FyPKza66xMkwZGJ6fbUwA9cmLjQOkcDaoPDf+f4An5gHJ
m7jaoPYZRa3YAmBHf7vY6WCOVJATn18VRJAni/nn7x+nAPwDi454tJmZpAPGTrcO
hcKoitftiZreNN6rw6SGBnrxUe4pfN7nm3PNTZMrj6KqQe4xjBvd9PxKWTYv1UVa
V/ZsTzbzFMgQBfCpv5QqDRtuG+uD5FfasuGF31ZcS/mOG0DMsiUxnHtJOpEUHGw3
aNa4ixhWoiWaliHbB8lM4aCROWMKlozXdTKqCrTnBff/EQGoItTSsdUSLswQXPt0
Ts3i5xSS9BQmFyAvFYo8YaFqNf22+nufKdwS+CClZEfOcv4WVTPU+0rTux5ELH56
3lZMu0uyYK2yLxqCsZDEODXwIigyDNzyekSnd0BbUPZ4ZGd60QIGA/CRg32210vY
R0G/0DJidRJI9mrO1Mg/I4Kp7Y13Pq7Wy16dVZDfAK7iYQGaRFSutzSwnwiawlVw
g11fJWhnh4WHSvUTgZFVWru9yPwSP5i2Zj+LUmRbynSv5KJOm62nCGfjsCZsAJt1
98ZYOOal3/1S/XJNklPh8vMB+5AWOf4WFt62g7OQtMsrlb5jFtVwlex8g9s+fg5s
CugzcjIOJvfMGP5uvOG/htUBS2oodHaaYhNU7nvexeWGjKlsLtWGQRlvZRtq9VkV
XsrUpxEkM57IAN4DYnNSZPcBL4iv/A3bcxMBtjxAm870/BdBEQvAr8G4zROp2KUC
GcltpTq6/ctXcp75mLyzccglesPmtT9JIAgIO/WsWZ6UdMz+lhRa1g8Gr65bDWbQ
LvINeugh39iKh/1H3J5iRka1r+2im+l+5XgIVBtYQXDNW+n+D9qt3U+iVN6Ypevr
cmgWs24nzTvhl6OlYitRTX4343VJxxrcn2fUnij1AkEl0gzeQXkv7TQZu+3HfWOL
xhSzp1GyMC2ripNJ8SNfrhcsnpBSe9MBCM3OWJi+Afce4LYKQCfjFQVSuBTICSIQ
6CDteTGFzhz4HngURVDMIBs5Dx0pgMr3ghQwOD4/hhfoo3WCePWdlH1W7nHLAcPu
EwPsaqzAaeRPRPcpFqFsMNoSVrRpMjsceprjI3WpCjnytbUxqXeKGqwFyiyJDWqm
gy+n+/6Gh3rA9l8GxNGYUrucEKKMmjbGccwRZRFcbuVGuq4pNtmRyC736eTneMys
x79S6+j+0shly38BZSAOHATwwsnmEpeEgyFA+Fx8g1uu5/ju9IWKUomezErP2KEO
mg3ceS3rpCXSojJWz+HnUHFSl6Nu9TmhkRqHZbVHqnIUEtLX1BLDS9YOMYsU0I4Q
c1cegLiYqx4TqKc1aZX15ya8ZqCZ5y/b1oFqvuo4mrZkiZ2RxD0oEBimQGah9KZk
P5ljKhGTs1++7gG+q9pTT2QJvLO5IFDxvKJu5KSnDM6g5ZT5EY6T3XOGSIXpf7i3
yXqgLdgIwsTNWWQwB3GCXtxPsWoqmA4F5G7K4LiZvhjTxhYKVIutNXUd2qqziamL
3jfxM/hn+nRQl530EHBOxNENbYwzwTP3wxoSOobV9/WDYMjFaXiJewC05VtgZFGG
uh/H+RIwpFkOCeIG10ZgkLKWQk71vnTQ6VYgSgfgfxvs5Cl8vjvJwHkvm0AA4FEF
oKmHJICeEnAkiurAV1crNgWeSGAhFK8kgr5280/LwWf+8XlEQrIoj8krr5eXH3jz
AWR9v7wi9JSdlE+5RXo6kCCL+WO67V79DIe7/yNu+w4E0Ae76nClTRLfrgPIuHLR
dKUTE2BIbFuiq3R3Siu57Ju2qqFp9OXL0jJtOlKnwM5dEOfPjT5ElDDHuBfTJoOp
tL6fM7WFT9tri28MgCPQhtHrAtoLh3/i1MupyilQQih8LZj0WH1Nk1It+XxRXMOP
/tmTYlxucR4d7AhDKo8tVjkXUhPjWkQps/carK+1ozVz95evEpchGbJ+68dCeNXP
6GlsbShyszYu2N3XSIlzZMlQr/0d0APZQ0VcbytuQflaTllWmEGCOTQyHOXP3pa2
oi81Sfh6QFhHBWwg5RFw+kDhcrOxkQxFQL7j7Duq1UJ7hzQfNTC6vmO2JpoHngtW
FnzMIKUZjvskK3ZMXE6BZf5LwG5Ghety3iTVssYr1CA1bM6a4Iw1Z0z0D3NdYu8Q
lp5pVqiZd5f878Nkh9wiaSQvzdQtYbGVerylfuOnrHbp8WpvxuE72NQ1tWT+6aVx
bcQOBWLyg6YwbSa1CpCFnBtbN3Oncog3ganHLcAGG3+/4cb1E1AOO+8gHW4UPIKa
JrH08dWs07Q3Ten6/WOsW3WmVeHJxB5ZmK43qesb2VPdxaXnhX9j6HUQpCj7w6sU
2TzdPNLEljtV+uA+3y3YAbQoGsI2DMLsFw3+9zXdViiDRYEPp6kA6wMOzjsTwwgl
Rc22MoQlB/mXeCyQRtYd7guWRrInAThDopoV6noNay9vnOVrHLqlMqh/diIinTmb
rkeBogVYHYTck7GaRfY0r28PbzXoVds/jOhvDywZGrIKOR2095X/BSXEoTfAx02p
pIu1IKFeNnfCgXwbK/9jsOUcI9XQjat02Q9IgjF7vKNOYDST2lYgCYyF4koWD8Hq
DzoZU1Na+aimhhVf25rXQpRaZ7XVyGfVOdmAs54/3SQLKRe3BZMT0oBRpIs/Zogm
lM8YyPfcr7sLIg66Fb2PGxY7oFG99tArB4f0fNdAtgvm4U3IMjIcJf4Zsh6Sl3+D
eqDBGntxQ4i2t+gXzRLhyBAL9ZDdqnteVboUJAo91g+NcyF2wW418SebBrSCydkd
BsJ3cFz+ctJoO8HOnSFz05AQC0LnnJOOC9EERhmRADnBHnXaNvLdkdb7ljkQZn0c
q3PPFWYiruc4OIyt2R4WZJGvjqtWKj7iTu5OdBb68BXKZ9UkvJwrzjsWz2UpcSVY
AgIa+dcnkblNxqdKlyudUsCfycCuXGBA692+Svs6NQbPuRe7zpXE5a2zaa5APWz1
DwZtaH15yRyJUgMQ0Ckp12HXeeFvdnCzOLPuCDdkIOkN4a0DpaLeRu0CbgRF4a++
SrT0JpxlD+BOaRz37QqZhnulgAvC6Gk1H0D/nwh+gjkef3RRCf5rBXkBBmSOEhtD
JI7GO4nHhDZ5qlTuV4HrAAIMNv+2wPVEC0b30q5lFSzhkGA9VzpNXiVnR9SmYZ0m
EHGAGcl3E+hLWHFSSyyLtSzVpjWjMovYuw0d8D7T6x4XD9PB/eWgqfwentK+sxsE
lkSnZx5NG6856adCI1A3OKhq6TP3wDzu0c5IRviRzQihym1v73zzl5Ka9qOTPlJA
mYPbA8O1ne2ews26vRsxDKtNZbLIBHpVrKqW8qqfCSV9VO56OFtc+UlN/uMvVZfD
uFwkPKxCPxp1WcZHOnMNp6zpjud/lT0x3JRI31xR5biTNtTH1roOJL+s7jD51OzY
ZO2D463zrrKO2szXAUeB6ahpXR3tmBzemG0UxhwU92TzML/kjfq2PDMLkCQeHMLL
E4QEgZXwCtnyf3d/pwgHdlKwig/rJLaEmN++JjT86VaMD99XFckETAvOMZTzyXlm
fAZt8PfxE4B7FnLwEVND2jysDHIdCX9QrByvpmNfGjGSEyzoCfzehCU/S1OGdoOc
L82g49FIwK7Gb4ewKroWVuO2eeGpu0kTjrlvH5nNlfTTUBUOmVIfTWsNLB7GlPFf
F5m4sQnsr9QkPFSsbZ1QTYtMp/x531aE8aSMMsbdc6a/0J1i9sK78lfiUahfa9cm
uZCGNR7jFaqTsDVvw2xelbnMt4rYQiodw/2VY+IG6AQs2PuZe3emDlhF+oibOas7
UHDODWOL840tvt3NZLT/HRjbj4Z6vVaZLRPo7bOyYVsZDEq2lZQCRWsL5/YcxoJb
E1jtOwpZSWHwvD1nrw1vkdHErWYQLWXjOgIjT0U8zcR7aFpWDd0iYSTHX1yizmO9
qAzAA/TEl0iHTNMZfhS8IlsWrA7Fbhr7xRCmBZOdWgCYDaqh353irLg2i7c+K6Jd
yN8+1l/fM/wgUffMYnIg07oN6f8A80uTys0l2WuGI6FhJUc1rHsxuHq9WV65AeTx
Bq2SI/RDK14KJFBLNJYX4dK0OtkxfFFjaQv40CYMHgyluRQaaotytZ8pLo+vIMS+
3UqwWTiD35NOj+3UoqpCIOj2JHBq5W4Ju7WdXCoxB0+kA5p3D/eToGEZs1Hem1pI
qqNPjQmg/BaCk6VjkrdS9/byrVJtDbHj4/omYKSz3+60Gtj3p9rNlM1090ri5rqs
6S3sHQFsEuZWQjnd5lkXdl5I0q+uJBG0nIuKTtNioRb6D12pOEefs04mjOaLxbHT
nfSIwEYkOcir7xX9bkR+fF4QQ6meyTnT1ls/eXjEPlVIv7ZQQVrlVVX3QH0KHyMp
VXJV47BoPZgMeey5dZIc5J8ogFieocCgaz81DZqXkwlyX9nqJyQ6mnoubxOajhu9
7eZyRNYOVkw37g9GtjjLryFU5yjQVjBfmlpZCRHZ5/FlJQ5wVDevXInECmhhCrpD
GrNw5Qe9ewWruuyK9Um3mzYX1o0gBptt3xWk1kGF28QkTwmACk77UQxmqx/Tp6eH
no0G5h77V70WDKiwF/RznjK9gBL5sRHrt/iO0CU3vTBKq2cFqYqo6VrwJeK1bN+A
t9vA4gkfdU82ohW9FNYjp2xEAkaUG7hXyqmmNtrPvf6mzPp+6G+5cbqsT22NQxc3
zSso9nwW2cn53CqiV/n1Zx0ptZZD3o6HjELCjq6J6V4hNc1NNjl4Vc82Vc4ebZNr
Zh0SI1YZZVew+zao+XkWNlaEOKGVH4qaQPYpA5rvcKpDtmpYlNojKa126nXoq/MS
t8+jEPJ7n4xBlNN4d2Mu3AcBaZxe0BEbGAqaH52C6dp4i1+m3nty4dNZHIN3qp7o
awQII6LrnjCKdDGWlDF87/MCEABBcl7t2HFJmDsSJUWWCvr7RHvAtyJyBWwMJKCM
PE2LXVfyr2sz2RC2b/af4vVZXjWpNWuwTdSbKegfOgSEUSQz3CcWm5oOPge5lgMx
4lV+1Vxp1cw7UJJNe5I0i/w9vMr/ZMKPw4zlJepmn+MowWQpy4o3fgfGXvjl8yUs
v4W1ZU1aol5A6NSLlqBE9ls2y4IvdJQDf1Yf6v9CB8wN78kYxwrb5ufCfKbkSD/8
NKXDpflFHxIoz0owS0pJ5BX5h0uLTCyfHifQYWNbLEQI4bnekGcR5POmxST8tKXy
qr5GWOlXPR16PYLsr3NSKC//bY2E4KtnvMfwYItqzYcVrDi1akqZGgX6EeLopzM9
IwpzztYvh2SgrqmndvLzT5gcE6q7y9PUpRaNR3b2v3Xd8a3bCGXQ9sFSLDYtwsiL
bnpc/VsLlAt09b1X5GKbxyQSvtSrUbq4IWq2QRM0jZ9aaPKoYOnn05+druU9YbuY
2ISQvo4ETN8E1O90zde68pxdBQc81ymh3vYVe0KtiChxXA356Cdp6vNqjWVW+1no
lJY/demZWtR6RCHF328A8zW9P1x4t9VEPo+X2OX2+OWeafVQ4GRtUvQVAUQ6MSgW
mH8YOdNB3BgUhnYQRGoGquvjLjHV+xZBUxWWXW29qtskew3nrg6J0VedVMQM1/Zv
YRLjasqQoWl5JWTpCjrGbH6dksMGuuC7JossdWv3HiQqkeQo4E8h/mSIO/taToLR
GCu8M/oa/isQ1EfO6Z89Y/yO22YoY/BsHsEOAhnuXtkJYVFFAO2MqtpFc4oGFu20
OvBodX2Z+tC64YirEYoM7qGHu05s6pnSZ7WCCp6xq4ZgNG+xNWT5kibRkszwtpym
POGZJdAVsvrzxrxPvvmhfIY9nbFY0UctchFbJJDO+QP86uz9kG9MT/VTl8cNkLDF
2gj/+YRzV1VpD30D9SvmTBZeCLM955hrgopJ7BE2yx2i5pNhZ4JMLUAFyjwTqaB8
heZ6GnS1zYdv/LOyEjf1EDxhRmn1Kj0TrmO/7gBZZT3eeq02EMn/mAy3dAtuPgSs
dX/4ZUeeovbNuCRiixDThJ9/gJiaLeEHnbDRlLflmvUpnr4ByqNdMKCPhyiGtMPJ
TJO6zygEPqrW0/eVRkyOIsQ93DnH4L3jfoT7WfnFRZuWsqOufDXBriPCTTDWw6ra
anrSCuP3r5DjZjBU8uTWHJvcuK9C74h4KYXE4oCxRsLQias9ITsMxeb4i4lDw23x
nz3+pT9PoFzt8qO9S7GoFk6vCGTDH7NleotJ20JEkKzgYfbo4r8/nH7pnxVN0NiM
ifiWWH+YwJq47+Pj6lUWFMrGizJghoVrFjBQUdKw1L48GKTcGm84RDKPs5Qhd0UX
DAW7CW5iw70GD/OQBYwZBqjxIcQ4fb7QI3xs08bDtRibxoWSFdVpCJd8+hzJSJ0S
gP46d5aZ2RQHSlnoifR0wvR0MeXKmESl4Z+wlUX96wGXmkVhrFOX1dN96n4O1FhC
kItk5Lch6sC9tzoOXzDsyH092nf0VZfg//vnUThchrAibu0k3wdcpgr5iyJfvKXD
NjckurirxBpszT7cAFDJR49vnhMnFlBCuZiWZNvybAk74slXXqSwtNZ9wefK+una
SwbStQ81lHalaaZzSmXwnqClQ4BVPfK/SVejFOtUrx2TlPGv8P7NoTcrnWmEAq5K
fJbFDQG7EFPEdV+2T8lpEqQVyKQSQYdZSTAEAg55UKfUbmgwkgIMS9VmcLzudns1
kLrBnCb2mtjdEW0LaiOXM4t7j1oc8m3GsQKWSlfNYQscai25yiSM+e5OX+en4ALO
3dhGvwL2pAE+q3YUPrLvzD5TS0HK3oWMdFSBo2IVOf0YO9M6cVLrX+h4Y7BRLN5P
zbDSQIYYMDUYPoEcbbc/nGYZDEar+wgxjASmq0pRRexHXIAcq9tc9nCpqTUz+YAz
lHUGXLFOUM5zIN0oL5qULYG7OMMQAQovaB9BW64ybcYUafqkXp7tcWDxY8zBPUmo
BSsVbu7Bz5if6AWQ7/d6rmX0igvl71yjDoX5tz29XBKe+lOC9qKEK5RTJ96lboPV
IoQJ3FLRatUgwkAk7TwCs2+gu9OD+IxRcGi341Jxg4EuxtH3fiGcBEaXqaNvUxUd
Pmu57t1ef0At09IbcX1dKDpBbwbwdK2z+anKDQZ7RxtN2kCrTmzJ0r4NMlttYEQL
KdTwltIfSyR3GuOOTU+V/tdoGN4NG5cT+GJhx4oYNcQQfxB8N6ve0fYDNWUU+g/k
mLPMLhk4+yanrnNQ8Qio0N6wNSrxk29Z/guWAeoJSNlul82KAGssOdJCsxJk/oYe
IIgxWJJRxGaZsnyHuHnaEzvrZAJ9Jo+VARJXI11pnN9WXpDkzshZ+Qw6EG6A8Zi1
/ZsOCBpivisqo+a/AD4rJOJBdTDEwLj5dmA7Huk54j9lkyjdO7enO24mTT3KsQhG
lRkGri6O5cCd9YeNuzoQk/+fcDH7qQqYu4HfDKLO0x/wD7vVCxEjiQl9PYP8nuQE
Lz1Kw1VF3NckzpfaHaANc/cDK9uafYjzO4Ev/0Jrib6BnF7/cLyT4e/lQiMw6pvp
I3+UHlqDc5BJOthHvGxar9A7wjB+zTHsu8IKWA1VpV7M0i8WArD0fcA0nyH5Vj/5
lRxiJTvSitc3r9ZeoCOhx4TWxpidYP7zwfdLlgdq8LN0FQ+V+t2BjOOiA4QLzOUs
Suz78WgpzPdvwYrUDpWtXdf1LE4Oyc1ChilBRPYsEFOYMdmHF6HBjb80cfXag8MO
k50rddjEKyJsjFERdjK1WqwlR+DUVtRhEqqiyCMSF8LSHqhlItFXqWQPMfputlex
JH3ziGlb01MMpCi/Lm9UnFjK18rY0Bg4W2eKtMquM8+vjuamdLG0zc76SnvuSRV4
Cz9PtjOVVO6MKo0byN64n6M8hothvtctcHHrYqv8ddw4ZNDEJdpTC0BoOvum4lOh
HFa6dgOzRZ0h5o06MD0jlqNJTHCeNT1TrebdCtn7t1hNMxHsOsgLF5V2D+n28Fe2
3+u/snNA+T/HxY6I7PGmNurzKyn7xOyKGn3FoRNzhq6tq3hdG0ZxKGsHmfBvt1HY
DiEcKSNxILtij2d0UKd6DFXCS2IQANY+xKsJHRGWQfASYxjmG+9BsFGcStZMNWzl
1rWv07r0dHZVeDtJFV1ZxC722HdVmTJ1tJ9k1owUsjim7ct1F0w+S/71qnZuXUdn
usW//JD7ikt3It942AMX2xlK0DDKU0hmaE8LzQeDg4CLAiNX2gOIoP4/TGljzxST
tyCM6rVHWmOnk1LkYdEVllOprc2Yp81EIrsQ4Woaj6cM8AaYDlGIBltf7/zW4XjI
HelI36naD2d1Iym9F8wzmv6RlgNQ/gJZFNYjD75Unf7yrqyLvFFkK39Cheib+cw9
5ycdtcBD6p7pgNiZuMkyrwBG5lqOGC518S0wl2Kd7G8TBwMshEzjoT/b/QMNHs0M
stZ1C7jDxEESmpC+CTPWVDWo53A5MIGiVvss/ny1v4n2rJO+HSVpJPMrWy3c0W8U
TrkKQgQp3B6oq3TZqhRNDhpTWYdixQhkLOQrrzAtqsicvy9mxCRkDPEV2+vW/kqH
IWO+fsGcU08jYQJhvHk5EoDzM5pxeUTtPX9hEMRNt92cFd6u0MC6BMejEApN3Y+N
EAJ0qewFQrhmHtip3rCJrOpli3APTo1PauirmxkhdchIj3HNYaZnP14ZqA3FaULV
V/v4XB0HjOybeuabNjiPGcqCpwd4ghBGU9CLeC9x66uv5newQuGstwQFPe+3Gp2n
WpLZvTT7t0KVjEeddgDruR0EdESmY4TcPJOmNSr9TsW7q2y/yCbP+dukid9eRZe4
J90yjzNf217gJGkQwbiN44eWyJ3FY4+v8mQoBSPjn3+e7H8hxz/CCYW0X0YBIEza
v6i+pxEadWhIiJO5cNdGg+NYQZ5KrA/fReuhk8zOyoeMGJynBEBum1+MQkAf79o5
bEL7fYxJENC+RTK48yuFhst+1ABzbxVkS2Qj/OfoWLEYSoPR0KuaJ9n2W373+1Nb
lc4IPlqBFswkm9tuQu2L6vQjv3Cc+8xdci7MG/17b/asAxdPMreDl3G9XZU6pJst
nai4JS0gN7b6iBEY1GgyukFY//IWcOEys11v8qbxp2vpjk24AtJVlIibX2VOpKiy
MJYXs7V830sN2gdpBv3IrnRFQEoB54isOs+v8C4R035s0TeDLPjcHBtDkayT6S/M
5uWr6EZJ2ZGk0HDmVQMGBSopHbsAIZa24tgC1+/hx99ScVMa+jFTtD7E/ekDvxx7
KCN8YbBGJ6SbswSwtoatYWlv5IqtJ1byd1+42ZyNxCriD0X9DVG/zcpWI3Ux1OBh
41wK23hvn0oFmQEBZchyyXwB0BPHe/aCQUY/Rif0lU3Yaju55L/2GGXzjX1/yx2O
vA2S7lYK02nWXSxVi8sU5gRcYMiHZ67TbKOeqB7/UCOr+yBU5MynRkd+lyM0gsTE
yMVmsyjW4bunPb1z5eCLZzCD4DwnlyozukLlYmra0PyDiMoefSyOXxAIsXo7H1a+
Qaz0+mbyfiZ5mtdvNzOKRYMxHzMq7Bd5Rjkh+JECRC5IwQ48P4GERHqR/Teftfc6
bBO090CdbCg4ttbCTBWLtPMPcXQBL3OOfVEGD8wrQvoWFE83pHqLhZcw97pS3uz9
jbCW+h35nFwaZUABQAzhTmN6rEvNhmyqX+7FbJ6UtbGMXqulgck2rdk715dLn2ac
61fvlKZ67e5XREzm9PkAzcf6ybNel/tt203S6s2kgUszDKe5qi+YA9juVRaTG/bD
DQ+d3is+FTzz9ZBvjim22eN36PqlDNCfSX7kODEpni+P0gdskH2UYWr9a7D5G9wF
6TAQAXGWhCL9ORn5kGLPPMbY2krxnUOHBjcjrv8NtZb7RYDY21RagfGRB9TyvQS9
ezRAvXy6MbDFu5t0dcNYiHMfp3Aw3V5RXmqo9OAcW8Y8Ca9Bryt1czGA0a8UK2z+
Tuyh/7BLLOR6KEv0ryS+YTrL6khSGMiGrkMRxWj9dWT4pYy+LxFyWUff3y+vQu0C
nz5nWVGtrBE/+lOkrxVjqJbN/VE7G6cDND+9r6kZnXQXs3bSq0qfGvdy67TR95q+
/ulXRRnLVrNY5CkV3fj4m9QMEe/BO4HVZr1fpdO5/yNm7yuad3FNtX4kejiNHFQl
9k3bFeHpD2YpTJ00m8tCsBiWF6NFkwqCSzj3XUdbtcMU10IvbXFng5qsfKvyqcdL
O4umqzQRDJEeNPpq8cmHei3B1TYQ+tkslRZVsemqr8ydSG2etQ3MWdE0VUWhYZli
KL6/IBNcZvynAHy6VQn8j5747TNRl0zSkKYMoe94FzmxAbiIn3KzzwuH7AOAQepr
jidSW6Uf6y+I55v+0rlUPpzlX8ryCoFmOu801G3Kp9dLMxx7Ytb9Xk6EJ8BN13na
ayvujMCNiwCvmgt0342dtc4g0mkQMc923iezBKFaY51+Fv0XxOLr/t3tRDgMIc9S
5jetySRFSr/p5MEhw/kc//+EpVv9+isFZhBdRauDehWGRYFaaziMmEfqNRe5V1g/
+3SnH8WDinmw/Z6RQgXrK6wzwea/vWtvTeq5eXKCJ39KtKUsi2lir+WRa1RpEz2J
wB2gQmOVAwioGOBpHx/HaBNST9tf4Sv7NKeyn69HJMIP+CR4dgwTGQInfEeUIJGB
YAhKWT9TN1D61cv1C7q96uaBnNqGaXwND/w5FbTKw24kDyF3XSFz1ZgfzvcDTvdo
LA9w7eXflOorlZyRyuEq5DKAh4HhCNOG79c1QW386PH3BEMrwI7aJ2wtvUAznKeU
MkHOG2ao6qvaoR7bd3oXspovMiJmynQZnEcgxI6o66K7Pp7DV4tmVjs2DFyL/PlK
R9R5dpo4YKvFVWCK1E+CuDeJKSFdNhhyg+Rso7i2lmXA4jwKITEBIVbf8aNRWn8B
PTNNekcdZJ/kxuHiS8qfnAk4pyQZQwEmrMhmanvx+mF423OejFovr3A4Gz4lNpZx
wcC2DPR71Nnxf6POLHsATXB66Czbrly2f7vTheaMypezr+Jul9ytm1R2uKN7cwsK
6lp0+b7GOZ61Z4/hJgzazj1URpgRX6jElleov405V8Xoz9vj+NWcBWo/REdCI3X1
iMSqvyvbKrE/N3GWieDIZg3fw2nrYndH9fis1zuk5Wv1Pi2APQrXldCIjuM8fvia
9i9H9zeBdar53hP2sfAkwpyQ7eYHTHW7ZrBy1Ljz0GzRadVgmyV1vitm48FbMScU
aBpuvYy1ZiORfS3TifvUXSXaJA/8wVgoco2IUZJbBdKpK0nCAOOm8cZ8u+WezR5k
SR3VOWKum+8sU3KEzWtn7SDaCPdnPbiArK7rOoipdzH4CZQjJawESo7ITg4j5ic7
rjZ32hqR0vWfstsm5A8dk7Zu5R+yqR6S5kr/hARlGLvvcxDOtqvoNma54E04s0l8
oVdzoOZYgP+wy7x0yD9dQNeZSz6+sgfwxLKo0wyvIpi3bSPkva8sP6CY6lhe/EPI
ZQlusYlaosK+rg33X2Do7SWvFPSYxXxYzQrI7Uet6Z9wHBSK7Cf1lQIsUAqrn4mq
VVg9Un0p283GRSMZQvKRBs8ytta5WoquRE6IICz3hgfrTVx1O+2uZdA1uotiLDpX
9+8SKSckQYVI1F6p9KdafPNDC0PQP2AEp96Tmh/2NDPwKDCV9u/YNYybIcOwbjnW
U9N+ny7wjaLB/qVWWZiEM7J5vxBmD6O8gWSLslMbftVvtVllpFPjQ2GZGIX4CL/T
E25svykVoXc0OtoqKgR2j1UddSIyx4Jg5ls3s/90tdoHn0KCSNahI6pPA+XdUykk
c+d/fbJf0b1Lq9KymGyaR6nkMBR9QTbzy3cNX1g0oM1pAgTsnw6Tr8zRk8CNGLdH
MlAp09JLzO8l4HcZTkBJufvL2GnGNaIa4YdeNGgb82/+0IIbqsGAjHrm4qreSpbo
6bGLsCPIiFJJwGDT6PuLK9NrHWPN7QkoAKg7vpwsQuP4+KiVLuqHPYOI1I8jw6Wj
U/Y51NEKUQB2BsxsoACA88BeS5E/IbDxiextMlzrnxQjlZ84L3HNCswwa1+FQKh0
gkM/QXbSdYk8KjH94AqXMIzF8U8jO7rGYQ5Qu+EWn3A9ShzVxWewuLy8ZybcRgf7
akFMK8vm6qyj+yHy+1MNNqsJazRh6Oy/8Hqy42KKLTosujk7lHuHf46/7+fCUq7z
1dPfSx3yCAoLF0HrEFPDhEGuBK2jrZ/Kyv67+VH4qm+KuoY1GhLFxxNE+wgF1sAd
Rc0BdMNzOW2xxmvL9lFXiNogHkOl5oMY71Ir1P+5IP322zKM1DpghnnHqsNDwom1
Q/rkW8cxVqOg2umUk09DWUz2ROapcXXHEXTiJiJ4FF1pSmOvT10VVTlJW6h2xcWK
VFx3y7aMFv6vXkNlhS+WDH4acc9yD9Svp2/S5Q8vsbCYskUVIWgL0/ax/Bwqeniz
hDhT7R/DCHwZxZiEH/SnknZNOKq/dd5qGKCc7j6NGiziPYSqqbdHUFGok21TnaU4
OwZL/ve9ZSbFG6SB/WRhNqhWStl2NmTL2MQ39hlXPXWNgkx+3T1BYTmV4KjKOrYH
c5JWficN+/tgBN3n82U0R3uFhhLPKLQPwOs7iN+Lh+BngRmjTfScJXTg48rK1uRH
1I27DfwCbu3pqKDMoSV7gxPy8cSC/qPZmpnLfME0eKOSBVYsUMV0e5zpZQMx8xsp
qKoMYDwd5bmRGon9GxfgloqSdNjCgSjBRBcH78wbUDmkUbtVfAtiwNXP3VSDbQeb
milTZwuzftFlF3koA2Fd7mSzI5mSZ3v2LVbpMzqnqK/St01pjsiTDl4UfBKnwQUV
Ge6qfbVeDiYt+AOvjmUidFgd0VnJ9/7DbXCrID1lzbQRIv908Eo5UueD8dcW3Pt6
snXkFBPd1HfcIhZPQRW6J0OgoOc10i1iy9U3Byp6py9NvdGR+rDsnyvvHG18je0o
iRvmUVC73v5UiX4JQL3o8+ewLfF9m1J3edP8YiOf0WAN1vZ3ldnKAWYhJ5V8rUro
VhBdr1RGQluOQaSox2YWZaxoEGuJp+HQAEynGUezbI3uPH+M3VsNDxRWr7e1opx2
IaWZ5Y4oilZ+hhRMDoStzmUePFRz7nWoSCdWr8YygtxS8uNYag+5RGg3e7j7c9sf
vmQcjU4dZYSUfrgSW1WLfg/qbGbPUWrxMHaYumpQf314VeLQK2ZAhVHRVYfq3HoA
j0TYMtmzujYYJ1YN5e6g+d6j1TYU3ZhLFLrNeE1IHOrVrxciKo3o4UAwGhcBYw/K
QwrDAdOSBEFalEl6q9hxn3jLsYXxJzm+Cg4nlZ99kRwJqDFkqkKO544uEQMoIp7Y
6MqBl5HPhABp2mU3q0HUkYpfKvn/+NQwSvjLSdzr3eDT8yeCGbQrvH8jPpDmOFOU
i2r3ZxyIlS3BxZgQvDOUh6lqy95+EsPifCucvZsgOO0ZL0uXUTq687m2VDJcFHpE
7DOEbDic0sudB6eC5ceeP2uximZ7SwnXOqhQW0wRNw6hgKL5ZYGlMMc07SOUnm4A
l3lMZ5N8vA9wuhmCs/w3G86hRD2min3E+3h2M8zgIe/oXW6eE1rp5YpC/ITR81il
BBtSwASGisMOSNfn+xW/huDjisnOZL5pCVODCghpgwXFqT88OAowPRP/HZAuzY6J
cAKRyq7XiS9u6iXnxToMKP8jfh9q87TUIFeY5UcTKa6PeNsM+vlg+KCRXHQNR27a
pxru2xjdQcdhzf9FviB1uVlYsJY4mQ/d4i4Qogz0tKWGfz7wdS2FGGvQbmOKeBGi
ZQWGoxfIjAGVur0mMg6YqV46jeRAdNai9t9j3itkGVGVuifg0036czW8DT3qwkKN
cpofdOqpjsn6xO7qSBP825XLL6ZxbsnyFqU4O1AfLYNMZLWOe/lMJNf41OQTu0DV
UuYlGL76qU2XEA/9Prgf0FacHNi4C+VfKBFDwNT8oFo5tzZE00Tg+BMOLCcLMyup
H10lSyBvkIzjeHEn8urs9xy+HAgDdmTLkhphQXzw81zAVD4bmgp+hW/kdZIbiklc
tzNSiT80iIFbhMz1rDSDR3cPaygWHddAxwycw4Lfwf6bUVltKMKMAp5zDLKvb87s
5dTkIBhFtOoOwNZiIr3atTB1ld+F8q3t71pSeVvVKLVAbIX+YAronhJuP2eBXCUY
j41c0pac5knuRHS2oR6qPHJIyvseMW/50jwcM1cC66ZfVnzUBQxWxNZHAhPIa5Mg
jqaMcnH4/0cChTBhyuP/ghYSGBiAMYtvd3KaXHlBNImZJa3YTBJmzX6wIqPYQHZh
XIPLIyS8Y3YNdFNGrxhYAPqAnBChcNqhuut597ZHxMuVv9c7/Dwo2otY4TAgkMJP
dtFYXL8krXC6I6eLxpc06+ZBs3TOt1L4zxEt76RLHX7ddLKbiPm3O8jW6EJXPLO3
hKZaF3aZ9E5p9WgcjirGmbwTQZkOsa7EZir1sjdkUz+MbSSUN11eZphHPeeGzK0+
vVKFWUyY1Goe15FKuRPG3JdwDn8exEETJZe+YNoDV6IEh483EAtZrDgavtSXmYlN
zUO2yqeJ17gQQJ2FOwa2urSHSH47Ma8PeOJI9kw+hUYa666/OsWPv3c1a8clwAqs
bsMkAZCPvP/IGfbm0cwfrAx83m+0xyESJoDfMRrJdGz4axWsg+oZ7dW9g4wEuJD8
DHh0keM2W616sBKhxM66ZwhxT0PjBy894yG3cSPgKbY40zNwvO36z2ZjNfhvG2Yj
ItLqNPBM7bsbk6n7+O/xfWsVACr3wqwpCigV81KfLMGpwTDnZf1T+giKv+a8q31y
hm3oj4FP8rOqVkt+fJkbDUMXJna9ml1qHAug75shkkDteflxC/daGtUPKX8JVlA0
adAZoA+K5gniJBAyBybAwID4BvXWi9zsn2TESc4/J8BWUyumVOyWNW+EEgbbVjq/
gdkhyvU9pms7hYBASAyieRru05LGOXaxDfE8E49M/aZ/3s9kk5DVs0wULUDFeaAz
kEha+oM6M81ku0ArWwfb2RVDevCAD4iF1DcgPHK0wB8XVM7eogaqD14or+iMNsTk
G8CYK9wvpeV13mVRCReM9vezYPRA1nd4IXowNCXZ2LxFaucSRrprJ75WVMbMB8Ka
w3GPot6/hWyP3SFGrc2OhJRLxFwXHaNYWBNkAqsZzvSfEHruMfvTf6DEoOnfTrbj
PwuxSvzofKAoeDgwal6+xvbCHCFmH5SQzFfVjEPb4tzn2UZ066Q+RpSI4QwAtA+D
YkycYrO1P6tpMBoovdvRUaSFrB5hdo3xqvwavMtzZr/g1TwOHaD2ARqGndZW6qBt
LAwB+cRdJe/chqgeFJBiVpGbrN+XeWX0myIKP33IKA11kHSr+LKNG9Tl9dEBABuO
4c46kDBm9u1K5ue867cO5eEYZ7+siSZ5sI3BBSyG2l1ANDhGTel3uSLIlGeRU9vQ
St/1202oVW7dzRCPRlLCY/TVS58fLJLzwM5BBZ+o6c2jmz27a8JdEHrgiRNx4UuB
HF6yv/H6fh3oh3apIGd24GTi5JgoztsIUParMmNi8XSC7sFRu1HY3gH5OY9jWM5A
7UkqXlU2RtGAte+C1ovhklc+gR4o9e4QlVUQIzWlad6KOjzVBmW510Uw96ZqJpV5
YzLifpfTOaZkPnG3kaebwzk1TD8ryC4T0AtyWjg/XRgAPCH8GlQepYRcew+x8FxJ
7NRXx8JYL3cqip9w8whWbKaKZ8REDccQawQAefTCmh8pZSZs8BhYb3eSPRgipOR3
FTe7ueJFeXr4cZ6koqEyzO4Gns9+J51gcVjCA/6RZcX8q/DquuomZYgRpHi7i23L
NxSf9WECpa05tvqxMFSqhyGlu7eTXB6/mdcgKGShLqODw7X6UjRoB38CWzV7bK8U
ihT0vEgYzrVgVFnaGTvJNvWfRbFE4Ej8eoXDPAyF1Bm0hUHt3JHxFyPMynt70SjE
xzVubjeV3gHkJ7suD23lGx4tKm+GMvhn18+vIUEz2v7yoSdgR4x3luN0jvV3whFA
TmTudKieBCeYZgi27pL4hDaM+Xe6UbXFY8Qvqvd8uQFL4m6+tWByLJqpzUs7ONO1
PYIrBD6eYLkAIqXUwiKPLtkSIe+fkINDeoo5h14eGwpVH097dSdDmiMCJAGjVZoY
5dFLKc92qgpXyXPuU7vHj8O+7O7fR2aBbVRD2I1WAORy5EgUOfVkrWxdvUzWb0rY
qD5jiS5MHMxWgV5P3BZcW3TBOGxKM50Gpy+w98PjHbVPvBawO6OqnsO8YhRzAUBL
fVSrHsLAnbj5tEXSzlgA5ZljoNzFW8pKwNSEIT3O7IJ7Ud7CatBdKo9eRZPW289L
TrlK2rY3aGI4PRkGI8AyPy7YqWuypwRkeK56AxX85rjd3tLP0cADQbUqFP5G8Zu7
l5EmXxADNSiZQuwCak7ixFRu40kWYtrba92DizG7IMg01XOoG8Ty047YK9HtrSmA
x45FJjkUy9Mf10ujcxyHyILBLK3j0AtkxjWdSKDSVZ4ojT11DIHb176DjxWEqfT8
nKgb5qHPYQL6GcQETQUEpCzhsTu+zZrJnpk3CSnDwRg6kJ1MkDVc4fxUHhcwOR1A
DdcfFGe10sXb9B9kHRvD+ajFqZx1h3uaBUZ33a9HhC/0d9vCoKghbFBWZOlpZR8A
eQy7tSFMfkk98hcL1xz6he/WLbCSF0dLSDlYFdRQhxxpypZ0fwBTc/gjgi3DF2C2
aZ+lBBOKQIn+arAuD+TWqmFkjZJCYPFcgIJm+JPNvll1EL+a3gUGbyjV8lxfeZwO
7M2KboPQaIW1+YNj13RqFwKWhIjMxKgOeQnniraxnYKkhs8K+l+sOgNLUanS/HI4
XreLa+eQVZWOLKckA+jYHLaLXxIOUX5HPWu2KfGsBhSD2npWbjfadxO6us1PrRyO
2Dj+g7y7s3YFq+TdHC9BlGqDwWiUWWGmdhXlp2sTEuxFU+Q32bkBFYSuaXHadigj
KJdB33dblsWaArUuSyCdhl/iJjg5X+dCIhcEbMB4BpKHUS9PXAtBF/EcoqHuG8hZ
eqzHXlHibLvnjskQShPpiMo8g3sOATfPufMoGrL1oH43c8AvEqU0Rx4Ib/JFOSx6
ydaa2iokDFp7fNCvuJwDxkTEJVehqgRs4DgMKj/d3pKNGhHJCwYqaIrKDD3qymhp
NBOJ9xi6d96gCN1fJYsoiGl5RxuYggLVOmG8xzyxEC3qspe2ZEpKtxaFat6LoX8R
0E9EJsn8QLVbyykpm25Skw7GVvIs26ovEsUG/P8v4dzWyaHOnOhfSwAdEbhBOJLF
AtSX/8/phkDUgU8oQZaWfPHZZeDDIPwkNQuYmatcpNeuZtuEXVn7oVQO6bXmh7ho
eTKjVTGsNhuqEoUZyrhLnJr2hlwXru0pp6SM8juwcIaRS64QlRiUUOvOX0OSP3H+
Xl/oGbeaJn+92hyw2vWhyG3qnhCrnl3EMGHDPfeOh/JtWOvtwseQnWfoafcO7ED4
Lr1i6+dSkmLZGFp8al39JtYKH/iOaiz9vlxrOj5oNqPc/kdMWOh0cf8C90Plbxgq
6LW0oAzprmOsC7Ka5Tz6wMhjJwfeNgbIG+76jiyb5/4Zh3D4L38CKrEz+w72i18N
JK47CB3xIsYRhH+6tEvPdbftsrmu/LGSpPDn4sf5llM/NB3b0+LpFmhzQ5xU6oDb
q0+SAHz/FO0M/5G56jKu5tjxgbElbyDv0BqzPAVEUR1VmOaQUNRbhJYZZ3c+WG4B
PGPhcUZ3ToaOjVEHTfoY0+Gz7hl19AZGaiY1aa3A4udjHbljZAa/8oDeBS2T5W73
dkQKRuiFoWSUdoY5eIH6QMxvapQP1DDRfmMeJ3UOQIUrGmkjk9Y9Pimygjn91YQo
MShVqQJ7FIlVArh5tdp979JHAXHLun1chAKPSuhUK+bOCYdzVNKrGZPIXiGZsKrV
UrHmBI3Yu5pprdzkjFsrzbXFGMS4IoUYBglg7aFbvw4t9MgOAutcaW6PgAaVNOq+
cj9CpSJG+fJrRSQpeAOwUvyxGJEfmC1yER4FPBbG7+e8cK21oBJJLxFDpZaLigzL
rsrcTFOFly/XE0e2X1NeWiO3CsBlaNsdVykvQ6zyuirBaI8OtDvVi21txzALTAoW
XacMVC8PUrAf0sHfKWgTMnaOKMKwuwKlNeGQhV8V8pwNFndgFK9yRZ+zTiFuf5ct
S8Sqn0CpYIn3UQ3hkqHnokbJVT3k3LGN8XW658FNTKEk5kbqlrO6pw783kVi5KF1
Mni5e41E105G0wwtXBB1mKSqD2NCADiEPsV4R1lnokH4JIbqfTnuEm19kg3yXny4
c+uNp/rerHkxSMvQW7aebGrYWB1ggOnEigAUYSWXM304+JEhs/66HoAWkfv9/7gD
qbTMrQjcxDkc+JUikIdnD+jSReP8JQq8k0bCnm9ZX3wH+sZc1I4cXLLmfI7BnlNG
6sk06Jw5QDEwvcovN4YVaYKwTjlSFkpzPlmCMmBJCECUfZ45FRgOQVpDvxVsh7d/
CR6l1+axpo+2VIOhiH8LW3LDfVz2rww1b32m9vg63dhwMAKH5g2Cohy3oBBiL4zo
Rv8t9ARYgRdO0l9v9unlVLSCrhhEDZHH8Lswi5bIJiFv5pm9n3o5DqFZxzaFy6e2
+pLpL7vlxVNNEESLOzeaEW5HtcZ3u+rshED5IBL/r74unm4ZaUWCmKbpqPJslpjv
rGZTzPNjpZHEcN+GScsnLbuhBOYfr5sa3BrDAHVaKk4TMdvbhlNdvfZApPC0kNL2
zfYOGBW0jxUZa57hs8kk4G2YzYedatyIwBwZjY0gm6D8wrxuPymHcgW6iD+9/wNf
LcvImcxrURqBjs2bCzIl5M0F+OJdOOK+zwE8WhJ7anYxjOVffBhgTYBQLwFqAQeh
L+2zh2UcmwtDXuKk2tMve059/crn2hm5/gFn6cacm4gs9xHrm+GYVCJ4BN2ZHi8J
E4Xka20qog/n6DW3wkkjWhLjwg+OW5zberSiaJcnvkszd8iLS3oVxRB1JyKS+Eqw
50QUX4ep5ERTDCn79i4W7ZObXsut8bunTRxyt4DRc1xo4m3hLe8IRnM/J2eiapDp
9+NnaCf+PIFNdEFZLcrycWXggcFOHUj2Js8Yi+SsaLcitTmIGZW5lgmOMAB41WBX
Wp1GNU1URWlqSGJbPXu3lMGozQKwncLz50K9IWZFw79qnlDYmKtwVmq/YP6CiM8Q
FhC/50ncMWDSHAohSpxD6T1P8NWlItLu7+Eb9ezbZeR1Y8P7HVkHtT2cqI6pdNKb
EKi4wWTH7w1UGX0UH8C15e0RIaS1cF0ckm6/GId/evS6EsXsp9cDd+2RruhK6wX7
YIwEfGlUmA2FhER7gWfF0RYUQFKak46dBGZKI9nLr+04Qv5AKNRGF3SXuBUUg7pJ
9VNIuPof8AYDOtccB3a3kRcwag1hjcKlJv+7hBisP8BgClNreOinUouuwmEmowWt
MoKU4Mi8+EYV9co74LMfJwDvCsIsRSSnc+B6q0gS6la487eF1bGZbwadODA9K5qn
Lsfvk0PhxBITcXVO2wNdeGNox7xVNi4eafLnw/aSQY30ORfciJ37sB6S/mYReVSV
hrKwu1+SIK2X+/J8neJYUmaOxf++ehf28hsLW5cMNyake4J7SGsknA2KGMeKeBDN
VSPkzWMueLAVu41daLh8TWvun9o8Wn28g0Y1B8ceKx0EevXGBNDfobwVIVr+dGfh
D1ijoMIcFr7sFHUaCIsOu6HpPEhvGTeNuz+mDw2ndBhi/nBno0AqT/QEA6zBtJwu
OIs+9Ffc9xyif9Z/xQ2EZz1zwXF75tqAsrJgazkNuDx8cs35htgVmAWfxWURjGOh
E1jlzbwsocR9tQEij//80SqHxVRDtbKpLK+5SCY+VsYgac62VfuByvz4a/tALQwI
8uFVP6vULhby0J3gE7R2tsiOlqyQJiFL+SdcWMRVUuOp1jtUtLioU1wcFE9M62gK
0mH5WzrhAG9+9QfO3Lg04qXd//iA77H8osDYcKFv0/o7+MyDWYbOFuln3EEwq03I
9DELhHhSQxxP6uehcnXQjagbPAzz55THAXjqQT44ix2HQelkGMF+DxuJ53I6leND
PGTnzHbf/X4hXfmmxFP/hWEsMBO9Gxecz6TkNOfMvdIXOD0+JGWppsxbduxoYVua
as7lWS4r7oyhEGseA0uQqFMShqwpw2q9qZP/0K7OvkMOB7I+MOUQ+u6UsV4eorVP
d716A7ONKuxT8LKIG5KePH17tNweWwQsz904x5O7t7KEsEGBoar+xaTStk3mz6xu
RKLpzZ8WJeVFADTLfcDYkQWNCPwL8MmUt/Wrp+96C354q1SQv77nZ5rNmkwbKTjk
4TwHKJbs11R8QoOQmhD0OF6hs40wk3UMXm8Dnka8Zsemu/EWwH7+UAef+tmoK4uJ
4rC4aB3y2W9XcKYjdfgxlf1SwjRl1SHZKw7aZtrH+izhxOvB23C04fTU2w26ZRS8
wQ/EpncjTEOo+/bgGLDZ8eYNlnUOFW2u4Fquob6BUKr3dA1u3dFZtGJAhsy1GXtE
+eNIjTuHSao6n1wQFTI0JoJMJ+4AXTg7RPOgmvaWaRTFckw8w9j85fZ2B++d6UB2
X3u8jsTMetcmsSvTa32fIue2xoTm/6/rUXex7L7eYOipKuOxDYwUyE7/kivAEkch
dSA2hFswiwynNeGksPNx8STVFknlBp2Y1ZH0yGPCbdMu/coTHLAkd700hn2lduqu
bLKLdptWKCcBqOxXuIkiw6uX2giG6CDa2YPgQBgenK/k2Wk3QrsfaoE04UFTo+UY
MZkEPtVEdmsf6m13SLRQMis4YEEAT7nvbmRxeOmyEHb5wkbtXxeON5E6/sEFOHYD
4e6MVjtp+IMe9e1Bk5Mufbp+9tQmfHV22+H62kfaNG1/wrzr2ZLevuySPuK2qsed
i+DWsDolCwaAAEWPVkjZoTmB50pxG8hn0DdD8Z65JkUd3KqkXZivHiMdGb7w/b4T
SHDQ0rbPpYvPdrHgLjm4KiseNQ7Gk0FKjGpcEMAGVIkb1H8NFHHBSJXJD3hCe5gk
i4JTSzMXsxB2BMPq2g+ZtV+WHKgBmRKExsV415kdNYfqPQG3+UjeMVjsf24dIHuT
DFy2MkS9toSNrKB1G3w5+NiJe84vDZ7bE7kqT9Of7HUvv9aSa2a8PFOYw7RJ3+2z
9boY2XXaDChLz2xmhYanhlu+vc253t7PfgwlYjX2nW0dvMmHhkZ7rrqZ//+acvQk
o+tdlP3Si8RhG3GFzyRSdaRCHrR0ARAkJZ3TX6det9+22/veRcyA0e3y/BnWuzQQ
aHIVHKC5/vzo2tNs8ZSs1mxiGxIyIQmf4MGA6lCU7AJAGQfHr9GtocDU9HbYejx0
BpxzMZi/1+w+CRd8G/AINz14bV3/LNVbZRDVDRdN3E4rre8ViEqJm/oH3JSI9fGW
yCMCJ2kuNtTelqtMIv5DDrV4sq3wqp62tdqoVKJybxx4yplwK6ivgus6ts6VbuGb
PswuipQUEumDcgkMBHLamnOGYCu0/3Wl8Lm4jzWLKpVn6dbaoRtBsZ6jG+SaCLUd
Vx3BG9Cte2plRTsrZ35C02R0YuNrrLw8R+40RXKNB6NF27kGTEhwZPb8R5BKAEoX
7h+pzJvzW3inxfR9wvJN98X08fNjWvZQsuMQrgZ6iCze/Gp8q6fe2XL2JXNqLhT+
L51MsfYdft6WIQnKlPzv85CWBkc2jc+8oIfHoBBl+iSmuvA18KEPuLa1zDGg6pN4
p72JWz0hNXfqaiwG6r3v0+Ek1G1vW1i5TXMi1vm+2mfLGPxKYBsE5UdXV3GTVzDH
LYEvTPnRH+0aGB10u5MpDgr4kBrLk8sUd0qZs7KLIhg7jfyzQrJ2KNj7RwXRZEV3
WzP7cpGVv1NJfC9JPjfNIldPmC3QNCeCUpR43F09SoK7amxl/ljK9Y07BTS4j0Gv
v7oeKkpGJYCOSss2RaRFZdNqtpS23tStIpde0+ivYfVzekepaQzEms+07gPkDXvb
N2ZGh2t6JYkuINV17eLwos6YLnsmaFikP86u9X0TyECc+tm7TZNlH3uQCA2Tx1eX
J0CVz/D9x90k8YUeE1NExeArWQ2h8xCRlJA2te6VKR+oEEos0+Uj1k5Ry3SDM61I
11I5QGR4EW8PWkzmumNhKTxFkHn9vE48hv+7Z2/hw35xu45m/Q4pwlvI+lN14Q/u
PU2TPU85DhubmRAYxpIhTLxheTlaH0nz1RXb3NZvCE5DPTh4ipTtz0kflYLR+Z54
HCDnVJyjdOBiJNujo8EjO31w2Z3NeYtFz4Esf1CFzOcoCMBdR8tOFp7NKAjIdLYR
p49+woFtSy4Ad+jjIFI/KvJNbbtro/ipFeSYYnLI2ic+A7IdqFUF7D0L5zFYH7ml
emPCxKC4jDrKRBp1NerpheFEpAbqxAt0132DIVNAo2nWYDyYGd5+zJAi4qudppXh
ISUZP4FzMUPav1LeiugLg+jw7nTyRNquhSUCpGWFRQcENnTnfKw92KlSeKC841Tb
peo5IYl7py3IBO4bFJ27SilTnzzzL48ZQ9Je0q1SR3TZ8ryTZ7VuPCAo0aWO2y4M
CkZ+zNHdosYSJ93by1OKeW4AGbhciSJqRTJoTuV4gos0/Nq2tIwT6FLOro3kmFIc
WdR7NdwRhETSsEzQgP36cg6xKqgmDI3dYZkNT54K4+F7Kahvh92ZHPgWZYW35eOd
olSFz2OP41GTjSJ+LwBwMyd+1BluOc2PJxOrkk+KOiw34knZ+c6Yc3QXc+70Sl4+
Rj2ywcSYvZmTsXfEOuSbYbYqEAG5RZPPGGXN2dpSQd31vTEZuXJpcBZiPycAQHi8
MF4zjw/q8Pq8/0PpE/wV8TF0jQM/AqQ9JmOEvsRJhBknkJaGNwLx6z4jnKIl6YpH
AsRyl0rnGZ7QkCtXpZhB5ktbv6qq1+L7oTe2WeESPpPWgaxv+6kA3VU5QSTPyOLX
M4omm26WyH4OSPxRgUUWAtOf+iwLLMKnrcM2jtNZC3o5Lkfv+UhOwbjVDRVpsQOa
TuYHDs5VuSS93BZvDZhEU3Ldd2MuaScj75ucYtrBaFDII2/056i2B+GfzuaHsvN7
/S0j6Yv9TY7arc/bX+57Prglu6qcuYZECR/65YYJJYIN6tLQBdxj0oQuMsQNohUp
gfDVA6AbPd4jrP9+eXssL4OjZvFoLPN3cYZYeGe65GbZizrTVi7jZZFztqa0T41o
LVpXPf+JbpcDWaav2vqW+uUtA16Hs00Dl8eOzBZVfi1i2rK+u5rx66jWgp5fGaVL
9r8ghH93DNP8MLYE4fpyPonmZTzK496RG5Kj0QWJ4omr+O7EBqSGCHZ4wvTRfdPc
mtTWDJ3FsvDlNhBk5oAIRvkJQGQlIuKtDz3mfj9w6HBMklpmVeMj0wpOwlHnaZCV
dKYr5cjtLg7Tk5OHemzGfKkGwC1lVGP5e4ajmnHSxv/XYRjJkkb5gryIWPUEQnBS
dKoCJBccA255v1ctRnnRYV4sD/hdmioYti9SDYEzJhDR7hg7+bcMpiKbxxceCmJo
3SyuX7gWbgE2SUv7icEtaAjcUdafv2J49aZDDJoL7xdoM3bW9MfnagNCMoIkLIHy
iX1ZcL1VNYAAtHkANZ3+2PTCzUrSRQYoBo+YqWpuYqHl94zahNM5HTq8KwGQLj0Q
t5bXTAfa8r35fwLWqqdsaPye/HBTS3j8l0L/4O0gnCTQ5kzgZz7Xid1LHMrz69GV
Jyqtvrt5wX8dOLWzwUx+lFm+8RWa9w7S6M82TMCLU9dEfesGU5DIrDPJPBvUayqD
lVf+VFC7YdfdI3tmNvtTJZgxpoRAo7C0pvhBOjXweHP/rN80WL8Q0b6Y7DALK8aM
d3+l1cSnVFlX5WUrngt7FZFyDcN46StKptPqDtJ81GV5MNe0OXS95YsrZUHztV/R
qkEUIMp9cyYTbqCJk8LuSQF9UaVTbmpexJ4uNjwSwwttIDapcg4FRSR6DDiTUrm5
p2zEedKKGuAo9MFGxBpI7dj+KnC5RgK5wNIQYz1hrKCK3nac+utTW2qbFuVma+in
r/gRwCTv2Am3+HJCC52ARsX7QQu6tPmlUSF/vyO2GlwaTz48S/+GhLkk43nxu+Xf
10/UNJyTZt0/Lq5HkrGAjr6OEcf2sd9+PtfG7KULmvrcMZ1wzn7O7RcX6aApZ6ja
7DWcj8nth1XEwcjAL7NoG6eQcIvD5DikRYOX2N8r8mloG3vDIoB5mGSsJQThBvck
qEsKUkDFEC9cf/wULePoePqCIVwVM5r7LKUa3QlilOEmgOOe5DZ9p7vHF6mPj1W6
X8XFtyr4rmYxHoDz5uPJfd2eEPp+pCimTt+VSQUFbFmjAPBwuKrZt/vQxCjuU0rh
OAgrrg3IO667LV7mJ31E8DWKfTX7+j51RrklPaHsxVZ8eGaYFufMMS+wrVb/C3JQ
DRluMhYU9ctO4mNdveZrsP24/PZzmgBsZaj7PuTj1JQNhmGUnzgszSesFbBdiWXC
qiC0tthP+MoWUoUzqmOGRpfNQbbGROay9jlSY/hBFWBa2Iw4PVEN2r6HJMQUEJof
nXEdjYwYSIKjpE1aEGnVv6rLXBG6prTLOCEe5xToKh3iMugtVLuMgMRsreX3qE0W
V8wM6yCt0+Foj2MilasHOgFnYaWA+xRdtDVZ5lJxfdYnDnJdXuppA/kN8tczmgN2
QjWGB0oGSsOVJ/soC15+vvcaDQ0WuJBMePfT3JCpAiwtGKX5PZY1ENGnFb+fhhkf
jk0wv8Nhr6eiaS0h1Kpip7OAPH7486BTxCgo14y8wATVQrLxjo4nia7+p1ruhpnR
TCQu026cbdPxYPL6fLTFuoW2hfzxTUGyMC/5PKNfmyq8REXQZYSv3eCNbrFxIYUR
kJZ2HW1eKyOvEWJ5j2KvJIzJn+rgPynTx8Fol4BfphFa14/MaSSM5cPrkGYFjMrc
Zk5cuivG8DAlKmDAJVbarJ/7OBTAByVsDNnY4t3RzczvezySxQeMSZrojWFMtB1B
pgLR+Qhw3AMWQWX1k72cBfKZw8SE5FxnTvnYukyeI5Ti2iHdW/ql91R/pJOqlzui
vfG9OEdIQ5P4Mtexuoh44QYS+aQS4J0sWaX+aiTa6qcbR5iz++1MADmgayjt4YlE
C7pmmzBKAwiePlAOm6vdMbhgU915hcBJdF3SkItWrZnO+hHgEiwXQeuwC/00nQH4
xq4y4VokyX9g3Dw4Fprj6dvRYjQvJzrPkWGdylsll1Mjo5KHvTIUp3nLxesykxjC
vpziPrUXZ2elQQEwJPwYTWvzmgQYyIsLbqR9Gvj9yWxHhELzJOb09tyX14H9ex8F
CKOXz2XY0H6hDLzmMSWBzr3gEAxzfCA3gqE+B3G6EmlfR1SacWiBeBpB+r60K3mm
hn9ksRQXMQBlsUJ7JT4tKWO0qceQSWVPxXCZg3aOzzto7IIoXS4WB+DUE/PCcyD/
dqY8vcUd/VvQ327Gf82HCfz+S9V3oTfVFbuaV5S1PkAiIvLn9r4Mnl9iRkY3i5bp
YSCf29s5wuNfDt1GsIbl/FBLaXQY5aze0n8Ct0TcP8F6eTr7MbdUol71SZk8EdmP
5YxCjsW8RdV8lC012g/06fYQH9lvOd5mb5NlbAJ8O9kq9svzcWbRkMKWzLhaKiO9
jOEOWboHq2/iCEU2O5LWNaLOg4TbmMlA1vHZBKn3jgja5HT7pAhM1gERJ3xu9v1k
O8lhyMJ7yAy60S4uQ+gHF6B8938HJVYAQbgp4t+nPo5riGrtlP5hudMd2Dxsmw4y
j0kPHw+U+zmYd0AOU/vWEY+JlDHeBrBH7jTgGC2oYNaSFVa5IyEmEYpIRSyZlpR7
tLQD1LGT5wHvChuuoMK+QSG+8EYCd4ce0NbnqBgOw3t77H0xIy6aUxT1SzbbpOvU
ARe1vW8D15MgAdpJpmvqAudWU1eV0GFBtXHcT8MjsWD3fVPj7jcSMH7GUs3Ktjz3
XoVvt6YjwyxI0smUVTXmQMVU68SZ5bM49dYtpohOB5RysHT7RLOXXp7CU+2QPi4J
UKHpX9nKjbE9e1uY5SGBEip//2E0ORf9JKAggoJFzGwXRO1uX4r7Ur9K7AcWWrL+
INEU4ARDMvICDflaRcTG1UCzD21eSxr4Kd7DJTXuH9ASbdsjrPv/vqHKxc2SOiYo
jor5EKVROK2Ia2WyuVHu+cF54cAuXrADdcio31Mr4+lS6QTLr+wvJJ7CPmYOwC9G
gV2kiSSyEwCxJDOqjW0Yv8/Zwi8vMQJJ45mckUoFHihfUIsoYj8sP8EiD74gW6ZZ
8O4pdlxLBv7HUptTx9lo/CWNDYEos2to1/oLbrYPETDE9RBacmLFHNZezCHRcAQC
BXNr9x+RnhQL07xld0ItP2yh9x2DGjP3Lu3u4Z3RwQA0lukjgrC++GZxg4LU9y1S
IQXaGjLORrH9K04ysdYKjvp5YDOl7xY0475JbJ8M9AGnFj5+G/V4Gox/tEnIxLUM
fQzpbMG63zqQckDwrBPmgOlxRf21L/jpm/mdsRExdwj16rXn4/ZcAadJqhyiOeNg
uDCc6DD3TvttyOjYiqYjol7K/l9U0ecZJqCGUrkfsQgQFXm6oMKfL4drsJ1GE95o
Iql5MD7B+BZ7RpyiJALWJNWkRQGm1kovdxGGgppBP0seX0Fgkp3/ENIcgAaaYe9q
cwyV9BEk7FXEoT2HLcrIkbKg03+/zQj8z33Y2xC0dLhEvM2gumORUNeL9oPVE+u+
62+IjV1108nNFwvrrZyg8xPqoEqnzsIQVX1PcuX3rVtx/2f0aWsCh0aadmeBc//E
nn3QVTBAq+nQXoZLW/iNGTgvuO7CSo3W9bK40tyay8hrrm/YxVACiASXpolJlQ5X
E1rTb+hkrSvwBW3G/BDX4hqHFugc2CilqZK41Ze3cRPBBJy9jKQxAsTWXYugAn8O
8XZ3kK9J6ZQMR9cK13xmFLXmkqnjOQwDJnU0QdHR2Dx4DURk3tvqa3Dm/OK5UC02
3LC6hdq9nJtkdNkCzSNaXrR9/9d68xzwUZIYT6Z0aeQBE6GI5gDpgSBO/wgkPeWP
LAqRC/dKH1huR/3D0v8fcZh3/wOOuvcOoHO6FaXS7mg1hAdS2DMM024flUorjeCp
tW4LMH5pobkUpPepMa1R9LiFNJDLP3+6BzFkLN72MiaANp/7YYHvnzGQEjPX51+X
DKBWbVWKZZzrWPO4iMXXzUVeseHt7xm2XQjhVZcMT5iOb1ZSaY/858hwUv6J8GMx
cVsJ1LYZF8SKbA5bD3bPUzJAHRa7EDGwyNn5G2Ke4YiYyA7fyoSCEiAUbf55wzhB
oSyU3KurC8Nc/fQi4fmwoIbm+iZlCoCppXNsx/nUR3ya9Ym8aVyQGy6btD8BbD6S
qxjxC5HUIChH52Kc/1sLoAL7BaE1ChGcPKyx0UlGoeKHwxGH06bg2Q7Ou0sWwAwM
sEYdyAdoQbSPX6JWqgH/4Yay39qPV+VDh8KflniXkCiG5TYPyULNzLfHoySS0PoB
/fSDhisMSLqUqpVffbMCLi+P7VXGTMTP4osXJG+MX/MovUxmxfc9sGBoMyS1QW+5
zn91GhwGteSAU91ZIcYJkPuSdR9D5IVDWei0nsHNpeP5rTqEW6DDamHapJ7lNJwK
kc8Rxilj+JYRJqlqJomWsVWkmRjrhPsktLRDZctv1vidIfsDjngZOjNCP0AE7/mk
b6zs/pb4sDxU+Q2K5pYfwu71Qrf3IX0ZvQNAYEk6y92FnqdB6gR7a9I2b1KPFoKt
W3olZupiea12cbAEhTV1G0Wq1V5bqER8Th1kvfvlraR5madFgQdmn7XSdEgznAq8
GOU4u5WDs9B1NEggkPk09SbBibwnfpZPDifvkUjZ9b+QOlZh4PDgIgQochZor2LN
y9aGZRjtvFeSXcAqWd5b2IsgQUTS25Ct5JPfKKtDvjvhqwleZaIjI7q5ntZdVsAh
p+Ctrc4M3te0j1kfz3wvHmWLUxGN5Zvu6+j52UsPnBgG8Yd1b+yX8eLbZmamiMKd
W1tR29Nh+TeW3pqCnyMKey7EBDiTDDecyPU4mQVLBKXQBFNezjXdwgjiK3CJZD9b
XUEB36VlEsHMMnR2prR8x4IZ/oGnpkCC8SJxYJJHzvaS6x0oFv89bDhiKUkv4KDJ
1Gs4pPHDIFPYEYnPnbDX4TDn38TrVnktf12HR8twxR24p7Ei5dWzWYLCUzp8LnqV
IoIqWjxlbQuS3+jCjTVexUCAd2F6YX0YjBTTZQ8Hok7TUy7oUQb0sk9kbf6R5Vfi
Izp0eQMBG6DnpUPdlbXRGoQjhtKCu625U+2MX9UbT2spvWPNElbZrem5EM/quitn
nVxX6MJIh5O74Qc2lLYx4aDcRrrY/AOGyG7HdkT0Qs+NKO3m+xmFodN+x6opdkjU
o+ICn8aK2bNpl6fg5cATs4L/6Zslk7YbFAXe7IyD23gpGxoym1P+vL/n3whrA+0D
jctqQ8ZHvUPl0mCvWbXXCURVdV9hu8dkYV2gHNsI1y5y39f8tRbVGx/xVPtGaFto
QWRDYMFZaxf5D3DDKl6Q51Uh4oOsIM9V7LCZhIlFDoOwbrjJGUt0nbIk4n0U7xmM
oiqDkHez3n4zMc2ClfJB98iaZ1ju1i4BXc8CCarhQl8AIotOpYv81RcdnN8U54Qv
PiJ8bI90N0ruN/dE2HWbGzwEMZIWpkZX9aFIZ8Bk/mo6qnyCSHiq05Uh3PoEl17p
67+ANgGSzsSBs2O1gfql9nXMGWK1Tmkv+qnBIk16619csZEHHLX4VTLxdxNjfchY
vrbEAue3lZM1iuMAiPelQDhRSKukauY6Xp/CCBZrX5K2tiyRNB2k+sfvq1ejuAFn
vU0fj+CBVm3DzEcNlCIMGgLquoEmgmdN/IX4k5Dlqgh1Mze2vqD1YI0q3pOWlqqH
oS0vI2OXgLxfsljTgqhrtFpQ/eLMFuaYARXYTGIFgk6PSjZD/worz0S2r6OsRC+h
UugVTo3BAMqlqyEDVbbdcGDfUvOKudIJcKj2nym7VBJEXlEaBjXjFU0J/mg9Aswo
sLrNa+9chEj17FTBwOvHiufgRqmC/z0n0jQ0n5CoWm3UjMF8bosUmgs8y6JCxLI/
OhnWNA5mZwK1ldstBDHmIs6trAFm3ZESJ+IJ3+8+JgPdZMeHAEFghKUJAbhAi9kf
wxLAMod4YoWr/7QNjB6nRrqks0kFDHVOjxx3XQWw8TXiF63nUP7/CS4e/WY+afnF
PgUYgQ9J3FSwKbVNl7wtQnksP1zLcRy3EgcNPRoqbH1+3bdgMVxbFkMItEnWJGVd
xdWt/vN+Vf30CDpbHcGyd3qdrH7KnEpFW1HH2Gr/DVq1yKx2goOvt9fijvtawlh4
nGgBcMXWnBZC43u1rasoALIKRehDRZd2oxgcNDInxTu+lWKzG+HfCPuvfk/oy2bC
VrU+oQWftsLm/rElCGQ6nbhLVEYpjJAgtLQzHPbhaeeVfv8fJ2oS6tSP9WFUwbDe
QsIzLnSVkF/9aPfMxl3ZvPbLtWPONr3qvJn6ZBHdnw1StFFal6z6yclmiPi0o7sa
EDd6EzDHBoTvD12edMDL25tbIVg9put3+3duBKtgiiWOePv8Tp6ulOKOOoR95GxS
Kevl5Y7gvOCzvFQA0NrfvScAfI50EzrDafAWRiJCl1+agV/uuWzV+jIOcunaH9lI
ocDa7Z2fFvgp01bba8zFf0QLDLeHYGSnXqxTbTYJ3LeNx8bQ/TrWWe8nm1+dG6bM
SMCV0SApCEKkvCst8Faq8M55zrGrHAXoicj3JJc/rTgcz3QaaVutfoqDo2Zh/E+l
YSW713LlC5O94WlPHJG9gyjpRRewMb82ccKYPlDus4V/XZL+Cj7f4yDUoNfKVwX+
vtXT5kmAD0ELHot9P34bVwJ9lS+vi7EcReXy5g8KOnQLvDj4Pci6X1zzcO25TqFp
XiuCncXwCfkl7O3AFRwHWbNtnACpMWwTiFHkIpt8ocDDE1UVviWd2OvlrzT36dKS
WdAz3qgNUOszlrN4PQVzZyFLrIsAwuJdzGdQQOa587/3tHhgVXblffiMUr7757wo
wK268wnm0Qj2VGRXwW0iQcP0Gx8AF7nBELZ3ceZ02C84bmjEEEqpuYy46eA9TNwN
/ZII4yOp34xNUWGwzvIDinkae9GtJpCEctsSje1KgeULaGdS09YTshUbIo7Vg4zQ
CtVDc4VSryCA+PYrSVQ81/mKeKaUTx74MAu81Q0920/Z/dNRkzrGzN1BbVyKIrnM
91bN6M/8J4n/0U/89q1xOmx+21jCSdK0Cp1PJELx2eFxvKkM0bkUIuFayjirR3JG
JriveMhS9gIB0oISg2SWMl+idbcjmwvCqydBcYPKyTpu3D2omL2OLmcqW1+M6ZFw
NzVqrIjVEqAbX4C/CDPjaBTu1DNXMzkA3DK8Da+9LdXNgHm0C+UGHdD7neBbKYTL
gTgQATz1g87e/ZMxLHxdofUwpAVlLYjh+AD4lwOjc8rJMSv0joI31OD8b0xNHs0G
1CXMOL+saZCh+FXWGHo0Q7YOfm7rHm7SVQ7HhyzEnVV8vIbhC89yt2BWw3gNK1b0
bTGQ1FX/i+4i3WGBr/GZbYBal71gfU+lVqUQQgvKEV1rtGCGY1QNebjWSriA1BN7
rN6VH5iQm5zuJ9Ui7cAqW8JcdhutRvSlBy6m3z8z7L/AuvH1lNY6FWbqJwXsilEu
yG6yE10PcreqkDWPW3fisAffSr8Blrqv60xJXSM1z1Q6nLy6B2lffpgOfCFzVmJ0
JUePojRj80i5O9VQR0wvjx9N9Pte++zEuvmOuN6XokArFzsFVv4SqxCO3CtCcNMq
wsFkewE84ZbqXZpLYb7L6PeXeooaTmAim09mU9kQkt/OylE5YOSZQs6kXlGqQhJ2
xElJaVpbX4Dtjud5scHBVXZTKHqET808YQv4Ub0Tbf5BsuJVLXX1uzXzSx3E7/F4
Wa+IXmIr//roNAjJ5PxuMfpEGbdjaBRi6kuOg1aVFZ8+NyRjHhCiARJsyYt5uua5
E5s8LHNt0nL/Vjc0AGAyQz2ogY8mmOR+ZSxV0Mf2dSsmd0oCXJeu+BdVsA90gPsX
7jTkYbUdnizoJrQGSXnToW2jVotkzJpuwot4+P661fdS94eE5kDYhlWTHgmqM5G0
mvQ9/ZclZ9wL2XmZ4j3U7GXYyTp2Be4eJEdXVk7jj8hEJ0ES5orBMBlR4ZS3b5S6
pukhhwtt9C6sdSpRBu/mPyYJlqQPsduV8Htb0xAaVlDwJTLdSmRZ8xm7tcOtG3RS
96aisjsjW3QAv6v+fN1/lCbZs+Pms7QFJOJtv3mi8RpfQluuA3P9qMMMWwgZHLnv
V2as2cVv54lpEuc83daq0Ds12LYHW8emWYMfZhbdh+GRNrdJx0CpaAhht9uCNnIq
4OXyhKRuzBHUCDw+EFWusDcpW9J2m2/FS6jOz6BmVnIqS74wld6+vZoBMkniZNRe
OVsBf5hQmc2+0+4rIuUK6iXxbkNPc0OHO4WADK96seDGm5vb7EMiO/j6hEKvvBup
/Lq8NeiAer4FkS4gooucm3MPE4MWuXi0k7Sx2L+dVFe4VcLLzexXxJfivv2vVMJV
7YwO8HE+GZJUE7BRSxq5SuG67lnnvJocYp6prSrepIMf16+X+OmxQhUQ40cVRSxM
U3KqeaEnFBXIdVDaS0j/lFFOQp0PQw93bC9eBfcIFvdn5YDzFpB0vl++TFS8bIRP
X/AhdpxTSjHV16hOVTjvqz2Q5HgsEpZKbH3HqWsmX168d5EYRpB4b8zkicnpcOQF
C1LQm4EboD06BPU0Gd7HTEpjsqrXL4UsHgqGeWkjwycB7ED55WBjJOD00LHY9JI3
10oI8hq1okm60tKJLGc0eOruJBuAe/GrvhX+0U/ZERFg8FdkAANiiY9uBlvNX4TX
2WiRPkGbDWIecRAbxm6t/CfzRmFaYaXHiVlO/+cNxHBguMCEFzurPPEZhOfiUr0q
+5IcjBP6UAZhFSUF0pd6cjhBALe9uC53rifg9QU+SosFdoO0ujFtBkHaK0lNPDI9
45dAlJuOX4aVBq5BgTHvxcHGGOYhNrMrrSkmkET0k2FeclVcp3a8BYVtK+3nr6xd
mrug/m8dr3lq5+Ah7nTPmprI80vPyf7lzRcxUMJGyaRjsCisok9VZZ2G2XntyvV9
alVVKnjWdmJjvg+WYW2UAHyTpGwfZspB7Jk0VmEe8HQcSYwmjZ+OdY6kaN3W90iD
IRvcNJJrfgNKLikHfS81tl1JgDzYFVRhdDV/jttuiinyFlzrC0faWXUoHgs1tUy0
NBPIak5X3/L2474EvCv+9YcqUraJaWeizVOQRbYLuXWCjZBeFK4F2yRSPZvL6VKE
LIUL2lGASJ0eRvPCgQ4IZKbIXLli1HqDnKGPyO8t2CHjSzcCnzH2ChQOMq3SiDVi
vxmLGLTmUpTLvVK2jWRdZcOZ1VTSDeaRcqy76BFJ12zBrbjudtKBmp+QN6zHTAgf
sqBMXoX28Zz+3heTSP9nlcFcBzOV3kIBeeJzVRHc4WYG59jwEbL+Ujl+JDkLklma
LDO+0jgzAFdRfaBlwF3tBNncorJ1dSbsN1pAQT5FFO8qtXu/udvFqVA/It5Grxnh
53n5hGJmppIYvG5EBCTxDgrGTxs1LZgAlMxWz7IQQLhSvIS9i8CeP4VNXZEptgYT
RHuUMjyFqvL1I6ErUXpONrp7246SwTD4OBzOTDbgnhzQTTUh/Dy0D9zWgcQcgm1H
jqC0vjgXvOj+1u2qAs6ij2wHLICfb/wRxdmMf03/ujctGx6n4QjzYWiMWxcwZk+y
ROveLradAtK040tcENLC+bpM3WzmFanvZ5uvVrO1TACSF43mOpFx1/KWcGVgjRZa
5liYw0noQyGNBoqpx9K9lyb0/7i+sx2ZEIdy6JFRrG5k2K/A26zWGXmdNZQb5Vs8
0TJxok0IQMFpxh5Q/KxvLeqt4aUCo3cWwUXb/Ug+6zxX/OXk4jcyWek5atHMucK6
YzUbqI8NEKrh+K19XSJT17UiWJmnAv4qMKRxNgQtFFgj31ectqPvYOX0nmdMf2c9
o/kzX7P6NLQe150DwKblJYX6+MrN1PpPdaGx+qjWJzAbhCbbBnmLzYmdtqIjYFEM
kqb8Hf0oHm2jlIhR1mNQdnwIJ0Fj3WO0RMbxOS/M8qNw/xvQMJcNHXpB1FZQzEpr
qdR42ZPDO5lq7lupf4vYm6QpGRtA/i7tBDkwC6+cOwE2HgeHkEOv9wLnfwJEr2gW
BMkoZQGd/CfzUsoFGnidXhiYGjHGd/qwfxCPzIao3qNcpHwQHrEJLAz5WT4q/rMR
PKpYIrhVH20ekl0DApLe+n3X+LXg5rqjyKY7hbVUcvmoavunXO+kCxCjC3Bvqy/6
dKj8ixl8G+wtg+AQD+l/SLLUCTuCBdOQYKvFHpRZlD/q4YqoGhdUW8pu6vLpImla
8lciIqBElVbS88Km+Y4/S7lwyZmZLhU+rLvWU4MGwpw62oFohK6acFqr/zvogi6U
Z3iuMgNcDSHm7BD0ixj1V58/+xaFV+YsW9bA2OPc4ST8W81SJ4Wmf/pCe5DuQv6L
/bZOSdJ8zgfzEzNzT1AfxBf4rQLKhxNIxVF0hOOj1RbkJiIB/s6aAAxLlGT8HyxM
+j96nnWNXolYyaofhoqizOyLrp95oB9W7S6kxGzLX9b+UGWIGw2h9EN7UsdANakd
xeUfLNuPhI2ERXEKeTXdEz6mAO4UAG8V6ZtTJFeC4lIIsN4a33XDle8XNDXBpQP4
zXIiCTXoHO1clPePVaZoKY6kwgj+kzdDDLV1Klgis5l9SnUEPAmYQVNZxemkZRgP
v4yI2OlyeE5aUrlP9vSCpypTvlIIV49adiASLX4YxifpH59cthf1aWAWOrHNtkPe
TgpjkqoJWBnbW2qc4A7jeStYAxrVJ778R5Sx/sV8Uah2YiHFycmRElMSucLJG1i0
6YpSoGctlDp9PzPKCeScmOOb6frgzVNo/NTDR5u3MWaJyGdLKNoHZj6I9ozJpklm
+J7Pz4tmKk47ehkNNHNOB1fuGjclWU/HF6qwvEOaopjRdtfeDvd/ZwEUdh0+1wMZ
v2M1wAxR/+IuErWVPKTD+HWEj83f1ttLvBNesm/qnH2tRc/vvqIbqnwlpOC8xept
57PTTCJW0ajvYcIdSTW36Y1CB7tHVQ/1DCqzPiN82UiihGlDpt6M0RUBSGVstjQw
HLmKZvVcsDCakiJ16vIWcgIQz2zY40i/Cn8mblIbxdZ4gVm19C+0VqNgmTaJDpj5
10I9y1UqbmoSgd3le8bOIrq7hocFSyaRhxY+oWVMZf7SA3JZnYBu0QB0M4wCxHgF
jrluum7lmq6z+BRTliWqnkDGZwzCaLaTvdSTWpskBrbLvPx/x8Nw/wG1I3be5cEt
ThwATl/ia2ttf7KSEYqcM57UDzPcyNsSlq1hs3m5C+wLI4byUAHl1WwriDZuQqbe
d0JzcnNpGr9lw1wKWHwxWrI33V4vBHVwW1FSB4WDtFtmaALkEaYCU/LwOyaftPAZ
uNVKyXHW0EidHTvxmegxYzPBB/T1l/CHjvd1TvunEm8URtIvzQN6nBvJnSUZzbV2
ZlnQ40X64Mc0+6HHvf0NAhusqxaygj+ghdIPLBvmvS7Mt9kvOeGe9Tz6h2J7O3is
F1ztDM4HzjQEsM9N7yLRZOM5ekt1jmiRCCByFKfQyBxVyHx2cR3ATZmCBVeLmXlx
7OnD/HRcTHKeQCmONM165GGS3NGwArZ0kCZK0AIgu2Uc1HIu+6hUsF+QezRmdAPQ
CyLtIkXUdWpQXQm3mt4ySCzpgufWcbHM7RZFU6BjYD0+LwwMYjYtYQlDpw/AD+fE
BdQIME33Cy62KKcUS+XCBFXONYJE6oFyAUQ00UaLHeZ8vyBPpeljwRjkUvzNIqqF
wNvrFzzKuKDteSg+PJlBpIRQBJAwHJ7t8u5uWNiAsJr9/INIqOXv+3ahtKb4LA+L
Tl8kAmzt4BDyV3gi8PwpKN1bYsz7+NgY4vnVPX8vXdbNoyfyprzQmtQsiDcMN1/s
cGS31tWnNKyc+QRmOYIfEeESq7kQ6lap26tQt/i+QEm6Yx0rr+Fe1QSGBDgcpeaT
nVk3cOJtzouE6m49d3OKtvqFTPUIZ0ZQyliYNE75SzUvN6H37budDT0AnMI5e1NQ
VRLO8pZOaxB93SxqGeZy9QvAvmcp7usmMupvGchaDr61wEU7prvWkJJezIdxXLcX
1LHYSjfZbISyj3SO2ccEYt0qJedA4cE8htJNxfMHZK/f41aZnd7Yr2bNZ20Yy/fP
Svsb2eNDMBtU/MlxOxK5CAvcOD6CWMkIb97nM7hDo2nBQz6rkqb6IpJolkp/hP1j
GkfisZrvyp27UJeWiIXNKBEUf5oKfMmyr6WnD+T6OJvYLXAdfx4wa7n8IE8FIc7j
HpbajVri1GJKbzG+gFnXoCocb7kTT+uQ7gEXCAd8NvaGzDkGQ+gVjLhZPtQGUW34
SaZM/qYDLaFdNakpWLwkibA3ecsMqXupycl64b4SJGtIrCv3abPBooCrWpFDdlWT
4NNz3fu5a+8bzDTiZJZxGn3HGrbRe+5tcATJpMVrQf46OCszjQiSabyKo9EaUOaE
B1HdKawEVkDw7pH0O6Un0OMieJh1/MjkGETyS+cntJC4C1nER565Fvdi7n8BZe8h
d6xBoMuiYYK+nkNmwdCYuyPH+92jVYi+7W4b0JKwSp4JuDtCDxqYjH75TfwPxAZb
6y0wle9swuHF38bQKGoZ31YLXb8JSPVAebmtcyMY/Pf55HykhDTAasqjFSK5gABk
oqlRFBL/eHn1AjpW2vrKp3lBB1F60STvzQ7H2yiEww5WkXfhqbWKcg1Fy6pXPolR
OC3rcxo0l51ZKTVWvyAOd/vlDGbM06Ir1W0joTDSNlhukcAsI8MjmjKSICnbvQJZ
RdKva85JUx1JdJHskITMOl32qBUk/JsrzY+pzFtBD6iKOkEsxqZskWG1XZg2bRsk
tFNrA0kr0DswA8qV4A3Ba1ScTLeFoBYl+WJ5l2CQtJ1EnkS6d7G/q2htjgjqQ/21
fosdbU/yLn+1iXBsLe7r5Foxf2eT13SXmgiY73O2DAiyrkweWk6C596krRXm62ca
jBb3cUS5dryQyMJgOQuLIpPORNq7ks7qOKSy3AEmPinb9PmSaaoEuiQvW0tvja6J
NSPnQqD7nILVOsqpyFPeyRYV5WqL22NH99hy5faU/2kApCaVwx14lFRWZRzZTJPS
S/xYo+C3NPp19nODkJpnIP090T2BgZ5AvaFknhSuOELmF3wx5n5MecBRL+u45PRU
LeKo6TKbvBjvwlhYbiepo/ll62/ilwprTru7NHvEJZDTnomcydD3cqTf5/Zgsffw
yZXZk2Px++sBuidtZOV5xl3MLryBB8Aw8FvdAJTXq1fWaPQO0h2jQXwMEpx2NI+N
AFFqyXzPEoE7Cb9KX+jCHjP/f3InbGJFPY28nXWXb8mlkAAIQzz7+5hsVk6D4XRW
AyeyNCRyh3TwY7m3M+pte4FNxJn/BOs8UeMr0Zgqb754uSRcA1a9uAS8vshkJCoU
5umA7MWQscshutWfdIAPazI+YRIKTLJlzgYtMJLk22qep2iio4qPEi5R2yI67p4g
jtvhUs1yBlYeToz8Qmbw8tSV0WowN5HpT3neF054dpwEE2LEW8ERg2IQK11y53bE
mCvRjxVMBCe5YXeNLzwQSWOHly/X3EakUPbBToFAkN/sOOgW44KrAddnEIRm8NK0
iTXGJdxi4bIjED6bl5YX74kqsBRyUrBpneeHWng7L8kF1Ofe4tMbDEmVbC1yyl5H
Ia/A/vgOrWGpIkGDJSD9SIMiSIPrX5Xucip9r1oD/xqN5wVazk3vRw2QcoztXZnt
rbk9MDTcdh/k4whd66TsE7yVCPxQeW7rfoqSA//DG1X6G0RtlciUVoPh+vvr63PM
l4y+ISQqyoKgi8Y5S2MNu/zvkEJMa0y6c9NhNVw0bkTP2y5Bs6xjDik8FgY794Mo
AbkJ01gTX9/oAu4ljWXktH8cR/3pQGMyBGkeMvDLcVifaKWiLa5iRW5TkXt79f5M
eY9fCcKiCezxrquD+fAbUF0iP+LkugBQMo+19y0cLTtzqvXysCoUOM0wAx8yLWW2
v+i6VW8w+O0hvALL2ZLtVjF4I5Vk5B7TMZ9IWmW8+lNTPZg9ordK+zbNDRlMXVmk
srxPc0TYWdLIsEO77W85TfqQ/3JoXC2tM30cziFkj83JFXI+BYkyI4yysED339ju
eNRbgxWutjsxKhlJGjQFpbZ/vmxUpRpyCjpS9QFTZNyDO8kFhnhm+dMnkIaiyh8l
qXf/vlUIectpgD0kzriBHa/1/DO0WHJiN6dngzT1Av5j3r1eHYYm9z5xlrA4hGgJ
O8l1IWjA6o7Buer+3hNdE+Rfg//++ejT0ds72bUHL8exuuEgi9sqz8VYslf3D7v+
iToVsgYUgzPbQunwqLZ4sFUzq64v9ogayBzKe7ziyjCjvlKJ5kA1qKftee5eFTxy
+9ovVZZIi4QdBJl8M3cEw5xeuLiUi/K4TIiPhhW4RtN/4TiWUn/0ejtziEW9Tzrd
EniErtrREVjrRgoWAKXDKnGVuRVy/HPRP7/MNX3juvqWGVQcfcojTg66k6BfXnQE
6cTWX5BEhDWAZL3Vw94fgQfA15vjK/1peAZ/RW28G1wQLz1AjnxJ2x6EgpeNMwpg
dwCE8GgHkg5o28JtXmE4JC3Y0jx8fKlVLVpK2IHvML1DprXhxUVwjkVHEi/T9m9z
8o517qAbuHmvBPtUxjmykTB3WGNgTHuehCmCVQs5p2InqelJLr9RNmgi/ya4DHue
i1Yi7asUoscN2aofiJiTXi92DAwdtZX8R5Qqp1OETaYZCblSe1E6BusZMaWPB/DE
HFBvGlKUAfPtHq+pO86WnptHeTwbaMrux0z6vKeN+t1prJMkAj4LhCs3EqXG+vrb
ulXLnUdsxzpYL8fjnv/MNDkg75Tn2U4GuT15LnH611ZEmHzRV1TwYWc3pio2pEF0
h9+XOS4su9iw43CspMhEVUXqR5qAMp5az5tjiXH2TMy4/p+qkX270GQ6UV57693v
nUfVJtYFM1BMnXBKpI9uk0Enl8u37Rcjbyn9iuVDcqdIKnDUv+/spe1a3i+io3nU
l6NJvCRjjviG4izpJxxt8Sb3ZKTB+F9wPHHmvVADVr0ypu1QqA+1DoXPEhCroxt4
4XxGcP6k06UYZUqsVxio3lcJxOtEQ85SwODJifL48+wegMtw6ezAjrOyQCErHBDM
6xEZXfpdlMlQfBfKpF2jO+OJz7qkj2UEYDzhcMOeX2V+zm19qzBBJkyVFrZ1c+cu
DzcNhEhCJTBlLAsJCyn3WHmC41RUxMn8wWVTjyFGUMOEHGOG3a8zQlWKSn+ZNAYE
1D1M8b0RbIkV8yeGUpyAH8s/KEVtgrRf+saGVUNbx5zwisgEGlPUShMXRN+RaYBU
jeS18isjXbAhOMsbTk2bz5gGS+ofjTquWo2MO8ufV60wP13S6EXAJoGrwIR7yBgz
eQ0zgwJ74ApMFW+F9ZKaA2Dp86TNR7IldMH+rEQJQovAr0hIO08ErOY9YgY9OLGj
4IpppoJuOC+D/1uY5L3f6Mv6xVlWjwWPC54RImZl3saocimFte6BxbXAoldiesAf
GM1ateXNE+D1+W1OoLRBZr9rqyOD9RHqSknDZC2cFKqi0qC1tY22ETdmRPKC0ANf
ST/Dvc7LOF3fOYRKdVjf+kWdEF/rVK98FHsYdlIFJgXOhwS+yKkVQ2pHRNVCRsC9
i5NfKjTz4OqyEUziyKyP7D/EengYqfYmgmVMfzwU8KvauGgQdHl6J/7DGOfWtjQA
G016BKdFZ3SuMysF4MnaN9UpFDDec6g+s0REZYkm2AdaJTO0ocF93GvrtKbJQpdv
V44FBry+/0JT52RR1qfa2v9j1CdEuLtznVm9qVETiviGaaVzNqQvD6q4li5hrlc7
xJM5wHOth9CQOwIVnF8WHqbf76cKJ5UYGZaMXNsp5r1dEDp50kMPJiVhPbp3TdsH
D1asWuWt7xhpNCICgu97X9ZApmQO6WTUxNaWJmnkmiCaQOFS8she3Z1zky5vc0fr
rUCatC3QsF20sEepA2DFIoxMiyJdIs1ZR45G1BtQQCCykb6qBgqZ/MMhQGmfMk5b
NOB+HTNok9ohmWDXbV/u1Ezz4NAlFRjH0TLvJ86AmPsjbmQv0Kxfe9qk01sHG4gn
g/kQ0Mpl3aJYspUv3S+XLmf5XrTvontNMw2AKB4+iOrS/j5PKTkXsVnXqu8sPqIC
8o8H6ZbrUopR8DQ3zGr73USQ35bQa+dVsdq9AUbJElBAPqVl1Wn8uUmNAwkrq07C
7pHwv/HZx420kAp4g8/4lleJkOnj3OFFE2uuHlqXlkA8gu/AJSW7SJ44apDUeUlz
T29b4srgs+nNjB4WyI3pCQfws2B0wp8/jfswpMPGpjZtXXqE5JZKHZ/Q6hSCCVX1
Si3rsZ8U+gE1oG+2Kdbcn8Ibo+/a19QX+REF9vhrt3poKH5DKRGYtuS/HSJp7WbK
fQ4KbKTNLGjSKYZdopPFYPVw1UgULjq7jHZMLwk+s6ay3E6sYR4bRrqppBFQn2qR
vXJBbigqafvF51MKJN0b0jQdRv+bF2QOtW/5/xKMSPm1fpPXWq+4hgsckDcBfFjI
MRIaP4WQpJ7rAsLn7hfqZTbnXQkLqbWOPhvY7DFh/ZPG/+IAkAgqRSJGKPOXQEU1
4GaEBTDa53igW1nqwzUKLfF6ysb3lKLa7xG0aBZ/Rho8DihCAr6OxqK5Pv/BwN45
qmlxqpP2Z0gW2eAsJMCbzIbatW55fW3VRHg1IUA+BFSKaWZzjvwYi6BraBhyt7Kt
IV83oV2EuOqRlbljQ8L2HwtXqZ1GHTr0AgYC9E2PEOO/RnpD0z458BJu8OgdJJtc
e2B/vgVVVfBHZdMlMSIUspXLVV5008uVU5eHI3CqwCeV6IE1r3Vqriyy7zFgi2bf
+4Ylhl9OFYhcZrdImjstZDpWJxEpezLd07FWh3rJJ7fkgryWbteqKTd/38s1FX+5
pLFktcwAVCXCeV8lITH7cc4wazNudg/9D2oChos/Mpm0sV+bv2LGw0+u2h7xl7av
pnPq3PzhE9GKSyAybh77O1fDoWwCnFgxYhWsUQ1l1Xw9zvgpRO4CvA4WKtUAEPmw
rY1pzbtohwmnFM5Nuld2zpaU5qwAE79NLPmm9Bxxs/k4+0mhb5NkIr421JWtGGs+
JAsfegxGhPfdVebCwh9UcPLUiJ/MQK8bHhDwVhEfIzu5n/Dz9k3z66zr8W7F2/ay
uFZe/QB3c2ELz765tJGZ96yx2ry5bBlOekw57rEeqt5eHx/zoqPdYzXJHPOcxPb5
DQp1jVH2xZ7UALR8ZhG7QQ3tLG95+deFN0JqwcnumtR8T/UlYL6b0slNwlSLfGHY
ZjYqsNEqxYP0D/U5nRworGPsxUGagEn3L6L6JV3lWHm8zx3zl4tHw+V6Bny+QWyT
3M9R+a1ngiGocNujWnZr8qJjTb0T6D0XnciSLs4hWgL7BwKa0prfvx/WPhWJgsIM
oZd238iaNgGbmzpW2kXjU9Lv5c+2kjD5O4NjReZy+ly2MlYGJJPgBBgoab6ujqax
HJto3hl8wth5QlzaZZQn5f0eaUd7JLwe4CoWMexvELMLotNK7B8JNnTVYAtIupGB
uVpyeN4RAv6aInh+066/97PHGgaxYjR2L7q14Otc+NXqJOa/uJPoKcKD2LVrwjDi
IWvJugb5qLfmXoACN59fBmqfOYye/X4ZeCxLdkgFE8pbuCmi6cmRYZEUIziXBqlU
vu1d3pA8LL3h59fImnGPMn20rxY+gG7EQ31PQOWQ4+gzxujMy+EpCh2ZaDfIfJnR
ABncTx9tOijtjuOhX0YpcvwR0K5YKhSn5KkUsY8J1mE8kN+/vZqJq/jCDvf94n2m
jaDeQvoWpS/aNNVrcNX78Xj9PH9rLYksEQV3MYcYMAMdXT4LEmEQ2XR4SfueQImB
xvgTiwTW4w6vBPo9XBZQ375WEDWLBSUnkqV00R5Agw6zEDr9JrpozR4kK9q6+EYK
RpjvzU+YfgzTM3OTfU89qy5hMG2Y7g4uaVu8kccdoSmEV12wjmBwel3kmVrJ8lFC
egAi4LsntdKdM1iV8GNchN71W60fpUklSRt0YV2kgxtR/YV4ZInLLR1mbGbBckEH
rin6U8jpiCUf9ADuIRT4eQr7pQb4XP+Dq+tnO/oMB4/fWLNYaal1GG/xJQW4OKai
6nLpjeedt33T3Wk5PzW45bxQ+IHhNFMhI0Tfhf4jMczsFRjrE9m6Rl1rcO7/IFZG
NcsoCZwJkbo70RVzP/gvGpmTINnaKRFHK3rjfBcKbWKZQwvm4zXCb3c3zzLjKeUN
Ckl9N6FK9ItroyWrqf5eYviHYyoi7hvjzgTSJ0DMSfVAArDEiHgdMOOd3Fq0Mk4X
oeBgHUkSBks9dKDtV+UVcA==
`protect END_PROTECTED
