`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6ZHvnsIC7Co8gZXEUWVWIsjqLUjIQDRnCaFaDrGcu2Xm5mN0h53QNA2g9c75WoV
xyDgB1hAquH8EPRsD69PzuexFgvru9Man29W5F88swUplWfPsGoY1WmNeqRIS29S
SjtdZGcGApiYmfeskSD+Mi53nWUg271iBg2XLk75XkMfdB/noWp2vkW/Oq1CrXOm
1YtxrXT590+zfV00UJR2rNf+BZJX+sG4A5AxoKFmbGwTfZW4myCi5lLRL7xqOj+f
CPp9OnE3Lv0O/KPCfgr5VJTrkQp9BAeNRtxAIr+ZCxLrtBGwW1FnrDgTCgIby99b
kt3Vbmw9m9DM5gNQU5M6pQ7WF9bgg9x0+TGqWQH5QQt/UlOWxI7xH6FSogPO4+ll
BREH/p7TeT+V7PR97d8hI9ACI+NCGCz7mxlJ9ahCfoey0VX6Rrgsux1AFP/I/e7G
vuBby5q2OlQNg8C8aAyTON1a/evzhCNaJsA4O3u5URoldPHj47bltyr3/E4psmAP
O9JgWSci86i0vMtEDmR+hmIS3qoig11d96N/QL4uuGiKncZSXWtabTzlc8ZyrL4B
xaKJtQUtrwIdryBrvYjhlDn0coivroqX8xtL/YeFHptfYf2rpfj64EI7nB5hBeB2
csSDa3AF1NbFUwvUPBB4IS/6mL7rl7vtIOCFNvA/himBQJ+6gKgZgWAwXAYxxC2+
PbNicU0umH6JyOvkX/rRucQVBXoB37gMRIaPgo7QRhuIG08K60IY8dD3G8nds/LX
rTbGinK75PGJuMYGARytgW69O4YmLccIjKnv/C2ULI6ymnM7PR3Ax5BP0pSEU38W
Qh/PG8XHzHpkPvYfNI0pr+IpPK3b43rSGO2xEfI0wQTj4wvduuuzcjcXUS6+NXM7
moFhTy7kMdol7Sy5M0P8KqCZ4aECtOjxL8a+9tOSjijp33/apgw1dFAypI9rsDJm
PAkVZW9gFS3vl2m7BeuFD1MdCk8Sqa0Vuu+FGdTogKLdpyT2iMyrwlED7prvsPZO
Wclrv95V1tg+hl2GKi1tUcFLxbMyYPthsfoEKFGUDrZItMg2tyGK7Px4uURj1lBM
8gSexhpPv+NYjFd0YEOkj6XDgZG3+RnPsgbw8MPby/4bWMIUbvt9ejvqRwDE8ziz
X2F5uEW3scVXaIsKRF7XLxdXanH+W5a9baS8lWJJ80HkaeC78mcqDJ1qH+efuKbZ
O1BByAOKMY7JH/CZzacRu5aKjKzIDNMT/EnMd6tB/tTKLI7DC37vDev34darSeME
aDQWj1bxYE5zwz10EbCa9nkl2uSMytRzd0MgO1URgCpl0urCLGgID4UCro6PpvLw
N9yafPqiethJA8/LL5wbnLjE8anPxz1mCPVn3bWlBLu7yIRCv8L1/SvSWHWKU7ce
SmartrQocCuQJaxuivsaUKir/hy/crRmwyYwycEKWoZitC35i39ZS7HWOUh62w0P
5gsEy/KM+gelh0P8OyllePlP+iuIO+wl1lMrXr48BMDMapOP1mg4qSY21x3vIAwB
GMJSwqikRiQCHwz//+s5iZgs/YA5ROKWD78Cc2bwdOh+pvzhNpeiJjclYl1FUE3B
dF71ixbHnImfPAZxBOT246MOlI4TYaPIlhtBSdgLSioVXqy+CEaQIoioQBriDfoM
RTqoTXLQATXB+oNCm4rpUiCxpss0jZs+WELEtmQsYxv4gl3YPgXGbnJtSwpVBjlb
fHWw3oJtGQ7EYcyBhVXb5hHLlcQKZubFUMaqgFnP68WA29yE3nDHkIt+C2LRRdv2
s874Zo/KKfE3S9BLAwUPJhGqQruGeoT1pajvt6Ojryoe860tVZ4ar8YG5XvZrWRD
6Usj1Ss4b3tivSkq9lu9kq+HZJmNv1V11HdhPHZ9C98SmJNPV6yUZPdDScbhzZiQ
JjipxuGLV0fC3nzmiE7hr6OU/f6CnotvbMfVGdg47ArMS2aLnTm7bYxS5X7BMXJZ
AKZhYS/MorCOOvEC76BOgi1yeLS75IMsoPgED017Oirs6eHwu5DT7mpMq/DyZSa0
Mtc357tt4+uh3YO2JvM56DO4pwiICcPWsI+4HByE/VYLCdqVVM7vz1H5G30L2vmR
Rgbq3LIWNx5vzriduG0vU55d7bkse6OG/DWvqBYhPDMnKt7nkBIozBc0aBkLRnmm
YEkn80jJJc/atjoChsLebRKVT1HPyt7O8qQMbJlZmN/rbCOYaKC/vF+FsPwNRkVe
iIgCKEIKxk1hrq/DBjp3t+aSioU624aI5VmJcdgAO28ayTzP7oMt+2FZuaNAMg4a
wBs+464hIMHXdbaAs9h5qF0EVdNtEOrpaLqPoAYhzCKUB58KBwOyMPTsD8VEr0G8
VaQNn33PU8MfMLowFbtuXJHvELC34g4v7q64qBHsHjRgDqjeMlOdMijCHRj7X4mK
gsvOb5L+4qPxs7cS4IgD1lx6BcWm5LP7suC4zMPth8TxI87KME7CnISIM/JaCrC5
X4mg6Ep0aaZ2dxu35HrAxKMZkjjshj8DxuvMwoFbj2dAYz6c2U7I97GoepQgssb7
xr9lFIzC4olUUsYuo5SepP0UNAKaOK1SJMQUrea+WPC7mLvlxB4WjpJNQ3DfMrl5
pd49TVc1N2Pa8bYjY4JhPAfLPDIDLEfR42ITOSMzfIt071inzDUepfyVUCfRFA7D
OLjF8zPs1qoEG803K6xdgMRSNVT9t9HNn8vSzD1g7JXu3//xAwN/dfkl9Qwx0bXh
YL1qqjDakhcWmBiDJb+3pybFVo3L7/LShHpmSXXXahD32qPQmXGd/UxkPqrrzDBZ
jwhFY+v1AbG222nxQMb/cnzJgGW0EgFlwoTXhbaWV66dY+gFZWHcOaTs1H6CTwb/
p4byiHbIcI6eqzOsYggO28TDZxHMof0sd3TBDvxJeOb0yU0TycWXjiUh+meCXoIM
VXbYk2cqNvdSd4gvF1MAGYxum7uuzs80Qkp5urKaNrYsKmvfTRWxtVkhqc0Nfrto
C3pzCCNg0ur1feKBEArOMVcXSTVKHT2ss02I0cr9OUk+5gypRSxt7CV6HWieYQ4y
Wzl4RXw4zHmdcggp2POqipl6Ns8SoWTVdminMtBR7niSkg3FKQ0Xvw0rNA4XQ9pj
pnmw34zMciYXDz/SznnWuaERHz5n5VQr72ZpbjpKq3ybGrg1h59RcQ42X5ecWfyL
kn+4hD/ofW9890TSW2HY+QpkhGiz6J2DO99fzpxPdtb/QoZMncfoVDVaBhSaaBXJ
zhB48bSeHDjXuFt4psiSVoN7O6VT15gq0qQK5UNrk76RDfBMUgONRmfP10SomJoA
nD3Tqtch8ptzQ3cCsGExzkw6XO64ysP5JtDGT8DALoS7CZWEK6y0yegkbg5CT67G
fX0wARtyTV/aU1sfZWcxgkVWKYogkcHbwewclY9mwTAUAwVWj3MWJuaIArbNSmHe
dvTU2Ffp2u1Y8w7CEgWK74o9dhp9FYMMy7gLEBRDnQ8ftXHwNwYH6dUQfMd6rKYV
3pVnlnuwCiWPRUUh41KQ3htOls7y0EhXMZCD6wES7EMPYw4ceDACDJ9kuwXTdWGh
jMfC7wpPzu8Jf07QNSYzPyFqU88N+xTfVncGyL1vuEkmIIyqcoxh+57ca8V9yAEM
Eoop4s9qf0Uf4Dm3V9FHMlvOa4WdpWiiB/gWdNtWkYcFiyDCMP3Yik0zED+tHb5P
sC5gjbi7796txk7JcO4A2+90nn2xQXLuvks2mITLPUQuOZrr5R7ffzidBkNm8Pcv
79fpLVvWcQYSHkFPHNERLPBC05yJBUMq4rqFeW864Lpp+0MR3tAk631A4H2NNOMR
bmIu0yBqAWI5dF8z9xbj5HYg2V/g6M8hejbTXJ0CgNqyFjO/H4RNxz1Opkh6dctA
dwC3o8TJuV6jaUSVFdT8AW/RBq3WILEBwnwS293EdoI9POc49aC8U5zdJO5qWoJE
5jCPYCHgNZxWEmx8QyIeekDtwYhjHVLfntsFXxBRjo4UyiDJsvzCOZFXDOMs2llD
FN1aJKVYivvbh9ogglSbZqo2SdaGYCCKlohC5Xkxp+LDxlpwMZu26rcEdweN25NQ
DpUMVAIx7YUKflcFfdQNUdZpxgJo/o74ipH6FnKXmipGllI6m/fHHVj9jvLAvJHt
ZDT2VHLxxAin1lK5NZhGNjaAI6IRHVBgt57O2enUqeG5RdfaLulCp4NBt5oQA2/C
WSzrLeZvsa4Qyl9NWZjlsQ+QeelLF37DOS0vYBbMIBMIPjO7Yl0rzDYAZiUmOKa5
qCr7n219SAfe5aDwwzOGOx1zOfI5Sv2wE2zHzVOmIyiWiKwZZ0wOnvWTtMgG0m5L
vjPFP5z0LU5kxUrjCocgShg9Izc/0ASt29cFUUjM8CpHkIp+J+qYs77kYWwEvsRS
TcJDqJCuhCj6LqA+i0161VC+sCavsRludntR98UgP0UKgH7iyuoc5h11zooxNh7H
VMRmqPuFJ9Q1joXOl2DXtT+i9Fu2pHeP2jNghZeNDdnsvoxNKuVqEsJrvYnJTy2o
JRGYNHU8vTkV3FOXwtT24fKYf/euR9FVnA7bwE6+QAfM+HcGxUjXT2zTnHP7PbJx
1fql1KGxq09E+aEV+9nX4fvlVp31gr1NtcjL/FWj+iUoSwUPyP4MU2TW3thZU04U
2qCIsy53mYJpcH0kQWjvYGpH03rvXqmva9ZB+HAkxi3IeRqvvtTnV4m65k5P2W6Q
4lfirZhyOM7SoL8IyhZIbPkHw5xy+011BtwgygQ+FK7lzwDMTH8Ll8G7fZSDw1U/
91G9oBSs0+8wLhs6FwpDjZsV3jbiZ0a78Sf73teO6iGc22HPyRat/FNFkuKjSJ0Z
fQKRGTK/5nE6hnJbIB2NRVomY+AeMlucLP6q0DHNyVDRCzJyixKn8hgfOqi0DidP
OeFiJqN5CFYYD/kpcnKSp8iayaqVV5mBLRSKi9kcayQWJ6Q3+Jr9tXhd9XmV8amy
1j4VkHxNN+Gb7ycaHyLXOoZ/MB+rM8xmU1glKXpdmU5DM3kxpoK1WuJAF4k3ABc0
SKV8tgDZDN2f7NadKEbBImMFY+NFC0DByZQzfKn83Ct2zYee86HjGrKRbxctVivO
9668KLSW4Mmw7OQil/R24KGdBz6TYq/4z5SKqZ5FN3G6W4etg6fak0oh/Ka5AWzo
xQjBJTTR9wk+w5c7k1YrHVU8Kf3fW/F3Zj3NpS6fUUcPE07EKVz86ihR0iIYtO/p
aBhZ7nVoA041ic0bPbi51VV6S6KMVfqrFWPTwg2LdgnmH0I0VFoqPWGVxyb32Mhw
mlEGbaAdDrogS544ugTP+QLj6JEGvOIxZ5ERQQF5piT1B6p0qCL98PF4r9Gv6uSM
L81RGswym2on2RqS7kmExCbi6ThVFQnD3Dp7MdOKlrV4PyYtd5dL/NHEsHwbjxvd
tO9/vfnsxCDaG3tlkm5CAIHDOcQNqQ2/w5cEqbhMQBaNsWddyZXPUX/qYUY8abyx
v6AzxCFRlA/ZlY/dS4fA87hTFOPE7OjSfLS6wM2ULPsWraefa/iOSZp+PPjyH2r0
G1C2+IIuePvXI4pPMesh6x9wigJ9KLQ6UYV5fCN6Y7JGdKO4ther1m2RJx41v3/X
i0AVY25WxgxdZQCqhbcUkrz4kfDcZ2TJA06jqosf3C+AhM0IUf2jvYqBb2aTErSN
RolyyLXMo3eUu3zNkRthJRnSeoCja6aLq/UStQaUAON/ie/VQJiDSJtFySpogueS
As0n4GQIXltXiB7DdlQKKNI3loa8x15ZBPpFwquVG7rnFGgccx5FX6f0KbVNHcRq
Bx0oQYfHEEWiZucEiR3X/nlKN9WJR2ownJ17FvJDwKkJr8fsJ1aR3sftgkiwA9Ne
vGOfDKCut97JPesiTMXEqpT0/7hRp9cr732lTy99XVtq4XP2Ufa8dLlLI0/2hzIp
AvtU6VwXX3UNOsWxHoGNfVbhY76jXuCz932b7Bqzn+bkM9veSVVG80J9whS4j6se
TFcWcOif7KwYzo08AdZ+KP71cmvG5N1+4dv/pSQWtiBkCsCCykdv47jStoKLoOMz
6o/+9XeAp4AJsFVKc3OZoPddk5DHUANb0tU7a/9l76LG93lMKhEvIKt0aNBDz7Wy
hs3h6uwbkv6ausZ9nkX5Ufu554b9SkEAoUfuy8XL+k7l9ZDRqYB9RYf5577fLRjX
/hMfGITVLBZOZam9bjVNYs9cC9/4RM3TqKxt/i4Gyrtjt4kG71sandY1uR0q5KF8
rHCuTmpTL0SFNNMCqIIir7JQQiaCyzlOwC97Wvy5qBjRxjk43iCuB/EVgiAlJBeW
qEFlmn0P2990PidvPGJmn0q2GQwiO6fyZb8EMANeNSzUZAoxaOSpslh4unIv4xJq
q5CIAK8mG1890L7N/zRrJT0ipcqMahCzcr0vYojMnbakUlsQUsiMC37MqavHlXvD
QI8Snb8LZNkxloiYYP1UxGzt6QNcZ6pWNRMB49JomaRTmad7JvyZXZlciUtX+hQO
hnUNHWD5l7FFBL/fxSYrovYZGu0NKbzDzit74ii0i4JCWQwIeAw2HcCI9vCSzcI8
pW8uXF7mB82OZ8yGkEHNY9YsDvoG+0FieGQTv86FB5GQfxjWKFlbrxL+LbkXKiVH
pXSj2tYh9W+LFVyIywbsSO0hG7+xxlenQdC5MMwzW/q9P5inl6OZgNO8INJgP8Sd
QHjIDL7QdR6XL4ARy/GH20h0L7ARmP6EDkdZYByCRB+FSkEybxzYZo8Sapc8SYmy
7qsNA1+NJRmCvlsnY5yxlgOL6sQJaTaPJvXokdG+uWGLqY/IixC5ad3yhv15a1u7
ZaOT3QDTdpQE1V7TWqxs/kxIHlvojaEosuZRhFy2upxC/aY5lWbYAn5oSeG2eFdp
atjRwKWRjybV/5tR32i1ygQ1JrXXwBuF1rR4HiBtoHVfFsLGfQmmKwZ3NXuXVp4K
HGjtv+Pu/Jw7nbqfx6bSInA+u6vGI+xIKcSaMISHgX5wsDzwB7tQ4BOGETXGlC02
R6ohWTqtLPyp8oZYUlM1+W2N+Vc4o6nDKVyWc8ksjEbdng2fEjyu+Q31SVlnDMrm
4vDRawVPtFB/5wm7E5Hk1DZSoQdBu5x1Rqt9svRU3xfoZckn4eGVujGfxQ3zY9Os
30au8GseKOJuKK1/aKGWbDFB9pqDSC0xEhYwcGLcyAT0SU8QJy68RNbFyTkTBsBS
Y50myoorDN+gtKHG2GmSzxmGCgdBskeza5AsqysImIJIwpecnEVlxl3tpm4vuiRv
AFU5WA9LDcFGywcenRc6ugW+chbH/0pZc3zkfVQsZpw=
`protect END_PROTECTED
