`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mji8TZmJfldM6NMKqJMY5Wsu28ra50F8UojXRZQ1EAgR5fjUprfMgX8Py5YIHOoH
kZC5gP4FwIUk3gmvgKNPyx4fAz0oiOP9PKAnYOowZR9yK+aCJ2BxdKWnOu6qoxOU
Vpw7gdERPbsReLTirihsjwxtU6EwMrwQiktKKZAm0JZPFi70DXvi0TJaNhT3g+Qc
QDbz1G0oPdap0DxAXNt1WK33md9nOYmJBk8sgxptcNsMqAN7c6BXAx1qobA5NqC4
Ritq7no6c+lw4ASEizRySJLw6KbKiZkQ1jBNhsmVwGmaeo5ATPnQRUNccTJiIYI4
5opOxPNLoCct44pqmQGsFP1awKbRg7pm2bz34W5OSh2uwe6LdGS1fC7ctwTnTuFb
Xhiw5cjpjgujecE7I3y52XVi6pfqdoY5LVBDC3nBYq0H8Z71TCAcMTnhzwvzABFt
ty+erglcAxWwSH48yFaIO+zkajZZKtgtYj1QfBbZmSoacfnfLTKAvJGuJ+B7QVnb
yT0fHOecxrdwIc/gA1kV95wSuXslzVMz6X6WFGBlj1TyW8YGRfLvj2EtQxmIjTdY
Na2/u+vUr24iCHE2YDUrIMjI6gOp1xxS1BurG5Xhr3/XrBzchXsA64qPZ+if6MiY
V/5Id+y7ZEEI3x8eSB2TF+/NYD54gXFgmKGGP7IVYFhTmhJ3lMUB6wKM0nMencdw
3FUvPAUwFp9GZy5IIjvhjWgo28a6VH7SFfEd9dG8rsmHw+q+X1dGIRPRxFZZvRIe
hfEY+wseJTYC9lqshiaDeL2Yj0yODPn0aPFyujGW1BYLqtop9glCUMlNpfukdIrO
bINk+NbD8sUx1XojHm8aCCku5hQixoduFpcNrjAQTiTZbgR7qjbkV+yIMxhv8Cpv
ufmb3Fp7xMZQhgGY8OWlS9We1gIU7t6GiwKVjNsEYArNb+7dR8i3KYUoW7vM1v8N
qQoYqWbwMHb+JF4USMPBnVl4y3Dr1JHuEuIpCHzPD0HePgLpZMRqRu+RN1LTreDj
evIMcu5kmnrrS5sB0jOTERccxxWdMpumsvRP61I5j+sVzjFgElUfUzeVw9CxlYxb
pfmbvsIQA+GVF+Sfp3TbimnD/UMfpjR6jb0+hGh6HBZWirjUezp0yUSNSyfMtz7G
8zLpaqj6zwwPHsDWqL2itBLCAXLRdta4gDonXKT09whVA7fu+81yaMJQoF1LS4br
DKiOrserFWP0pX1h6+mHbghVXxZUTkPBE3xS0ZFZteWxH10w8O2G6OAVHOs+v3bk
SM+NvSoX0bdFLDz5ey9w+MtP4ouqwKfafGw0eoXCK3wm+8LzyJbFzdXHj9bP9DU2
N5Fw7KBqXWH0w+HTDx/SL3/oUAIGIBL4qna+7pwg7gzCHYRy2bX39b1XojCYojFX
qrg0vRJL58aL6EtK6tsxdGHFzRsxQvU2P+aRnaYG2LdyctGBQLF113W6+0XvrgeD
Lslxhx74TmQJTsdwwRRY7XrAcIPqoXqS1D5PA/pM9F01VGQoAYcoODRSk5z3hed4
lWJVxo7cWVaq5imVyl05evS4e4PqE8BCAYuaa7ETrjO39yz4XHoZVmUaoYuYUdOU
ceiRQZTkDeeiw7XIHV5peqau21QwLP1OzVW7nXLO2TVxjQihZ6tx9CxOeUOunvdz
JQLwDrf7CAWhLs2/zgc1CJ4yLfEORSg8/B8/B4TqytL460uABnVKaTmtZcWminq+
FuatrwO9sGKK0drpQ+/gUqTYpV+FJt3i1v78DdXtsEmQeqZFdhNQmfE7Jj5gChqY
S5tNmahiQcRtq7kCTHvRwV9eZdJHkc8igbi2ceSc/rmk0TlJYPXMLNub5HDmnAVz
nPY9LpQdHur9QppuxopLpoZ8q5Bsvioaco/kSR2YyO3yD6gU4Zis72mHSXr74/wT
p90WFJPh6y37nRerGobcl/ULhCsSskttOEZ00CYjpIIKMqJWnQuu9qkjpSq3necU
5DF6JFhlwkDtJ0bY5fKH/87C0heMQJjY5MmEJYJTnDvpOkqZsu53zURX/eI2eqoX
iaSwEvF/QSuozFkVnhq/XwnVR1Mi1WHSvb4mZpBtOFGpyyvgThb5ZRGNrEX9U1qe
dJIau0RSU2GYSEuV6QYSjq4VS4W3Hx27syxF4xaChpjPNww5HuKG8ixfDaxGp+lM
JL4G7w85MwhAV6wo90OHdQfNcRAcZtpgVSH5usp2DhtxSttRVjzeURw3O/43JmWc
I/7r6ZD6R7fiOM8jskRVp766WfMQGwTVn1VusHDdABUUTYiYEmtK9/fnMASUUtbs
QZ1MqpGl7RMoIBByaS4m3hsUYZ3L3UbljAFxGF2JSwuW6A9AbnFlKN03VRhZ17ts
tMMZCBnJF8P5BroaB719G8cdq01XOGTFcdCtoF4UzEdubfU1VcUsRZgcDxobAFrU
g8UHtKZrmsamIxHS/7/yYTPlxIza+kNcT8GAn6hYtaPbx4R88EHOcqC9YPCSxOHn
uj0USNCirraeMgoZNyiwof2V754MpnwpdEVqaqLrurYDlOUFAE8SRSm7OgL0l1zd
nSDxn/5He8NEGrZFPYBT2vYtzhhDFC6FqsPIJcq/PM1mbVN5llUFcAc7XPZwkJdn
/guM+bPrS5uFt93FfHaYfTNAaS+t5uLsduwh2wjvI+YmT23bt6CS0iPmhYiCzf1I
gFI7juQWR9sA+QUz739zLrqxPR/8R8jgv/kBRkX0XdTTiQ/xOlG9GhfuUnjEFvI/
IziZLt7A5S6ASx0ntnAcaeGMNFmQYwt0xsT4erDQEAc80xphgBwhcuqPMnFfKTBz
rD1tEQmzAIuMPmR4xL/Nnaz6gQaR+2HcwLDLokwfr8OamxmNqJlRtKUGDjJ9bp/f
4ipHxfbHPgQRstVihZu4raMrznSBWIEPfh81d/tHspZoeVrYkJoimlcVdRxaupwp
ALpHhQgZcno8oA8pEuMJybVRgxr5Db7uZZDhZ2Q8mZM5Zrgfsb8y0NUx+vReYZRc
3yzYQ2k0aKxVlJpY4gw0NO7+pujbYoPwmqYr1GFSqGMLiIT+6ucB4fpiIwWeTDCD
HZKMIg9h6wL6uomwG2M54C9FvbLYZi7wX2F0h++LK9H89zBPiqUQzUFKugNU2T/M
jB6XWpZFYDVZVa7bZb/frz/rQ82Sv9+AaZp1LBL5Ix0hxESrTfMMujtR6h1sMrAC
TjFTceoovtMo+W/6/8TafepRmoAIXsvdFT9sOItOHVwngMEguOPzEcAXk4xuqYY3
Qr5ISrYZhOYICvDC9VwXWxtubBdHMCddyvBioEi/BHm7lRQRCL7do+HTXPG8Bptz
g0EDHfyfkgoEDN8petnzMy4R4MT98aJChpNQSTghstMIXpQK3day3wSR4pp8u++Q
dffTkLwJaOmBZ311XdlgZJfqkR1Fer6CjYL/3qQNYPXUD9zgcraFLvSX8li3xAGr
Eflp+hbhdHhptaU3UcMfVxobFSWmkpw2+nKeouLbAy3ju4tVbxt/ULux/VSDjFyB
3X3gCOn4m3oJlOSuFBbAb/G3DxMY135ieYbJgW8BesH8FsZwN2ot7E0zpC9F0jup
jJ3XaKQAJH1LEdyjEIWIhE0DrdNXZvUhYKR1QSkDQc+NmycxYf5YnEBk/2xWwn9S
lVda7Upe1U3X63ylvy9zRDKOmw0c/l0BFMQ0NUL9tWpubDCOKTs8IKOppurKiZJ8
kvi1z3hIs6RQhDZZTPPnpmY0bGmPoIj/zusDKuC5xpMm9DcrUfaNoiPOMk9cIBSZ
U4eni2ClT59KtGjbIwIGVjXL4CR7qo42/TKNqogEEpGSX4rLEHO1S7UO1ci/TxcD
NZnbjbrtCAWHOcTpnQ3ee2lW6q4PlOl5CJeUU7t6B/WkBkGyIjp7iZRL0UX53EP+
z3vnn91ogrz1TvDvlhuosrKZ6lCcxeJ/322C+iYprft/5Vxdpa+BIyGx1kOQihlC
8y+LnJu7Jmxz8Bi9k9wFzsccwvsJIkYBbzxVa7WNQE2Y3K7OHIZmA3qYpkBzv8gI
3JofJGqBDINbuw0ZkxV1J8ihMnG8XYoF1wTtPl14x2BLKkI8BZAJDowiLkamao32
V0fJxdFBORLj8wQOn8xkvd+HNPNKUnvJLfnddKm8gNTmVQjMa6nHq9xKQ4RF0yXY
Tpb06UutXCTI9EX7TX1kC42BTQf2rR/AMEElqyjWe9A7VHA7Th9uUhhprUyETo/S
SlKLYylA/vTeRTm4dWDrgnDnmQQGYL/I3rAoDJ8tOojuOfR8RAzkHsWeyanJI4iX
V3P8HxpzamDgqVYTAXBNLbYpKy5N8kjoSs3KgwOPf1IA0qT5ek92uzkyl/pdhFE/
AQ+copYseBgnEQ6PxBg9dImAuwUo1pXQsfQ/va5/ak+z5KiGJY+lqf124iITceO0
hNaN8tglFP4y8yUkSl5b3JTxq14J4SqVVnKO3LKv30QsSyeFJAm7tYTzmZR+lH/G
yg0I96v3DI6MRBbJBiC2wJvQf+x6u8WzMEzLqMt1RjpUTrSpWDZKzjhqtOL6oZQj
lPkQkh9FIlJLrQ+/S+/NfIJlSrKur5LNKJmqtuSJG/bsGziioJOOJ0LOB26nu17Z
oDDStZ8FuWeJdIVMcV5sTWNpAKD0aZpWu4bwP86/dmcM4N2OdfNQ06rf7Q5zXlDo
N/rAK8zpAxMk8hprbiys2NBfdarW/5vCx6Inm2S5ZIqvHdOFZKMZ6amaTXz7J5gI
UhAOagYbrAKoIBnhq76g0JHUMvDcIYtFNAE5/4fB0B554aOvwHeKKa3cisDQkpou
MCDBXdMpIOe27BDDnxNYrOiJ1W72jSQ1hwSb4CgZPuSQKTF3UOu4DRO7AibEXlAS
kJRP9nx/myfmI5iw5NXrbRWs5PBzh/qTXi0cmS1TQ0V868A5mMwhY50eKZymQx7L
0n2LueWFW7XUbYy6I8dYhuwHWj3tVktf60/G/wPLq8YMqwb443XkBsmCpzrxbcYi
tFnwv3eAcdNZ4KiIeKIFgdX5Bj+PnP5ESwVzTP4YnTEEukwGtroNYodeL3I2dUaS
liZwAfrmbebR/aUPHHtUK6a4jqo4y1XWtCydbKLK9F0K14voYJmBzhqwsapukShG
UlEPWIb6gBo+RWTt/Eal/N5789nnWiA+8/cgh2cg/1TPeYGkYw1Pssh+Y4DlBNZD
LjZsNvjd++PyG9VJ1Eaea5SYyUIUKzyfBwPpnCfEOnh58Sx3YDXbkrlszzwT1FpA
Y03bsNxSPyBoh0CBu0SI3zxxiqrwe11fEWZ8HMr3iK/xIqRT8LJQ6SYsym4jMDNT
uHyDmgnM+4DgmrdZN0YubCUoRWGhq4nYSG833mHjq0qX4enS9L+P+z+rEus2razp
txPikbkoJuR3msIGOcUiIaDa5TSx1NVA0bRs1sftfuKupCOzQju4NM6JG/r2sNa5
QGiFVRfozXUk7wQWSCK0w+5JfB/I0Qk+7NDpF6pYZxsSbqEgMOaHJ9bMJeBrLNXQ
ErRvTa/MBh+JUI4Vvd/iO9OhWHkQyyDl31JCxrRVltvj2+wggwoEk+b5JJXzNAha
TkKi0qVrGQ36KUSaQm+GAmswkY+bZAxea7WH/RhfMlvOLLpZF4hPAPo/11m8ZlZk
IoEJwjKXkFmI+ZH85YDTosYmUieRJk+AlrWTzi2+YAa8kXL6eZQ6VmXtuWBmR7NU
XvfWTYrkAdFpTXPY9UG1tQ5aIE36355U43hWV6HHIxN5JuJkstZBfgcLVQALv2/i
8uU5FHKba2nlo77ralz4ekfEbPOfRvY7iaSWY0PjemDOiraEgCk5VBp3XYhBosr0
naC/DHxZ8ohIiqOtf6DbqL1GD959kMXuroBix8wgKVhImli9MtkMUEmyZCZERKmV
YxGKOYAqybO8B8CtxtugtaV/nSRJZ3FrJSkw8+4R9qKMyT3CxgyocezOwWU5ek9p
5KkaEQAXFavSqyQnms+oZlLPUYPbEbokXyIBoQH0U4tJOLnpLz6JRLuQd/enMs01
3X8q0D1BILCNhqc37qi2UeRozcDxazfEpaiT4+m+e/ix8s9CBxte8fdalvnci2Hq
cdeR2d7xo8qvQPacvr1wWfGD4jm2k7sHenL4JZAkMmYSmVQm+u+WzrEy10q/Pa8w
WcXxHfBkIqtvQY9TxnhEV3iWRQn3AF2imhYtF9qHBozGRLvEbha5Zs2Bu6WAFhOy
Yw4OCBRTCWwIprU5OHpve23B+ggXFvEySWDOvXk0froLNTQJ73Bo5iezwINTq+5k
2NE1eFeYjM/1JBvYUHWBJ3qow2UoV82FLadvsTKJoQoqLalD9LWJoK0TMxa47hD3
sDpUqexzyRqhm5uwzuxHLDEIQiKWzw+LOOzz4C13CCq1Ecepkjf7mLsjlJZi+XS4
TH8TcTa0gCX9mzyPL88NRzw1RysyvpdD+8vFMYrLARa6sQzeukCNlnXxWTeyAx7U
R0bSFO3hsLCd3dPX5AR3PFbs5+V7zrXicJJyXsLIO9jl8Ikt7KdGKyRp0bPBUqwz
f1qCIOhl7eWOkTsn4oiQZSEAWf3KlqF2zPKR+FYJggfxkoxIo8x2L1ML0B0V6h8Y
rgXcGEKPImGQ75zg3cq6uI/ELYNKYET1G56sOqs+oqfWHSreXVbn2Vjki1XzC0A4
AvfW1gVbCTx+57hYdQH13fjrc0CAW6059uyF/h5IjAI2hWeZmce/bg2FLg111kyt
6mXuF4D9wALYzz44hCP+wjbBhtrLrh2xlzgFjiJ0TsW1o5aL7RNNiaMN6x4SkxE4
3Gu83BLWKdWCKh3KQHlFmWj5N6DktG46bF0iuinDEO43lcvGAiw4NcFvfAsgMYXq
QqZn8MeVA90Q9PvpbJ1z0aVZk6EFq/e25aPhMRZAg/u1ndDYI8c9GzHGWg1bs2Qu
8dnTKUR9Z4sM4uvlWKsznoXB4PiOeunq9KVUSvohcvQqqpjueWxH87AXUUTfNDXO
0pf2jWXQO6U3sBxGhgNbCsQbEV2YeWfN6Lmfc6OS87nES093HFXGNXbMvUObIW+E
2HICrA4NOdvvnOjB/JN6Bz03xhukpHJylVtKr8/aundKoSA/BJ1bzij0/u8tCeEC
sXQt4artX9pxeIHjaBEdF/7tTAXCWBwTuAdtYvGW3BFRZD1UJmKtZeHw/ytX6aGF
GHpHhtjmS45zX+u/s4X/MRQQiKxiXYjfxPGqE5TJcWv5aFLgDEL2vdWoTex+vcvk
RKyrIl87bE8s9y4OHYTHyCw991vGDfW+XdVLo07/X8Ukw38OXNHF7cRRGoFeO6zb
7PKh1gaDPwJ8dUH5K6bUIeenavOldWxK/AS4j7NTr5jgXH7kq/LEeIarO72xy0Qd
EvcIM7LN64wyTruNE7m5OQxgH+gkNGRSqQTx+uv/EAkAXyoTRzs9HQDY+nydIzIq
X8IU7s2flGtbwZ9rEGgQ7Sp437Un7ao5Y4Xr7UFcpor5D9AM0K8Vr4kI5O6pnjsT
02lm0WGmbvtlu0RJ2dUpylmyZoqlGIZycPTHBsTIlh8VBZ9tg3bffI+e9duVgBR6
RQNuf868Pcgll3gaCR3ZcTvDQy+SV0rThgv77HfjXz7DD85oKQG5nWrXO5DhFa6Y
c/KD5wWH3Bmer9Bz4QB62WBqk5dewZ1ki/3AKcn3oGawmCWcn0/z4CZLvbd1cmE2
6nbLfTWqzfl/trAPZAA1teYaDTtaKBYoZejOTBw08LwMW3YiBVMg8qCjtHwKBJjX
ljlnZf98R2ORze2wwlRivDyBdHEzC6kyirwF1UovbLiNcuN3Oy2MAZngLldVC66/
aGTkiuuxmighEavC5fX4sEw6n8pofTx/YIO2q0qygT2Nhw4ECloAmmlCOaCxtBzl
3ztJPJtjH4DbZlAdWDwHGCKHJf4YV1Tnvm3sLriKgSM/pqURLGkbcXSlXtmc55XO
W4wJUyHtKb9wTHbovvnSx2erdY+LSJYGHjgucrJw6igTt17J7UDyedcR54cBqapO
sly5a/DDV6kVnEyY8u4MdQj6BIF6zsBnPomL9FiR/7JIWiZTxRjjyw7ApyHXeGji
b0PIOchsqI3QAUMNAL4uV2Q2ZFj3dhm1XOC6qN4OLhrPYJgvyQSRSZoxVuLgel4c
WRyM48rWnyYSKw0CbJ7jyAMyEb1UzJpxQcvIjL8xn2D45VUUvp3/JkBXeB3ZX8vQ
OYPsHIHVpkDWTN7qZ+4j0qLdQDiHx91s219PO1aO9efUmAXVGGIcaP9WQvs2VV11
mwZ+Ian/usUqe8Kt26o4Xm3gHwZQWBNSUy8+ez4rU1ljBWkOLVVMmhyr5h6As5ps
QWTv5p2O1WWl+3eSpfTnze8FMwfkD7e1bnzN1LOFJEIYEJ4ffncAcFZgiPDnaWZX
D362GY2Vwtx3CR/+zuFejNnLsPlmgsQ42miqido6jqwnDIv7AwFPepkZ0ObAt5XX
HGqmQO7WVi3vjXKzg54eqLngTGw7NtgHNBAjPXHL/w5BWEx+IidtH133MPEIAXUb
YVzYzuWkpxdoYrzLsQGtvNQSrGFSvxpgCY5yyAGBeSwTiiI+Mk24ycsbqdege99G
3dAmWGL+29VJZuUPUcXz7Ga+F+8TO0YZZ6UeFBwjJgK6awwd8Bl+5dcplzoxjH4Z
GcxtZeOoqFhen4PJGNH/9mTtkOtBe+l2aBrOxSr19vKIJAeRZ0Ktv9T64JO7NaZH
bXWqqAZKt3UmrEEIARwYngzrh1YNh/NvS68y1shwwwRyt9EQh92bw1XBblGfHaG4
rijJppez2PIw03Nmy2TePVk6iJWXJmaDqmXOI97tSbpC0nWhFLWrOzqY2Myuui2E
uIpyVhdyMT0AYE5PI9OJqtbEnCPmX0qq6mOigKVS6l0OtWFAmc4vzDWhVrQhNSMu
2Ydp7w2UHc8IIrcJIEkhiB2gtm87w3o4PzTBbfnE5QItZl6ugTeN3vdKxBZT143h
Q9VZX5AX/3JxZCl7XDIBdcwTrXBM3d8w39mgdZREL89L0Oa6aqF769d2YKy9JARg
NP31kOMvEfrLVBwkeGFVHxwIBZOgoeabdkt4dw0vVMi47tQE5Asxf1H2DafEmjBs
Ga9pAClOev9TqeKsTwkttBizHNzKOMv51wxhARg+YA62tJPTBfAfqme27HnnomkE
Eo4ADGoCuffZxLSQSX7AX6ZZQWvqc9obg9IIQVzS5SSQi2zO5CmNd2qJtJWUBqHC
xjcCI6MFYbMLQiu/kc2Lmn3RQ5/GE6SBn6F9/IoFz1PJzOt7d2mjphkJ2J1E/ODZ
4P4G+6h2M18NcK04HPfE44iMD09jownkRk5P5XUV7iEAgTCOFv56sZklNM7DOmZL
Hb3Gh4KK1uPrO4U7jbscM3iWmfFJDbeVCvja/N3Ys8dJwQr5TdAt9Z5maIcv8A+p
qq3RPINDVzmDCzNtRTYQGOo/GNCDm38t/cHHnAdo9LjNdO9rOHlkEZ3RW7JzxG7b
uPs/svaUJLSBBVDpOexoLmYM/EWzcgV20MFyr9oLTBs5RUZsCD0JVgX7nnNaOZlJ
DglBT9I/iiWEsaKdqiejU2muU9l/DVld5BkPR8vUm0rxz/ZBTJ7sor4oR9JpSmU2
fES7jIGe/lhlSAFeRSnndHtVdGKi3MalK5EArYFg4c7hOp5TwYDAznODkVm+Q44W
9xiQNB+iKrW2fD59ZWAPBExDqqnJ7JfrCOCkl4MurX8advRgjNsj4t+Hi33WLaiS
gXOQkD9Cr8iylbReRmUTpRXN2vm6wKNO9QPVVa9BixNV6t1hxRc5bP9EWKB1N6uI
K/obGD2xsocZ7sYUWYV64JYWuDhdm69HcF0klTc5l5s+p9sg1IrkB9RgpgNc3VF3
iBJ8oF4LnyAoU7pIslq4NVk86SNJqaPE3irKUV4gsf5ABcYMD40WJP6vXbdrjul3
JIoHhLsYzOgBPldp11LQGITwPRMpiYEcOfLb1BVHOi7NwyD2UqyVSdSUrp0shyuS
DUkqGGWuqJCFChQFM2O9JeVqpBgHAiBqL35kPAAEGEXMk7MHr+pE+tOc4fxoVcyO
LaVLmm3PBl7JnLrta/NtQbXaHZ8Gvdz7ei3f+7u9pjhiUXxHtgpkH8HCAQzC2ivI
ICCkWMwm6EOCiLzw4l/93a/WM+ZwrwUxNIuadOJfAuzHRvEwoY3k3rmtSagYlxdu
o9tSbTIgW5neTUW3WeB9QJODeugfN9KcIcc4w5aAJbgUMoeA0q1MkkcjIqR6IfDJ
mfTISk6lVx8NBiKftK2tsEKWI+V4E87quc2GqmSKHweKIba6fCE5Rf+d5FuWwk5m
uWbqlNkKPvYTDAwripLou4XC0kpL9hKJoylLVS6fnZa6hWZkIjbrI0H2rnINrJWF
fl7PWtLxHDXg0DGS1rSaG9o6r79v4KT15oPETyZNmR1JGagAYNauG1dneCiURqV6
2GU2rVYhDwuhanQ8In/B3dPkiS77p8NgHxJ1oj7keRZNG8zKP9ua3r0w4xUO7Jt+
Yy2ibWnaNpy6s7lx7iOrCKHpnib1LZvFmlgDstkjX3KZbybKu6CgQhdI7GpJ+1uT
HSxdKaLQhyhXKmPpyt+0IQGuRV4UOMh7IQ7+I4jU9GOaqycPu6hsNWkoO7oLv6oj
vnOqSY6vhedUjbkI76o25C9HMPYB2ewRMOMKVjGFX1awfu46Oy3AIO1QkXNn7kwo
zuLgWVjvf1TyIut+ga5iFsjQahNLtZElTZ3tCY4ICrEU/JU1UAGKtDHMifSKZ2Dm
3QK0Vps+w6aY+7zrp6kk6OmeLsWSgR2/SMurSQykLk0iqh4t3zlry8l4qaFpOmw9
vrkcITjQPDmPvivtPz2rk3gsbMvDnieHpedcxpxbvkwvS4Owi50HK0+NPTX9dVzE
9MRs7yldNsF0kFEesNOYd6atXb9IJ9P97zFEvvIwrRfdZI27NRosEQ+1X0umCqF/
ByxLabrw196IgONWyvnVznSf1elnzIiqR2vdffxTxSG9dC3LqNdL2ARG2j+DbXVe
4b2aYxcr4x1NB4eDtE9xBLMJdTnk2KnFRTzFgXbl9+8l7orMNOJEOtMuWePXEskM
CeU5wIxjTT42Gpwp5YFSgVhXMMM4XHpSZ0+7NnN2X3/RWdW8Z+NjE0XP9RPMaJ7c
+1Yco54wDOw3PGxU30Ac9efxp4QYl/vqQGr4hUH5iOu00w3QqCiTc5zIEQF5WKrd
G1mLuoM6wjBgXPJc0/22oFCkv36LI6pVwftjMrLfpzKL7riAxUGwGGtoZ3dIsMfJ
PfYhzW62z1I9tRq3p0TnFnVgMAv69HBIZ673ZK4RmlbkpM1sIqfOehaSA89IlgVl
SfirsclQBS0inlGj32qpqHCiqt+wwsLeScj9rgQ5BtSo9S9wYkqPNk+TQGA0Ru9s
gNZ+unzoKm3bGwOfMITxfZWTXfHm2ax81pnRkJd/0FFPJn/Id0VrJ8AHaHeieHye
U8UfAkuvqYdqj9RFGtnKdYy3X9GJZdIv9MsBzQxcvoe0enhQC+NBSpqTJV8/RkGH
NofMMm9Rjveyfz18GYs4x2hEdJmRehyZy3XoZPpdJ1rkKDWLnLXaotYtKayMTCTx
FIWOOst6oe1TpxoWS0+oTnzSwLZ24ygAF8OOHp93h1tSYExE8LnXEWHM9MT9LN6t
RT9QcDxJY4AoRJmFKJxgZQhWWlRmHBcZ0PVpt9Pf7bPGa/XkrSMWVlLKmXECXPgM
bGu8Jvr2l73fI4QcAbVrd50daTxWyBmkU5k/JQkLOfq/Cr186ndBldkucs8k20tj
N9uG1ID1waD8zlkgBsXfwh3JfMZ5efUVgs7MBVV56ijzQM5/ul+ypEpLcTw/fge5
SB5nqW64/e+hli7qBD70Ur2cLIxcXyZT6p0lZqNfqzdUKALpB+yIAQmajMyfuyMP
M04jnridfC9RchMpSEGq/Wtxx9lJ+05HYPNckZDSsJQJ1Bq4+SNR8KgQgP7CRZMh
9R1mPlfaY8mpHDX7mds9+lxh3rLlBKS0Nwo8wucr8guhzDoQQi9rG4gCg0FFGq8j
ALtfYL/ch0Kw067e3zRFa0AAB8oteuFNW/BSlKsMNCBU1WoBmQqa2iqs1ainjYEo
63dhRyQydr/2olEekW4I0x3gTJvNhRz6yCA6LmZS1tHSe0r78JYiLyURIawhJ+5k
o9WVIJ609d5aL6O7GNI+i4HexVpth4A13vCFPLMR1uZsFLd1a1VkicrYFhBFIHlb
9gCP2s2nZdmeFhIDuAIX8DGKyqQpNqHGX9bMiDvfk6odM33MKjaFxEyNrq05VkQF
G832+3ks86bkqU28zHy5fF4p9zwJ80wiyvanA5yndFLxduJAggkpWi2+eDTFDLoz
tggLOiCOvcA8GefWMarrUWlv+u+VgSoRZoFA5UBk821dL6PlIgG1cqPfA9MmXDAE
3d2NYWd7IAgQdGuctM8t87BkNVLYISa/hoHo1q8qlIoGfd/A5pwr6YXuXWF1GNxH
/2GQQquVT7pAI5QfE3mMWjVerKo2DGCXCoaSz8lsFjEuMCy6geo/WH93nL2fLWQ9
hPcKDhs0U/a7Y5kSX89bgTfzk6odmmzTViCAC2wQ4fFWxYXEVauyctvFNPN45/2p
Elu7e9BReVl4z5N0bkBfiqmQJs/OY07C2NtACHjLsGz3o+TKULmKrBsTbxrB2eIy
x4taU21JWARvmEYJsvH/xaS7C9u++DaOcN+dug6T+fQp3kHe1prGm/nN0/xIS2mb
OadVfUUj76uQU45g7iE2EiU/ruDf6NvbWLoxq6wIEsInZjs1mMq/fdA7sa/weZNK
qiThAppVjzmRZvLupkHtVMcQz7tLHIbiozKfpANded5NEPv8+qDkMT5GXDceaUeA
UI90SVVCIVZtjKL1r6vgBn+NSVdnfI2SRLyRtH6FkJuajk6CCQoQI2/ZNh/Co1KG
x+gP/qtiq47GVZWATuPagAhmWNLVa7cCK5mibXTLN4XbmtDlOJgx9WWdOE7Ct5FD
+ArNzddHxnfwL34amNX2qT0WpzaESQHfmjnayVvoI4RJd2Zl499pPqz4OiHY7THM
4lXBZ5YEDhLnu4BCeqgxPX9WH+HcvUItvdNduxLpQAsoo0GvZ/1zvFpwReaPqna9
nizC3fZsImL4Qv5yBHel05t7FZL6z9hM5cVGOQZIN9tDqpRBOu7c40qVeiBJcWhC
SYqeOdOJ5dX/fgQJZQnkzqj5+UVuxvqUDKzWKVkuys876QV5WzyfjEpyOizxNSvX
T0gxVM4n3P15J7N5WRixnho0xFfIzhmHNCAohclgMTSaSL3iaQmbMcqooJX09JBu
lcvKLWAZRs0cLBoKMoKuC48BlaW6rmEuhjoj92G01BYKGe6a2CihYuEab95EUyh8
rZU5iZ1awY9qGIryTZQdqhGNmh0IkehPPayFLG2wZMSrJr0aQQSrZ9sfHIeWRlun
Wi38RnCO0kIRgSanQZs2xZChdWlqdK58abA4hKNIDbOqwqO0hQizGgaQ+U1MOOkg
sIYE7osdQYL6ukCATJ/CHaGsTUaBxC4geXcEr99zBCkK10RkXj3fRRYEpDiDlMT2
/fWZVGuHal/wNgNXWALVWRijZyoRZCAXWXjvLuqGQ14OcxkGZZzxhDNAxn+phU9O
hP5o5vHIJUT92opw3KZbcppXj8GRhpPJbpZIWFFhbo31gmj/kBmQwv4v4M/MiXqS
dEKR7tjAguT1UcqpPgLvLwaAzl4Kbxny1oYM1Q3jY3WLftCmBDGjBJ+uZA4F86VU
O/6+ASQQDQGEIaDlcBeSvrgNgxCkkb6cB5Y7si9rKUHHT8VBTBtq88fkp/+jgvpF
JM6C6kAFkIO0QecV7Crle7N26ki1cIFrt3fnHNqhLgj1K8bf9ret0kH6SEJlO4ty
NmiUAXR/XomdNFjiobH5rKoHxCCzq3OZe1qW4BTMzGG2w/zwDvY1MzmlZX6hoZZH
VQuxQu0J+gQbfmJDk2cec8s/IywJZ8PxBXefFkSxSZFp1mcGpE8YE0u4b2drpCvS
Hhv2/+RVQ++1doi6qNjBKx1Vf6cWDS5o92uZKCC5G6sHYjtNdT45NKWRycPJlRPH
bfdRq0W5kv9SNleF9vq3PNhivbudxlKMkNed/E97RNfggz+I0iFNjPHYzkGmMTkG
ltfEM71ipjFv6vKRJ8IsF1D0Koilmz8FpG6hpJ74C19aq3pbwOWsTWW7HC+iU5Gt
01SQSIhURIdAVlh8HikILLxcrKehmI/PEOTryct5Q7cGH3x9MTYDC31HkX/uW2Qc
9ShwjTvvUMKK1WmYY9D6aPaMIOcus++lUVzF8qFJJYAUVs8158+gvQVI3puYcASB
oqfwuyVilZm4B1DASFemRz17MoHucZ5WjJjxz1u1UM38bH2CZIpQ3SJoi4OVNzMX
XwN50j4hfS180SkA/ZbOKfUeN7dvfM01jXZnoiZJaBed1k/FVHUFhqpZnz3RFXDe
gClRwlU8JRDdUghfAcHviBhIWcCo0B2uiNiMzxjI24+H+G2EjfiS/O+tPOYo1IT2
eATQt0ousRJ5m8V2/imKRN2BU7q/B8pQX2+LUCVtYBnpjL2uNCHirUaSu1EMpE/1
NcMuLA4hSD62x0j9oNYt+sIn+2V9oqwF/fOq3XZSnO61xP+tHA4KEBoFGACEbUyd
w5jc2dPl4Y6zGx4V7mr01GGAqQjsgBgG43zX131nTmkbHpYGbj60Z7/NnGO7OqD0
/dw0f7WNIrRGTM9QKWNJ8NKvkM5vTpg1rthMM4OsJ3Uifa1ZP6ZIvga0o/RKIzKK
or71ogyuoAHP/CEO8t2pn672p9FPpgMy5JjwRDSqLZL/F04idhIwBcIRvG1V/Ew8
ayx6bJsw5TZ5aCpDFRCM5SjP8bFyU61/fOUBtPSeEAwZfn4JRHnvrjRSbBYDDiPV
b2yfjS0ygSstwucv59iKHka7F2S7XwImBkG0g8kqYmtEF76eLcQPQyOQa6bHr3Zu
KkWEXPWGVA0cRdc+QMAqx4DEZh59auim6QM35pBYbeIZqFQSf86dF+Vg9zhuhGwl
hNbk7WeV8+W8x3xDimO1b/noZ9ldXY1UWF0vZqi0nuoIrddig1xABNBwRwdzQmV3
9tehQHb3KQ2d4h3/RZN2ngn7vLjSIAhnCP1ebZ9jjCnnMFKkhBtvdgE1MPOYWsMy
XPwgQPIgMbvW577PXNbb1XhaC0th1QNpH7eJVQv9M5+Cd/A2MyMr+fXIeQhe/bMc
XIcaOJmYOvYYNVNfSGiUqJTx7vIU/ug/RX8UzmcVLxa1vpoeEYWy1r/m58pUiUJb
Zj+mvB1Yttd/kqUZPzbHlcJdXUyyFsbdz+l+crqe+LZDySTKBE7pTMngkLuxk5g+
WvUtkK6mbfiF92Ud2xnpskYQWi8VIkPTvVhnUr0xj2cVmt3sZyzEcUyhbLLh8qUI
iaiNmQgqUSrshvEZiGyCuCzcsg+xvUNbf7on9Wcyl+punsbax1dKc4/rkz7adEvm
vNDGsx2MdJ866jN5bWN/IOANror3H9b9fVd7dA9S546bxYhXGS/IRG0sWLjQTJKq
aKhM19J4KSRpxgCrdzbiflDEgGJTGS555bP/py/gCzohVh5IM1FscPyHIbIxS4Z0
LYRUORB5zx355DF3/DHG374YvkHimPW7ZHyL2xJGKbK4B3bnl/JWpTbKtTH00/Os
6am9fBcjUdqUORpx6Iy4ustCDt8Nj8pJaaYL8TgVjWycRfMBSKyQaBptfovmyQ0G
lLRUXuCPgKeyHK4c7++L/iejepXBKv0PVeBkyOQa54ZvszkEjleBxf/oKJDUycEa
4EdGGSPHpy/C0c5hrLQP49L76bUZVATlvD+/t3Qtk0v1IZgHucgKQZI159p0QLU5
0rd7E0FS8gj4D1Bo0a+Lb46kg/EmpSto9nEx43LSr1Yf2BFajgMpkoEY85B9jd9y
G1CllOXl8a9lFV22zxYgi24OR1SDKT/4bLRZy3nKXr2TcFe8siDcloJ/gmLNNqVC
FrXWaFNyxxoNh330Q/bozJy/FWCkpdltH/MzRRyrikzF0gQxlJkSHhNjTPF8DKeq
t03tMx+X+AKRnKMNEGqqOTwWoiNJxXdmIA5ExBHu/2XnhRiRKGrSqge6xu5THLwV
GiS5J49sAZVXg3KsyW6xhiMAWAiZMmNEdB3Yo/KV66rrcyUK+yA5vxGTdwJTkHns
8Z2Xhnjjr9W/mw1K6GGU9GoFXwQuKtyF6ivfPY7kSq8IBDp6KY26ph3TJpgtr/tJ
sU0guYotbfvpqozwzER9uV/QD1l/gbxfurTpc8hqAi2S8tpy/8hvjneD3RVkV6YF
OACYlgqz1IIBuwtLMt4/uLvZkJUQxrFgBajMOFALg96R+cWzACFdTjPWy2f9l6X1
cGhjsKRDZYH6KsGOgon5+P5/ecCHR0KVojAdKYsNkCai0JTbWRYvq7b7PD9mE0E9
vFUMxVUNmzLzOqo19TqXMVjIeRwZHQztCoFxl4MX+nFmnR799x3R+3nD2t2OJXFj
hWhrZ9u4bQtWTgA1XCfQAXLkcCEYnSyPDqrS2sG7EBXyIOQF4sc8ydEd/SsAk5Gq
AQWRqxF/NCz/3dRg9i7f4ErE83zuTfLSQZL3nO05snrcNxePObkGclBVmLA9PrDH
ZjNnmUx6JeZTv1B6ONnsoBkFbZjxHFwNrouCj5BQcDzG1bbSbzRRu7Mi7nyPOvbH
UY5G/jGgFLw61Wo6zWnLp694dy5Kerj+ThA7PG8G/htst5JBYafNhrKniUuOr4g6
NAPIEmPw9EEih0CGoVuhTG70D42zxdKtUBPz0gQIZi2gqocDgeV1uR4yiepNytHY
Hfwq8emogcg3F1fi1VWpIuk/coKMJjxpBoAedxd1quyUMMzmkH+Mqroy3EBeKsv8
ZOWKldEDXVqxNUVjhhAyWiSel9wVY4LEXT5QaTSEziU9jg6RAXkMcGoMa3GBXVWZ
eGOI8WRXHfobYVKWF+O7eeYej0NNxRcc73jD+fY8EUoK2awg9iqPJIrFESzcBfsc
mTkKzh0enH85PE13/b98rDszKB/CkgXBBwlqYCsk6I752txhUgUZvjrlmAb53mD1
4PNkJ4vRJniyhqYOoRzAKLBsEg7dV6pa2zfAFQdVAxi3zhguRQSlyWDaeWk6w/ao
93ra0R2OKMg48hIbmrDxAUO6Zxql1Ep3wO6kkOCby7Fhd68koX5HvWrlnz/sSkJK
IvumnlgGns8i8s6wCP/C/UNE0zHu+jzOmFS4qvS9MpIDrjo442qB7nnH/69LD19p
XVYWaX+zpDksQVX6nDEwe/xSvJ21LmrL1+E7SrmVeD7kGeH1s+Y3+kPwsf7+YKJ4
jOaam1MeLDTC3OVZvNK47Q6RhzqFkdzz4szzKlnUbSPJRoVhIqzEgs/nUGcIpi1D
Zje0/J6l0c3fcDOMxfMAz8zSMB0fBfgksVXyWMkcC+KKutXLSp3n/u+5MAjgNtvF
bUIp4i1/FnDFAOLh+XLdL2qZmgTz8HR5gY7gAcKe+27d1TdMAYtLuEuG/iPo90wG
LtrvIzYFWZWXxgXccaf2ie06KkbvVh1zhDsfa5/Q1tkKfDOCrfzWSAsdLIJjNNpC
pco228qQV7Pmd3JxcBc9Yh5YC54dmlqq7l0c+M6LKPS8SzUjEkx6CNntgppw9MAY
l5sR2P7rBhJZu+l10DSZtDYf6P4kHQyKJ4s+q/LKoa6IlD48xZLhX4jSUTfQ/G52
2s+cB+0SjSIavnO2nDsktLSIYgDfGi+88+mOI/bkD+r6USn/QEoCHSXZldw28XC/
UnBk4GLA7g+koY+ZtTOOL6xxgD0gEW2Vy0UQ835cP2eySd9IqiepUV4oMS2CYSF6
2YCzL5A0FY9Eatrq/UNIVhdGCvUDKaXL07X5iD4bFG3A6rBrw9f4h8tGySfxVAOy
j7MROv8zgEa9SZ5RfhiMNJJAvyEPnngg6t1wyPcfLQSn2wYRHDj66krUFYfoRp5e
sn1tbJ/JCIt2OrluWeZLyF5mVCZUPvqRfxd8y+dJOvGUcdZ8R4buxS0FaJn3NsPZ
lfxQh+IYQl5kjpiU39KjxhAuwJ8Y+QUSzyPSMSEeiReov4tSxaTt4V1ZQpJZiI4v
VDNZ7Gu4TLqpOdOMZFOZyA1l9vmz6Yg0RWfCuFLqqa4ZdgZ2rxl062WuOaCOKj8G
/7Gf5evkBN7UEkTV6Jvev+7eTFdzR7yZ7hQ+npc6JsCA3dHZ3AVD/p0PfArSR4XU
huI2mzXY6Sq0gakuDuxX9Ppi6dxh303CmWslddyUtI76sPgw6mWUou0j6ZqG4UUt
MM6TBlWJL7lGvYwh14e/dIByOOsjsDAfrBFYfqIgly8ljyP9SlIurFRDVsg9gO6S
budu+YYvEv3XnzQtOqMSGNxkpY88wqeJGkQHQNE6mmeyWA/B8WH2qqOtO6j40XZu
59ZpSrtkbw0tliwfMtsd/3bm/FU/VJQI/MGnz6NJ++AzE8Dk8kJ2y0vg9zh/xVgC
5kQ1KHLQJaXKPLuOSCKZ5HN3RHTHvEpWIAKvwekVOQKq7cxg1JVfM6q69Bk1yQRX
2D+mfloXZ0E+6ZiCDQ/ng+AaAAgw7iRV41xbc0oQ+XoWunAeRzkeLDTf0Cd5Ux9Z
MKN4RdQJYPLMpBZTUpAt0m6xBzgjtYWa6nmx/EXXLC5vhBUcBTxJTKxeftt1XLzg
bwXUp1uSQ78R9fZjdBlsBLg8+HoHHwo+pbM1jbLFAA7UeHRoHSmhO+/IJo1YBwVF
0WaqqizCZWbcAAB8LMAN73ItcO+WaZIDUlX2OTTSykbQ0yTqT22VNihds2xjo20s
I4lCz6jP89FNGZlzLppwW6Nh0n+x0lngirTAqZWGdjW3RQZK/yC0ZAZAKJwLYY5U
sZGfkvwQqRj1Th+yPoC0UzupAXOyxGjQOYz3hdtAPB4QjRqSGnKcHOW+v4EHgavp
GMd0uLJpCaYt/EnO70sHwh/uCWTsIZO+Z9vacEQl+uapl4GkwG6h9l5nBIJ/9fBc
rJxvyJqboHBvgw9NOvlEdrEO6lUd2mlBh8SZSOzIzkqCBTUaaJII8tzjKD5q0dNJ
zwgq1LaW+JdRwaN+YJEGPvP+3ObHfRrhN+DTeF+ta29SdzLdiaTuoA1zWP58YILC
YFF858V1ybUpRJKmGrPSrugECHOweOY3mROGNp5vTvdt83OZcSnX2xelgx16PAe1
VwpcHgIKMoLl3lMBwoPjMIMYeAXSBKLoA88NJCW1pQ1QK4WGbVJZV2uTx4uBs/Le
TkenrL1uU2HDNTYFR6pb+vztJPk85gaQ6De/+Qi+c80MVRtOHOdh71HNnhEAgSPr
6bQpw1qncEnUJbGbXVop/Rz9gVmy1oV9plRGgjpNTvOPKIoHCCfkhOZ6l+m7jv40
twQxOOX7jmT75AE9sq8DVMAM/NS0WmQGPCI6AIwiS++9xfDvlLnswJaTj75pfxT3
4fEtQgZEcdrhVU/RCmlyNGhmk4w3Jc4nlHZ4Fch82ZpZGB5ZvLHi36thIpdvsndm
+wuesEC5kkNq+3ZPzWYkRv/opA6rvSS7ZDhIlWFjnf+FrJp8NbX14lZbd1obdKOI
UC6bqIm47QSwVGSy8xYahfB3izTuNK5dlbO8NAfxJDgR+gtZZGBaLk78WSjhuFJb
yz+q8qqTIE6xD9THTiLX47NfVUUjGESd3fVbCuC/QgNekwD4gvgMKmHJEFRqX1uc
bBeM5B7Rg1O5TN7HViQkGQYV3VM+2ea23EjLvh+kabBTWGYW9Q6AJxRi44Pm+TGo
zEUm5YJY3oM4QzfmwvalXMtNJX7wBMJyuLpAOpk71pUxdKNkuctVfWDBTPKoRv/c
sAeFmrA3Fhx0I39hgHLIPWdFPG0nrZKNzrZ6rs+f8va5dojlyMmMDhtjUtPBD3OT
jDU6ohRwKlS+cSG5Rx6+692RvBUNFxR0vOOX0XUXo2cmwymbD/ecC0yTNDX07pqb
zx2yCHlBHyl/Gs+BipVv+YOcFyOWziHerQiA/26gyF7IB2uL1nlSuZzXsMQXpAnr
uMougI0gJy+WSScNjUH5BF/ytMByZO8w5+jzGToEh62LqT2w+YeWoaK89rkxHfJm
BEejAo2T9cuxkE5/djDeQR55N4MVMpLiQ39WAKWQE1RxdqlV1gxC8dWPKuZrzyCT
W8L9THypFjTtZT8uFbM03ZDImBHG9RrIdezgbYGJiugMpV37S83K6K0M3V/z3lfd
bZaZqKPF7jHvY/grMtGZzJTiR3brRQBI5zS/U2zENUBjMYrOfrurFnESBwuwGUfk
bvIav5zv4qlIaw1Eli/HWah6cCS2HnhyvPu4GxDGI2Kl+7tiBjfQ8c/uYDzPiLUy
4E0dVBS0sFkGLC9q0qTLnptOD47tuFxPhglWe+Cr8wKLAiKBv7Xka1DZYfIm6TcA
c2e172LQTYTf18dbKGk6smxUc7LT0NH9p3xpka9fDdjesV9eF4AJdY6WjAev1m64
BHkyrWFdA3Ew4C7DH3yMQm4dGl3a/4FQWkVXCYQsJCaHubc5z8wBVvvbZhkbiEdb
CMHBynoo04vnw53jzNxo2Sfarx2USoGX2i8xVgxYY8oJGdtUM0d9D7WohlDeuK35
oyQxzhM8KmhR9Q4WNyrv1HeCZOOmtjRC4VqujLuE1tI4gdolPdiBJasUqMIIPcJ9
KBQCFGSlEzNd5FZWEfOFNonU4q8T8XH7PsbOZsxu7DzPjW26aB4RReTlRUeBpgxG
0MCBWvTLGpHgRjSpOCG4f2LQq3eTetACcVDkJ5RVHUkyTAZlyImqed5vLPozCWuc
w8kbItdR5sx7Jl812/OXTzV7f7DVnFsl+uRokGBFcpkuUjAcXyWkSsecYIjW5Z0d
uNobicXxK/pRcDqE2m2cAVNcWSj9jkS3RaI+4MBN8zSgjaAEbTJOilwWY8hE8GN/
Cm2LXvSsINdIq9Ex0jirm6yF73SbcGK+9NisMQF8Iv6lKnyp7l5N60/6COf4xT2e
uXXyGS0EeF17WsryDZUXTCO0Z63DGGCYzC1YwWEaooKAMJVj1eH5t6uxSGyN76XU
G1JwvFrX7xfsMmKwy+G2QPsvO811M+LA4LgdBZz5kdlO1wVY53A1MOzOAIZmuGa9
0PA3b8A7E0ONVZZZWilMjTeSsSkn0p7XeDQql2g2zxMEuevj5mK91Ovims7Poh2v
yOqtuGRSmbktM33Yu+GlUrR4YjOTx/Upr7IPXUiFodMJ1s2ZhtotR1mOc8r5BE8t
gQi9UFngWEHrsVGZhyNe3QpRFU/yB7GYsfnEdWouaE88iz05hX9QN95MNAVObZgJ
em0lD5C/CiN+NX+8v8tdjXND/4iCvhpvH/VYESiuthCT5jiAiL9O+m9hhEiLAP5g
qyK13WCgQl5GT9NcTUd+7xmDx4JJXadYKpncSeBhHqrYzrBJsB8mGulHPiny4OyC
xmFPvwIwUGgysjmzxp4Di6Ebnb09xrG42ZlJMi2fagGsHwseFNyvXNqy+8JZftvj
UIGK8v1/xWCD+7zOBRU/TalCxDfMeyFH0uj8niZiQduljlt1fym2bHcjuDDV90Y2
0odbYYMBz60MsD9CtV0tBoGgRr8YNQd+U0vQj/3qDdrWMsrg+J10n1zUkk/GJzOE
TRLrz76dSK844IWvOS5ImJvZ5+Kd3Q+GCPgXcSUg3LFDBTrQdFRKFxZuzfDx5BQA
oqlYlPWG7sfExI+UciLy8xyW70wCObS5vSd4fZIKX2UvuI0rW5A/La6av4gmUGpW
KJGzRLKxczuGg5pNt6WGsbR/QoEH8xVsN6dSu2uPogH869Ay18baWeuvWDdVHq0I
pJZErFJ+m/W4ASqsNzQK3Zl08XkbVv8UfS40lTDNpS7526QOJKZFFq9x22gVO+LU
6A7rpTyNZIomY6JTqzPwaj0+vKXLop33DSBqJ2c48Q2UVEOqvKEkD8/pO1S/W++E
Wgods9nm3neKORJN69iq/hStC0A2EgB93zArKODKly769gcZGrPvCuSwoIBGb2u4
89mIqVFoWToVk7cPLfSgXOJxRXwCxXk+cVR2wCehMyiT1BvCJMwl+njxDrvqwwMz
Y1W+N4PlTnZ+7FHzsTYfad33SlEVlX/M7R9oI3Qd0D7kh3V42zHgHJQQUSo/qZOM
6gDj8T3e+hp5PeraFvETifCyBU+bNEcegd8LYhr2cM0T44EH4iy3xIIqp4tntsNv
WXuHLZCldEljqcgTIDTaNVjgPuRwNUbfkJt46Bi5FqDs16jPFJrgVNU/ydPxYHvw
dE0G8wrgjISqeo/84OfB8Jzcj0IOgh6VGI5AV+ZUEmybMkAuB5TaCbovuqZOxMRl
IzFTEOmIYRiY4vYBUIysQX3XsR/sTiH2R+pzr5UT2isa5AHS8DPQgeE2h8li9znP
yWWp6RGKW5/G4teK1q5bckE2Krsvoi/XFFlesasQAeACBFCs3Q/HHM3WywDjhrpx
GgYZNdKQ3Rt0QzNOb9/Goyzk5Ywzk3M2ZXbeniGfTz154Y/1e3Ft9rvh1d1tPn90
Z7pI3nWDbIDh4xYSEN2c5DLbVNUE8s6wQB/hC4R9q+iaZx2yHbNcpUAkbyk0bYwO
MMDD3CxJP7NVzuVOMi88rJHwyxDsoy6DZ1bjMdkvJDmUIv2I2b7Y81TwYyF+i0XW
K7A+fLE/WvA9ZVT7BgRw5j9l2r1ZVXe0S2NOtZCyZlxaOWMsLdO+lWoAv8pytLQQ
pEUGQr4cI64ZfD57x7BVr/s8sZ7EUp9tHFYXG0SJ0quNiEYfW3G/IGexo42w9b76
FjJn8Ciez8WrT7xneo4ENvLqdhfYLZSE7ADPvD6duFGUob54ZqhmOBUNV44YopNh
G+7nz20nubj59glUKI8eEYRS4JLtDsICiBhwIOl85OZ5cHOhKrf+Sqqk4oDnOW54
WN1XQcvYLeH2X6cttQyfK3Vz/fTP21CicLLVgO9P3OEbpqHkfe0ioNGNEgyPW502
3NSLxyQ7Z3LGTzRCBl1DBhwHc17ENKao1EUPfWtNwKojxBCZb+oFTL6QuWjCIvwm
6AT3UrSaVzE0/K8RgYtvLP6mJvxTJbGAuXkxODVbI18IexFWtpzPR0pv0RftzN+D
LJuRAIQ4226NvK6lcMhh0baK8UxdhBz6jKV23yCHLuaEmi493Qj1rW3KUd2rJeDp
Xmb3uaCXKnH1ha231MYINvtFdTGVYonku/h+CE+ZF7HSRpWwIV5KhZEsqipsn4TZ
gkB01zliJAz0ddXSeoAQXC/MOz2dsaTQTVQRy22mRA6UYeEiUEMDKc+UQU5lyai+
qyExz3n/TtPh2DvkndgTfBUP7U+fXgOLEpr2MCKirTYnmGALSB+41jG/z3VXGOpz
phq+LudPiHSS1mFKuIJR2R2fUc/n8CNXL9Jd+Ck4wiDM8DtIkFTDRxbKhuG7VQpl
PNRR1c1LW/uoNGNfIMnWtlSNuLRmRX7lv3Xnoy6KX8IpZhWN0IUU/E/BamK3OyCf
1Y2CrTC6VWiyUYebO9v3F/i2pGlQ/mfIrcYgq+cX1xoe5ERJgDdXYmxpvqrfu1Ft
bDr2gwOVqQRrO/bj2Kgp4DJySos5NG9KHB4VVDjQ7/ZaOTGyBSNSk9+Sy9MqX9g+
1FVGeICRwmTa4mE2hRPeo1p+4swpIQgDikW27A8oGCfvoFr4Aj8OQfVkBzvlV0jm
R7zcHRbWuZrWPSwOEOmRIYViVrcdvPPa6oreqNiSdwVICrayI1KWGSKR58a+yHqX
DkgYVWvkWYOv1SympSvf+mU0B0N0a4B97gkK4BNnGkR7Q27Lsetlh7co9qMleeSM
2eLMjUiYbGSFIbRuKJkM/jZ75OTOp5oSdewfx0hIQbHPuMGyM0vsxUTSdG0+dUq0
Z0I8TZAseoWtU7+fzABmOWy32ltxe1VlxT2SgmRAJszUTeZFx9pArr5I7gpoi/w3
TzCU+wAKui6SK+DbE+L4olyTK5JdO4N2d/0+cW8Uf4wj9Su33qUNiy59vvqq1/oZ
RrdJyzT679CjsYrDX81kkM5KyYlHsGVzikYLa7jwMn+iqgCkSXbgU1ZIK+tatlrw
0bChWmXJCjxHx1uGo3Foj8Q1qbaYSPEhmmlMev70CCcVOOPj7fg3NsMmM5rtKJeA
sfbdQ/C9aeY5PJdElEgrYbgqmO5mSVpLTVfB3uRPuNRiO3OQo/aqbUqaYme57o1R
VsgDQ09SRwXYTPOTtsEuiFj1tTLw2TWLNP80fjkqiQ51p927NIOZjmY9v4edl5JT
VSxCvpLVJv5KdnV5NyFUxaVBU+B4h1ndRckgnODTyUDpEP1pw8XdME8JtdEpvmcl
mB+0vSKdN7NurNcOjZwIblWQhd+8Z/7vqTj8WXl9op8U2x0MGK+PlEdJYs+z9fUb
a5xPfBlNPmB/uLspNEBrUKhqsgw9LJ5Lb/ze2brN7KljcM+dwmEW2oPC0RhOrxmP
fmxKIosjaOUpaATgqzyTk33Ua5AAyZI/HTwb/dyo2wkTjti9YmsXpoEhUw9AbH9m
E8tcaYj3M3UatzpXjtq7AeGULNa1O8O0B5XZFL2HJg7d0K0G0pQQMXIcGQvzl5A9
ovRq8+4N2qOLwcVHlnjprNFxdfSieESCyDNTZDCk1dQ6A//0nTjT+Fx/gf25csb+
yNTGb/zyD9kOecT1see0g6gqcd/XPKULH5hsCBMTjB1UER/Mc07vRKidMdUuEyAE
qCLniwjqYpIOabEzuP2k03tytyFwWN8XOr3THKRQYafoxi6/j0GV+9yy9uA0LV2v
T3j7mmqCV+uTy+oO45nl3HCrk4owmJHnqi6ms0FholmvP1Neg0QG5lceHEHyVrAu
meEx2HTIFGNk4XK6A0ioddvjG9/f5p3sr7Fo30IWoF0Q3N/EkR2NJj+M/my2Y84c
6TxaVtNMHj3O3N8ok7Xgx9/JOonJvVkuDt1G4s4peXRlcpWP7govjIC7xYW1vL/V
77pGBchZVtaxZnfyrvF0fGAjjJ5pOlVkdr+/Wc6yxr31nkJk+bqjS0jFn2CP5Kul
K6PQDYIQp+TtIsxv28+ZIRUte2Xzn84gCly1T0jiV2VnEJnlpXUKKJGTGREcEcib
6G+nCUF0bD+c4kwtX84km5szDEfZuyzLqgIv/NToWdiP9R8OkDtNmNOmwFNaMQp/
GaQVZxXWZ3KISqJ8kYJxRCPIJbaXjXZEGqOfZ/YVV27G5urWdcI7k3F//3P7el7w
D3iIoo+yrUI9uK9MCo2XlZwUOglRxll38s51VxRZCkjQ2xuQUTbuzZK/6cBgtY53
MT6iR7zOxHdVKewPEVJvzQwXPsDAqAaQzwDbkaWG5XP2+nlhrsDgpdldZYPa+5wa
ifsGhSnmTRHHJSUlrSLiQ2zNL97CYJZIHNrJFiwx0ScBF4WhfoPCHgLHZMO+Aop8
HcXf0lbI8Vw7utSDdf/uE7hkm5zOjA1lhCPvRKVECDWfkgMpQbLk72TYm0I5KrV9
jqSc3wZ5vbbwbAT9vxo/Obx1CAOsiIlSzBZ4JD8CsNfFgzZRAO2pniNrpET/DXnv
dftpo8+8y72a6GQR+fQzEisU1crbmXBZobAKq6ZQLe8M1xSpUkRoSgoT5g122HzG
8kzyYSXAdO4TEegfZOjW3UkRSMret6hxPAb7HvsA7mEvE2dYqVsef/TVPCfNdlmF
pqB7ZEsGcEvnvjpxE+ZE8tkVBvzMRHT7BeRSXGjIM88xKM3ou5OZLn3czwwvB7mw
2jZM5TT/HpdVEzJwa9Te4mzbQqqQaUOa5hPCL/C2zbJvlVWoJSJ+fLBpvQqXkQLj
YqQ+jXmTYOcoMUyhu9Pao5F5SZwrjxcBdeEWCrmor922s/PE77akh2uKdL5jF9LI
I6CVVNnVULJYIeWzaKQOJcEf318I7g+2+bIG7u/C/PRCap+d5E+nR1gZIpmI5lWR
xarhLa28k52aqVX5u+fU12m5nGhApooXVk8RcV6+QS+1qsa75y1UL57z27GJaJiP
WMThStlyDqEEszqW3wc9LtEh/JPsBrOVngQhtYP1zE+SyGRPLEv/XWQMDt71OCey
vegnJom36GLKDsO0OhXPAk92/1eiS/4vCC2bCphasf6FzL31aBuGqRlU4vQu/T4v
RTQI+tHzWw8gqIJIDKvRk6kmXDM1fehfwbE2hWSr4/uV9rXRRutMt/V3jvRlf4J+
1ZYSyyAERgLIJipr1MCsN2488QwocXi66dtdL3yO734TGFBKZ0QibKVCL695xUJq
bKHnYTV4+h3ZUucFJBh2bJggvRTnidmshBAvnsQ3B9lgOtAmGpkvE19aXoX3qnwz
g0M62FH0CAifPHVHqzQPKOwfXHsT1iRIHOpYmx2Dp0J7PxIngNBRBEBdg4vWvwIu
rSIk5/MVblW/VaqSAVGKxmWaazFXDci9GnoZNSg4rXh+cFC6WVMn9Ja08VYJPTnm
PeVvy7icECRW8Ahr4ebbnNTHTofNQeGtf+qEoowdR9ITkxEHyaNUIjq089MypIun
Uly24S1BpeaJfitwQ8tgKjczfb7ncw5d8QchV4W91Ucia2lqyLSFHtNEJtjtkLMy
E3FO0Kiv5a8gQc+jn8TmNTIdLHbbmJBdlDgB8AkUqWftAtG/4BqilNepzY+Xh26J
eAdKYxdENyNCV2PHIrf+rzzcjjRLKyX3rMxH99clme+JRZTz0l9tfMt1Hq5gJrla
EXJLsRytXj+9Fs//j/MkI35HR/odlLFFiGi5aycSTayItdGaMaixLCkrfnUyedd1
Zsq3xOlb79kk4ZpZD2ekxe2Rtig8YBKEdjDJboKZtucLWps8WQe7H8fX1K8C2ng/
fTTDR7ilFunCmFdZQ6z2pE3wCGKq/QE3Hcp819J7eFPNTnSiHZmztp0mQBWgs99e
0GxAyrHTN/EONnp3KU/okBzLHiv2+EbkLnPbwtsVtO9KW3Qp/5+Ioc/8D9Estm3m
L+OgqBh4i65t3UTciwjNlOEjCn9HSAy+Y51hf38+0tM4NR5ANXJ+02BGcAXC06Nh
kaT7MPwgGs3QekcRg8W4WXOqqJlD1un19zUJKgZqa4bylxJ8+Y2ez6gRbMOPQhIb
WF+jmqFKG1MWYIYKIIJ8DTA6KDV8pjiO9QvDbeT2wNI14l7q3JoolnBtGU0qAciy
JYsvZmr/935wX2NpAGU+R+pVasqvZKZ4u5KQO9/cDbAFALmssBLGryF0Bc9+tJP3
Ca+UuLUwrpwTM0KlTihKPb3SwyjPQIo2dDMWgwuMP2WU0x7RP5RhFgQSN3TPhmQ8
cu2SgZNv/WYXDKDY0WQbMcC6t8rhXJ4Xcc9MVMCQuSiyiSU0aBz2HB+YbPxApqEF
EO+mMzKKmYEN9aufY9irPrI8c553BFBBCjFDDdyhWLvBw/lfUz9DNjr1k0z2gMpT
bCELHpczJxBgywr/YAgB4c3kIlsLHw8EUZeUSp3h6Ke/C+r6eTMjeJgmuOzj4qoc
KC6/8ZE9gJuID2OhPXVtDmbmufAFUPixZJ72Gw87YSOlkVUE0nLtw9c6QPa0zH5n
dE1+AaJ4S7Qjm5Xq6KUPTszUqDrfijKkaEfpUsPPlpM6WG3O7rM1tqHuk7Hq9I6L
MuWzhklQRJr8yPelrVFlWo/8xEiwi3VL3afmrWPL8BlQyrUc+KfuRvLj2VulyML2
7pzwYoTM1xHE8tIKn93ykKcKM930ZzlGyGNQFCHrU5qzroZ+kRrmRlvIRYFXmURs
HhWK7jIoHDSh79czVi1tLMiy3VCyfvUyFRdjE0xbxj9nfUodMzK2IoUDWJAn5zPT
a04gVGwL7b2Yi1IIAIQ+vD6D1fywdny6yq2QDXo7xbKPSMQ72bvCGDA7G202s156
HYsjhb8OTePjZyi/8bSUiXvhqHjPWBfEvNMMaeu9EIBpHtXgUb/n566o9Xvv4ZZ+
7vmKERJVMc6Nhp2G1C5mXOYvP7aX6pS1/Ht14XGMH3uIow4XRHwnCG3rwNIzN9d+
o5jb+rk34zJsFD05qsNgL7Mm6NiwUMim2t/kgb7vtXhwApPrXx6kHl+M14AdHXp3
iwDqIEFpwZSv1k53VkxvhouUWZZYB8mK6pKL4xBQrGmzCaFcWFziI8RIa9LNo2dh
FKYGGig/cR9FOdjWoDBQv3EFg8VuXYFWwnQujJVEE/yFmPGb7xlQ02gM5LS3zPXv
rPg6hnvVPDDtPJySNUSxosM4GRfeLkW0Lbs9UvlTx/QLlO9s9ZzomgMZuKv/tR/f
vmJ3q2W7EMpAPRu+iZbz5iEbx1R4JxnME1Q7PbUYFkKbd/0BFhBypgugjnfd0zLE
UKSuSXJUQ8Cie5aCYcaEX9k9T4KFhq1Niz8LG3YN6qE3xh2kBZ9ueoh2ExFxwjZN
`protect END_PROTECTED
