`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Du6Gs5IqgJAt5VNboMyq/HOo6VyfojY9pF9joklQt1qapyqAjJgs/afw57ZTmyk
F6KnHmBRa0v5c9XJWewp+2JJpEo2wa0OYOI9XFoEBCg7QxlVK6V8t2AZD28ukQ7N
/yHmTa+p1cMkb5qmuSljyFoV/jywPf8JrZmaHK4Qz46VfJQBzDkEBdnk/rdmYDWL
fWTwmT8rRAkG/8Z1D6bHkGzhBOpRZcY209b+RMd/dTFX8Rxh89oxrAkGs+4DLn6A
eOJ6lyQFqsWrgmhFJJWdDiKXUX+zq1Jf4iXIWL7M0ajzacBR442W96HRfhPSdwjb
nfrDjylpM28ZKa4a25ctFDuydokD3g5/P+rtREuKQ9O7BiyuT9e6KR35TOZyR89G
nrLjnEMvkRM4UIz7xf5QuMvwF4nU7Nfs+SSQF2K0dDKDWOG9yGX4gU1aNF23DlPr
jahNvjjCzkPA/ZRvenoePltEGrDkjm7H3JIG9As7hndU020z3QPp+LEC4WUL7QSM
Q6C2LApz/Poi/5j7aehb4Sn88FPadxqIiKXGPKYw8HlFr2Ie3bwjF+0v01cBl/Da
rrM9T1ASu6mFDzLE8RBH12wHFUY1JiY2/PJYG1NgN8b+IluhfU3GzaV3NpVv2GVN
/6niX5AwxMYrckshQK7+f8eF8cindrq9/VYK/dn4wdSgycyQDtNblonbFhdqOhjI
VgbgibKOSWaYqXSy2SDajQklntIlEZgqJ+sRKuQ4yAM8MFNVc+eQjpOIByfpngRJ
4FTVsQ5MtNSFcqZwiFWFrgbXUNyJQXnSv98V351tB2SsCwHJfDkmgE04y8RRmm5W
w4VTdzwgFupmNl+eRTmxZR+Zw7ndHJ301cG4Aj5yNmbf5Z/c6gl6QIMg6YL3Lfz7
PVUkHRnIk1xzZlzFd3Zfbxk++rtpKexPrPnWv69AyTHVmgE7Tb6nynPpndTFGWhj
Bi069qQhgmtNviqyzZUjQhVSCv7inUyUdyb8SHqdCi+nJUxOQn1SlB4ncji8zKN8
ucd8QEQqiLLqOWOs9aQqdKFoZ9xuhdeNzd13UC/Z5X/aB/9xDs+APNWiQwTtOS+7
TBzzcVwfFSEwkCNIVGL3ZvIKGKyb1m2PN5cnWxKzkILfVwGz5yJjc5h6tN+L19N1
N6kHRtFclPXmCt9Ax4NbTF2YL2Je/zLunKo6iYGw/Ii8RoPrHOaUZ+Z0WSwdmBQk
bnqAdCtrpxbK3Dyg/69ZZBMTHjmRZdhY7ly8k4Fj/Zvr6jIG8ulSbOGk2D3a0fXW
kR/fnF4cTR3OLr4EvfPK4RMOE5CO37k5BVx+ceQGFAlDluOLQOdK9m9eVOrxfXXl
6u7v85OmwSZgkEOTqmInrMRpdzb33g/vWVILsPgEj6vEKdD0bFZjfb4obJs3rGfp
5WTst/CQipoEKQbub1lWLca2la/LOWm65bzW+IUdIOATOZt4P8QvVBrNErSuMJ4o
QNwNlyJdaQ2N4JHnGQ3kFfshS1lG+d1jVlhr4bu5B7PCDENK/aEcSICpOiIfwpv4
m2iT39dGCNnR+mflcAsq2ektKZK8wI0jp+oF7aCBI4jeh38vEny5lcZbxshKnM3y
uIbGH1rCN0juUfjheFRjtpElAbM8V4TdLxAFqC9ArcPIUFGTrrPop3Yw7woZXYrR
NpSSSzay1k7wvU3GI/MkjSIq7Xs0kFPhHO8M4TDDX8Al19MWrA4ThQmq48SbemgS
19XRBzfp5RaqCudXiH0bEhI4tZPePySI1b0y9GhcDNJZWz+yOAe46/Ds+PiM5fj+
4dkG70q5459JqlXJNBWWfwq0kYhZND+uWB1eImUe8glNKnrCq97Qxk2ZqihEOJ6X
Rqb8/irkHmlcDCyDhnlxb9UZrRQsWS5rpv0jTTgqcd0A9e4uzulHtB58hR1LruKF
6lnyJ36gndUFVCDgzEybyhOJY8nm03l49IDZS4Ht6ia3gIWCrilCcGUqHqLoop6q
qr/ibDkSoKx7oG3i8QHhxN5rykPaWIfxwyCpijDUkhNZ6HJ3mVodWuilst+R98W2
eTLm9V+LYVGq6ZDzGaNFt0RLTroUGG15eAyvHnd2nDpzmw1jRHmM9Z4bP+UqIH+1
f+c1XVwwsm1Q+JmfIBbxqviEgjNHmHtEvALjGyU21e7//aWyOI4IWvVMgU0NDDSU
EuGgmUb6XxitKJJ4cTDRtHl8HvYWhIYRCTL1ee4J7PX1DkG8dLRtL4I0IazUXGUm
ptARuEy8vY1mwPG4eaQxkQ1toea75+wjl1myybwJM7WmugqV4eAodlnHpTa/IsMR
zn0DI225MSNVfAUmixIHsWsT2V8K7bkkAayu3BISZc8Xn/007GekVDPWTl0wBM8g
xxKAwdX6p+Vx+VYjIY4jYAMEzyzMJ6zvfZbYFkEKCBSr4eososcH7H6SZcIrv1ti
7+7eoaPLscF02L9jTTvw8FA8wpRNGpfffoldz/gyCw9niM8mzGzXqxnAwu1wM8DJ
3esZ4kMTqXc6sTsixlyfXTBKCCOphnf45jpEtkuS48m5gf5Wiwz6RkYYe3Zbf9zl
112I4hXK1JftUIE+OcPtIBpf0idzem1PP3ymw5jUE0CVi/zNWq510lNH9W9I4MkA
hdNrU809DwWfnpIz4hDkVnQO4zKYV94Z+Su2AkpNVUFRw7jJVz8/PeVImczs6RJ8
dCNEhZVN5B7f+ZD8jKNbc6+oruob1w8Cv6zJxGkMiUa5bZuNy2GSiRRreqrEHJV/
gC1JbdHcFlXmZA9W/dYU4Ygf/LMp2uC7Bf00d+XOA1qiGoWtl4G+ETjSUKeAq2LU
zae0iFwHLkJ9xHoIH8enpswynFONpIpET412mYg4VXVQ8zKvVlmiU6a0LgIA7/LU
9lICtNYCAN30fKGzS36jWlMmJzRKa26it1Qrf8aw4pu25xHEi6hY0ZJMGwtSv6gI
Ep1fSPjSNDufbpSGpLZfXmqHFOm7JlSsRQxkDXut3vbUB4RXmrzaJTkDPnmZuWnH
rKxJm+yzXVtTwYtx5Xpvp3MAQXWM2ucV5oIUwRmDWGXBHHI7gnV229teLejYRmvW
jk+BNceH8SRKcS06SQyKhBx0eyZ9Kk5JkJ9rVDiEwJtDXRqCW3o3yE8ms2cI4+bL
PAD71/NzpRdfJgUatCmqYmVSb38le3NBvYSmmimBwceNeLI+IK5LsGEWjp0Kox1c
U0PR5xKMQPQKr1NOd5NQBd2+nUpwt7GqngEE5Dm8D1NhVh9OFi1Mi+NSkjCedn01
9AJss7i19Ug/MLYZiog/elZbyvDBRgWHlm1c7r0k9i33dnnmq3SUznKKVPRlAZya
fuxtwwVv0F3AAbvpIwKNwKWrMpxwDc6mJcrc4W3ELdStpyi9TZy+I1tHod7xCKyC
MwYvp3OqhQjzGBkoTkU7vlWhd2/u01yMZjg0rSJiVJ7k7Q6irzVFqklHH/rWDzqR
qKOze+/IB+fswoblAWqYQbLoAKwVEZC2gM6kOqnRJB2D9E3S/TKswLsKBirdGTWv
sHYVdMQoE95rz2d/q14Emp/tu53S31GjpCkR3AAbTE1FnhtUGQ5lMURN+y4nJhqa
1pQ66BmL2N5F6jpyZQ6fbMRNGVtmwNMLyMfoMl6JEk60owg7rCQUvUWXiWaTPU6C
WXcVecJMUA8+BrMIVRohL4uVeS+dAaU7PZ/J9KCBrNCxUXt0lx+wnQ+nHG0RVlyv
tu3pnL4ee/F4bn41nvJgLimNi5gxYqLAYL4zxAW0DhjN4o209cButKDsMILqD5se
AjChjK7N84spAtOdfrkduvdM1kxwXZzJjiRc9x9D/iHVX3b0zX8rlaeWZF5m+P10
gRv1QUPybUk1bJDt9o0pr5dmS4PxKCQmi9cru2TmiktnRPSq8duLtKyOD1qiE83S
plYGwRkWJuWr562Qj749HeyUsFp0yHd2LMEXvNo34hKb2kX5QPAvVe0Rq9p9utTy
QzqVfx2Q2R/Jlu1n9LLWEzFs0ugu1cHuCLGE3DYT1NwIylfhqHCTtc8tG+sHIKvg
uViJfu6B47iyUnkmfTR6mfbvArEdIRX0JrBijMvVrSJZWf3uxedjYTV1nP1wToNv
Ts8T3NmoQgTc61R5PXL5K2FDsFBSQRRPH+WoTeqiLynCGH9dVP8U6BZWhBrqswa3
O6xd08S3XnwsJ4OM4JT2anKWMp5f3och27HLoRJgIs2wadYR664tvWshBLiUzuXj
uSddQtgl1s7MF78ZIqfxclAavPTMY9vHlkQApfi/inPtYINrgtzHHCtxHVTj/0vw
Pa/J2/oEq9D0ep9YeGCXOGX15cr8X/x8y/fNzRtCk9ZQKjCqrIqHiidq6sslG8FQ
nw6f2rTIomnaa+xmvNFhou0CvLOHWaZnEWL8M3++tQc1GQJYOkjFCgz/tiY4QoRH
T6i/EoaLm6MJwxw617l7G9o8g4UQfoIobQb0Qr0TOVuGV/C/Px+jSVP0YAM32XpH
yEw8TZ5h9eVCup94vjWwy3EuaZ8JkWFpqd0NUxWYwit3GdRKQzdnk4mQYldvQAqc
cj9iZkvTeSC4NAtXRp8ChAhBubRZQ4Vhng9UxVwCuTCPSl/xFTNUAw9HDBxwrRUl
ks3D9cLvYrVlV0bfj5eQ5fSG7ichB6DhlpldlOJGiy3lOlaUFObyQF/pBZFvz0iF
8h3Bj4Xu9EQgjOm62aI366TDhxlqY4XIci6PHeGwLmm8S+6AxNU4EOvfsvVXYme2
QS3CSPX3QcLTgS1qQzEijwa8PhLn+dy2cDqaLWmGXO1cGLU/KuaS+Gv2mbHVEXxZ
MoAcjl2q66B4WxYWE89VP60QWM61Cy4O/xVG8iRVWs9f/X1fwA8POsQRWVoKYJne
IPftVhkwuJSwFiXU7Ea+w6PJfJrvHDnazhgi9lm03ZijixEJc2dVvDOLL1OoLTnl
Gf0QHlWGHH0eMrRTMaVGdveL07q9KC4z0mjsXC5NveqhpfXCVZDnulua/ZBAFQGN
Ni5w+lyqiJd0aUDSRbhkIXdrfqyfKl6vY9bQxrgo4pD1qh3NxsWF2qv0Nk9ya16M
HwsEDceM8p0UeE2obDdgfOaxUOcFUvebJKfPB4h/T2hEYpd+1jzoeHDDAkuB1EqZ
CE/xOjpY0k4oq/VQmp3A4ulVBLFg68ah2/3p1AqsKvwbI9n2oOe0yuE0HuQn51vj
6yRVTrrrpQOgGzS2RnPN1Bl+fDQIKZYpeS+RN5vZNg6UKq/qopAbeA4kK8LywhDB
ArEATm8mu9ulHX6OgRqkwIneKtUMz9xozPrXkCyVlYswqFS3wSpxHEPVtEA1g8d5
Et/HPl8QAi34Ve3dkr6jqSW2erEe42uct2zQT66LmNjSX/JjBEzPDTYq9/OVgsBw
90diCLvWYVUIJKnkuOheDjrMAOQPQt3/LPki3Xy4wfV4qwj857ijhhyYy1wfa9kD
UcM7h9eaTm9UQqHNA0pxpsvmUVStRkKv4JVNKKlf/oyZaqao6q9FxDawjWIUqwBM
NnFMj+MmyJ0vhlcUeoDsNt/xnlundUDKifVYxVLBPgwEFrcu38KV1HYGxAOQlk8I
ECUzLImwpqDwfukl/dv0I+IwY4b0Np8zllLCtAADFQfOudNUlfVwDSNYBPu3atf+
kEWucDuh71bHKg1QX/JfF3IHu2qPNBn1eKF179BMq3GeoRVuoQTfEB7CPSOLlkUj
ODNIZE9n/yGUm3yoRE9cLMOn7gjqE5LTRTLRRH98rjA27nDFOpI5oZBFcpQxpqye
QDTnA/+VwcB7CLUXkt4u5a3oyaoEYvywX8ysvUwrv9vlcu9gcnqHzoYn/t5/YZdI
uVwoaVZnE4heiI41WETFMb8CWzJjDmnDyS1VC8cj43NMJl4TmvuB85AJUJJQPRwp
O+feFKpaKEKlW9sBSiZBdqHS4LB4rCOy+LpFMRk5orHqupI01s9oLXhZj7IRsJF6
ciuY6aQpRXIIyXczdEsYL2uf1tJ1a12OGnbVb5ANwBdGn3yulYRvr6C1PQdpiz1P
0OY/7Daj2KbtXM5Muo2jPDTNkFXvDiV2FL8s/b/zI37dQN7C2HwVdZXWJHZWFwvj
zYukkdHMcEEFfCveyiit6AeNVQg0ney4aFH7Gc2k90g6QAxOtmtFzju/xBlRC+yH
SohA0+SYe4RYM+Dq1WJtckZxtHx2odsFbTLWYZ5XbHK4wKdLT4Ar/P9L+5Z9TPoX
+vZWo2YVXUHyOYVWdm7pQfa0y0HwTOYtAp+vsFyiWbO2rjhT1WmHRI2I7sRfsl1n
NCbSLs1uC5Lo9N8gvUvJJau5c5uVpc3rvKjXxh/hXemDtnTQWhzY96zGpKK+VXDp
MSDGe4dY5gPMkKB9VsZdw+VS6DBD/+bU1JeqVkbAnBKuqBPv0k5TUotkYRcKMGYN
lM2xssruZ29GvvqTglq7JAmG2Mz+wb/qT5Te5rkGX4DWmFTuVkmnp2m0juCpEPGB
U+SQI4llY0qd96/b9SFIFl3FpcVYp6dkqb99XdefDlbbwfyk4HA9y8cebCvOTsOg
OGeXNZlVwlRhXlWzkmzdQH4/Ik49WgLAhxZ75RxY/dp6mHxGROMwuzqbDR3kCTwe
kax5QIWiMBZqFCWyPW7Fe7bOHRtNQTqig16FS2vxcJ8fj+hu0otXGrCUq4oqAkSt
F+tLFmV59hsjp36eaGaTevpxqPoafCNZX1A8v/K54UWGYQ0U8vry0GXDbE9pN7Eu
Wwg1uEyuAC2y87jGKIMlvyAct+yjP8Ycu2I60dicP0ltdJVLC5Q9NWzJqjjLNgKf
hzTzZcmHT8IS/nlPegnYCw7yNhDd9/w1ywxUkLWCGjhhCv3nhXALx2U0SfiYnAko
u8vFYWZT4tj28t1tjBt0BBJ8YXPEyzXOdVjX5dAVAuO3N4EIqBe5+8ezqHwRto+a
6Ebjs0Q8TM61WJ1A/DAWuS89F2HU5Hu36ioCS+bGygnYHhr2WP8gsR/qQTH9/w+1
l+5dKXPt4YrHkbtufneVt92qFU0CNAeSx5iwp78Px1UJLcSbLu7wQyZYIlETbo0D
cArOhBmoRxM1m5TpTqHI2TI0UWrkU5YW/GGH2eVQ7quXDezVP3Sh1d1fia+vK7h5
J7vmXuusP4r9QQogc3c3UIwJ1VC8FP0lbnxMMXwXbjuUs5cvBwdg68dlw1k6VDmN
A4oV6b94aIsWoIOaqrccGr2A+jHWST4RbgxhH4qUBrscLW1hzhPKglVv7tBrqW/q
ZhDeAov4Nysox/YkbUzKwf0c+7FS5Uc5cxQW53v1DGp+SbrP61RypJwg+9Fyn0we
E+0MIhmQPL2dEHCqlQO5OjqF+Og2zSqu53++1y8eUfeFTGtWO2pKLeofZRGu2SV/
VC/VEAIjOFtRDLd7EUcsZL4lzO6YtoLclaIbZiUESf011U1YMgFMoyQjWkxq18PX
u+ApH8y4S2+cntBXiyZ50Fr+hZwdWy87gzALKooqQLdiCaayk8+J1VjNBBSbipsj
nm7N+SO7CbKtSiHR3pwUQdDoZnbGwgJQaKqO2XbEsZGsykqO5J4qmsFOkEhtKc5u
WgvZ+mbX6MGt99X6zQ5bqsALLjIC4QZSDtHHpWbMmAuFvV5DaUraJQUgtF2qSTLQ
RFg0WtdqATm1vneec6RjQUCbFsqwV3v39wDB5MOLyY4Ko1ykchE2y6PaZvBSAQ2M
Q2ulf5IKa1MLFjQ26XTKrAI9cNqQnfAxeNCdjoQA/7yzhXpfzyyRGjo/XeqF9Nfw
Mtuavgjxloh0uzCbfFBSjtavpyEHkpoeyi72cLTcFNjKrXaO5/IQEVOUy9w25Qyq
7TUGuPVZyEaCE0tWuEANRFqDHribAEzwJaSXij+1l3/qjXLi8iydkFTdhrK3Cw81
RiNTFt3e7/3qkAskeoFJyrWoee4A47K8lQoBQYz2moCarsXsWxOxgT9sO1YRbCJl
Kr9uE9C2rTCiaLb/vmKagEo2u2GJzEcD5Y4eC1R8esl6I1xl4LlCK3aXl4T8Ba+v
GfS4NijX88Uu9SnuJRr2VTAVrJUhCQvgy/nQhN1RqipWYtvRw56t0ntxqJuQI0AI
STMksS1nwgPHxh2lLCnsLRO1XBin+th3LoAG+B0h7X71cy8JjickT37ZbnrD6S6Z
kg31kxnJvzKzQCfDUyoT98J2RPtWfsrbtZp6NQmoZ3g9jen2Xvd/ISrMVZUYVHfM
nYi/efBFdP/V5SSnvS9hPUZqQpC8MnhHZLViJSKOcSKbgZsUzFxv0SN6psgEnV3q
3+PGAgcSO5IMCAQe3/yjzJ8UFGlpbIRHDxcGX0p7BfzQEYUcm+Hvs+cA5/1GZsCq
b3RGl5quIXlO/2n3l+ofg2rtkciugtVhXzGOfxQilgaWPTNPv4K9yXYDPAzCf+ZY
0igdomJ41Pfg1gD64/uHXfHs4oZZs2NSfRHvG09tsI2EF4cCdKPp5x7CnZaoMCd7
BS7DajLKHuYdgeyPo/Og+/kVJ9KlmDZhcMwidokmUZJtJvsKSKUyBN8DSXGdjvWu
8paWnFbNXYy+h8Rn2t+93KBkcBZqP+s76aGbEG0o9vVopppLzhSkzsVH7uzg8x7+
NdTM2OS4cmcNvGmmPCvUniKG1R5XYCcEZwQl9rQVpllVX76OUqBE91Tjc+uoAMK+
VXGD65jjTqEVUxxBZ25118RLk6L7BbsqFVi46eGh/PMQT1oy+YvSfOBd8VEpEGze
m6iuJtIcWIVX4O9d37vTovjoM758ojYLbAOXALzqHhnLwNwPeeedLvH1a5rGy5Qk
k5l1bruTt8D/Lo6J1x9ZHACo+usHKLjHtiLBz0IhfMrS8WXs5hHYOWyXXz6eUAJJ
8iRcSog/0JUE6LL/aQafvzXlO3Xy8CaWPRHdB2QLFr5vQ0QPLC/W70OvPuS1lPwv
C13bHnLLUVv3BYqPdcyonl5OJAOANZLjiCBi1kOE82Cbl5ZaKtBwBO6QN7CVQBIW
Jz/E8Ue/BTMzevlvZgKtqcf/jDjvl2+W9owTQxEM15nH3rMdRzBUeA9jEczXqZSs
hCOppJ8/1zli1qj7JRZvnRc3K5iFjrEgO1LOo0meXXlbozKQHGEq0Y2oLuJ0+4xj
vDXcTGyu7ExZJZ0n0An/OWoRRmpdUVPPo/oYmrkxNnvsab2gNfKo8hA7duvjNOcn
KMQfT2OFe0CORq9MtZ1QfLTgROJKyemWowChMBOQ+AhGeicGcDDhQrnQZC175OS9
tmjq24Wp6PZXeASpCq/UTSkmmPEva05VpHD4+dh52wDsDFnSBvXGznusXCBxLsG2
yTPW3bznw7ZgHZnFOHLyOKl4dPX/hTacEKq1PQknglQxM6GOSdHv3qrBemwGbflA
24IXhXgbo2/xweq7lIlQu0GkSj/6FBJcztWMxIII8ODjDnNkEZyb/s7ZefcccBij
N1UvcKwJMLPb8M88V+Ll6zMmOTyqIFf86fpuHOn739taN5YzSPV+CTcO5xlteymL
6BOl9qJB54QGbxtBbyh96Ot64CvafEEBaDAPE+gon2IO89VkPNVDskfGxTj77PiD
jBREGh4WkHSgPBBy+NAEH7r55zaYHscSzjK3Ey3+MZEJvD8iOmBahC5eF7IK2iQL
JIkgZ8rcU9++I7jv4Egq9HLubsIYj4npAe8eNXay6FacUWqwvuPrYmSbxmyaBFz0
bYlG/qHjFwSbv864dA2uSjbICclUykKIyuSLlTvLiVq+q5FCN+2vESrqIFABwVgh
ILcy1HcH+fBHI3gUrMNlUR+3clkCiBoGyt9fY2wTCZBFKx871i0XUDIrZ6WlBYEb
lAIU4hlhiHmW5e2RFAM/ypjxx8mRiD+1ewSO54ZeMM0YH+OeRr9WVUHhdPzHEppd
aeXCIlAzOFbuO1fUJoIMaGGw6u0a2z/6Vm6Ow/s77fYSQ7T7OJlQbp/mnhAKn0RB
8qLzttHeJDFxIwe4EJfd6CadPy8mze1qUf6T978e1XM7QnqVdtEJnacae4ZwGqpQ
YkBaSqqmxTjOvZATUv3ZB8V2odAtz1NmGBRaKnb48/pK4WLl6NK8fHVjW4oq/YPS
g+GsnSNsd4fzt6RZZJMz27qfd1Qk7swxLaRCRUxa0EoO094EYHm2nH1N6em9ZJkR
NYkEl68dAtjPZ01ayJY0+jgOet5vVBXpgyaHaGE0k986LRu3JVudzG3vYEfzbUcV
fK7KNNsmIsKM9V4HUXfuRaQJ3RkNGMxMowyC5RrcRqIrv2Me7L70qVcqs56oaqUN
2Ls33qcDdv43Y62JeuiuJlW8B+uLhqiDSRprh35z1kUWV5Vd4GYpS/5W2X4shw7Z
CaMjfgClxMXYYH7yMcAOPPWY3p33MD2w2fD4lifYN/0zbRPN4fvR297kZ+EiiRl6
dh7fQ/t1B7aF7YF41n4H4zAuKAqycn2kq+S/3hzzxgRg48volPB+l2qmDPRztJAe
RM9MP8V/ERrqmsjXuFGdJLs5Qmbbbs0jrtZbUDY66LaXR3SIZk8ABtq1N0yVieyx
DxwlItCz86vfuHMykvECsHIrbecPA07+2lW5RcoqkL9DO/bXiTrrDn+dthRWEpgQ
fXE3o+B5iSFp6MlpN6u38gBfL1DrYQpiHDqb7WUJkCjG9IrapvRO1Emt7h0BYWVF
UMF0++/H0oTEA1rcwoOebClq1jUHuKt0RvRiJKQgjAWB8AgFzL6qg/Bl22lsScsJ
mToSRrsS/rnS7wVA+vn4h2wbHxCJPKi4wLkJspjKJ2f8gHSh7DxKlU6A/ndg4ekX
ElFHH9YfrB3yph5uY6cNTjyjShVKlQAglrx8jZUyZOQca3FuiqX7lj2hfs0gGZtZ
t60wXrJUNvMyUcc7Knh9eO06e72gW1IeM4VuUqYbtaBGhQZVmDIhPgq/EhQyphb5
H8CmpyUTc+tV3ujsZC34VzsDK1jT8oRfvGiehnnKhesjRgIU75wlbZPZEcIAIm5Y
0OPC5OeRnq0uJwrPXE3ToOfDB9o3fcbdcnR52mCt/TjYmxGbQvdP7pYlGvLpgobf
+7HuW65bY6HXfBxdMa/39/u+rQz/NMgPxxrT38rMhu/mrS9X2f6ycSN6FzB8gQNU
MyGd/lkjtYGqHi7Sm9TxZ05rVHq1zTdEfOZqol1HzYafUPJWPF7yETjShuJG5xry
A6P3Ekhcm+PUYzWmf1tG5DAUgzvus04jmnXuJyTn6F05udaj4L7QyyqdsvBRsu9s
oRRk4+SW7DlIXIRWTn7NSJvTR4m4plT9pKGuyE5xDLDxN9KRbG0ohsqO4HBkdPCa
onnitd1gC0ryCy4qdWIQwruinWSVPffrM4nLPvSrEQRA/TFCOrLBSuPd0ZsAAvFP
tgeDlUxFKRpGPBGE9iOWFRnARJHrbu9z8qPa0dOAsJCO2kOr8COp8GlD//PJ3qti
m9tp4xy6UkRzKfUPICIwobTfQ45iOcXfSi2CZXDzeMNbfH3W8o2xZTQ3kI+ktKC/
ywTrf34h1d6rx2xQmAYx+0z9Pq0zCHlskaNT5O6UuGE/eU5MSFlcpOOyjmyHXm59
JK+XC4V10mcyAgZxbq3O+X3k/slI2vBm6zrMKYbAs5QzvLndHt+UiOYi4NnVyRgT
aWQCLiH0eT3PKNKActJ+QW1V+WIEZ3t5MrRTZ79c55UvYn4e5w3j7GDgp2XzRAzP
aF9l6KvwgmhwXVb3HdBM4twlBXpBJE3aZPTcbCvDYQMyFA4hLUIrLMEDnWUPBwUz
lsoVMa4pNzzf1FFDxo3vcflivskqW/4M+gXHNR6MDj7yF9jrACUeVgH7TB2xBXqy
W8JjJVnMqwujlFCnx5H71UDGrDEvM+bT6H5ZIs1ke3ghW8VCs6WWpw4OdIqJXcqy
y63Gj1QWDRldhiCyboAUVTmkc+QRmahimoAcXl97M8FRT0f5K8z5VqBDXJrGFV8t
8/LfnWVZ9yw10ocqKQeZTL0h/wEnPCFMGJpcBkHVMWYj8lP0u7f5BCP/hILwo/HE
8KrNegxnpoLh9JqAcd9C62zRDbvkykOP9MMtaFL3BJhovuZhFXO3UpwQDgDi2Uh8
ft3r1YoLozeFPYVcv88f0fTnz7DGn7BcpddDPZsTUEVXp0om9joo533LkR7BAOqw
Gl4z8skBMw1ufVLfOnFyUWkcUOyBLGWzimYYm4ovGkbstvGLtLXpsPwkth7JlTtC
bJet78p3UxM5Gu08khJKWhtR7GmUE9sVo4PMuLy7ghjaURepaan9YBSNomWMz+FY
MjGbETYKA8HgArrfD97F/26l/LIo+rpsqkZdBxQHmALezHrspn8HK8l4CAFODXUJ
6t7BUN02rL9w8/Tf0X1ZuUAwlTmImyOumudmDsV+r+5XC13LGmsYOG1Wufiv7wlQ
jHnNypki6/ypOP4e9gP+e8DH7vsh7zHqdFNlvlYidlexA5kOLgWBrhc4S9xsUFHw
sOQyFKN8kcwn5S/ntxQGj4/44fac0TjIiDd+JC6g126mZr+uARA5Rgv19nHwz2PW
hqZ/+GbqaRSUfhDBjuSrt2UdRZE+ldz5+dAKwSQr81QDnDIxvb6PtSnFbyyAlM9Q
Jrd0++So7TwqYg+e/YUV3NXgwzyp6Tj+Z2uVGCCdJ9f87RAKIVmTVkw9Lsc76ca6
8Cja8lwyPScxBcJEmOtl/WKXQOMeIYlb9FIPo95BlpXQKMcY1jXUbxAp+nCko42J
scAtkreX09ZAWV5bFML1MNdlCyliXK/X8fppI5vT6T92L+nsJOXRy+ytX9+Dq0dU
E7tqgkbvQF4wa6sitPiGoL7FEJCSJZ0OHsF2mVgVfT49ik75F8q2Gmc544qrlMaA
m2Ifo2C0zabOMuyf6OBqzUsEGKjQBSQt0xBIMxj9Fvq7apGoptO7RN4P1nBzJY6w
w2lnEQYq55WSwDG0dGm5Kd2PQUCpY5gRVGi1495lBV0IntJP35G0DKBVVBqkp9s0
LPmahd7N3paSN549DXiY/8mlJ9I4izgjMf4ltV66Owv5a0M74SA/iD7X8nTDrB7w
yplNd/upJwXCpTogs4Ez3CP0uu/hP1TlK0CyTI+vTWm9WqUmaK73pKgOS03KbHBG
t5KO2Z5WZdSyT5T74LzrJGh4blELcvUmAuRsq0f0A/b6zIzPBb8MQigG7UgDx6Hk
Jlr86Mm4omT08DfDplrQAvhxR2N3P+f/x1edySZExH9/bzURoKPu+JZY+hAlz46z
l3gdD5qBlAGQ1ppMOXd52Nz1HXp7WT+bObbNhXz+GE6diJ2s/Y5ZLE6lsQbEjzGj
rBEA9Pzw7wXGD7PcSUwdGjyNQjRi6N4t6uknAyKj3pFNRN7dmdlS75ue4rp2nZO3
BKGZB0V6rqv5ikjVEPIE1d+4Grr3B26qMGR2k20okPYKkfoqDWq3jbwrfHIrkLuk
T7x7sUzzzOTsmnpOWr/OSuoBhSdvcEzZ+XCnyMCY7ULu3DTq5bWHZqqmWYXcCnpr
8kuGzrRLsayajzcGC33FLPsTLcU8SlhHfPQPkguQPdNcgmxcn/ukDQqxuRZWYjmm
PsfE7xCVB/wsvY5wRMoZ0jrnS8tl5DrcKe6Bh6yR1H72CkkvzbNimJmbPTeahxHM
F2F1XmFtWuSDbsKanZJB4mFp0nSHLdHXqn35+SRLlYTHc8hQJVs8Ox91xD//qmUR
ZSbam+bNziR4/aMkFzvhWzI1zaMD/pxzMjnXNVMigk59/1MXUCRAJmQeXvk1m5eD
SNzgqWZPoiGERe3RbRNZyu0xWtGq27rlKtQozDoSHKj7x8PiPdU9ymhcT//01N8E
ZpzY+Qw62MLSicGQjO6eVqZGlLnm3pOfM/pCDkpHcVWR2Gk45O8pQeCig/y6HlQZ
ProDfDF8GGzuAZ9PIQ0H8cKhXJNnvKvtdQY5syfehId+WtbdGNzrJ//zOLYV1grT
rClawEfFYKbREc8b+sg1EYiCuofT7n2FkcR+GJBsNBnCcc+bQzEQXqHFPjXcCem6
TBC69hVeEQR4Kw9wqibDY9JuYMzR0WtR4Vn5SwmN8ZVlfwa9qZWNC64l8OnOZeke
0G2tFREy3m9LC/3lRbIEyA3zWI5DOPfVz6ZSYBt6Dj1mGicuXcl3CeqtEBu8IEMc
C+DIlYnKCt02ddIDsWwl4FMjNlmPgms/V4NTqCD/f8WObU4hJ8FL6vAp6Qo5Fk2l
7Qzh1bpR9appmMWobR3AqpaFs7XfS/d4nNDXJdH+xMRAj0VgDjdFQiXSsRN6YhVw
gwi/Ad0YHlULksxGxJI4tz67UXetHe3iYF3bl7WO1axGo56DsdzXlwwtVspmIuOp
i2BT2hMcAf2vcz6ONagiy6GlP23ImQd/ZMTZ//MruckOZNuoyc+Gc1AKx0zuPmA3
SN/7Zt9Yoshh9kdcK89/J+/OCoL5msZvv7GKGFW26w83GGIyo7womXeAnruShX1N
H1hNj0jXpzoYkpvmkPTZK852wYA6EUzvWwq+KWNVtmstWzsI6KoL05wDitkwd0CD
U3ziOxzOslchIBrDIXKlKjvfN/avfa0QtEjEs9kaTDaGHPkvMjqw4+X1HYzx3dXT
/lSE6L6vrnNvfDhdo5aMR+AE7ZQeLAvIfgVDK7yE2HqGsLrgD1wMl8AQaUP+NSty
eApaLUH9hFIqfc0h8ZjcosUTIvcjIGH5R5WXIM6hca6yTJtntNmrTqEhPw7eScnP
UqFOY+Xoc32aVhGvxjtdqflhKXxThQWW6+z3JkiJe+0rQPIMisNpSMqqKQc7LwrG
dE4w1ab/Gnyqs1BjX5lMZV/EZdHRKw6YsuuPclVBMKQCawV4ALVQxAjDXeSmhZ0A
Wbn/nRGl18JDlxs+4BTxlgjqtDRuOalVnuwNYXofnhwXSg2Lq5R+/rfXfj6zE1sg
BfmCW66efnBaxgsj2vTd3idKN7N95b5WooaglozPD9HVlWf/5IehwX3Thf6oUVX+
TAptSVHBfH6OJhZwhMptqYR4rZDosvInCw5nTDQilQxhIxW6z8u554ldLJrlsaII
0+vzzOiScVwmc2YWg0Gn8VMrVkZhvwo31N/V2o2ZJjwjT7JEVsnMsJJ9JAeHBZbY
XM/wuvfDGKYBbMB9eB8+D/wqsDZqTpUuaR8tMZbGgA/Pbzq91Kji29fMtBcCQAgz
d3VOyzmyoV/pRdHwtXxzAxmImdR+W7KWMUrHBn88kvZpL6JhVuTDwoV6PTaPjgby
dOQUzkBHlIEdCU/XcQOvo+pZ0qcfn1Hn5F2CeB5lG5G+ZtMj8iTID7qEOphK0gNq
z//S2TcqMyK5ITYnuEaSnQz6/OGic297M4Ov85MEqw4N9N5VeX12eMAGSuS2g5VQ
msyYAfq9mSqMdc8Su1MqrmzkJx0Lm35w5LIX+BNdnnj4qSDxaOrVJsG7ysz3yOw3
uUqYUE86cLc9FhthPXQGpD/Aq5jV76qwkJplW5lMAXw1N6a+J7WXCekk0IZclBEU
xDtn1tN8VgbC3ShjzybTUAeRSwyCXzFxcdqDhPITKJzC/kuUPmvKPQQbRT6cO2e3
sNVjedfo89bd167QNUWiV7dOxumjCyHd/NwoM8VDr1CGCuXGvXzQX/CWWXITmyxt
I/Xj6wC1b/S3iY+6j2PoSDwnNf31PRXhHVUB9Q6eX+fu+T+iAMOdBEO2c+9Hsza9
TwJitBIt6zmvYnKqj/ae1Wkkeia1htxRG2FnR2JO4FuOAGrd5l7g0oE2k8UgaFFR
ZjdyXC5c1id5Q1Ku7ikv/F/MMgIn08yoXrc/95Od4XECIJc9xxaP/akm4dMSFkcV
JzkbeQnLNbTNTaYDSeuyvxUWD+UqCBwrQ21OGOc6v1Sjv6vZ8HC8yHBjjHUkxGNa
peFPLrbbacMEV+/1mwkXQf9M+DNwef7vSoN4xMSRvFxpqLgpFRMP5ZtimbtbTCGl
mIcM0q7ebk/B1wZYmijtUi+FOG7PEv1WoPSLe0Spr66sIqwsby/qO7xbYvnw9pHS
1CX3jMFVdrOmhe3DPkHv+iLW1fnnxkruhFl8jGSS6P3nMvIuIAFMmlE3QBL5786p
eRSOEcwzRf+x9yeVbKUubdRD4rublvbj2LFK2PDzL2KlcmHDWFfqemOchpZ5YitA
sVYJY2wMYzk/gsLyEhGJYtwZEJkKzs/122MJKaN9VyC5dkNfaoIsuhR8XJ5fpZ0I
VQpkHSg5h4XTqAc+bP4i+DoRHNGdeGS2ZW2A+heqk4XTM6EoHYozkEhwiigaIYjQ
3D2NwRgd1Ouo4Hvo5UznLdsBglVNCQMHNUUK9V4eveLykDm7aSoLXXZrXRExOOIy
W3BIrgCM5YAQcrCt83+NLhleE4tGWMjmdz6ixdPQLxCPCFIuZLkZ7b1agQNFpyuP
TOEuclAVaGXAv3/e2F1FoJsrYWwQoUuflwl98pgMBVXtn6ZUGEbiFE2QPulc7yAV
tCvzC4J3SbTEc333wOOOn+KwHftZMvun06y8ryTO9SpMui54RZRBe13bUK1SGkap
c8/v/f8dSS4tsdM8MfwqsCiLCiLL/pEpQ1BpZY4awA6ADcL5s6Oqe5dqnIuEsSwj
vEQNaar5p9o3ITch2o8YYt55Tqlfa1ammnW02pjviulnk0umA7Co2NYxtfEgI3hL
YtCksrdxFjpZqcC9l0HnFhy8rFQ9/kgBABKYl4HmViFJfYVhwD2BVL6v5qO7prUw
x/GlJZViWb60UQv1MPlpT7zR8gMk7rRFdW6SbrJmGwBwh5EY7mG90tnmkmhbY8KZ
+rLElr25OCXVN7LuIukpfqPFCoz4tnVh0G9o8RJiy5ITLqYqi3+FXm10K35wVFtX
RNcjcOmUh3nSMmFfOyZV+ZC7xMODMJYb1+iybAWKVNhJOt7DyTbKi2IMWlYbxOIk
9s1Gd/vzT3XYuWo7rbVaFY1NFauZptSqrRbP42e1tlqAys5Zpqe//18CM2u44Gg5
ddcQMYsVa76PDQkKuUjIdMfvgsWX6nIndTYSmq0qlvLXVpKMse9nhkLUWEuvRDP6
OTI+vTQ5ufvcwCb05QkOo1Ab5aG1xNqP0WXuaya6nXzS4HNqO/gFgCALfO44pWcY
lR8Xo2DZC8STSzA1EDyiNVnT6MTm0EhSAU/rS+8wqLFWOM8LYOmM2/5OrxTPPEaA
iPTpOciuayR9qP3fri6ViPlMyr3BAaI5ST0EEpeVuXywOETNTnsG3Hj8qcFD1Reu
3jbriezngPnwf2y19mS2Rwy/MxRa1eIGMNrFt2IBWGufMLARpJM3aScHoH0zozSP
EdeIEDNPYCHBHxorr4KEU9Tmx8ltqipwgmWE4SchixT80Y4rwzb18+k2L9laZvsB
GQRZqlPhM25ZyEdJf1M2XJbOKmwxefiJESPI2m1eu316dmPwWSbWUA6xwFOx6+Vq
XCge9Mu5PGfik7gHadMdk34sLTZg9IM87BMFJO8acHcH05AkS0wz9+ZHXwYjTRQb
hWRqRKoncPbPKI71JMqzVxLZA60TsdkfWztMxDWuR1bzpuqJiD8EZUfMugdw8Raf
VMjE3XxqFz1RbkkPAH32KBPgvWK2hPVaWkFqQaL+oTPEAEULLX59CPUGnDp++QVr
Ol7P67tg8TQJf1GsOOzKZG6FfbCiHIsjITc0H5dViS0sxA7FhePDzu3nSOncideU
INItVWvKHGVv2mYy/Qhv/ntcVszdPQV3XYmJcgri1hwBed3ua2mXZhqxXX1x+Cl+
IxSkaFJC4oeYiMpdBOl2F+zvgPDY8MA4mn0pE7RSES0/z/DtyWB6hxioIxmcAjN4
CV14lZRd9rFhBJwxB0ZaDhqDaTfvIJrcciXxVup901wg0LH4qYp94t3HRhCRfFHy
yR2Lw6vZ+AV3IkUQ849jiNInlf5l0r3LqhyGXVO0qHILK1uL0qcnUepysUBcQrce
TlNPG30XtVjZj0HskIvlvHA2rGvCCSjMawtutpcduPP1pnwyZCso27ATtIZv/3mq
9QUd9kJ95fJzBK5t+fp3/h8/jriW61RKOXo9cVSLWGYJmweTAiFmtNImQ1rJNF+L
ADRU/AVKh7SoaNLxuQ2Tmza3unzEKdOTYvTUiggpSVbonOLLhynOu1fy3IB0dq/f
+5GSIy44EoWLorrKDQqFgvKas0L87f4gSKfKhdpuupug6tJDlTly4Ud26tmygMXX
7sR4U6UyqRpHoD/yoZYITUYKOo9TCIXtum+77b7qk2cNzW8x51Od95WIDR4g7aeE
aoYK1f1VfcITWdMFh4l6EJMECy1vQMtjhChE5flrQuZeKokNsXnaPnKpQ3t9m4LM
YUkOOCs6NUbnJTQ5qVcT0h9UyK1vJee1IN/fecK55g6WUZs/iZ/8BP4LTBZsU003
IS/rc6pBv9SG2NxsEd+0eDkh4egQfSVLiQjiBFDxPyS2RCyUbcWQFtXJLGZWnN6q
5W2GK03etjn95jAAYZnNVXS4DcrCps3eIU0NBRHxz/yLe/EVhhCppiOaYBd1HyYA
TPKIb1D6jwaxo4KBT7gab9frAnnsqdq9BtGiOxrUWSf/RMyMeVgZkCa8oMcv8NsP
Ss2k3Z0QWi3EBJJ7Tjwlp5tBV1rIA5SSIcUeVsWywKihvq7WVhvyW7SF7FjFgpOS
BNWZmqpZTEoRZtIvjk2XeSmPQPpn7rV7VFcbLkkKvQk3dfih/xYRt3a9pbMMfAyQ
bER4VcrRQQDL0aPcnqW3T/ojcRF4wIVFal2VV/hH8Xb8f7CcyZj7HBfkIOBY6T50
iFIT5IkxpZfz3WU/DdMTIWVt/0L3yn9C1KPCB8bnXesduvzZ6NoLtuoqHLatcMyN
s0GWzvGZGyfY6/MC6T9ROOBChzkbSUsBOlozXNVYpSggOMtslAD39UJar4haz4wN
v/mlCf67y4csVXCqIQZyLkSjsPRhmCDaLd/RoDrid2eiqQXPyK8zX7fcGuxyg/b0
L9nHkdU1Jf7eJlrxbBrrLFXhMI1L8sWtJ/A7avFu0AmIX1Hu/RQYDZtEp9HMxPbB
E1188bwRVRxetYB3vs27qimjbw4wIFnxQOIh9t3qRrkwClsYgnhFC67J0YT5CuQP
P6ymTFEmFOdY3WCvAj2p8nQ2l0h5TTFLFT/5mnDX4InR4w6Lrs1c1IVUvdGYVTHL
s7Wbod851G/N5mSBbJND06Hw3FxQ/CS5eUFR6hvfGuH8w2IqXJ+QRp59skMwK8q9
QYHwf7Zw1OgHl4Qm9t2XNHpshiKPxogpxTZP7gWfx95twsCBxf79fE/x35bi9IKM
p7+LMOf0Nm1T47KUmMdbib0Xe3wVST5AM2jpq/bAbgtYZkLOJ4rorREKvQWEJJBX
RT11CrzdZTQtNLOLYk4HvZhhhqeSzlUNWl8F2FX80//NhXVLDxgSscIUBq3yfbOM
SkRR8OeGE1coRcgJ0VLQ29zxiPebovITuXvrB8oklovVX59vIX/6nRLQ1ENwTdw0
PrPMSoJt4IZRuxRD4coblUZK6AIQ2T6jYaxhox1kCVuMEwWWEroK4W2ceanKrj1A
zdzs/bljN1mAQYTTv2492dOtnTb+P2qFf1QGsYLAdxakVb2KyVRUstiXK8MDdjAp
t7ng4HLBfvTOXUXZ1NIBfRsdJr/7ccVrJrmZDE1jMBOHRaAA/NKW5cJaaVJ6oSyy
jfik3o+ZvmaUHsvkXvOwQ+tVDKn1KChxBGGkJBQDpkkUImY4vN9bbkVrDlQaFVsw
/PdqRz116qgRXFlAS1dGbZ7icWLS7A/+9wDxzMMMCWgeXnggcyCmWX7mQyQIkfR+
tCpqqQ1oN/08jgX34LfekCI8hZPUwiWSx528k0hQ9fQx5AqZyOzV8NHu711SXQC4
CDZOFuqy+P6pkyF6/eRBulBZ6XbpuShTkAnjvialBPRRiWamdTf9IzMlZ0rPPb0c
K/S1VUFWrwf85MUCWsGsbHfFg3Hu5l7e8JYrc+hZ5oAbjiJPkX8KfoiJfboeb8UE
`protect END_PROTECTED
