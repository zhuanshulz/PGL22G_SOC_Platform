`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2wqxnsV3Q3DTOZPZjjq16HUFOXgagOC2lcBw03qZ32r8IAL9fS/r7eF0taycR6p
niuklTHF5G+ZQ4z8T/66TI+z8v/Rx33neADXPpg2rlA1AekoZqfFThqYtC8yNYH2
DtqGXToQCz2ZUpFdDx7A71qKfdAI0mDwg0KbK6y57Wmm7bCp2tDnzMrBBHWdX2op
aZg6AWrZ9GBLGyzWiELlwvnhhjtbBFkclucQqdiEJOUHnbmCIZfclwa/DFPi2f9V
w52gVW8L7sPI3sBDJnQIAbsoWBZQf2ndyhdW1MABgOP2MlA+yMFMP5hcmWI3Z11U
kSK6Mqu99q5PdHcQ+7kAl+7ZgUwjNPnsP/YuzTmp2yzAxyWSM+nOoFrEJa8cxK10
P88sC9GOF2GL8Eg9VKYlZJ03+dd3lHEAdXF05YyfT8v8camivaPSmiMwE8lagCXV
VNwz0c6RoMecQxc5oTK4bQh8FVsFXPpN0r+d44tSAVvoEa+s/u4XJ0n4hWY4J26H
+veFXkLE3Tr5owPuREUUgH1DpBzdnGbRdyQC/bcV8S5Tp48EWAxziQ5vhjaUjFXr
aOR9tGGUUpAHprVYv+xqkqIpLek7KyUsQHboBmAM85nHBNQdakH+jRP84eTAqujV
guWBqLyhridyXY6bkIHaHlVoZWNQHbEBjcQFwzH1NrfpXo+dtMWougT7kd+zq7ai
QxkFDeETbbvSm18ktmAa7WdKWBv6GgOMdcrKXuAcY8Y=
`protect END_PROTECTED
