`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vtpn99S+Tq4W/fRGLz1hOTfIVcFHDwyIysnF5Vn9A9eooPmEt1B/6KdqyQYsL7Ly
rW5jcHbYtS/UDNOpl5rLj5PDhwbNhwEWIXgK4/EZXmrxUhaxUhRKVkZlZnxsK1aC
1iEO3b5vzAyc3JPUcsfAtOAlvAQbJBNPpFHInIUIeodZ3pNJzYkYN0Gtbz26rWaS
2D5sZytoV8WaBE7UlMEWlWkKsLCXgchHxng7QJV39puPM7iJ7sAKyQJU3U6nu56k
DJVaYVj0bK+nOPPorLrpIfO/CoNIFVtzGGrvIJ8xmhXYnVBJiumDSae9sv07RaKL
1XSGblZ4bOgUQhwS7Do8w/K1nClt4r/p0t0xbqEbBAy/WeBJvsr2l6LbxmQcoOpk
CblO9tZltTwC84mXTYK7cDuCvXPdRe6+gKr6gAZPXXRBKYMLYeeO+1puy9vOFri2
CLX7D2h8VfUfIBUFn7DbB0G62YZPy4IEFQOCWliadF9XdWw9cbsIncGaKfNoGzOA
0opF5lGV3bHWCHLKw04TT4a9W52bldFZsshE5vM1tEWAzxnz2kv3Mu37JrzlO7nb
kDTCUtRAFyRl7OeILt8qRwsgPqvma2ZhO2KgrS6ADPRmEE28EfvKSy+9a1jdWYRI
+SMH/tUeJP2I0jQpqmkdJOBOwA7TzsodSmmTWKse766GDPjSUyyf+yb1YupHPncB
q5D7H0eYICKaabBDdwZWbUMdh6qBK5A8UZ9KJAIvYZ9k3bOOZvP0hHUVJCVUjpue
xkfvfI7EnsaoSUR5Cba9SB0HfusxlwWBDKnwH5VPikfwAQbNpcK9Hptdzkm+W3Bd
`protect END_PROTECTED
