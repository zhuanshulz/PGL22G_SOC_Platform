`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jl8OZMmNRrqnmnGURlNY6Wa+cOBxibbvo3indXGYJ7i/CV00hedckwYNMh1sVYX+
d495+uAxW1KR+F8Wh4KTPTf38A0dhd1dQ8pbT2CStCSRFpA2OybrUGcIaICJhyoE
3NRXHr6vS045CFmSn7gIfxZx9lIHo9SOPRfhhQo61yRzrputONF54uBupLgHBg5e
5Yw8GfZHcxnFRQWdUDh99oS7FPxm/9cYjwfjHFYmwkNH1b7QBuvTgQApqj5J4nuI
8hhBk+6eAXnBwOr6WhaMafVwFdZoNn8MXrfq0KruoaWqhjvL645uC2GXxtFdiSy5
uYa2jjoTW5rJVqXFs1mr1A7xlhVUSSPedCBtviegySqXie/Nsf01mfdZFV3NR2AE
dfAmQ3d6s3t799pFNwcUpGjrlDZbpxRfmb6YlwKoc+jhfoX3WzPQC9eRi0UKqc44
OwdknD75wlPOF4WLxtaVvvpP9Ij9pjaPxnGjZmx7WBEEbcxh/OEzAluajB2YVPsH
vY/gLse1Y4DWQEjM1zPZsrLvMWHHgPS9eSTEdC2xYuBJtqUG/BReqExzbFsRd+Oo
4C8m3hn6QTat/mi7elucGAMkq7hVH6xkH5e41uj75M5fdwsNIW/ZZqgxQzB5dNA0
MDusQCoVM8cLsQE1EnKoQb6FJnekCBZFzPY8bEnX9yFcl3PnupzGt6KZx8/euHOk
RpAk5dPVP0rzpqve+bDjMYXwcAFdC18TRm0u6qZw9aT5Ilz9dbHvHMPFYPASLFjd
8vuU26Zrk6BHU/djWKtN45CYFkCH5P9zNhTY+QXHb78=
`protect END_PROTECTED
