`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WATeVmf0Lq8oVIA5QL9QuwrP82oI94EN5DyRhdIjYveITNTKGYqMHRbusNN/PUKr
myj2FQ0BBdY6lrqztZrr9SRc0eYenxK20PFBHrKVtRm+TbjHEXrx5L8tjaYPECCK
tIW0et3xbr++UPj/Tnr5fliAd6e642l00kCjIRFtMUaDcdShXVPzKnb51d/vHWLt
kHHu7MKdyOIuTGGiGRW4lCkQEzi4ZZlcHfNQj7ikc2VGSl8AD9bSn1i340AToL9U
M82QO1SRTm9+s1NRkzoqSxomcmczUqp5nMXu52H2340ohPHidsc4rpEXwUIpALnX
cwydKP4f5U/5lKQhoGpkBB+e0KtKf4WWCQt+Ws4JatSynuIFHJsUU2ctq7EhMeua
CehvM6s7Fx/FB20t5k8yJw6luZ5ri7IFHoj57Hflhcd4HwVgPhHUBbclHdO1VCBY
hoZaslZrwok6eSYhWaUWHayjZ9u13i7AzGTHPYQ1VR0=
`protect END_PROTECTED
