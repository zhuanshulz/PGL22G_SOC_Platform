`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGxJK85Z/8IiXwW1VW7XD1wQneZ2v0B1dwrGsyGSshBOaKLbXe8wyhbgQmgoEVGk
SPr5Q13t6JRxL43obohjddeXrgUC5UxjSyieoEj/hzN1llFT5h9LXpyUVoHxjIeC
rMK84iXWLy6kU0SfMD7pxWJoOi79iytWxq2A1OyIvA1L9zSM67FocqtyrXvEQzvh
ZmCxynTKzy0+1DYQM+Z5uNVPU3Eap0/bBQC36PivRJ1m5sLFoUUDBuIZiUGJoVxE
I9XObSMfNMUeF6bMXqI2/W+GLEnMWgJZCtRkVaV+iGBTLnteFiCB0RuOUwj1Hsry
4golJKq1HjMFP/Y4crwKS7rkGDnAWfYa0vuEzxp0696lnP4jODAxZ6+tBctW2Bux
HYb3YxnLAZlke+6gjtfFWi7IRYWAaateBSY1kYwWy/JZOyjiTPrKSqXipwMb+5gl
j9Ma7D+EIMuUcWaF6pRNtnlhB7PzO2FCmYIuFBq23Ml7OIHxxugvgOJvGqagkSqw
GLoX5lbGej/ytx/uNnwtY88P/fFT2AN9bm2rx+O/tW7co3ZY5kbR7mUGPSCTwMOJ
cUxQzMQ9dAKd7isamumdOipzQzb9gL4W9lC421yzhQqnAFqCpDqrst9PJMtBaMuk
TV9TP/aQjaIbvJM1x2vjUldQ6hRwiVyNbYEed9RjvtuyzkVzck2JL35ZTDc0DO21
EUfETsdx8AbBH/WlSk5hoxwR7DEcrHGNkxPwwX/1Q7fgYHRTsIHYoXnK+AOFU9y5
C0+Y9PFv1lr/5CpAb+m4vY3g1HdmPECPjSNNClOpwFP932aJ2/lQqPPKEFB0xGR3
bMBwHOec9YTLd8FWXGNHb5S120eMe+DJlv9a1lb2rrU=
`protect END_PROTECTED
