`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXAEHzHrPR+DatRG0EyQ3UoSmW8JpofpqTZsJPx8AYHprXOVKQWvhLThKyJuBBen
tscXkrHrTOiHTpvxLH25Gjb0+C8CpjyTd6e9qr8ICl4kB7HDxqA0pDEQq7M2PdCK
H6BzL+DbF8cl1EQogwxExYywRiyq3CK9h8y0J1VnRrGPqvpY5qr3tktjC3QAaSdR
R7CzolRo57BUVka4v9XHp8j6HKRHDSj96YjAkiEuTb41S03NAfh/Y5O3dCumsOnQ
LqmSiwrPkpClG8LyoBtcZMjfI4NaiQpEHJvWaLCcnqqsPAMCkIpCoMvS53KsE9w/
hzan0EzM2I5IeXwDVU0p41D+rMZXkByPB+DkI5TI7ce6CMYk5jNdOkydz4w3IKu/
WCVUYDkyBS9JHnL4UaKXZdyNK2Y+SZCkhLFJwmEPDH5vzJzYj2zEviaOz0GFI7eD
5pUBF8js3Uoa0jY4V8akRXJ3YfXXO+z+QvhxROmRh8K6F1i7nRerwNgumsAqtxO/
lfsjuo+vs7cEnF5r1umDpLaQXWbClo9hIsjiZX+lYn61Vty3BiZzGrZkfaq/PK1V
ft73ene96J/2VdCKL/sQNKO5ZJAqrpv2Bbj+Afh1kBasfFTVbyauNsTr9drxYObF
ZNNvbvs3cJ4ftU3b3/JxtMI0DNEalM0aQ/47tJ/NdNci1aWvjAMmHRCCbUY4n65N
9KE9Z+0V6VU/nYQFLVeoh1/JbGTsZK+fDFGiAGVcP8otVcy+U6PR/Ny+LB/BxnP5
686vePcESiakygA6ezcGR4h6FP5wOxmHFQ+6wS+hgLbNrTM2qcSkCliT7ywwBb+s
i1prOwQmTHyyjyYJYBlSj2Jzo+QTfJ90EhCEM1RGuy9L1hA5Ka1MQaMwmF2y92b9
EwgMQLz2c/Jbv1p059DSkPjLrGrp3wzEMN0rOAmICNYKOxH6SboD35n3T3MxJXgm
1qbYv+LnXMVg1HUXA3obz6240WVRU2CatlgI3HCBCV/uXuq7ERtxVHchENR3OR6M
/jqPMcWLUQ6rCU0JxDhmxh8niitUn0kzYMLKjkrp8kwql7VnZe3Ku79uYwkB3WU9
lagRneYW8fq7DHzWeQfD2YueQ08TjUA8uUMKWcCyB/ZzZf0AwLOhiiIiinWNvG8C
lpPQBv99jGUwNbyUsHVJE9cgX2nTCLCuWXQa1K7rIabLu1vwzU7TvKBGLqFhndbk
uwJMq9+pyffssFUqJM4dLlB3z06p94xxdCptCBSUWXZQAtwKaGRutzfa6FLv5FXC
BgEnMhw5YV1NdqGlCQhbK+Qmci05OGhurwJxBUrti75+87XH6Qx91xEPKWNmB9Kx
7EFD5wBHEGZ+Rb4mX0xKZ/LO552IMI0fE7Joh7jJcTUTw89B4cXJwme4iQpptGQi
sOb+ZrX8VwRx5Gl8sgD+OarR+TvdIH+SK9kEqXyHuaAYC5zQvr6o5iltV3OZLPiA
ndCJ/BcFg3HgBc8SNFx6V4/BYJYEfzUiZJEkDbL/WjE9x3vA8+eqyEVMHGcCne3W
xpd9QzzRPz59bbI0UBldnChh2Iz/1smmuLm4zN0k7APwOBVa0F/b02CiUWaoJALC
sMgM4EnzfUp/TE6X8OpkPGBXJlesgSc9K4gseO24t7FU0+xHmBIUVCNy9PiS/soz
c/3PMuDXHlmAmgGT61VdW250I6bSu/LWYYa9USHD3OwKAZFL5oiDOUKoRufndZx6
fUBDewhR5FK2zkHnPXwGdOj8DhH0stL8oSUoTe14xtKZRnNTNfOTlAcVl+9A1cqD
SW9c4Ga1x4cVKA5heL5ktWYShaf5kc5IubQt/p0vGx2+r4zRucTVQoRIiRaBpl1G
hiVDI8swKeaW+rYKlGvYXBOUShU9Mx8f3+rvlUoUm7XP9cl9jTXxnvzdS0WRJS1G
k/236jmfavOuFqL1k3vPoH1GFYAQ1nGEZQNfAv3Bwv9MQKuujn0kq2+bHdDS9aML
yu9eehc7p+xZAp+KlIS5aAxAnBH5yrtuCn2V+LeNhtsw0026xK6fpjbcgwZ3OmMB
`protect END_PROTECTED
