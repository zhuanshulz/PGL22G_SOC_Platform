`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yww740/x9u8J5fPJdJB7b44QT0X5ZJ4SLUUPFkmZn6OeQGDKFzrbVP5BHr0HsQqq
bAzhtoZxlGR15L1YmYAg21O0dBqR5ZPC3xjr99UWiGgcd/Txg2DolIgrXAEl3HjJ
E+274aMO+T2AvfLHIxl1FUXJVwGQo1Qb/lvyQ03EX45sLQZFea/xjZJP3wN4u1Un
vqNK+7W7xKLoeOnl6u/Zd6xVdUVbtIeRsdv3ah4Uof+cMohwqudI0sRWPoYDMBbK
T0Ev0GdktKjHK0Coux9LCLUuNkAF/1VHbJDRRitXND1hOPGSAZLQe+/PuBKMPSYu
u0UlnjaKY3ZIGou7WnR98nckFCs60OCFmaX4/KmGr5F7vRvharHmUsdIb7kbfPIM
V+2ijzCtZfOmt0UaVhKIfvsgYFlD7+LIFqVkEAva8o/sVs3lkWRj6c5LGVakN9/X
0AuHWPOFzNl+21HxhjqDTLX+1tetSOewB/VK1pDzE/lSl6bZC9TasdW8ZZ/EsxjM
0BZHfIxU2egQfmWVLPM1WzIJ8Y8e9VPZOPG9dBbCzow9BKSbS1qxUlIUJ6+pRVDZ
4lnHTTOIGDoYnEFwYpcIR+Zht003cmIynLishttVy1UcE4dGyRWQ2odf5kk0vQgT
yIegf3bBOis6AFcmEABVdgJd2Sq8zB/8hdzRGLZDiciGXEwMm/g5nhvagpbIbHPe
GT0O1zWZeZ3jgFZa1w4i5YWy8gu0aVBYE8s0FCwAOHtH/UN4P5wqOCTJAs8nOtNz
pvX8/ZZxnjnOgP8K/Qum5CG+nJAV39AEtmQwLHIexa57XuaYiRYfXS1J85IPD8Gj
SvyvxnvF/dXngrdsJ4t/iCSQ3ltx53z1ZdpzkdxuWRvmZ5eYk04KM8Sr/Mh/rTsQ
AMsojw+5mUbVubPqRmfFc0l7WjQVf+oFHjLjVsouijP3genOKmQ8/bfvQHBO494j
mPU1TQSuoJS3ENfJJZmmcenWjtUNlgF2a3kVxWcEnugHU1NykNDzlJm0u3aZUWfI
4/HwoCTbx2cfqZ5GktXHn1O5//s1zlTJeuu/yZig+lKZVm0JM2wqKsBVzoppgO5m
9Xwz7iW9Dq2+SwZKFZkIra9BHvHdttfzwPHtqNEDRfcTR8+EdYI5/gTVt3m6Zxfa
z0jhcQPO5oH0V8Xbonqb41TE0Z40zlWJNc+z/grwJotWKA60CH1QncIvM0win0ze
TYjou+xi1vTX7hnayxy1TEzsqs/HLLRbWT4l1f5BiEXG1q1mRR8ThSY1f6KO0u4A
788pVJPjZOJyYPVMKYfSakUjTL3CDnwNSI+t4bQiM2s9gIkwy2EjfVrZ/9y0s/NV
VPje2MB4FIIm37BG3K2StfoDdHMPB2rii2UXeQT9ARkmjqjwB9Mz0XLoZm8gc0wr
RswHPJaqGSmzmEGDQO7Di8cGqmO5bfeXoOeoG5KY71/a0iDPHlFcOFNM/QjUya4B
DA9K8gL8s17HW1Va6V2EON6waRzewP5jcWxnE0+MeO7m3WZVXl+sC1LS3DVkdEq0
dBG8cz/7zdHT+5IW+bpF7XeUvvGYLxDa1i1+SMyC+LQ7RYPbt5afVBsNDr9Ep7bw
5cBWJOy1Iq5RBHZICIbzUoFwo5LrbqA0bmkfWkFKgyjD7cwnzxzybmZS+TPDxbsE
dVfyeeeCek7rv3sI3OorscqDm6sm4y4C++W/AIuXGgolId88Ggc7Y75rIHjz/EFh
lLvhUl9TN7r1/tr6Q6Xobdn3z1lB+tJSZY7M/RXGrrVGHcI+S5xEUvfo2me/in8F
Z9rIfwjLXpqlUb7jwRI+EieHS162A+YhIQhcKLQ9KhZzs12uSNVUos9bUjyqYTNJ
dbYxbTx2TryLcWFg3WDBSSb6gmsOgHvLTidqJL4uMaoZK3XWRtD8U4GGDw6FMUMn
40fb4M8nUrOEIY+dGS/A+Hre1IjP19tLl8msluspHIObjW/6698C4q/fGUqDOc4c
Tlp4z0yFrbcJ4QwDIMYxOWd7MsbZvaArlnhdgLfqy3tpxRWHaCHi1l4Jj8KrhIEm
TxeNnxz7lBANyujPyJTncsoOcFYi7oJXYUthf+Wc9U/KmXvbNTajl9UjpfaA0PEL
50kuuRdYr9qsd4jpgOfsUntZy/eo/FeKhZ7rxR7VbI/z+sp+JINjLFKdIO6cKDzW
RMrdCkR2mBPzpzxHQ0HmUNBkl0DeotGz1A2TvFlUvBmxQVWdjiIgQ43n9TfBWq7A
MO5d8sApPOORXN0twxWrjE85NClhx5Ag8WwiADuA1ko9SuCIZt0DsMW/Ee+TBKRA
L2m/uqZpadozCWsCFCWE02ilGzb1zG6sWjzltAU5mQ6lWP+SipRp5YEeYiV6bbxl
TjIMU1Xd7bFFFwpllL5o7ETPBM1aw6i/h9PQEDwEZybS6QqMT3NpboU4cGEpDezJ
ldmnF25v2Gg8e7ErPryI+W6EJnM+WpWRHMwYsT7QYAAnLmapcsZphCtosUjmuOJh
QpsgztEJoncrkf/XrXBvsfIAfq4Ah0ivDqXYzGhKM229fOfqGHjT54lG+kbl52NJ
IBWKG5u25oUXTI45jltVQQIAEMfw9bqa0vKSwCCOlwq9lXXsRRKVZudKwNd9Cmgf
lidS9YlGoQN4Ybnbi5X0N/2kWaq6qyuSa5K1RJiKyCsfMEpOlWczWjjO3lWITzyT
G5NGrbPb7GYN/jD/ayV50AIx55bEbPRa1PAlAV78zrCDWPw6V6UjPzblgOCPKt0G
dQAOSzPGYkSAkQKH6andf2OmPjYrtfSoD6IX4LF9RhwecCdwkLafO6zP1sLjMPQU
7tXol8Dp4v7eCScZW/WTWHufqiTjHfdPp6dff2/vjjYEY1hGrEJHqIenZPzyUAnQ
2TnEwTnFkzJ61i+aq6yg1ptgMkGiTFLdadFPlpm2WuGTJq6tmIzC4A/9ztnSXamt
VHz1xIOABlRkjJlDlJnjVWE53SMWy9zWx0aTx2riwjiMZIg8dEQ6s5i0SqBk+/Zq
jRb/YadROqxdOAefQNFzvjlJbh75MxBYQYi/94l/bB644KhiSxMmyTfaxGwnXv3j
GItoNkZULhEAm42v0l+LZcPh4g4tj1Oy6oEwvUaxzW/lNCbHjZxvX2MvBszQtVRF
AIBZBIpmbJ/hdylzhcqBIIIrWsD/gCfxpwzhxCazqPPMoonCyZPVp+lI68lfmTcN
2rfBHpqsmabRWH5pBr2YNAYg/hTa33yOPKU7czGJInShx33mBlAVffMhu7WwJzPT
VVZ/tDsWCb1CM1MHGjZXS7/eChgJt3WvQoaqoet9Mcd4+lLUkWvhMDN39SERvmwb
+9jnvjxGcubKTqRm9qvby0RJn8OJbgluy0km77J8viIt42QAY/P+JbSgGPIkY/2A
gE9YfraygfR7VvO0Fnugak7UAh2ELvX/1gLDpLjjR0XP7kDRFvQKmnqFLlP3+S52
2BDkZtzBWkuKqNAh+WR8lmh4sdYEmadoW9LgOWEjo3zHQDR5wedizWNtPkKXbR4s
ZVWEIkVkoQWLRdNraYR0Nypllw/gPKRsTq+fxa/8a9f+nTijc6Y0CnqL4wlKAc9d
ioJEWVWqbTKPvgOpQ79a74BdE+Dj+EEUe37S/UyfvYPN8jNDH4FrrXwWjGm+QMC6
9OG0oB60QJm3yVtyQu38MhoMI6He2AhMHNArUNQdwYRfHCpyVQhi9CwO/l0mKw9i
vF927/HXs4qGEn6l9tx43a1BjUuLdAY4HmsM4cBZ/3kLpJ+Hemu5go1yNuZC+v7B
Z7oFWvcEFFcNBz6O2naCgcClrDVtgWTiFVWt+SWGFU75fEo4ZcFH/d1Fl7TVxO59
nSiFA+16riTpWAL29rKSN+dVVgJBNA83+tPZygEc6AZHOmsbkp6YSoa2BQ67ChjZ
CAI+BRXtk6sljnOSNPT0GEVjLLuvX+9TZL4QcFtPWWQvyjqAvm11JmR/VSrEb0K9
IeBdlG0BLannPU+Mt8gIOmStg2kDdcado4GUu29sASAB/O/pva0PCdlmCr8UJiZ6
QhKJUCv/j6MxKMTrE0VERQPSuWr8iipbQ9XkLcuJmCGo/UekL3MtNudaO8jms75u
LxfecepDbS/7reWTdZrLgsblFU5GNY4CQM7nk9oXH9b48s9TM+iftgQUP4AKC5T4
hLJHNcZ3Dx6X3Bj58RIjuDXpxr+0lfEAyxwcqGbHc68TwlIPckn4XaYrZb1RPFJ2
OJ63uqpXF7/XmLFhauCZVmgE0w2iiux5MBKNjpT3FdjgAJBzuWoxdaxIOWXchKBD
tENPyWww6a8e9cBTmbnGSbc8R1VnoREuHMq7enas9jJzqkt5aAZhkYF1eKIZ8j/b
40ZBRVr4o7vi5QiOiDMRBvyWw/X0B73qZrWUkcoVbXNNlxbjw/v/XF3XXzhGER96
9oR4aP5G0uHngCGVRVI4wwc4NsL88px4aIS3AkBH/fVa9tdRGxTtDeshdwhJ3qw4
V098IXX6aLjo5+zy20sWh503SJ34RKruo5/rBW95O7+uTfgTESiBJUfBksmEQiiO
csslEzeGjS+qdg8gTo+aHxyZBWhIvEinv/dIyR7yhZ3Q0SJoLvwUhxGiPL6qLVdK
P4CVQ0fwhVjOsAt305+QB+uC1WPOwiStWIsYZxSJp4IoAf4D5anHFrl+EG9cKQUg
XDo9Sesq/pDoBBV2fvISyTGIDzhrF8UZWnovpkNi82tSs2bJ8e+c8Sd7Ci4MJ05w
9pHlnOhl+PRoURq58HUKDEUdqzfLMUK+SSlyhOotf+DSZOaeUPnXeJlqZDakls2S
1ZI0DkudCy4zOSNO9sk+5YwioIowvLCpQgX6818k7TFHf6Ps2MGmyyGcDZCIYbt2
9vAnL8eOo5DO8h7OdR7t62cL+O1yF0cLPQqSMcBOfMnLDaRmOPce9aFkQq/aMIR1
QIKGAtPrDBDpdaSN5EsC7oN3SSJ6LK8cWueSmDiNJk6/647LtJO9RT/Jbh2kJACe
7KQfJ5/Cq93LdFoL57JLi8ZGB6WbMG1HS7Ywd3rt008CxQaQWXFvZQpacZTSw++k
E1l2iX/wI1ATFCiO7wraS0ykYvKmgPs05yATlEYmWlvFt2hu8f8ccvG9lTLHEw0V
j6vXrXG4usDfoBwOvuj1G8xL8etf84BdNtS477Az4TEU4uYAw4hx9tm0Hpo6TtGB
4w8pWsLt4kKSLIiVE/9s4WCoXX1jOY34NuuXNPd7h7fRy0+iYhDCRjthuNIk5NOR
yXyyfhXonAqx9peLedCCHtigYJmvGqJqCf+c9sNhOm1IRY35KFwx2Ll5/+hJM1VU
kJ9URkm0JOekrFmcPWC2NpPSP3YCFPIVZR1X1EzGaZwHNZ4FN2awb3PE2aIbse83
mtfKsRVqTdKilNni4pV+/r0jws0o2oOs/A9/gyAvbaLIEFE1DkEFiUpM/TOTrgwH
abVFMMDWr5up74nhs7OR9p3pG6HtfjChKsPwN95QcUtYHdtzH9qmAF7Ff7vFidgp
1N3Etn4JeTJjjh/utmdw9iVhshiv3Uh+2m/3qx8D3sRFdoPYFylyjG7/LxIsuduj
38p6LY1VDepx9L+7QZHXTJvW+oSVWXc8kNCiym7i3BoTPdvEKXUZB8/FTj9QxcQR
t4werkhyE+9j/icFa5NfirAq4vA1ALP15Bqq6scUTvZ0u1pBdRkv6JmcJFcdTIkW
tbe7son/4EbWllXKC1neLGvpF51QNUD+saznJxDMJQR0hsGbHQj5vIbpzl13/DaO
tP2pymOkrz2fIzJL5ryBAgswlIwNWfB1apzn2clOrjYY7XgmYHSXRy5WcTb01jA8
owy7Ke8fjceJ/WTil5gfNINqAU9Xu5s7qvPzSji3kZ+pe2DTSL8bB5RHOOZQLBw6
1mPZK/4ij2mhm+Sr3syyFpBJVjgtwm9qwifVXVtRH7liW6RBxCYwfDicw0xi8c8J
WcF9lAj2aRmch4ho4Amt8C+NgwYcIAM+KzgMY0l9ZQNrBbZt5Qe1YBlFArTg/6DM
jmfomY0ulMUO5VwsuxZ9kabmESvr5xLl29mIRXddDJRqtT6tUFPFOEarU6KM5ST6
q+Qr/qgTTh2p72deb03xGT2Qx+jJbGrcVOmEqe0HtyrgbWYWe7NCabp7k8CZCU9o
RE7wh2CpGfKGeHvO9nKnhCbQ7g5uz0OJqRNkqViySybx0zL6xOiColRgyn7xm1xb
Iylp+KsVcCazZoarmHsmlCPUizzf7mPBX4sl2ocfZU20dfwrDBpcxKPJRmoOQ2Ob
zhnW9/0MlueS3R1IWl95YbjTm3gYgTUcoyI2XaC6f7ITMW5MT2FG3LlJci2ZccgF
ZbOyU0YK5G0IJ5ZJTyz0WqinuCmYfCGfR96W1kDRlxeJdui9Ln0OP/PuvGLA4W97
ftBL7gPvgC47KW/uNcX9+0+aM4SDa3bzdeTtHE/iRqorUoP034UD/Mc49LLoa9Tu
hs69T/k0LG/WfA6HxXkk4chyIr20HSkRVfS6yWNKYHqRUE3Z6byF7CJN7SFCv5j5
jc9ge8fA2j+ZEQ1Z6dlCWEjXfXglrp10dKA6Exg1zVH6F+D67vfM2uRMWKJV5Pg8
O/0LFnxFvMW+FlmC4eSf1+IvB7344aMuLbnzzyeGhdwsvWXpuAxgRbT1t4X8dseg
kOymJE5s1n4BcqX+nlCaU784t2mFAkHR3QrsrVOQHfSW93ZzIm5QszagFyYNEcVW
YDFl8SmODkoAst89UWL6HQNwuZINXEVbj8Bi9Y3ogYEj+dk5S+TOaa6y7F+2sQD4
EeBAI6+2xfr5/evQlevu72kk/AMfjAm1EDBzO7jkxyq7NVA+mBfR2TvCax3Wxx01
DYhBg3/AI6khlfD+VviSLLEz3itSMcK6GeREwMnwqUOPwhonDrXjCAr861j7h1dh
QWrqPP2nbFuAgaF0FGZGEuwN6m69wIpKuwmHhPEh7dn1bBC2tGuqdO2lKG0Gg13W
bHb+eTJHZpQWaB7tNCkMQnaro5hBgtCvxWZNVwomEmkqfaDpptC+cTIab8X7owbB
1oZX44kwqUv1VheGKlvXyNEEzZGT/jEbYnGE21R4a4kd6vip6Nc27jgnejNfbyAA
IZ/NO4kwVzfTlC+PTuHBsw6bOQ0jhTifwbDtr6lQk21EjaUFg4U1uw+FNQbTMPSZ
qwQB+hW+TcDKSHpIeK1hZZujkxeG7RfQMRbhbC0iY+wcB/Mwxb85u7q+VPZ7EaP/
jV8rHuhBO6duzpPK447RVoaeDlDo/6kZSkZWTQSwv5MAYpJL4caIgZ1dZjC/SXsk
fiiOwt0Cx0IngbSavVwtk9aUieC00pCDHzi0q/4ujwoLPUlewyMy0/hBrdomAriN
9z957pCKxr41zbJep9eEBbxxWz9ISjMH8HEsdr6uzbe/45ulXr/A/Yzi5FAnyqx4
9H1czjn/jPP9F8HMDa+yQPvt7S7cQH+0qWFW7KicWj4jqgdEUh9YG1aYBf4rfrJx
bYCOgbR0d5M/9keGwXnYyfmiKZZcEqr64u2gxamF8ddz/SLhE1f0CNA5K87gMPdU
TynvrMP4jeZHtNT/moTtL5FntoW49hDZ1J6xD6js9n3fFbd5wR31oc/MLaA+1M5m
29ubSFVtNcRBjDJOKrHq3nNwtdyj6125NVQn37F59UEP4j2ZN/745VAwglMmZBev
lCvTRXMlisyaCqZCQEN4C72flXDOHCMbpUd8meKCt3gLIFAYQnL35uQ0ktQc7tja
nUoumV5PNHj35h32Ajrcxo3PgeVR7xgII/s/qnZ6ZIxDleJDUU+CPAaQIoqUJr1p
tVvlkFa04nUpq/jf3zSJFNsXkTPJy1xpng0IsGFtBE8orz4SNvRBpbt7sS9QDfW0
qAOP0PJIwvHxO/kFXOtfkJ1pqacEl4mWgTaIG9aH6xej3oYVfbPQJHnlLVajraoc
2fP4vp00vWJygQNOMFechVD6JxXWGmZ3nKNfvJgTzlR1QFcrSQDTbynwm8PPvTv+
x5CTtapL/Hm3pEaejHlM7+GAkn4y8GCE+VPVCr2gXL1+4h1MNdvMRaKK/EPRG23y
PTbE39t/ldlFgcWt+qL3DeBC0IBsXuwCYsaHfqwdoFmHmo8dAGMLnKDdM9PrxV98
GDzBJDj/Z4R4XDbZtgDHTgP3kWd8Kuj1rJPDNg0LIoYXi8Ug0C+1abCkP0IZgr8L
0/ZMuJRg0rCYJLN1MieBZRvdrgk3WaWv1HDT1sgFo5JZRx9Yt7Zj3CNm7H0JLihc
HiderQMOfcN7QCNJ05P5JOZLDLbK4O8oMv7CTMUKAgMw4GuO0C9px8k4F50hbGvJ
zRSZY5qKC4j+EpY6izY9Tcq6i8oy3+jRMq01qi+Bn1mzU0TFDXopObZtmH1sXgae
rErOKKE6hldGaA7ZWZx0Xow7kDoa7PzD0qcm5H3XjJoG1BbT/ccdUzqVfyhP2Qgd
BzI7et96DWqVzuoMYMDXHjXkDK1pdo8deouUF1KZGWqH2OF+dCoLpJhBGOJDvRI+
55WIKrNmNGMYIJl06ViuBX/TCPrdepL6rsQqquhi6+HAazzkSXhajTvkCacRkeow
GWLKsXsFlkdgQn+2nDC06O30X36RuFj5iHB8StqJqj07JFgPlBO8g+ZDSR7wQKTZ
kvpPA25SB9bBaYROsu48HaUjvrdhYHGquPVYJ4npvEDkD5zwf5/bCFysSP8shHV6
RkdEcfoX7HGBFzxh4Hc8Qrj4ObH+SpOpcQerjVr9+tDKNLz0BUqosaD1U7noruFE
FP2XJnU9S0T35IaEt1iSoZNWNYfSqcQ8lHt6QkFiNVcSp2P63EcuWxZYb5vAghTx
BpQeT0Ks8jERdO5YR9jUzkuQIC6exr9B0mS+hej+/2lg3v4QAVOU1AfRo5IFfZXj
0nnto7sCfeYq+DNpmnLjfJ+AdaZZSFj5jOvUa0PlOb+ab5ZHBYisnnj73xaW/Zz1
iazvstDqQz2DHs6HCxyx5woKfVe0b+YHKCeo94fYdDmlJMv2EQafaWT/LqpsTPbx
CAOJhITn2bDKWAwXLGGEYeHmjrWZf+k7TipCeErPt3/9Ka8gKXSjGlbKeX95QUGe
wxo4uoz+29VnYvg6w7G9+9aZrQWSh/F0Q6Ulc2tDmMVWW44iwsqKh4tpvL+6BkLC
fUk1PRF7EPaqn4JTN8RY5Y4Vr12MoY/iebotXvhv+edElNwmuEA4kVVn1WJxkj2a
QGh+3YqA2o/ad6XnUByQWTk6dGmpglgtpO+Eq4Rm0CABY30u5ip3mNSvRjk3zYi8
Yu8UJaGnC/u3Pea6GhyQ7zbb858VSVJmHbAqcIcYYjZ0YO69XLJU6sL+XxOiryuz
KYUA/za6mGyeud9ireorSTD8iMw6e0B8i+LXqB6m0wqe6GvRjDTJ4qup/6ylQsoG
3iSeSAy+cdVOOC26yyd1t/GwCJI7w2VA7TFVcvDGlYTedMy6hhSlNZolYHM6+PGx
XxuoLKBmhkH5z5Xy35LQp0uo9Bq/52VcpSIbry9s4Y40ZxwshK61dwStMvnx/arS
uTbkoz1cgCuuUReQ3t2ntWmi0D5EL35o0IP8hcTSuMoOEgFr+xRQTqUt8sywQOOd
HhHTvdDAPNebdS3mvtuzu+irL8A1WHNiC9dfR0qLVVAs3s3g35ZmdKWn5Hkd5ly/
fAZSZMd8YEjs+qDXoNLuwKJ56wKAJcMBJ3YltHOm/MobLYEAqsaO1XY1mAk/zhlD
5dw/Deio6GqjGNBpuRY8NsQ+mcdJSif30I0/fwcDIrIqKHWvV7cgZtsDcaF0SH8l
Y2QH6Kb2Ftm9c7houmlxImhWUoTN5YTaLTHAvS3Hf3jQBgRHx7/Y+DkS2ss/DEJa
vt1wIQyCwfpLhtvG5CMTqpoBHDzAQzfCRUk2z/ZrhsWIubQepsB/8r2ZH/a9cT/I
XDwuQ/CPLbmOk3Y8g9u7NRPi6KQjXOLsP1dihbwvuL5NbQ+aaGCLr3uCLSKtcTcb
/l13kx5znjG48FCuY9q1OFrQ3ANDy0ygvX3Q25EfwT81tOl3CrgTcpa+uEeIsC8G
iqHH9WphMTtgYVzul+KbGaJHfX1jUCzwRqvKuDogInRcErs0j49on6akIYm0m6zw
aJUSxeTJwWjimrU/cXxtwqmaJQgl0YEj9OTyiOQ39Uoz8mOJeDLaMeBv8oNKqzPY
Fw2Ke+rFO4qw/gdwYwm+wx+PZIJdrb5ej1EcAwH5dOIPWmkeU7iRhw13yr+lYA1K
5bUiaMXl+KlMSBu/1+gqKXnrMjwAMWcR8yOp2Ioo64rTKbXRcj9lvEpfXgG01K6C
9SGa3Ah4nkP90Ujrdx3PwpiTxOHZKINIf2epEjeYEehWDFYBmRpk5dW77UvK+ytZ
Tnte0BlpdD9xbN2DePNeEs4q8KTJv4n+mKPabjMD8540qbCQT2oG3S6MKF7IrTmn
WAluzHHrqPmohPFBbbbu7vK1uY2C2ozJOM4IlxtUHzcrAqMVTwhJe7sa0BpOEaPQ
lqA3B4mKBTLp/Gu6Uwgg3Y7HLDlIVRizFzUbsmmbwhy08f7jxYM/aUD7m/Go1jFP
FyA9FvAwodeZaqV3HauvuhiEJkQJVB8TxQvXi/pqdZ7lT0gBJbXQWVjNiPV7rCet
tNSkYtBfyolIMmY0ODqw3mkk3jVMpQDY8H0SVw7sTQ/cWoGaeyNjJZ3oV3RPXBpl
7FnQmLWwBRnaDsrVdsW1rS9GcnyVNdzLGqDB6vftBEu/W38AQxByxdoENzTati4c
FLml7+Wg4LCx8jI7XzRuIaSiuCpwUGUo75OQwgwEbfl8tNXB6vLYH//YHBeA8Fqs
aTzHT/IHtHqQl5nrUIdpPeR72/iGSaMgZtg3S9jLgtROWbnTyWt9MrfgMmaAwTVX
S/Pm3bfKXJa/pNqjywUuwUnFH2tmk6TYSn8E3bzliEC60j+9vTT7dUorSEBVi8rx
dMpQubmd04i6mR3/NRtWPns3mAt2ys+Q+geQkmSk6veLqGu+d2fGTfmKxSefDyl9
JAZ3GDrBUXOWDdx8dmSq+WbtRlHBDI2fpypWexKyHx1spWxpjMLPDzc6kMkBgNLq
LamsYi7yoPnbbDUXLXjirgGwdI1mR3G8FMd05HAGTH2X98fLxMEFNlYwQ1dCfrnp
HcG+FAmAle9tkXsnC2jiI55fCT9jUv5XSyPPAuetrfnWyBAxl5+X1J0MvnazOTHx
dOoLwXemfl+iTaKt2Zz2ukH+2e4o4bJEcvivi9U/OKBycdXxufONG6UDmBBRLdhx
SkGB1LygGvcLuej+X0H8jradRsNjF2zNypIyp2tgBH6IvJPQBHV5iqw4kW4F+2lC
hU6XoWy/c/zTLffZY5G1if11mjvB6fN2v0j/xJLXQHf5PvFQC6TxKPcQ7kTw5rts
e9iqK5DqkayrLLMGZMUxs1c1Zb9NBr6Jard1WuKB8nL8UuD3uptPurBUsR+E/Qzj
yZbFGPKNI4R/aKXFrg22HkQNEDz+47N44xR//XXsuVnIu92eovYp+MPTbhgckSnU
EHa4tnxFrcEYSsClM6LzpnwuIdImpbuKhCAMLe/q93oYKwvbeWEusf+3SPTk/AUA
ol2BhpoBAvTh60UZ6ja+/4ZayPvqhxsL0FO4GPIwaPp7KrOrGMwhDyb+m84WQKJV
6FMyOAmkp1HXI2YN032nXV0Hqv+ZujuD35gmvh24HqNCanB4JTX9WjGp4HQi8j5h
F6MRLT4849Xf/ru5atstuNKSYK5lZlvuLmZMAqIungB1m4WybKRi1AKIikiE6x9U
QRYn7R/+YjgX98ibACznpG6LJQoExqRTMN/cq5qo+RrY+CP/ejc+R6N/h5QP55G+
HCEBUxQl5k4FuPsThLQVLzQxku+jPTt+Zg21QQKPIpy9F6PCiiSt58BO802YQ86q
1unAepLjN/RkGAstW2KnpcpVljiE8NxQ1u47xDiFupCKeJCzmZMURiLq1JTrTpGQ
ZAU+EFuyzCTtXs/sQe5LmeWPL3PQixQG8EyXGPJxKWUeXA3In0iBOv5jXygo5yi8
MLjnYiHv14VAYcxhREUofGP9U0GvUvKBva3WD1BG8diWNM995ndvS9c6lDXXaZ11
LwRA7jZ+bMLfDMUIierfT4jpWvJkRpTr3sfJPw4gFp6wVUKM82hPAzhbUBvsj/xd
JQBvDJpVjD86TUUzCDyrlwI2nqMKzhkrDGjHy+ABzeIXDutMo/bsGhfFt3r9zVBZ
QqNefM7Y0w0i1LPFC2RB/g+9yOBjC04HyzN4P2xEnQO3IdBPbH8baQdCZkjrwao6
8Hlcikd7VD60WEv+xRSFJoix/GexC2b2mOOOK5X7KkCr8eh+MCZQpb99Tvrv8viy
BrCdjEziNGrSMmP6HIWI3wTZC54Z8Y6sT8e1wTHQGRz3Nev+JC/WgZRo/hQMtrEI
87UldPyfgFDtiES5zBHCL1uMusww+eiAjYlvp4Rkx0ilOy4lOeMnZMit+MF8tHjX
Iap8jgzUgkz71fKgJS3/NzIEQVIoEFazb36XTLfi9PNq1AiZrJFjls8ohHfTI6Er
lhs4jK0d2MY7Jyzi8qix9iMSCsRF1QmcHmEPoQMaRtU4rdnGZEXo53MXqVHdFBAq
w2KaHeFBvKAH1QU8QjT8TCMCMc+UbXAJ+sUP+U9siSCyFPSf48Rq58DithY1tuPl
bRyi9sSYpJe2XBA90VChzE2vGr6v4ZloQDsXA9gO0Wzmj3kF3atpyqGalc3aziD1
Xy7e4B5c5zB4qVyOcR9/0/VHbNWfDeE2Hl2TVZYPxYPfbJ5KP8SP02U6rRbZ9aa/
6GNsttutAGkzIBLIX/KLko33HPPO3I0hCESFPe/FUZNbzzH+cCjeGSshazoZsqsV
LyXc186MBpDdCU+vsyVsqFhjCz74mjJDSHtukY++wongHjlA4jyfQguMhvAn6dMM
ml62A8KfOcpz8HW+q+9cSPT71jZH/WvtDVHwOzCRr7n2E22nsiNpG+igdTP10hF4
grSC3piK/8BDBG+sawP4W3FX7SyyfhCDLqeV92HEQ+kLwo6F6w12ZLDPL9GfRf8u
sFMIyDyZylLVCa6uuR7qeATdNp35UcoFqzSYl0YsZlxMUW3uM9wXlPkRojSkvpnh
h0HEFI1/N/SeK//jEA+8BohC2btTeXvTyio0Hx7V8Uyy37y7qP5LE3dIOK0fUkFq
zKmsH2xCsOX/RcFm8wAi3/o9cAVOYnk4SLnUPtfCMq+8DlRuesoYffdyOHa3bbla
88nXVorDNnNsVSQrGMcbiaFdbTitK/F5NH5Sm/gsfjVXowlm6KFrUNKDobIM8PtA
s0Ge2ZzKbxr3DD/5xfVfHQEwHNChy5sYif3GHRWGBOqHuEfKCcLG8euDwGVJDfOE
JHaHR7HceK9zyJAWEFtELaElGXKqi7X5qojF/taoQDLSVaKVOnHtLLvHwoDzT9JC
4/Dblk1+/3mEIfbCJioinj2n32CmHYOLJONi3pWFJSspZgbcltzlUKgab77bBtaz
jUbLF93DyCbZxjbi/OxSBBRC2yPiumajBi8G8q7hG8P4O0Y7lvtlI9tn8+me5hTQ
5x27zYE2WO0PzWgY5iziDJO/U39NrEXZ6tpmw5Hf3VKwLjyVx2r8eZq1yCoOuTx3
Xv6LiYJHFKDYOGs7JxBKzdvqp6jpcdRcYWKzJI4w0A6gWtBykDAQ64wwytt9bVee
jJ3MDVWqjLY8/zizjHbX1IHsid4SBTXXAC29bTYN0pstA33/sHgLe4fKs6e7X8Xx
4L4HEyN1FeDBstV5t255kOyU4YQSPNiiU9P/j+QSkrMwMCLZ0eyF4rwjeCGWbpIF
LE1MU8PjlTTJq2Lo/c4LQK3dGu2H4TH7Zy3CwAfwT4g=
`protect END_PROTECTED
