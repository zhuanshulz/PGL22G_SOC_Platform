`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
md/7PmGR77ysub20+NKWbKAs/rkNvId+C0cyrJcqofKTIS7nxYuLdWKldoH7ebwp
ADx4F5HkoKbGufY2cOlOVPBSY9c8P+bi8A6ENHuOd7bA1w7yD2wRuEVc9iz9k183
I6fMd72b3+tqQrCiYD2CUfEZ7HmZ/fL5I776K6Bp45O8+/sOTlVmL+uSYhrbgHct
ohozAMaXPqC+sAiw6ElCJtjH7QEfO2BtCAvYdqAdCr92ZIAUIXgW449PtWJDhDgC
V2Cq6NrA6+FshDLv6UF7EFkyKJeyVnIdtCublJBX2zoyQ4r+EgG7jv57x7SiO6/I
V77pqhska+lDvUTLKebVd4RIsq8tcALaOPLoFXGX5LjrJk4F0TbQ3324Yo9H9GbE
+WkqA/+g3exO/fOO5+1rcg==
`protect END_PROTECTED
