`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6Q7+7NhrsNqDDPkHJHl4W5fR38M2DjKMB7A/Gsn7GP5pUpxbKASg5WyzkFhHK/L
X/CMGr0gzUAzs353QBiWurNtd0EguBRFZ5T6tTA5h5Fn/sUa0fLdmPyuO968cYJ1
tj+z9bxTcPKV3aa0K2XSPPkzsfUD2d9winGS6DjXuJagiX5iTgT7Pd0FwZFNgPie
TXVmZ0YXDhkpvxt+Ar26G13X+7L3AGyHO/dXa7D9IGjCbR0SjB24lE4Djd33xkJ6
1HGlNadvEfworsIfZohozs9wI+ypfILObaTNFVx6WCXrqK/ceq2kSWkxaVr0vAUt
nd3EssxMNwvuuzuTNU6/5/MG1TnhxhBUvvUfcKb1bJAHKskNya7M3hDZbLj5p54A
1hTLz7E9i2NIhxZ395H9sGhpHsQCwZCXaswrm9YeEAWtczWXGovhraOqeNvop2m3
Sdg0Zis7R7ol7KYuEYqAg8hQ8gObsiWtS0cWbVNdmWRJlw+AF2p/xsCWD8SCAvC5
3ABHhx3/S7BAuXKrz1h3SXxc8oKWLQ8DSn6waJcq2Bk4SpXpDvKsSewr6y6YhDiK
U+quZaQCt8583mS/mQD2hHS8Tf1E40UXuQpy78bEyrEYcLaes8hD2WL8lwCfUVK2
Wh0mrgYOr6WXfg5TWNk4AHtlM4iRvbspbvYlgZQiVT+I0B9LPSc2knf2LHv1KziJ
Z7kZdotA2SJ/qzm4KgFuhE1RLbe21UqV8UHb9GNzW9sCY+/cVOBRqznVVepoAHQr
Ib+4UDdHXppo1B4Y+FAUSdOoy+jOBP0Of26LQPON47f8BjUhcortjsoT4Pe1JKN9
q+Wkxkw0iKuPmxv87UtG42p/JwNg8rl6yUPdU7MOn9z8BOVPX5ccXg5tdcF832VY
hh+5aZ3EGZqAiTqDTLY7NPR0PyvahtpNAL9OxbqvD/Hf+LKlrE17KVPEHHtH/rVy
9PssYbVe/n82kS26SwKj2qHvuxyroI7ekE28y3+VSObMRSh4RsujSkqBqDn3LbD5
UNxZZB5py1JJi3lmbL/Hk/Maz1/QGD3cW4xmRpu2v8zR61siejkCXz7OBi18NO/B
rpHeslUtd9JBQUpdKJsJWzTHbz5fdGBCDPZDw3h+xUttjBzfofLuIHUwcveF1zvW
r4jK32sy2NwfpI9QcTcFuoVbXagOVc0MN+cl3TfVTfm1iufSq/vOVW3aawqB2ru7
bPtvj69Y5dJo2TUm+T8tkaOKq8FKBNZcSwlZz95Vfue9/tTVAuVDioVsUpJm4w2v
`protect END_PROTECTED
