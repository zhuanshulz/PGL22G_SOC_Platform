`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vbPzDkMqrYHxSL6K8PHUy2Ezkl6TNJ7yBQfEUpvAPToe/DfXPb11nybdQ0Xuqsp
BwX8k0S5xI70NUEqRQqKuu4QAk8wJXErAVlNHyht/HBfA3quJZTZgQXVWR7FNd5k
cbhV0G4OBhVloJU1ccWDLtY8FRaB6sQiG3AZHnuUio7xre4riQS2E5fTf5wvsh97
yvyJiyCXID0rMQtDPBbc60QXzkV1AMEk4imix/QyRcziAbrX1UiWFuneW271+E7x
rvN7/19HiHqO4XoVsCZrNf9K+pimH+tpQcb5/pep8Z4Ny/a1O2QnUebALzJsTlGK
EhkEKFoCHCFg6/RZ8ahDWU0jJ2FGuQdsLAZ3cyhe/dpVFeeqzAiISQG2OuGbR0sC
rPspnIg0aL5CYvh83tlRJ39cepPk8mSItNk2d3CAVz9djozQnrQxW6ylG4yS2SNp
Eh0V1RlQPUsGu5t80NJHh+TrKfImDbbQF9H4nMepFvSyGb6f5KMYLx2/RVWZrW4Q
yCbjNjuwDeG8mzJg/nIAEXamS8T3tFWnJIWU+5330GbdeQNUHUhyQ2op4LKVJ/8a
AyzpmozeFZJBGp4iWx1HwY5dF/1uTq/4/kTWd51XRyggfZnyUOHag89WImxFP8PT
fAOxvjjX/q+yFjXyoFgg//8y/z06dp8xiC02Lyo6yirMovcF7eBg5b2pNLa8POIo
CkaCVKd4EHtOPkW+XBurFFzGgksNGzwpwy/Mvy1aLvVmfhqYDnqg4wndRDPXmIgr
u0BQhDMHcnVYrdYUmzg3zETFWEQ22mVJ8Q0x2KUFVBF7HcU+Mtge3Ib8GJd7Mywq
De6UfUgI5Ao8OaETNcVuyU3bOSjVhlcKmNXqdbTpdDOLv6ryC0TF9+qWqZA70jpV
/2HTLHl4U1M3tZChPuqsbAqWOoPNsaXJf8h4W5Pe5lc=
`protect END_PROTECTED
