`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gYmc8PIGOMMcdHJzJgiZeqO0W/WOo3Q0vE7GDYGjZXJlZv/8+MPnlR4wNHnC/swS
q6TOtQYLUOp173bu5XiWP4A5M2sCPvzCaNL3vAWzGOpMMOqzq0njJgdy8blgvVHc
AAPoFeFyHjpChBYSZ9wZmZar2iRxtPHeqlg9p+YsQdf9s1yMfP7W1zPCn0DK/4EM
YvQXA7YgzkuxbmmmQPvqTLS1SavdyBin7AWHO9pn7L2C05aYutE97F2TWF3tzb3w
3YwF2Q27eLWwmrgirgwKpX0cY5EFiO+9U0+YH7XLhXf81Kyg9HfgRbXZ8osJ+7Ta
bFytUW2TVjMCCz9xGQlP/UO5QMO4ZfICP0e8sOA0r3fqAOS3A5y0OtbrqJpOUfXr
f+D84dOGqPurhOlLIP9w+AU74fbgX+CRYsvlUNAcSbxcNN2dCy+hPz9Jjyrd/Mcy
+k8bhNpZS9pMXLFm7kZ9pY24Lf78C3g3Kk7L1NkB8A5EjcsjLchnJ4nX5HgSYIbC
NqS2DyH7PsrflOM5g3WtSA==
`protect END_PROTECTED
