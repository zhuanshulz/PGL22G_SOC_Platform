`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkkO+VwdtD/hXMy1POpt30J9vGcHe4eeMCw6HcHbp+JuPkPA+ypKyyNSPrKtX5Gx
6desp8Iu0ucBNpl+QQbYXN8toFeB7jeFx09jbx1eXfwOHCnGbvXEtIdL57PF7q2r
vq/osF9y1PBPxYmVNb85fFq9Qa4PjmamC/rlytcng6X0npW8RhWEUiCW/jRtba6j
c+Kk3wU5+t/7dbaTymq7DDBwkey9F5xY/b/ao/G1atXQoIh+MXle61llG4/wRXiu
yJCttk5QA2IozCdQVycATopOmuMYRg9YLwwAH62lRH3o7ylvnF0vgLBVvcUorUNX
vpoffeJGUX0nWRKjY00htEu1Jl4gxAPTOpV0W5UbK8bsYr618Y5hfaPey+zi7mrG
pkGDoFGkzUWOApsimxVdyEqpZkEKrP2F7z8NHbKDtjgxxsJGCi+F6skb2da1tfOe
DYyIQws+u+EcG6QH2BVGLOIL7n3jskkqKF3UChg/2wDvHtIfmY945be48+gk/RKp
4gI2ks5i5uYHNJY8BVUUoftAYsbukg72QWZZJOdWtF1hDGiaOpQKR2CLtuAe/glk
d5mqi0KSjfoirid69dlSi95byhYpsZrHck/NBAfNJ0rTgwedqMvEmaYXGhvZxra5
//N03uDREo0TAgG7U3SyLI2+d/vsG2tW7i6Se4w2bM7LhcLGpmZpXN7SjFskK5RJ
uvfSRylL2AEkHu11hyyWcTxtHEmQ8vjoMzrM2JlXL2Xw0YFgBTcyTWI0vyvyHDNX
BPGIdDkphK3GGneBe5ByZMxXnAG5ApT/+Jwaake92wp5Z1iYERIRfy5YdmgHNHDg
4/rlsP81340VOgf6xTchABHNG/MslORONLUhmLzFOyrgQz9dPf/+PT1pOrDpYsLY
cM0QuO2dgQnuNyCfs5+k0FYsdvwC+znnJoV0U7APfF/B954tPEexmUgzvdpJMM8y
Rkax2POivExDZfMDnHwHTpMLsVyLsiaB1ohDfvsTH7xvnBARwuv5vyG50B7sQUDe
YhIFlZEH5yws8T/jB0fFbjyNSiVsI0MIPfMq3pWnunaVtn1bylRWe78FbrgRF9Dn
qzYvshur1U1x5b6ievpOje5Y3I+ZlfZJYzapgQUeon/7sSfxWV6UgQWTwT+aU+SZ
N11S00jQpS9awH8ght6GI+QvqVW3yUw5F92t6AA2NZphfsmoQnhqVfvbgZhNbQZA
QH/IDQna33KRBhpac5pzYOf0YTLSBRTe2hz2UjlMGETna5CIz35Ax16RmWgr4jlE
JsJxm5oo1n+q7iSstLaXNlDX7HffTeyx58wYGa5QfsjVSDY1S47rVP5FhPH/FZfh
nUraI+IGVGI2iuvhYgI3/bapYI7OqPBusOzicTzlNhV4ws+yROUww7QY9wrR7pRx
ji3u3VlspCjU2WUs5V9u728L73qnBOEcIFSaMcpvDnHeokxMJRnBavoFtBZZzA78
lPrl5eAosk6VX501Ue1BhakQ2HIpBWwVTYmIkg3vXDCKnRfyxOfH8uvINTWqXfn1
YbdH88XcqLkbrVtzaEiirkUYSRLOKdNMCjeZ9RxQGIryKoFvxnn6zP55elB8LXb/
4gah2RLf72cboUdHMF1Ak+RJ5bunqfJEYwm5rti9XmrV3Z2iDuadvvLSqtvJa49c
ZbjSzl8seqdhXx8E22pOwcGrpm5aqqzouRjIKofv7jnHY8tIrDkibKMji+Lo8YNx
DCAq7cbp5z3V0UV1lClhXnIDjg/Ns3YHOKoSpNPIZpUzc9RIeZFzFj1xdMXIWXm6
6g7SvyjQYE0fitdrE9lC8sJF7a457eR/1jNOEhESEaoLUaCkaV8PkqSr+w42/M72
DKSSWrPnqm0C1tdSYGtwaQ/cwMEVJK6KcBNY0TMGiv0r6+qBuuCXOoM0vT4i39cq
DzrvAbpvFJJCG6QQmUKNkcT8txtDGppdRQz5lRuTEYWVgrhCm9HD+AEpQzi25QmY
ftKwn73w0FWjYwQFCEguyP6r2wleORcUXGsXkSSBMrzteMDj7lazqI6QvaW75Els
/GRneX8c4O7qQcJtFXI2t8IVFIT2I29XekmLKHuMLimNPGtHUZ2BuxIRWgSpLNUO
6TLtK1YH3HSlFM8Mvnf80A/30dVTU2jPB/+RFgsiNLmhHNsPqbmm2XwZM4ZU9ana
WIXFna5Ljxk4fl/lC6vsto4HIAez4E2vogjh7AcXugsKtFKkhU0biet/pYgN+nm1
uZFD9UqVyyX+IjzpQ00UNNZiDHW7Qfk8LJ9O+6gl+c7ec/5tzoQYLQfMhNZLc3GR
fFgS5A0eL1TcIaSc1ebLW254tfN+STFtdCYsd03IcXl+ujBq650LTYCulRXbINGt
nYTktGPb01a310ZPHjiH8oRwzYMZCSIsXPtQ5mrC0l+SJJ9o3HokzSllsSLJnQYy
3zQFpUeHfSq5r0sZP3MuMFxmAQC6BcH7IkM5cGNDHKJDhCo+HUFm3Zg5OZ2Bk2xq
Fl6mdL4Wkzv6qib1UHx6mUMQb/bdS8pU+Dxbj6efGRdMq4FIql6J/Dd4JVnXpzrj
xWNAgTvrsFZBgYqLno0wkw2lxVUHSMVBVXiXL2vULzWqe9ZDUB9f0HGXILILA1D8
mivTk64qK7jpclkQXsUTBEhiTBCiNbGwh5a3rfvbYdfr2l7Th+8RIcaJkT9ywdXp
bkHAlNQTYZHyQG4zUzQi+Dbr+wDa1tUbUWtCxPWsP4zYmeXQ5GhCwC6rCe4vnBwy
9LUK28XbSCCbJbilugps3mGiFLC3H/SmhCGFXadkXxCawqKh7fQKqf0gDTE9ksfc
YQ+qMcjjJ4krZ+/q6rtYfHGGMPogTV+8A6Qh2prTZlVqYhk9AyWxi4fef+sIBEHQ
zYh2ulZCTwjC8ZftE3NXWc7S/SAQrf3qRghQ3f5BJ+00AiBnAuncY4VMtZ4Q2rsr
WvoN0Np2ihsf+43z70yXlx/wEvGFl1X/Q8TExGuhvQf2KEE5SccJHPy6lkeu+83b
82XPKcZDo/S6dKTW3OFgJfIMO2sWwY1Bx2EogBd+dMcxuHoz1K9c3m95L5avER6D
QY7rtMIlnNn+APEsETAKBCBGzlGKtPRwvSbNlnU8x+VjxknwT145jUkTdi688K2G
ThfrHN4/b6UP5HBaDhYJdi7dDIMJrDK9h6Xl8lOKLAwW5UlYZCG429zjFVOxC3BI
HD4AHHKrtGi/CoJz3gsM8Wvgk3iTGjluVUy1lgEc/ufNk1arGwhI90E8XWvgv5vP
SvtUG7pRUJclmArcOpGgkLbPY2g7b+CtCXtnkyDpMfVslLlA3t2BJ9v1kzfhNwtf
jtFJPnZZAijzcrQRLs4cVmHVdck+TBla2P8e4Ke8IiUF2UI7U9S7mp++MI4nlew+
G75tYYk2a87MstudizdI2eKbQPlUKN8huDHJ1nA/aActP94eRIrnB1lnELixjQbr
4ZgIwSlrShoWiaDAZWZgP+uNnkBCyDdT0PGaCG8oRu8UZPFH/+D6W4WxLK1dUgNM
SKQzP5kpFDLYfF3aLpmi933CI0sAfpEEf5WZCY4vTgyTq+57ldIQ6gI+3oU04yzL
SovreX2K4YsAoX7/ql1GvDNF02pm8Wsy8GXwU/K9jZT479ysP1TQ11UgV/8qxqou
TnrJmzXN2LJ5LVhMR/O8Jeyf9tVnTSDFYZ9tDR0721NWFp8vVP5BJ8gjr2NHDGdI
shlF16W5GFsM/8h5HdfQMCjBXUmnqhboxAyt9zg874yWV7bqbAN7cdUN/ODatzOp
4pUlaQ9Tm4EdwtXKuDGE54hZspAlOrsh2rpJsERd/HZLY5+DEh7SZ1wU+OIv8VmY
aoDcaa+uMERJvrk63Lzr9zAfchHV+LKOkVu7NCo7XNmGU9zJrEXjKYFxuCZEFMyW
ZIvzjbVpWGtMnnCz2HIXUFPfcEswCyxaihHmiSTkmixMxEUBFf4O3nvbtd8/xKIu
x6W2ZmGuj3ozU3PsN3OU2gihv3NLF3IZ32FMWnih2xbxGyL2At2Qls7PBWML4mOU
xsDZRGPC+fnT5PVmBQm35yRa1V4S9S8n6Xrr/BNzSeUnFM+1o21VH4u/pC4I7YdJ
i9YxcEV13O+3cYuVpryH7bKpZeaXd6aW8MkS9OtpI4v+uhNxp8Afgz2WNyjQ5DHT
7fVaFAELqfUkt1oqlRyLBkxFhOZHXBk8m4I9L2B3tFJOl8dEXTqz1mVA4VkwhRVP
9PwlTSY5yT6xEAbS3mdf7/xOgKDEeJkQptkCo3Zg3L+ZwWpfjGXZhFzPeo2U8doX
DEg5CGgrLKx3V0teH1C21pEnmdGkHAnSR/n3jE/y0Pju2cQAemI4QxQgPnmzfqpZ
XNEwGbSAPvjmY/GRR1OLElCmBAOGwVHhzJ1shtfmGfErzB/raF99nokImTV7zvDY
bDgeFIs5tNvjE0pOC5FwdBldIjiH8PZfD3JZg4sYx23+0h+Aul9veduk6dLYcgUK
mYqqyksMoAliLlR1zVZQWRisj5T1uGGW3XQDaASbEPgwONYWcyC7o55pUC4/ASPy
gQ9OM5dNA+I0wDMSNygDzVH0qu6hGfDPYqSgP+CHkGlWAbOHN+gthSbLo24xV/Y2
uNDIbw3f6KMBATF4u+BmnUDgjTCVKJTgfcbGXyip+N+PhIDQU+RH7zIQ+LW918LP
Uq6V/nMe5UO/tyyw2bwbh02yRLC1X5ywKfAwxY4Qb7GRJQ204PR8fw51DlZoTjgP
7txgBJyKiB1vanib9nx2iDjO12LgA3LbaUa/YbqY48Ctwg/kRyP58kRx8j4ROJgt
GnuiX+aaOq2v85M03RRY8hy9KeSiTPSrc9CYXllfnptr/mg2TCfslFP2m7X7Rn/G
ktcHFWX8a1RjxMFQY+zQ+ZVUniG6tM35DMfXuhZV8MVMqVBDED3/nnojBeNPmYT8
86F4CUimeR9wE8E549tjIwJvpE8o0TYSar9ZwLQM/bALZyfI8+NCgCfuIeP0y7VX
Ih1pzI3K7uqHeUH0/+o0P+fxJnvZPclTS2/RgiJmzRpvlKRmoCm1h3qr7wlQOen0
QfODQhkOlTYO4KAcCrELq1wSd5xerRwK66QFdUI9pTjcURhra22VF1Nh+fkIO8CY
I5tvkNDH/fDoKhv3FPaXYPFs3eR32moFuH3Wdp2a94gaIkhMxP1wQSeBAgOgasFt
P+7jDjQQMqyZtMkDDN1nMlGQSyoPS5vpPWOGu9KGH+xVyNbUuwk/SFXQYvTrxVBU
HxPmvqSCTIBX3BqMJa4flpn0uwp/OwM5pzHvthzyyy/WtaGwyOtYE3mkndW9BdXb
jm0ns3XnCfcjIxEl5bkt3CQQcc7yFV8FORah73DP6YmHGibe49Tkb1xFLtRgYmWm
iIpLXDLNjbOd2N+GQAiKGlIrZGYdByglia7b4/iBJZWp76y9UehOmKtC2uaqGpOR
VCrRCviQae+Cnp95a+VXLu40DgUoDuyw3L87ytDg0w+uRbdCdNtMvnefj5PaEKG+
seTxNyUOLp+OeHNgGdkFs9ZE5ogL2DCrxETNVOyp7AMT2fX4TKGq8UfQYjK5G9oE
OO1/ItoOelKW4bv3RoRKA/zmTzLF6Usm8TQcCIdGGTkuKO6gypeVfqSjvGyv/COF
FaMZ8WMhYQOcScHumrGB6zaL48Sx9sfrAgVEE0uoCUMGZfeIBb5hKTniKO7qUn2G
6RTUkjUnrcqFoA0cnikx3dF3wOXvW7hSrJ+FDGSsr08A59B7xmmySiKC0+t2KCq+
9+lUL50MDmo6WmPreElgU1S/kBmdWJ9Qq0TZ42CPctoTit2uPgSsPBHvsa+4qkTf
uLOhPZ0DosTU7Kgwfuu34rHm8vXSVUq4QZaI5Y1YmiRnPnVs45KUmW9Fc8WFEfk0
fwssUppXGXiWObYhOrNQt9mcoB+J3Felhn0QjdisJEBLRX//k7G57ZQl0xFAvCrD
AsPEf5k4BVoi/lvqp4PtFwtvBSn01JVwtPGySjTX078xpi3+0PTgVl2HWyiYE1lX
T527v/hzWKZsBTXPPK+tWvFRtojHN3EdKTpHhSkEcWn6lawKhfSw03sXz+XDUESL
AFYxJBkJKh8bG0CQiic7uHiuhKiSlii6IMQd8q6VYFtSbSBof9MTWg5Ldf3uIkO9
U7MOY0AZ4P7zV1+wVOVRuw3aj2r9yNEDOOXjwuZSt7PuCuDFHSCjjMd9cM/hzpFF
VAR1A5xlLZrwrL5xO45/1K0tEj4CWmoRZUNUmJGEgBJwf5dJD6gM3HTPD0MkSGjJ
OBRQrqmhkVjn92sPQIwE6V4/zA4vF68NQCRgAv1B0FI0trHIhfr76IVJpIdhdHs/
9y67V/eutBtpiZ2BIbEaAlHGy6OIrGctCRlttc1mp3OYPRquSUAmf5hPyPNzNbQ5
XcE5LHqWrUiTIDmnDHM/FjNBMVhSGx1DgmeKwmb0dpRWH5MM25nW40tt50QZcsom
TWtPvlEPk6XLyUh86XlAN1/qaqwvyRsVuJyZJXKB2WRIhDzelSxzB9hT9BASWmVj
ZBmEcjOEPMOHU5YBgFfm0zrm6l1O4btnSYRYYrxOZWrogVeeIGjQTTprBIDKnWTD
3o9OEFaU8Zc54en8Tj5qcZ9SMji3HYIMC70qF6V7brh31ofRymwDHUBHpL3pgvpW
mpQpUiUCFch5prwr0Qku0UUxPihMpYH75p7l6EAWfpuhBg29ZSA7hRxPUo9Fc1/f
bursJ8RspvaZSnfHUjjWp/FLaMmhvDS8ZLhc5euq6sWr477gtHvOhVuPhhYoikHA
DLpsb0xen3rbcpUdBu7bzX+fAzey/yUvDWYi2VshbOQkFCyaYEOnl87lesk3KPeL
yrbqlnPwLThU1ADnYvEvmsj0lQSf+mrUxxytTXGAYTyWJD93sj9i/RczIvckvBYi
HIpTLeilmE3fOAO6viSaCcnwwsXlWdSC13LTs/iGaidTnsRnwfjau1RlV5+pIWOJ
LERaBpfbhqk/oTIW+9CDVpZ2lQhgrGF+NdMiT/Mqpys26DNlEw6ppKaiz+68P6UE
w5cDERzu5qIYpf3t3RkhN7d6G9j5VrJ6a7WYjoCUWhNE5XoeCIt7WLwG77AQae85
glmPIXGz9lfG1myhhzzjFWgIlKogj0hhQbkmt1myoC1JZsAVHq0MO382X8sFe0dN
mr+2LjRoNHpJOrfnKuUvviGoDp9yy5+BBfgFELGkYoSaRmy08Q898lYM3VpQ9izH
sWcSqV1fIimrLHGmhwAkUwIDa9dyFxIv6sB6kMRPFm3YMFTrkqh45pbuE6Vzk7RF
Uzi8BsdtJ0Cmxpt5SfoqTuD13/SdTEc0eE4644w6lnDafwWkFq1F1QlA/n0c9pgz
/aZpH2bg2Qohubo6gmiSiVeb+2+LiMlyHLrleoZY67lD8EHCiR8DVDo2HPJQZhfD
D/rXFkw6vz06R4sjGkOn2D3cIXbTnxfKSXBxwsKc6RyoULFL19V6YraTKl4hWMjN
5vtXZ+y+rYfpLmCv6djT4ZqdlOOc9WdgIFo899Wj0DnSv/IhXvYwDA4xki7tb2JW
zJEztbPdRD4d8E2bxJ23dId1bsRd0nhpyv5I63xWzOH6jT+GK5ABMnUBzDzh/u4r
TCC7N+EsrRicaYYTMNDH+PdrrxJOkFiCpp8b3RKlFGvP+UJXvvAkIq09MjbadpkC
Aj9jPhYShZKOfEVZe2sSr3wjaKCz9lK8ow3GYm+hzfZv4WQhgQ7c070O8k/XekBz
Hrf6oRd8DXCrlJaNxhrWI+PnHqiLzngJgLOcpNAokbl553VuL5Si/9qXOoahEFEQ
hn98nLaHE5O5FTJLSXy5S7p2tsqgdcts0ARfXaYEaSwXvIhwhQUq4GbVK4FVoFqu
KkuUUuzU4gUdR6Sf+7qNx1x8A9SLYzyd9XYda4XrkU3807Xbf9ZC3M6oRwd83DNE
6P51PvvpH93ysDYOirRtcoydMBu/QaUwNtt2NaON1PPMjnqMBA7fK/Ruyy1DpFjQ
RrXdapeRXxETnSr2N+m+KgDhO13FP0OO9D1KP09a1Rs=
`protect END_PROTECTED
