`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aCxLJH9cTJzJZAh2QBzEC79NclSEiCWYuvuqDCC33lui+5unpmtRQ+LrXGE2bY4
Sr0K8l8G5RbzIMv+Tnhjfu2iI6Xyi+fJkeL7C+NuMcko1hrKjrgQsrz9bmSNwUEY
OSpy7MuJKR/ZbcKvh2zshpoYjZotq3YE7ZrAloCCyzdAyWgwRV4nrr9z99LE0yyD
UXbK+fsP6TruR032xWkEGpCDbx35UHrzkW5Sutalyf3D2A4Acn5fz+E7QstFj+7a
s9RSsBVJLZ+O7tNOyWKHif/nHo7SYPzEh5xzbeSk711mswnphZ7SQYW7jMtL1A2M
f7mGfqTAkaO6EqBCylheAWabZUOiA5H8sqIlRrpBDUDMbiElls+586TOJrOS0JRO
xRelexd6aNCwx/bAqg7N+nk1Hqj2uw+6YXHaXgiseQSsm68vQPPF6LRr5jmwy5/k
Het3LnF6vwxrgbq5eYOKGlG1qihdO7RRfxnF7wuxNVuobhB6CHkqryJxZu7Jd8Me
4nE0G0FUv9xH770wu4WvjTdOFKFWb04zB8O2w22lvTRcdQ/6D0D3ank9X9iePlq+
l5yYxP2tzzivFhi0aUO8heLSQApS2M/Dz29jmDYgZR49o2Lalo7GZNyoGddHJSZt
tRGPAtdP03pXTfFdcY6H51mDSYR6NmYj+DJ/PId92l7uwO/FtcQrYkDlLsNrw4/H
G8kXiYPR7Bwf2dRBqbcp5XW8g9zWRVTColgeq+Erkcc9t1H5HAakjXiE8i7hAauq
Ax7c1BFzv02bDZCJz+V0wm3aE4zwZvQ6AH+rVSmjTy1hMRDgVuP1ahB8WX1EFCGl
pMNkM8BzK3sEYELmP5/8F7o44SbLTlXys9sNMdJdi17v+RVeaVxTcaQ9Pq2k+T8o
dJJ6Oa65h9GMbdMemHMtOPc630P75AoM80Wb/D3EzuQir+jUYORVTQBeVjkxGYSR
oxQ4UyKj31A8WV44uDU6hc69/cKDqdzVwiNhETIRKu6xLuTMHBnTyx9mvbG/mZtF
9kAsP1qZm/Dcqz2L7pNGW61htjVpa4LbjX5unUt7r781HjazIKGpq5Z3Ybd0PNG/
Pa1oMrRkUVlKX3Sp34uZezQdJgExm7L5dHF/gSCbYmhU6zhPUiywLgVOPPVTe50H
zNohMko1i+gBfrazTGP7KUrNLNKifa6xUDg2cN9cGYKMYcFXPWzlb5ASIC6TxxhE
JYxHejhgyX1tPAtZP0Ayi/ESGegEW5ZhsXKqZdoJNaLdlVKy6HG7bL1EmRwlgl8G
Yi47MjVxezxE4aSChvimQqg1FBkN/st5z/0yWEaSY83HUX/zpKbozL7irbP7aalY
QhMi/QAmc0wxyrR7AhAzGD/n8jw9JSMY0o8IrYsGo71kwykSoxgeonwHwrsF8ROw
rqZljtNasKiPwKqBqvNmluDl1OwBuMkEX4VIdAXeuxqBFCONI8zk3TZqiiXVuvkI
NP2DuJMJW/YWnIETZm9bveDZi+vTSYP5kh0mP7bozZKBmur+++u8/PIm78hQaILM
5+Ora+ORIZPzy+SRGVttIqQUhnQiQWG0PgocwFUKxDiBvOyuSJUKseSCb2cpyIlr
hmqxknqmKY9303YVf1bXO/SNvAtlUwWgB8E9SBIRERK++vZh4A3es0q45y1k2o9j
`protect END_PROTECTED
