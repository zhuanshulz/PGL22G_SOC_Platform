`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l1Ro6a53M5xv+RAqtcRVtbK7gnEgYzUVpx17692S4CO9eZSF4CNgFra3Gys53jyb
Yv46X+xl+Gw6NqOoPNIMMdrscNXYlUcYdNyVMXtEDredvZhB/fWUfHwPhySKoqAc
xX9dLROuWKac3eScQgoacxT12R0CFS38KTKP/aspCuqjuKb1sWhy0O0NB/vfE0SQ
TBM7nGyeBu0V7Z+HDGE77eoo8wTtMcCzvu3VXk4wJzLJ6AEEjK3frLHIGwOTpzrd
D6bAuyRKsj6SU9K2PUshRROCuLVfU0Q8KiCrMcmzxRpu1tyufiYl6wdNXTWTE7yF
Ir47Rz2eGonztDUGowsnJpR+ZEsG/HyGmu6oDBFaE5Q7P4GBm+Tuj5TxHCXJhPCG
dojsC9xIiF5IYsE2O0rSOfGvfUpxl4IWgtZHPMotACKtpLKUVvs9tjf8h438Rq6O
9dIIYS/1/xV8euIwK6xZj6PA5YON8wfS1pZ0fuqzESWIRO88kUYksyYbpNX+qX4V
0+xFa2KSbiq1R6vQxvXdkNoSQBH8su9ObVByMn/gpuaVOfBG8lsnWuA04aVYuWAV
izRrbdPkolt6u8r8oR+R6thPN+lHD8WR2+wZtuJcxscIfp2AlFgjL2aaCdvpf5Y+
Aoo5J188acBGKSp96twnNHOnz87CYioRaGJj7JJt7D02RiBATFiM7aZdKsl7yRAH
zNv4nqrxBpQB2uzAkcBq3agws6i+BeI2xUcqvRXakv9XMBv3Bzm3GmJqrj6kRqHd
GYKxbP1K/OCaHgmIZqoDE/bim6jhthe/C8cN8fpVN+4XhoqGteM1eQPaHbsGaTKI
J2KvKzJeU1jglaJWcN8NG9fBhmkNjRwA9oCkp7m0bzVR5BdtaBhmJew4j1KdR1vw
pP8DUvyhXhxxgB9kzE8b2NQhcUSFN+82geUwhGNJBNmj7JbGiuZabVeoBtFQ2AIi
c5T7Z2r2caOI5T181ITIiGkSVm4HwyFZvv8CBLoPap7gLw8zzXkmaUe4s4IHlTAZ
klUkHIqMcwpnrTy9ueo8LWmmj31xtVYHVhgQ9XF7FH/asBWT2XOp8NWUt8FI7HbY
18uqP+rXtqKXxqo/s7Gsfa0826tAu132Zi6tCKc9R50ByNLOD2HRY8a7Gh1uaHun
wutznY2gqJbxmuphzyaDVtHE3lZMufazY7DT4Ypy2tQOSPRKsZZQa+x8Fngqs2Mm
MII6Y+ActP5jlHteqTHiUvlFBDM8V8ikPUe/0ofKAlvQPuCoFL6P6XUXCyBDIhKg
SHrqDLfo1t3QrsnuEovqdaCZb2Wxv8MAz1JtrmysBPM+mMBbwfXMoD8YP1k3M2FL
o14GVjFtnhk9oiKZWA38A0gshzH0Fe1+yJkes/YG0uXrXAmI3naytJeHFniA3t2X
p3YDCu+vLXER9rLH9oRdnNxdA3fKJfY2ooVg7RpvWSbNGeD+cijhQtu3KtFlR+kZ
GqPa+yk1SeENnGYIQJAW2CpMzFYLwVpi3eYyo7zPow5/bzUSvkZBPstoiRcMHzGb
zvjfAXKQsyPAUJINjf0yv7W6U9HaWujluzilxqFIGiVWEboAQaWlbiVR3NeUKyGM
YMBXOxaG5i+PF7pFkqTyld3BUxuGv5kIA4xYKdBdpKqzQKkyKtSzLqQYCVC44PN1
DUO+XoWH6ApMXa3BoCr4lldCP6PRCv5XC7yIG5TCeDSH3ln47XcasUCzlKawLorC
SZEh4AEzBMuw2AV0biBOWa3KodLW3UeaC+VqlmeBHC7OmPM6AS1nA9dRfPa0EPM0
aAsxnj++dwKaHBEpnIvml1iFQfZCu9LXTA203hcQ5Dg4BDrJtlv59h9a9A3NeGB7
o/C+4VUbnsbKSNEWYu0f58MNYjQumWm/DJ5I2fERPoBoLXw0RHwpxGqjCkS9fSD+
GwpgT52jRgjt7EEvKjd/gA3LD2HrO6muC7UBXSFicYJTzerd5i9g7poWcW1AZuyV
8Z/CwPYnVilT72bW6KQTb0EjRWQ1l40W1iHDhBT+5DL1+eOWlFgPH8SYs6/DqbEv
zgWa39MoB6RuEPeLvXDexvC8Gts5fJWcl3Em4/7LO/U+CaesmD3VUVq26SjDUkc4
BphjUNMcpFMJSEJmK1NaYSJbx+moW8Hlj7sY8pU3NKeN1bQA23S3Mj8xRrV4+wbE
j2IBq4fZi1P29GMuzEwGLaPL4vnQVS3HSUPaLg3yaSHnB5OA0SPmXyo4fPYbZ0lW
Q1wyeny8CuzMdDSTKXHv4GxXQv4xgF3pZKMPT1SanlVM0O13nEBbqOaC/FeldJVK
z1dAzOj/5YtlCvJ1HPWhXTH2jvSyq7N4uz4VLX4EbSYCsb36zD3TqaiKhT+avgZg
Wc7XzBXNeflAB70lDWiD0K7EwvRxKcZypYnj98yf8Ll9iUyMwn82I7yH7ewsn8A2
dNfBiRur/vk0Pk7mTWbQYNOF1V/fM/96v9ZYi5AUbdELHTJQp4EzmtYTFhzOqswl
sF3gyE3zKI//ky1N1G4QZUDblEXc/FoD/zTdXbWbHb5e0s9Sb2DBbvat7zaNVX4T
As7mr4cpsgYOQLl4BWXrrr2kjv7/RP0e7s/COvmSnHO0hAD5vKODGZf7iON/Wc34
YzVApaCaOGC6NYjCUO9Q/yxec3UClVKxFsDHkLG939HyOXOusfAEs/b7GxVu7src
jY99+4UL/ER3XldnWshprO+/lQIFfP7FOWpICQGwVjHL1/+Jnryl1pqF+jvxfuuI
H93GNCB3GJkdC4+hS5igS01woZTPXkfAoc9Wqu/LiHA9HnsmS8DtmdMLQEqcEzHT
xvo8xtC8Tb2bbtIJG+61YyjJB5Qo2o6foSTeUtZD6f6SQJv6BOKhorVk+epz7aFD
zaJEzg6GbpWLBqAWZR+uY5Q7hl+qWYrJHZCApTxjkM/ElSoJOwNPljxlSi3zgDgJ
M19NwCivxHRk/SQ42ObDZuLBfAA2qRhlq4h0tWh+ImVNsJc0/3z3majYi/tauUEj
FLyA05/cZo2AE7WwapvA+g3vo3uBzZ5XnqU94ifECJpYeAE7E2AKNv574Urtcswp
TgBpn10lAXDTFGmqlLmLKctXNqpRwrLJZf09SwV9ZOtmkkh4xKIYoICwJhnwKuHR
cz1tLh8LMR60a1TWN9DC1AwFw8um2x/+rx5r35Qrz86Jbsps3NgJcoIraIpSfl1+
HGM7d67RpmSGc1YrBBGch1y7rQ5ZLy1obAU+7Yjk67SC/jCt6KTW/WpIP15FuEMN
HljRMrvPMDmLgejBtXevb2OhmGEyKRhxQF83FTaq9oznEURxVwHERSyh4zFbHprG
VU2TxA0UQqndwHGPFYhubHKyROlbvjXUyp3fpPDSQy7ChRKjtsm4wBJEb0arMC+Z
VnQBkv8ct2+nv6JTealIW2h/bmiOhzaDebhttYPP2MRMv2HaB0RFUfvvtPijPeYc
C/aN8wt4AH3flkgloD8l9btSe9TNRSzmWJQkghXt7SuEG2P+mIsYtI+bQhjNqPXn
co1F/MGt7EUimo5MmW2MN8OIQrxTL9vs1vpe+d1UNgXnwP4LY2nqALQ2qqkaYmof
F92l4TTS+v0ZUOu+IZQNYQm3pPm9L54RmLauWdQLHen+LKzyVD4bLhSrMB+Ig+CC
RMRcUvPODt56DK5fHbchIZd0TyFqfzrNSo5FFzVlLFPCs/ZpxEccFyTgmZippmWR
LSJ1S7ZNJDEAaag1NAo4hTuamnlxYhZVauMvB2LSJ6KVoYHFI+epwIypMDFeq/lS
iNRh9zXeCCPz37BIInze2MWwPYofNwLXv3OshdZSYr9YGw11lfqYh6CF/GAIjNU1
SOer12XwjDADG+T0TjexSw845clOn7iTQFzOn1yQt5fi0T+2opvumXv50zs0Sb+b
ljzmSFyjhulHtju9YBqt96Xq8089sknQRenOduCRswHzn9QB5x2fslJjAGsVGB/D
N2z5RV3S/I7jV6AGwguyYOhONek2Wi14JsOjVrCj6vgDNHR0nBuGayA0SvqwROmr
C819LUbCiQT1eK65VRmZ/RvI+yPJYnI2Gx3r+UPCKnhbTjW7JzUPTspXRRucLHfF
xAbVCY6i3dSX5+BMb6mMPrhrWkIIat43FoJoKdxDgD7Ma1dbMqzs2IUrxqLoQwtn
3o1Ct6P+CPpCbFsAwN1OsXI7HuAECAykJlKnG7OqMLiVrLEm/loqbIHWrxWqTwRW
m2NSaT5mBLbt1dux0aEy25gMAyqr1EdMphBUxiGnzzh9CmGdGHqWyAEOIR7SR8jj
Hn0i7BLvw4yROqyHQUvKgL3o5kIaXAfc+2XT/r/ry0rZUQhztEE+Y3TJ2fR+qTOq
B64LBfTtvLv9ZE/YjGQ+6Npr7gzzewhUDj7SMlGqUfK/3a2IH94ZpQrxLPOlgwHv
acxJC2S1s7dmcqOCjjvPJHsVS8fE5VRyhcvcjrBWJAQiFaildlJMKl0ekS5juOYH
F+fYBO5o5HuPn2jtH1Qt/6Bn8aLjOqPj45mDLAREBHtnniIA5pPxnIsgu/+uFGwo
665MYF+4mZ5jWZcjUk2v4aMKEw1qwZt0ayLM4rtDAR0Keo9yNyAvsMEq085Trehh
4DbK7w5O7JEDF3+ZQHvrCrJ01yMDvINjctrz8Pfvzy8HhU0aXNfAmYCpg41wC4xh
EDTOwrNLfGYlSZxjO0VOv6CgKyHhFI4XCn2h6ehE6Sa279JIiRG/0O+MurVE1gLj
ndnTGzToqEmdnWVHIlIO9S1GzBrPM3fFJOvVTuqwvqWFWTyGG+9B3zgSdx9TLxa6
AWoTRaZ53CMiyDeREq2BHDi024E17aEj9ZrjA+VG5f/P8ykqnONqA3XJLQbrEl+z
1tsvmAFcOTUxUnkqHwjV3E6SaBeQB9qX9v/rRc+KijORsSUp0k68mA8AtmEH3u62
MRbvdXCRdV0irM+pg5B85SUWBn5pLB0UXio835A/SGEa50yeaPsGTNFy3LjrjgqO
yoCxiWyBo8v5fqD6cTDvveDKHi6t275KmWC83aEdopdwXUR46OaaMmWqwLgZLtKc
XZtUaTVMTHV0rPmOXUtjKldLKGcFL/u+mD07LGXTAX6LiwXti6rjhoFN8uW8fED3
n2GPQf0J74qTBHnAwvoum5D+uhC/35M1KuXDQ6z9awW8a+XkPzoHP992YufytCcl
X5eQOLlGTduGXyF+s3SeLdBcVVYvpRHSQacTwA9DprYgLfyHJToMxuEpK3QOfct9
jsaUz3LbbLDZWn/K23tFJiHly7N/Zr6QIgg+adCegLG4oYvHaDn3luRZhJXKpoKM
dLPCraCSEAQ58pF7suuwMb59Ku/xAYcWUUpAtKlgU6LhMEHpXUKz5/PI2GE6et/n
Na0Y7pwVqFNcEx+jW9JgqNzKjNHgNW4il3trgZthhq4LO6gs2Z+pADPu90tT0ngt
46NSHCgds2YdM+wlppSXfdJoFbnRp7SArvpZt2V6FM1ryyu5T2h0LXOXztGhO8rJ
eYd5IBsGS8cPL5QNG1j6QTKnF+eZjNLZkv50NrUCY2pQLzFT9cMwOcF+HPzU50eH
XHST1yOHCkYBCPOOBtWIvEZeGgXc0tV101mVKVhrr++3FO59mFr/5tbFhofK/gbD
N2smPp+Q0y4JjRs14agKWsWrTcpzImxZ+/YXaRzaISqpmtSjIJ4Ny2bbt+6b2Ona
IqyYCMOfOid88V7u3Bxk/suvTyoQx8VBZMC8DWivkvry6FwCPwW/bvOdK31yi8AN
pC4bXtJ0T78vmKo5cuhYbmNMQ27T8Pn+CbK8HOimYfNMVcmjtudfK48rKVax7vsX
HsengIeSNK6zVPOjDmjG14fd9XDoLo1+Db+2xBsGxy+CXIxmegWCmes393CXPkAK
ZAHRC+9DXS6/FTJs5BTTQXVjFp1B1mq0nUzncYl0AOUDyHIatfaqBdRDvammak4x
WG42S4vx5Ij8/hWi1ZSMiUbhVP8yN3zrdK7tSNizbf6ORku8kkbubp8Ub1a6+rnc
uEPA/s+trzBQKqskQZhj4qt8sSGO3SfLHupD5yaFIKp3FWK4rqZKODbJ2WJ8NUJE
NqWsWjFb+vAYjyJRnn8btMHKK0UQNZy1PKBAj4UNHNybpEle3Wb4f7Gc0HCKLylP
AgsAzuPNjr/0LOvIi3qzUrIa7bJ42VI2yVEWFrzgP3wiGjLjp8xW2WSr+6AmWno9
pjjOASDk+tHKyX+K9psEWZ0N+ML5twNNbycZ37xsNhPG8xT4Rf3u9Hi4jS82oUq5
t63wSm/3mSguUuntjLhNyUi+JeeUCWEBmo31wTrAuXE1UWTWt4+R7wC+gnFr0zOD
57pnFDHV3orsvUOsc9B67Pas7SpQK6PM/IylbuKM94MfvyXQVxSYYfCVmJjS0NxC
uQmgPSCJVcbJajuQ8rA2E+FRoRRLCPkTSyYtmGZbpdeFvEmKhz1ltnDwiXI/bY9i
skcJVbLGUezt0IGo40047o451wASq0LWNU9qHc8Vo5FhZX1J896P/RbY2Orme2t+
EJSvpn1rAlbIM13v4n65S066ctrfEv1m4R6L6az/YIG8bDw96eDjgz4v1+0cuogs
AyD4Fw5v7CUHdn5ZHCODU1ndnOA5QRniIa8Sk7OH6O7Zym+nZBU6ug/oiUBmcWfp
7A9EbZthfYaHJEVbz+LX1vIIvPguWUy+m1PXq4VrQyHPLC91Z9bro1d9MBTSoUtQ
9Jsl07niM/neu2ytfl7TEvowNTL+2Cz7Sx6GqVv92x34m9KUoDcBqdTuWV0gXU/b
3TJDBHHK35rDF0qIe/2/la8K62m7Rot4cl1d0DdOtpk5th/SLajuU0woTgkydVG1
Zd3W4Q1Qky6cm6P+nHZG1T0A2C+7QZVYrSLHSrLGC1CDnUrs6Pk5uH6AObkM2cc9
H8Wsy7m9CsoAChUCw5TgKAW3JW85lqWHeAHl67O1Ni8jj0vjWzH40ZznggE1ddfC
Qb8lC7L8uqwizH8QO67h/oauXT7uaE4yCGjR/YexMWHbnSGtDSfmA4BbtwB5CzSX
fLlzDaH1gnris7w9rOigBhmzL4knG5kRM091PJGr42ggTlexdVK3KEs/krHnCM/k
KRwn0ebR+1N7TqFBQ1WaKVOawpTwLFsywkmNrfLkO1f1Djlrr4FAPhFoO0pWuN45
uKEdc95U9FH1AU+eiilg7Nm3TyMRCNRlrL2osMpZOzVGOVlwaREuqJfUGNC6N5hJ
MaY2hJsHwoa+kccAVm4/94hPGiibdWpeUc4gLdGL8kpLtubqB+hBP7mdiiEfdc/f
9nT6ierSAa8lWm/kEm1UV7pc8ZkNMdV6L/5nFqNbynPjiC9VYhsSOVLhMxzPMKRd
kRUvTMybqEYSPCmOfmLrdCVvvkc4HNVVU71ZZpYin2oYJ18jfVnVXqEXPaKR0kbG
vrJymsZWxKDXtGDGW4VKzG/3PbUFGr4Lt1DhsAhwBtUJ3KZ32heOigfo9do94FAI
KeMg0WfL0OOhnW8ru9fD1rUu1F6f1Lp4rhvKBlhUKo1jdDi/NPt+h5TqIg7+5qZE
j4SYQxgXI64+VoYx/MvWycS2PDgu4BYFbTK+me28k1vrT2cDtZVVqjSdD0wHfCbP
TRcvWagdlo8LgwnnQm90cLkvs4O8Pj4CH6UfvYIdxhAzgmEspcjbu4XrA+/BCqvx
I8+gZe4Le/JqNG94IATQJ/vztIJ/t21teQPAKIRu/rMQVRmiZntSBUzm20qWBh1Z
nCSv7yPc61bEaQUyp1ChiBEqRDtISLFm+tcjFoulWUg+OHV6j6Kl78y4XpD/Su0a
v/c/oz0q3BbLWrAQWyQQlJ947JMXdjy3mH4ta6gCC4raqBUiJpNlRHWm3tWL1nuD
QJGJL78eLWEjrPAMmt94OQSg1i56NMAlzFlNtIcuhskPcUPDeQ0IC899yyhCJXc+
LSpRLyju10SCrLSNZLUfhl9l2dTcu0SFEiWExleytQhSZCxXTiOyrMtB44iinPVp
5ZCwwXnIIbgOt2l1o6AzwqJ2UIm3MFqheAdItHUL6ZzfV4nVe5vZUayqbwv5QaEv
iYTLbHUzrWQcRDcYA2RSaJ/QIRfQBIMuobyIjrO/ubHHaagY3ejBgDb29L076Sec
6gTSuaJvQE8AzJV+VzUm2fsNRmB2JPbnMpOrarplhTsYoo5g6+feO5Y1lqp2KwSu
bw/BHPygHSF0aweDD/rK3vo55rDnA3PrNDQFn6EaQyf4VMDweJIhTFBZghFqTS2w
+Rgw+R+vgKvTzJTulq/ckEGZUwjjIgGZgbKqj14Lt6WK8Dj7sccKBr61b3zukbqN
TGLJ50ELcQz9BeZAPYaV8RWT/uGYE7++S5IHxdBUkIJnsSxWPzb+epQhQIBwBVkC
y5FNQXioiZpMGgxHj3nmyiljqjqbbh2R/N114t4C326aUFWyRwBeQKJX3phkJ04f
+4W3YxhV1E0ddYkdiTkqQfHbp20p+BvHFOQNyF9XPoumtiakpTUfgJP86+G9tyYw
xf6XSDioVKXKNR+tvCfAdThCL9eL/WQBwHG58bBZz4bXsTuntSATalvsZRLIpVe8
irvw84qJkXz1dBcC2avC/C6q9mjoAM+iSyCFLaITCGtULimT+9tr2bE1uGSK5J1X
QVO7Ht/o/o40CgUmiVR9JMgNB9xrqAdRxx7iXeYxjmYdHJuVyiw3Dhc/fWaC0zF7
f0daYLRvMZWhdwwxfR+ee1FbiNqRUTyhd27K2AZkdgGxLWsycIVsGtpnoflxkNpB
bjDVJE7t8EGk44TNV3qsIRVydG4YN9y7hwVHCcYSnPVtjVFg327i+V0Xy4A1u/eI
EvfH2SA23RInsJVgDB+SfpTrDsIeiCh4FEVCfOYqMOLEYL+hVtZIKa4WrZDbioeT
aQgGgcWYq8TylBQiP+8nZLg04Fenp+dvM7TdqEWk1EQ27gjgTPjRaZ9upMdVK+/X
bkGHOUaJNDykBxM/EwZRUXaKUTcws999O58nrPYSaV7BxTfHBskcoh+ICvKpvdkL
1FpxqR/ZR5qYH1qwxM9Kv84Ks/QWBocjVDP/6/TscDvaOHEmQKsxJrURo1+GprXL
FlR/nXhcxVXyGzML8ooYMRh8aVSypnYPL30GbxQtmU0gmxzJXEPuxTk/Mu8vH1Cp
VpXQZCKFgMpjHzd3zdRMonBOopjyx74GkojhpmA7+DwxC3pJezdCuSPt4yEOQvMA
ipSBpiC+KdTXlp64B+6jnwV+MahtDU46D/aVa5/mGB84tj2ruWXpoUaY1u3sPs/r
97Qjx8q/1TUG+1iZuSywa7G/bL2GCnGE07zZSDBvJj1YB0ndtKrb76q9pY26xiun
fxQy90AGZEN70l5L2u7eodBmG0aiZo+Qifz8yHUVsJd1DBsASrme0/rwcqq+1/Rw
hCtZFVe8jKbZVmW3z8VjS3z1QhfS0aJdAaLQZMG3Y4NkJNiIvDkvqygi7xlLWky6
ElGg3nocz61xT3BGQ+ewk5oNjqBHzAFT4nCwN1ts70rmwM70efgvQ9YR4JaAqXuJ
bLm9D6buAa5HnCY43fCI/kOzDAOFpXyHVDjq9J1A5jbBhzcWc4A8Lr6EGWie+X7c
IRaUZjlCOi0WRddVpmLIfPQFcxU8RfElkExF+4Dm6iz0C/AX1JEIev26EUNvYXaC
2vaJRvircCUJNTndnKjPwtk576r4GZzKTpjfNAEfkNI=
`protect END_PROTECTED
