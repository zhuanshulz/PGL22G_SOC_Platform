`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tDZ29FQKpEmgYQWGLq5Iq2cVp7R2YUulFs/qyIqM+lqo+0senw2Suek834DIbhzg
zpLuo8k2wjVl2uBgqkcwyScyYX6Xy/igFnZyIndP8or6TxZe6tt0AVXnlGv3OBJH
rLVd9Qx+I45tX+Gcx8L1G8BO2hvD++GVz+ckAma7ipiET4fvX6x77isut/pzVBE1
74Rdo3wP7WuzxVXcXZsfEJIKcMLpQyBmDgLXh2937N9R2DjPZv68xX0j+AWMR/75
81VWzBn9Jb+2ENh4h8ARcJ1DuGiA91f2xaNCWZ5Pb4wY/JYWTuto7w/yRMLJr388
fK9+Rx9G7VkasR2B7fHNdafFv1h+/3KbK285qp7zSH4n2p97S5jKxguSTDg+NK26
oabiuiiNTbt+IC89tvKI395+AI1GKR411uDEikSK8ktQkwkXXFj5nPEX+2xJsYkO
zPqKil1L1pnowyV8ScUNyqRjAAAnm6EyjDjESkWRXxm/DoP1FKsIfAs4BtFabfo5
w6xl3m6nw39yyMpb/i6+fg==
`protect END_PROTECTED
