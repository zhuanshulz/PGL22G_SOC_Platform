`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1BfhyKxjObELQj857KW3HOH6UTYO/uPGHxnYA0PD8MjcjEO8zvRRW2BmoSQ7Gat
PixSGbRZ7p6QFQzxbX/PqWBJMjARgILqvK5b3nUOX/B30sTZoZE6+PRAex24NA6y
mJgW4nX3QR5h7G7VipaGFnxDWvHoD82lgS+4u1jRVLDURz9RK/MkaRiIBJ8y6w/q
4S1gq0P3y2NcI0ExtUpg9n4dNANEI9DKdccygfP+lCSs8zV23ycXNryc/cA5yALK
ebdXRFd2xrxwRyY76imsHg==
`protect END_PROTECTED
