`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5hzjINEHIO3AQJWSTK+l+sKPPr3Gf0tkkGddFoCIzRA0J2i1eD5EoB5AWLGpAHdU
vmS3IujaC/vddrxApYHXfXwC1cH+boopCr/EGX+ra+U2a2lIUwv+ttjbNOtc+Qc0
Ax62eXmZXX/yrcN4Y8UWNHQx3NViZ3/1muOqD/bcMRzn/NAucl9pNl5IsfjW9Rjn
Xs7TL74vcHfg+1nAa29IS+VcbqNyWSIDvQnnlS+IpuO5+5K2dHOGlQluexBQ5wn0
inZaOeeMc857/I+HJa7FkUWBcYzOoKiizhZeNU9pJPYYafuFII47x46fJ6Ed7FVI
B9Xo7clozAMWBnhT237Axd6GpS8odkMoR2xkS1Ri+hTxY2p0J2iYChYD9N8j9jh3
F5K5991fiRfLMf6S+/TFww==
`protect END_PROTECTED
