`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p2mD/DW4eDNYVa3lPGhiIwWQ9jwKyrFYbdCH2naY81Z9997q5CId7ys6wWon1AMS
z6H97SLsHtuuhriwRvhmbI4r41xgdCdCvkNjwLdy5elTeRf5clTz6WDO9TO+38NZ
/39cG2mjj2ieiZyMiWr7sft6XI/uR/5sqgTEHAIfVPBbT9So1b3nkfgQCSG+EUfP
TvMGVMOdVJFrRHFh7fRJ1eYmTjkZcW/60FLZEGjI3ijKPWkYswRvtek9HA2WvV6Q
9HESMUavEI83GTTkHEVOzuhqx6dP1tMVWjF/4L1XmwOcUW+MaJs5s0fb1w5G5tdz
QxH5I8bpPpV3C5Dk7roAs/lODHP7xNo7tuh1+kPwH3KUMPWseBn8vu8zL/D2RTCk
xxZEelMkj8Zxi9K2mdDib4QeTyUA/DUuYZBHfpkS3oSc/2TWPgcukX39w1fcaRQj
wDA3JklJ8ZFPbuj3DYfERG0owdmD07MRzEtfeem9LCEoZK5Nx0XL+1eGUYbo9CYr
Zc8iNi2YJJ8S59Q57AsiSVGyJRIJAdEujmDl77yXbTOzwq6zaY9KipBA3IxaX3js
wlEyuVcTYLOGT0REuKI+P2z5qirhixRSVzsiZnhUvK4maS1PujlEARSqhBIO8Oc2
i7zvzXIGxJvTau9WRgZsVEY46H7bZM9QLEHf+9YAin+ksYsy2iEl/0R0Ck7ulHRF
CgJm9aYvxf9WoLqEG18a8r6jnhiiEljeBtbOdlUVMlWN62G2ICE7f6zs01OSW0zq
ADse3tgCeL7GiBN9OKJIb7ZpqQcw8DBgdTBeOksuxXzlSsS+fvj/QmcyLw5Ql6aL
EH2803u5y8IWRT73Okn0RjVHw7lajG0egg/vk4/BdTvJ3AsXa/8YvXKhz4rsPJzW
5VsKhvuo1VwZPUmOBRCutr5uo/kdluyoNjsAckOT6dtFKZt+YnSpf2gV5tpMRQMv
gUasiTlbGwtgLmndloZFyee8Mv1Wo+1a+cGuBzdcV+yXyColYmvSKAawMMa36JKO
9D1/tau/NR/Js1lNiEL3yiMlpyznKsFvd4BgAGQS8WvKm+gffmAWItO5RTqB69jV
+bHPLGEyMuNyCPP3JkczDpAPsResjapJomYYVcrocT7VXnkdGaoOKiLkQRgurecl
vZbjzdtcUG0Mb+t1EUz+fJB4bmIg5Zu0t6wT3Uh40twHTJ4MyG9ggjv1Whi9HWLD
GekFpc5vSYOSsQoxDHUjMrhQ++NlNh9ahk/M9mA26pOEZlC3l6iwEFtTAgX9CwTD
pFeyobkJyG640uC1vtM2uyyZJrRujGIMX8E1a8wwP4Tq9g1k/VrFqKGehvlMZsSh
7FMQvYoI1wAeD3zskNCmwudeUXA64OgwfcaDHK/9zm0WCIrdzPidvCxqaUoHKrYr
BnbWa7k/WLF8tCJnnKHqjo/wAGf0xeicHC4gWna8h0HzMddkKAwMvNAajcKw3tX3
`protect END_PROTECTED
