`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElKjsmCyj77y7jEcJFd1sgPeRHnUJORKHpDF+7Fv0gjaB5iGpw0/95hQ/85OKq6N
6DjGOI0YxFRCzcz6Z1w/fYiTyyVpMWBL1NmJnMgxVrt7yvp5uOjZJ3mBQWTNLKWN
JyKcCjCvEcQZwL/CxS+EyPSyXbGH9V+cJ13xR/4TEM3RqrncD3kUxnHgB9nWliGO
XKRgLBBCXVm/Lad4laqkUEUG0aExhyjhS1XDyD7yL1UX4pMhSCvHkU5GfkNKk3FG
0WA7XIVRJt1Ut3S/V8t54QA0WPi/PfK45pW30hwh85NzNwXf78pessUttIk0ZOqN
2xPWn1GYlPrw3MIz9sBpR5/2OmCsIB7KolFbxVEhaLkmkxUa4Ao2hRzqTKKh0APd
0IrQiih5cP6wYZKrYHrQrgYq/xrKHJaqLyxGLBIsKtupNbh6zO2Sr5NHA5wfE2S7
25avtZm6JVVv3E6VmV5CWPzr8uwhidMbaDPW82MSFttYcf+wR3Kb6svMEbFx1zoA
3Yv5GPC347w1DPo/LkO1o26cjjOgThUsPrmgROhR5uKbrNeXpspQM+/tqN86mO0I
DPb/EEdfDR3d6xTceYQ8TVzxBoa1gTZ5OVfYwcGARnbORojxppD+svQ5qVivqLRS
EH6aR2H2hq2Qyt+wjmL5KYQHJirxacEG6mttZzAcLvdETkcNymhKNyohBG+NS+uo
ORJGtFQQuMR1d+6FH0nQrzWL4c6xwoF3AuYDxrqGu+t9Xt/x5e8APOTRtuXPzMyh
cJCi9ppw+jQG0EPTZ9EZlJiruPZbZcQc11dCiJ4+2DtdUb6JPLDhf2+b2Mejq0Gy
4RSg6XxZbELgNznKrgnQNmnMzCiUSJ/bhpvi6xI17NNcgQeZLjVNm6DH/OggT9CB
JZnlNeNz6NbuDsScdHd7UQzzYW3+ZwAuGkeBd5/Gxef5LKiKftXsA181j9oNojqk
utuhFGbcjjrkQxGtvg2faMLOjwcY22NqU9QiQqvfirCvtxSr8Yh63ukoG89x2qU4
miutMd82am30Pl1CSjkB6fIx/OLYL6bdbcg9KoEtmGafzdW85fVs9HKUcZ6IQxjw
0yuVu7z4SIM4Ptg9MO2lStL1y25FN3yimgA4XgQqP/sa2RlI7ktZmSBUgmZ2Rkyo
2bicZjBSlyetyhdrsrt+tPtCZD3ShlCr1jq/dg+wE55NyC0ZCGgS7kamThBowr5s
bEMPrDafaNvTnT2fHkQkKufo4iKFodXkSru26seqjFFXYxHIdWWqSoEcC4DBz/k0
Z6T6w7zvebWnd7smV1UdKUfHbu/SUr1in3u9QHUyLRUO1ZFihhm84G3mEKLb7cy0
HcHw7llAyHsq/d9zLStUVt6qu7FxfnNhM1DtHCIl4f4EDdcTOaBMh5n9UmU1ZfRo
mfN4XAkPX2ET5fHe/xChkaHkNe9ztM9jMYz8XDsRmzEIm6354/QPk2TsgJajJLFC
FiMXvbFFCHpa3MStolDxVF7c74k8WD85n5K1D85WvbWkD3TX1KqSZd/vAFYhS2LY
XQxjJ5VZuIT//LsL9WllVPXB1iJ+NNMr1VIFt+lRD+wt3n69xKiH7Ye2x7NcYfQA
c2ns0PruN5AKmcxFrv0aDzKwO283vSXDRsZ3RpZuL9qUtGRMs2d77wPTYxWl/L6f
70fDO8+1wmmOMRLrPcg/kh02/i2A3Q0pDtm7Wqfy+Wc8ZkAfyglecG2K+dP/Rhpw
WXxsyyLYzLAjbOzCRqHHp3n22r52mQe1SoI5mXzWrlnFzVur+F5t+dqEXQNgEDfb
fNV2ar+fnT5T0L62ZkAEvO/JSWxS9FFLhhQpTg7MfTgIQqmMTYJnfK9MT3eO5dGB
`protect END_PROTECTED
