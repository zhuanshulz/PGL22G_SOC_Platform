`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xa81b+62CBtSDK18yrArj2n4dGhAp3312mzSHvZjteYEC03UB3u27NE+Yawba9ju
wl/BmSpGfPhYVSbjKOHLbAshhGn4NSfrox4ayP+8O7fBcl9rrfxoegwDnsF7urCM
iydPKyCCgWt7Q41MTr94xGmEcYhJahvv8i/CwEG/YSdvkojtFBS96yTIOgKJc/OU
cBnrcAnetn8wzetelsBcTbUXWAyqVP56XYnD+J3x/fcFyx/WMvIkTcYoL5zzCgF9
1sLq6qK4wMLRlV4AWz+NePM+L5xzCkq+LjHoz/KXnwEyXly1P4xiuppwf+W974T7
9DwnhHjcR7XjzxikHZQYYwWQqo9EPe8VXuPxLoG2JnXvZd1Ly8i6ZuVxVyW+WOac
`protect END_PROTECTED
