`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWw5ZK5f5eKcmWD/RqzCE8xpIPTQ10pbMMOf5L0erWbhhf1wwmhceKbZzghBuQq8
RBAM/onvCwqpOzCSd1E6LLP8nJAgQ5QhnlSUonNdLEBtZcrO4Z/0M7iYSGtNSw/i
V4/AGt9ZjUOwSg5nGO5Mp7qYeIa7L10V+UQ1lfEj4+b6gaHYjzL9XYbfKo93lnAy
EXDFgFl8nWkNrP22Ef6ahLKnlUPb4X17JmGjSPabIroZiNHutrii4NEs8JsCW6lX
52/a8HJMrm63DANA1Vu53Tzi1PLRLOo9kZ40c2xSCWzvJnegNKBiddcOptwSOgWY
3lfrrtQHEmyIy79Ijy51JRud8IpMulNT4lpqGvLBCIlgB6LNIbEv6ywc+7Y4WUWL
wqdZghOxZ3muiVUooZNK4B7z/aEFUuBC4QGkL3GVzMop4+Vc7rNAJRFZphFY/eF6
TDU5ADAXlrd0GNk9BXI7oe6RDDXRRYea+kRncPEQh2dPD8XHfPAIecvekbXmZJ42
9mBuDwhObxfkX1TqktX38vK09L4uxJ7QdNj1tsM/uduggezisoO5+wnuew1JHRp1
1m5dn+OhW9Pv3yYtlAJDAZXMSCbwyluE4RoSl/s7B3gv8byuZBwMbPgTs2hYWC9o
pL/BqnneMuVqLImiDJewMhIhSf9ZVBtl7GC5jRNLl3p3wmcCncBrUUISC97iMAbk
C+f0ZgUJgXu7C9oYCuPYnToXqiyrp38w1Sghdx0DUIi3W+sd37WFQWNHMpSBGZA2
oK0gWVHq6V8DJ5ba+gjKcjmKs2dg4joQGXzfdtVfH3GAubx8cYpt29l0F/gffyYi
7Kv8za1FTqPAoPuZ2Y/b6IoeGRh/C687qVqUmxpC/usVrSWXg6jRCndJQiRTe6h7
PdfOtB3vErlT7q4akPiX1W4Ua30/51kmIyMB70ejOmBOkPno8n8xXYjdz4FoWd9h
DjU28zJMzT8fCCtzgYMuD4R3idICU8ENmGJusuX9nEHfwDmvivRJ+fhOmxZIRtr1
62a6U9y46LUD4atf1Zjrzi/SdasBierBw2QNvRmFdZqKbcDoKRdhZiQQ/j3AMR47
X1BzUfkdyxF/M2fU9auhSS0VYf5pqN/T+zmGwlcmkbonWpniiScCtznvFtNpvbsX
W2kAPuOQVSQXnHlUbJjs+u/mH2lFqpaq/Zr/C40sYfY8kcxSDF5v9Lhyhdtq3xNx
zTHyXQ5aeD0FBFQJzwZ1xJqvgbhvjBMQXX+XvdjYpLo+F4jiSKgWPxtmU82DU0QL
NwedY0Hv9GDXzFv8zJV3Cp7CYMVUBOcO9MvnDNwfc1pmST6zl8hf/LyKrVmOzqGZ
MNNA1rbpQNrnb66pyodlxYcCIRyLs5sUd4ifPys2BfA7/RnpCG8cFfqwEwNEZqZD
TNcCnOrfjRSX2Dt+NkYjqkBI1VEEhHLb4pg9FuS3yn1dtTImBlyrmSSzTWF0E8jh
BBMrOQU7RgflnU+0xlhQL/E3XD0lzmHiWReQxnuwova7v5VhNmL7Wu8fMwjXxiux
C4tPS/uqjJ9sPIis/ki4j0jT3/mnI9AbpyyJmYVqQ9pnGiEZIIy/E5gryP4+39/S
mM6dBtatnUUAJypHPp2lIcgTqlvNGwYIHgK1AFUJaaQdpZYgrEGAZgqf5LJnZBWz
uH5hxXVSr1aNr7Y8KXZdX1r2ro4jK99+9Pk9OLuemXeEwlJR0GleZhaJbCHjMfJG
cgyASBz3RUl5Ez+XsE6tYc5ymEXoEp1wJ+FYJoHxeI717t64koPqePi2O6BZNF1h
lanObpax1XxSGnG+ZuOgczAF+661sW6GwUqz3sSCmFWR/JIDSg/NigQEeJOSiz9M
`protect END_PROTECTED
