`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZC8pX2UPrRnbKYgxF3h40jUG0pUFOEO/N3y/w8hTabHrlysBM1BLK/yiVk+NJtJ
BQ7b+o1Ua3QYGMnCWP0zrX8B0Wu9Xw3fG/1GowgQk2G+uRiGVjGRXPmztAzjXmIW
pA+VP+IMlXQIvFhb6LBiAQSCUho5j4WC75c+BnLhXBSmvEvs0Qn4uGMd4UOte+Ci
I/JNfyvKc6k12l67BB72AofP80F2oM5MVLAowWnIhCJe1WupCGacuvCpX/sEhsUw
slz3xucNK+mRqJGZtJmivVK/gDF2+/aQGn8gFl3ODbkI4f0oAiUdvxhZw2oswgZz
CttOXlWXE/x4OKB+FOraoHBX2/16p8XSmNNPeIovZ1gfi0hynPQrX/KqCqcjypcq
aJaD3wjWS8bu9u/o/PKpJwB74rfZXuHSCRME7HPOI0rR8ntHOFeJ7jPZRQJxUUzV
pCE0nslbsOWVIaKcPTvyNps1NhaO302e36fcQm4kqDDzr+XLzd1t/xTeK00+tF90
71qh3jD87SiOZE73kfSGCKD705IR36apLpIp62g2jho=
`protect END_PROTECTED
