`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrgaRAqDUECJspIa8StxyFU0ilxWuj9OHu+EVyIDNcdrZPyNj4PfkEr/fDnua7sg
5f8Q4NPgJaXxaF96cQ7ApifVKXKGVN9Z0A5Q+DO8OKsqrJ+lPS3RLDqnRmE5dG1V
hEDkS+hP4e+cyqfXRHtBQ9PNCGpLSvnkSCt8MPm+Cmd7V35AU24H1weF4TKrmHqx
3ADvnSK0bu7Yrk5HzM7yOPefs3hV8rDzED0M1s+kWsGSmmg/RyGSh8vS7orz2xee
1tCOzCAZ9qrGze0rIgzHtuz/J8EMYKf/xnOakkb4slPl1g/yW6UyVtwePJLGROMh
FtbJMC80F228AfA3zs30kr6hTETW4l/NfmSAiUZ+BbztOx+uLIXxTL6j4b31Zy/m
JY5rgAcTKp8tX/7zP6eLE9/qn8oH/BMNNUGBtBhl+jXZ1g//oJXi+vN/NlJ29/yH
E0FLkNWKFClpSD/UHvkGf3lKM+9iFtWUuNZQioZEUzH1CpnltgB9C1jnf/fNYIe5
eSIpfEJxNrF7iuQlBFw4/BQ1Uf8Pe8RA4Drxfy3K/XXYcnuKhLyDXfwj9BSXZXoe
SaVbrfwHZFifwNjNJ7XJu6MEaFy6nkh6D+5lYxegVxUlhEz/Xc4A1vpViFjzkX3W
bkv7bC+aVNIz3hrZunimp1z4oaq8BduoEZTxXeXAJ8AotoruBquQQ+CqzIuRst6G
8U4c4LmB8HNmCWRqY5VtVqZ5od/td5PpnFDUDAPgGbixelWqHmk3YuTwHqPQ1v4K
AeZ/LOBf2noDe5mELUiqU8NXV5OyMrel4isMw8dziqwAejnrx8+J+fbOKGMAKi8g
luWpepYXY6/838Lm278cxwGwhW+FH+P2cjgehW05J+Fj751Nw4bYgqOlPeCDk4/G
Z9CInbcGTGD3//v3Z/DzRahFyuCArjE55g0YE6s2CZlbuC3WeHez5Xk60dJnCt9Z
ypL0L1r0hWN90FT7e6FscOwJhRoKS/FIEoX0h1szzOU+JokQ4KZVIgKHw2pGRjti
wV2JH4nw7ib615wbmQI3yEzKieQWHB5u031kcc4SyAq43JeYhfkwCDGjFYBL9bHE
YME6q8NfrbRRJxChOKtcNnmRT93G8UViHO5zSBilt1ruy3PAWkYWENfk//vviBdu
iMYEqBNI0Ngcyz+gekbwq6lrWwvFU5Bn29SvIGhEuXYWfUKfg1OdR3OQL4Bp72N0
lQVVySNA6uY/8wwBdI+ucOcpT+LLVVp9b3jsksb2uKsvJSgp94L62PvVb9JFRiNN
pG7+FZB1EOs6spiOdTAwJLbAwFm3hGgpyq44uq2LZXTyCJhAt1OeRp9EpkQyowVE
9yPwETyaLz4r7K95+rVkS2E/RfGhTLs7VYVBgNhUSZYZF28OiCl2PAOAH+KyXxY1
vqfWM3AQ6H+fMFb6fcVrGDfIiP2qk6Y9ZjxqLQrCkeVnRUE9I6zITf08jcmzlNkC
BQ6GjNQAOlH1zAZ2wb5GtHMs5azY1ocWETcL3w8cOqqBfMBPckT3mhGos0Sf8POu
XMQINffeAMdIKrbZsqSdngRjhOCH7XHrd7hoUOaZnh8R+WHWaStkFTgKh5oKi2Us
OanxrXQ58J0kusi8EBSSqgESupC0l61R1t/zi8RgBHrtonunq1plzCX5Xxy7o5/O
`protect END_PROTECTED
