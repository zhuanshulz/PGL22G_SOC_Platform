`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
28NuDnJj+TV2uDmVnZvS+IZa4h+R/yhbSet477BiBwwScT7T2v0W201Wdqe8NiB4
H1gi1RovEPtcUGXnzJvOqKeVY3NELVq75UD0iRypNb/ggYPtBn+byxLByZ/CdUoW
Z7Eyv0tKrrdnjy3v/wGA07whAt/sCUSLJddrufkxyARloJYXK3tP2qnmez5ncc61
PP8egikNCyCeowWzReCLKrjMQg1aWC2NXqzkHas0+PsCauB1gZejK9ZVrOIYyVSs
eoafzHMsl3WAFELq82gUOjPp40QkCIy0pav7hosXwjC+PcPumAx7IPSsfF2dCxMt
wRcZvKRebK0V3WYbu1XlcK2JvRmLt3w0VGH5LDreMDU7Sok3pq/9VnLDCKJvA+bp
I9PRf8NSnB00KstfwLBN7M+i32ohtvsgNZZMVEz3aV4=
`protect END_PROTECTED
