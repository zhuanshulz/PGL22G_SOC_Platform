`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
srHUFOFwRbzpdmow23P8yi0W8yfp8T0yJfMpFJKP8+49lRKKTOcFQmhxdwCPKd5P
6AfzvMHvmkjDjYovb3oo0fuyoSUphBRBr0mThWBBv7SVT4A5oA0f7zXZUQj5ukCi
eEKfd6Fdi0mlAIUCfq16cjf6pdtwDidMG+do14X7WlCINsvdgURRqtydJpe8iCNv
Wh6NntFr27GMaOSMcoOhN1ekhmhZMdvcJ+vchVFqHW1y2lYSHs0GGI6Bj0MClr7Q
4x5yDUuKSxepbYtrSw7/Pse4Txg2U3QxB5MtDxQtONF433AFi7rlKYCZ0qSRF6MF
JdXkyglMwxN51xwJ7q6GKoQVRbnljQm1dL03rUsRDMYDlX366DXuH99krI6WWNep
J8tY2p14INWIyd2orxMO4HNNdCBnQx5k0ym5K7zDQ677Bbgwm+j4+d1TZ/WKzfY+
RurB6gh83+liRQswmGvZolLzJge4Cf8Q5oUaJKokG+kEKYSSBNcOWbt0PaAKYxn/
v1nvRO/bbX/Pj/j67nDZwGAYW2FPZ/q2LRRYKalv9yHBsb8SMkyvRJe6bZEymbvw
oMYNBHDlTm4pzXIF4otgxXKJtUOFqsHaP44lKNGBDL5g54fgVWk6ErqZNYLMIZQe
fd8Hp7Pye1IexhVjAE38H5juNz2qUdZIPNozh4rW2Oky9z+eybpFnFK0GoI/h2i7
lmvG+mq3Xzk3Kq8j6AFtS5MNFIpOOi4dJ/p2ue1CruTsdm7CLwjYtXu/2LMo+TFR
azcIHkWKVlo0wCnkJK0IoRt0bUbY+lqmb/MhN8NXQjf6WNh2+JHsFEf+U9TTPi8k
K0gIQk5VBdtvY7tnA5s56kHDDKdpiyTrxJQ4aNRG2faHgnzh11umLtbBGFFIgAIz
NfdiQYJcbK/uxBEpcV907zFaqFEuZx0prSfCqWnp7te0zMOkUqgFdMT50kPwYJU1
Rt1YQ1w8Tu4oIA8q2Cta9LFNWn5J0b1mtn9slSTecS0QOziBpkAcp66g9KlNz1JR
vN6JK/WYHLUPkbL4kVw77JwyHHA1HwV2hYdnJihwN2htShvPfx1sCIlCJ+15esTY
+RWo9wmpbwC7EzUoxwvJArCb09dVad9OrDOiOCjL2ERoAAGJIr/DoCxZ6T3RWRQ3
gklKSRMrbIGPWJ+ZDGH2bg8VixBjRB2W+ucFpDrrcNajAAR8BTA/DS+0yxAtkEmX
AcKOsRjbemtVMbqWQFu9bcoEWdwcUBddk3G3m6zx7HzXh4+bMCZq6I8PMa6aGhHK
Rj6V+SLbYKECXQR5p4tHFxQbEvDRm4Xa3MV8rvKdj2xnmUHh1o/Tg9hgXTzNjOTx
wx6bhY57AZQwnDmV1HOvpiglOC+vvTlxpj73XkxiUIy+KxxVtR1Tho8qYRfOLXKn
NTUowXHSQhCjfc9HRqnoOo6+iPDAlvrZyu8+M0b/TpeununhHLwu1cuj5tuR2Xgb
z1zm3+nQbxaIrJ3eDPyIi9+HFWqV5aBy15694uSrHJQ+3GnS6u+j9Ul8XyFKb6Y4
Kh35XU6Zvx3l4VgcLVgDJC4zFuEKL7iLseAXT4jI2KRk+rLJ851z7AtQGxZv7vVo
Fb/iGVsehhT6MQUfaI5R5pdkBsbDJcB2w7SGW5Qs9w+9hNz/sXxHO2yILCVM7Hgk
qWCIcpuH+sttBZJw/Aj7lPcFQK43wiAqSY3Oeb3Pzg++nHZJFaaC7FwIGCSz89FG
g/j4w+1x+OUMpwacI0cosY5GpwyhaUCZLotWJMl9DiUKLxiQ1wzvGarakLfrxqaV
Z4dE7u4YVwq8lFwtx1e4bula40jT23iyy7ST+9wUj2je3WLCn3gdIAHYSg05VOQH
qLfvP9s1RdyeNLnZ5x2xdK6AR6k2ehMCCXiLcUxo9Wrv4mIg0aAajtWu32YzNIMu
YWhL1uJYGEIelSDoNldmzrli3hwm5wIx6FTAcRupU1zhgJSqtET5x6/UQMlu6tkg
1rlpPfT+TtYQJxjRo4/DBLL9RR9LBdDDcRB86nH2HKM5rV1pUBKutawW4ZmZqBDT
Wt/h3L/AdL7uETjCJPWxm+f92WiAKePgyD8tNIZVGdJTZTPemfmJlKmMkeQLoeo7
DN4RzWAXfZc77HpbauqpDykVHMLwxdilD3aNhUyUwcpAZIxSoQ0gBjSVmjqHjGqH
d2tIYkCDdHFp0HZVGwGnaLCQf8d8UqzCAR/YTscXULdARFA4ymEV0COkca8a7Hlk
3id+PmiGR6EocVUesNtyE+FHS+C2MptxzkM6jifaNVoOBu6/CLCbCgPbewgt2mao
Q1QW7JZA2HxLowskEXsfagdhU8qatS0dZX6r5LrFGD39qSLMHk/dCFXmdX6PqYp6
0SwyyCo+tENKzngOnf5ONkFjQH5gtHFXGZL4Iu15hoDUNnsIrySKJIulKr8mO0Tl
M5kRyC7iFEdMZSH2XQp0UJ6KhuudHknEfOjzSiYfjeSv4UD/fHn+XMlkCaykSEFt
AjAIMZncLj497iwJQp6NjNukVqFclkbxo5s8QJ1VcYN7ygbZ3JVWypDP9P1jIx6h
`protect END_PROTECTED
