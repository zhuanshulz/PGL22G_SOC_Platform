`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YSAxwDByaVKfQxMSQjcYM7j36akMVztc/wC/ujkmvK16bed5r5ACv8Bqc5yZ8Mx
EMJOpYbHEFHA7pU+bAlnC7327ih4NIpEG/Ub2PM3dshIcPBMIDhBtBiCicHggAfA
Rj6Yzf+B9h88LNwolgrJg+mn2TAWuSsZOyMBws5k7EIwlT7aIdIgznExPIeN5xAR
qcluXThLbLw9EO66QS+mWe0cBlvcXTk0rG6etYzOTYq5F4Bl4w3K3tWmyDpNYb2w
bCVV72QfYG9RS/jqcOqnzLyAZiDo/ARccIc2WI7d6bAw35rt8vRf8P4AgcqdnRCG
GxW/9oMr07RXRYTu0LG9yRBFJHmfrZD3DR9DyCHHR5J90UEVx68slzOsLD0vX9I6
CBZ78kXvHtS6NNpvGTGRVGypNk5uSJsPUGaQdHZTH2NTub+EqQuIYMfWY474OpzA
GYth3b5AzUpKq5niI27lCkXD1welL/ux4PD8LJBdIhxWSgMUmZcCppSgoR5jIuYl
fpW/FWCM3i5tjfhY0/KLIyPu9aBTmtVR342jwAlozcdgoWfXn2efnWuyqxY144DB
d+agFTvbdHmpojFoi20av0uF/DJaj3BNUiFdAAT+HCLqnnzFMhUyu+/34Awc/gkF
9Q/Zv4i7VhzLixADW9AP9aZ8U2yjsI71joHqyz9rnaxSde/Md0f+XnM/eupe2DEX
QZEyG/bboK8Kzaj4fLj7Fuo7E2OXVn/N1zjuCv/3fgg=
`protect END_PROTECTED
