`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cV0HlD+CDNrUkZtBu6lKTh50hfBxetE5wTAliGY8A/SG1kDkSkDumoEu9flaSWZG
kIgi0X/tIBllQ1z5kHLd8gTb7rFrzc/6Vb7OBjDaIdsRgRR2WHFdIJgBLePO0g+t
aGqHyDdN0PvBp8NKc3H/DXcuscx8z0xMGyCWGKOTU1t1f0emaoqrXmCk5dR/anCl
NeWSwEkfkygLpd2XeXBXis5ao66KtTZoG7FHPH+/qIE0tODwy028Onlmlg60kciu
EeX8B3lcNkQ9fqqlaQwvF8OwTFzkl6zwHZVNU8ukzIunF6mQmzmbdjXy0jWrbGzt
X3wH7z+/K4KMDT/g28YpAUfTl2LJ079wiUo9ophRz5z/F9e+NM7UlOqB/G/ojkr4
uf/GxO1LENhMtucq86zGd1ctn3zJG/6P2UnjwkZOZ8+TXpPIEff8u4bOqSCV0Z+N
8EDDjxDwkmfPbU8knxse5vEj/wQZPL3cj4YP6eADlFE5Q0PsRrfrHHTAciSIfpXY
7jS7X65FE8d/FoX1hK3Sy1M/eH5J0e2pkPyYiBntXtiMdX66u+kmm9h5AyMiDdNx
hjNBp80f7I6IK2e+u7JVmxwaRe4xsi/RR/VEmkbbmG+tthW80KG3sRdxN6P3F/Rk
Wm5VpoAukaRVOPkpVz4DW/DpdZmvxscQpcf7gM1TjJmvRkeV+eJVtfBwbJCJU8kY
JC0A97+jesyQVo8/87OkwhJ20lpbF36yTv9k1fgNAVRIGRUGTKAZPSPrM9ROQ0Dv
aW8Zo7zYp/m1BhhR/5YA871vtOSdhjJbuhFA0Y/X6toOzQKTHfSbT3Uopk+rL3QU
x+EedE6ItImwICq3w+lcFOpXMCZ+57OrmO4G5LQ5clTQJaSZfgNzr/Ng+rkAjbGp
LP0MOYJbdZfh0vEee1rJz0PAla0eVS2aHyygVytdnNJrAswhR+wVW9IsclZhfEFe
GyjumhMWHMtv+OJlIy50xMNB3lKIRfp3OzBcObhPF+4znZCfyOdmbhX3/UAvVdFf
DMrxvbX+WQFYSeX6M7nJilOJKsigoGLRMcdUDvwZHZ++YCWPhASAQ7ZR56X8nE92
cDx8hc2PBevOzw7PhiHp5g1xKCUZrVqNgmcHCsXXwaUzJlWI/mYkK6mWfEnWYlPA
3gqJ6pbZQNTsbBniMzVqroEudURdgiUmuxajeL7UyvknaJKWmQ4DHOBhKAlduK+b
pCGBNBNeVR5Ird2zvWbk5d7q8Pz2Th4OlNw3B9gvgYxHvA6zEOcx6I8Pn07pgXyd
NZrTGmzQVKRtrx8YIjnPSZM7qsGNGsT1s6GZOCNwjBzAqzjVMAB04Bt5qOkz/Til
nnn1EYHi3XlM2Qj6lVFB7YMJFuJ6rOsHRGN6ArKpuYw1Rjxexx7qkXjVr8rjvSb5
YD2ZCQdF0owLN9b+6Hr7+AGVyzDWaXWdLNfjnI7xWFdobb9JKG/YAGu2JeTXYS24
au8mF9VyGAFoUQzRKUX0XZ9y/0OCjn4Gl10Ci2G2sXnb0vRGf8GkAVo5K1at/AnL
wcUNaxLDbiFzN1nGzHEAAg44NQ8guKIbwjjEKI0Q0UDkyxVDukoLQ8s/XftwVSWn
voFkTuzkwRSoCSflk6mmaPFdBnKxFz6aCdTg5JzYNSkha18zZ3hyyoJGxZ5Qe6VD
N9nrYEB2DFWlgS8/18xDvKV3FkfmgeqhpAD0AcoDTz9x7yMiiwxqj/uGNGorrA6q
6/jS1jbXStJPgSN8J1/cFTraaS8zhj90VhtCymqR4ZmXCjL3r0j5TQnNGSxcWdaf
DUquYniC1TkROXJld6e8c1OtxiBErRSoK3QKFkhyX+WpeaHQnfXAeg9njZsnlUU6
JlsHRuzi3ES7fPM9xX5TkPpmsV3tc2F6qzyJS4QCApgR9Pv9MjacDRoAHDPPZveR
kX4gce8Md8WSzEVekelyQsEw1/93iiAwa1qACIAzikm4c/FB5JWBi1GD+cYufzoR
/iDBEznJ0pBnuZWC++zELkqs6pwka0YjI5oU4P6F2JwaIMxFSJT0OoahpmARK5iY
qnLtvDC6gDNiUHDq9bUTV4buU7GAx0dMaJqLLGuDH5aT4GKZG7zC3onRB1YCTrtY
jvk4FSQ7UaC49Tj3uwdhZGN9FPDQHmfl3AQsFdDQW7ur6Z/Sc8Ty0wn0A63s7QA4
N51RXO2NmrqxoyiphU4TlrLwc0IwPZMggtqUiAenZMpvQSzda377kum7AXN1O5vj
G2UoxwmYW/kCeNg3jdbX28AhrAQG+a6+6VLvurz53GL9tQfm4D1gHDefbfyiBqvy
IEUnofWGO+76RyLy8/Oa4o59mYGLqKc5yCBJlqafF+ATnCZycOlvTpkOv8okq9Hb
uVAN6DrWe4AxbopQxF9BDjL/oJc00/BNn8hzTi5SGLKpJYT1fdQoiFgZzHgmYmqh
0EQh+rOhLJZZ6KWUkDnmSSFsjVF8xGRqXAwmalOU/B6+iq+fUQkHh59Lf/kafIQW
iEFbZVAA0F4sfTbfOD4lEIp8PtuGGCpsFqaBwIJkoXZI2/ui1laybJ3J/6qmWpTF
1uScvRIkAyzvCZtyQcltge365nkG/K4eKxzKI73cpD8=
`protect END_PROTECTED
