`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUPsWzZMY8eX7auiy6mpKv5F9qtVLD0tic+g75pXpLfVqO2Zd5COm77p72Qd0xkm
G+0Oaf14c3YV9mmaLns0GYb7fbbVBv+Xoi9wsgSVGXI6gFtSAABqf4Yf8SGGnmu1
Bm0MTACczcUlkthBUNPAXuRPpxSoVl3AlmAynhTvAmscqI9Jo8Kguq1GIjD3IRN5
IPC1WHwTNZi6LO/rzLAfrHDgR2CpknAtMk8e5kKYqRbu2B2+81zViG/0FecsaLAB
/Us+YZ2OQ4lsPkik+pZX85eP/UbvRqrcs9jpXYjD5xgoAC7KqgrqXgX/KZl+lPlS
N/D7WgI5TTk+/JOyo9Gka6J0kR+LR8rUNu42htb8XAyqA9wq3YQsAI+9AscLmMQ1
jm7/mnmDL+7UxCihFx/X/BNrTOgaZd6IEY4tR5LBxXoz+InZhGC/58sT2ZvdSBB/
2zX4AxPrNSzt0g+SQ+F04vfjsHV4ksOfw9M+n6yp8l2VQuM6YB2y4Rf50Uuv5/ZS
FBeqXTv9Op96En7JQxK3C6ZsCvhrans20RZCdTRs2bQSQnial1dJSek5MkqtM1De
nir4hwnI6PWX2zo3VJbZy1uIitdjntVU7O/1+P4QESFE7FowhAQ8JLQkYKWvQqDD
dpkt/MYVOS7U0wumKzXEYq1RKXqdJXWREa7JEImpvgArYn8SUUL2vovTyE8wF/DY
/y3CZFFynll1yX68D6H+keh5lJmqnSVF+7gp0dyYgHkkmX7dAwjKqiBh59HdqYKZ
YV04fyzYh7DqdctW/b6ZEBKfzC/zJlqnVHIyiSB3AyEf7abT3Nzftb8bZHztMMF3
HtRsnz5q1pfp4ySR/clUETHxz2NDfqz0lb7HZSJiXl+PfMv1m3HwkvORdncgDkEr
fWX7Gy2JKTQCeLpfOlIIO9ZuVocVlddffZj53pJ5J5L6kOMDPSe6jwzCe56U7SnM
Yd2HfPcZdLktuK5e9gFFSBmeWECmcycbqxq/tvM9GehqUFWWHmIpzLdmcldZ5rc5
UvaAa79x2xViNC07r5H3J0X/yCCljxN4tROkjWO6WMTan6hWC8CbZK1dRSc0l8dT
gOq/ZDna+9DVpN8Wnn8N8ORDI2SsxJ63MM2iXrVEadoABp69ee1aXocPM2I2hVy0
0b9yOJQjSyTQ167WiOjP+HCKIbIuwh+Ah6F/saayqqJFfotAYH6eVufJ4tJGLXyc
FGoF+thkAaSYX8ma9RFRMJRmp1xiSXvJqpl/82cFbwihavNpRVP2A76OyKirLmKF
ZHV1IVxxwRizqul1CHNpfeE29z/XVn3PsBX6iTnSCwW+zTtvJtxHcbkcPBLEQv5l
cD0LWj1hBWAByp9T6PGlxzG3eus/Onq0YvSlU124v2Fie75NuaIdNRyZL0BPst1G
xvI34iok9JtzHsGcWHjVNLHmcUr1GyfEYk8syNwEb6ii/vtJexuEmv++4byi6xN+
4AHRC5Ibq5MSmmGgejXqRU2jb54qq4/4GRCDkkedQ9jwRlGq1ZK3ncPXlTN4qnsp
un/M7/SXgt2JEG+Py6F5K4cyQamOUTNjK6AUmTHP6cJw1sVJJqccGfYxE2/eEOyj
ck7lqD3JuziH3CHVGHi0Y11T1uXQ0cyHRSkpWe3ybXDM6Xgfd0qJQzgNaFKpQ5GP
Zk16UsRAexLxM6q8kQfpGjVVV34uk+PEfvHaQcFEMB0e50rkDE64wPxarSC20Jqq
UjVseD8kPfx1U8UFJcYDsqXATWT3XSEQZmLU33rjpm6lLUOqm+Ezj2IThNjtg1VN
HUZiLS/34S7QfaLsDNPgpYayzjESsSqs4xcZ2nApRscALIwc/NpND2vaS6Ppdemm
5o+Y9G7a0gyOex2HzMdP9DwyUTe8Aj9K3WW/8WmKPaKJjocabN1QdNrqoz1YBww/
m9Rz/WcBPR5GqopSELZqXRKgQlrpZn/mXtSnRr/5thtuUtEbmdvV25nL+uB7PZN9
NyYmvkMWgMSl98umQIcu42rAczi9I5U5A+b4MphEX4BZJis9G0jQwQfxKq5l4puw
MuLQvxYMVwBv3rDrrt7vEz9qWUcgeW7bdm3VJ6L43IGhhoKOIZQEPXaXiI86c3NK
QZXTjFXMaAb28R9PpsSOtz0BUgsKUv+6eLlqFI3G39Okt8PqSNz1wA37UwT/P8sA
xkMHnuGMYYanRk3pSToSMdZBJ/XFy09efodwJokJVWGnVKzQKxdbTQFryV9ahBNK
HFnIdk7b65pS/oUo77PSPXfTQoxK9+r44iqGn6cgNS9G18k594G2QGpVjEFjVlvD
7x5ABl3lmysUAPcrafPrp5seKyR8Y1L4iNZhXFrFk14NcwPxUE2tozochuwab06z
hrbkMCJghK0n1eM0KT9dNWGb3VSSgJIjjn2WON9rMvTLvyrcoIb/lAoin+cJa0GZ
Zw21xTsV8uangV3iRGBjx6HHOIVQwJY1LaaupdPt2W/Gai1YzEHpz/6vd9J0bljI
0kvJY1NhoiDm2Yb6ac5PAmF7rrmPxZ6tglhNU7UNW5+XSvSGQIxrvniHaPYJlqNL
MqiEeR9AY+cz/veaQcBzrk/ShnVjWSIE8A52waztbqKmc14Rj2zjnS4X5l0pV24M
geW2LJ5mwvG8P3Bw/FrY1rVpAKnoT/1v5kiY0SI0hPI8T5s+hHs6uMvjIyGWjjtC
gjWaNW5FgOgVSEPKFLcvL91ox+r05NoLUW/yBY8Elomqsb224nCp7psnQebjv2TI
86pmAbLzQDbgEI0ztaC2aaDgzY+Pht02iwPTgxBtIXFZL9pi+cL41WFtH8vlnxnZ
O+nr5kG9Bt2jzkuibe0leoT850AUVAUD5dcwtkg6X2FVDMCp06Twg3avXx+BH0eC
H11uf+M2+LfQtBBVfLVLrjBseUlKpNW9mCKMyjO/oYcS12Kt9Ajs7IQ8/cKgSPdK
ECA7IH3juHkSHpPMm2t+1iv5FllyMgyeEvhdv9BzDVLqSvKvmXwtsKe75NG6WWmv
Gom+VH3a1VHowydI01qBKWTAbejzbJ2lIQHQg3o2+2sYthj05WrWGgC/hbgGdFFA
UVDQ5JPlhv9YL/cwH3xR3PBaKQbZN7E/UG9FURFzoEq0fIQStMOZotYlhru4gQzf
CKDCmtC2YKpKN29WwKEo3a74P9gukf6G2wlEqr8ZR38+ksi6QAK/J4Ezx1vfA6mA
WYQgH9rqASGDtti3b54jERJjGy0qFCUnwg//2rZI8HmSppfxvH9MZ2MzbTtccFQD
AZ4FB2OKynNgYbX+2SAoRfQ2jvVe2TSLdoCU2Jv+R8EniRDNlX+WROG/1/F3uNmd
lgjsZPfc1o6qOH5zUTNoLGkkdctGhbUZo0fby8frukr+ayhjolJcbmKKs5UbqcVv
t0qBjSah6AE/ywlSNLWuGr/UnasdsWDtpMTtI4bmOeKVuSq7Vk39Xlk1tJJEE8q9
hzUAkl+P2o0quybZ+kRPZW4JO9baOnMO1Y1dOWRHgFjyfQPFPkxVwai0x64PxXw1
+xTI60ChPSbBpKk5LeEClVOjcSUk1hBjb/Fd2DvRPf2WKWaZWG2boWZwRenJuuSu
/ygiTdK/aH64Xj+2Y1STHjVLnaGm5y0AcBTXoMsm8Zjl94xN1fD2Ijxx+dv3I0u+
RHm1dPn+tF/G7vIj/Nq6GsQaNA2XedOFoOLmMUmXR/vhDMGNgTTIg6b6eDT1LZRK
`protect END_PROTECTED
