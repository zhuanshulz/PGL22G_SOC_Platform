`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6SkIOgacy9u/IprfvF6nEpkkMVN5+Pm7aeIMIl7PPP4csX1p6IFazcKbQCpuigJ+
CrG2SnNsNYXuF7y9l8+KR+2gvFMVlDXq4FRlixgNJtxeNXzXkjhJjKAPcYCpODhh
07dftZjEYvefO5KkiCryF2xGlCEikR1YHne1wd7qugLmJj8CiHtviOkgxJJrPe1D
DC+6Xk0apHYNxovoGsuDJUb2aE3gPsVEjQjVWiZm1+Kz97ODc/y1mbRzYh2Eioul
uRmgJvyhXic0t9036Ez6vl0r9PxjYlSdwdh3LGDDaVVTezIUCl5YkRL7ge/J0n7L
oIPSHo+9uHrN2NiYqwVc7ISuil3r+2MKlIkcyne6f3wLB/YKR6jQIc45ybe2ZG+p
bck3eoqbClVoaEamV6uTuPrW+bbtsveRP2IFle5rgNolwlF30oYSP+g95ua4zJ5N
RqTBLE6lpkzjpePTS1O8RmzwMbd7u0MDz2WvfGFvCspFN+1EhOQ2F4C4ClzP2N5d
UCKAoN/jQO6yROyjD4TewXLPid8Ywp8s/MWg7bx4v2KzsMKJlco5fCrbovRRE8hX
c3Q7LjX/FwO95A1PVt7x3H0ZHTVuLb7ilCSd8pQrJC/ef2m0hWLvsIGZr5Y+2up1
Pnx8WKLBd/WqY+B5b487tMMoE4kQaI9kWErzXGG/l1m7/BL6wMVhJXyVSZeL5si8
LaPfUTO0OqFU22giHQsCM2kApcxHZGF9dmjRx2WCzgw+BuNI96d3fXKGKaXM6Hy2
XzGGmxUXtDwegjR4hqExiCtvfDGGnXwrHXUqjai8Olm1/8EiFGNIwgIc9yQwJ/N9
4zQgxTb50RyiIAhcc1XRiiWfR7+59JWmJ3VFDkBToM8PF0f+9WDIW27up82PZ+Nv
OLq+lE7DKajHPR57ZmgPcIWHCd35dUzzeO1tnyhNCeQ=
`protect END_PROTECTED
