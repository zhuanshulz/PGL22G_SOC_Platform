`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDk/b3eFEPjGXrBqSbUvbakvRCGCO2QLGND0uMYdcJMbCQVpWx0LDFkTAYx+C42q
Xbklt3s8MUwE5K4chBKDfxXbi6/ZvH5B7ImojUfDvLO0IoL1R9TzEVm9iubXVHI5
eQQzbApKJgyzlRZYGHnTL6k01QFwa+oD4F+q8o14JND55Yi4P5KcUsc41+6Hj9q4
7aAzdlUzo+44PjZj3SiSJQX1Ky3uWbtmQtldJA270fEX4QnL3zlHcFB94qiSAVjW
7XkHUuJoajXIiPCBessuYykuFJz8oTXkm/ZsDKliHxkCTnpu5pAh/eiq0oAjoCUj
qNQzkf08btksd1gxtpg6mlLJPj/7pP9Q3+0ZNXANFSswvKY6g3fw1FQ0UR5aaOAP
oqTeVmasJ+TJOGwmHSEDqJTl/idRCJBUStOIWlHiAks=
`protect END_PROTECTED
