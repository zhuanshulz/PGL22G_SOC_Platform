`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGVbB0zgBuZzdLcWJPM5Bd7Hbn1udqV/YBkWrlIkH+y2vw7nX4o/ybFIKMAgvhMh
1mGsuiFwdUuQrZX/pe9U68FTUpouXwV+uKA4eN2QEHrQVZjY61m1nqqbYYoBdTHD
4EfkZUf1nRDuuMCzh74ypr7t1caHRfUU7Yqz6wwRhIgB+3m5d2UhhmJG8RQOvOiL
xg9qNN/iL10K3BGwxCTu0ah5NdUo0Nck6evvuSFVU1EV/YowpN0M2R2azKavtYKY
NyhFfGwOewKkOVU5pAbCUyD/mDPMwItYCsqwQBMhsrjgbf/SsL/f7lsc9RfLOiyd
z5Pj2p3fkCxRo2SCA3U7tRCdba7PZ+Uu8Y+upRu1Bnqxit3U394mC1sCITPS6KSY
qJLrJDuG3670Fm3NiofU/gVNkF5Uh/eC9VqrDNHshQARzGnyEJLA5XvmbWSq+jgp
Y3Tkgna79YRpfbnFowIJZ9WVaQz/80FCjw5DN2TdLmUlzjPhhHrYwlxz8KiLnxTk
qgy2ER9krHJhLP+bdjfzgbWiFGxLyffasBPxUh8/9em3mMO3ciJDczoyGSmw1ukg
z60dvQppObrJJhkRup8w+Z2gBHe3ObfLndwTeLAqppujKNm5KeMNh8P9tQ4jf8PF
noS0nDiVppHsUxmhdYbGOHt6E3JsWwYQ6yEWME1uCWb5d0mSrak96uEcFkb0tBcl
hl8OJ5Z5FRqM3PQ4g0QMghkqxVP4JPAuKbvAjr7XqUZe4MSFJWml4s6VR92OvKqr
jmd2UoFBqCxe+CUAifhrWXuZeUXGXQUQ6kZ0LIKvE43dtFjSvS0sdYlvcdlI5FDq
Q49zjL3g6VRyNLD4B9LWRUYSPrf+E5o6YFnN0WHS6KHC76OKJj4Q2RJYf6Fo1jaP
GWQcidsf+9cWwmNBn4NEHc9GeULTWyTgBYgZuWuMtzob2+RGIWule6kf6Q5iAiMb
o1j0tQs/8rlbscdI6bKYeSO2n/nwRjK2N9Y81jChWTnygkR7PK2asnYfqIxDk0ac
O7fnnujRCoke16vE2CPj2HkWKkD5SGRKJbcKs59iUWyM5e6lr4Fas0JRYiPNh7ex
f1GAIUAWAItj5T6MfbO/cvkyJKNKC3KX6yDiwJFEcI/ePJOKdzLmcdYshtRzj6cD
UGfij2+RbDwq4JqdGL5N8y2r2x1ZitCHGu99Fl8k+eSxywQYepsmKt8G5Bg7QkWy
xOC5spy4ZcqTQxsEbTXlbozSR5V+i0dV+nsjO9uxd7ElkCaTQSdjezh/MuIqQQoj
T46eDZU0b5Q39B7CtCfm4iNJVVlIPLG6GhEG83JDQ4Cl6jaf1m10ZF5DtnybJAoH
Am3BfOvAG2OyD0akQfsz5u3o1J0ncN3naY0Ij8Eh4h1gZlqWApTEjK0Nv6q+hTz6
x4c2cQr99EsxmrSyrc7459Vn3xPhzZ/r8GvKWqYgj/t2RVBQ3Buum/aQ+f69r6w+
9iz6kUwGCh3Otvod7lGChATjziUN7hjJXJixZGzI+K2WxW2cyUdKmK5eVqnYQsBA
1h5op8IfQ4gFqS6D9xRqjM8xG7eLljj8l6D7L3snYzzw77W+FOAH5Q2q7Etfqp9o
VK+ugsvhYc0zrLBXT2PKufdPG1KKgZ8gu/2XycWnNN/x+q28vXVSJuH07P4GlbwJ
DXWc964luCi4zpPOvS1gUXfI7dm/PfdYiG+gRMfru6LJptmN0dkitMa7R4Gwt/ew
kB5YiaMxFaMiq5Pyz6g4gMsGEKj5GslpBohWNNpdyeTydbm/nwCHDnX6jA0LuyKY
smrxAO13uUgUNogX9aKA9+06sSLr2pDvCHyhxOssa89AtRJvBNB9Cscqt2QkvVmK
`protect END_PROTECTED
