`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/LTvW0WMGCowExyhZnF1wtX5pmwvzK1uMFX9rac/g0Pbc0ulhgJmBQ9QZL2DZy37
L1hxSlWEJVPQi9vJjBLshLhdgyUpYLM9XrHXZ574vx+HtrXiKk9wnsSiKrDzHKJ9
EJCzLVHVIIerUbP3Q23Hj0ayUVlXSfdCnoAFDAETC+oa6y8SV2wfG7pWpPCEl7zn
uc1JgYyy637iM9djlmh1iCJCJsSC0dtQvIfU3nMoUK3qJc9+hFzIaREZlgzUWeg5
Ik7dYi05Lrf16jtzKf9uzVuv5YPZfeZKxAwgiMDl4KJ5B06rZooWmNTZ+EcmuZjG
9SL4CcRGf/E5HkR9rP0Wus95BYAD1e4dPm60JtK+vybeQYXdoDQTyw6N02xJI4I4
bvOMui3+68eWL6j4N9PKHLMxb/PQ3g7Ro2fGimuE6erMd4q9NgaSuIF9jF8iwd/2
VMCc4xkX4OHMm2ZtshF4x0QNyVfNhSW/FWggOxc7ztGc68mamUTXwHqsTrh307DJ
9csBSlGK24SDlA3R1QOOWs0TDZOuuZyMqmchxrmManTgBa+aujJU9vm+VPGpBXFT
qdtkL38ujANgMdzQxIdszqKhBhH6wrgS7mRjCdf6fp/I/47Ouo0+JbWoDyEW6bfY
crZNTshyaMD52Tobd97UF1hOeciD/f/9bdgnpfZ/IVtHMG/ECxSj/cCj+MdJju/p
xpSwrFYE3jkMMMd+bnkRIIMbIdRQUK7bxqSSmWoNWyl6btYRcRnCQDq20dVhc3mB
`protect END_PROTECTED
