`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ITfE8/dWKX6xNjvJRAMXJBi4MFJE4ZQTRmjrckF4IdozRDH4/6awvwpGES1cGupD
RT07s6hMbLCK0jqQkJ6DHZP3doaqRcZGHZFjJ5bgAssAn4+GpUVUHk3bMn5Zj6XT
hqTMKIZixs6Hh9nJc6LG1UFHIjpSetdqGPaYtg9ejXgfgnn5WvWeuqyGoNq/BO+A
6gtdAZsm2SyhHjVQ85JEJ6W+ENyl0rztahCinICljp69EX20oEFfPJb+1aXwXxLZ
n5A+b5Y0K0fJbxOHfu7iZRO/zRAQ8KbaalcLiNg9C9Vc3o/RaUCH7pJC3ju9Fz5l
WQr739MS2JfKretHyCsPiN5YuKaXDtmu56Lw2GSFDtq+yPAlwNpZ4a0KhKmlQ/TO
oVNxhfF4NzD3OtXDT8kYtOkOXOnjMjnqXZQzrRreOAFw9KYHoeLiflrvJTwZpKho
wsmO6rBN51wmz8HKGnzt5AJMJ2SMm9SOsUh+WN+P1VZsIVt5w5CjDsjhPrjLRmNC
KzNi+mCBWC4QXFL8nvRynyL4N5SveLOKZq+eEI9VIf/Fk06txptw7Z17FQt9sor/
QJx0lEDhxXq5LefkDGRZj0YqGac4CAk0fcXcMYEpzxkrKI+Al7Izgw5BTqudcMQx
71F+rDf70PSWodNs1y418wSb+WweZ9pmC6i7QCsPqMOpnRfADnkNLXBW19hRkkgj
fRAN0C6cQAJPYmRDRljCD3+3TEBuiEREQiPwtim8oL3/vjrutFp5TWUGQkOOq3zs
kYQTKKlYFXW9QidW8Z1LTugh29iElyFb/8XIVUjxrpglhYOtoV6bDWlOH5GU7Yuu
qt0jMMkkIYCZVSAL6yDQID2aOnk4jsJjv7EVl2uemBIXuWskvsJa/Snv/12XRYBZ
m0vTvPzGG0piYrfLuT/qhOmTEnwXJAUgN71icuIQ1Vvd6D9+V6G6lUyxE69qC83j
VM2MByc+TTi9nGP1WRJsL2i1ydXLRQi6syeLnWGKH3Pd9OZPQDQi895s/AYnzRFx
sjuW3QkCpydZ1ym20SVn7CKdKLZXGtH79iokz7FiODK5RNC5QOr3xg55xd3yhEQh
9jBgnCbvMebM/l0Hf3g6L1Pf+n8JUIUGFElwpALsWo+7chHcMpADkbDABpS+I6JJ
hX5xNaszCnixaG48W3FUxw==
`protect END_PROTECTED
