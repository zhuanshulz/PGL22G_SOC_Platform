`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZL1PpjK+bHayEjdDFrwVm8WGiRx2Gs8QKj1B7YF+NOrgX/cp1FnSaOYkOXzrStB
oBJ/0ZsNWd+RqAFo9H+VRCNjHkbgSx2B+bs5asxe6/bF1CovCV7cRAfzugHStjDn
Nlx2o+v9+1fyE9ygXezQmnMuBPv4C4tn5UyNYrCVYaFPVaVMEKYN060C4AjEc2XF
NjRliO7Lz+hcLUqmFs9eUkCrc6cULna6nzpVsWlPGvREldnSH0aQ//bILWW8z0Tq
gzBvmYFtCSx96C0jFvUQa1MMSg7fjm1Cl9lNgWngSmDNGA+mwDfhBXfJUaPdlqmc
vMCnpQ1VOyvip8OqZl2dA4QQgUdzHcLGeWLy/BtUOvCIE/vgO48RJZudNWDJN66S
pkpRK4suJtrP/fzlAVdbDw5UCpgfhZAwDHM11WaRDctVU3hiKoLZp0z2Jm+DQjBB
5sukUmzPE186UGDmugmWGtMbUjBaxvYtXtPoOpOjij6pbuNErR/31uW3sJAhP7cJ
C+GY0RToXW49lOOeCx7pVVpSBE9NPPolKS6h7+zLg46aPpGRHxaay8lBMg/ciGDA
y6TAcmoxqEOe7nnevAhQMkuCkPAGEWAFRz+iua+kJaCN4AdBoC1Yb2hS5H+hFFQu
8f0XI34D9bq8PWqQ4jIRLGb9Hb1wC2YGYd1q35YUf3p2sL7Gv4n8TlotMhwe4nt0
m1FqIcyWGHXt/bbuofNnP/UHENC2Vgib1gihlTsyIDjFQDwguZ/1YIqoN0ljS/wy
S2IZ5TLZMwIT1gnpyLzNaS7LYbbnMKRL0Nf/h8LCx6qkg77erK8sWC2pb4cqnSdN
tBTcOUXM4PShsC22aA6xhkUkW6GG8C5r9moxesRZFnqXBQZp+D5IyrLblHI6g/ew
omDr8tA16rEYzvdM7tLZxcOmo6bxX0XogjHwhkETlWutOF8VRHPwjv7BpWqRhH9o
VdBqVioTipRXPgKLD7IqKQ221tVDk9a6Q+YU/lOTz+/KRH+sPH/YNx9WWF8+0YqV
Ur5nBtpdpI7GO8f3wUYIBBX+4a1BrJJ75froqSLtYGVj0AuuTRpYs9NI9ee1Rd73
EThBASo7Hpu5choyxbimLtrSI02BDqg3iUQdERi+qz4ZJ0ZrPSOZ6PujRsYOd062
THo1yT2jHHS36d5vqS0cRBzHoY2Fd322YCOvjt5ORYc=
`protect END_PROTECTED
