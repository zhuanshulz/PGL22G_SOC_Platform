`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWj3chQZN+H+V2YtC1OjuMPi1T4sbYHS463qPIzS1DAJv7uSaBj3hz0VIkPBQuUM
ul2genxWYKG4LML1WUZB2nop1S9CslR4Rt0ilkOXPlmn2q6aAou+O7rNw46rBOH3
/FMv5H/ZvgVnnbHB0b82KEd+yAPlhjOt9QMC8lwKwI42xNnuBv+Hp65yelLQguJ1
MyEcnWuB7kOJKWVACuslN+kyvDC2d/zB/9xup+y5j05U3AZBMiWsEZ8s54BuFA9Z
mvvtxqHLn1OPlflnpDLi471fHnDJFh4Cih7BiZGPiL7T7lGjda3yd/LaA9si4+Zy
7edkc6EIekU1B2aWldEmRw9t98wlLmtobqIfmxrSe/3vpiTZ7oZMjGAXtffKE0mK
tS4N4e7K2Wxtfy3zCqQQdRgWTCWsWWWfefyKOznBOKJYZHnfTqxun1OqQzqrcMYK
DroRy25mf+kP5+5F1f+zlaRPGEIwTzuHjrNvu8e0tmURbZxy2GJBWaRcpg91yVDU
GzBMRrKxnLIj1DmbFLCy8gET2ySpaVpVrzUnE+5Je0nHg6s0NVod1iM8yZt66bXk
JMZiPrwHjTiVSSQYAWLqpsAikopghfPOe/96s44F2nM294L4Kx1jlWIBXZaWIZnF
rH+LGv+j79Sba85hpkgzxjjD7Z5AxZ7MUYJ+y1zCaP2Qa99DKMJz4T7/yCQXIFhQ
RwLlqokYd52ZW3/1dgUVPsKBdWvHnd+PeLC2+UbxQrVfPWi++44qCgpr8ushmu3W
MncsG6F60Oh8OSuVnHzxkGxcVJnQDwtjo/afaTMkn84bISnaOb9ZA/5NXdgCI3Nu
/Oho2pquf2TQOVOAcrrYkWIn8SEZ2AZBiplE53dSqu7L4Tm+KIKiGSZCQdATTXdF
fwEYmGJmPOi8Vnwws+fRHro2RmP3Mm9Mci+G9A74At/ZAmewFL+Uun13Y6M1K0Wg
73x5kjyGsUj5rf5I0yhrZxsEuLNXIvyl2HVFJyQnt7zF6627agxo+YVMqa0kgI5a
mGRtgnMgDmuFwJfA+GZkgjOng2sgIO2WyFtHwL8hsBbBY6HJ0Zw8S2EvOkavHXs8
VGg2ZXNc+w1sKyqU0/QrZbOT+YncjLh7z/sUq9uEdg53jmoMFxWix16G0etNhTIU
w1H81TlAPYRemINY6O9Yd5HcinMyhKMVQpNjpQ1Z+QqbxfEBRUTaZ+swjBfEgzat
Ed0yciDFzWPoRR1+oJtq6QmQQtYdK2KdgkSAzJGZaH2QkiUe9Fdqv9jmPFVGXyGH
Ucsfd2ARUmLkYxxsP/NOT7W2nwg3diuWV0708lTkdshTU/rl/N7MZYdpxmj2Qsa+
atmS5+EIVQFDvjxmgO+RkkHbZhEDr5MaTGO3OGX+r2IUeVn5fTIC3vdmw5cFy4yw
0wJ8B172c+NQTZsDYTc/t17uoW5wTNGMhcmBqyYwrizHo5nSlW0x4oktMczwcvx6
zluvhIOWhaoNXtrdPzYn31bzMWUXFBDxsg0u+GXJUIZozWIzseHAtu2icDu7tUzI
RGqXSruOPo33vGYYHHBnpgRzjDGy4i1fJF8Q7HPg92uDhScjJkXKOmfvbC6e10KA
WKm0OKWxYrfLEbjYnDuIa6OWMVFSZU/KhOIlj9YOvxaoH+dFm2VJ8CKdIvi9NuIQ
PaFOXkmtVR9oIjAcmAVM6TZJyYcUOLpHHR9ewbuwdi6XQBaHadl+zXWy+UHfOk9m
06+EIOi48BaxT0rAaqY9KhXF3r9gjJ2J8BZ8eAH7sFWci9zufA6gToYB2pVUezZq
FWKVp8N35oXZNwhSbbN2nWJbPob13qmyVMR/ePQZQyaWd1Eczg9a1xq4tyTRJyjy
ztiJMArWpScpx1h6iK/zT1svY7jEUbJaGFxKZUv+HjUZjP+CzEXCsvyOhzGAi9ge
N2eEDi+QWhZ0mzdjrUatOH338VEbLY0+u/vjxRD6Z57jLqBZu+x1c+ZmRozCRbyM
7Iy+h98UQN1dCxLAx5Y0j3JEjGma7YLoGSjgbf+cbzbb2Nib6rwC8et4puPk5qZM
js5KM3kTVlvAWOrA0QrpZQoD7xCnzHh1iqMpaJvplRo4Ht5pPFSNIU6KWnBmzwdG
VvZEPc6VP0xJYuGXJ6W0NOAK0X/7pEjaQvPgsbZptKOEeVOCCxtQDNJbuE7deeu5
AEAm/cNpDhldSwQXSWOkLmU9B85PjgEVjvP0WAspOcHMbyCWYvnWtRQMbfgW/Zkd
9D/BNnzdn01gkLoymIuBE0Y/9fQCS4pKFUXdOpSvFx5V06bVRdrNP+ORoS7L/WJL
KtQv3on1OdwhCtiJF0e8qnluOlHWcvvfVvFAYY/1vfRnWG3866pvztMsXPOEg+21
ZYUgHtux+U45G2qiPG/Lg1OzmxzYzAu5q7LPRpVWw9LeylS4zTOv76kXlIv7TNPd
2PNYfxlr1pA0qwG0CWTkJiUeXdhOPMO8vg6mGEpy5ll43iiRIKSJqL4JhFAg0i7J
2+aS2+uiR2aBEBttCgGG49V0yAewscnASitCxyjgTCO8FHXXVbHrF1u/CQTg37w8
cl7Pyqdd02slLowvFPgClcuSYGHnoUyeQ+p0+EDUtbQPCA0lofRDW51EI21OvIVK
G501dhmCKvZsuGIigj++DHcMV0yNSvtheLfy034sQWMs37sY8Ld3ceQ4sjAKA0OC
ZOfVlcr+CigLMvCILv+cfqVeB04HPGoXQSM0+tUd3n7gTB4H0QoJEq0YatgCmtwm
ANdIGHSKX54L6bowucMNoPyOoa7r9yYaK3gZkJQ3RrBYZyfZyxfji+JjngNpbuuq
NxgK8eB7Sj5H1V+FPOdagdROTOux0caMVsZbClgy+L0dfaC50Kn9AlIntGE+dO54
2bBYpa7piqB6g2bsufG6fQ7DqCrxjvhsgcJBd9uD056A0WVpR9PH/C2z6BTdgTKr
pzLpPQ0WdPkF7uIoFEKOgeM5W4JnLjhgKPa6ViJ0bjnNzbHs8my1iPq40izAGaBU
tEskMLmNH9U1t6S6rIOurbe5Bfo12OZEpJLOBrul2kKt+aqrLszwZh+iCm2YidiA
nHx2DOoli1Zw5O5eXfHvN1UlKQqIUiPiKP2bf2DHD0TjZTsHf0c9rGUuy6t5cBCk
L2EMi2hW7Xw900uof6U3zwXJq6daZPPo7R0Hx88KeD7T3nN07LTWgftV26nvDLAM
qmS9zBB+V5gkvCFkQSloRDR1l+c5DKeL/gUEmpCtPXT04SeBC1XC6kbMGGj9aZfq
FCPwvmoA+lehtOQkqiCfS/s7fv7JMTSCW+GS9etICtpJbIKi8IA9G8t0cD83D3Xg
CJgX91AzwyWnXLGxwn3au5hBKMkc3t+iZwdeLpbDsntZ+9KJToCqZszJ/NjA32zS
ucaotnmXvkvdAa4SEKIyR/u35xL1Wr6zZsYUuoNkWzqVID0583SJpCOU3gqoyKFC
MsDJ6k0hbkIlnxgoAvOUJPx9PzaCgnTK/cx7DprUksRjU9fJb9A2dGXe6jUrf4xH
Gmjpx59a+YejWhs+qM0w8Kc2eaNf/eqJWMamcs+srxc/zTQ/mF6C2TyFaXezVBx7
8GnANggQ/R16bMOQvuc+amVufj+9dJn/BzBTA9e1eM16cfQRmOMMXB0v2L0n9Eva
zrMIbZjBLPB8tZRSoGwZWxU9o4aAaWkbvT9NDrCt+0G296hC46vUtHW187+WvAm5
kiib4X1zyVLexfLI5oOmDIeY9U4/bMOPi+6Xhewh73r/784H3X3HdGx67Yj3jGfE
u2J5MqoDV/ySWCtwLJApbOBC2lB/TZdVK/oauTTdWcjws3PO8FdxALETXUukX+zE
Y43VV3Yo2E5vYGQ2JkHBH9jkZxdQe8y9sr8pRrITdiJunesiwuMWPu4m/o+PtoPP
`protect END_PROTECTED
