`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
usMu0m7+4T3yR7E2GekeqRbPFIz7gQuyVrLB6kHm6HJE/ilciTuXHSXFCai/BO3U
w4MrDwzheLCWm2L9eCEx5BT2AxV5s9jxcsfy2xMYSNN0RWX80J6XnxDEcKvUO8ob
ULbjqKtDfEcIZ1tuNsVaOuovfIu494z7y5CSHPBhjbhAx0JpL7o8Xm6Y6sZo4Pu+
RXkV++PhYOEmLTaHLo/LiXWMyw72JYGGwjYf1Rspvpo+aQ02iG7vPSJRx5Mzz1lJ
kriIpOeH3SXsKoYaIZyywq8sNk3TiY+75iSdG0OqrH7K/BFT+AkfXmPwvpOz+ekL
1Mx+PJHgeGiIojnGWohIQQmNGkH/AYyPeQvkAHIimDIXDj0VPxKD5a1ZQ8voHBQm
i6I/RFZ8s7J4iCqPcjX7UShS3h6/g2GVthaoikDvnfZWs3TmEAJS8ZzDRZkza7Mo
ZKpQNoii2FA2dgdIUwNxxe6v0Eqsk6jO7TKe10nYKyFEkF7cbRnX68pru7cBOCkw
X++ukfIImL+qznscS7GgPtS8+Og+xyDXq2oHTN/8lTkJXGyfj6tyjg84x/3UlEJO
jwnGJMuH6q5X07AzpTcKYLBL2r6zu5WvAuYbb6QghFnXwsuPu3RrsnzNPPJGPRJt
kYoQvi5ywkJnaGalPBKV00dYS0d0dFOXXxMgzsdH38HKzuUQgc9a1aBzKDX/CwcP
O8Zn4lehvBtMZeK+/AHEp7hDJIH+JQ3LTJLOs5u7qzIvPnrIyB8qHbL4tfwtyaJC
wKA1Tn9Ibri62M0Q1XK9Z0m21Zkv5IHhc1b97ZJ/Kt7xtaQvwFgigOxvTClNgSIp
bgzOCviVr/qkUtSKD0Ak+n8KxJVH2NJFsxoIXZm2wukZfzR8UH+zI7NU/yIr/A7T
HjNxl6xOcIpxx1QbzIuSVZhgar7wbWOWnW56qBai0JrrxDz/4mQK5fyExyJgVhkO
8IOOAt6QP/M6zLURFfab5kzfgvPhAI3oVERadBYjfi1VqqZxhNqjWDNZzqiRQlG7
rbb2kE5/LBC3HjvOYERCq/zsX1JN3Eh1TaPxf9jlNWDeP/whKDuK/zmWZz33tz2y
3Xj4InqqhET4Hn6wrR+ErL+oI4pF0YvDrit0/3KmNtcHHMAD3INw2s3N9/oXe87j
m7hVzBDkZ7H9RCfkDY5bDw==
`protect END_PROTECTED
