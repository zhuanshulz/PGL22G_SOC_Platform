`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ihL0PzZz8tP4WdZSqArWcKzsB+c66nofRGL20GFmaNEV3XIrKVGd1pncGnOxM+6L
9TNf9OxX4itvm62iWdpGAT9LfTsRqTRnRktNFa0jeGC8yBR3szePyZv4n09YCK7b
XyW+/L4FwK6QmL0yly7vSt15neOnaHbCzyZujPArSdQDwVSzgp2qDMJBUat6vuTP
IPsfblh/cdzUfN0ZCD8kkK+vrS84Mei9pJXirbbdDxpcHZLSCsoQ7r9MiE72URnZ
iOBgxgfL8oeP6jBe5bv+uVC7GklGsxbVFZqudRxy081+pW5WRRCP6wqRK+jVONWS
qexdWbckgMPSRJSVZOtRESMGsfzTuRe6EFkaDf9dH0wg0zseHhiRdOOlK3ljc/cp
ZphkSc1J4mMbGOVKYpn977Qlju90lZXr35xuSwnBRlIKLXdLOrozfUKSdqWaWLFH
FEtj/RG1de6hsTu06RUiI1jbWvYrlILzW7hH2G03ECSO0gmxDeN1Am20Eo918YZq
UizdRLzryXj/1AFyk3hAInAqj+5c7KqNnY1cpeJx9lnoqUaoy0n+uNWYpJrehPyY
9VCELEvnV8BIaVDwe5t6tQ==
`protect END_PROTECTED
