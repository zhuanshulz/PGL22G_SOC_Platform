`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1RG2em8aNQKrpz4Rvg5NKOlhW2DnAEHcG2a4PLF3GR4HF1bzy7peYhLnUHlQghs
mIhGehAILelGCsXEWn+z0DiiHVrunhCpUcMgIRksY2Oxjk6inz4ptjUDVQHTiCqb
hrKGRDWhyWLlEURPLqZZ4bSwX0OyNRDPDM0MU1r91KlVcW91AU3yJ9+TY7AXWi0t
IDzm989PCmNUFazz8CC0HmSKQpBOqRhtVLLPc+FOijKvUR4/spI1aJvGI32wTuHH
PyIWI1oeQoub/6GyigYiCH8dBKuCMMV5p61+rwFzdrdW2J52V+ZbkLD2tDFmjC23
Dy8ry6XcFhftjDbHW52SeOldemHcc3K2St11CBOCj6ujPiYPA3LW8C/LgpIUGHjL
TxkwlQ1J3sPPPFVGOjccG9IqTFhr5TGKyEPhR0GUo9sWfRHv20jOYiq83DX4yglF
q1bTbunls0WWI8ms28ildVOIl+33+cpHK0qiB3C0zWFr2N3wPeGeZovIUgmGUeho
XXUNEZqVl2V7D3e6Vn9Ba48uesKq3mEcw30wYw+vruG5dCH7ma9oDB32z6iUZh8R
hUZNtvi94Se3Ab09IhmlYk91ftZbhTQcy5eEOCcPqjo=
`protect END_PROTECTED
