`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+bGJzNJgZOiu0gev/SINH3nfhP+nHLpVcKw0XUa2K2yyKmp6wM7qjSE1lnNfaogX
xIMmcNAVPuH45SC6OyVwyLeGea5MZSuQFC667XyiCFBIVN2hy2Vs0hrPhFuK448X
uyQq+NqX7IMCr0MORZciVinZ9xpdDWJR2mZA67G4GirwQtO8yHA7zwlsgEXWrhD2
iNy+hjng8dn+GQ9OJNXKsLvvuQpK43kXcrT2y1aICaaFZMeKOwojMfpw3mn+ZIUz
tspoB5r+cDcD/rTzeVd7F15ggP0a4IFPZ5tMHZPxQMOQQ52YDhJ2vwmgmi2h2VO2
y9QLV07x34T+CfbzQJ9tpZBUyICdtk7umLODuv1jV13isySVvfq+fk1FGK0dbr8W
MlBjU7jZpbPhXL/46JVzLTqGNRXbaAtrtNunADGu/L0edKR5gmmDibLBzb+oP10x
vQsXjkPYxknNXOoKbHXMooiR3Yg1PrWtsxWw02N8hIou3RSgURPmywla5QAcIcNm
1fDwvuC7cTMVEhEo4WUG7w==
`protect END_PROTECTED
