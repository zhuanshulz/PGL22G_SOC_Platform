`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hnAK1FUKPM25GNJh8r4ifgVMMyhu6YiZ/4iVrgySAn8SNHnbU9cN4O3R7SViB4xY
bEGpGZNxHAd72csqZasybvuLaANoDM7c5dAk1bqgYXLQ0l0vu4C5nyzcdVyPURvg
sUzb7KBFk6PjQK/i1PngFFAYq6PRiBhYE3JX705bZJouT6VNLfcMqdzvJfJ7g3BK
IA4CRPsp6raqgh2S42bYRnc1XBf3HpAS1UiBYU5W0Yrsgui58z+oY2R6QvT9rIpZ
tE/EAMg6/4N4RBBBAPgy1CjoE5eOoqd/AVFvT7VeGNvHGMT7J3KZalgW3iRvlj0x
FcUn4gW5IqyYYouQwOOvUyyLjF0O1P9jLKaHK+5oxiLXM+hqtvz+RgTr0rQfbYAu
zbgFL9WgMY9wRKPKFE4I6bbelN2LdAwFomCx+FICGwKGAiqRkZlbV3GWqvRjXDm5
NoJwaT3wkt7QBGrqeoVj7QU91vEvm0dTmWr/I8fnsr1zt0t8yi/OCr1uiGAFMQgY
oZTSAvZxmj779p5uQJbcDsEhdXEqtgY34SVOBSig4dl6fPRi1+sq5Ady6Rd7yacw
K9yx5uCN/VUCe8Rv6gBzgydOPKpfJBkkHxraGTkaqwO7LHwxtSaERzhirxuTmCsu
2jdZcoVDk71xSStokHarktOUs1bYVeBrZWKH76sxZ6sZd+Mq1hieoRn+lkikuel7
7oE2OFN6MN9uO1BoHhYXqfHFdo61P0GC1tIgxkxDeKywqk0OPOP4kaHUR19RLZar
jG3jfFfT35dpPkJi55ZtabYUrRi0Hx4SfUNdzjT7UgQ=
`protect END_PROTECTED
