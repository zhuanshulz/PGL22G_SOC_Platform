`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iHklkRmL9AgFkAn8p8Q9dsg/hmiv+Bot3uGOcy4mX1VVbbZesA/dXFCsK6+Ja5Lu
wbyjEct+PTfvSg+Bjb71hIAs4jUsxMu1zbS5PrQ80XnGU5dIfEOHizZkpu3OF+VA
3pr/4IEFimWkThleFCQCoEXImBI71bibq15NIpeZ/v+8zF7Ia8UiCEUEot861TIx
SgDzFi3LE4yyBAl3nV5FrDhnpvGXfC7ZBpxUDtaf2z2hp0bHZTkVhjOYCb5tpr6W
T83yKpZMpkTZvr9H7rx43YaJPpQWxxwPNVwWreK8As12oSFW+Rr5eNd2VK06TwXM
r/7D8Y4znVzI5rDRyKRhgtBtPJMIjl5SW6QIlWao6wBcBqCmTtYUqsVS8Nj1Cg7G
nUDyiXm5yJWthxLP2jZDHGGbCtF7bVvprJD3VA4PBLvqqFBruRyc3nd4goj2lKpZ
gb+R7KgUxN2hJYutq6srWTZFOURUkWQWkrsdK01WpMT8gTkL54enXrVOcHOEejc8
PNPTq7sOk6IPPM+1HQ0k9niUNGGpyuEwwgrox99QhEv+mdHCrMVHWpBazJLRDQSI
+VNnsC5xacct+T+9d+xzJOcKEfznZ/Bu3rb+ooDSPiO/iWaIh/HrMiG/56u8G86K
dINch2tSTzGzFF7s/hzi2Gl8xI8awP00DKp7A9mJjid6kRIUL0U7ZExSYY/1XPR2
jw2OqPaT3BN6ziyah8w85q/5P4nXsKdbZ8RTPFZWfhUYMI5grNNd68xJX9xazxo4
jdKl7+ywj57O6VF3hHIiJL1fXnFrKct933FueE/rV4Gn3LBy29aeBRWFO+vFCxdC
EtsDDU1Jd1hBgpdijg3ARXAVJdyRnAxh3grJmZo8CkwfPju6G/coH+JJ0q5CTcpD
AJwrDM9YnWipWQcn4aShQsIXSVtHr2p8SmCI/G2scqNZvH/1W5OIKOtSINDzU/Dx
VZR41N9QUTXyOlT+6wvPUV+NX79BNIiuO2Z+WjUftRPzg4bUmJKhrKys+3J6C8PN
lREeXv/9PLOgAnaQLIqTaQruTCFIttSuGu7SAW3RMho=
`protect END_PROTECTED
