`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SKDvkkQGFOMbsgOuhkNZCLJX8ZgSzcJxf6lEmIpFcrvDVwQWv51RpVFoNAGH9L6
vaH50km60SewMSIdLTsVM3xQpc+m4ICi5KvMmyJ97I0oqZibGJ56ki8ISno9BG3E
fTaz4Xfr6g3UOENqGFkgEVDUOnUzdwwSrpaZUInMbppqQIHY/yrlzrHLDN9NOVm/
uH4H7iGZgvknPQd5jP+XMzVI4/FVRW3BdCq/XmT2Z2fDS/y8UgAefITYHNE5TzYH
ZXxt01+bHOJ90+aE3twHtZJbTbhXU5zF/cDNSne51C4TnmzpJXqD0/amPBSkeJ0Q
EEGjVH7SNJQHJ6r20vHK2Q8RKFz41I5GgShzPJJQ43wfztCb4j/CcCWby+4KRGdK
QdcikxYERYHBCacanOXVfnnm9D0yn0CAJuf/gsKfp1vsdBYAJyduW7nxtTtlErRN
jZ0wVWEzSZTCnNMdubm/Il6TwQ6R4TM65IfufLIyTKFNJj2eiAOYOjyhqdEinVPA
P6ig3PeV8sxLEiyyCywmqEGv0L0m17A4w7UwI3he4xlw+2UxM8cVNFKvf8Vq76eZ
hdDaz4Wl6ZZaLkDSCEjGDSCh1DF9jDNFH6qew3TEzBe+PqtrerYigVT4cXDJDB2k
E0XF080ggWGyw2gjTUL1LeCcVHas0tcDknjAwNhEG6KDs+EYembIUa7j13tZw/l8
xi4x5/wPsLv3/jxUYvCGgYSTPp+eOq3FnB0zSSMtLM5YKgoMNxLbQnBtS2GspR2L
vvYb7jy5LLf2HuX4RqLZLHD2JVaYhmWhFOJ6lQfLcf1xwXI6y4VXpkQmtZLHWpB0
`protect END_PROTECTED
