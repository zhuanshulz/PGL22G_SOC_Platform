`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/u++l1+p1Nn7vsDvxxPP5Wxv/AM86UsXwfHJjQr7Srt811fNeTV+t2r8hbXWRkcn
+U9AjDr2xATlK+kcPTrMOUT6hzQwMj/AjBs8Rdxmf3ZI7rrOzFqDP9RmFKa5w3kf
T+3L41x2FAJmSAajpYYQJEKnsHtk1wZtWJmMIGmiFZpEVd+wejiueB2pHbWmZhM4
iH3AeRJ3i7jo5on0O8EZjcP8OuB8yy5VbejJcbH6OuoBGndewMjyD9jnGVyqaAc+
/SzvmbfxRln14WJHOQnLFRG/bVG+f2vMVz8roCBEwIynlxvAvPm5LmA1fsuRFNew
ItCrmR1gjN6QN8HejLPrVz190mnD1ZeGNvk37930kKR251gTMcNYf44tqO5H7cqZ
IqRsJvotC/HqttS7W+72gk5X6A6NZH54d5zUQ++3+n/JPGVflVymkoj8WF1LWZ4U
XIO5oTbhfZM+x9HdGG1UwL5bCoIXX0ArzD4UlLyxSsI22G06tcWncwDSPmfsMVkJ
oaJEcyuUNm7LRqkRq6itm91RqPTms/CqhZBb8Cx6HhS4Wf8VMxUk5ZXQsWRNyyhl
8nyTZi0Cr39AYGx/tUB/rvbGsJd2CreaxXD7sWV6DdGI1TINy3oFnFSXJOzz8r5m
lw1tj1SZQ0KtqgD9o2eJE+ZHwVTQ5M3ecWafnBQ4t34BWcmDQI1xk0a5582o6uIC
2RqMiD/bBdmXOebDoFgi5joeAadW337lOKtXDmYW9HjdbyXo9ArD17RxYq/mSVwn
eALXLmx0E/lQ+VS2i53LGYZEWIUkIP9AAUneZw9p+iM=
`protect END_PROTECTED
