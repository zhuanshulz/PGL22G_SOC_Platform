`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Wg0iQOnypOdfWxHjiXxZ+JhoC+OdxygleSpteCfIB9prNl85U6xRCHOFMa8Tgz1
BfFAdGdWebc5ifsct1CSfsW7+YQ+rQL70MAKmZLm/rIqb1EstkTfP7ajr/RU/WBy
0usGFfhfaXyQ1cShaOQ0yW90G311wL1eTgvNI7HTjCyYT+JJPYJcEssPjntn6QP5
667UAcsw/PVvNLgPcwoRs+UWNxKYy8jES41LuVkIeAHuD7Q6kIDqEOFA5q92NdDZ
h44pL8Fr6bpOM4Kcj3OVnMwqOJZhwWCUTP+aN+0v7OLGeAOkBi4BRVQZovHZR6l+
M2upm2QmFf2pYyLVbKJXHR3sWgX6cC2D/5lWnf4fJwQ=
`protect END_PROTECTED
