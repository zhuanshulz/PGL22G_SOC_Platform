`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jLu0QE0GBLay3LpJJfuVzRubeWnrtrnQqPq0AywP2NOC0BLEZT6HB3V0o25jqr/
1rUj/ibxh3/ZEMst0pCoj8flRw+8jclRoyfuxAMgezwytFo4wAAOT2+4S0OK+MwO
eT3wwsS2L9bGWRPbv7iGVAImSC35vfFnF1VOeqsZeYjpmRPnqCdL4ZrF21sXfskf
nj85Y2/fCUCa8fImeTzPMmPDaKe+1L2CcgAFw6qcuCws6fvsrd68g9yl568fQkkB
8WHmkk1/c9qktcrvpmPwZTRa+p6CqIMbc8pT8bBbTMQYD8Y+NjO1APNOkalt2iLt
lSf8c5CSM8GAb0UVbGgdGq0o9cDjeY1t5UsxfNPLlDSBZvCRLObQCG7A7m8uglfg
dJK8kX3BE+/UwQjwGqTp3dDwgQ6L8ncYioDRjRHUiQWAAIdRGKgg2eIDMBbScoLI
efxwu+Zv2paDsMX3nMp92AUpzJnaSt7cICut8LjUDYDIrYdUnq8B8IXznlQRQqQR
p+wdrtSgY/e04G8/WG+XAwuolnzLW9qF9BSLWjFnF3Rc6YeKtKsWioJnx63lS9EC
OLg9usvToPCo86dOVjJf4YIC4Rkqe3lw8W8Wpg9K0qQuGv4G+sg9aKQ/O6rc80Ly
yPvnGukcWX4XmcY2Bk2VzJY/tCQpGMs/z98ilI5yfKl/lI5HtCvgpE/f20hINYAb
BSKDi+GiwBYbgth09mqpoTI0jMiO5/Cb9y9VOd4XdJfcXDTp4HfWAF8Eg+oUvz/F
1f3zIUFMuZtOrpBhIbl4OQd2FwZ3s9fsQ6uadQUHLkXaHTWC6Qg2W2+X/a9vVgP1
/C1LIkZBCH1P1hm9n9u/Qfg3T+A+dcznd2mHnhClVyELlWNsVGjjpTfoI8aCA7bB
gFFYOTyAmZs9OoNcEszsWzFgpHHol8ROVyuKMyG6DAYNwWMW9gFfjMqbQMAlM93U
6TYT0chSHL/37UCZnHjk6FUOaLedanS4YP5JeBe/8Iisa6FRf9WvcBNrVpQZ6heK
gE49O5fBc8AGsaKL2BneWGRf2b7jgho/kyPMyCM22wzJRjiPfk5MAr8mfJDPRLcD
m92kWEquYj8sLrJ/wdsJ/QvjQBnzHQG4VE9spAZwB4QO9iOcjo9lWSbnf30FrcZX
qbgv33502SRLsybkEv+rv++1SyB1SX+od7Z/BVLeQGFrVnWSu28JIX2iWAkKUbcY
OFeCo5HjF1zU0ytfEwvYAq1iIvwLnAhFJ1m/ju/5KcPxeZn+iGbzH6L9qHUAJLAz
FA3zOl/l9H50ZdcASt14HkHbHgeJTCtb0iqHfMiaOY4L5KZ+jTXOId/YCmQPMUXp
uMYR5v8acz0dRUnyRnhp/wg7aQSASSXEoMzcLVV3r2Y1CkkdVC73Pf755OVH9aJy
zSuaxQdvCEkgCrizIzD/mUBCLBCGNptBD0Lfyi9RU3UATkz47FEuy0r956yLxljj
Ki08zkahuQ6w40AYQTXgW58Sh9/QOxrjkU7yvFl17ZC7z9Iet3od0Keba/NyQMtN
+XCGtGtZoi2fAnm7XPQHFng7VHamLIJ1EENasDUPbV2Prl7/7hQ8yc0CXmCVfl8f
X5a/2O8kxUw6HGATV16gmg+nEapVYFoTRrUWI8bjEaraTgRLLBPLzJdjo/BPXNyd
7v1ZcbWetk7wCkXhqNNyqFArJk19V/424AtYHfsvXPQOCjfsOG5QYVPbmka4lrh7
onkGaI1pNBAuL1tgoiLoRIt+o/kRRB7Ogcbrr9XfdHuQb37J15Vi9hgMyG4owou/
YTdZOK08YbpQnUeI8Iae/DOOTHElmJ9876iWQIpJdE+3sG8ZZP+J5JfBTSnxiQtR
QVxwICQcr45Z/ZkR0lfLnoN5QRcYk0jTIXirAskbI99BgNZabcTB39jmSpWSVQ/S
qpFb8t9CuxP3l3ugxeQxg14hdVO7Ua55vJO4+12Wa1ASEbgRgf5+IqYcxeCuNdOD
g0guUajG5mG4k001DMBSGZVLqqaAjaqrwVYrn+1Eu1oUf1kDlQ7m/2Bjp2KE9rPP
BwEUWehFoPDrR0rYwd0b85Dis5vjl9t0ZSyO7vML/iSWb3Z5in8yuST9EtauDjso
Xlmobe5co7crUZTuh9UEbvF28X98SZq+WnkokL5Iu4z7yLxhIuWZ1S0EOd3FxUOb
4BMAxPeTYhwk0FYbDxQl9mdNzpx1TdZaX15ySqO0t03ELxoIVUn9g2ulzzN2wXtO
xfPo7Y8pXaUjeqCf+QHH/AaIVda8NKCIIlKTT7DPvr5y3Dc4aDhvGNy+m5mcFo9c
8KV7NJdK4EhmaHUW9qCeKOeHLT1kPkBOJ4xDEHCzQWxroEJRdK+AaZppL41JNq1B
rAYzNiZT0QgxuQXyEyMmRjLSrmUeB3IfUg5dtQ5EY+HBoWb0/pEB91y2ekm6BfB1
CN0YNClLZxzeB/XIWLft/anLlw7ekDL3ca+TQ2Kv6UlHq83cf27Bxdapa28uVgRJ
6+t1/sQytwa4cHiyjuN3/xa9xcgtp+xsWfewy05LOdyaJBJkicGODQvatXTJPs19
upLzZGRKSQgGtt06hzjKZ42Wmj+0cTVWMmPJ6/pRZ4IEIW1yX/DvmXara61mtMyK
RoqgQSCupZjPyukVzwudAVk7xRUnxoGkZTcZoV/K+A8=
`protect END_PROTECTED
