`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asAyM5DbmetrHqY9KSQ8DwBYI+JSEpHYPBm5YO6EReguooB590v0MakBmuQiooiI
A/SegTi+/TfmuJEdSa4LA5INTD3j5ej/+qw6oQ4/ileuT83l3WhbzmmKObTDMaRl
bYMaQaU98p0EvRHVD7K4/q9tmLx930VEb8aiHyMbcPdyfYf1tlw7ct57TQeahE0Y
NCikxzaLUo9GGoZrkrtl7e4/6f6MQg7tvKmBogW2e9aBVzWzzDfBvreEmmQOconT
b8kFtzluhR9OtbARfj3JuMVWxUE+M322+zDbPxo9rfaYWw4FUJf2mCnPvvRR0kCW
pVkXwnvUpcCP3RiGbHF5r2GSSBWBxmQTEybDZZG9BzdM6BLDtOvw9e5vTyQ9eHBh
C5Dd0RYt3F53KaEX9zFb4sgGTmv/x+JaWsvyEPJaxDjPtlqGQWHDxlJ+EHdSJJek
4l89Wo5vxXMIPIeTQcN1MFh4jaNemN0AD/go/i1/VltW7oFPzeRqrxdDVd4RklJf
YRnQhxoZrxEdGVLZWk3tPejIvIpcoV6PJBg40t0PaDOrCwRId4b6o8CJkqxuOXOW
jlMwlAANl92W535OGv2Z3GOW30xvIRiVnHZSI3mdPBAMYeJYwHA2BVYpiODOzT9q
44/9n+12Jw/JMTs2hXfPcbtRgWW2+sIsDT0kjIA9GI8GJKmreTzP/z+4oUGFCFaf
zSsGpRcFbFaej/tl6bbBS4Pn+99NYtcuIVbiDUT51Qrk7lAiluzesrssnoPlS/d1
hZqSCdruACHHTK5FRh0BuNixUXi86rPy8DWVM5hZdJscqw/vfRrPIGvJNl2m3UcB
TBW4Qcgmw8sw4aIsvPrM7Pl+Eca5DQ+5TqC24zngMg3HeNhQPHvCmFJ0ka+rmq7A
aVCG0/8NIyOhn78TXy0+VrGQUWIlKpc6VrtEA4o9piajF6DYo6hNZJHkBu6mkXpb
bq36+a8PN1VncDFpZVemCglZonr19MqCtuLJSU7amUArFCnUyMO910t9NelfEYyw
wVRD9WWZUNhRBTCr1btGi/hW5/AnjPmvflq9xt+qTa94UHbSlczITZLRn/Vqw+ku
Cl53jKlnaPaWrsHJ6U6IC7QLUvse2vctgOTI+TklpFGjn83BwH56RRaDaxgF21rP
TaLYcbfc+Ur2oagsHc9sIJRzU+GyDMVQ9DbCI753JguE68aQwNYlYPyjqXvglk3Y
N1i3JAe27/rgIFg3Dv/KPHdwDWfuATPgDcYJBDXWUqNl5DN2midM4K92Ip3rmktT
1b6DBTciS4QL1aJctXo41CKF37ZHXsSDoGsz1/G0QGN7nVTCcdxyCWe0V3Moh50Z
WeoHusrrYIFvPGEAIDEJabzHVWYoV3nk9ESkIec6Nl9m1svvUNDIsG72Se4jp3EP
OhagSP9Jl1QFgYnE8AOGD7y17PbPUowr63iY4zAAkzwXx5GWQVg2S8HMWRIbAuzc
A0JXyzFE/wsYbMHS7u+syw/E/+BDhBkX/IWCp0IgjPtxspctdcsscoLnh7C8yn+z
cb3dVETRvhIfJcK7RR0FQt4SCFJY7HEp/drsovAaUXd40G3r4I7xqgbxslvzZe+r
QELrUH8ME41uXeH1W6qc+KQtOOzwiAYd1ylWkPSXupWL2150zL8JASU1o0rO6+HM
eHoqWsrBh36b6Wo+fN9a1TqR3TORWLv5byKsMZYtLnJlV4BjIfb+SfLjW0TA+7Dv
H6Gdf5IWG/HXpneCmuuvT32C6AamEX/P3Y/zjylaGoRdJpmP/0W08xvBWnxpWkkR
TiLF4vO32DQpMZz6g1dA1uUAARWCUpv9eDEU7a7Ad2Qlrgjes9Ca/VLyAVKXW/BH
3xsjeagj3hEf3fiMuafV0srNpEa20+Qd0+Ldkp/IShLPdFNX97sRheFhn8g190DH
BpRauElAcAbQxfOVfGOFANqOOlaEgY4UuGYtHdJ/5r2muOtFDa329IsDKb+Ti68h
Ehm4PZFmBM4IbwtBM0xXcQ==
`protect END_PROTECTED
