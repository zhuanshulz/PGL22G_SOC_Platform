`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b//ikblcslQvD4ciEblon+Rqjz0nwOhal3ZOxNpY/+I5GTG0pRLmN1JwaLnLMwgD
/4sCcVbCC4Npf0LvS6v8hzUK9pQvvUWp+0qV2WeW1nfkKb12yKaddxnB4tVB7jJk
hqwqk5CbQW1rbLp0HQU2H6Heckad2UpxxsNyjnA72ABh2VmBvvi+oUfOGknKsHOq
Zw+Qn0ZBpyRwfhHzphL7fCbE05a47FPGZ8CW+I8XiuoKdVmbk0nzf3gNRQ52baWe
PT/65AJqER8xxDvqRR2pHfiTiVlTEDO/LjWXetRr7lZjn5lTdFCEqRSkDPFFYGnl
NMj/QuIspvxErHcenOYr0UWrS50m6tRAavZlC/IFi9lWg893tU7CUT8lwv6JGDim
UoSmrssBMIpPpkf0I0IcfETt96l8ds8zQwUu6zx3ixKy0F5dko+MZdH8AMEHCZR6
e8aoKVZdSasj2zEzGKAMljfqH8ZPk5qiKVEjKPhR7pZ51ByTo41rnWCXPUILQyrX
R+w3wzPO4OsENIQmkFcdBP3ltJc0R4I/Qxe3BowFOFTB2TCQC1DzsAKSHnemEtee
7FBHHXNSzNzFiejets98skt805qbrXMhrfNiMHyWcjjhd4DTDgPOPIDQQ8FxAUf4
`protect END_PROTECTED
