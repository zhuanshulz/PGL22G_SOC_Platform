`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
COvf6bRdV/Y5N+fydGT3jB/q9EyS4eiKg7/e/PG19dKDJixWtFlTxKMbh1tWBuiQ
0nk0U2IgGEcNzlBzP9MU8cJh2t0q/o5ETVk11+kMP9E7/0xnWC7yqb2nNULod0Ju
gKrA1Lak9oEmuDudO5n8P1xWA/Z7UdabnER+HP96X2/BNF1tqDQSY1hVS/UJvzHV
/UvVNzQErVar3zGcHrivBJFBPc2Z0ZlRAFqrHTQeFWu4NaTnm5nJGYnplSdUZKbU
cWDJeNcF36KxPxP7lOGFYq/peBVfBJhl6/El2Udm+GG3nZpQwP3cVemHlCeb2Px0
qRQ/Y8YzYH7pkxMLR7hjS56AwkkwDtapsk/pp7Vmpgyq0bwPqDgZwFAVuB18tvl+
XPlq1tnMFsfl7hteSl/ARmmqDQupG7IerQHNTHV3DPs6CM5d7tc6CCW/SRQSmPai
kvkdMwW9lffHP6AZEGCMxBTyTcYkSBmo+7tlZh8RqaNmCChZsAfhqj7RsuKQMHtn
sB8fkR9fRwhGu8CVzVjKX8ceJugNBG0Dp8FzoaJlfVwWxkiUgWkKJifVr6kzprk0
2Y2t4Cj2tsbYLbUU/Qn4gTZ6YHjvYrnhHxZ9/tsBMyB1lk6IYN5BdnHKwvKbWYPM
TAazFiCwV49DusKVAwqdLRKXXXkI5JNjGAf6WTzwKl67qEWJs0qzZcen7EW7UGNA
ORsEkfMU7qZZFXEpURaGqmdviBz5La9hkhHf0Y9HJIOOPR+B5MO9Cbzz0LQpexXO
4HqdEYrLhD9rFCzsj5STAHrhajcR1a0LSnRAjfm65Yk=
`protect END_PROTECTED
