`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
86q1cWfc5ArUBwOAJFisdnkP/rJ1JYvGgXmudlHOWkN2tEL8LIEYFFskhvGUdCYv
vc5PqHfXIMLeApW2wsACkumvKd0HejZJ9VeiIjp2uvbqa/vThreRixalGckb7MZF
TerUQwEzy9yS0Hc8Pt0c+Jhxo3kY7kbwHrbTUIXxHfxz0MWjaRnHcXAdtP4VS/0G
2RelDUt3gCxcAaa75W7Vf7tdE7E9RfMw38ugQkkACeTidP7pgiqyIAOhSLXT7xQr
1MHKPBw/baQ77jBRjG7satz08qzTUdrrOE9MHnyChZTxryt1BWVus5tFG9WU77Nq
gT+2ANsGvacmF03ZmYeX8vZ72w8YQNbCcHh7t47zOfjLKO9U49Gl18hUMxwIZCHX
nFzPPu3/poseoiNojfo1uxgnWAip0b5/p8jZmDvPO4k=
`protect END_PROTECTED
