`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RoHITudqtcHUoflxulwiOn/9VR72eU+0V/vj4xx29bJpBwut5oe+rdR/1usCrwuR
HIpPoFCCdoS0dvT18nehW/ETpCLlvdWFu5tgiF7jT2pI0FRKoZlW7CT8FMm41JXj
XBQ5B84DwoN61QtvhS8E55R0vdk6nhRQ/kcw7ZpGxcJNKJ/lNO6BBFGPfbh3t8TN
HUDW9rpo93efeqAsztwPCh8orqVLneAsrc79OjvLOASUT14+HtnRY+4Xks0WoXRd
OU1wU5TP9qAXD4JDejOM8QLu7rUh/bJqPS3xhEc7KOtz2FfEb3E1KdmPZAfK8EAq
DhisfKii4HrH3wlzXL//cGPZcvaeiQcb7M/d+gFvRjCR8UEqb8dv+wZJOj3tBaA7
e6Nc5gnkb34co8sKfkXe7AW4b8dac+M3wAZaEWKIeofLycMJhKGIBj/pf1piAnsD
zgrshycKerF2mnzzeOy1S//JOvARn08ZRqHYU/nX8z/ygPiVPF2oafv2owCwb2gJ
9wV3K+3GZgtGK+4slBZRlHMzJf/kJUh9Vk0o3g9cdbQCr0cfH7NsEZJQvD8nQY//
w/VgHqrF0/DrXON0EPD6S60+yv5ZX/kuNUpsWgaQktAqXR3KlM08rhYWOeV2j2v/
BpoVs4i9iu/qRo/G5FA9/DMBe2805zHNOf06CDXMo57zDc0J+vKHyDITBb7vgL2R
T4uzBLQfTh60DqvDml+RTtVqYON9Cy+o1aWP9vuPQnQXOTKgl876QCjSLxu4FazR
NjYRIQB2DDjtG2LwDtIjRxj4FkSo3zIfg510hhKH3KbkkC/l7yZAPE+epx1UcGWX
ozgSF0AWdTu7GKsIVzqA3VPixoHRtywlPoPrGVZFi3rsmcxGUPeU6YmKp0wmwaUV
WumJJfzVS9clul5Ob3EmbdH3WMGvWQ1uaDkYXn/HeXACfxUbTmzokAEo0ADSnu/H
9Y+eciIrKUgBmzqQgMeO30tkf5pnQ0IFJx8hOeiLuQigGoxjEVYejJUMUA5Ba/eY
sOaGZVjKKiq5qcCOcCZZUNgpHJr/PCDUJ0pli5JwHlpnTgGgAL/1GH3Pj3bTpv9A
4cfRlEIrK9v22qErCBwdLzQCI71Jl5ZsroY/19I1VbVeWznV3PQSUSsg6UYjrgvS
merge7RjLq9YSxztENoMVKiiCn42vzqb3LbjVcsfY3UzlItHxrN5a6NelAbAzr6F
OpU8Fhj0GsJiZ92j29b+Ks8yG6wPAeMKyW1jT32Y+eDA58jBFzTrSCfBxV/cHp2Q
/8yGHpIwSpCNBW0tU7tESWwbYqBt9Jxq6gQp+3eVkeVGAbmm5AojbhBdZekaMhRD
etlblmk4PqbEnVqL6TnAVy/s/lUqOFdxV8e7SKUoc8VG5mDoNTDKR3ggnE5FiwuJ
/5pk3cf0UKZ/MnC9gE4cFP7hg3ILrr/eDMWpidzcl/5jKe+taR8nwMpetLLQp507
GyxxNE3ndLTp1BOUotnpAhq3tsWRe93EEqLGPXo8c6f6pt8xAZ2kVriKGCLi7ocR
Bpi4e+SuNAsGGuv++JQwZQ0BRPK8/OOm/O/8gSNkcPN5lFZhqIUyWKbofMxHHzXT
KcAttMGYnO10evM1hNvp1lBWpuzvuM8DQpsnsEr25PecrlIYrTrJ9KXbbQtKbrSf
Oqp+ONKt7I2N7mO6CiQjNoea8BqaABUJK45Z5oqsBDH+piQj/h/Td/6CeoYGekQQ
Vi1TZjQSJbj1OeSu9+imShWb89hqZrVXB6JNcyAe8qny8PZCDc4Qg/VvMbj3RRtH
b16/o0Qk6kLXusWJdRwLNr2bpzeY5fNcfdKPxx5UagF2bl7fMjUUlwaGaDqfXp61
6ZcWkMmMEC/96CbOjX+E1m3sBcNiqEsrUhI5OqRM2ZX73zMDZWZjxmYa2ieghIlj
sCICD1Hg5Vom9gD9W8mABIdxNiM2PgBHu1C+2MSweN539JUeDhdGlPW8EfrdoYNk
IKNs3d4fiQuALqOjIN5hoUDV2vb3HU6ILQBJkaJ4122/PPD02XfcQY5XXA1DAEmD
EcAf4664GBp1tgsc1limawld00/RYukHPr9sfOgW9N9VRIgQkVGK3PTl6yW6EQks
L8p8k8nrASjqZy7PyEx37eeNkRQZ8zX+xdK9IaEMA6pFQ4XybmnZH0KZ2aIuv0bm
TA/OcExYtNlA9x5hBPMM+cEJT+AI3SPPjTuDmrY4nYpa7qVGat1vptT8J5AM4RqV
wKH8wLavMJc8TDtm6sOGif0EAYt8I696PbzkmP7288NuyL0R0UwFUejI2AFZga4Y
BSJO5pLiL88mhtA6aF92Di7RPhw/P7i/GKgHP2mpoCoAkI7uZXus6e7Bz3jeVk0b
7cWCfFSRwaZ1vr5ICfVWB0HKQFE4gxSLmwg81kDx+5BgjOkM+UcO792oPxvVSd1S
8ksfQpXG3zF1HWHgNCsVM/XJe4H6h7bnygkjTdMM5pavqJz1GHUWOhbq3TgC/f6S
PmDOWPXApgNCz1lvpdc6gvJsz7AaXACGvBu9zJGDmaxjc1JTOC0b1HxXsYA6DnC4
EE2LH+buTxXwnQv9HeBr4oZkYXY74T480AN52jiVytj6bNoiVMA+/bd+EwtMToGZ
f2yS5RxUcl5YBaNqHcOVeksUzydPAAQlfTIc5XGYzPmyeBuTYzusJzsX/tbdcQxS
lu9lHschF4bBh5Gvgj2UqqeUEzMJ5Nbhl2ZBUmwpLproIeINODTPyZissUdBYL+b
O5Qqits5L4IYheV/86Fd3tef+nFCqZ1WsRHFb5fgpowA+STZeSSs2XE6JGFv+Ye4
JgF4UBvWlF/PlhIddviTiH810gGmLeivaVX/RDl9unB4i0Q9slS7Y1EMvjdSF8As
5VzUQiobzOAz1+3/HW8ivuh6hI+fg0vCMuvFjTdv65EUCmvR9vLAtpdlL/6edlTu
3GYqW7nMeuyZ7oSmYj7I95EFCB/Ih622LO84+oyr1KF6WZ+Fe/bny3MUAQIujCZB
2NryZSHea+owuyu99TOvox6XrJl6HkxZuolaDDLVZEff25ozru9Wnk565FUyd6nY
flnrmntPz1FWu4Q68nz4sr1dNeEClRoHzoFsdYbzLUAmpe7+DB5xj78fqmz/nJjw
UNkhQa3GvSW3nivbKpvhbPwPUm+NBBzx1HTy9h4BZvn8Na2lyRXEPtNMgJi8rvO8
ucuC2ldnsC+Hb5Cn4phI6D0kGTm0dz5rcjVCG+YwU2uZlqVGyKzgCDUVY/rPfr4z
/UW9hogEH72ZiGTADex6K2cl0FH/ddF5b3200zgZfGbb2VivBOdrqYMkyrP9I2Gj
Svoxxw85bwk7kpfMTKMv1QrYbmftfre7f9noVBhddxh+0B9+OP3+dyx7zqjbsVnp
ucjswTsoNUbGYJpn/p3/6mp05wdXcTEuITOgWfJTNfArOe8Bez10jpXLPM6Uw9KN
2OrDPuZqkBwrHzuDEVGKZlNVqMY87i52WHFXy/AT5IleIc3DJzAgcsy4Fb7s+Lhk
bVKEZ86RtxYgHRZVqSQTAb4usW6415olw4+W99v7w8wEtAlSUEGybw1yB3LTTnNp
cRXLpcG1K1KbJI2Yu5Mpm51C90YJCIEg/eFyqYI9CKuvleBbcKIA0aMdMD99QVS3
ISSnXg+iLj9z18XL3gxd4yoaoqgFyQHgUqNfCGShaPkID4qyWbODjgjyWiheGb2o
HwLXJUPl1MbywPWujk4WSTv4TFeBayivZ7HlM/gnlo+BQ4zmPkzFTCtCaFKGjkFL
J3IWqUGMkC9Cuvj/bURZtX0iSl+yRHfbEiVEccLSuH41WiZbqRdoeyNNUprG0lDF
V4NBANoXjdXltbdmE9E5+Bs2WPyYA2SYOcWGx1UPmoTQQKBjNCqHkQbi4qVz7dSr
3dkCXLpL0WOzzG16D33dRYEfg6eyv8HRBzSOuYuUg9WeePu2neU9l9lNySyFzgtJ
IDM3he5oAe7rZYL028KWpzGJEaanvbLj62M+EGNDM1NZiLz9tmAOIVdzUcuUVVfn
/Deg1ii615zrdVbGR5y+U5bg4ccn0UVKxkvgKMpfYcJqzOJXjTg6hDDPXDs2JaGn
gFOKVU0amlTxG8bGHBCw2i1ZDKOUc9kKEtYUq9LQJZQ9CCQnqxlMG3FiD4xSCyp4
6iNYveNa5cBgFFQOnn33KnbIKj3UpSFODTdnsMcQxCZgTs8sZz87veZULA7RYszM
mg+s+sEy0VjjxK9+GshxjyxQDtWYRGO9p5ffzZfUgwdXXVrSrWVJKOGSJae5xZ2x
UKLK4siYbqowzxJoALWYbpYQwcAu/E+7fXpGsCY/QUWInjN8nDt3D/UslRsc6liF
/AKOQTXvk1B6Mg/V09s6rCuXOJ3yM0XA0zghQK2S9Am8atOnK1Bq3SImy1xxEIem
zUFhTfYV1LuEDSa0ca0aTZ1k5YqeRx1/nby9KzvSoczypJRHEWfk549z9YxHaYl6
KaS4cQa/5KuQTsyKTUINmrSB+38wFLGlT78ejE2uyssMa/4u4TeLsxPYwgkMYps3
1dz32fBh5ozBl1j/iQWi44ijvdaqSULzm/lmIc4HEeWn4MFI6nGXeB+ElX21/Kj9
4eK10b/cWXk2rXm5Z9oT1wvE8Cc0dGAbfYrf0NcRwiZZcGfX+acKGeIg8K6uomN9
c3E6R5nahyX4W+B/jsZlC6BUf+JhMFkEvpx+JDS+SjzB+vUz4tI2wYeEjyYJ45CG
oU6cBtIAaXMoz+OodN1mqiZxAkF3fKQrNmSEhW60sJU20avY7ekmKBxv2xt4yk0F
VmPqqjgFK3fH9h6cgTeMf6UUplaYXQEL/1Mps4FSCb+gDgHsiR+zg4cZvm/clIbi
tEPNju+f47X3lKv4vhBMMnSg1lmgiRTYEIKM7J3EZhO8j5DC3p62Gyj+IPSBVS/P
KC7+dHNveEvdKRHXMLsdJLwOhDAtU5jR2FoxI3j3jopizY5VSYOtf46SIYLyXhrS
0UxgEVQ5iIxxIJIhLkpDVBbY0TzcRgxJpiavJemCkjtRS8mLQREv9z6XCCnUeWqV
C+YQPU5KUK9DxID90PanOmfIB8biJiUiezi1cBwlt84bg6ieyRJ3YYyVeJCXisKe
LXguUSGC7SfEyc+547FsDvVJVwR7hXKxRXa5jO+Zbt0zcjVrfGC/JinCkToSU8Kw
FiErk7cQZGhlsScBqmr3UUuu8a1HkKXf3fNxPnZP1AXEHELG4+p5qcTe0C4AXQX6
g3dPViL7Eg/dii57HxdQSJXlO4dwOVW8j/vglkYWI/r8cxXryOhiko/l0NHoj5lz
HmaaDuRCrAm17JLySaNGBma4gJDkxUznehJGFK3IJOwcxJwtyn9uPpsJO/PgB47+
sjMpUlHL0Qa/Q53VudF46WZ4ahcxCBcMW6f/XtQGNKVlmm3n6LM9HeUUn3wos+ny
9wZ0WsEmOX++R1BnMCg6fJhk82PxO8jb2wz0/G6HOSCYJbk/dpHAyJriBpgJZxFS
+LC7NGiG9omd5fXJC6e5bH6s0nGSI7M+PMGEocmGj9UbR7SAaKsMV7D2EIl25obB
JWGwUHWWX61qIEthkhRRKKKQj5qVfMK6mGW2aUwrGdk/NauRNrImy+C/66soUFfr
GCFuTeGfC3FVUs5zO/NaJSyJjGE3sjj8KjF07G8PT8gwjH0ZotHZ9iDGtuu9FOUD
sRe9S0DreYGeigb3unvME3NNAZHDgsh/BFNf+3fUevg1Z/qiQbj4OmMJNDUQa5q0
IbpH1ppguJCP8cOOhi5SzCMFwTafeslqIPJ1oDd2cB4hP7Hg0+bqDShw0L9hPuB5
6RuC/LJ0sA2OgK4HN8vmVBsHQlMC+lfxBpmaHteAVdISJscswjXwBeBd7DlXZ60B
KcAvLkPJmagdMRALwNLsrTCUKm0+bGz893yC+GTcIZbTuUrWdlTSLCatqYnbVW3p
8VZ3G3ohpl8yXBoTdZMN9eVDr9NRK4Wvx2YyuedHpMMBukdurVbYQgU9YgwYpnmk
Ze7oDsrtLKCzC11JR1GcQAJ6uT4WqlS2lNM36fli5GL1ReojcPBhAVIaW66SlKzp
doPdOVqLXEO8bbaQDUgQVdOqGjPm9zPAdEiBHBGvw8XO7UbZxcfQhw+jMN8Ffrby
SwS+vEd9qRDS+8Fdmlst6goNfZ+KpnbHU2qPR0hCJS7K7d92m3DVDctUBrKWEfyG
9WUqZjXqihzrrRB8RdMSeJwSxs12SIo8Y7gbbHC2se61hck7xfG2EHnQqEkzSiCS
AIQKW31nOzwDvZ/Y72cBEZGaIyIs3yJZpm43scILyr4w42ce75pOYBfEVvWzndJ8
tUEI0IfkWFMRzbveXw59c+ai/KUh2DOry1eldUhUBjy6dVjMZ7sY4TaNso3jhxl3
LCWDrPzFBZgRVlV2tNUP4ZV+QOKoqlfj0WeIK4gZxyDPk2UlVYF/ILvtsUrsmPkm
mTu2h2YhTHlOwf5p5aLApTl+Wt98SV+A8x+GK/2nf08qHLH6EExgQij2f4d8bN+v
xuW088HBr8GcSc4bLlUJs2GqiYRqkrKt1poy0Y50Z9+vEHHjK0YnUhSpHRmUDJP6
XKsYj+XiHG8kzkVJxUYYhhbrtOXsl8xxd7ph5FsRZxDT/ApedeZ75baypaLReaSm
i9YaaN1JFQA6/sRs4S/Ff5DPyGSCj+O/F7flljr8Jtj3MXC1QbUqAkdorf+4DPrU
xHzfKGNGEZz0oHwYOTyociNVzZ+Ss7hM7o2+TLsE4xW/It5G/vGdYRnObNRDyBQF
yPqCXe504LauVX2ttMSVlr9IQRBzgUWL3mW8GU/qiyo4+qE/m2D00VJZUzgfwczS
g+1eXH23ioJW26EYzbR1S5a8dgU1fsc0M328KePO/vWNe+WCV7Rj7MEpCwtgnf9p
T891yz41UcKg+PGDUmKoDxIfXqigYA6HADV2qurr3z/U/Mv2/8htwHdnKJ3fh1ES
OxX+4L2IsqhwjtuaYgHJXxxmTlOWxxwWlbxD1pHVXnosX8BbIGnVRJDFkMIbPQZm
HynvhEf9P952FOVZtRwgKPx1TuLOVmcj5+xTCkSFVUXwb1/SLrZ13XeNRu/LuqFr
1+XrO4leI4T/eUdSn5KWhnRmHoAyxDY1AEc26mRXfAFbHrBUCwW+0lv1jcGinBZa
hv/3riJAKS3UN4N6cYCzfhcwdbHGej2dFTzkbo0kO+EiSz6tHk7g4xA8qja+WYpY
X63BTyMCBxI+yyEY/6dYxE14yE6eRQnxmvBQC9CGf+ZRdZW8IkGzNzZmtoTwsWL0
N/kugV+jQ60XBJXl/BKVQdjMpGQ20KqYtAuFevBFIDDoGABikgid1K5jGkhGfx/k
4q7sx4Msbm82uM5Faa91GjvSqrS7od8GB9hzGPMgElI0EqwHmSPf7lB8AlYXe/t7
JEeWyoR0TA6zfAz4mdpu49JJlLPVh9mzUR1j05vJ9BmaFtZYwwvF8hJW+ZGwMmsD
USOqT1rrGPlnWFjRehiEN7wxznslDj3bbEV3E2SNGHeXHhS2Vt+eqPfBNUbRk5I2
R+sTTDjXYEaKik1TDUnXmr87I2Wi2gnY19HiQgCePW40hJ6I78J+LfuvFtPnjcFD
A89lijVHhP8vlPGIGvorTw==
`protect END_PROTECTED
