`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kalfiu6A9B/7MrCq0T745voBbwOiF9px+e3aR/brImxT8Sfs/tymAk7cXUtKc+Oq
yhT0KiXuJ+hHvnrn2Bdm1pzUQcQOcRVwQHj2y3cZMc9bJv/3YKdbUWDHWhIZRzxQ
jFn8tCiTH9+5qTDsFzgV5hqqTyirSPQqs2MgS584Thq2cxRN594IocMVFyJUL0GA
Vyrn5625ql2UTBAfvmXMeGWFKu491HN0ImWZEzldeUdR6q0ZU5UG+k5AkinUBKig
8HFZkJFfNoDa1HEh02WtEN3+k44M9JT5k5bXuKNJSaTbxYgxlTR9TOSKwWBleugu
4FTFYzJDyekeColOBU0j2o4ZXRXTOEZuv0JpW1MVbmm6e1LHMJIQr/igq5Zsq0sv
fb2NUo/KdAHPv4cw18b65GuCh07gaTsOOgdBL7qYGCOvxqxxIOuWd/AytGuS8bTZ
AGRBPxUrvkRfTuMSOUJodoU4FTm8074jNP43UTT1xxSCfCTc1sVt9tBIqUlUxqko
6kNPjs9kh1duwBy9LaXfeCzj08E1Tic8WKLtkQyv7/8V4m3CmrYxxN35uvHKfeHE
3leH+KqLL8zNtF/hFoKGACFLr9ORdmIDH9za/qHFoA0L7jFhvqTIXxdn5XNi4f7c
ThSMNTboj4A2A2FufTximxOLBbkgQFy68hHDJ7wUEviLz+DpU2R1sN8nWgeebNZ5
rLQn2I+l9C0VIr411fMKZIWasdSJX4pXzTyIBFmcy8+MoIdp3W5KKdkxqjdBWCJb
tZjK+CLiGGZ52fi0scBemAt1fk9sYS1yjwCtHi28Vu1gsMjsHlqK4FbDG4H9PgS0
1O7e8eNx5xgPGdqT58AmyPnfzM6LNenaIT46Ztv+XmTttqDSsjVFSWJZPpbNl4pA
hUIRgtXEX2U/oZB+fPt6VHyrAgh1viKLrEda/7CQFvm+Xmdttw3H22rKe11PznWs
GrULPd/oJF0tifCzqgr/Hk8tmWBFI9En7de7uKdG+TtExBkP1y8mFWZxqCoguQSr
qMjupP3aL8ygN65DnbmhivIGuXrhgQ5d/2ncprQKO5gpBPU6LFI34iGfUAYpRRnY
eHybPR4RRIJO0SYBDrPTIuwscRAsVAf3K8e6WR8s/h96b2V5scBbjd4jVMmbf+uJ
aziXn+ftAPHidpRTFf7hiyFFpXXvitOq4iIXL4gKk65ochcfW+8UtAFn1NdiAfKa
RjUNZJ6Sjq2hR2EYEk5bN5Sz0sd9kToqq8Lhxk0fgYWM0npm5Li8sOyZwstzu87r
Mh0J9KuM0gL9bsJ4vJ+gGocEtvX2wsu9u9s4MUoFVF72LXHOdS6BOM4jHiAlDwZ6
eXeCP01penkAcqdNzXU11qQ1lNyeMfZuac630HPfwwSYy2IIYavS7f/Ilx6/5gBB
6Vu7Q0LwXVwhVVuZ6aEdPEXFTpzhN5B2qE7s+Mwt1uIsey1NBYLz4CUNKoiZg+OK
InQXlnLKQNGz8w3sTHM5e0oSTmXO1iKcloCfwM3Rat35kGukt8SQ6dzNKD+fGjnp
LfkeoOd5AihP9ev2WT2EnRPfcoBWKLQK9LjF6mjfezKAVg9W6deYHiW8Xmph7rJ9
0VBrqn6heO0i3jg30l6Kp8zwgySglTZ2xNKY4dCzfZlPz2bF8FwCri4jwKKMBCGJ
A1DxTzphrSaJwj4zrI7E2BR/hG5Qqgbv/KiHxc6nzGLJZnt81M4il9+xY4H/ySkD
3XTaTrruwdasWddMxATaxrYHOH5T08igXBmgmQ0zN9zY+JmgUkfBfbj3FWzbWz4S
MbPBkpURGz6Wl4CBZaxZWKfLLjU9O/eaeTWB147hKdRW9e4VbYbiGCbsEXwthd0p
xFJWov//E6CtEDr6X2tYQinchd+2Yt231WIe7Pd07xCuLfEnkgZHIA0G0mNYh7Gx
Q+TPfoY3h4Ni9DQHW5YVAMtDUu1DG51FpV0Q9ukvWeyHl8oLAFx2iT35foSKEkz9
Tw9vcOQGFMMFMIHhia8E6VLskOXI/jrLPWN+DVshiQZzOQSqOcVOPyqDDk3Fy6Gu
bUpOvINYcgmhYWptwWfHTI6lkrmxPX/oRgCo7/r/yw0WanNOq87xFcKeMEZmhdAA
PGoal78Db7i4rXSlXxXlk18Z/y66iNmHzp7JQgNRlm0budBFhSCf7BCeeGqjSWYa
OZirefc5Ug5FX2tt+CsAjqKaK7+wb85pKzYaSHk4LnwOXm8E6KuNXW5W2NmrW9k0
fG54mBjYxWIONbxyhXElyPy9FgeQvBTC3po5wU+PFCDQEmlX9NhF+Mcdmh4caUf9
jkwKk7W7Lio6dd/bkB63Vvk9HUYDjgtI7PPgwUkF90obZ7SoIXT9UZt8SLEUuWiW
UNIoAEmnyCILQ07IzhkhFbc1iXSXlF8CUcQsBxKUK4oSdzV61yiYz3zI3YmQ5C57
B1G+OlKgUl0J1CL3cNgMW27TaiV7cDUQ8hFRAgqxbmA62V0poikVMQLCpo/R+jwz
nO/eAiFmdLXlVCkXuQGG4cDYhibUFYf3Hlpb9UnWw4TjKKrazZofHcSbWe9yTBw9
rYoXfCRwLSwYi4wXYNywwunHjMSZ4mcDYaxPRZ+92f9bEpgOZ0kOju3DAzxmX277
uOYbOkMzZ5wceAlmLdrOpbcRqt7E36I1r37ifT2ZdnT/nvfI5OyxmHTRRlUWH+Fg
daZhAS6LDRnys14quiPLoUdpVMp2FHU1Jdr5Qvs7ll3hyGSva8QmUDEfih2GSY6J
`protect END_PROTECTED
