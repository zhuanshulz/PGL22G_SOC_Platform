`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oLI4sQ+hzWeH6wUA2eQ9ih5sUGSEio2ySzQ+83+ih63WujF9hADTPoLJPhts8l8y
It8n0iy2bMvmMiIIOSK2uZwSW5rQWFun2HFX88ac5UZI6ArO/wm6e5lK3zfYClJM
OL4piXzw2XBbL+vDsane+D6CMNSJ1lls0C8k767KvIA3VvB7oQzhVlHDyieqUBj3
lRoDJVntzRySp/zibRIwTry5HfUjYelUOysrhZg/9dj+0p/7aZD8y3fR132ujjih
pW8CIr0ATn8r6FKS0GbdKv8fjtAALZKNsRwtpKh1YNOZ9f27mK14s98fYVd8E3jw
eKTswRLz3BRqcbCgwNqRFXkf2d7u+tNf9bRMOJdRnWtVKTyq7uM4y+0RoWGYnO1R
d3M9Vnll0eYtvxM1951moQ==
`protect END_PROTECTED
