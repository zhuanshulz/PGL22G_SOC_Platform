`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xtfeh1+1e4PuZrT7bXJFstvsX+mMFvxF8jmrSgJppXj4krVbwFVQMVS9TQr78WS0
4HB+KQNI+undsELytXcOOgpmZVoTPaRfRTVbcayCBy36EBHXIIrKHJu4AHwx/SI+
YRWKWpkOPrwxH+ZTEpAuCA2lKefIS+ZXPaWBGUUq3scm1kPhfDPBHRA1jbokiJyY
16CRIQ6dODg1UAutjYrivo113XR6eGK7x1ZmFFxrL/hzpNKXO2IIWSM4/H98yE6T
bCWw30maiKR733ULscVcf/FxUTWaOlMOca0DHHlHty2a7n75mUKnkgQs3NtSuZIU
YbO6eNANwoNz21HkMUTFbZzRm8QjAgAQDekm+Dz/usqMHBB2iv/39ma7BW0kRjy0
hOYD1i3GPVkjlCGTi8jW2/X5OaaHVy2vG+x/svyDBtMvP4tatLakPKXKbGdDteJm
W6tjb4CypYEsCMx3xuEpeSmCjkdXJ8THnV+hatEtNdS4vwEdx6rhppn+FfMWVm3x
+aB879twcmSBOZnYdwTF8pj3dILgTo//NoUrdt1HaRRkfjaJDsvfeKI8GMyheYvD
LxsIr804VLy1VeWZmnxfwwMW3RMf5M2gYcUynRjWHCr+Jyw1jiXQET9nT58U5GLQ
cqLkUu6nBburIkc+0QIle1GEpslKS40+izwMlmgX+in9AUuEL6J0OtPns6+uJVdW
UxMkD21ldEfRIkVDVw/RQrqu4FII1aWSq91xQCV2KylzUOrNWySJoZyG1UGVunXg
afD6BnE4avkM6KuQPHsNFweUaIZOKOPU0zI3ltx1Z4yRqojaYX/Vs05a5WS4k5go
cLfgycNqPXACGSvTzuPW4GmUOvD7xkD6nmj1CUocg/8QISdakQfQOs05jXqJw74v
lFmFOTtQObjpH0V/+TPMmECJeRgKYGd7ifH67wVDj0vpUAedyschE/C2I4BR9LhK
nGENdvJCW/95O2oany0u0u8lX5VTekE/PDrWSBXY+s36RPj9Bw6s9cmdyg+VnJ64
HzP0Hi+/c9NB2az8H0z/iU8ypXgJUYHl/zeY1DT35NFgZqsjEfSN42jac8RPRT0O
K9OODgKWKVrwpVIZ5El43eRO0x7BH4QdMtqUx/Z4bkGtJiK0V4W939QbmyqdVBbs
jBlMn8JL8sEV0RhKo8fa0XTeucL6w+vje4A5VQMAxu91D7i2Lw6TcX7AxH9Xc0Zw
JVaNr8UNCSoqnqdziQvDzWo2oftkQbfGTH9OIr6yv4iH0AA+GLpEcjY1mLCBMAHR
3JJVB307Nte/iMaOmn1thV2TI2w8QJ9NHVI159zyGClgY7yysRhEFVoj08guckDl
Kxf6tDhrB92JOTpRjHFZd2HaKfxJVbgtnSzFf82D0+V3LrOoHIUaCONiwzbeAjXm
5VC0mEfMCwF+eoe0MazXVr2/NgJRc+q6WJNOZY4jNeBQgPeYhPO7MAgFDCqu/ern
eRXEimeOfyE8cU4pUJFHOlnVZO4PZ0LGR3W+70c014T2ltQld9Veima1dKuGR8f9
Q8xtl51Ave7/KXglX7ML5UG9z2V7aMq7m655asjwckM1zdCbADz/b0XqCrtE0EWe
7XjMippNe/c9WAcpBp2SNqEXS1Ak6chLbqJ6VkWjpUIzqGWId/FSQI/5lr4IMzkT
aQeCedoRISWHI1NcljPujHNXvJgE3I1HYtyqumWIh/aJguHqa/3FEzs12F5nXKCR
fdahFhjg3sWdV6AbiwcGh4sCMjE9pvo4rA6i7Z+JE1OttnNkZ5SO2hb2eiLvXdzU
veX6FTgMqbE5MYc7/XjkF48eri5/85AUaO3c+EI0gFBP50dtdlFeEeTst1Ylsckc
i8DLaRV2PRJNOntnshIdo3hfK5fYFHRoL0QMace1MrOtn6jQWoaCKbiA444MQ6gO
M6j8+K7z+53Ti11js/2R19MNb6PDxnZJb7aMXoJEAUMDou7xM/wPaKxYe4uB8L8u
wesGmu06TRm066VxzwL+k2ka3Scpi5wsaSa9yDR+2DOvcneS5ZLvdKCGgdA5OcDZ
K6Ol0CwD5pZeL/3yK3RVV7W/J4U1UvOxcCcItmSXnE2KYYQx7ul+cSP6z+q6CLNz
b4ydMJ4FbQAbnnw035HLNcFAHtjv6IsOPi8kRD9zzKlDP3foyhlp/Z/fHGMfX80D
verCGSq6SD2crQpH5asFz54x8J7cLEvhsNHBQcauF5X+5jWZ3W39EmXp2F+edMbH
lrqSdR/Jq4axXl4PmdN8mVW5A01fgquIaNvCpd8cZRQV4eyGHMxMrjSEGW0/GXgS
zm4zMPu1psdohVZarImQtDv+lVZvwWYgLM6WR1LE7lS4sa6W18JoWHuElS6h7Shz
wItFcFAV3cr4M8ONENpnZmN8zdcvJ/1WgVFfH5s5zWWBk1HbEoTY/73hiC/yOdWh
yyWBROI4VL/bCI2K07JDFNG4piOifm3IbDZEI6lqG2V3wL9amtYUMf+YWkZ1o091
DtfoiEtP6HljWq5acMZ2UlTFd86Iyf1ioYF8M+nsNcLXY4n6dIZxSnF1suITHx6J
+CanB2LsPYn334oaA3YMtZWsNxbAfoUNQw9mGtHT1IuF7Z0vsR/+KUpHwy31+QU/
DwVeaclvGcx2J2ljLhatMox5RbVIbRpPj2NaM0VquHh3XKQtYZCRUmfTyhGRG1zP
mBysEwn75B4BQXMnVXqbrQsapEID2Um2y2RwQXIvenPqofe5rw+3KXaKJui8KtdK
8xPewYZ+Bee7JxY9r8Nrnn0Y3pv6yM7rvDbHdoThsVpvLt/9PGblLEm4q7Gj8Ub/
kCQoB4/Q0ayMTkHdZobkJA3QNkucUCaCwnmmm+z4/85nSVunmOGcRbQGAhg4tUzm
CffRXqOw3ugCjrRWX5DFcq1fJ8+E5LRkeNeImrK0GD4FNzhxAL6ya5eB8hgrApTT
fsSPtlSIyOmWca7uNEfl+qntgVcMBZQC1XsdLrcqU6bbs4qca6FuT8Qb8jng60g2
9O/MN84MvY4zJKTFzFIxf70aakmvwpgX/QnE7x8UP3MvkSrtWnfIa2ymdLvMQvId
l4Bov5wJI7VMUUSVDlTWeQJqyydi7gab8w1rvKAId1t9LC5HOUm8uYEIKHPNYHgT
RI/I+WJndZRFh7aWqgAaaE1BBYEMFTGPahuga7qMwzpA7gCegXxgd3EEfD1oskw6
cLoJUXGD+6txIUtcVyEd1FjoH8yS8eJuf6O9jJZrea0kRuFd4sYRjBaRLvIxRVCP
90LUuxmjfI2eJacwvMw4OgOJwotlYWDk1o7QVB5vSN7rANQOjdsI/x5k9COp4tMD
+UTG5txTR2e4ng6cKiFoYGz2hujbQdDY/IBqmPsLjVyIO6hX+QepFyvE0befGebm
7rc9M5n9/XVpuOOtMgkgI389HI6GRMXEi6sNako+H2WgdiSzVTQc6ZuP1lZjGmaJ
ULfGFHBq6fmPCsnnpfCeJtwviUyrNuhcFEe2bWZYwn/1XL9jlBNElG6jz/3aWg4E
ZzDr0AeMi0WEdhBbe4C6YofZ1mJflMuD/FytPeHZLU2BUWxXh+xnXJBigV9MPA/h
xD0jlGUNFlRjoTQoHOSnV63wwBUGjXsp+jMgtaV0c50x3MnLjThXvJ7tZN2jerk2
jwW1xzNarSYyZY7DsXmRtm+Lu1yYv0Kb3XU0jIAQPk+ETNYtuhx+eOumW91svs/b
9E9g0jFu7ysbdXxiE89NsCg+HKP/Zei57w70PTnm36ep452oMjQHc2BdeePp57dk
uqv5fc8arvDsaRQAfyHjiUYBTZey2VDmmBj7UvT5etxCfeNKOeDZOC109r79N5KD
iucuS20Ww21LHXCIWz651vzNqbq8A4GxeLRKuzHY/mrD86cYkrjzEwnbzktxQPUn
psOYVOxMuDC1G9DSR9oOlz1velyDfABIwwqYWJnF9eNvTCDO89oovCqhzxv/L301
gu2AqL+BRIHdlYIKFslh4Jm9IUVkw6I7xw7dx3xlMNohCPocBplIRyAbevruMKok
socFfBtJ43HKF31ZlEzAil5Wc2TIIRGL2lhTxQvmIGIWQNY7lFGyxKPgmmbgvxiA
ESitllKmTBUgNccUG5aVdGvUKOiI3WY6Hyu2+pjqvczjxE20IoeDozw1QbtDahmk
ApxZlj2YS5HOoQ3q2PydS5hyS2xS82P2b0SScPgiamBQbhrHdssAxr2O4lE5+d6X
epIz221aehCn6uo4yzVjOU/H542feSCpMYA78R9vyBpoXZ83hMFx3HAZjbzo2Lya
2iNUcd0shAZaXCUJA6hzmNIcZUPBw6okrjk85lFPldLlvt0F62xdV/ICZYLTTbiK
cF/jKyCzvXVM7BMxjuGDHYJlC4W6brnbz5i3n23ztLnp/vosXEA0GUl2CaxDIV39
U5QQFPPI7MOAG35xA5D1JdClTeggblRQicfx7tIiaOW3RK4Dbu01WKRfysSVHwAP
DArgX1ny3xqAxDMItQG48JykqGzAsyrYjNOZ5ny3vvTFcuoTls0tFn9HujPcW/Nc
BtWPsC+Ogdb87EDxk0bDgdWAMfcUmWV6RzTMIsfJJ223RbEU1cUro1gfI9rHQ6xj
21mMdqWgPlY9QzL7Tj+Bp9Erd//HQ5ydxhZuvYnXFbb1kJMA8erEOvtD+uw11lAU
OijPAIYNbPk/Y/MBMshgGpfXSnb02pxCA1mPalx1GFGHWXoIz1wBgaKZBVSYYGsk
uesknVzJMGc9ShraAisywZ99U3xuQrDCMMkQOsTegWZ35hHbwD64CMZMqORj5XW3
rHE6cPMK3QOJ5rNAVdJ5dQLIMVvIMTKxW290560m5A4=
`protect END_PROTECTED
