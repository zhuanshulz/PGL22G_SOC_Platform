`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cP2kwRxTYI6m45hieHaJjtqoNQO3BA9IyWhFZL5YFuOfV0MYkujac/C5t1NllDzH
N9YaS38HydETLS0qJDJWDIiDugy+zhWoEd1TWOCQY75mDgxrmQiWa4GSvQ4/RI83
GxQVCZ/ImIYVcpIgTb5bKu1JXkYCa1YwGyGXa4ntghBNy3qBF+laWAc3sfHcR/PZ
bsOxaJqE4SABZEFzKkFdXtd3poi60l8cA6xoWUrROnhMgfr8M4S4y0Bg7egRh3ZH
7ggBDgvUZDfKaEiKHz9N8ko6OKJHrc4LfcFDq3EAPDY4zMXkVxGxZi4UDWxKi8U1
VJWONv3RP6M0WM6zj/AIVtpFxz6+9VPb1TD+lBxGS/3poc+eyRFCNuV8cCPggUxB
QKgU61wDKv2Z8JiKwxe4bzEZ65XgrB5z+Jrn+bQCKiiSjN4E21cV29Xnt9cbiuNo
FeioD1rc5CsJCfCxAdS7W1+5AE1lEDjkd0/j+GtZ457Mut/2+2uVbsCjfWSShHfW
pl0juVXb9uUT+TehLfcQry6a5ubYobtPIojhIznTeRbTndEj9kZfpnsfoyX6IOca
jOi0lvod/9Y+JTEAIrFEEfMQuK7J0mCJh4sDi8rGv/9bO6Z9uKRPAuV6tmPRMfJx
4LcpMGspaSo7NOCJTq5EtuZCQO2iXUr2pb3gtqIVkf2enbAH11HnS/wKKTRMmHHs
JMeDRosQ//QwJHO9fO2573wMHC9NSd0pv5cLomqSx+FT/wl6wKzphReJjtIZisvC
+rmK1fOuoSVJj7u7YCbVv50AvFljpYu2Lux9iZKOKUmJXDgnSYgzlTekd6IPVIoo
C2svM6M/m0024ChNOhdkwVCo+wGPPFD9r2Ff4F7YDUxWUSA6/ShT+aiolhnP9Gvg
q5lU+0zfv/hCHYjBpfOGjkwq41+AANipiWm69fVBW35F4eKdeHhyP3WkqlY9hPIm
gMExskFO8h59EEB6QtqgWRU5rQGiB4mqIHtwFX5YzLt3bqVjkMQ9E64A2VpoLCRa
eBgub9zuROSLatHzUy0NdymzI2juC691qOtMbO+KlDqvfkxXVPAHhz9TczboEkxt
ips8y+yFMZp//GvQrEk3capM+YZPLVlee6Qezo9EnVmc+KIRxflSp8dkr3NQJ4g3
TLE0OlE16u7ufacX7/Fm+DIUPf0W+bPalOuVLiXMF0FOl3knBZtaHxwPd4EQoaly
MhijZaI5d+/li7XSYkYRqrrMOU7HN3vgavjQmHYeNK3JL20Dlz3TGpmi/sgSx78T
vvqWlfpeqA5PBH3qOQZ5O4gv+z1Kmic12+nVnLGVl7yBqmQS4IhlkDeXSpcK4Wdy
byMna7xXdxRr0K9SK5SBG1eLTvn/EbmMbdoaT9X2s2kIXHzj2+R9M3zCreWsE6Jh
AFhCS50AB05SOFXgk2ExinBBK9SWdCyXvBu1OzTxq9OdaKtuTvJ1dlwMh5B3fq6x
jCh9WwTW2zd3umskTSlQv8EsTCBOhB/53kZqruMm8mHhYaZThRYXqGu6tQkZj6bO
qZwTjTSHrVnr8xdfMrJceVE38Vn43QC60MLJfO8xNTx9/IyC58hkaltqAPhp6jSb
IOosz/HoX8MRGXUed00Nuo5kH/H5H1nVIhITDbcmI48qpqjIjlxjJdt6Udqgo1to
nMToIzPmoZOfdSOviiSM984tf/I8OTd8OvuYmnN8H3i9TDdiezEahMJOu6NDtOo5
9PZ8bTkfT+6FGZUUBl6BmYPmpGradTl1HJJ8e64NMzeUpTq2GBhEyqN4LKBMXtIU
eziuhtXg/cix/fRfkFDkrAvi67YWWRFDbfAM6F5ETMXHBDPGlBrXddKHTjRmupz5
d812Xk0s/OeZpdWBgVWFYJyYu0ZFTY8S0mgvmH6WNIXCh8PJYAOcUeJh73eAIgjX
32t/i/qAnQvKMBwp+QA3amsa3Y1y9bpJ8tGyYPLE0NykUKs3viLblkjkcNtfa1T+
ihvOMPOJPB1/pZWCRFbbv0bURU0t5kwiGMeOt0Iz97o7q4y6HpfaB4T6yL/D1fMI
gjXpXHBzGj7+owYOPZA56YXFEPd4VQmAFIN6c0ISSyx5ApjncB1dlffd6NwQehxP
VX427bHcGRNorpfy6oV4E+GrVZ7F0I3UtLkmT+TtVFsCySWCSIsHp9oYm3xmVyKq
Xk48QgEh5mmqvQ+ldqSxkoSkyQI8d30aexMJ2mXrE8M=
`protect END_PROTECTED
