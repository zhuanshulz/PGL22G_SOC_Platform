`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UBVSbM6BDKRP17vyYQ4jhvLxsw99zB+rR31vNdnh7y1EWLPvJJSxh/kB/8Grll0o
ZODc9kYsySa8l6tso+zAhb3dywjetHvL7u2aPXtOksOgtH7vFZAn5bX133yLOrtF
a2iLRoiZ0MdBVwvi2JH0riuGla+cT2ye7neRBxfnvQq3jLkzaYV2+g1A2t04TyX0
Eu6Gc0kNQZxTjpz30You5OEUkCZKekWsVPtNglytsBVHGRbZN1XX7c5XTrNyjWZP
UdMfMjW1BYBUSnM5Zq9xLdQYhTpkLlN6rVVu3KM0DWUKNPoUm3rXsgTHUpgK+MBr
MGQqhUk9HHvdZrCcfzuXoQu98nyJoHge0RGJzGG65WwJZ7lL8jqy7x9JsSdzK/ch
ZagibVguo8Fv5t8YSeo3KGPFoGXBjH7U1GKN6aAhzeNXqvHh/DXDXe13kve2csC9
NMqCgsQw3a5ONt6+yCrzNcbeSGYJcM8Cd9HS3pQH5Dw8Cb4KJzF9fd3uDBZmUTjY
YVul5GYvnKDAosNHkkuXdxJMDybpWqqHqI9/kPB3CAp4AR6l1f3tGzjql08ovXSG
1uWjkfOfi91FIw1iUMMIkUE/6z1Pxbb7RryflfBYmOLKvQNZ/Q768mfDC8J9N0Xs
URQxB1PqByWhJzWP/qziKw==
`protect END_PROTECTED
