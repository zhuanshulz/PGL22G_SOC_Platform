`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuSwg2lrwDvmVfYGL8Fa7rJUoOD+NMI4xmTGAFq+0UqHXfDlKPMZlh6vMOKGZBOH
jd4O7NKMI8EJjsFvyLpQFGeqCCUIUI2YKRQPulFdMxsgDk0sX6NfBO7jn43zPdzI
Fv7Sw84EQj0EOlPF8BmXcx1bGqN/blXtewfVosl9YoXDknvoUyrIcv1F+vsEhI1g
5c9S0+cm2hXn6OdBSnMHo/NwGGKJGWlVwjJjWXxsKlRt1a+sTsVqm8vf7CCT30qZ
ZlKtftRXVL1HKLlAGX3C/vmXFY/4gjmlbMPwA75llBOUgfpQ1/pZiGWtzZN1vfRt
9oMzEaxyAiKtgKzfZ+8Rb3Ks6FQ0zmF4Vzv7sdewKG14gom3AQ6txbHRwMp0OMWV
Oewm2knIpHYabzTKvsw0bCSxkDP5yf4+QwiV+yl/w7V4phIZCqYNlYpolJwiJrGI
nEFGQ8oodSfZZW8NxPUxz9hVXApXdVDEX8dYG+P0zIrUpmrJgUd8Guhmv3kcywUP
FDybpbh6dNaRvAktaI65sWv/6BElVx7lAtfKLpwnGeWQau4aJaAlsS2LPd5rxiPI
PjdqP83/Rce8IbZpGo/HbMxn2GpDdFslCHxzptJTQlqBJNJHlB59bTs8MK8z88EQ
3eFExfTrHiTvjbNn8V8ATiQ4vMQqdJWpAkjeeho4r/vIBEXVhKtFL0xDDTdOsah0
sKcBZiVqyMVIE7kS4nNrxwhlFTLZIW1UWmYCtAr2i0e76BBiQ8U4pc/pT2GIdKwI
olFXrgiLCi0LwKzudI6EU1iryN98cx1HJvh+M2a3pMQ+PVG+KuE8X85u9EDb+eVC
eopKJTWl9QD5bWiPfSOZpjZpuEKilp6s7lrMsQkr+9nCYk+FtOvCvP/4kE88LBTR
2ZxRux4g5WTZZB3hQLhyHW0E2vj/ymfKHrQsWkAcYSOuGcI8GY4YiRFyNC6QZPtO
6OuA0miCAnlGGNXUuN/qG2eK5gualOCkwhIfug0yxkIwnrtDr8G5BUgrUwncbj5L
hMx+fFTzhdNxeqDh41oj/4ebTW8gzwYIxOwSeijEhOTCXhZbwbCgqBTxux4c3qIo
z1HxT87oXUjAOFwvR5g9ZAxjakMl0PQgnM3ET9XbqzVJnbt3getJiNpXRs9GpCqx
UtLBHPvwH8fKsK2x8vWyO+ESzttFkNfFELLGZik7m5C6Ta6eRWzakujfmTooBE0r
djctWoCVdsOCn9HpZC+CZ5B3jBvLRS+o0w81iz59lj/ZfviuyvGGLlHeB38qbMLh
yo6+XzbiEHV1o51aLBxyi6CiQGt7UDTBnefP7Ycvd1d4+3Cz2AHSq3hokszNvWYK
IecEHN/hBCSSyD6+0zqST1jts8r6jGCO0GBN0ON5xYjtK5S1Ayj4iBCOJPKh565P
UP9l2pGAjcTFa/w32bUnp1LJduhQktYPjds2rmX+oFI1ZD0292RhVFmHKRb5uphU
0m0AeJPMcLzcYA90txOtpmcMwjts2TpxgE14R/8PvV97jlN12SlXvkcVrRopnSpO
qyPXd/L9l0ENFck2TH7XImJh/mb/F6+v5AtDU60n+bN2zokKSEa7fT2NvywxsQJh
ViOJ+0jS3rylVHhf8h3DBK+D7KbKHv8uk77lk73qbtkwdEhap8BiG2/5HalVIAaE
uDiejb0nKhSctaOlWP2jDFGXV/3kO9tel4WXkUMHxrShnyDx3THastClmYy5++wi
cDCa90agdA4RLq6pmA+rkAiblmqvNPyTUho9NU0HGRZF8EB5EnyDxi0A+v2DGldF
DGe5LYetg5kpBNIX5tO+weoPrDpKUVSFl1dLIHKbak5mdgjE4BbStY+Jjg0srlqw
SKiqRK5I3hli0Yv6/ge037PbYAmLYTwl6TPyXCyZ0nfNSmKvTdr3eYmFNL7j6eoE
+3xNZblUJqzqT3uBCzfm6zj7vdkn1i2SzFvfD7j10vpKE2ek3GjI5YR5IvqbID7x
c+X5lqbYlSlUubANcgCcBjIhftAr8qR/y7nwxVp0URcUTYV2M8Hnjq2zHWmMiigy
GgBt/WM1zZTR6K9+3HHxRDowD5SKhQDpefh7mz107VcumF6esmg7D4YmdrbCyEju
7Y61mSfVA8iwSku1grPIhxWKd7fINv3Xn02AaE8ijkHTYqVGsLUoEybOElmKak11
cTWHaCon84QIbKxApUvDK3o6H+4ytpaQgbmRut+sw1mW3Vv0SrIwkAHSr2NSnC4n
3hpLtaaoSX9wDqQBw7KyEh8bOT+bFhC4daqiDsp3nXCp/rjphadk9YdanPRLZW4S
QB8X/KVLrnip9SYMNwSM6gLp7ApARo/6KgNNZd/tPDMRg1c8a91zelWsuy0xtbc0
kAC0FXnu5dSdQGLlMsd5A5/j0rrbnd+Cc2YTPMTAWqFm9BixYeausTdGb1f4UiVf
U80f6M479FyJzq97kiLTJFYvRXTgBxWdi1HQvovZWklW2JXykHlVoXXXGUgEhOqd
KRPCZVHjNXzAgs1iy6Jt3q10YlO+jBqBp7KR90SPEQYvQ0wyr+c7GPTeQjFq41ox
tm0YsaIAReWJRbcOAAt3cia37UFXvQ786NU2KqsTAbmZMhSfnfjOuMjUE0LpbMYL
Vq4QmJMbvC1jP72vd92hL64B3oyJ4wjszJXbKKFZGs+InEI6KT255Q3MxLN0VKA0
71jrYt/wIaBr5/wUmOfuXTLHkOd7AATI0eXvX3VBTIk9rAth+boa1tyzZKM8+6fj
kp6S3qk67rJlWDIzs/r0hd5SoUSUstC4Hh4q7Z0aHHst1rA9y+juduXSUVgSCkz+
NERR0kbxpjSXcVlw7gCipRFf74Ercd62LaV7bVtU5myc4l7x1KqXDElRunQn6Dhf
1KBaB4ZiGM6v7kRK9pOqiZTZZ5ZznWhyGCsUGOqeQToNWoProbiDpzaI0mlpjqh3
jlrZ86tMGcwxC7o4lsRRNMVthrOlRGvYSyXzhsdDgFJa9MobvZ/m1CUcxn40Ty4s
a+jLij4A8KM59QeHRdEpsg1xcI2Lm/60I1Cj2NWB+BW0gxa0VEigfFELN6j7yZD4
mh0AIk3VNHsm8zQ0DOH+PD5KF6uKkampaWdWa+GsAt22pZBzS22mi2MF5jMxp4Nz
KU5qSYJB4LsNlMNbGFlCpHElAsbtIXfA9602Ln8Rj/PcUc4zQvJCrC0lrSDQboxq
3uy1YASz2kA/wfgP3qY7DHMBAM781nffky+IgfEA8QfwPVEgTDpP3ZYzsaHGZ6tw
TZ0xIu0vd35O7W7uMNBtUI0GybeuhcnhZI01qLw13UNRvV1jGfs2BocLflLEnsF8
4xN3dG74k9lSqClKl1qBuu+eSS4mAxZH6QwIHUI75hirUXtdRmOqvSkCQcaj4LLR
E3fquf1Pdx/5+esbYqq/8jvQR1JfTf9Q2+KQtNnfE9URhgqso4Yf9Q7a/XsmoTW0
o61wFwHo3NYhgGKjUr1kTsoWZdb1uzxOfREU0Q9KCokVpEzB15rdPS+j6RcNvElh
Z5hOl5JA9XizZGmlM0H8rDANSd0oH9lZ05G+zK9EvFm45uD5XzQb+xMl0/aVan2V
9IL/1+4GbMAhS8OmCBcE09JNhV8Ld+jiGWdBjCFYiFT3jZSmUIsS/xoGzqXdBz0Y
sBvo7jYhFQtaNBOYNRksJhZH4VpIPOK16isr+Jb5XycJkgkXmUk0LMUyOAJfVXsX
c3oYvehFlJOCMQS3pIGyfb3jw4ELcj5Fs5awWCXI/mZv0piROXhKLrZ4JydjbC7o
Srem9T3IdKHr7EWlTkzcKXX9KufXUp7y0qiHWU34g44RxvetBU1JSUEjQTHHToli
bWkvQLHq0MGkkdM2l/tbaFicAzS0IRDtYRf8xFuIW2cs5RjCPYwaZHVmkaD93Bgg
PLgTAK/iPghtBwTJXcDrjYauiU92vICjhggz81PaoY5pI4PmgHXqU/69hGNfrQF8
oM6dluFw2QveHjdB18sX7s/yn4MBYKCEOj36rGes7DvrFehbA0NC3z40q6Y0rylB
u3irYKF+uXzClR0a+aoxWTo6ngmCdL61YdZO1CqvaTUVsq/dVq/kXoBPa9bJ+qIB
YUYf10AlXRzX7IeTx4w+Qx+CyZLY8q/SjbtEQC6AuRYZfnFqYOR8q9hUw5WTl/jG
LUPfgwPJQFgj+DN5a934vkNfz8k5vdxoo6xugO3227po+23xFZSEuqjyQzGS3t/o
8Isn3OzvYdTwTaWu5Ioq8jB25UqwMUgxVKzNwT2GxkEpKREFZr45ArBNSWXp8rEA
eRTlZKpgWA+Yy65SR2RORXV7rRhJMDAOMRKsKm0Ez7GMX2G6anFK/ZoO4xEGgDUp
Slbult404ZVWDO3UwACILEIl4MceSHHiWWaqlivQCsDZVIxmRBxZvq6Qlem8nDzi
SwI7yrItCfCyKGS+r9UYfF4IMOTnBfR/AP5NzDG1Q/XXU3kK0Bp4fjbAG7qhil2K
7BCTXHWkRSzCUN86UI4ESEvFqAsfCeUiZTUcgntKQOfwV9YPVsoKM/tyVtvr+Qiu
VHQ6o5Ubr07+CwGrlCuiCRRGhGceKOH33limKb03J9jcZ3z2OLDWnaPkRiemTebw
cKibv9c1epivHhJ1LDsAk5CNTDrf1PNrIlHFSH+5kc15nTzvlu++18bWocA1bR1Q
q3xjbge5jqTvPNARSYv3gMe95Y4rbq5zR/u6DACdRFodi+828f25kmfVwta+7nRX
guGBc99gg+HcmRnYmwpQr3V/4qaVt3kIDJSywyPetmH9UUfAFibivDHL2jzGvKyj
V9tAUzZpI1jUTYR7m6pnSkxltDcQ8F/1PlkQMznJTC3J0ZYX/pUBX8PVXrZNpWsl
McGJAocD4WRitCbNTjxaE7nYgFUilTR49q96f+7grZ8VbwjiQ+Q4ix44vrkUSxRR
Vmg7TzGin6ZxdzO56etadZ37ch9nSVDzHkWFDtt5godT42EVyDZ+OrqWx9mV78Km
2GzxruNuHUINa9+aKS++pWn4n0VYPY3seSwlxF+Z0z1gyje/inXFnB23n7CKekY1
y5i5WQHKCJO9oZz9Yegu8RIetWULFyjAqbRcO/fpQL7jvvHA6ij/fnX3308lraP1
L29lrJ0pNA6wbnvjXdsUQGHkGDCB+gx/QOzfVnNBdUNJsbYYCdcTX9Ouxdq0doEd
hNKgc0VoJRWtVAczjp9mHobCxaJVjWAdTRaCXmMWdMmnpQrV6dVvmiJMjaSOzjSj
j+zMeCqmkCseIWodTFOJDRwAG3JB9HwmMiFWDI5hPVQ25jvvZ0NmqbZhX2i5i5kr
ENcxgVJs62bt/1ZoJ/DtW1jQGb4diCb/or7hNJi3ZeJhXBURpjLVCag7C57eZiKC
AnsHp5J0sNHBgJ6gJp3cH3HDex3aJsT2sBJMarwQZ/jFHbUCJtaBSu5RhP4XDKA2
XVNF4jvSRCTFWRSGk6LTnh/A0rPwbnzhCdSxda5pFxKzOMfRya7KTPb+FL7iths1
JnFDtKn5z01GJRYCUZ1UfwqqH3SyuoBuRJ7Ex9wftv4abCzkOfpuAHs0u8G96F8r
Kn2qLcaNhDTmlpuXUKQ9/nymKC1VzrpXbq3paBW3ioxETaZj4yiPAuYHzAi7kEZP
MHzdjxWxx0crlZx/D47kimKbgbLeFlNfhE8xyvvG+Jy8kiHZ8cySKUME/rREyQO3
D7KDF+HIMPBop5t1/o/GuezDaCfiLdIWvHKMh6fHvoI8yKfPIushIqHFwTxp/AGp
04J3OnguMvR13sCJK9sXVp4kWNelWe687D7+yoEX3wMVTgbd6TZoxxy/YY1nb8ng
FoAxZE4BmGl+S+iGLdf/XZj1eeQtNNRko0qE6+4fNG6EBCn8vxX8p1YqFABfyjVe
EYS9cX/2jRFdPZKpWGEhHAJGQJ0i6bp/qP3cimXu3wbEm0aqSqq/x5wpyaXdbtqz
zIibFFHnIjcb3CfFCewHJzNmDfiCDn/LnXUCs29AUvoOmNqd1cryX1CgmQtdmqMk
IZTUdRL7GLVZuVwEeFaPOprdkdTOQ5sGEeXH5uN7AUCC1iyzI6ESDIaXnh7mUETD
6oDa0aCyFHVuelHMHUbSSzP5B2dgrrdtEkNML1+gcW/974ZDdIsQOjgaG5ryWgM3
V6vnnH/TVjbzHv9qmdt8k1LreXljd1R7OeOtNHG03+t3r84UfeEWbHNX+T8tn50c
Am9CpudQBc69rqp/oBM2gGRdjKI7OaBVjcYEzwJx3gh4IaZqPChki7qWiCOCnlo/
8a+Ezcq4Wqj/qSUNxDDGUr2vNrf9hMYX/AFU6CQ53o3ei41B93fmHjReLJIbUoy/
Q3ASUAxED8bHcriNWjsvSXJvsEKDfHAM+niqtn6er5nakzI8mCOGA6pvSAnAKTeC
Nm63tQ6+tuG7UT7ljULMOLpoVTrFUn3AfxneFEqLrMamdcIotR15XicXP/Sv+wQp
z71ctebX+e93N+sQfUFKllXR26n94XroKm3rRZnJauL08Rf79y/YRCkZsVpoC/Gi
J/ps54jRoQFJkWon/VfoC8z6/erSD6vv9jJMtoatZClqVICEbrL0lI81Gdu3odZM
Bf47a9ni9HKKa8QPXY38AyVqasuvrlA+imYg76/nLL0BfmFA2HtdscHI7ToEBngS
X0vXykDukP6H4KCwdLxlkhdSBSvgiJ0s4lHjfecZTTQHBGjDGnTXTjAjYmexubsL
KLN+iHZmapP7c9HmZmDm1z/Vo3BdpgFfTBo2VnvACFGE1T+S8h+w+v3f8QLuQQJI
TLmBYOoFqQ+QfW/YrlJPBspJ+p/2EPOMeztnjZMAUM7mHTheUeLwexHLQmjNTuc+
sZpQ4MPjsuT3FsFcO9M72csReC31AConRiIuW9tS1CcL+WR9cH3fq2nebzIkikzh
/jM2do0THWGQy6UBdtHLDGn09gAFv+cxDkGf6OFgF7t17Csgf/vL5dIHfR1Qqemd
0xB23lzj1FBLZ7ditkLkPiWRA1YEy1816num63Y+f1TSIJ/ISLjeU715ScZ01nPB
4cbbXJf460rX+uAbKN0i3O+R2J/dIyVUImrvVl2aQp9c5s/MMEbIvNZk8gGh6V12
rpnf9YIJtJ8O828BgQfcDtLX020TknSXRIp9sdO71hyhNBLtx0lHzw+Rw/Huz1XL
K6JSqljhqr28apU1x7f6hbZSa+7FyiYj+DpyKvgI36Hmi/lq0nkdUgqt7HMlKQ99
G0a11L8GvnUrxv1gxaDeqAEl5MOdIryEFcAptWAMBFbdWAlCGjLM9GDcY704cH4p
qRe0rjtyuKHK38ybFbmSPaheO44zh7n6Crpn4gwd4CvUxrXN+g7lqWWMK4xvsBF+
zFCAzk3RIF3S/eudYi47iY6fYERIT1x+KBiVv9shzK/3V7KKC4FlqHoFIDKpvpql
U2TA+Dj5wf9cuklT/aJ4/7Cp0d8eYU7vpRTo44MILBgRjQ15qqaaA4wiHCu2A2M6
OOgEaMflbT2nEO9hO3VvH2e1bs6fFd7+DbBSRSVPnJWrG6z9cgNWWWYMA1e1YJWE
LvC+rEw/Q+BMKm2bO4Y1RzbiYJLDzn8U6HbwTM+Qt7gzmcI5gwtJdev0eYuMlbJd
ZZwYGIIdCrTogThlWip2mCbMpStdh+lU9GOumgHR01lRGNfSa63Php8GNUD+OdDs
FF9NFV9hopE2pXTGWJU8OMGvVKqMhqQ+S8LNGulmxiBZ9wm0QCgCOTBrX9aB7jtE
rPGc8BaFYmFTjduBKnaL2Ow+7cxB0wNEA4Zc3L/fJ+m5326e2dX6AycGO1vODdOQ
VZ4ndC45c2dylvKf2eSLLMOCm35rrkYZn2/Y9s4lNDP/GyWI7WMdwuzfThmGytB+
vLuSiNKAEkPn0ddiWhW4MdXqTeRreb8LMxZpBseFElXsDGRGOEzbZAicclaMQwDq
imxVFaJV+a9x0kYlJIMMPoisQOi1UacvcmDXXjCyBg1urF+yhdupWdjsUmk1qFWl
MvxVjSOpgmtLIIgacbaq8iB6pFtA6x9O2to+srh7JgaX9Mx6CekT03I3xg7rye9y
NRmyQsKDlJjykE/5lbXBYJaO4jYCWTacigXAk6WtXXjTQsIGtKnirv1+Nyfa3+NK
fQpcZvgIMWlefA1zZOEBDUoiVcLFMSnZggx8VrvaPQEULkBf80MBcQEWwSXssJ5b
3DAoo3lwxxZHHvQFhYNNUubkFXVg4U0/8gTrrBeUG2yLiETOh9MuiHlbGqOY7Nxq
G0ZprYaeuVt6Br2N/g9gZcqIbZ/PwnbcNZWCHVTfPliyF0AcUPu1b0LIstTv0qnX
gl0RnQRq6UrJ+6BrPfZwMUsXsJzNL8j7gQBHOOICpnFzK8oikbrKOwy3CTDIviYR
0jIxM5qvt1y3HNY6tS5Ak1o6lp/+o1jFyJAKQvXl9Sw1L+mHJL2/Az8hwHLoJn2p
uG5FUDuJpkqEcHtnNDw2vo859YlPHBjBan/sbEG7yg0gWb56etz60WeiIcDjoN8u
MhjBMmmfVT9rDqB/fk4zD9HTl/MMTbvxvBYjALW0uuPyiokf/WIMbYd1iE8SuVP0
nEIFBYnHIuc3QnbUvH2q/9pY/WxoY1p2/3Sn5BROfGpSfqE5erfN3WpN8f1Jrpcq
jtXFrOAz3LDPGUSe+2EP87hNlldpLPL8Drvxtq48Ws4Md9F1Fl4UhkfwhOSthbtC
qONFPr8EmXHIe3wJLNN5sfsQGnPMJyGTp/Atog9xlKHuCUrNIe/rNbKoqcBRgGAI
EM7bK/vJKPh/KZZrt5d4QAR2ZZRX97X/3V8kDV8lD7AmVTGDiXXOCbIKxkreNWKM
yFPEaph3tEF2ChfK0vtSoLpxxvjyc0NgAnGtZ8fYTnyGdB5Hct/Sjl4yKTeBnL2V
4YJWmf5FAYVjDhjC9NrqjA5wHdT68zmXxjudxDTf924YLvVgs9Mrpfy+dZZzOGId
8WzIcWDsZ+cXG9M+8+4qXKOa6u0R24qaf65KPhWUAJq3UThAIio3Uq9DMwYO0ALU
p9BtlXEjSKjLqinoja95YNrjqmRHll3BcKUqviybwpQXlw9bc2nQHYP6twW2u23D
21HWHIAYqartpfLmphzZyfsmbeddsiQAOeMs26UwQnnfShRBG8FY06ZByJ3U/+HM
S+2767JDwmu6/g30uAEa7gHhdmFTh9Sdeg/pQjVyrMZ+/XCGH2aHSa1seqYLBWZQ
oTj7niqHm7jDbAc/I1qD6jLKIfoyrx17Um1EV7c+OBe6MT9aKxtehkFLnL4Fc9JD
P6hEk4CRHDTgXK3dxokWP8ct9xUFA09TsYmcDx0zHm9+mitoI5gI4YyOUWRx8Pn8
F+eU/Bx2F/jALxvbJxBtXu5X9wszPMkRULWZAB+B0aTyN5nHE1oBTirE58vXEIMk
XmK9cnT0gwhI1Zjr8irCDbvL87gcKPk1IqwrSrOkTakWu3VLewaESP8nNpK7ax6a
NRWIWf0h5JCxYDco5LeV8mHqHkOgdICJYk7g460n8G7mksu+NECUe/vj0iFImnZm
00kLATbfgB+uWToW7/JwvWNK9P9exNp0Hrviv48eUBOLNb/gaiK7HgG5WmzK7lys
Ib7r300pNfLJAmBgmY4J2qGfyvjcb4IpLo3NBt/5PNICjyIrNvcdWp1ko9WNAV0b
5J6h0L5KZEzAwZjH07v/WJBBTZhE7L8Tzfv9aJv2A3A2k1sTUYuZu4wPEQrk46T8
/kwjd/28wJV7mzlQX8OcmO8BXGXrmCmUUxiK0vilo45T52kHfSLDkQgT8zy794p+
f2nEPBuNK6YQA5wEfclK0IoFVEWgra7RPyk7/soJ/6ZPlIgTo2xDL/KZAdswXmLI
S5VEEZSGrN9FTDyQXoYaQre0csaULo4cvU9e/xPlWTlXoEn94mSsb3aqEjs1tFwZ
swejGLKflRRPavw4wIM1Z+n1MneBENTAff2webTw7I6sO7T5E7tXYCa97PDOt7qV
pc/FvioabBT2M1GXASmNJYMoMQGLRx8Z4zq+jlf4jd8hi5DFJO3at6lXYsXXniLC
RPqEgVoLGVgD2Xjj5AhmanNnBGNSOD9MFfgLbE4a/OvYi0c7QQSyjOIT/EWz7l21
HI+982yvEho+ZXmQtoXrA2Mtam4lNNSPqbR6uYr7uxPwvddGy1yNHiYoD4mFUIJd
pdo4kJWJsxb4itWlFmNHEHTkyY9r0Tjgk2jioFTtFgjQrW6Y80yAaE696DbOdrOW
Kms8S3XnrHRLkIoVT5AtHxgdCXWqzlN5nZwarzHDXs/ZdlYfki2G+8uc8BULuk/B
uqy13QB9fdM9sVsxJbFdH1wr6UG/1w+C0PyUFuh9qLw92XkpzHKQp7PamL1nTIJt
nhm7whefmpl13zqsXSBty1qBTxJTSv4KyCAQkB33gHbjdBKah+P3V+g5Y/PALkxq
Rmmxq6BSX9LvwpLknL3X8lfIDRoFtCgk+RUCZFkpDUSQQ7oGecamEp8gYEiWj863
rNN4utqPLKwZYDRSibN2vy0jln75Bf+pTS9MSvciOEEknz2pUbJpLqDzKgEGKY3T
a35PUAngi9rRVetwxOIhigApLSjvlLGOj6oidPQg2U4l196YoHEZZcre8oBDWDQz
AtW2qKdq6oCNRTQjSGp0K/IB8dlNkD4TTiKK4ZrmLk0Z7YQ+S+C05k/N2CMRR+sz
Z1RvhjAUFQx6LgaCys73W9+LZgp25OljDAakhBGg79uOqQYcZAghG5u9vaIo2v6U
eAt8pkUknAiBhQ2LxsvJLp4w7VsbZzz+o43SHICwkp5X+N9p7NUFXtFGY+RteYqh
9aH/NAa6ibtAn9FoSZYIvCKzoFmgKhrpS6D7WxZH+RCj9diVPuCh8oOcM3vt+4gq
g8U3ynDzQoS+FTjmBJiX7cNiijyCjqwDTKK3BGqBwkJmXO9mHhJfm4V8os2oOI6n
q0RX4jvv/j3+rOv+rGFXk2k7ELh+mwHgMTSewVY8TQAe5qA8EoKWHcjou08EIyO/
hIWC2Ct4iXwyVSt1JBPVectW5FNPjsfXMF2n6MNefPFlbn7oGuNk5kMKLilXaE8R
GuLu6crAhHtqZDIH+xaltLouPKZWvEe0cpNIaGDDVbAOut+bVrThJyUlarOg7xVH
UgbS236Fw/oZus0WZ8rPKtqNHBCWMw68GHe9HWhuwB7RlxGiMmOQRkmX27zF0O7j
Yw60z+7EtADCAsQi/uj8U3PUk+vWKeL6k92Wk5PxALDOPM+ljlBTbyKHbEskjGTD
b1ECAp4FhW0LTD9lz6qHISfQQ6+/T2OJvrFAYnn4cKK/uzT9DOQ0+c5JkYcQwStB
fPMuF+mV3ogCa+kbCAmSMxMpD4Fm2jPuWnnYyJKrVxWnLKtUIbIRHh3N4j6p1J55
WvFFRxaP9aMGk9eUXCrvWLqb6hg+W7EHYd+ble17VRqFasmvFSP9G2oWXnSQtUF1
TXrUw+ab7KxgELNNcTMbAk09WVnl0b/NDF3NjG3sY0piSF8gB9sDUyAvYqoIvNSq
sE/Wgp4KMBlHIpz5mvquePQdRJiesovsf2ZeIXiboDL74K9d1RKHo/rD3NK/94/l
vmMizc9lLZCH3Ow3PWEKeD9Mcwl/lR2QUqoxpK8hmkDsu3BMEr9D9nbwlQjvo3iP
TF7J3PQ0vvTmMEgc90Y8VLMKPBcfe7tGksXTCYtsHY17Lw7frx0d8CQUl91tJMT0
EXjeKT4qg0zVCChNrTprmXqyHDo9fqjms0cGSvDFoNr0fMeGzWhpbotOMQWIXjDR
mdV5fl9H7ABfanqT0C60aT91dlMruKb+zrVh6nh6agrvMN+AknFfqHypIYMmpmUy
ner7Rq2fIafqa1W7yP4Lj/HeT496+h16JOl2l8rx6fCufe+FG2CdRVSm/KmxSnpN
ZQB6iQmFdscX6/lO0jgGPSVvqhR2qPvZJwd8HqrYp/gvAH3VeiwF2gPwWue0V6XX
jVBXl++T5lN2CVEi26dp9ikRRXRNOXV3o3R6FizonsP8ul0KTppZupGSt+zlX5Jp
y6RgT4JR288LP8VmxG5e2H691v2VV8yKHig36VDEbetWC5hrlyMEA2V4/OIvFYmk
ry4E+F75elOZzCWymaO9hMiGNjeMHxGXcfZefrxWt17QBj0mtwEAqyCli8S9eT+F
Eyh+rh6mBoW7TdKOPQsG81GNWecTPr1Z40nTbt1wIUQlWKcaA0k4vvhMfPFT3FD8
27AxaCO7x2yiEPWUvdYnPY3hWTKORPD30LJrVdW6q9RoBDcUvG1+D8NzZT8JXYFp
vFTC+ghf2V/nD3lNXJB5z3A7V8rO0nZFe9eu4sHLP4UUEEGPKn+ZZl2XN3C8s+a4
eKI5S/VNrpwcJvg0Qjtkq1Rn0RCKCusPT4aXyO35g16TpRjnw4O2i2y+mW7mi4q1
f6I9QwY6vpPJj+nlngGwpbosl+W9xuJspjaJ1l6gfOvvIsB1/bWeaRZxC/YvLpDv
q8AVdZRIE/emI7zeF1ejKawe/HUtdm+oDN4s8NkbwCb2GqOLO44g5Vq+ZH4Fm0b5
sTaX3/r0NbuhihvhJdeQUbFauMFwQ5fmV5X/2fEc6IuC8mJvaQyKOYR0D3atpcMD
gi18gXfn7o0hGAuknn7YuOIIO4FxXw7O6EVIG2cQt7y9PlE7RhDfEr5x/Opc7B1B
97aTzSF4H4XaGDG4keLDI8FtZMj1g0I8MfoKVWplkojTb7Xu/y4/DPF0aYn7Qnba
xlxEfwnw8nbr/GMFA5OJm8hoctyTgCDe1Ht4PXMEyBR5nst8EgHzqL2g/EoFFotw
jWSZUL57WnyYsBJXmCsWkrIVo2ZWGi1GiqtxKt7OKSbROOfot/TpTjBNUlWU5kjO
kc53ft+7GrvVVNAMpbVVRTvNnTDk5SZM9mSvyjQjoDIxwrlmEwKVRfDR6vDdv0nk
NljgIS3lKmdFcEsbwDCz8GrYlTfx6YCmNvspK94rX/aK3Us/mTcTjALJgyGp1zJT
SxU+PNHnRML5JKtsdy4iMbXoNDB5Jk5tfuUzR+XY77OZ7LURom47cxaqrU2Tw9Gu
ubWHxWsKodNs9E2IyHVzwBUiVOkZF6pmzOZ4LWhTgiO4SNAwMs5IiEcf7i+t3VwR
3fAWHDaQQxfjfVJurcdt/retuOdfbHSmgLSl13rcjdR/cbzGDjFZNd2Dkc0obus+
3rWzAH3WLJjhNlGwRh1FZ5sRgS484vF+HOEa8XGbvvbjH+tM9p0tZlKI8xzrcOXg
zlbJU5J1E4VDvluAL7DO9bblWzUj2pjmPRUV5QBZ12D22maZmWePe3DD64bdodw8
hXsACGBz30BnSC1dZXm7Z6NMZw1G7jCi9LKLeSos/3JM4mZcKijxvPoq4lk9blO9
pu3FHxfh+jfEEcu6dJDAWC1S11b3teGNED9Z+D5tnaB7RBG5r/9o7Wak+UpRtPng
XTYCi/86QIYQ5J0eJ4U4InVuBuJbZmQSZvftWu58VaDkV9kpsOKJWILFDWqdMb7m
w1tVQNtbaMT+HMA4M+78TcfVRxXxEAMGXtSEF9tFs2NaAoU95Tlbf7NXcObvjGwz
fXin7yfp9sNFJGR8zRWZ2SOSn10wIETCLypOAjbdlD9fhMx8lxfnaD+u0cySCSPJ
+0eiLUn9qtWaUSbdQTMDsFBCPz44FpPtWN8M4Ewd6HKUE4WBaIE1nzKDMhxckojP
erRgei0m4FZ3XSuGpCnjVnjmE/xJJVyaX/q8CjQtUraYyF912b3hQhGVkjtigsp0
RDdGf4lmq72b8m/KKu4OFdXKCT+sEYJR0yHGHZl9xSFptFvOloVNep7a9eoELER6
dIL0+b5dbZ226vW89xOXfNFI2ynOWlsMzg65wb8eemO9AxXTBV6G6dhlU/FVOpaI
QdPbq/1bOshuvERIVbtlecUEqAQuE/EPChS4pbA/0Siq989RC/iVgkQ9WdSCJfR8
YTO0958DGncWjOPfPgB4U3E7jX8q8FSZUpjJZxS4wrJjjKvF8/u3HLkWp70CQdDe
1qlFkZudbAfWc4cHOUcIieVXtSmgnRVKpfUHnRz1Ke7IQLadbjEtQfmoVcMAseLU
3QvF9hD+cxxxJm8FOkeZHEwWOvbYUR8IOwFerJjGMoMytJuLRY6+NgoDDujR7E6n
6Zr72t4DNj/qtjsWTVYFpLu0tJgmg6osPaUUmWVuba+DAT90FqHLXpr1QkKLtC6B
OqZdl+WWu5Qn2I5NLwo0lNCUpISI5WLZKjNmZQayUDg0h3ilRIGG7oK2RAAjGKW1
NM/hlH9kt2oL4NDy6d+ZHFAqG3WnwfSmA7DJPxMWIH4Dimx2dWFgpRyTRAEqUcoJ
fmMdAzMZUhfnW5yWfEC/EVO7kmaYhwQzkdgaKrCglCck6KQ42zG0t6fxZ+dbcVYb
riV6YF9wqm+3MVju1ecE/8SEAOwEvdJ3dftEIJuEWT/vCr2DVZkkGmIaUh5zH4/4
U42V/57U4QAgCC5XmjDVPmtRTdkvljKgzWizgUOqZ1Muh8+UxnhkHaS1l1cYx5pQ
wKK7o6B/i3XvgwXYQ6w+En3LsVUAiFqiVJeiBusTdzeA7aAhz5bvoETXeVdplcdh
v3qvZ9hZCLvMXhGF29dpVCKxWxFMFSsOdU2zHJQ3Fdh44fJZvyDBpd9KvsMUVR4P
lY38qgeL1JPlwVLQUybUJ03703V4LkERQO/5QrvRp1q0XSZCsyCb1jZDW0/CQs91
jpe7vNg7yUiLbsgLL0jmZc1YB+689bfTBxsrXQcCnEb9Uv2fw+TyOGNlRko3FTK4
e3oWiZsNh09AB4WASVAG0lT7wKJjjGl6XG3oApstwwls1Y3S02Dma6pYwEPEtjK1
4m/jZpogRLfGIhKwupOxYUhRJhmHZff5xtVw7KhjJSvGQJEg17pqU6EXzmQU5YNw
9HKFQkMgOma1l2WBws1w+Vbzn3lBKBJRsOOfAC25+GuaoMEPFig6+k35pGLOLUNm
egNdAWB95oWFEIgSkkZcoV0K/NQS49yQXgk2oqO3nNrGX74tRtMJ2ZFTAxd7CQmV
OcJF6250ZUPywCbYUB2vvr3mqicPtEIe4Y5FC+eTPlj44sbbXVZAxCPR/Rhc56jI
4fx7QqusMhJk6s+ip9EaXSnSbIBvky9PYfiCBQdFyQ0CeANuOwad2p8bz7WeDfL5
ihR+TE0Dp/gLBpcY9JEF0sd0ehkKhXnopdcAF3tuWphdFU8rOmdxE7cauL3Zyhle
q+LR1x3UKwY1VVuVBYI2fw6NMMw/FhKVlnr81IwK5ohYaV8RS7dk1juPbw3zElxW
uhPBBhryIyIXqxrXp0pgw5DF85s4nWswBSxDb+s8zSRRc+74alkUlzQr4vzjRqYQ
J/SxABq082gJNCO/2nBQ6Ota3JF2HV1vtrlFSpglRLyltQ3lNkV1/0oh6DEjrXHU
d3Yl/eU2ipEPUM2PLEkMVLudttkHsgcgSjgVEFagKTcpSkBhNtmaB4nyBNRLIIEU
13NUaa2Fei16+BGfIxE8kMlPHxLsgP+wX0eNl0o01Daf+JBzPQYrJbHR3oOwOwa0
4//g2rRR6//nxhlLnGkYyTz4Gps0F/nyJqh/rXIqHP5kCK1a4ZVBJjFEtdjUhg3h
lwEYrcDo+jazlTQ3avVC/vVzwXgrRLGOEjXpdsjQmWTRhZEuwRp4AFS27S6iSGHi
eZKNjNummsrnNsCO1T78CVOzET9aY56cFvrxlJKFwCtTuOVt2M6kVyM2AtMWVpEZ
8cMOj4XGc6gIY3KgphHMDtsY1JsSVEO0cwCCPz2D/zeXhP97rRTxw4woKBKesfzR
xRAIuIJrCl2x52WChYdEb48RYv9Hs/1ykce9xzcPHu7qav/YdyXMta2W+8mBFrKE
n4tX0GoC/XYAflYDZ+5+WA+lcDH6fccUQWEJmoeKUSSGvxMYU7H7EqxhXXgJOOMo
nPR9EP0fhwIQDzOhOh2TwhXzhqfaegJh5fODEWO3HSHGVIPiDNCh+VaiNNnRgFFA
NFF0j1QvlqmBr2YPbwzMH2wozLnm60Mg5jf2OOnpHs5/y2+eKqsmoG4HVPE6V7xL
6TJFInx6nBXzo5+z617+uMS3HqA7v3BBcqYHMsLMpAXJ7kvtQqs5xNtscxm+lKLt
gAqObhR4xrj+aAFKYkpSHT3Cope1V8p3RLjpf3FyflPwcpXwhPF8FHMsRs5oircW
Ek33SzmhbflxHWHf+GmkMwdwEtoTOap+BtBF0Z4AtNxJvVpfeAjJSZj4I/6Zl0xf
S7fLtr9ql89gV03ONOi4c8s8NXDjqvs0YF50ExCZjdXfROlF8+qHDAAWjGqr34sg
GdB2yeQG0LgEhgOMmUJvysiw1FDtudF+kmq7kcoZfLni70kGt25Aq5Dv87AuNZXh
3OR31rG7EdhUX5CPr09e8+119PHn8eNwXjyneM9pK8H0Wo3EZdedF56So2WIp2XR
A9rbd+TGtZ4VZZej49nkEoFxXsOD20DnGNmvzXHr8bJF+nDrH4D0SAKWft+dOdvv
zcalkqegEX/mFUw+KLNMFyTPf++FEWh8Eh4EwidJi/MpQgdOZQ3uPhZI+uj9hzcY
roj/HU3JQDkD6cwbkgHFltU2+VkCOkGDbIAn1m2ltMhLCFdWzZK+d0GwJHtvvYf8
EW42Dz+F6cGhv5iyjjuDhh1KlA9mrM+UXwrbLKU7A82HLSTspBRvGU9b3KZ/+lnG
VvYzIiimeniB6xoh+xyHlgNeKVtq8vb7ZX2JTL/fB/6p2H3jjWs7EQhfqb7VjZyH
El/tZpTjZewbNW7UvkHCpT3ZG5kp9RsK6FVZPXApzKpZb6PIhXCzMfQWW/mBckKe
uyN9KJykx/Q3k/ptyOZbgwHb1J4OWEdMGLZzQ7yIC9A62Tmu4fJXuGIEA+fKbWAB
B48n1xzKFeIjFqcsWPA07cL3JxqAbj/9MXA44QfLZP9o6tgD3qzhHdJiHJkilSiV
838j06i1+fPnbSWKczBnezAjKI68nKHHxIE9AMt0DJ2aCjJbZnHBvUXcbh97yacR
CSM9Bc1wGAMYcLUqAJB3YZJuuCkWAT6JMFe8PcTLmY/yn3rdtm/j6fsvIXDHbR82
vYnrEK67/WiRbw/KWqC7WuWiPe+0/XCskcZfzLFlog5ecIbT+u2Z1bnlqXmUw2gM
QrNF8u3sfQXY/cghr5zgQwYgLYb084xjfQfE6Dcx1/iyM854kVTdxcIoHETxuinN
qVX6M888m9nVnviW136QUZWRl1DHBA8lIq2zf2AOxSMzsZcgBCNt0vPF1Cfg/Gdx
Yl0IkImsoVp/2Z4sbcDuJvWgBp1X0smpnCpsaFGV2MDKto5PmI2bmP1Eb9+/Fw3D
NwDnBC3uUx+OiX7s+WraZWjRtnGvJFESZfyJeiRmyPP8CqrFcgJG/otW1sVo7IFP
HTDFyhUm6jNL+WCez/DO664KrZu+0jH3OZAt5HkBWLl57jLZ+kO7IH5m+GNv845W
4IB35eI+RP2hEl7HRE8EKLU7KJD9d5cgD6Ri0c2NgmE1+Sw2UkHxOjsltMZ92nTs
NVG/uxPdIKVjyc0SnBGjyZC6IgelVKqKPk0wCVaJyaT32e3Q1hKvPR7NycBUU6Sk
NJmFEgoYNRN3StLFHeKsVWD6XNYvVme6d/53YMEDGnFL17PXOjXETXPWgH6xki1t
bSSx5rmqTGEbp9ziDviRqYcNM4Eh0Sdnhu4Zb5GfV5CkT/r6PGk2N9eSaGtaYScb
aFOvknefZEKJvxVplnA1ARm3DjfGw6lsathPSj2ACtmHH1GC7qhGxxefK9Lr3ETE
dl1vr5UamQ0gIU/hM0Vue9YrjTSTnbIjDIeQUi29w+X841gpgO6l/RDBQR5Dlbgr
tpTFKLd4p6XtUfiZSnrsUXGHNwWtgIbQ5tTK4pO14HGbNoWlxOouzVWe6bIbAjxy
Oq5304VYepn0GuaUgaMLL9sZPyx+GfuLTrB+/Lq9rSCLrbKkFXyo9j6vT4i0ntc0
a761gmoH8Y+eFIZzOsWAKsQd6WXAas+L44Rhw9IClgyoDAJuokZ5u4yirpJEZr3d
MfTU0qVbIzBDd68gkwoBf16bLcrZpyeCbCm98Mev4lV6lT85pnOWABf5PfOgeG1P
+2rAcmWv7ymdhRlxz+auJpajvl4srF8iOlVoQ1jL8qg0ye0rGB3i4wn7eWM/CIA/
T5ndxlso+xvxICKTS0iYIgOWQyx+gZTAZ1vLQShrfaY3VF+/LbzEnRa+G24JPhyJ
ka4oxNYJyQ6nXOMEB4taTulS7sI4YzVpnMgFfhD9VcemrzLeFFKDu+zbMT8YSzmz
9MBxksJF7ue7pAJo2PFW+u1Tw52WOL3O/zl79NEBi/Y0wmPXv3iQWKCufskPIP7J
j2NUaxcXq/TQUVMUAGYA2QKNY+28aJihzS1eDdjaf5mMDx2GMucs3cCnUEqEdduT
xX5H/3iZpdr38+s8cetLXW3+YUSU1SYObZa8OsJaPFe9D7ej72FVllNTY8GDEdmt
u6KBhyoDfhyrd5k7KXh3LjjvyRfAPwcuuoieL/aXiFyetccctCCA0m8zgAlo1vnc
zHnVvDOWdf9nCDuloGagNSHMIerRKFxQuCEhQ6Ht71nCOhcvEnck15GtmysFIspf
FrYy4TzqlK5VCx9bu4+pgfJqsPhoz+WS/sYtf7FFozfCIpvumzIKPl8PHMhOHW9C
wZJniDCXwQ1GpAZnjJtzYI/YwLFGObd+NGM7dHuR3AvzJLz9udr5UrKSdP3Yt+Eb
q4m7UQvi6HTADApVzgAc0uh7l/I/8qIq9ZtClaRHJdZiaz59doQhikilHDO7VkzR
jLU1P/cIf2fW3OWHOiE2iqk2ySm5ENYmmW/gZ3EgtEgODqNbUuKIbYaUSCyvlVlB
ZZnI2Q8RZYrlxtv11HKO8LnMsjqgyLg+pDgJo0l07Oxi1zPuuyuO6IAhVt9vpbgI
MpODKTQgJAKuBzDABf0hfKWfvWGNPOA0x63fel2dZzvgj0NHGI/I8ZHzbiGm+7fz
CD/CpO9RW0fwD8cS83CpiIYr5kIzaBEONhB46NCXIxl77yAGzjoKuILRu3kJy4Nk
rcmhqxKnOpgp3dUH3PQQc74uYlaDdOjJCniEK8BBD8nkc+Bt/YFX+o5lk6nQ469h
ahyMxnwTbCMJpVbyAzQ+g642BkbrUAdNYhDJIy3SEJKP6rh3lpffOvPtmIyaONbK
uO4qgVRf/rBpKcWFFlzCdN687PS8xGH2tVSckkCjGNwI7RqJGPJtGHfSZA0ptOhY
hVVdoRzXgtZLT9ihLxdGPHhtQjl7/TDKdn8Zf477xK5t/3VEW/Up7FWID7v5pTr0
isnvDzppxnm7xL53mKaAfkB61OnkSFUOhteAUaIaZ49ojzughEk1+QMtsCj1LG7Y
hbJEvv6hypmQ81dHZTyu+RtfrxjXwGgNUSVsT+lRQT46swdzBIUOdUHG/KeYRPI/
lmPnzEc4ZP/8cl5OIDxXKpi1q2LBom4pBvE9LxHeRmVe6rRgI5Zhn/uv34uY4+fJ
sHCT/KdeZIYM5hjebpcey39AOcmBOMuKBkORvKHyv8PNW2jX9GDiDz3V1kXgM20h
YQufPurViH5CNEF2X1vjC9kfQvIPyrzd7yvhsie7U2a72pRdwP7ZNZPTDYSjoGxr
PbzuydpZd7zmVJf/cRHreck3vNvbQSUVmN7ufQt3RXLaSHhdMIchX4T9RY12d4AV
ihNsDVTCkD6MiVPd/vXKTu5RG/ifAaFeafcntwK9gp8zcDu6mVkbrmeYj1jria1E
AGpPtWbSr7oBa0Q5uNd59HuvAyhw0EaWgY2pjxgunhqYnmBeOG9eBvUfvDKU7vXR
xfBuO+xOeO9xTj9Box+2hXqBP/DC1QD1Qz6Y3yDSNJwNRoA8DyZmrZ+bXOgP58IW
YZNN4I02UBi4tW/8rherghcaMrTnmPpYgg+4PFcqA2Nk1/Lz+I8+GtANEuWZu3wl
H+BtWRT6X2z81H9U/bpqYelGY/GvcLylPM+1IFaIwmquoYyGy8W9msKciUwg/MHi
PTsXJu327bYTdjU4XX3H8vGon9HlhHc42wnFiBmVorvukWhzCaI/0Yi1lGbe2naw
yNoF+sj6L7k8x8J+/peCa96xVS7IP6IejILam/loYB1s3RmmXUi07EJN9vwVmgzJ
evATjiYR0+myHJ3SRo6u82LINDI/n8JQ0gdJDrjmt0UWErCqPjYXGvsn8zbcC5Wa
7ChlOWFg5sEMMDd8xjZ3O7fAp7VJ9ZjDBnybfcufCvuHCVleKIj90uE3r8d9hAw6
54zg+pXiLo3oPOOG7JvxThAlKRJI31ZH8gjOzjLaQ9bbUakrm/asyRet/Y4d3qnh
XtAwT0HzRHnebocwK7olvozQpUtz5iUtiINdKRbfEY4Rk82B7ZwSXXsd+NLMJ3tx
iOyjEdsfJ67HUifb+lvwGmS3NZJ7snXMc34f01vA9pjuGcPjXnAZ6ZwRvkPHMy3q
1dOZ7bFRqO2qdeHa11XZDg7pIX+DSRJ8BDerpEV0xFy4fJe8VnF3PZsdIPz6cQNq
BGL0ypdgh/qmZ9xxQlCfXPnt/y92q0n6WZrqJxqBBe5eH9owvrZcMlCeU4DKWLue
rvIApsYltz+b7Qk+ACC5Gzjeic+AFOzIgrSQYCRf458my5oeKcHNEScTdWDES3Vj
T49dKIIV+QHrSfo+i42i5oZd4ezSyMfZ+NnnYjxmu4176ww7lEsjIHH9jbYzshBk
uNjVvF/mqr+MlHjNz+o5OPIzXv7o5q9EqmpOKkmZcxIaX5dCdvB5x017QdZu+m2+
YeUA3ISmhtDQJJeRt9dph9yS13MhvrKJsbyxr0Rci2fFag1HjEJGEkEX0a4oUOqE
IJXlhMXR+BQSPZIJsYXjPAfthdCGNl6wx/uQZ4whzLFKZ36/SNLFahwfv0LBV3nd
VFZPnzMdzbHOqw97+4te7WxiuHcPJjX5VcZitkhRpWngrA214PNSfvhy6fm3928s
WvmGQscuPTQRrZ0N5Z+5yuNb7/5GrKu0RPHmOzPippO6RKu6hw815Mf4KVaSRY+c
B2DIubjLl5nMHbQE7L/omZnBgvRTuMO3ePXOG9hPiUPNU4M6fXWOxfEuoLDKD2QA
AgELouHfNsl1DtSuHbXfbXQtCsRc+vRjvifzAVmHm53LOwExsYehdAoBP0tlash5
YMtqxXzBgHmUrnoCXsSdmh5wWtR0HyjH9m5nxzV9YMSf6AzJpZUJEenv/4z4JwME
tMGf7D0kEPebKkc6FgmfWPMW1KthTFO2mQawjNNYS6NlLk0Lv2krjEt8+4TbuWL9
eIfOFQ8ZKMROvtAAg45nGyVAKz7aYpywDmheW99VgDzblW2DhH1N14xm1Ax3Rtwd
IjGGupuHhfw5AfB9lGIKgdp97Pi49Va/4NyJL7ZFvhIB+6MLPQ1N3eu94pyHZVND
41GFxPLIkj8XgXM3k+a1jhHo38CAjPQajBNddKnETodQgumdQ0ZVlE6Sk04IA8QB
FeDyz/sATBNoPUvDPE7Uj9oktwolnEd09ZlMKkfrgE2W7RTGRb/mvJFB6NCyaHB4
05ws5YtpZZbSqXbK11hFMp9BCtwxg1bC4nh/AIFNul6Ij6pC1ofzOJShVia1a58p
40+cWsRzqifu60VHrCUxTvgyBhRxFc69hRz+FFwHEddq0ISVF/1PnH7XV6agAd5R
8mc6VqYfFxFfE7HnulG9VpBd1tASwXzk01hbxCe0Oisp7EMblRw7pgP7Mv+cw2yZ
qkGYZqPLUKx9Nh3IX0neubIlJ104pCHOmKM7DBNbJZoKyqTfjzMyZYuc3PiqNl5z
8km/Yf6TkEvp/o0Av41WxXqOWMOLiBaOANuYqf+sL722HtcmFFBHXzoE1x8yJDr1
w0v36uK55gQ/+7uyBYSQWdYi1/X8GOGt0W44X6GdePCtFR4BQImO3wdgkmkSsnoF
d2gH5ZODidGnPNpSXMlJnEqti/psH9q9CBqmdLiMgLGZUASbP+AH9Gg0LKJkhENy
7V7AI0owj3t14FLkUiMl0Xs8Q37ClgtzXbSX1H3ze8/yiGVM2COiXhrD7w7nBFaK
COo8w1wMHJLIcx1rzPjVWJcPqEKIW2GQvUQtO42f5VI2KE+LpfW837DbqK1EkHHV
ZcS+wvwdrpNMRQdaN1uB4M6mGu+8/9Qe3X3WMAJcBPzvM8lF98tQxkcS/uSxwrjR
sPNbwaa9oL7Kqrb30WRkMfaV6miaLHNM476Yv/F/AisXqPKM61mam8x0XbyeNTzP
77nrjTTVHXFio9DKM/zWfCeWwox+n9/5RsTNGWDl1sodAM5t8MEWYNZS1blOHKiH
vt6wu84GItvljhXiOoJ0Hol0Y4o8gdgo+NSfG/Yf4H/ajKQrCJgNI3Q8EE/BPqhX
NwPslL1sgBrXfx4ly1/Km+/j0Ec/lFhCivzS6mUtvz+pXWUmP4MGnhxHVWTAQ5Xa
2cr7BHBQMvBxYw5q8p0XUuXp7PnkSpDQ1AbSsZJfOJI3AxI97mRLVW6M3JbSSXlX
UhDZh3E+oahc01nfuKbTaaZ1P73UbI94ilgygtpyXk0JCxsLthVjrXdjagyRATYx
zKo2FSPMQZ4xt5hCsfZO3+J81ZqkmWGBN1Hl8GCiERnduTKJAJ39O+Xmkiwnot0I
bWtMxinHmmmtPHwtjEQKc5pM4mjO0FBMD9nORePaooPltFFgczl0z5EMMYefM5pw
ZHezV01EewIlNlDV9BV2rKcECPs50S9nighb4nNKfdmqYHu3g5GtZrPfEfEo62zw
wJesDeehIiVCZwe6vuzY5Jj70tpUjVj+brUNSdz3NhxEMHvhLD2XRs6uK/Txn92n
6csquXvKU7opQuuiJDWVUzI4m+66Vhb6RGhiBz9K5un/2+dv6e4Aej8WRM+bfzeW
iq3MYKYl2iF8PVnu/ZAVHLLw/K2PvuzbNLQgWgkzAeCFQbKB6KPy7NpBxIUQz0EG
zpEHGbk6Lz7vMZD/0hxJrLsE+9Sdjehp6Cl5DqllGPmz+Ojsr8Bt1NF5/CTyMAeV
3H1zpsltYbboJeYzQG8uiUVfLMF+e0rDM2wnvBSlxCgt13YNn7KRIefZLFPUEp8k
z1nkMz6UL2ZVDi5t8MNPXyBeR8RayCAuULRU0QhQOOzidK8Z024FhmeOeaFStq9T
Qrs4c3U014xfnw6dKp0hXtqAn1APdXQBMQZfA1OWbMDLcMnjweNmvnVYTPg5w78c
d/3ekSBuH7iXI/Dv2Yaje5WYfVHqoG1JZfRym1i0YNkN9qI+q8iTbm891M1M5rB2
LSd74VYaobLRH+bIjDDKjmrE/9pB79mcz0RJIKl0Zqujc6Ef1trs8ON8WfLNhfxG
xaTsNB0w51t3u/6QVmbE/2Ov73u2t0bSdI3vwUFK3XvOETt6kDr1bA5n9N0MYSa/
fMCVXftToaRUyXMbvTrW/vHQYibTFgjrS2mJuhQ0AIK40hOWNT1KR2Df7yal89SW
1f2E+JnCB2hBw2PymAoJi6bAZG1suVX2CjAiKFsysq8Q8BNynbAD2uudGaH/FLd0
hxJ5o230omjNUNWplIBzutF+pT2n+x88IA5wXWB0nilOF2ewdyC+udpWTWZ4DBSR
/OP4mWr/kvddQTTkNqwNwc4eqYC74qoBOIEileKDRlUpveh7SjvI6h4bkEEMnHl1
piOA6m/pPcUvo/DcgvgXG3O3JXFPk2J89m4+Wf1ONc9hLexiee3ZaUBrsqrNw25V
THFHeZ+1IsCVG1gCgmaSdNOzLDegr6HhqYLq1iMIxX40FEwjUtnvP377qtP89Rv7
w3pBEQb8wIFkZ3oh02UthpD0Ek3cVquuKPO46m0ZshgTNjYUbv+x3QYzuNwiCOVj
whdFKvR+Sv2LoXXrZKDYv0bmwgW0swGhvjVgWGJGHDLKd7hvfhfC0LIthMbX+Wqt
98JF48hUvow6kyvkju9leKBZrQr9gkrJ4ZNojmG9QbgRpBhI3Es0KgiWe8d2d0TI
jBWNTAbw/LmcZC0X6SqfvJzqcSjto+x879Jna5dHe0lBl5Ni3znB2ASaOTZ8g04A
POmnr4Rrar8FkCc5llQ/jYtsywogtArFUNWugpwv8XralPq+pCB1NvKLW98kIV5d
p4Y/c8CsKJ4X69lf5BGbcc4DZw1zTbJagix5fd3EkTZbe3bjRr1dcgUJ9Ag8BErJ
iI8fKiB9VQo9y+2YtBV0bsJmKI5psExv2suJDK/9IUaBWk9QlCYEtb845xan/e+e
C4pGKNhMV7padT/z4XbHu5s3O4bFUepcg8EBu4/yIhC+B4RcJOA86/jR4s9gi9Jg
8JRc8L+1TKUZPQmV7hfaDup6fIWVihvCaKsRep8j+e7Bew+6ujcHY00t4ysDB54i
R3XfFNEDY/26WGFS6uFe2fvxKYM+pNDtEIw3y3aw/8I20iMTo9y1c8zTBHDbAQkq
Uc7+Q2b5uUQKuPPiggoiipGkWqW6T7C5NM+nEDnvfJ+9vAGIExRpEN921qn8AxMV
amnS4JbjnvU19KDLDBzjNo0aO8PGAlXKWfSHu/K90zm9zBQL/kGPVWPlwVFi50LD
LnyLrtDJXsbG5ujvnnplwnPYS0ruJ3PMskyBRIcnvC7CpfozQnBcmzXjbKVgAYVO
wpJEs8RNlHFCRtPEE5RoICL/7KTVxYIz2IdBd3oDqQUkmL2O5np3qXb+jMbMaSAD
7kOHn2Glf/8sKlikZ1Pq9OunZotIVngHVp0mWqU39Ae22V7u/Ovk6VgqeCt/b9Vh
F6g1+XVhVXGMofLMPuVzGKXq/dM195t7K7aZe3DpklOS1erZFvCLQMNBTdRfNOmr
+OJ2c4zoGWvbIQWgrJGcZI6exQxSYy7WzFc9uoP0xuLmER6bE7N+DuvuaN+s7zum
orDO6NyiD5tPfhkOuOzq4Pm/Z4PkOtaD1vxV3HirMbWTyfDwk6yG1+fYD2o56UBL
9Ozz+VjHGqvxjM4+3JFJ1cvcVN8oStm6qjQQCO1t6rOAJDwoQgQGllG5uZFqe5tc
grgwtswiK4hoJJ1WSpV34hoX+axsY4qQ4HLkYvBBKfaiGy0oWPoQP96tH6aBGMhs
eA2E7zB1xdI7ANpm6miZBeBdc5FLRccIRKy2dWyukhqFN+gL6ddrDaC5b5THAX6w
2A9yoby4s4CpM6GRfd83u4Yyc/7x1CbaCILMqRLy6yW9fSOYUJWrJjISDxDQnaWY
nepQputhzuzQBQ4saaRCKKA+spBheRKWhhY7Dzg0BFmGKubRStUVTM3K5Qon8uTH
gd5UBTskaPetwWzCke4re4oR3H3scwZM/FDFApCUzPbDAu0nCFjB92ZN7h245B/U
n+rigkshjKjrbUgLMlNJcew9wCBoXpfkOpu8H+AEWWdHWR/iYBSsHaW7aGQUlGLH
en0Qnd9Cjs4VCRpscxt+OEm9PALk85xh6BnQH9NyeWQfmUaNtOlKYk//vOq5KOXs
6r25ErFEnUVD3EcCaGv7ACnKCtC2Ru5d1p9yAVXRZ7VLhBMXYokE+SPzYJ63Q6rV
zfgmaSv/pVKUoOgJfpAGDERDrUT6huysqwr2ZbhuUxc7V7ZYq63S9gBPxnGbrCt4
2S34td1O7DZmS7JEK7ghkl2+Qb0NJp5s+aJ9yiDGwJmP0Moi8Wc4R2vcAPijZgug
IR+EuTsmzlNwWDBlf6b7sf8vhKq8HiNjftJ3Y3ji3V2BUqBrQIzz2TogU5Gc7FvX
iiQ0A3OP11u/B9uO43SoeNjpm9HXs5jAR7VopLP5P6zpE2Ie0SfA3VAgfGRmTj5Q
JFyaTQk0J3QGyQgl+vCR9SW73BJwNED/PUV0Vqzjaw8qHrkUIUOyq6I4MIvxuGU5
sXrqTBWGgEb42gzNSTbiLl0pN97c53yXbGJCp4TljZOHpGNngSJhvBAsS6SJzQb+
9scsu3UKJ+BA5Yqsxn4S/ZwR6PrrmholR41atcwQ1s121DUaJ12fKeUgI6blUgHj
ybqwYfaF7T2TSuWIr3apEgbfkIfGUshIxiBBvrE5zyjkRIEgVzP5s7ChqX20jCDj
7NH43MOATyIcG2sk7TgRApzvS3jwu7sH26He98sfUGOeK9j9cTA1tIFlDYTJlIki
TlUHUBQdXVlxOoWQOQ8EKqTkuBYQZy7qEdF7NtFfVFySQxjF87qnirtKKo8yBJlB
3V88mUKlAfVZyG51J02uiurEb8dxc4eXk8uAGoF8DJRlJpSqJmpYnSbQk0DU2GUI
KPtW4mZSqg5TfIt9R8h3ca5SK/PZJij1dXKKJ+xwH04u4sW340uXlfwCrIyXwCfP
tJlWHC1fS4ld/tVxnmkhqUSUzslWYdkJKRehfbskzVT9QQgTBVPeoVoa7ee7H3tq
tvU3uifHzpTTsTM7SE1DFM5urCemoslDRxw9y/J4JoniyQMtsCuEJMddmIm7olxY
Fg+LY6jeTLsDcqnxbGvbSRdCFvbVf6Ze2BnB2l31vbEw9XPI+11GmGZ4KkJj/O7e
Bwlw8Zn5a78FCLg/q9NXpbd6HVi2WSaHnEg3R5SDTku9egGpNRAiqv2J1nCj12UT
xBQMGXOkXNxTQ/qWpE8nOV0iiOOMXFzYnvLs+JBL+0qTom3gb4mB7LEIpN/yAdgP
kLM5J0qwigZ2TBfqvliCj1lPDwpbZarscvQ2w+SBh2yTdJg/WJVGZlxhoqG9wtiL
sKviZJrsjZXjiJl6H5BMAPbcYUuyecpx3ClfHXPzkfuA9Reb3iQYWeujEbumfDlQ
FxlGRlIKtHOquVk4il/+3vXmIFPS5IRA2cYAjdzriTRZyykmiRTum93s4jYw61jg
CP0K5AJw2EXRWUwQJ4Uxke+D2rXCGUeIgPf8w8lY24PN/ssTxj1Wqi4vkcIi/03J
W1grNrpjO7eIy7K6Ja1+HiTjIvTTI6cWge0bZvvGZzGL1uK+7lzgG/xTdqv+DJ7a
NNB71bxWpitkzjRE7FUax5GWkiLxY+LaUppgnyE5fsRkurkSh4H9fEeUVLXuFc4W
PRVkL5O0DY933W5tIz3DkWhvOvBcr9hqIGZKmN/1pCIwL5AI0FDp8ywwB7+je/wT
vnvT7dCtoZ1Feki7Q1yW3dnhWP0kxY55mInw/epgmf1zk8+ttgSB8qqmsZR6QoF/
0n18KAh1GhXxc+Hef7rxayrOk1Y/zRee8br/TgFUvpSrOKYL6aQQwH4uQnutEOga
v+ePrlQBTBRu3GUx8QyIty9eBvrn7BCoOAr5kS04H/UUk3Y+y2dXK7VXA8zE8+7t
/MX7CuAVpVgfHoJ2ydZ2/tfN7yfTYsX52O7CaULdLY5T+uZNu33YKYlp/FAQCFH2
p8b7gTsMDfHKcDYRvQO/S0yu0j6+HHQi/flvVJUgrdNbLabgQ+CWIot0XcHmvShM
6L/NUO1sRlBRaPUAASJIx2dq+XY2pvvIXKqrdLYBBmns06W7j6H2dha3omSIaMBd
Kpr5wqbgyUO2u8cIZF1+2m0k21kPo//YCH64SU9GGWx2X+gkQDnXgY4hfvGwN+yI
T6tH07DU35QREhModzSaJkCzLOqyn+kujh7526bDh6KBdoBieg7yYZaFrz74tbEz
V616iDFmtS6YjwcG2x8oSQedhhSt0st1XgRdGdFFx+IOUvqzth7LLOPCbSiV5p9B
zDgMCVtbC3b0wZd6n8Oc1gwubb/2lev1HtPPxraHw8Bnoek5NhKa3atooeEPCSO3
Pc4qg6GjdlNC2Gu7W24HwxcskmdAIEyWgfZKqhHPUM3htVi5NyPD2Zqtn1FZS95x
oRx3teIw+L4dZpFFtbrPCFy1bQ3s2qVE1bY2NSV4dho80H6lseOKRF7L6cYrR9BS
d8lg2d4ActRUbFBhZKFkyX41UyTFRr8wPo9SBIgvh3rK5nJdADmgO462jEISJmka
mQdUlR/LFuMne0DC7EqcfjiMhLtYtmM+p5yaPPJq1jzbgbjxlCTucnnHAa+P1Xd8
XTyw7Qjl3DbwpDxJAlNq3NbuAxdnEwGRGnjiNqdEHAO3HAjJN5yvtX657spdPbKf
lSg74kJpqdPiZJw6dcGsA1fWnLLYJTesTMF2bjJgVQvcn6ykVp60r2agpka7hbVT
LjJ/GABqYohAiHEdFl+aeXzGRqHnT1VqQThJnFso5JtjVC3y/9gjEoytEwmMvgmz
D4a1swwHS0KITsMa3Ipp8/3gU1/sMXaEH+kUvHdtgeSj8MCxswy26KxNV9J0lw6F
6MEb+scIY+zfGcKxLDpnmk44Ul4fywhMPf7T/4zf3M+30UKIIIHMWfvucKmdfVtx
UcK8hvC4jLN5qj4I4zzvLRDzFSWEhanHmmosGHd8GLSPwPqDTAGWW/wCbdaifJTw
R8GqHlbttqjuOHcRNtp+dUjQ4AZ1917w1ycpT320jkrDsr7sMjEjr3fBVSP45yzX
SHmQ65NAnL0G5DSNCHczbJTb7r2Lwqz0rJVCyTYPSU8zgldkcCwFdva3MGmHqjYj
5XsljAs2YRmm7yVjjKm2JXxUSfzb+YvfkyN2+czApqxK5Pub8f+nPt8Cj7N77xH8
QMHB7euBNeP079l8lYhQ1r70AlYJPYUXfZR2lvzkQF1EdoDrErDl1eelCWO/w1ji
hkX5jw0EP1FTW/vx4Wv0IIr/1qaCKthP/Y9lGLywWdfPJlwpbOXH+1U01+GP92EB
4V5RS3lH8eZComtOuY5kaG4tdG8nfK4dxntdQGuhgmGD55hNQIkC0bcbNQ2a3DBi
LexixRIw7NhF7hlVbQKVaN4rLGAwhI8p5GEwpP4MUU5049wDjCu2dq6eBjfdR7GX
oMhjTrCFvu25s0ul5QY8HB31pYGXBb2DgBPq0ziZ1FTAK2yK3dASw4OTulQCQd85
H6MW0740ClBkkzbtg6g0LW+haDzUoeE8d1pxzJGpFKtbwR5gjK0Pvovo4dR045Q+
MR/w73OLGmGqqcwEf+bmrQSObt9OjTWlD7X+M0n39Q9raEeYL3EktLrvezUcofeh
ynk0nptzdAMZHWD/Kv3CMpwTGcq3Bp8sTdBVtct8m5RXfayQ7j1SAVTlUvot2AU0
NC9S1h0Axfi67eCL05eBYkB+3sXQPkqbXwIaOMmYQPUQYSp5z/qq4iLwM1fbWKg5
vMbgjIpo2HUoNlwIOgi3U5kkgeasWqDlVL0W+Qi5I1LE07Tl81zjkUMwVjdnefJI
pq0Uur+cAOjI8OdjO149IWODLtEAWbaDp43JJHo6jw5GdP4p3P1LPLMey0P/m0Q2
6Je4F1WFz+qtMZziNnPMaAc/TLyI5njRdUWhx3Sl9wSoohCHgo5AKUly5zy+81NB
hGrJbKJay92OIV0O6cKLBzMvK0oFvns/+skR56yQaumUWrsRrc2v+wGT0n5QJF15
pvtEDoVouXVSTcrPj0kpgqi/QconYT3ipAef1N1EcqeqxEtQpPTlrQtBRvaahh3B
8KivHjS/pMMFLeaq7LcZyaspCfUZnS98HWqrX8OP5RhXeC2HMCoCQSMYTBeiIShu
fA75rtFePrXu9Mo8pBvVGNtdplOzmB9ZqMGyv43lJ1X1cxCY1gFT5vfPULrlMtva
QiRLcEJo7yTgnyISPKCsZY6tsAzf1DFH799PrJoq+HzD/oo3haDO1N4GmJ0O9ryN
W3LODbiuAi2i054VCGvdRyfvgASlkACt/CkmntufPm3z9tj4yIp7JAZb7VXH9tjg
7YFq+TbtZk9vf8PPlzPy7m0EcVk4jZ006H5Mckr7LbxRH6EbilC9N+1Piiw5FySI
r6vXtgcyo88HbgnqUP9xpRknSsX4DQHokjbuIrzN+dHNtDvOxl4KuzzLxcnPcFtM
n/C336gzc5+zuvcK7FF1G2dItOZD9/AB8yG7ZBafqOkxAP09BF8UbBqQzlijwRO1
CoLuggeF1DR4pewTLznA2YwsuRbD0l04eaQi6f3epvS04nfNCdfvRjFliK6payy3
Q7E/GizXuitvoOsle+O7B87UblCP4ShGp6w/or+BtzTIpJX3zi99wmrcgTq7TG2L
T0Qo+amwQqIlILWsjBtzGWtPKO2ljcC8SWEGXILhRKu+beXpYyRDNZSE0348WlUc
LZ7tKE3iE13NEjOvg+E8IVbyOP44enISlx2Wxav02Ci9xGCJWDaIJDfqNAadfaYu
zXLaG7MpGUoDMfR6PrhehgiL2HeZW7AN56iGqQfPerfuMmxiB4nmGPZ6Bl8AU+9A
38D9CbTj+fPi2BN7M9wnMye8kJo9oLMCDPfcy03knIV6aGEOeXNbweHt1jjZQyrL
vHfhIs17FkRXYB2kwXlsJTwW98Z+5IW1i1m2SjbVNRnXOCDhvaRGnmR3pJCGghIE
iFuR2qOOCaTKg1hwlchkqRseWm20ktgS8xq7EtCC+bTewV50xXSV2VWcJjmAftZQ
95minSXiUde6IfYBxxjUBtIxMxAHOk4WdkLTfWC0Nj4nJCYLUjCPj91Dnw55i8wX
4IGKfJVtV9eI6bZQ2FeDKQK6z7pp9WnEqQD+HMqhAw6T+vaFfVNINuCiVo8NQSG2
CQPiTGKVwMJ8Ba3Z0+lY7YHVMoWpcx0bhir4NQXTH/kyD2yGwJjUpxC1eeUlGqaj
BKKaAft5Kxnk5eiuDTdDpPFJtd3JY85IXKtzgqWs0zIGkNkPRcGcsB94XQZnS4s/
GxRcoZpytBuIPmnaqDMOQ4TIVJf3CI4nhe3YEguGsghZgKNsjpvKWpHEH2wUUXg4
yNN9e2ThUub/OH4J5w85eHUJtrTENgQ1McpJu6z03sk2k0O8n46oBGLEv7jV/76g
Hihmf6bwB7YcFES+fVoLSq2MayZayOExelo416HvizX4MxXS8aQoOcOsvgIBtA4l
OMhrHEg1mfGhtgyxO83v9AtkC5kkYEXqITEAh7qMjNFvPoj1E5VPO1+3Cdx6lwAL
COTrfIC9caiALuFw14STcpnlcP14VR0lPjq/vEkseMsKko9AdCTa6hxvXZjC6+Wj
I1exvnSywhLU9OEo7Jrcf6wLWpqSz3oapA2EEHnikV4Ni0qOKXTSxTZyT55Rdu1P
hHY6Ags7JVuUT3xKstk4GNFHfz8KIUh04Kq7tnlLrBasilbVMmluzZzkZByuuUEe
ES74uJ0/7WGPosUDiOLC3VRj2g7xor1q1/aGmEvqYAYrQjQQHsI+fuVHj7/jCS5p
PdIGeYDDeeydZp1tE/ziYOHIn43zv663AEp/lxxikD1caP7DAvNskmRlOpi/C/SI
3kgnQE3DMNkCfYuPRceywMkzWYdBiE3O1Vdj/EbnEJg49rudXn6iTMInnwmCLTop
NPfBuN6t1FkX4TxXWRv79vDigGt3M4HuUBHgGYoVReScI307OuZ0HdR4fB6anNI8
3RMF3Q1GiVZUYNrMMkA96u/d1ZiSArpJGYgUMvF4wRpgg8CbM1TlYp7VLclafy99
/y098BK9LMoMU2Ch1HC32PTlCMrJ7JDUm5eimqFryZkglwKEkOUVKKIWX2lcZDac
lXAlaGHv/vPUtso1SVVerufdOnoF3JrMDH75VFIa6p/31TsrabMVXk98uqIFpka3
zry3lGkkDDm5k9lfN9OquF4+NF0YB30s0oF2w95onmYkoEIXo3fkHp6N0FOEO8+G
IY9WN9QUzPVCGrEoMZYJQ2gl2N+0+qvWIj//BpP9nw+CNYleUzDg8fhLYYTnwvwf
aDy/YF/Qm6JeOkf9jqjIv5AgQK6S2umtYfqBRkQgRpPyaVTevNXd4VeJVvVIhCrv
HKSFqYbNgiNw90pAcky8j9Wp703Dm4prm3MR3mjM9HEg1h+G1dcb94QgIIpJhfwW
FtLQjw5ai0NYdN+LhLQrP3KSGNlVQXqoWF3/lYVIL6u/L2/ssX+Bjb/+KANDUlbh
l3ZZ8lcz71QI+6PHgjMkPItoC7V8YXKhjanXK4B7b6ibCHVWd3CF0HtxkXDVNY6K
Qb3VElHRl6KcgBKQojVtyRZQHDQNggcLtW76NkVzC5c8bHwGx5UgEjvK4Ho0Zrgx
FQnrnnv8CKEV3k7PhxkPlANRITuh6LweW6Mj1zXAi8TTao+U/tef5bqMSIZ7r7N8
a6gXaF7zk/OsvVOIKKhmay4B0nisQPiniuEF+HVVW7ZwNA3YjsejgChCkHk7HyRn
vy65m5wwZOdXDDWuddffGnywGr0nsVFP1pxSzfuWrULF0fU0HaiEW7FHKUKH4y96
EF7MXqqat+GuB8kWY9ZCk9Ii81rbu9rpq6sCr2VIcYH4mU9uOJe+J9ewn7eANR51
`protect END_PROTECTED
