`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0QPMvkQjWf4GgAQEExXJa78qrZ5j77tgZWxRIjD+J4zXpD2I2ezSaxENIDiTCeua
/3S6n9ux941RClMnYRUk1So8Q6qh010qzfGDEXaqx6pe+u6ggTeQjXdz2sNwKdc6
wgxGPmoFZbCHkCYwqo3rkEq7fL6HxiN5bHGr1FmlEvyVxWcJ0d76hjNBhSCrhCgx
+DxDMegvL9VV8226MFkF0QiI8pb6Q5Dl8SoODa+mfAa/0Fu62zPZjMsSWFjyh39v
b27wt0Yh0m+XGbva70LSrEFUvadsjoUZpa59POlkhxS98W7aqgB8fzkextGV1m8V
O81/I7P69tiu9xwuOS9Er6a0mal9zMEmsoP50PIlG/kAHl8rah77DIgjbl4/U3o3
EYAwzdVmDI0gsOFPurdssBdTbm6rCb3nlx50e60sY3ttMkL6DpWEK4qn4vQbJCpu
U771TtdJlzBbFfr1gmCkxoV/D8NTJsLeqD31XfpFVCqy7QzekjGXOqEQPox5SxjX
wiIkTxqFbIpfscDwbIxGB6RcppKzblzAqMqWd78HUImK10os3yxvYjzlt4+fkLdU
g1SX+TDty4bfRHxcK5ZgkVdDl7reqGdl6jEhoCRGV3QdSLrG6SsO3kEE97tRctW5
StPdlnxLPsOHq6FGOn6/YmPAvkD3DMrsVldZCLt50ezqN3KkjpK2rywU2X1fdnfr
TL7WraWb6Zy3Yz3n8ZjhqxOu89WZYmPM2osm47ocRQQmLrnMOwBZHLZD/lvuckty
6yq3/hNJkyodyzN9NBiGB4A/ItexPdabaJrl795ROXh/16jqyuIg+J0XD2tGdi9Z
FpJVEeSYL3tFoRCFkYwVWUTNQK9ULW9JB2liHdoIZ9fh/uLCmOmUy5iYbfNXeC+t
jhK1HpZ78W8rZ0jxgwxgHIW5ky2Zaz/7gfP0lXq+YbwYHHFFwmP2UYyciLAFAsNg
tahCdut6OGzOSpnl/C0h7jQP53hyCYETZjTNzFzQ92e5dFBd/h56rIcvW2TxQ6fj
VMuzoUd3nXcs/PRMph+5JFHE5oHpYnf4PsnVwEmkWSkOVn7od5MzLJWhwBonCiCm
sXskkzZoB8iLSTcg5v38rRi0E8aBoaT0LoG/AzaI4cArDvTD1QMRP7ifQWkVwBTc
iImPaXomtiZzm5NedjmXgeGWmxK66q5c0Gi0qhH7ZqLoRGdGuZxadfrmFjvKM2tL
xiOitG3sYRcWwE60il3KKFoHQ666XwQMxPxU5deZILrKKkeEmQby/Kq14qxBcsn0
4UrPsVBaG25aetj03sAM/E86zJ+v+MnzxZV3jgJepKTvp5GOmWqfvqf5mh+IjWO0
TZW9BnqTOLBf1HDSJOX1aOcBlS18QkGc6yqK24tRkDRYhCHM0+e4c0ejw9tVTGyC
k056uNu8De3PrhS2YWal4zFJ7V/Zm4HlqI0vXcOdY+bQaW5rrKM2JqibS6U8ZvBP
RLuORX+SOFHKfQ5NsROMY/MpWOI7ldMyks4xa694QEuSDA5Df/ro2m4pU16URYYf
+w/BO22thvab9n42qWwdmD4T9l9WDKs48Z/SofkdhwtrwyORuIqH6+1SO2Qfp56H
YfvzXpFpQXj8PqpMGXtxtU4X5tlKkzC+3AtFIiD5C0jmejWRw73vJOHJXkeLF/HS
Xvo8XM65EOBlOGBXZBKM8eyAAp8QPPIBVBjevnKRlKebTOExq1oSKI4fyGvAP++E
ANoEup0WsN2W2pNxsxO/IWQczP/aurCGV4RZJRAzMIhRbjdgFVQC+ibOvbU+LUwq
z/MiuJv7PUXoypKEku0fP86hrC7hLIfrXyfWvKMELJWOZRsMcCN2m6lgjxeo1YFh
5loA59DiQVhPJRRDfCDV0BjBy9HAdJmANlra7CzPcE/0REIcGBB0wxCeaeKDHtrP
G7Dhclxc+VbvoOWm61UVNUNSSczrEg0lLzHl6LbZcGw9jazh78D44VtepCS5nwIM
wSNGSDf7sGLtdX5W4y44X4QjNtfLf5SYKBjuGIvcuL28EuINbtxUxn2+FrHC9Vak
OvKH/0cHvVJnQS78Udb0qfNhny3uJBUmA/kTO0QMXDlCc/cltef48hr26LqZG7wo
EnTgjfuuTqYRJ9YHHX2RF4YRQhTqyc8qsQ3F0gUs+/OTDe2OsAcS1blqR3Mx06Wt
fzKcVBzDlPVBJtFWNKWJf9lHNi+EDtUO3O/Z4BSRjWoSi/mQY+5iNzkD2Fuo/OQi
lVcoTa7458lyjrrMtlxPuFr0fJU7iec6VyAOc8G7HWItP1iWvPMWXeqvk2fGTPlR
1dCH2NXuqgmCI2CJC0qJZFQF4RlYQT7SKiHSth/fJohsc8rD5P9zRv3m0KUnlARX
uDbDh/RH6SJa/E7DYMU3+hpd0X/y8S1if+IUYpdKVtlt6ZdbKzNnNoyZqcFCt1aE
CQZpzCCyP7+usskx6RHe/umdur7JgYNj7OvV8gU4e3qAWDmAh60/UCOt51WGYG+G
XJWPDC9AoRK8Pgg391VzxqrgKFZSO5efPl5q1kwBTC3P+gYOuQiuf8CSPML2dVAO
0MG20zHXPwSlh/h6GXH2kyenUM3NMuyriGAXbw+JFSLI3Ud8szQXH6bhhnXUNmT0
53iePylqp+ZZV/ZeXt8AqN0qIiaJqauO2WCot9l5CmLbQr2fKwmdL8noRyN+Kkr/
M4vWzMAhLs3xf7uGm1uXu9Ew9TRhlerB5xGLcyD7PmMKDRXP2pBf8ly1TGaEHuGl
+M2Cy3qTuu3G5+o9n1oxoO1ZaCu0zjSzCrXKUa4wzL2WoeORen88BQQzJmmNCtlC
iUC7TmbTjXu/R62Xr6px0vKL/kPaMh/9sQBdHOxyxyggXJmyczwt2/+yIvAGCqFi
++0JnqCBU29XtCAYu03SLd/uM5Wnjav/QmSDbUl9IJX9CZOHqxAFY2Yp8zIGjsOs
K6OI3Fz3mi41AqRd6+8nd4lcjzwCToOGjgABYKch45Hlpd4Q9vcSBR0sF1nVDFrU
Ff9lx51vM9INC3N2GlDXxv+h3fAlK3NlSv/JZCnfwrPSlIjfikksKCPTtq8Nf26u
xJQgdiVLFYF5WvRbfLnK9dbkqXpT5WFrqY9Ap19mjwB/y/TPP6WvWmmzt8hRCTKm
xTc1CI3KrU9x9OMMCABzHcdzPOZa1EUXel0v+G6mem5GnY2tDo1Yx6vPsTyU+ymP
fkpPUmScvTcWv7ly0j8Wwrj8nwxyA4V43tOMXiw3lCUkn6rX4KYpI4VRlvU/nIPl
SQWWUjMEakObLGEkBfPhzJV5PRCG5j8iC9hr9EDlfMXBRrUllVm21Fm2G2S9sGGw
qFG4wv/Nu41UO/j8o7BsNpIZ3fU3sPWxbd+UlVGs0oxsZFWzfKa6M4ZhAlZwUFNl
s8+oDoDir6QH5q1MU8Ms6gVbgEhXEaNkNYxP7fl0FkmdmNaisioUKO/e9ij1PKa2
KIf4XIgZF2DHPG0u/rk8Ky1i5orfHgIfgMXPbiilkG1bNY7T5y/1FxWmtLYcemBW
EDfWfUW9gmZOBI4sw2y/Ge8K4Puktw1OXnIduJvZoEw=
`protect END_PROTECTED
