`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kbYmTAUM8cc90rkQb3hFT/K+2MgXvUe9xwSkyOX6aPNKTFWfI7H3//5GxEQfb1D0
xZyXw2+T+cp7a8oB8YtDT0Ykh/5prmtEuVGVZmTdisio06cVfT1ETFeGJSlZgvmP
Qcr/JjZy1xaVGeDIMIExh6Z6yJM7w2XNoVcxo/kl9LxFTYRzvXnq1PVU1s91BEcS
JMagALtbRb+ky4N/rdkKbc02y30NfRBjcl1RiKfj7zVcEeQ8N7kTYAIjQpkjNSFO
sWyLcLmXqeZf8EuZE5F5/euxaX1ZOCnpMTpJb/ICS7yi4RN1m/lGFsAxaMByHZH/
yq0sshYBYxXme4tQUvWDxjnQX6LbwUPfAOT9niGM20PrYCvnoA/aZHPeKUepbgXe
xJHQJc5FRF9CoDKj1pdUzjgRWEMZDCk2Se7ZtXnS31+eFxezMohQDOHsGGP0T1Y4
xLUtAlSCTQpJO7ByvVBpNHdjsqu2qdb1DqpSPMzcW1rhZplcxwNR6/ZQnu8giEXn
YTvvzHPIjVfnXrd5GYfxeg==
`protect END_PROTECTED
