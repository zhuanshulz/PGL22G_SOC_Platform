`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PPmudna/ZIPBijGPPgUkXr5m7Ok1RVQyzJmTxB3P0Zgs3wIcde6/mWi1Elzr6Tsb
ufbc+HVyNShkn8CF9b/TeEuyxCTbgC0qx6y34o5zpt5O6CNCdz0wgVzGgK7UcP15
8u4wu72hQkT8mej0s2tKMAD0GLb8pRksLsfNq6pVCRJtGhTxccVkYRuXgrlWVVXs
L5bkfBi9XvpKdZ32JLO3EUWmwWyW0y4xyOPA4mfSZuW/m/I3f+U18ZxZZtqCR4PX
ZNjyKEoimXEsoVRFg1yTpg==
`protect END_PROTECTED
