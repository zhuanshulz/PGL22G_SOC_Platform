`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpslK0eWo4QFe1fReD9EueswUef9utVmQMRbahhRkIjtHhL1hpfMy/jEUCkjgHTd
d6E11s41qeipipIaFKnj15o6Xykup1JHJ8pZcsQ8eHZW/ABSteoXtUtvXuUlQ/mC
/EnEz+pTAfn+/MIC1AfQyPU5D4QRmj3a6VlX/1JzXsnFFZDZi/KIKDErLYF5IUa6
Y2XC8OM4EzbZS3o/5vxvloE0vrECg4VT7pPuGUzE885NVRi0m4qoKPhvaHmd4pUG
XqESSSptKMCWDI2e5c4aqdzles6Fqby6O42Wkq9EmudRVRP+2Zt49EB2Q+awGks2
uPUmgvYPVAm+RMGWfbWmUbg3+sofHbh5YA+l1FA1GylUm3cyxHOlr5kFaXCcNsIg
871sSxjsDK59huckWknpTjyQ3SoegncWMU39wFDt1QE4i0BdTRmdvmv46eSIFvr5
uRf471ejjnVrwC40oaY5A2E4wszx7VfYx1zARMP7tJWgTYAgRBuGqGAm447773+v
l4nJXrWCiM+rPDQYNdmuUN90tUKmCfwpMOwIdKiIOQbS0jeKMVwZ/S0ch08Scbmv
BnJZ4zttxqDAx4/WhD3kPAj6Zr6JFEVyTmEaAMOF1ThPqTooX/S9E4cDUyDDErcZ
Ti2Xm+lMh9tjUqpyzwuIA9s/liWJdvvu9oQsDTRVcpyne62u0BHqhh/j5fjZ9Wvb
g0p6JFR2kUtWpPaScxzEGqUnMhFt67BQoIELk6C/U8TSoVa9cBU41Zo3mJOWZdGw
qiaHsKZoDwwZRTRlqh82NfaUGKv8Kj202J1UUQfKplELN3sOmyeAGlWshiNxRnrr
TGppgFOQx2gSPZPIpKhCoJ7xWGrIksV6hUp90F9foBLhA7HR7V2Y6bvBSrn3GZdI
NB4V44IlGj2NN6Kh4bAmNAFU76Y+5lWoXTYxvitfPri25xDOL3DKdSlfOHwTUuvN
QVNWAp2doRK8dgrz/tvHTqLeUPS+NPaoiHo3qh7BW607rfCnGxLB1pq7Dccr6do9
8F6uF29gw/xUCq3Aw0CW4REQHn5ib+4WbNrCKnfsZIWrAyM9zB+LA453Vmz+zS1Y
2CEqbxLx8UyVlQnxU41F2pHX0o7pK1R2DgV1iwVR2/nt5Lu9HfXNcZC4YnNElChL
mkK4wfegfKAN2uiwgsomvp7iOG/tAF/8GxQ3TY9BokzQsl/Op8/IPwAxMzKJIPKo
4NJ9dgwXITwrmfwjxJ7ayFweYw8DenCcTbHC0E8E5snc/tnSsfkzpUylCDkdiB1e
WVMZgoBN/ZuYG1Ju5lO8Z33dz/l5p2kVfw2LpBh5a1rCAAEHd4wNUvVNz7p7BxVd
BZbmYKboMQljbMqB0KW3HJEyenBYdpI/FwzyYpJBI3cMIkrZBSJEY+OypjNXjJ8I
MCic7LLY1/g017M6/p1oXK+Gzr9Zf01xqsegIV9BXf2b/rAP8JwrvLdLCyqZMl6H
vyFTxrdosX8Kuw4+QeMXw7CWRFtdvye3Z0HmxkV9Xqvs6Q1V/ihL9Id/Zt1ThXzD
o2reaTTKD42rik7dlFZ++YUiG44g9lCVIWIdRT0xVj4cGPSWoRqmKPPchZTfchDg
arrxkSV2NsIPpU091qMYI0NGji3JFK4xyvwQjc+xzIDz65ijCuwzjn7jAQd4ewRd
vH+sG/C/nsL/cFxA6swPUTDPaNUNaCgaDANfimNBF8dsBerGPDB5hpGoSyC7BFON
yjhTV3ktsQqNCP8Ba+FDiXFaBBIwHZba8+5pOSyrqovaW5HMawk7v/PdBIbUpxSm
OY+CSYNHaShb95fbyeDwFhlEnZmLBKHFl/71hHvTves44FlGgqA/UTJX6cYzj/RX
kql0Gp5hCZgDbpJPKhQlhm1Ywo0hy10Lk9KNpEs20o/VnO4GyLYS+yhffKH8x96O
VLDXO2FtfMaKFEPEn4OXK5yaPS+BaHxkKerrERcyyMnwph/aaHufWJpep+vaIf+z
lr20Ggr7OlzktYCoeeNYe0JNdt5/9pzWYJC4aGNO8fInM2oIr6hXOWhPSin58ULk
LUCwnAXZeCdK6JstQJ+ZtofhmEFRWvaxCetQZ1f2HQMPxOdL4YhFMglWM9BrsI7y
tddH7p75XiP/aSL+sL3pYQS3+FVQT0KCcS+Bo8oDXvFXV4i8trVbQecOGYURQ+9+
9rfFZMO+neekMxRC7/nqcy0c+PMvO/lQ3ACLoYWVGrMlowvBv+otred39I6BCzgU
ydEtzR8Vgn+GbMU9xT48ughjXFd3TrRHkROw4Xvfho3YeumIMmYEXlgdad9p5wAP
HxLrtmAkeME+xxCX73HyW2I9nZAvQkp9uYgFSh0Z19vJgA4uHgCSMVsjF9cl1nPT
G7NQsuc01R+To56c3wSaCys3YGtfKhoB+SstBFFwlXLc+H4nRi4VdQrFCxg+VAIL
rq7SjRWNEwsIIeIOmzus+YLIgzQMUf6IB1jvSfAzsRYyUg+YvegUgZ2Qv38hEPZp
AUkfumVFly5R5FCUkKl33IyoVlJM2uUmmME/KvxmgYTY2hIKJYxVzlwtwxHAZ/pb
4ocyVBhRX1cY0LD3DOdYlYV90T/rPcJUb/vneDWarx3hAzNWHYmYvfUwn8H+eC+A
ylMbt0ADcAFYZBQPorG1FgQcekn2ZQ0fLAkclnFOchwvTlQgLJIovMvZKrAblg+j
ZHC6QaFNFEFCvwX1dtLJlRE6DKXISafDou/JlPk+n+f5Rh/dzUJV4Pam6e77i0EW
j4u4C579FwHLw86QblPKrfrz1R+hvjANxGZvkcTphHCUdlPjsgj/l31H7lwQJ6Oi
M7g2LuPN4EdzAdV/QipizqBKVhUE5UZvuBuNjlXISqsdlmlpJxOQSe+k9QJWW5Wt
bIS4FbQagPUlM3ozEK/65GoJF+ToZrmCU8ndoLJSaQ2/WgU43sCemNJ8/BSHLKp3
MV0V8+DxXfIbW9FCe652ruwsPpG8QUYWUny3/eQu+JHHf6f9OYqwfQJhMbup3odw
//zQm8c53qRl/AdEtxBxXfVxjVu5RP5bGnNuGsC/q4FISiSu/vyUxUgcQz5zpP9J
U9taDmYMYJCwO7sCEPvqHSEUt344CC/U10gYGbKTiUUcTi43wb7YUJ+7CDVfDUzx
MX0MuVik9eHTgO7GDbSzhu5lN9y6w+BRNLaZ/CI7yoqyyFmKSGcHeE4MSgI1fVHv
NE4u8W7CPKBAfJr9CamYfTXfaNPH3IyvsKMJG28P0HzOG4bMZCIk/CuSgRiSR13n
L6DCpfk2A5akX2w/JpNtOv2oPlsW8TQ6z2iSaXgusMz0HvkhaWiNB3W9UL8bogyR
WiONVQ0vTAajgGMxFZ9sjmnikI7GbOI6nYGSXpAT/ULc2GtpLPeLeNRWpB+mGoOu
nwv+T976+dJOUQ9FRcPGyVRfyk9PGlkxzKP6KhuOUMgpDGXawC1cxVQ4DzBivoUL
O9Ec71fvRlW8+tYiar6LmNIJ9kLKYK3mlIokCSOPtIJe/AYsQ8idiBSFIsAeljOh
acClV+qmy1H0UT/uvl94wg==
`protect END_PROTECTED
