`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yrz0J/soYhyImNi9DwOci3Zm2Wlx62zV6QDVvn0llQATnbA/nuVJjNZhNGuvkptI
LokWXsX7PxHyJXebxA8GlHpQ1RSzZGIvL3/R/qrIwBVK68crxljNZvDu1x8nXY8P
xjj/G+WuMpeeZTmY+BtcZzqyMR+WVbAoYMsl1Y0CGvI5S0pQjikE2VTvExr7ojsV
+MgQMBuoTk+TM+PYDFe2dd6jKfBzJNFECQVfAigl3yKqC1w27gMa1OqOaPRAznId
JMkb4Zz1D9Km7lGex9MVFVskDTtfG3YSauMzBdx6wStlwAGN+gkdxfjUPEtNGSxu
+vttluSubNA4t6ZYRtE6fEhyyV9ju9VbyuA+uz/NbcvcVE9Adm582awBCK878anh
+X2GkJ+vJEQd6hy8Ykfl8eu0ftXE6mdCqhMejl2x7Y92sJc6kHkUvbPkqWS+JSqf
KjGfc8P+KEJN5rR1xI1Nz/jQFfGy7eo7OeIh12CoyfWGm8qsQLqIMU4TBp7Ct/uI
QzjTH5zfNcvz1ygAksMQz6p8Mhxd4GYcbwoVbclsj7Mw0pkJnhuuwCX26sJPLykI
Iwcv9cNzgtvYN3k+/a8ANCJJK53ieYo8IxV2k61JMq5TQGruY+R/x9hF6ZmcW0t1
ugydJZdUPBHkIErBSwxATK9QpFLexhw0kWQwD3ZwG028snSMYk1GfUmx/aydY3v1
dA6464mbxXytl9TGIhchP9ebMJYChnMxdK43jeOJ9SPcTmGZmjMSkfod26Cu881z
tN4bnquNer5qqBjD2RfMYT6SOzZ5Ym2IpLyzSCankUDIZ91Jypmkftbppl4z7wn7
gufJerbxvOSlPOU5KFEYuRT3KewjYV4SgGE7DvRGw/7yyOv2vr56j9bgMB8FH14E
fqChnWevsW4wuE3GmM+UxG6zoDIcNHtY6rIqRyCYBql6GmM2yez9RfVvvLr/Gh4+
/TtVkLwe8v7F3CvEckpVi1+Dfvua7/gw4SshLscKo4IwK3UKcMv3Oqf+yfS1w2Y7
Q1Ae/ZL1mvBF9xo7W1YPLEs07bfljjWBRxW6N4z3NElgRBmYsjDDCevUM5qWDKGE
+DLDccMROUxFevVSLBG/WD2Dj0km6PHSxz3J/zuxkvYXmXkSVuFA9Twx/7ChcWvb
t35wKAjG43w5a/32QNTIGqmuaFi+cWVagaAjLim1f0tdPNMHbvSpeCntxE4tPPIy
0qC+cLhq+VvqA7dUqikfmgfuhW47US1YBt0K30SitISYYu4CnY601aUDHmgtRTpB
nuJVZFu7FPzURQjN4L1MAlYtRZ+sI5yxHMz+/7HVKx6WOzstG1Lz56SDZ2YqS3F2
Yprx6ZKj+YQadTBUC/9nStwXNhiUkacD1F4/5expTyMxJAW2BxjNvUmzAmIvoQyn
jua9HtAbV+DoJml3RbaeqxkveH7buHe1Ud+0GXcosPs86tbN6w4GaSFGRGsTGE1I
ZNLfuqhpAUTcUFZ1Lia3mVzw6mybgY69zaXhRy92wJHH/WjwgDbRzafU3lPTCxnC
VP1I//Frsz67mQKBPgtX2eAIRfxPpep+TXVSBzfQ5sHl24vFfEmGkCGMuAsQ1UUr
AwV34QfiFiBFM69NXEO1VQR3sRS6vXws5dYUPUHYnVJW3eOZ+5aNHa2gw4RoowbP
7bejwjjTUq+OgBmAn7B1LZPX1iWI9LKP9FPuPr2dlLWO1VuZOpXXt6ju9JdBQxSg
VJW2RMzq3sDyl7rvD0jzMPn2vxG34r6TvHq8w2NZuWmCtqgEG+gbzXCf4AXz/fV7
Ivs5MO5MG5HQtpANQK9gwFpc9hOUhoohPlLioyRzIZ9z/GrVZYUxfL4yLmiJW36i
8M8poPi9WxMAerk7h3nyFwkmN6cgkdBNBiIx8Eegrcg5ZEeEq0Wyszbg3604WrS3
+rGzdP8FPKRtnwj4J1PIc87if1svmSOAPNWpVkamxGMp/zoLHouUrII0rD46UA2u
bieh7osLzCI7VqiluAc1hwtWNauxO3DKbvalY+Kqg2ENvwvGgAx7exO7vu+PMCNd
EfDc2yJy5/KyYRqGkXaWHAwlyaXrWak1Zz3eAbr1BlRqCZHJgIHeC1Un44Y5N7gp
G8pI2+/JHTOu8jYGBK3JgeJGVBJQ6SkHU/xOm0PN1D4yrMK5sjHIvDo/e6dlhwyx
XPHrdyAb52iIOqpL9DQnn82ibMhDQVTvZhtQd0IZTCeKkQRoT4E2r+fLTVw5XiFE
v9RKfsnFqM/4jjO9AXKNg5egehLzqLIXxyMcXVgTph1x4fscKC/Ik7kYb3P53h3E
cFXnFjlEP44MLPKM3vqBqDKWfnsQbY/v449cHoSmRk2Wy5smieNIsvzSJPicGk8Z
ZOUat3Afezf79WlSdfLb0WcHILO/DiAf2C95YT/bYVxRSYvEZidEcUIAXJFTIxRF
kG/8ecV58am+ARK78vDEYjszHpPmj1lmz+2t4ZYQB/8iHXYX6byUB60/S9rYNN/R
1E7QJGbFKXgeRi+cJvTicO1IAWn+XcfspiiJ6uVU7gmmu7EK0fz6YUxPEmSOBM1l
90B2ZnjVcHN3clpsrOyiWc5Sarei3kKw7QTeSMnN0rPlEKkkmu8sm8nuwVyJNN6+
nMw8vRu/oQ9+Mb7/W0nJu8bwoj3iA3uDA7mehmcNOAyi7ZpYfoPGJZTUsgWBFrkI
SXUcNQJsYoRRqDVLXdQbyDuSAmUzTvt0GEc+VLWDZs7tKf1qJbFebOQwH7RGxVPy
ZyK695neKd+Zd2tseqzyzLtvY8kTxMKiXi9ALSLnfhKlwPGyh/uNKRwqe7TycKQb
7HQiPE13OIRII4+lHmc1F7CaDL4INv9y7W4UCTftton+8dfGhduWWzONk/ytplKZ
DBm798L4CU8tFc+qsLP2E9s+86HoO/QaRjNXw/VcX2052FTx+jp7hkloLncbdaKC
PhCdHF/GejtHlqpKlyqykjypREuY9yEPNdXDvRE4So+q8LlypIrNbBQWd1mA38h5
ashvhBYVbXPm7+Us6VWdDlD5D9acSOQSPjxBGYo+48w63S1+11aQibNT79LdjtK9
x0/xAvqSj1bv+03qvBcALgPcI2qEYvCe2G+KR4VEqDIRlJKcrEHYmx077UWU+u2t
03qcR0daFUV5StDjRXAYJMMQifPCyTiAKAqpLHNmMrsV4sos/GAk8f7f09Tuepk0
FiGYr+mrktYkNRBowqqlQRstOsYltGoUQHmOtI0sKVeSkPJYd8tXYtLYJpu7VtSV
CfR3OLicC22sHLnw3J+kjNyt6c2nqYC/btFHlHezNQS8S7O0gSDDk8I0qUiyPitH
AAaM1hcBzyPkUVivGAs83EjThLur2QprMstnsHAVV9Aq8d4ccKinUSGtvEyOuh+S
rcAFpma9eJbQXLtMzkGQeNEbCtU3/m8ZDZuZqMK2jA+72iRdes63gM+iaExl2v7R
k5F/NoMmbR0SEIxfjgLbsj+lyE8Sw+RO5Eldr84fzdSCSv6B+euI1XsuZf5V0GRU
JUIn7miEwxIkxM27h+P7yS9boRc0+37DslGutMEi6kVUkfJx7g8GIwpkbCO4zzd0
1GGixeO76PE3r4zdXQqqkNeLwJIiwGPX7wzrirRo4B/3qGxi/xZ3uxyWWpKOFBdN
dh7hYG2zSA+R0edIGqm6XhChZ5rmgBZ8bwGp12hXwmDQP7xiWujZcWR9qQHhcGoX
IrVwza3kuVbk4a1NcYbPLfZw7xvjyI3aPmwwKjgufexlBd5ncZj+yMoTHrt1B1j3
rFN3DstGskUFCYAyhOGzflZLvcdHc4JG18GI/xUFJvcnO+GW1cHPefXI0z9DaLha
FMK+K74I7OEhH81a0q1WL0CSRKRdFCmBBkFVAAiEFNFHk/xXTSAcw47QEPq0sISC
zTKuROhX6hIUm/KH1iUNEa9OyrQWAmW2zwswGrqPMQ7TWyrUMUuhOxIo6gw14oyE
nGYcQbahsE8kpM8LjFEVEU6ks8jRH+9ZaV2K4AUnThAt67iGMiBBKnH3XLn9+Rxx
Az3F7sD4icAzOSMNzcSWgS4hzOHhX3z0NbVNgq4C2HiNulb8VIlcfbBzCSiUy/RO
Omzsh7uWVOwInQmi5bPLssPMWh5TE3AJdP8PvCQzC2NlOPh2u5/ndDrVPXxUSgUu
OOMRpXwRSMPUuDqriqCTxuWsB+hVoXwCNxR3cVoIYr5vG4NFW7+JQDSG7ZQnIctB
QItVxMklJe+gBELZ5igyBzEIxAclxu680uRZlEGWA7s9oizxV4Pg8UkZ/I45U7z3
c+GUBvFPGEMVUlBSqwtGHxvmOwypUUK3/LJeHZWejKlJ6T4Z/OLdH+wn4iblQggd
n6Jjxkc51tr6lCfdxZkdrh0jrsfWwWjW/EViO7pF/OQk+oPJItkoiFHhMA5el1O/
vfU6NZArixpFCR9PI+vuwQ3X0G8lciDmn+C7iugWwN2IInyC4jcwjJBbPlFJlG6P
vq0yqc29nID+qAxiHkuDQG2LPOksPGlBjQmzOprE+n4it34jjGUssNlSQ/PgV5NO
1hIm0fEhbLp8Ywy7nI9tq6/5IaiIuf0SbIxNaHr290Qg5O4i+v8h+FLCANMp2QYV
39k+g7/lahv91UKAOavwQyaoAEZVcv7xw6cJClm3gbcXxPF/TgKVtdQ7rr2T46fg
pe5q91GpJyfz1PycC1nDiTJkDK3j5olSp5KDKgzqMQce+FcOGoDMOdmceLSXW8Jf
Bb4ufLRnVRXkrWm6KjOn8ucK9oniEn/p4k23sP89hQzLZxDzuQ9GPmd/JkDvbyWa
39jhm8jjmf+PXquJCpvkvZ0K+SGmoaM7aE5glMWBGjdV/peRHT5EttUzNGxxDzqR
E+dPjnB/RrWKo/x6wC+1DIAGdD1vcEQFYEM7iIjjxr6RiI1JTmqI0idPMww7w+YF
B3Uax72rR6JbQEp3NnhIXULhegTnxsOp8eeShKNugf1UWoaIxWeAXc/wUJXBDhY5
nvIFn+m9OWLsCQZLN6RjrPUcR11HFVCXkpeSXcGYKYg9RQ6ASjXkjlPH7UUonh9r
6/8TFhALdGuIgJlu+B4sKuo61O/ZcwrM0fDQQSCSxmHIENTV74NlkLqAv7z7r9Xx
LMk8bZWtu5qwygCcKMI55uhXRZFFpyiXZtSrfTTFM3gQ1G/RShWWH1fsV0cSpsi3
8uhqwA/mI3sB6oCmvMf4aCoa6U0A2irF0vGmEmAKK2SoP3u1QS+hglNfQWtUd+Zy
dWAixbMd24hjxX/e0dcNjVTiKiAc6jUBl2Tetz9ZMHQ/6skIADIX3JslpH6+B/+V
4m/PUHMEml8i54IPtaJaqO6Z/Im9w0DhgvUdsATfWx4zZbS8A8kpiMJtNQMcJGcf
YmVRBLvNB3SVYtxhfdmbQndmQj3wSARGYp6aGthUQsGNIYoscS8yJmmcdT8CrKXH
BzytudLB8S7rC8Ct2U2dFy8SeOvX4hO1CagJDtscYnNF868Bg1hXhoEf2nqrNqs3
w+bgRUbDXrEsp9uhUvpWXYibQEDNH7rXg32hwJHXvfP24WMCtnn0O/uDTD1gkMM5
Y0eGvN/+9s6C35+3+QakRf0wGzE5cHsUKNs8+pED+cjYw+ja5nLDZrJ25BMs1UQW
BayxnRtgK+6eyheZObnM+FAH8OX27aueAX2/GgnQQuLz9fM3CDEINOBH/PByvEg+
RTuxME190DUGXvu6la4MCpnu2H4bNpXy1HpukvPfFvvillT2PXadgkkjIOYZs0is
6wX8XBrc6jcsrMmGar5Os48FXeiDju4hBl8heyUjvwS25ar12Ycn31mm7N4LQkzQ
Y+KldaereXafOFaiawJb89Cs6l1KFqW8W7MiNu52AcQRejU+nYzTSLmJL/OYJY5j
MrRNLIimrLNx6te0I/fNpx83pyyfze38hsg7RNRKM7MXFjJM4Cl6j1qDVf/Y1ced
RIbBhcqVRFYodFmajKAQ/JsStSmLhkrgm16bUaDkNd3Ii627ZtlXecp4oIhWh396
gJEGDU0ka5++VQ30QBtiJrAyd4XHm+FX+qEd9VqMU8Trsk+p7Hzd2UIVBCsO/Gvh
CPyRcT48zq6rs/OCv5Y1M6+S703Yi4VEkEt8gSQDfNZk51Q/Nr/UEluGAkBtqOPM
LccJjvIDfiaMe0vX93AMQpeTkAcIYnjf9nlAaJsCaPPxzPmkZZf/xHBRZG+SrLAw
`protect END_PROTECTED
