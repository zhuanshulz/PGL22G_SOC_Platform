`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytg+XGODzWqE0RB2amPUTGHG4De5IIlLZeZeKBnyPMD3W/Pelh5NqfV6TPaKfrmE
DAMP/maVDFizjWLqfs6lSYo9p7KHEHu32YE9gju6BqXrjFKytxAwrmt3quS59Pgx
YtmT55+c4aUeOhDJXbXa+sjN+uhymKrfuj1tCfYmNdjpYXXNpd4acdrpqJgBlyZc
AltjV+5zNGE2tejCxjNH3/l+VbuJpcSjDxQeKhV8ny7doJwyNKeUhUXyfenojmWC
wUqpeont5BZc9tPpotX0rZtpzCgeru93RoJKOEc3lP/3piBiTRfpe8zIiZ4LVs4O
a16LQbUEMZhfLld0OZp02CYY5rlTcv8FdnOnLeb138vshP0/Cs9fhUSqJ5dUDagX
Vweirgwh9rerDxIgk+HQAuk1Dke6hbleTN4Wmny8D/dCahGlQlJFMlljwI3azj3O
bbunV4gHdBcDeJWN0m6at/iT5fXO46wmkHBwG3mIxYQRVxB4DLp6GhugsiH8mVQ+
SorqQqRWmDqjDc+KfnLGVLUyburcKPMYpoTNevlfRmO20qgY5vc9N+aT9CjE72HO
AuOx1wSTecxBbPwgGsGv/KKAKdiVqYybI+482I7Pu4ALd3XDPee88GpJ5iPr1ZSX
jHgl9rklSzts1chasIqljDkYnMlqTI2beMeMt9Hrj9bhlIxP7mYQ2+eWCPe8ADth
3jM6pae8QbSPtuYsvpKtahnigSJ8F4b9r6SJzuvejrOUgiPq6kxFbhPsugKSkxds
s+R6g+PbrJ5pRJJU21ODPW9vUGdkEcZeiGOhCpnjnTuawp7GDnWIp7ECsy9+dVOS
MGrEpzVxhkVqsTYHB0PTxKgpukiI16yn5eBYJR9hozIVkwnAtfjS21EoWeKRgK0w
h7fBb9Sea7SXI1kK1U3/zrvm65k1We+ShsVbsjrKzB6YUA+QjDXvPEt+gs1zawj3
x+zU2fHT4j/6PZTvRq+xkFg+SLr95Cbs2KFOHCfX8ND4N0G/0SUbh4iKJaNIQWEE
sIoL+6T4zJMAN0QM5OLHvswyons73q4LJZXii7jhiEyaG0Q22NcC/Up069IPNwZN
n7hPL5ezWz/HUJBegRlr4/3XQQP0/vwSMDD1jkz/jzwx1cPPMi05dVBPLj5UghCo
wYkA7EW7SD/MWFAmq58HkFrgV5v15opT2X36qvWpYGgfF8KDlqOdGT9/EH5poOIT
IoBL/p6P5ODpMj2tyr8hoEpFpK8nwBpg7VoVNAeaqylSJoIOk+dmZ1WHfSRaJBsO
+f9YyxWqESMv2GnBfvhwaREejguJIsKqpwKamNTdyQzVDL83IoMLOLvNH45uvLG4
9fmglg98roS4bAZiBB6A0PnOGcgAMjmWtm0qubDwawp1nwq8XuUDEFt9b50Gv0Hn
6dqyP/O/yvYWmA2wegmFsR4mn6e3yg8ILkH5ntUvO3kjwXpLq+OwzRkBXOAsggtI
DEWG9eMvV0Yyzi56FKiwEsDl/pfF6aL+uBinaQABVLg+K698Gy39QJ5pCdbOMwkM
hm+AC4yfGgMMwt0da4mdrHO8LKvZkdhLgNfOP1Itbz1kimQxX7+Iy3vTKMvZvaZQ
YpyLOpF2ZgVeRvaKJWjQorSWvMoTo7GnoSP7y6KdDZI87LwdUmEqsrsUFTrUUxM0
SAVrj+iJeL/LXPLk+uK0EbTuccrXr9h/kBnrXdFGc1bydGkeQntQFrL5tB/E5opa
B1sQTiLoi9W8qP/Alhh21txiEBy8NU707Rc1EPCr1toOvWpb3F+7Qn09gQLNHZJv
vRuZ2dhj5wrH7HE1uX8f3rDAXOtSVpBhK+bDdxrhXLzSTXZzcRF/WgtDBzIQKWB+
wLcSg7gwGfg23208dIfItONMEwBPlpqd4Ett7/cONKqWefHW0CEi1E4sOqBjzz0G
Qw8Cc+ErnfMFhuySgpg4N1fotv2l5RpMgnmTR8NG0TGofB0MmQo4+MHhWYO5rrYU
YG7ypNEBJDedcDYenwpDnM79W4udNYefaQoIzbgamJ2DWoJx5KrRS+BXb360W0SW
abO48Adppg/p84ZO6pj5G9bKDqjXGRoyCVdPcx25s4bHUTbS+OqaDSOF1wIttWVz
P2y4/xOLuFcc6fGOprBhaO4/Dpa445up7dKnfZiAtk6MV4sNXazcdJ5piL7cEzx9
VDVh7/2DPKjWmhxNtl4BMQvlxYNKVXrF0St1fpmT2UT7oXzv12CxqK2uVErJfXb4
CT7/LW4FQdKCy1xNr9jIzjfNH4kGWt0CJsb+8mZOBqUJxWH2j3O1Iiml2aEOb7Nz
T6NNmL/LPXP4BHuIvgn1Q/zQIhfStMGFLj4CrsWx9k6fcEoo8ujE3DQQH+DSygPn
rW2yi72++vhRBgzcfqmGLf4DxnCoaXX9oAlpD61Gtn3k60eCnNEWXcz6Utf5boBO
yBYx2p+eNKMeUkj/GZ8TBO2YHxbcWcb5Ege40lvrovsdLROJbN4szDOez4qsDDCw
IdTzkfDpAtVzx7CvzwhG8SQWALCT/qXeQ+P9UkwVUe373adVE/0h8tc+q3KuYbmR
XmcWUVpSjpjhScwWLwk192VRM9+0TkQ6Hi6OoOo3XFWlw5PQMAs7jgGreUBQeCXy
BADrQ5WtNhYjiN74QweGeQTl/Icm03RAjRVPjhzI+9pUDONvFGQwy96rOdtJJKVG
MxIT1wGZqN6IJHeDx0Sqyf4qSBZjsOMlyqITcQc3V5TXOCq0f+PgHgLVXc+Ru6UQ
wI6Y8wo7e7WwduRq6BDNnY9DjAAdI+6QyCSRR2dL1suyms6cvhF4cUyeZvxXDD1B
sKN0eCk9XMiSSu+Wy6F3kCBJSCFjJCE95+ZJkrOciihsAwFntc0T5QODJUf4XK1z
oH+sVSlYDVP8F3SVJ3LJqsTCm0F5NVAoBFmx5+XCI5HBslakX+KLLhChMG6+FclM
9nhBFZcyAGei03qnc4vN50uE3E/uSsjh8qq9M53VljEBLNbbh/9H1161ihuH4rig
YopCuQRURcc+q1tW+Kp4EICIkeg0CyEttXSEWoBOsoI5RsHPq6NrbCwQYLBVHg+P
ie13gQf5CCxObobG/I8qJhuuBgNf1MjRrXql7gwASlc5j6wL4aHeOKy/K+Vqj8Ut
8yPYKKTCvy+o95xK+Z0PZBJtugo7ThBwVuibSdb0sHyd0TZ9w0j+0pMhqeVS89y6
OaeIv0Jjw7wkRUSABwD4X4iL+SuKkJeM3tJq9t8zSnEV7o59s+AYccAqC2Z5WlZr
6JC5MV0BsJPC9XcYmAjx+Oa/MJXpgvSTpPmz6+U9Ee4oPfkPy95sWsVWTikqeTzb
JLQNfZLwIO6slu4THOgRNrn1y/5dl8mikNoANy+9CUInsOtqiiKfE1hOhAzlLpfr
Mf1gJbbZ4mXLLnG7ZKKORofkAmt0FrBUg0X3I8gGESzn4wXvVjRzpEBhA8BW1G7J
zvmQZyTCtDLXCKsvAPvRDcV+pmdqcBsZSTavtRKb2CteuJ3qiFRed/zV1w8PZi32
oz3Qlw4cgR/Fl7nUJtf5tEbpR622pn+AcPT6MjzyYRkv3SjwGcwmcTimLWGnbeqU
AiAm3wKXrldGM7T1y7KWsWT5FgXkn0mWpXf2LC6UDDISZDH4tzIbtYxVmulNkXRS
H9Yt2KbeAWjH90lzQ6Cv9RYdsxr+tD5ji7lF9Xi2Vfsp1ihR7kVnTERCbMna5N2g
sdQB0H3arQeSwxLGr63B/LRdAIsxUg+RjwQtu1D32F2tF+ZumZSrXsCep1pq1W+f
7worlrr03NvKevMMlIpH9puP94zaRtPePuiTaCGAM1CBP/ETobfUCQJ5watzAVe+
2foMm1WSCgXcwXKvrlLHigVeea4oH9sA1922YyOj3ZlZOz351Q27CyEK40VfAG8e
e4PLbzq4B0Ul6FTkeDJX+4H+WNu7qt58QjtUHpqbpXNQdN4bZFMUMKxThIgjFyGA
/NfbdO+fMFCP0QXvHFw7rC1JS/v5gPhSvcOFyOP4z2SLtO23xa7NWa+V2vTX8uzm
38GgmC5tuLSwYlVeMIGooAniBaAPf4ZtrcJepPLZwbneJRxQfXkwR2/3KfN1nUCr
AWoFCdNyL3SDlGTUgIRKacXwu6EDo9c33cttKWS8h6AyNomH+Pp/0ZNQoJMgQNBp
NXGQ07i8LmZPBTO9OHEWoPhHBP2IBT/Fpqms/cIO8I1vicXKH0jipaUOXDmKK6C3
Irax61XtCHqL2QTO/E7FhP2JQA012LVvmILzJ1W4SNIsgxy4UdTh+4lggt5LmwCz
ZVw3Xrkj6VArG/1MjGSmSJzDkjYUFkcP/Li9UlppTke0Z4GvIR4A22SzeupaH0Ws
IHd/O8SRHBprWAl/a920rdhIfbX8J3GZIkm+oWdrwP7ECux18XfpAq3lEucply9X
MC/A7VaXALCyhhlKEV0YhAKoFK8d9lDiv8fqXDfxVcSIHnqjUYUrJdTOJ1yJhTSU
CAEah2sY2h+NWFp2l79urxI0JYZ3z8REL2xWvurjJS4rk3TkR9RVJgWGJm++dZ0n
5XRXCtAv7PyhBCzJ9i4WZcYzKk+rqHTCkuc2LJf2/E162uWkrg2VT6zZILB2zNTj
eHs61foacycuQYtLUbErNMawDICnu0b83jGY9ZmZUkLXVF/U2+Sb142PY4f4b8n4
oRkzJGYmS+EHVOPs15IGO4CbUesq7OgRq1Eh/PrGGeBN3XTAIwGBJkPs9OKwGGoB
HseuQuCxprzSBPgjdaQw/+p51V/D7ybAxJR0XpfQCR3Et6hs9TPM6eM3RAXgNzoN
Zmh6s+bXDX8W+kabEaPgj9H7iTAZnRUK1xKudZODRcpuXc3unJmlPg3GM45KcXTW
IjtzpXJxgXucAKXh+azjym6E8rxWL3tacYL/kppUv1a3G5WD+tbuAPbf1nUr576j
Zd5K+2u5voRUduVE5g8A5co8UFNIPgEM52ud1/YRAM0rNoEHqcG9IojvdgJ6TWpH
4vRElwRa3Kq4MmHA41WOh+z1f+Nh/3iwdVMsDWkpvsQOgb9BdLUmq90xt4SfXFJh
gydM8W1BzednWDw7mH4GtE/J43OhmCFKgIn6UVsKS0afimu8xNDr+2p8QrYjAF0O
xmNyuVVEgWrlUH+x1ls+w0yUWYOzDzXZN4O7Mgj/PGV1ei33PUTSie7JbNR8c6Lf
VBlkmW/OSn8zLh0R44R7fAmW+20mGc+aho+CBaRaY03AfhZknGcPCVD7zIsPj3TU
LgZcTTWeNaDJoKFgrSdjlAiMZ66ip5J9MR5vOOJCCOkYDmsCImUuBM0KjVbTd+LO
We4hwUVbaGbJYRhw+LHE828EOGcVDBJH1UU9r0u+Gl+2K2ZhBfccbEKRg2EMNxEZ
HUvaydpvU9yfzXFmlP/420KchmgmUaatuE0GIlDd3iz7jfnUTeX8NLDCagHbXsL+
aNTEB63CeCtWS37TSDmwB0Ulcq2Tk864tnm/ZIdl9/6PSDQp+Yhh++59aIk8+duQ
5vBcrEqJ0Kljzd9ZgqJg5UN63ZPry7qQ1G4WZ6Ap4ZU6l1B6zTxFfWe8FBiZGoqm
by13j3qtf6l2XCAzN2P3u25qo7hY7tecb9X4h1VDFA4tUOA/6JlAmbAGBmAPLqQX
PGbnA/zam67xeYQk/F+ndYo57yOLwDV3yralLj70EfegYF0zx7tb951cp5dcImTw
4ugF3KUhwFuMTPz0HDUTnrPo3NjAjBdk+uKfSVrm5iDfE5HzX2WcmR3K8ePkmhc5
C2/Yzk1ey/WUyus2R8LYLI2UZjbOhfWn5CU4LuipP73vDuUsMzqU4lc4Ct1U5XgB
ajkKf1/8cY/4XQ0Su8MXz5CfAuVUtkSMeTKoIraFwddUC7h902i/Gw+8ptPR2N9k
vgp+bxmePEb9ZwG17gAlFGkPc25Ufn/2L9F/J5sLL3CKX1ce2yh1005KlPlKmzQS
AWxzqxWgDLKGqewU8D4LKt8JzWGPkxbBszfPQRYcd4JAeNGeqMyttMkngnLae7pE
WebpzgVnvFZvbXCy0tRfYETbGFaifb0v7AOzvYdA43eScprVxlxfYg+p+ws6zV98
BDJr4+uEDtduo2yZ5B5JLhkPXjphLdJQPI1dAxF+kvJmdVtZHLpvmJ8PMhEOPkVR
u9FMzJwma6+iCVsxFUxdJ5tBHe8YNY3TGHw1TlP20/4SKw8/S+ug/N3htvUY9skL
epUt6BjQEXcqgV5d9YjPd5jbXAgvoTiQrn75jQXiAl/702UT/vmMJCPVA2XuZNpZ
JQ0U+x+MhqkWLh0gpeowqzCSHeVrUIyy+4JMxyBajCIi5z59u7R4YiZ4YsHL6Xqk
C2qErmlQH9Z1k80G5xupJWDdYpoafYhCQWiAws8bHxSgQ4Da2mV+y7SMQXVywDlm
IIo9gmynsGMCJA4ej0J7SaJ5GIxtsRR/c5iNHtLFZJSCOjnZ6SBnsAVFKHGbH1RO
cCxOEYNa59sKO+KIalYAohnKeS2nzMaDIen7GatyWRdaeltPSO0OuHnkDSDIWwit
8spgiLg/gIzBdNDxRyoA73pb86Ma66TXcFYG1edDBZAA8i6rQi5O5KjX6e4jbwtQ
V3jVxDQjJaNCuzO7/7MiuVFlHdPcXT98kUjmIPGUCL+Y24iKIO6dYIFSSSyeS76w
r/g1hTE8ySnSGuhi6NT7AqEYD1rNmX6oDAnDGaKb8T5UMEZc64bW8uk+mfllnnDr
8oUk+4CAayKmxWdvFRjrQnnbP79nOV3FbryR3aiadBWKEMP43ofLdCNg0Y4/sqXG
fRPgHK3Su4EucS5pjXxXjcNGd8Qfg4x5GmLamDgNWHMrQzqh8/g8LpjPeGPAKiNX
SWImr9oUwwhIs2Fk5kRLt7SQayVqW0MPzBU0fr4OwoJAQGwSVg6EBJalsUp8sc5o
c9KnWcws8XB7TEeUmFAWTXx7K3JxLTuVMvgqInB2PzOGxXAx9t+2ivtfqlubY+Yy
xS6Rxn2HThwuJwLalV/uoXozhGfDOeNdBKKyJpRX/3fmTC1JQg+CpsyVSGJKKXys
aSx1GtDdum1R0nMKIGy8RoaQoIv3Eu/mnE/WNkvQu54ze3WLSxtWPh7o6SqI91x0
f2iJeqX5OGM4vK4WUKNAt4LuPqZtfA71eMikT93T3NhJNblBd/VySevLEwlHwzvO
NO0XRLWa+M7IHHQ/O5d0+XWpaPCDT8Be3TRcGq71Kv+OhkyeTHkmO2VIbTAJBm3d
40BJoKLz2fpypbiyxSiS/zRguREQATqvS1t8kn/34CsZOcaHgzk0P29bQxcmxuFt
F2kT8TXtebdssfe3GPT1vYMdbzZDQeQEI0UyNePfQQ50NOLu/hj1kq5hk8kumYdL
UhS+DNVCUuHk2loQiUkUTrFVHV4H2xeFecSj3fT4jkxkNjO5UbI9CY0Mp8RN93Xt
AlO4kU8CqLcI6oj05TIXsej6c96/7tui+H9SygUxe4zBBP3frOiy0Qf8DoDTbJ0E
h8uO/lwKTJxew0qN9b7G7zMgRKHIFTbC47nj3GnXpM92+/g1UvEgGUhHGUvY/Ir9
jHnopjRigdNSVVEbsFw/mDQvFeGU8i1m+7LoMztsuai0Sqm5P9p7JogLPt9I+m6r
3U85lqZ0XsCV3N902Tef0+szgJ9L5nXWuLRU9d9o8PR7x3XraFLI2xwNjJwqk9Ga
cXdRq1zhXuFHzscuIf9viAhehHFpxBVLhzIM+CCWzSrWn4FOGszia0IKVxydby0X
Kp90YJ+MvyMwcS5TtEHh2hriqIa4OH3V/JcaRbJcAFaskrq4eLgDgXFpGNtLfzap
Jm85uHZlRH0Na+UUa2K5CD+AqSSpxgvjyfPsxdR/kAWvmBQJa2FrZsh14AWRQqAL
hWP18SKom5vj3TB6WGk+83xP4NaznOleI5uGYoK9eAlBjKFXEQPEt0l3CfEBMymu
S4vTNtxmPsnbWcqI4djwW8lZhJm7TLcL3v5dI92qdSoOh7AkIm76PDy/mFuKseLU
JHGjKQYVOkbLm8/K1yCFwvurKcAKtZ8kzg2i0SJp26idhJxTSC9kGrBSmGEMfJe3
qYsS0xDYGFs6ucHwW0WLTn8qm2aL9hj38lx/TKZSlYKBbXC8BPKQwsVpA1Kfj/nm
Vrl32l/rSfJtYI70HTQRZRt+dMq23oOfWFKhPHs0akiDUKk9uaXymnq/lFNMCp6i
qW5Nv0RBcr4mg5sZNfSdhD6VB0miCzxrLLPuR4E19vFSElUwNEY32pZpxtiAmDjJ
qYnRRa4ACaGZxenf6Yg+fbVPWGEE0txdGEkzTEpRRHwTbh+PMXoCS/zFDzB6bUpy
JwlRjzg8p8+4p0p8Ku2g74C3n8exBd/DPCcXWSDAQDSy8yXzyn/eWkcF+o6z48jG
GFnjDyRWlhoEXq/MXinzDQXKpPvseDMyTJb4798oTGE8MAO34MYFoDzXk07+HuoW
sGTM8RBCiSlYIwUCZaTToU6iHOaDCJycSHYsPa5Mp3a+N2z4weuSqLZbTcYNJh/F
3JuLbAzeB7SruCpMlBPnr8+LdDwT6Lkd7YJl55kAP5jl9ZW3YnK83A63KHckMT1E
yDbdNhVWkPDwgH7lnmNN/3z5bypr9WVs/Nvz7ZJow/4tPi0BzYUYYGDllU6zCGe4
W1YWKiIYUc76ocB3RxZaCjhfERGFGygn5Zq4cLyujWYkWDX6lbD7bJfyl7m9If3e
49biBQFIKJDneWTHVJphVxBr076/WTztMIoiaHfrFpELe5segxfIfwUqwmpCQnrY
baiyObEmWgr4GQWWnd/VhVozslTxbYnAgrXIfJ8AJlxVl/RJwOMfzX1IcMoUSkLQ
YlpsAYulD8qtuP7RYERFskcys8K8Ul8CwgKG7KVl5O08XL2rOj+t97U/UV31X/jr
OsNYVKN48/oH6RWdHf5FPvyJ2nO//KRzg4Tac/Vr7h74uHzJz9+y/dxarwdgPvj5
8gQSKQGX99XQ90Dlp5HG7RjdYFn9+IAe/QQXGXeu5rSPh9/MinGgCV6GVcJhc/dn
WWA9LXpCS8m5Q5QhSP8pJMNgUMGV/TM7NIC+tor2AAL9duJnKmxUSjtBaBNl6GlJ
mIsfUfKXgPIGlVCdm1IeKkH9WUFrVJxhodLnt2UjDrGSaZc2z3eqLx0ORaWp2Hpn
58eh4YTUha61td0k21+csEb4O9sGDLtUU59vI+wqhwBWqlUJFUCV8ZYZfujBtF+I
tmZqGfKmv9eBqDz/7ARVUndlEF9qu872sTXQzzg7Ol0iHlY5LlJ+mOOEFn3AjW/g
nz5xx34c3S8sT1/TPcYfSiBK+05rbn1XY2E101iHdIJX25jGye8yMB1/ve6zKzcj
Y6oh2bK4l0gMny+xzMbIP5lqbpn+QIpSMHtSyh4ZJDbmEh4vlZV7fZGT0QFCh9BI
USpQHbdPfdwpgD9cgaZNNSYrbjV+kBsK/hVYu6vrN3JZ/QSE0xkYIoBWxjiyo4uJ
eLSWyFITV2Kn8/3YhCte7XxR4UI3jzxHsI7WVwmMeR5JahD/TGfBbATlrfFNQZvc
rfwhRAaSriqAUueSDDr/LHNcNLrzbioi0ZNYr53x9k7MPtwBvK/3poapgSzG+sxy
OtEKCSKYjoew1eCdXtYvCbqsz17bgztar0koMC5AimCeSIhiepT0dysG/0TGFoGd
HzmWOrx4sJnvDbkR82Ovjj8VRTUVskkOsd0u6TefiF2PsMOSFSmvIswXDWapvrLP
VLHHFgt4ANFWnIUJOuUCKqehgI4MtHN0OOOxqzd76bP4c5bDpCr6WBVICe2h6Psc
bxSoRQriE4va3dL4zwidtFsUnsjN0NBnXGhQubWh4nugI4CtyBV5WYglM5bBLznq
LxUH2TWOdmmnjdbzPpVLwhm/6/OCis+MNUxr98n17uy4TzPVsHD4M98Wfca5EnOU
8wWY3O0+d5mUtVstxpVHp2QMkOM5IRwu+jF+ANWQbS9+d+q2VC0DBOY6+Db5As9q
AkCswSoy7ZaxJ+HA5x8sOsRNuNM2FmjYSysnZdsv0uaoMLx20szetfGbskD3YPVv
/NnhjWafEyLOaLNla5xG02tZvghpKEbnmxPlHREQS+DPS9vK5bXPu2SzQ7PZpOGT
U6TOmp3kHOWYanGCWqIS0SMZBB9UcVHfOaoJvWwGQmaLZpQCEe6dViF1XZPTAxqV
9IrnOp6JzX6pgciZwy/eo5g9mgk2Pv5bLinYSt1eGk8LfImEsqWqtdEdWAqdL5AP
3r52RX9dvp7NmHujXbRO3zObnLbxcPlvE3kUHWuMyaHREhGape/8EsfbCn230rsn
lYEHZGpEw795lKBoBz0nRE1D0H616wy6P8c1ScQexAz0s8SKlzJ5d6PXqJ9tWDSG
M3/AhusUDcW1zKqEAdzSggKt9oYyKi78Ib+mxNDjD9IEyU73X4pP0bP+mWN25Yqb
WGAGO4jbN21dsQOMLMHgP9kBqp1DmC5CdLZSAXqz4UMVmbAmKriAU6HAoa+9XE6a
etIhNYp7Bwz7PqlWTpa3USqL62xj0InZpgYzz6/lolVzf/RPMRGn5xsGetTpD+Qj
IydZhmBSymeRw74ZUJUd8R86bNKiplmUlhFhZuLtr/Jbodd2/vlyHhxllLlttJ61
ZQ8p3+n93lgDewWZ/ncIdMhGs1vF6ywyslmiwqJYN1Ahf930v5mlZQhrVAWVJGoK
`protect END_PROTECTED
