`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dw+VD0vB876arKfb5wJIF7GAONoX724QoA+LuESpebaYmicQHsxY0ZJR9Xrjj/YC
/0ZGTsQrXD80vpPbOXNTYVueedYp0r9EIgJJykOcvdsmuj40Q6mMXcHW8ROx8Eg/
4R2I5GFsTotzfT+DhVjrB9xKWzH+WgFQ6l9sqazslHPWzbjvUQdjOebiuDNZGtqx
7wtNUYdf/IiKhr+SgnYkz5HDw6Vc30HES7e9Y5ITA5u+lztXGcuPCH+XC6PQn4cf
DG9qadZr457F6F39Sun4OA==
`protect END_PROTECTED
