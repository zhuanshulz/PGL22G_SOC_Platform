`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yE+9FroicaWp0+WS3UVD66yPCTixscPaPFEYz7wYqckd0esPpGNR2+ve9zBEd9Sb
RrIyswW58yd4uMvL2YrdI+JyupXZgCbrbxt3klQ1AJD230I9y9linWumV2o3l+wa
dccRJDjEutYHiOk7dTkei71sXmcidb/XlvOfb7D4K2mpBBz4V3WQTZ9kwmEYb8ZI
AMSCqDP+o/BymdiG0T57ocDINE9yAc/qBeBmmyRqGVquLHEtDg8iaMT0MbTNFd4C
GYL9cn8y8ZFViEwC/boDI2kIEQ7qKdE5H/FZ9nniiApioJN+vJrNrziIuN95b8/I
PzmjGi0/GlPsqdrVKSu/vy/nVLLw5BJ3sYiNACsoLATGackUAHmuRIdhzwzHlWbk
iSsMFB917CaC1VFJEg2ytH5L0KgOxXu/cZxNuqgzs8mQkUMG1LS6RU/jn4YHP0DJ
/oWH7F8JVS7oaZusJEj5owU7BqfyyCOcPbrM035so98HhZwiG5oRto8y8EteGOBB
IEcKM+clNp0OkJIhp7uurrTXJk6S8eZ5h6Hjblw3pmpwsAIx+W5jiZ2ryKeKg7TC
57OeE3t+oIpgUyVaGVhgBQ==
`protect END_PROTECTED
