`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+mR5bctpUWjwNEnHChuICkNiG4nwRzC6Cq/XEMj6Q/IVgNrTSk786iZ6hmjzn5yQ
2FXhpgf41klYZjZ0lAI6d559FKyalbuuAHF15FhjINM3G84l0+TgQuV2nfvFPlND
G2IcDYWdD0VIAkoL8WzsKUMZesSHVgkzndLM/l5AUnfRf5dFLBBsk5qqsiaZvr7S
BBiXDqvy7Q37XYjmYfLA4FsmsQKuktaflwT/bPpNBHCtlUL3uXqMl2K3C/o+Qcs7
HAiGzYg04WH+WPIdPcq0IWnzlSwbxenAmKJMUCxEs6VmrARWbARJYz64541/V9Ka
pC15PHPeAdJIyX0Dfmg/8cpeMWyE37hs8GWIUir7zUPJFLiz82qCa27fnIshcx66
dcFG3dG8vTubeXIpssuBBBW1ypcOyJBARVNJFRb2fPRfUap0OkOODbFF7lDNEPBN
wX1IQF5ue7aKi5ZAI9t2RwDNw5TdvYd1dgxunDe6UrVXztGZg3SBrgaroYkWO6ds
h/O0tdTUtUNtmERT7srd0BOPbhfeT0g1FRuU3ivLKtiAeElav7QMnVY1dqfQUB0Z
lWiXqxGI1AI6en+LlkI0TEmrnBlld3rvB5KGPR6DHZ9YGy5uSZkhXM+JdBqE+oze
n4WqPg7y48exVESW17x70Rh7JwxWV5kAgsSXmBzZtON6IIUQ3kXfP9D+svNoGzkw
6/oiYoUfgFsoC0dZsQ1aVqyTSDT33Wv2cHpVOF++60VKwjFGF/aNXYjYYRund8jc
pAa1Xw9nZV/T4OvV5biypgqIjmL6iqKAkHVl/GRXNwyClN68qDp9PisqszxzEV5o
YWpIJVeoGK02JpSlU4R8aQWfMYY29GVdW3XOEPGxeJQOPQFlOkik97cVF1bkSmBv
MsvE3kXp8eVOc5iqsSO0PYwkrR4AFk1lTbRR5oPet5NAV189s5VbceaS4fnLJ9PI
RwapCa4Q48EJvdAPAmHT9PWlZcpBGG0PBs/IVzydZFObLwx5L3B2ZOMjRshLL1nT
5HB5AlWIjDvoTeexMEIefsqW4qqO60QaGSsdjOKfw1QN44/zklKHcJDZz1DeuKcv
MMyDuEsx0/dHJyF0PzGVeKXCkWGCLyUNueAmSsDiYoeskfAtqmm1/hFhSGMgwWDj
MqlGVN6/S0jMPFN/7SfwtMw4GQ329XXQn6FB1g6xeDOD+khNck413jb9g94bKaiq
kquh7agVje5khoZuDotpeBqESpToLgA19twZ8V8Bvkel9zZiLBRj9d4SxmERuG0g
yC0aEbrATw22+V5D/IpfoqEEHsdc1Wa+ja6/2I5PCBD2XAersERllQ+suAogaxI4
fMEY4Bsnxgb5hRbVfBsM02ZBSo4vfzz0gVdSV5wlx2mM68sTIxog0ni3zjD70QmA
PLtkDSmCICtprDvDkiYR5JrJ+BttCnyzxbNv3+E4oK3CvMgSfP1+VJUuR+4kg1/T
8UZL61uvJyYblj5053UlooNTRtM7C2ZSQDXbKjVNSLNhTFP8OMz+ay2g+HCK2BYq
QAglVxDTTBbRfnWsM0UVF5MtkOC0CLAYWPkiSVx/g+EXsbYO73zT/J9Suxg0joIT
eVH10UMd+g1vIYwD2CmZwKQCnsWU5+bGz/czRet90OET4KX6U8ITdYa+DvOnrFES
1I14U7y/JuPtQkwJIQxUW7+B7LVih/tYk+90CNnT8Qad5tpvVlBuj7Gf2dBt5Osy
Xwn7gZ5iv+9q0NnONuzuwJ5ICJNoLjYIO977wUtz+rOPxfNoBYCDuNxUdPrnxFv0
`protect END_PROTECTED
