`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqweNz+hDNvyLglJ8EZsFLDpclWQ6Ujy+YQvcIeSGhPOMS5XzcyaBRh3IV7RFNmx
TrtGc/NoyHiIueb4ZmNDd4qsbaMTXSzuuaXbugpDV9DEx0BEHl9nP9sWJRj8urR9
1zAw6C8wNjx1YBRemLbc7UmBfg2Y2/O7m+0LCvIShk6bJ4DGC+a32XzZhpYvnCrU
52lmowG+dHezYhu5kaJtlbjw1n/Ov1J6PCgQHC8Uk53hiiypkhTtAB2kgpKWk3UH
DWMX4dR1fje8jClEZJYs49sTgkIF3aapytTvwGExtIX55cCA1KXXnVhyHwbPgYQA
+btMtropAJgE9bEU9VCoIBA83lj3IPH9otRpX8/ls3rUzU0dsJVd0p2jzkI6tbBu
31j1Ip9xqddcTL5yNw9ukvuRdyNYSFrRvZQYvUGzUbRfAxmMnl9QQ1bYifvlUWL9
51TfkFZbc9LQzCQHW2gC/0IrEkYpyMMvejnXLFplf7+hH/uHSPCyC2b9I4BKaaXj
eJFIOlxgOzyv2IcC8qn52+Bzt94iHiCUgQiy4MFSCPH+xVFcSqs+Y9Cix5PFJpbd
UGLnsRG1WW51v8nxRiN3UUpM56D50sJrjUp74Aclgola+eUYOXaIpD+U7glyRVDc
GkjrCFkLunv0leyceYAYBlhfg+PWRHWSwvgTZanPZT+PDWxCWSf0lBw+jU6bnGCT
8v+0eOu33PmbyMAZlkvIzzQ/O+o9xrZL1dFOiIfFSAaKOyKAqnEbNOxi8C638uJK
OkEZ7y7zL3TCiHAWaN3cffvV516C6ymfHAyKjmX2XHam5RXb8Xmgc31cuUMEq0mL
N0MHP36WGde/Hra+HLNc+/9Fmz+vUvg9Cji4XHxQ9j/6OQ+SqeHkCvneHZ2avzsM
I8Rqybua7eIWQz5CLiu3n4sOKrPJjt2WYBMJGO8MBdMgUySkVTtxB5rA9DDqRFKS
BW68s/U27uDunR1D414Ej5afZ5j21DAxXTZt19+XO93utP3SEkHiXvaTqFz+T9G0
uki5RH74nMzG+Ty/g+0n8JoP1KfSL7TR/3s0WDwwb92T8im7RJ03o+OcSEc9cAI5
pEiQIRMRy/BIfoYD5bKBlIa/lDcCLZKXTaVEZP5i7k/7q9MDoB2XkJAGmglHd2HE
wt305iR7gh1gm7NOvV2drs4XgtFGBPBW+MsQYgpaGFRf0KMqljhPEEnGg0zBvIB3
BGrbRhcTcrFMsz1/S+T3fWNFtltV8+vGSUiTo/R3HjRIBYWjlfQG6WPxcLEBJzz7
VG0SdLiD5emEWi9DMmgitWfmha4Ifo3VscZfPerwLpYgGmUXY/AhkLV1Ph67Kp55
0d4K8rkUY3SKFyTLvgh60GmA5Nbr0VDCulfK7Fk7PtqRv0sPS7r0lanue0Xxyp1K
FL3wo+P4KJUR9cVDtQiZ0Hu1oSqUt+PbhF80+5PFWp89uK+RHwxhWRG47kJ4QFg0
mJs1b/21U1BiqV5W7dVQNslEFIvZ2iKFxsFPWrbXGGbMAiq4gRLQJ0ordSgjYorb
rhs0KAogf1AoT2EZX0xEEvWL41foWuKBQCzHbKaqfysT0OJYXHZUSr37egssEGHM
`protect END_PROTECTED
