`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AINkpbNxkyNJsP9o2i6n+sb7rgCbzQxdbU7K9g+I8h7ZW+HRteRgYexRuYI11rkR
3DY2BosZUnQ1J5uvRocJgPr/+y3WZDUjbjeHnq+EWR96PW2WkQk3pgt65kB0+gOZ
VOgcBIkcRpUBtCOahiyBZkA2aJES3ukyE626n35qOfUxZB/pDf/CiC1xWndQCflN
f38nge3GBxuWH3lof34WFUewqg4sNNq1+B8eZhd2oMpOfEXsYFwm4gcKCag0+n4O
U4d0hfZOCh+hkCQXwWmrjqld+Cwc8gwvaQHKY4fnoutYf+jZj6r1ycj5IHeHaCG5
a+SetjtdxgQx5Wi+RoiePMDCBOyaXNhtXGKLmVqnz2EDbxIhz716TG1EInYN8bWd
56FbF3ors4apj9NIr8rAeQ9S1KHbryB07A9F5foANk//ST0vKYURDfh0VBvCRyUm
7KPNuYv0jxUHcC4v3dFHboNXOf6dm9UiBniA5qFLebLzKK6dCyEUS8ejejiv9mML
N5uHnrDiDAOBBs8A/Mp+V1/X8MS5LmJjerqOVXMRcrs=
`protect END_PROTECTED
