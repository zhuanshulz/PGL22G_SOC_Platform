`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ObJSwtU7eoDj5JyJPzAx5nBamOgJcIEnfk+X6OO1ket90x6A56ZckLJspKwxwBoa
tc2X7VtGPSfIT9lZMzzZu6j/p1KaFCmCBfYgUcYc1aCxdlhWwtL3oW4myVBS+bi+
awiPlRXpx6Pe6zUW3NQRV2L4s4CGkxOaaWQaiKs7aVyz17hRdvuCTRP0+LvLExbA
uqM2JCj9HOoTra6zPKKAziv5FRk4szk7jr1deBOSLS3oRXlsvDj/uVO6nVjq6fFk
sFuD3wbWXDFCMnrrHXlR1nKCl33FvwwtEU89OkntBhTgt7wVIT0jmY/5Z07+NsM6
2SA/lK9dVaVHstGQXQGPfPnsOxQvLSKkv40tt/XzdsWwyqZXOIINcFls5MmJdP5i
VVOTaHCgMiW3YjY4N79GyYrMd7nIpUahV8vYCo2+M1cm+92OKDD5aSShwF6fYF+e
sRSGgTdmCuBvzDjlrhq8HUW6L5o0TovFqkF1F9a52wEd6LkBjuo/chcrvgEHafKM
Y22ubpjgnkuT9zA0vWl2sHxXbq6y9tCfU0VkSgm1coxGpVlZeg/1l+WtZOVja5Iv
91mIS9zx+nojQMqoTbbtZpfHDIfQYECBi+aSiV5lwwlzFnlbNx/IZprBhUqeq+Of
sSp0mTfpAfUZEDxe8S6VMenOcqPcSvQ3B04xh+/PkOrdWW1we9WekYe6Rh56kCyC
o6x5Lr+2U4Pv0Aa8QTsvT05+9LzOxEIccbvoiswqs4bwjp+efJJSLzxp9/fEIPSj
HjKSXSjl5ljYryt0NyfQSp+pX46k36QP9DTA31JMmlEliLHyiVURsavVm+stVPkr
JJJWY/e+E1d2eZqmtga/emWTSWVIpMrHn75W36B8Lt1cTisGaEfnbGUXhzMhivU3
fgDsOmGZT6wElmE0hQdWDl7xC/RNR3XNsfP93kzKilvQ0QevmCaZirh9gYcmUlag
bcJ5mz3BZ8mIGzVTqL1YjGaytMg31buixF7UmWw2e0nhgYwxNbPJoJ4AUx7JTs2+
5VP8XHZEe++Wv4kULyfjD4HJlz/dwjdUwRyy3bsJ5a4LDA4Af/1wCItQlvhDLeC0
Pe0lPZeKmiaGRpOie5wvvb8C09ASDKLAap8E1UONinMbbUoO2iT9CdN6P65WFa+N
pRDa7qeOLgASp3cNwLTrU8FonClLtTGx/kBoK0cWJLlwJpU0r39gZajWzI3rITLv
YO0sWNhZ4ITQcu+nimQR1medJ3hlwvVGzahY3j0xOoicJXs7e3nDwDb5Pzc8re53
f6VKO/2of2PFmI341RqQ25nOQceD6cVKhtiyuu2Nkt8/acm+yNlnbAS+KddKQKWe
EXU7Xz8etiJuaq3+qMyP8CUc05ojGUWaGIXYaDTMetcu/wZsvYK9YkRn04t9RgGM
Ruw3Xm8BFvDsd5vSuAapSjA+d+Xdq6uqt3cl3UT0hQhwsyEHYBHpVgzyamubS7Pp
dRAT/W7JSVKIOhFIUabDG0u/OhfTuAGL9Ptbfq7dzzOtKz3FMKLV9qIX+MW9cL3o
FRoq45+DRSH8UMikNOGeWTUkeiiqEnRp0dK2NQkCiyZWylCZV14CbR/dpPi8Uu3H
s1vEXuopdIgEHEXWQ8fM17Djxu3k5OUL3XXXDHpB0yx3MZmOcidJLi42CTOh2TUp
DTCvLv+e70wq0eupdM1TL1NjH488QWp5ZwojRz0t+twmd191XaYgaY99IsJEOH7G
IPNoDAsuHVoNY3k5JDH49iAF05LnES84QNRtCb/btAjmI3ydkVJGrg55/xSxshRB
Rpb4/12o3P2lnd8oAEqy9K64GCJrrF+Rd5W2+m9llRfi6A6y/pyaeJFdhw0BNtOB
+K7JXiRL8TMrCH1gPcxWXzMYZP3JnuLgCIlaYNOtFOGrrZnKLew5tA13KsOpcser
zk9d7L08JBZFUlrFXBiIo3FAgVtVfUUKOOdLB7H0snJyiH/AW4B692h635Pzhk0I
mDj96sFXpxYMggN7lQXsr7XFzEIrrJNoH0G5a1keTVilOKPl+jlC98biGPTV1bDL
s3/RNt6pnhQgdzRqw349TqFNI8hjO6G+HsN9dJgwiYeUTwkddpR9QIlENfaNPaMs
76nJ+h82FeBM6mkb0SCtD21wKLaVCPIEavbpCl0/+HWMvzLeX3zgNUpmCnYBcTEE
WzWweLatJ64sDmP3bpU0b/vsI0XkzVFMYW2DphdhW+atqIU2642kXrglJXKRu/qD
4vsEdGwKfQtNi/cOOGsonb4e92ucwltuQdfG/3BoDHx5tU+Y51tcNjT/kHqHJV26
iQubTpg4Lk8xj+o7q/cSk54Bbepdztwp0KUXp2SBY9M1LJ+n8yMB1BAkM72NYNvU
zxNpi5+wm/+v/+Xfw1xndS/e0KGG+Uj390PIcbZIFmAyu1Bg0lnTTu7DvWqPdyVz
pa1kW5OtHcRK9dff6dPVEjWkUQrvfNv4SjQFMvbc6ZjzlzU/tJDpIO2W6XQCikOy
wQDYHH4haR9Vag1xcSK1nzPadOgT4rIprjOuDfdcTAUwiqhWjf4HZtiCGam5KnU+
zVsT4atZ+4VbvGoXATtw58QFE9TvmtwfZjlOCvMmqe9F3TntIjr0RWnU5WBCG+j8
1loziXvUxbb0Ve3DS9HuIWbkIjXn8+H2S5NrRBQOm6b92wa6LkdIGkguq0yrC/kG
rr59bBR2/mnp086l4lJaUB4iv72EjkuscrloC0h546opox4SksIM3DzJpqsLqoth
YthXLcSlDwAZOrbhtnEABHBpbIc0ouZVJM+bHk4OfU90NEOAy23+50RcAZeXOm28
RiIHMJ+H9wHVVZIcua3ZYfhKu7tjl2a77fYMFfzAkwSXRXdjbepGBGNh1ZpisYZq
ikws6VqMSaeJ1I8f8+xmJnXvVY/LIUcks44U1bogk0ZnukSKwKqiYNrJdtvVy5/m
o0srx5fgU+16FFEzuufBZnIxZeIGa+LjCGaYoUg7bfroJnx9r2mD49SucLUuqKVx
+qXFscXiY2DPrfyMpTqQS4ZMWkzoLvhjFQnoE8h8R9yDSUByBskDDsRQBuAcbHxe
Kks/GEcCJuNGKyzMjBKUVTNUiOsfSN62pNr5XY4yH/7uRzDvPlNdhB+yNeLu61fp
5qRQN+fbhGqJ59616CKYbieT31g86cdmmU0LM/sbhOA8zgHIoXOwRDfYHm3d74ln
j2hl0dIWG9ysvAq5jrgyLmRWBwtQuCqk6bxQW872FxGrgAEZDq2MEwvPvHF+vAny
/RxsOPXA2NigRa359cRRUD2EUW53Q9XJfG5yhdIYanqUyeR9YLoEXQ5rE1kM9vx9
GuXRcPFrHdkRQopICCuL/sd2gfFmIF0MJ2dzFTsrD+sfeA1OhgsTYnOce9Px6Koa
5rfwgycXbhENE3lUI2awJS86UN4gYr0vn+SVOxt+TnH0hgvK5KDx6PL/xZBlHs8k
xYMBZOfxXVwJleSM8qv0JQh+jx96za90Rs4iEoW9ScsE+0pclNT7OeyKxYYPy6bv
z02oWXLVFEX+2FJUPh2eEOB97KxGQGMluZZOyyNJnV4giQTFzBsjMaEGDXWt1pIb
SNQXVIuIh8VU0EkVbsr/rGv+9d35K4I9PbfsYTufifbMB6z1yhopzPskd2GM0seK
Jgho7g9A5nQUKeiOe7YcipTEW/Pcum5Duw+dLeDmzhWrp7Gb/uN7laTOzJeSCMnE
pBVddcmhYZaRvsvO4+mYiH9UeY1xAZo1gWKY7fD5Sit9c2jnggllFqYmz/TgYtM7
58HkQQZyadu9bSKdNN1DVTV0OjrKKhuJVKSGkVA/heI=
`protect END_PROTECTED
