`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iW9cI897zGtxUMWLkhworDndoF141EtVx+F09vgOugyO7yFJ7JfdRnZFjaEq8ZHK
oD8kVDnxzQI9y8+YotrVGClE1LhLAI1IXyLgUSTHbK3c3W9xFlPCcTp64eL0yVjp
ZVF//D+kA5+8ieeiQAWdtmGh1xae1AsVMgQlOtZFbGxOIk12d4/YI5FJRoURq1Ou
K66Vsnj1BHqV04/DMwze9/7WkGcLWOkiMT33gxgAWwXy6FTm8iRW0LywU4fQ0ScE
OxyncbzIZcrchKo0wIJzw+thTnlNr9VCTfaqttiezM8AXKhqLI3yXxV1EkxIIdaD
LGV/z91GC+Zldxx6O17avkq3rwuIJ4HEYqTavAAOyOUp2lH9iJrAynzANMdIgWMP
FDaQ5p1jXdkI69Pw58WykQ41DrZPqD967YruA0f7HVDmGG7MHPxAFV+7RU8GG3/9
2bbMQBD8MmCR8Nl8e8z4AhfzkMUBc0epqYdGMrdb99qLIg17Zw89jsuUSdlREQ4s
hl8NFnkfhjGh2mpUt9t3ttV0+6zG2ln8wJVuNBwF1OqYelMcfFBaGwZTkTyG1C7o
3sScvvoclfrhKAOe99Ab/7eN6dbct3thrWBwK0qvOyV3dQmztSuM1PSeTDD4JCDk
8dNxUfCv0UAdURUQFGcfnGGR0icOpsMWFka9MyKyOYlXDoWorPSAXAzwLK+sKj0x
VMqQ5iHUuphazA7ZlteLhzN/Gf9LPCedAGbS3cg0kd+XowAkX4Gog1r+JM05qbcb
XkmPzL4ZAtgsjJJPuI0AiFwnrGKquykgcV+JwUBQEQ/5RTy/AmUejneZn50/4NBc
uIPn5+l9lA771a+vGhkWL0urTI5s1z6zjduUAauCE8UBA5cV1d925IhttWk+O45p
/wBZ+2YiXqVRI2oGoR2IpWD2/NgBpXG194cFkcIodjob/Xz5xjvh0lOdbzKgZnRi
5ROakV+MOynl8DVgwGzXb9mpdamXjHw6rn7eq19qeT1ICcx4qHq5etCNowvaRL6R
yiQqsnpTyUtjm5DTe47F6O/joX24KbLVLDBR8cXFC7n+WsifPXdNNN010phLe0Ga
Z+yCzAQ0SCC4vJUYwi4G6rKkjWtgFQfECzpFjVbqgHI2MJ4HND8aYa66QHmKm1xv
S9395SJHjX0u8EI+CilFmCnqZmjH/507WWMGeR8ZuywYCI4Xee3JMVrVQgTy3lFd
78QeLz7SzLXTu4LbMr3u2A/dfY5/LJMfq5in/RXfstZuUdDwCT/ZBZHGIQkQ4xJF
0fqI4UqTJByQcUa+MKqv7lBOrxgW52aCUPoB1hRis/VVKzT5DR2CMTj/u7mkFv/m
i9uqryGZnxBbnnqRzy1dubT+swQxh1hX8SFpli6GZAKj1b9vVIA6YnT7V3eT/t13
uQXnY89Lkg73biak+5orNw/+IZhtf+6DrAGewxQWKkuLfk4/FwtYKG4FBD1rOrWC
9CJtUa0oomOT5uEoXBJQkBIcZSpcTcfbBQrztnSR8+Hz1AQW3fthY8xbT9yJRY5O
oiCXPeubbSOS5L3X7rB7lHSioGmkFWBc/GNUgtrjXk6+8djLvFi/2sOSBw/RM8EJ
otVv25ddKA4vNW6q3miKJwYsAYq7CsugPEu1S0ZChYCQDhkNwHL0+0slys9AqpPO
UWZ3Ft8clRiKVdg7+QB0BbyjxiBxYHaZ7+BTivAGwW8ZT1EMsqRssko/WYYQmvfs
/Yn8J7Cfmr0tmCU8HYgGi3o33YrZPOaRAdhAlNwRzljzFfJ9g4cJMzksnGKKVi8D
48myi9tgtm4Yrvsxhd6Qo+b5Rx8j9OVoF0Vtk1uUEzdyO/2DrzfYsjeXhY+CCUZc
ozgUgZbs7W3ka6sxhmnP76E5yTcE0YPeMsPlWJet9vfWn4PairRwiiq4D1B/QkQp
YF6JJw75Gk0wgrE50AOmQGpn9kjar8AOiYG1WKXca9QyslrTRfVNUvPhMqCqatAE
Hw4J4qMu3ETRf8hXcsiZV/blJ0EuMZ1KNuujztex9jvg5+ww19WGnIg+pv3vEIex
HpeWBC4tfqoBJY84v1Q8S5z78CuCRcWORd4smxqBjNWEeSDSvE25kug5LeEbF+ur
m2fkSkx+4wuHuA1554uCzevZ3gzbLyJzySaN+YxRgmbbPAG34wOYdcNElf7b0yVi
VqtJlWAavirS1I27F15ZUF1eE642RLWVxa5WfUx4HFzK7c98xqHW7SBlRpzcC2Zu
Qlbl7olMXgs+VdTPhS+Spjvd9JNjHzrboQ86sTrHZDbXSRHW+42t5Ze7X8UcT3R+
reahLLLlxsm8peXdcAUVzMhyZexBn1YXxYh8RClZ65R7RH46c1JZ8WHMKxJDFN80
d+pgZCDL0tZifRhHVJZ9pkUkgFAoX6eZK7qIuGFN1GO8jvr0an0svG5zRdjShD0y
KjTcRwa1B7SHd9E1Yexi49vMb1gj2ooMM9FX0lGBE67ypJvSiBLzteh20OcAoix2
3l/js/mbF9l5ysqLUHsRlfIE6ILmxlT5s/20dVZtfh5mz24Q2PrkKGfee0lINM6S
TG73qnNyJOtieUFD+GdfH5xBTvHI8Opw2tse6HSuY5H7GygfsSB60fcCh5dmMh9X
re3zsLOtYZJ5hgdERyopHdLbv6GJN2384DwnSUTfOYP7vcAl/D10uio0VZfckTgE
g8ZxCPLfPV7BEg+aZVACD/296CJlXltMVqCeHieSnKnXbNkQqXN+ECsedyPicGBT
o+oL69xM5/H4WBrUORrHA7sZelDsXTeG7KH1sr+BRbM=
`protect END_PROTECTED
