`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCaRDzNreVc1m06pH0w5Vtgxl6eeHSOGrG9RoEHdSQG5Fm0aslGuI+5RfGTiqYVf
OOpeSZ4ngf2QwvvVTsmFMM6eivvYIR19RI92FgVun9GVcV+P2WzKVrkCtJbn++LV
itVUwRHGyVmU9V6ZQkkBL0LKtnWSVGjHNqdrf8RtJFEmoeDPlhBwWrFoObjSyNid
WzBs2/nhQMmVMkrbJnPXETQ+a/HuWkwYSOqLxTQLAEcLbwxoN6J1bunovf97pj2U
6uCMmmZGoyQMTIsdqCNxBk+bGB3YZwJTz+rq9JrkBR7j5imbOpSgjeIj9CGD+m4x
McBriw+nYWj8rMLN3zAExb30Mb/nmKqlJKuuxFR+0e7Oinwr7YO3JfsazWObw47F
lGgouDY764GgBZcfuShEHr/32plP6mNcN1Orrfl80xhZKTqM+smblR82SWw6OHZ4
V3mwdpi6PzH5P0K88e+5fAq5rXZx6nDMN69eRNx/ftgklglKz7pmTdVjLQkzNG97
bu1Ceyoykh6fD11w+u0oF9wKRF22RwWqoMpGuyc8O5K0AkVojEYZ9ghOPNyDx7iu
+tMBUZRr1O3AnaTKbLJ9Dg1fBrJfNd5+P+LIEbFBfXK59ARFxt6K6LmzVe0RD4NU
1q2OVylBSc5nKZeriwuWsUNrQDBaeEoeZve9QFSrVYOTKE+wSXtmdlOr58x7ktUs
1+anJ0jFazj+idf0/ZXofimHPHz0WTrzi6dyn39QpY5dJgpRSRLJufBMcDRJEcZZ
+4Kkcu75HOSCJc2LCpm6m/TAXe61M40GFLKIrMFw7zXcfrR7vCZBWm8AOakl5q+M
LWOw2Hi28MehQfLkNXP9Wt6nLQVQYspOIiO9KNgqbM6uXvXDqWsNtRTvmt7PwJvW
DbyxG7TNn1fDjv2VsCzecDSUIbSHKBWqLQUo6PqIjlgC2rng5xnlLJOeD8pN2YLo
jJqaMB5Xrl7Xilp9jXZCGk9cK0t/jeQHkUiXhk57TILLdukmP4GijgrF3uiwoqi2
HuCNYY8l9m9I6YlHmz9CQIfFE4TAwFU+iWQjGNlwiXtwLdNHVkvmfNhrhLXMmab2
NRBI68SfbcbB6NQj9GtZCWNdc0v+TOABTdUnYldTqOOTNLrRsaS4FytgQjCLBlaZ
x5y7YzkYUQx3Sj/9O7ZmVTPNdOW8Lf5YAUtykwK7uAmZQklfm9Pli7l2qhs5OiMQ
yHkszU0jDAfBziq+I8s3wmtZPyYOU30eGccoSRla4oLPODnisfbSni6OYDgJF/RW
5dPtFNspleJo26bMRS5nlEU2nA94n9W71007WA4qlKsZD55kxRQWsLab9M343W3X
KbwsjCjjL/ggewar7sVwuWVsA82m65U5pIRCCSjOA5kTyvpcTkeLkJy6rSOomvgz
7B9tq5sZBkY4zjg8NkShrUeNRZtOSCwHPTGrVa/pqUAdogFJg7oHl+lO4TYcy4H8
a1pSo8RJn6xmvrswysfAJaXvlnnn/cW3czoefpfuKWgekNYMw9K2u8d3Aep13OqZ
ze0/kBwZlKVi9PSZxxYUWwyKTyX4KDRFmbHYJQsjA9ARaCVlCzXfiV47ADO1kVtE
fYL16SaY+zzKduC3NeByQkyikcskzOFzXnEjDbYbBzeg/f/fg8n4O/tTDvvmcTwO
jltHNlIr1Ycwj7GSeKOAEnx4++jjxl2E4hZvBjNxsB6W3RL9XwEAgR1B0wxTmK2S
VHjVm2mORva6YDkyRLhzEQWOC4bmWKtuFftuGaoujfOcXKpD6VkNJD14rNRig4W0
uh9XIdXDqCzVTxfbRJrL5iClPSwbiouZsb1u3rGvpSpi6poa3ASmZaLj+IU33Y2x
FB2swuKd/02EcNDkWq61oTDcScn+MhdVQ3tLwWbhtKNKnr2VW6ArgpnkPi0onutb
AlHkz1ADYifB7gSqOE/VZp5RSLHs6TFUBaKStC26UTaGGX01tlgfBInwXxSuZg1D
DwL047uz1mecPT8bfhaCEFEgMALw8cxp8TVr61EFdQmh4PiZOgI3DT2r2koCgUre
rRXt1WulfqcdLt3sWRyoHT9UArU5Y2SLuu/g1eEeEBmJgcfYiouqzngkb6D9mP+W
i+JrmL1PhP7VziXhdgbdzi0GgbVPPo6azTQ59KagcJHJuhntgS5Wtmc+l5glH40x
ckzbUZ2kXeiXxjyu7K2y8NR6tfjjJN5mDm3UXjbLciOPZpLCd/CQuYnLfptNOUaR
G5+1Uzsx0wbKSDx5pA4OKdtMfAJK2iYHhCxHGaImFiPhXNPw5qtUSXvxqjNou4Cc
x5EtEaM3+Fsyf0Lg/d9wcfi2f8ZSgzQXmgvas8PiETAeg82oNYkHCI5oc7LvYVzT
2Pb1r5bwG+gFcP4lgsxYOVvgsVFLIz+bN/K9wyBvof995HSOLx7ibWxeObXB5hPK
Yn40F70p/xYJ/Vp4tHkwNYvF516gaWR7E6Id+JGRcUBqiUwOhC2vtrTF6nsF/b9g
RKnKKk5Kmghq0aed1AI/OdGKjJ9UWSRxkt5yt8sZ9n4j3wMRcAjjP2mej6ndLlsD
LSHp7maoQtFwoiAyzOJNFYEoo9SG1Zw3r2oVHUlSJoBiiZQDuH3pkjQBOSUnicMH
1nQofW9IVBDamHdOskXjHXS5wVMMtfCwGHWhyPsV5mE5Eix4vefW0gMwvFqVoCr7
YjgEq93QcJ/nQK05PQyolI+Jrsz1vhAuGxTwFVWaUZvsKtQXzNGiqISYpOi+9r/J
JqlXzN5wUg1+HAFebi8/aNt3hu+PoPIVcR3BUEolPfE4L2RtS2/64L27TqRKGj4A
tyUw2QnSdROUaJsvJEPRYOw6pMg1IzoGjK0IsUCXjjgImAlKrTCl94xqu8sA7z4A
zVkSEp2tYPwyiOZQ9OqHjH/hbJE4Nq1wMPBGbGzVNMN36C1Sayzu6+m1X/8oumwS
vvvqR71d3enXTM81hjsht0ExW/3jKAQ41gwpQDk1QAdWFThgCijGX95iB3Ol6Ocp
jmg6E7CKIn6n1MlwBiDnw0rOQReEx5jpQuzxBvI5q8OIhlG7AKbJPWsM2bQyKKBj
BKjdSIbm6Xr5chtQ8R1kyFhW2PooYW2oFIOIKG9hyr9G20TFcHOyqAC+35cf58Em
1loDmV+w8tcDKXmbf1BexRJYuFZGcP84K4dBEGFQVJT19Rx0oXXK3yvTBijwTDNy
WJ+Rmfsx3mMWW4ik1Il0UgoKAdszACWfv8ySPbWsFjIj2Jj1Ug2tprKtflPoPkX5
/iLckCk5DanwLfAVF6Gka8Gjex+pfIFCXsJp86l1G9k8zAE67oMjkNFbVbsfHbuP
B6if803JahOdWantIjJVzCsN5GKgS9YA35IjCoCTuuPOIcxaQSk9X8b3xQcp1F9Q
lDAbjtvMj4+8h+r+63xlz28KE7dyKuF/Hr5BvRoB5qIHNXmQKw/GnYgoahTlxP43
8Vo7kiBvKmhG0iolXkt5Mbvouhwk9NLR8hiErBr6N66j2fXx0D3NzZak0xLe5/oO
riiaIV9pkcDo9ueXGZKWULVqg6i+qt3Lzlv3jGi/cViQbySSc09XEOXBm2lFxyQY
jzpHo87OGDhkH5OGBcPsmE0SRTt+N8AGVCTsrS8SRlttKabZ3kmVp7e0EebMBWvq
v/ZysgEmaasS2OrcA8x/mGYQYEu2hx3zATJLtA9y+2e66OcDCgIijp4MmhQHzuSy
p2lfNiNmcMgbOIglIU4BhDyqASHMFr00rpOQKNEb/67ktfiXEnRFrhwr7fpCekOg
cp0FhcIa5ON7XTvH0VopN/taO8uwHY/tLBkpjgTJF570xac+4kll3tnT6eJeMiYW
GIvEb1CT/DAQ4pMT1Ci6SZJPUgm/XBSosY7tFbk+Q6JGpHveENzmMgWKPbAVHKuQ
+esbE/DqpEI5b0bc7sVOfh5xu2IfPFdx1yImdccwlKzxSdIV4sCgxzdaWzsIL+WD
ua75vHL1pLhl+9uLJyEjvcwxkCu1V4qU17e+ZVRh2hvRYAwJsH2iYDWEToRDFKlv
NVR3t/K/iJOsx5XDRhwPDrKWSVIQQH+eIHpPCqWsQ6TMg2iZmYAavBsoz9pDtyQQ
o0kBa9wP/nNf/V/L8IKzQhZezYO8XLzMI4dXA8QpxKlFvFUenjlsy3+IJNSNd9KH
EwnL2to4c5j/LAFhJXSZRxHhaqdT5CY7MwsgTB9UeaMOv7anwP6yL11ClgRHrJuf
H4V7N1YZXg4V1S+KwDOVter4GPG88HnIWwouTWzldocDkz6DIpsIhx02tCbJx7QR
rU4PPqAmtKkpwrbJBBVNP8RUoz0BpgTWSpN9YzybuYq6YWX8Y0Q0lxbVLi6gfOqa
WMy3ZWJxyE9SmFwSOtHaRUSQXe2WA5pd5ufeXaFpArkhqJ0lzws80DXF0qlsNIDn
utjtu6+1KrC6s8bAT5eu4+mEr7gbsM0PfRXYbranBEBj2Y+WP1ZtRn9h0ublm0tT
16/cFRRP1i4nWybGzuabBfnRRHg0cJ0jUIezkdwi/IPhYQeTowaiZbOS/MC5vIkW
qjCCbJ8fraZask+tf5xCCjRLYcnlUnE4hCX7seL8Lub8+b56oiWcflyHeilDIdd3
Vv1nKM8ykBZq2GYO8wp3NoZF4Wu8LpUW7zoUz/+ITsJuL7HmewfKhy96h1RokuKr
g5GIJE8/40GTumI3jrfgDpp7wHetdof6TuTneXtJ7rCvNyHH9M+KJMdlloDvEyC8
aeSyN/t56LH7vPUnkQjMtGdUujaD+AthNzSs4jFFSDT1v0OOyOQqpedAqrEGNq+u
lF+ocL/7NqLOXgYoscyJwdJ+a0nqcl2Kql+UIlsglyW4xJRY3USa722vn//8hVmV
CtNrQsY3lOu6+dP68NiUOlrwTseeMzJH6f51PTR3MZZvu39PtPYfH4pv+q9uHuki
FIBr+lPl+Mff8mbR/rXWAS7LwwFYRJQVZn9El21MYCY9HhBiVl7JxmPc9rfZq6sM
pSo/76d8wNmFTHJjEgHsvxuIEeh49Ur3o7fGu5/aBvVBGMU+TIYv17CMwSpL3Ff2
ucz53mibnJBusjZC4XWvaDQofM/pTMzQjOgJf07/6Uz6C8VeKnzu5yYzHO1siOce
3T81jGHlrp0yQy17k41eqVaLfNY/wQgRts8ITTtd29wP12xKjNOF/HXWmuHp8a2U
5xRNQTP9ao3v5VfiJAyhilchOd0rmI+Cj2KnC4ZIKInSEVhXe4IUWuyXVLC/loUh
hM7WnW7IM3w1KAE68ji0ae+BmRtI4SSFDqkpwVcud+CWPuSWQTGNHPV1kyanG2ap
EVN7vaR/L/gFPSYl8aGsCoSxZYOc2x8sbkJutGCZsUwH43Koq4nvEq1L5mCHxGaK
O4henhh6Y1OwgiOKIoLzonXw/SRC5iGmx6V/W1T6U4ZXBvuOLR4zmUSJcKT5IIOC
LAntY+Oc8xfWASsj8PD+izjYalHOwJlcH44VIT7HgSouyED9a58CqOb8kdETeyht
MoW+gLWl8ya5eWMuqU0eEtzKVzACciQD7q72YQnV+F8nAPLtT1CxurRkHM7Abm1z
0y+N2N/sacsz4oLm9L/SXdXl02W2Cic1kTRmC+ZNV4OE2ntVrA2onueT8FaA11PY
tGUZ4+puZTrn7QWm7x8RqoPr0OufLMd1ecXhBPpwKSvdju5zei96GgtsvlzpZ9am
iNtDvVBD7AFFY5i2kIEKKFLfbGnZ9QOMoGN4gkDCcIqT/055Z2cM3BkgMZ8FceRS
Ln68cqIzep4KymoLWEOLi1CebZjwFrx+7ftNLWnuEunmZA2B/2DUb+HeSe8+9h3K
kHdjQkkh9KIxUS876AOucDgDfFEVKNg0RVosCtH5z1NaURpPNSe+txIP1oCIopSm
2g9tBarVlEVvabQnpFIeHm8zxBzkEMY6PcfTEkhG/qD8s7RpqaTrlpA1NUpMqhGk
qSRstE3R713K9/avNv822Xz6PqUlpuqKIfKnvspOz3yYEqFvexYka6GmFWii/jhn
5Cr/HAXLRXZD4LlCDPhTpQg9D85vya405XWTgUeUAZCJI3uy6ALYZzIUtAT8uTTL
VYouzZ8O8FkPoYcelDKc3A+nvLYl128YB3UdFYy56bhU4TS7OhMM6BMOnu5CmsME
Y5zO5RY8f5qQAcg2BcjOZYGNfYzsGaWnJoUOHwkDm+iQND0eZfkKCynHM448HcNk
O0LodGCJhv0lIttzM03cM26bBdcNQECrZDRQZJyIrhFGoQmIJhXZJ5CW1o8vp45L
fCXmNh2wju2KqoDcKCt9+BL3ur95djZFtFpKurLd/e75ajUHMyQf/xuYKX1xXI14
ItuF3RvdJyc8jq4wLhvqEwv+9CzVCgHgELIrCHAkRgJ3VuTpT3xLc3Q7LUoa3pcW
6XjWopGadkRLRdbjHu3sRx+JCg/i+Gi6WEnC4ZS5UpSSpqN6wwpy3MwTw04nD7qH
HVGjAj//buXfJPhM19IuMHQmkHRLaGoCSt/CBZvgxcHhi06sWBpW2zQN3+lgmvVq
v8Oq92xlu4x4NhXh580xGoC0qbeHK2T8JdJIVkIx9cRdiJ0L0vnclLWDDLTzCrTB
yDauzKAiOXocR1GhWYX/aUYwS4TX3m6RvHCrvEPx8mKAw48+aZD5UIVpdWf4COEr
bryAZoouYERkbvGfQwvAlgu7GHcS7j4k5jN6jbSQ13cgTOmWpjN3eIF0zmVvvAqO
cwZSa+0z5C4xxRQChjYveQNOP0Ph2NzqCN9RGno7zVSV3KvRI2XbHonNoXxN9VNh
58bNwmVKI9sb4k+cejIU5sfJ4A8gl70pSncgDesqXMho6+6udfweaD/y2evA5lzY
Ez38RbNkqU++Y4U1iXQou5EzLPZXvCpE9NpPdW8zUk2gq2VZQitLuUGdfawV2srz
F0jkVWOCj51ZxYn4+7UqCB72FuxRDobIVCycLCqwr6C2oaqFXJV05tDVpY13M33x
//QVY0CzYka1gH6nbc2abggMEZPOiW1FtwFyS0DuKGP4jOBAAy5908NtbRmSYUAu
IvuROGkX5hkeRJNCMRrxHhQI/0E0q8OEjwSdJiWlTzT2AUvxnqDzGIUtvxoDORhR
MInNsTPavWNklMw5K19Wt3jvJLjVuEFAoaRRqn3meJADjKOguoUBbj3Msi4YMRD/
PL24psCsNf/rO15cIwpGfduKCe2GVuebeNgKPCQGvDsw/YKGSNkIbWnkprlbpftP
Xa1/GtkyJy951b86dYV1p7RIQUIAvWlR3Y37sns95gsL7Nbru6vfBgKdqwKMsVXO
2SqnionTn/RjpTwpuRWpF2xAKx6jqYqRjD8w8r9KoivUaWl/hsnS6Jv/CskQTX1e
oj1A3TF3mWYdGODZVEJrNJD9sDQYws4FrKXY8msmhsBgQ4xcoPQH5bxd1u+7f5Gn
n2GYpseI+eQULoZrbQMUCnTDlxLUOt5e63ViK8wyAoMVme8Zjzm+pTKsyi7hRpoi
S3zdnOak93aS1JjPA7ueIve1XhBMztkQ7T3vN9qadjDDsKVao4fl76CE3Sj81zUH
NbC0oUGeRDas9/DoZXQMVjvRD1HFC1+2noINGqRwAfGZYrVFmTDGWR9h9nNL4E2O
2E8dCpbVDWp+LgA9ID2LIt5GUSNW//gi6D081PlwF52O27R91ObqUYvUVYxm20n9
ZSOogbED7iTknmMZZk+hB2aa+OevyQGoMyCd7XkNyqEgysTKVZQQNap5LGvfPjnq
JqRQS0FbvzA4JHaf9nx53UUc/qFj9LfkMu+IoDFNo+USC8KMb7NO0nmgwvfZUf84
7ziPaKegT0VS01wDiF9c0xZxHYsqT+4bsP3iCBNa+aI22Q4b+b/ZmN2igar20evH
vcO0kq0LjNOZiYWX/Ft+kL0Cqw49VUSPzo4p/1MWqRgwv8SF6GeOEBTh8AZ+S/Hh
KnOOfICWgLfC3WKFNNrC77o5EgBA73cywcOzWGJQBvQMkmRHK0DnkftsbAiupIup
M1QkbwTkepy8+OMCJ1Vw1AolySQwPtd8U6MUO99M67sl/2ixmVvYJBxg1E0y24gg
i3I1szbsxAWymwZGU6BtFO9mcmOVJP6K6Iy66uPnCuxIw1WeJZ1qoz1GHMnGmbmB
xUblIDuW6sq+Ws+kbOpSvCODuYLlBIywgfPLoTrrLSACmtqgP8QCFNN2FmND1eeC
x6qWU/oFQBMcnAa9pQgtXDluKt+Jqc3R3CboYySVdOTsWU8bSaFfp2cXhGP/2IIZ
m4fticDXdQPPDYF4tFeM0myZOYXczWr3WaH/cIAIK5WEV7ssp5nGQHBAUnXDJmNR
m+KE+fAt4OzgaYoSe534J9emAZ0RkJKT5DIV0MPeSLQPsxw4s+wUWF3BEfb/rIr7
q+GCX57s6Bc7DP90ws5dMocEIr4xLbP4PiSPv8b0gHe/h4IPhl3Zs3spE4dAEXs7
zbIGA5sYJgzhsooldlkSI9AeCIcHtp8vyEr+tgHyzrbPPuGpxg79KgvaWOgouJDU
b8NBeZoIekNIoNBjsqG8ryMRf1MmxBj4BGU62wMiseJ91KddvcplSq1d7eoDAbpS
6dE+lJ/YLdAfbbJA6TfXrYcIOhrN82NOhFea9JFFLnatYlop0K2rp89O2PFtjgyt
txabpt/jHN27jDQF9rQRprt8IQT/AS1FROwgTq7IOJx6fk2avsaWr63VoRtif6l1
zPTmx6XXOHTQBVuF2ZnQD+Rnf3PzJbyHOpEIeiQaBBXD5H20Sk9xk1UgQGmbXgtg
oOt6Xzcy+DW4O7/YXyGeufQLrXrtj37pnypa0mIwj9BYDXl8yl2kBCuRKSXZd3gA
4hfPCEO8Kf76I6s3hbib6GL09p3ClBBpiTpW4JnVnU0TWwr/1lvN+apBUD6XMjyb
Jw1sW4Ros2jj5PXk87lC34uVDvv4zhasiYce0RZjjc0uxsB90QPgFXxg+0EhoOqx
a3HfQPOyOrPva62Y+b3OejJFpJx7fjv1py/P+nsF+TI4mvHYmbwdRKVNq1+C7KE9
b2Yv9NdF17SRPcaCiFMlzin5n45E3PlvZugDKbWj7An5Sp62UmwykYhx1BKBxyTf
D4X0DsSccFFf7utp02DseksWfyWgSBRbe3g7KRFyBIrn1VfR3IBQJCalUHWqYb2+
sJVG+EYMzFCsiY7Hoy4A+kHPzYJmBaiwhOMTV/81ZhVsPZCdOaGy61HTtl7FkPhv
XWTakXrHdgWvhVPeDU2BBKJkwTVj4gi0c4rUeyHYh7c4PL3xisQTXx1eZzb36FSq
v+FdRhvD/BJuYXt97f9rDII9AA3QkpOrg92+CWqI1j0VZ0rpiaRbToUKTV/nEE5e
/qIwkGe3pkbKUAbfMSMgn0euBmWgq7K39ntxj5qRC595HOX7iWkdFmh/ku3AXu72
l2kRH+lJx0HKcpTlsc5pm6xE9FNyAN0q9S2i1JrexeVElyfR9dVN9YpW//hYk2w5
Npd7ad1E8uH6tamvJDRQdQSM7qmTBeB7gvsmbR9tAbKL8OkyhDwOqjWi282vEu+o
Dv2MQid1b1kuGmN1y9ITTD1Yq7lBGr48USYGZbAEYDF5uJmLGNjlv8A0tz17uWn5
ZEtAz0W8sKW7GBJ+HChNKBlF3o6bJBnl0OJrGtoGJHU5IcfxHNraIHYsqmkNzgpD
ERtHrGrMt3pXlvVUDLsw5JJIZNhRay8+UvthRcnv9r/SS9GyqFcdAehg0EdYPTRE
dJrE4G2e2VdQYMPy3+FyPrNuE2bPEbHHLAk+pZoeimm8tkIUFnEpneoJgOGX9Ax/
FmdtKkiTxdVvkIPQAjqoQLtnz2Ilx+ADjqh7IjuHk0RLqDFtUlxy8wCpqj1/5s0X
ElT1SIA5xcSJGxd2Xn37Cc8NpXFxcZ4lwiOE2YFTHg8tY+fZoYnDTA6YEGRZyYxH
7c/rNr2ukzkfGqk/fX2BTKDKEGjjNzPKZmZRZK8sMXSv3gfxuxE+KTGdUBHjdDYK
EhpwGaCwZGvCI0XzrQOsDBLCTTjjw9sjOjGIDF/xYeguTMXs3Z1SUIUBkWZpAqCT
Qdfnar0aANP1A4xI783RwnaFmIXw/38N5AiyjsvVsTWBsVlEJZTSL3NajCEAHAel
hAnzbmixd77FeHC+FQks9kqq42FSz44ZB99TNrNo3890EbogPKtOOTyH5y6PI8dK
LVFFPE4srKcztdocrI6ENpVPsR7ftZcozWHP+mjQnUFWYp1MTC0KP4riCbmCErT2
UHSwC78dLAFxLBaIVMUQVTZdysMbJlesR831QXyf6reAdxUA77hoheqCe54Hot8L
/MHbpadKu1b6bH+ftCGYYt8RsvZCkw/bEaOw5HPskWpO545W3juGau7Z4WG8wVq8
+Ubg6FGTzl9gnlBGdtvxfcyqcLN0w4n7BpQj4SRS65ggbsE0/wRd7h5SbSTbl5nH
lkvYcssgJajgXOWAH5Ufp43/iCiZ1kULT2onWaW6ws9fx8xlAaNTqo4RaiL+kEoK
6FJRM7ziPWSASNt+Y+FZdp43gEAnahb8Ql9T0BZaTSiZheRdC2Qa0+O6lJdGCaT/
YikUJMVRseTBXlU3EBj5Cvscfdms/WXY3M4I0sZTISa82T77wNT8WCA2IedES0Gu
quQfkl/fA+uhMSDy3eyBsKfxKz/AU7tqovnUT2XgOe75Dq07LNWXa51d2OHg0H4z
bgGjVbijOSkeYKIiQ4PHo4oJoKdNb3TnKUjzPTcQYZEQm8oGjhKojzn8JotiGiyQ
1ZWzjXQFJGIsynPPKSOJ80X9LlRRiCAObeD2moTvCKmixYnjjYMonVwHQZJKwuvX
dkDe9rNPfTuFTfdnw9m1Xo8v14i7IJ3E3e4wIHGE66k9ONpcHPtdGIvtluo9uOK+
o+mBKRV/bkvmExwCH2p05GnOFrRygjTgYOClSdSQvei/8avZtaB0IaD7Sbt4Xoxi
TUohMMiLPZCJG4AOaJOdgP30iFCaXir9He37QGsYG1wPoBv16US2aziF8gWwQCMT
rUpMdlnyhbtFVJnRDhJz7fO8YR21as5PYPmXfau00rGuAE+bbedsqdlvnbmVgAFV
4FegRSMsWdKT0wHSu4GgNIQPdbKxZD5w4I2/fqO1ceV7HeZsT59qLqva3jVvXeEk
1MxJmyFthVO9Z5/3hjpPUgJQ3A5ny4umwhy1UI/cl3g/LGuwm1Ne+kTFtbyBSfr8
eLDBsAfKbqC7XxHJeoedd8k+v7XKi/st8hBPTx3yFt5rsoWsdUaWloaTuHEiLTLP
Y6Ks1oCIDrDAP9WaNfbdO7kyYYitEYbCgug/jsMZMmwUIGx9+/M5fmd06t0D99hE
OlEihGcLCO3GY4gm4VCvOydi/ZjemvqYuGO/VoJCAG0z0zLmfrPaL95D+8XcDeUx
ZBq/jiqqW4nWkVKxJsGAipvEPZvZgpewzA0QXveDNLuqxhW0MdHzwUatC53+hL//
r5VgG9EEuB9JP0T/pU9vvWfbGRSzmjgW3rL1OyvWx069rVJz1ysZOWkcIg6vnVFg
d1l8WjQ4MSt/DmtWF2/kRg1JUHCkbfzznA4mKYKzPa12VpwHvDbXS/Zt5YyBXG+v
iY+uPtnqD5g1TheMw5tsAxJEGAdd5gvkb90jg7pimeD4ouZXdBB71DaGghBTXoKg
MJ51udDHDlsIXH1k9wf5d5vUUkXRr0HfvUsLAbXSoM+GbO+rQ3ekHfjLbRXjv0Kj
1VFyR8pVcTOiZ264w3mSkRVZQGzskg+/2XxxtFSkBKcuwQmlpQVtQjfjr5HnUpMz
QX2J4MPTdtcjKS72bpsE4JGjJNqAgfN6ebBuTbxW4VzwcE3cW50SeVrff3SP78Z9
VA6d81Y6RKpX9gfnX1iuj7amDsQDp87R2qBK6DULfCmMQ4d2LgKVcW/e2/Y1vmQX
sKi0ZxoXuCifRFFdmyfrz73qJ97mrv6FbUSJEzH/GFVUmxl/oINv/zXTL/Da/BgZ
T8uMF9DMZNmL3jjiVtd1jE721Fg0f1ywy8zp4DkA82/M5wJDviiscxeIZ+aD2Pux
EJpsJTAVZxs2KlXknkMBBCqLiyWPAUsmj3NzeTTO1zD5LsAVxUBGO19HOcTflVIb
Ppq8baOZguQZuXs2MK3qalV+xMWPut1GnKOpIc/313QFvPwbQdJUrtXTCICxQ7Lf
LR2Ng4qmJEudsI3o1pli21BSvWtaETC4QVfGj3dnt+Ev5OSVOVSfQVmS7N8lHysZ
BeyJBewy0FYCTvo2BTfHjFLQh6VgoDYY37GSnWIiiNCeeYRLzTZQMaT8vmghYA4/
zXt7dcZuNUQwVxQmJvOnAeyWKBk/ma2wmPYILWFVi47FGfEn95EMWG58Ve5aILtH
elMZsHYocLEq2qBIS8dLLIv2jdjN/P+1+dlhKD39kUG/Lu9majFlu0cerC7EFLI2
sJFEsbyPrKT76FJG18+0tf0z5APkdzTkBzDNSIb/xwh0riID6bdtDGpEYWrxIzgK
n4TN8W29GMc7RtmKrUesm4HfBWn1XI4RNkpa8M8ge2eG77LTn4hlVjQONEGl5K4W
jCCQ2GIgEGUTsWDFMpZ7nQM8l+XNt6uk3WCWTfEsKFubiI8G5rHbs8TErYYjUXxs
HmiOeH+cd3e3HbxI4hYwx+qltEOV+EFoYepVRQ6+AbTetVGxcA+PqQJ8GKx0QtoB
06r/i3C+U5DvjqV0nN34UWYcICGz85Ct+rPYJEHvgcTZH6BOBcpLScewjrNX51Cl
J+083s+ChQhbscjIoGFOtIENWB4g1bJn76hlbFckXBcIoSJGx4bgB78TViorkGDd
fjipCTjY7SOZPrD6ELjLOGgaXEcUJRO4lBLGrSysP7vHnOaxavdhTTVuw6Z+o7LW
zO35/LuHlDy3o36+Rs9hoYutRTegKKllXzLvBGmRw9WyPrruU5C2Bsbe1wSw8f8b
qHyDO4l2V+OQ3BhZHfM8i1GdDx6ispTk6OsaFU3P7+22UkwDf4IXv20LbyXnbTqb
hcQ/5TPBpCdLHtTv2R+Ap518NG5UMqnbA6XPWOCnDYahWEIUWRNgimLe3UtGRhZF
cLYvXNhJQGTD7zPUSDCQd52LuXrR7PVjDeQw97buXnh9IORWD4TS7K0K0PVgJejk
EWiWAzWGg4Yu3kEL6skfytvjpkuOGhdrm24l4biYWg5iuMUC4nno+iyDRkADkKK4
BpQ4VrWsG4WlMYNual2L900UF+1KtdQ9dmfqzhnbgwLt66F9IKwSWC1jNBFGMEEw
o6d68BNAKMZcabINv1ahozsOIzppcs1OVBpC/yFngXns3sJWV+suHFsEuCSfhymS
Ib9qmXBUDJzlTgSJW8apf+mQZyuGEEKZtkMFyz9qs7KJMQpDyjvUEv00tWb6gVZx
LHpcrh3DTk70t6MRCUzW92SY2zaEVd/lqki6p961+EzEMl1+iEXa0uTMOnIe7zZ0
m6zVCscdW7Mh/h6AkvNJwYGu1Q/YyxZKABVjwXklBXctse0cgjKFvyRT9J4mQ7z1
lfShj3TTMoAxOAFvWFD+2k9OmYc9vZMAAAuk6Rpuhmwqa3gwUxN6FNVFo75ARmqb
RJM3QdK0NvysLJOd8H1gwWbq19AuChxwZ5BlOEhc72ndWL3hE/Yzrv0hmEFMOjx/
LQYknu2ACH6ez5gnEQPHOPcYasCVx7g78u53MFnZQAHptOu4Q9TaXDqeFU1tq400
nFWd33Qhc/8sSC2GJyl+L/YgDIKvCZ6CnkS6tumB71mLUu8v7d+zsh8yFYX4cFZf
E2NlDE95DkO2HMER7/umEDExnJVDUXpeLJIeBY06ln9wTSy+B6F8plGuVn8RQIr+
ivzfIbsDelIYTYU39H6i81W19uLjJ60VrwryMbypqjhhLLJB8z2lGcZQjIDSeav1
MJ+sFLJDidZTP+JxvcfjuHXzQa/jmznVGVYs8Pj/SohbswFFdc44HQqTpEY17CKl
Gx4I92C2l8w7gsT5Hwco4CW39bWBU/OhIsyUgFALax80k8kodcFIT7wizxQvGnbB
cNGMMMXQZF/CnMIUsgq+bo8dhEAmlhf5DYCoztGFsetay8+Wi90cIh685nG32ycs
cja/jygh3LWt2sREcGxv1Odm/dmmiso+Ix9dYdcf0DyWd1/clHjZlKdAlZyFHEUY
joBAuD0qvlBd3SvNWTYFvU/tSz57J44YtQ8ddm1e8l3ws7rQQvMar6TIQJuuQ4Iu
lRPmrTbL7CGIJwn082y9ET9e4jADYyaooyLum5mVmD3426dx2q5r40gaxt0djHzW
lDreXNMfAMxQ2WDmx4aFXav66InqnelguCV48X8shW1ubVCLAqTfx1hNtZNG1ZRW
uNTF26/U+yr7Dp6mXdkDuoRWPA7qWeeLFtiKzEMlINjIbrjQw0xc2ETRNuUyOZkn
zgSC/CDY90idAaLhspix9+UesRFOFCNPq5DLcd184mmAzE61ctzBn/+cSDLJNjgu
JQ48Mu1jnX3dEqhy8sUQAqPV8CRpiOfwhnxxvZ0ul6U22vSYiK0WGIWoAvNfVpKJ
CD8w6MMteCnIb0k6z2QEYGAcDxQm4mqOEQ43HeRo/BUD5oEyhabrErdj1QUmnm7i
4QENo8137/1/T3qSQoWWEBZYxiaQv1Lj2yYENcbiZnVfNEVmCXUyuviCavs/HXdu
Ib/3cCyBOT9na5AQYFVmdlSdrs73FfVZBKDCqsnZS7YyrvWe1qnvZzYuOhavSDRz
zrDnIeDtN/DaayR8reNHsrd/1YWocviIPan6en+8VVEy30UpFjZvOQD7T2m2VnNF
ifCtQHi+phWNcZcyzxR3bOSCKhZ/1cy6BqAt4VZeZTZhE984qEgrM041aMX7tH0U
o7fPMxtz/Zqu+DCu1D6uOIEO4jliNw1mlxJh3tXkFPTQ7ssNlFRx2pfVZP5PvxuR
mDgYcQFVEeYJED/PCjv5Q5mXj4BVrVOntb7++59W9HYgY4UofEXINy22qFCY36K0
3JTuYHO8IhSoN2yh5dFsDHRFORoPtUgpFkpvMkuRvYak3tmw68xJBVNwrxgbhE/e
PmCznb4CTRCeP6ampqnrxq7PBRHA6AJF8cGWpGypjbdGEazEIjAg3n1UTOeYIoQ1
+3U+W1vdQ02C5YrwRFCrh+TkBg5uEeTqHDCImb+Hbbs2moYeBXIJ369zAyNaIoQv
L97kP0qZkyzWIua0uwKpPdQ11BXwq8LUTAH0RLMqeoL3frNJNKmYCabxhHQQubp5
PYJ5HNqrtHuxobwgfDkB8/zf9l3NztcCNN0zx0Hmrh080lfiKevczj3irdbzRcFs
XIHcWWax6wHcG3ZALNUtiJcOGxEA0WrpgJrn6OcydagCCJ0QemSjs/yH1x2TvH8E
TLRhUDs2veahQr2Hvx2C73Ts2/nVdS9buxmuuBMvFc6iYqt89kl65o3m0inTRDgU
nwqup95tNxKvCahiaScjF9oJ200YRpysG9hNBOqlr6xf+22zijpWy8d+CXnNjmbN
/vsE+LcwCE6pBc8Zhtf9AJLaGeJV4kP8XJRyBjukEdf556nbM+GeFLRy9y5JPRWB
iIjglSviyO8/ARnHsNhFINmBkRUbK3B9HNWdIdeXjYKTmyUIZmhm0qMBRzsVqE7B
3+FYa1sDa5Cw7VpM9u5nQ82DQzcxwDQ0bZoreB7VSHRbUl62SEbuACJI+v/o0c4d
KRufe5sg+C0kksPAtv3N2Z68oto6BvvASX+uJiyMggKvGitqrEoX8ME2dyW7faE3
K7vj5lRS+w4+RFvL6TAD9NpnPQ1l0VoZJj+VL8ntagYomG/oqlfhW+jYT4w+1iTz
k0muFnOSAhuDlybB/QYoFZr+I4OplXrMAZB4ZAUIxCCioXSkMQdTwGWby0qQ0WKQ
bbWWuXo8egSPOF+Zo9enLEvKdJD9GiIyFT+Viq1esMoQGnhTCnoyWl1q6xCM1cs5
cgeim9QmRBm7CPPZsda5bgPm9migN59OHqoYdIgXexLqVITWUKdKIOITTghL9o0C
tMGZ7s+B9d4SiwMiZG0Z0qvAYIufqDvdXJSXn6sg7h3r5yJHAzoCHOptfnLMM02D
wV5g7Od1kMHPRLbslRch9V+/ptPjaifwpVoeBf+FegJW6jGzEDkQv7++9uKf6mVz
0cJ82QZ700o9to3bsqLOquwHxKPijrzR1jT72mCDunBIa+IPPUSIZgjbzApgMmO1
t54mhR5t0w5mVb5yQ79RA8NwDzzUH+7qMbaE2D3R/vzP/O3H4rXZDW9b6seBKycp
DlIv+Uo/C325dKavDs2GWdzqQHrOxVMcobUvRJ6XedF0Mjk5NNMG5vNy5U5RhhoH
BQ0FxBjVhpr44fckWTlOTpLVFPmgbmb7dueyPKNwzkUv9H8cWCl3LG772EvJ+ZDR
IPVD8ODspmo+g/7DWjkwIeSRFEsT8kSbHRKsAQEF60XLWj3va+TG1wOHXkNQd8Ow
YukLaYTEozjtUd+gzDl18KOI+dAEHXatykOk5eBN3VwNzxu/jAYLa5TdM5ib4td+
qe2XGLc0P1qwK7OyZUX6hcvKFUaGLD0n/XoPpP0veQGQTX5PfAEUFAMmuWmXR42c
xft0X6o7f+6y3jcohvTMd2wNdN4C6LlttT6WIpWmcIVoOAQLIxNDHPhVZ48/XTO0
PJVuKeiT3NCy5Q+bf1fdhUu8xmnFjQYgqeJwRc3V0jaWRlIZqwLfZHIizoytTtVy
SKkZQKASFXXhtYUXow1CBy2emRN/hZ2qZoFNE3GyQgsr7cdNoU4onqBoJPmu8ZWJ
uyzZ16g0Y+AeJIBOJnD3gfQBpVA0EZb2ZZcCObYRfpjGGxdB+h9Di8ELGmiU8htY
02hZDoL3HrWMzZrFAOgyaBPVUbjxAx0EmOIsCJNuphVXi0qt9TEq63kR5f/S4rB1
v37Uos3ILzzaB9OJ/cEInZXALsw8C04kuwdn+ecCZRz+q8W7BKkMoikaAIdptM7i
LevoeG1Lv0DFKmy3odl/B8kA0aBuJa0b5MrA5oME//IBwPkARbYcpRJ5oJG+xXJg
SWJ7kEqhNut7smyL76i7YoYM0pbrE27YawhTTC1xwkV+o+TqFQwNrU2X6raRo5Gm
z3aRtT1fMDU+4jQsIyVxRu70QsbCkPq0QUmzPmIkS6CrHM1uQIIepXqm3Qt2ZagJ
teBk9rN0LxxMA7bRU5cAcrIKg6YY4KYMu4vyMcfAZABrKpvP/TsmRVBkIrwXuVea
07TVASLdg4doD31BvBzN9GP8Aet+o6e1p3zWz0PVePwBDroqYz/gCe2paEPTr6e6
F5Ji0IQ73P5WXL/zSON+wB3Azt017VCnZSAfNLRidY1xQ8JfgXxeQEhqY0kzeVgI
Ua6nNuPVI+iGAxstZKy7F0bW2+NNMHYNx3g+cO9Au1jDH177Fd/vGld9zyyAOcwG
FNJvlVOPIXj1pKP1Du2agEbJ1jHe/2/oLVkag8H48yQGL9Z+UDewCAw/3RNTtdwF
V/mg/I3qFwZBSgQo7d8wlp1VhdSjLwidhMh5ChlKGmAVyuN0R8m5AwhexZUcOsO/
WJ8K9ml74dxJ1pqWpCun9vRoNz2urwvX6n16riLVF0ieKdqpOtq/3tiG+4wCcKKi
F9KqCecRvLbJxvcZMNDdFL3Vvg84v7jNRooswPuJCM1sDscXnPmfTJ0FxrsYGjR4
KCkgtS/T2twLHOu17exs8cFO2WI04o3L5OXxh1j/jdQoAv4jsY+ENufgy5aRMFZO
4cLB101zaoD9evdXm1q5n99z5X/zmbSkimgVJphF1EjzreR1jZWtL/M6i/d3gik+
n24z+3/dBP/+3g/8QKZbbF2fZhMR+7AKWYiXIlfiWRDaDFgM8VMEBoef4Esjy1bJ
StWhHOTci+hMp4UdtayL2CObzl6gxQlVGaCF9GnbDvCjf7y59i893IBq5w67AhDn
MyqCr70F5lELJ3plMeUjaYf80TtZD7v5hrwg/9PEtp8Qzq7FgTV0U9VTtKj1hSDW
TEKUSoYKI65yChxo2pcsTQQ8d3Fe/mKOrdvH2PTBX9pRlIo9AWycRHuKMInHQhj6
qMoNVx5FcpRQl3fSCk8GYEHqIxuuueLIkMTYxQODo7ayXEAmBKDVsxW2yckLSKYv
4L2zWWt3Q04mQHa+737uN9bivh3RuUGYa9QRlqO2rbqI+//i+xXQCZOmKYzGEXNR
77ufqDcbCJdOaUpJGcozVfTz+m3yFKMRlAOtwBNrvmGwexj82s+bc/2edZGb23Cl
v1g6IH7JB24C4FUjEliImQRvJXNA56Vw93O4htDmVBnlGQtTQG6T5me9/Wv/sAEJ
gPDM0HbCHfvrllJXaY4oe8KJ/b/HU2TEzWXvlbSlLK9vcejg3Y449h4QGoeyerjU
BMkx2eYiWpNLPuprWxInUdasRkdHNTYIhNZ+kDCykKLRlvXXS0VRFjNIpRxTABlL
V+RBBoV8Tw7nkgGPmSFhW4uxdTTKMfm7BsBp66E4D0Ov72zUQ+lgTAMsSfs0ZqXh
T4AdEAN7zSzdeLeagpiyMWCAxkd+7PUWoZ6eBjTmCRY3UjAjQGhzwwfs9IEQ57UV
2guf4WXDuAcUMjBpf1Zr4/EVBv7Lpy0YWcFBkwAef6HaRn8oXssM4oX4kBsDDYfw
HDVlaJpM9ZQXGRnPh/jLiz3YRjvuMC7BXJ3l2NG+5121oDLnPUBKU7qs9z9xIHu1
Wpeyy/E0MaFV90BGvznCWjMxq+S2po8Ghm8YB+Zn8jy5vf/Yk9XVMzJqJoororI4
vUvt6hrVsciK4AiOTcAYCcm3Xc2stGd07vV7BGUdxuPF6jt22ol84UPRtZO/KXCi
a3foiiztGynBvqIZgu6ZOWv83b/WUIePh6QS2rfLWL1kYaGqCkqGoCPemO8LZnVk
ZJEGgSY82N1EJP6dUtREy4ZDOVBFQ8obeZEUk9XtIM++5E73oULF4khfg25WFaGs
CxfyjyCmT/123G3Ote9GLR1cIC49uABeHfFYQKzficU90/49Q/Yhln94oSJHI13W
SkW0R1ErN+In6zDHk6TB/gfU1ncQhf5ZKEasGs963S75cpSWH7iSqqRrUy6SG0b3
jNTkI2zAvsF9gNUFKfXvBVYWpIu+rULSgu9sm5tw+TfO+KCWJI9hVYjLt7fLiKAP
+xafRlQAFjTEPQkBqyE/C15IYEisSBV85e4DiRJvNg1ndPkLK2m+1oXxlbHhYNKC
FPhbxTccGjw50OjKUy1qdFTvPc2Lb4LezG7lVRTXcwJZq1ttmWtB41Lt0K2xtuc+
rL8Hubvx/3OQ8fPfBslXrPE6uHvbvmrp8Ne0J9jFuGrZFiVu59dq93Xmd/8U4o7u
1fYjIYBrKCFsOZEA4wbi4x+iq3gB2NsWl8lpO/BRVv2UZJds75NQKIbqAvjBB2SL
36BoBaMnHzBqTWXDz/yjDz/qVPKqEuvAec1YTXtjeevDwR/+lfPIEIkfkusDFr/c
0BMhVBMlXfwEEhIHkpnnYJOHnClAYOHWRRrv9bCFq5+hqZgyV6lAQYPVc3xbw0vT
kyezcDWvzewxczaReLGWPScg2fggEJZGZSGSTcWYWLRS4qg/KzoylVpM4cTpR4SY
IieRnh6TCK0tL1Gq2nic8Rvwcl4+584aj7yLJwvKiDpms5Sj/8GsiD8IGY1pb94+
9qDM6FVXanFMAIm95+xSkMviG5AvGik+TRWlpckxg0gcufxzbbu0RBwv2Ck1/Jnm
vsH4W9Fbk5IZXdKT6Yq2ibN9wFNeQarCM5WzsapJ6VM/dPqT1ZGpKLFZ18EGX8wj
kSu/cdcFI072t4IxoM85RiEYcHjwyAlEcqdc8NmzSK9EthdZSKkhX7oZX78n52oO
ATVJF3R+d9PZceIJkCL4xZm2G15lDCM+3QrSnpm/Z1y4tgPfvZHhVrfvweRaNhEs
EGGO86k5hnvmsPVDR1qtLIaR3sZkrPvhT7+nYB3BLPEi6XPP01e+5gm7RVjXkJUu
EMGLd5quX78lxLj33tDqkFnrryIztrGM/VLZ9Ec1mWoDEnpTa9AH4E3VxUmGMTsc
rnYTtysmWjw64ldbUzLPiLcVqTgG3w6aGGuIlPIJj6BEEqPZkowJpBG6RegC61Km
9HeOXvfCsDo/16sogHBEVy7fu/aqIkZRRXOKu3TrF1MHYT2xx4l8uRNFnYYzC9ob
TmEyyjmkBuOQCUl/roySgSWYaarFtXnZdVC28TO3psUP3nzt0T/Hx1YKgyktFa96
QcQKbjH7OaQYfXBQZAfnZ6JbS+Hvq8VccCOT+F8wKnzS8PqY3EcWiYJ3gvNhkGpF
NOYx85+iLrAFZmLlObDerRjemOgL8eutNOJN2c3basltQX1cfpMRfkilWqfLxuWu
BwZZtuD56q5vvSzbYCKUCzzZv2OFCIO8Kpolzu039vIiC8c3D4fVpuamWpjnlR3O
xpYoK7KCGzvIXMLxWLQbAxVFLlZiPqknxLBF/dvDYnhf4WpZby/v0a8ogrG99dic
A46KgBV3iC12QdKDrKBbZICgu9VdkMkyORm4YXpNOSjnWpbIhJ6kvAw2MEXr8/Mx
Xu0e0sRDFF2CY/jLf8svKOCJaFoOzCUNPmjK6aJEQLtKyQePj6MZ8GH3A2xYN1Vj
zI2gMykhRbNZhpcX/YuBxtzxzL9v2fCJnHXPxqzMW6ImGK7TbzmJqyNWMtT6mPHv
ZCuNVN/csnB3OXUfIeLs6lgH5cVJiI81Ut64iyEYixOlc73/YMjcU8KEL4vxfgzG
bgfYkoKZkUIAaEiOeAYtQvbMO+CCmXAXrA6uRuuOJWnX68w/yua50JOEo+TFrGwi
VCCxzJ7g63BgUc7w4rqFnZtybTHoVg82DJFdeXQ+8/6B2UFnouDMEpOeCQpVbO1v
mI317s4Gk+DwV0tRDMNnRtUwLaIede/4Du3cpB6OCZiQog5pyHLv6iXl/mQE1CIV
E4s8Crl55AgEtSjaPCYb53ql3plBfh8Glvtgaa2rW1KD5QjYOwoPigitb2lsoNHd
s6XE0OfGuSvxYOUhB2NWHwv3rFK3fYsAziVyfws5UGTIMY0+U/E44+CUqDtwNbh8
TMbaE9KtCAV4Uyc8BGelkz73BlhH9trcYXRgxfXVIa9IXZBm6LFOCvOxd0RU/ncZ
7/lnJiB6dmgW4W63OzFXAp2FwbRNGQv4DI21eHH9yLVGNXD1KRSNT+yi+GhTu+x3
5tV+S9Gyen7iRZTQNL8TwxigE+xhxM0ZkOwyV9+z6fkz2xK2ztLyMb2E6j6BOrSU
TLpA/y15gST2WxvQ+30vx9FT5EmaYaQX1ECzQ/8xwkAld7kPe49yNQr9k62C+aaE
u8Ub8b2Lhpe5qyfLEgU/zOLKyOvasM7x2wsEz/i3iS2YMWN5qXLwR9OjonNJoKo6
aH5HE7eAHosAXZeeSKxI9m2SGPh2QlPD5DkVcQ3A3Mhg1C3Dt+dn63YF7TBXpBJx
h7dHv4+xD3BE6SORAJjen4ijSRnpU9muuWEl/9SpY18gOMdLxfAyJmnxTtuwF0CV
N0qparmF2RtL+9N11eFDVGFjznFOCIQD6a/4P2OZ5solCWFHcJMeh+mQSKm8ddQr
jxYi1x35k2icsFLBLBhvrG0W1JgyZwouIuf9IuouojH9tYGlQAPgtUs5O2bRAgoK
laYTkV4hs2zli/B0PVyK1g8cnjq+pi1Ivn+tii6ZsJR9/2cNv+otXkF7AnHkmKRF
KWgMFtic8YqjfCmqv9KPlPMI/BaEQSmTWq5LpJaIXo1XG7Ra/sfPA60TrskRnCwH
PAAG5ejxjDMsrUmWzBbsKlTPf9p7TbVNqrwchG95rXAK8nGQ+IyrxhPvXKGSWhMB
1WMO1cgWSUJqpvc9rX9jo0yJd+XzotLrpbyppzve6m73uJFldKvLveujBgXyVhf+
NtIId1BfQMf3tYTUelGHQQPOzP3rC0eF6pprA36qKl8WdzySWPrloGHV6cNCkPZH
zNK/88JxYhlXTTU6aFvS21bvR8TetGsc49Kfx/K5/gGv/jtyrUdnsu02WAaP2Ye7
h9SHDRK9NBj/TBGyrI/yMGHEoMpOTuI3jJtGLenj+uz1bJ8q0GSV5otJuCIrYATW
07Z2Xn5pOOK9D02CRn3qNgBaayEBOdnVXg7wt9rhlEXvsA500m4EtAidL+OIf3vk
a+C/doeE57HiBxV0gWb271mvaS8ashFtLi9SVSI9LWPAsulDHJVLdFxck1jZ46Wv
6Oqd5WPQr9LaiCKUTK+Co0G3NdzfxWuEzTzPLYebZJCz5ZD2gFcKg/U7nM1xhrpH
kp1OZKXnVIFg6GGM5f7bVqcjvYiQ6a30I1ZDKjY/LNavNmvNnm3C9s5Hht6W8uju
nZ7NhMPsa5392fm+pRzDIi8qDvIUFxT+YUxuMHBaY28qq0EhMaYC5ECwJ/R+u1U3
EKvIq1nUIT0XSVS6rr+cgZ3HQybObyuVKyneI4JK86KSM2m9yMu0hX2tbOuDhJas
wkh3VUSnPQPjJS0Bz9Z0mMYCeEEJEr3EKFJk5nRoiJSNu32X3qMbKHy7bVXMkYlq
iDLFtDKanGb/qeQGHp+bkw1rLxChu5g3tHcJjseO+MImEJ/lZo9zThQG10BeaMSo
5QemTmf1bjNqmFngY+jPi0vRooHDCK5LMa2h6gKPg8oVQG72etY9UmZOM+W/9bg6
xclA2dV3pOXfUwE5SBGaBzb50rmnKBThK9iZTZgV0fX5xH3kYboAn2l+bIxfxTAj
bs5XaO4uSFN3oT+HKMWv9NNfSKBbtWtvZ/U6Dcdg97PmpXNIvrP1ovfxw9Y5QCca
ysSi7B4sE5VulAVxDHiyYWZBcmHGJY28rRfGXQtqXQJOqiyV3u3yEGCEbOgRuIk0
Bm+0CFh28EGJD2ToMidrhnhD22KoY76fWAbGtqPvkDHJmJNhq/tIbe1gC/yMav5d
HfzXZChjkVdmy5WjYDgD9kT5375tSc19W+wI6kCCo1tZ+Z71PLtJ8zsOMSUneI1G
mrk0BsZYAT5FU67ZPVoAdg07L66qxa7BnH7JFqfe66em8QfUg52DSwnF6n6xUJXp
DN7pBv9EV7zxffGGXPXXsoZK/elT4r0nVpUjHiGhkwCOvs1iCvpEE6UzttdcIkWK
D/bPGm3x00Avsdc5T9O5ZyEaLsFxzAQ7Y/SQgeFxnYj/XCBrq2OIhqg4Z8pipc+s
dV3TkQyUQE0c1Ju2PUmeMIxbAxswRMIxqS3M8b/VX6L/9hxXF5sXgCrPaM4B+QRn
M+DiM/cOngmVysTsVdPsY+2vZtEUlbmhuhrq2p4Ej0KENgZAISa7jZWMGcVR/Flm
ENIYVYrmK9P422oOtnwvrzk1wMCmnkPRbE4r29AN474+3okKL4geXZRLSxC/cl7h
Gp9YHebnojl41DmD4UbBM6saYF9dSiXf0CaeFZUobwAhQdGSJVugerh7kbw+tYq7
NxnMbGDL2kXnZYhcUYuNkvHY06utdCXNjUCw5ti33EkhzNbjKDBuySycQv5YJrcw
5MAAkEvywVhZnNgXVyvtF2XTESL6vpvtgdd9ziYMdHxXxYXC+LzVOTB3cXfv09a+
KAheG1F5VNuXYeKFMayXnano+595b0ihYR4xV6cCUaC6zdgtNpJ6dn1n9xQNL9no
jLA27AaWpTsBnDerYwViFllsSUNB+9znwWuGm2nn16DA3aewBzcUfi677GuQShp8
AU/+OfbqcSdFUQEs17MV9EfKipBL2Tpf1ZAhOM2eNRRKBVAUTRrB4/0RvyDwJHM5
zPahdKYjBjcn+ILMmHPB3EX9LE5g47WGJj46iKQW1UAGe/MAQHXsxFgNvuSK3DrG
CN3Rr626f6MSU/1aM1YMgfVb0/1xtdmq9qxD/5YfCMKcqeoOAjx0j+Z6yzPq0Xs0
bzDzpZlk1zJhzTjLAnfhiLsjx8mUZhfdi5fZNqLBkq5sr2TP4HrKJOnmcGc/0Vc9
HT151MmA4lyNid3g0avMRrGFv3xeEx3tFudTVpY36lHhntkG5GpFxcKz3eyMq/f4
aXmc3WMfiZA6iHvErr9DIw51F/Fkb/KrGRmInOdfFkH1VqHKFS0s8K3QJCn0bpe4
JYOnZ9l/64UgZ9yZITOwGp0LAqxY/4IrJ8RJhauVfdHkypLn87TvBAW/mWMODVgM
0vB9Tb+NaWzfGP7KsLZE14FqIXxyvqZUIkrfapP0L9X5S4E4UBsSMcKRJnhf43ba
Ev67G1o0DdrmKvqTyjYVtCX1Uc1jGQS4Q22kC4DWremZGqLnn5gNhoWz0LPC3wyo
60f9xoC/79u1jnnnTNSE9NjsBbtOwh2DHYpP1GIoxrjpbfCduCZNSKBvwHxT+sd5
0sDzC2eomvrPyu/ZW+qiFhs1jndOr+j2CZCaajxNLRQV68sptvdnNVB3VEByh6Kr
QEiCNckEakFdTZKKSxLzltfPdLDJJp+GDVx2ccqLguiGkB/G7vu94LYFi3NI0AxG
qC6TQ/55t1orh3ZSEzw6UK/s+df8c7mhvevm4qzD8xBplcamMI8EV+f+zCaQMCuA
ozlvGUUPZVuIcOtIPHttLnZ3eZ1iJpHeasqiBrTg5BTIq5hR3lkxryvVp69BRVBQ
2xTUoq5kkPEGiX3tDiODk5jIdEt84QzkS0pLUj2/DPLGHOd8i6n3sUJBGxMTR1JE
Aw/MysHyBttm2bFIfd5MSe+C/hinEvKY4Cs5Ko3r+ag6Dv107DhjfAcfofzyG0zv
PDOE6u3MRMskziOH4Gw+0avHzHLEE6hh62g+EZaWlumvanw95RCu2v9Kfe8CZ87Z
ejbYDNktrU8M7AtDt3rNc9tnjLbwtUsiimhLUa2O1sSvZeeCVV0y7QadLC3cRKZD
EYUF1PrrGWYOGQbwmP6YsL0EwE1TaaQyFO1R8TG3fz/hu6ikYtssm2RAW6+fgy4F
aZjTailjSTG5iiUg3G0KJEGTxgQF5SUZ71sR95wRTFn42DGbbjcrxmLQPXaMzYCa
fSo9id9QYONBcWhJNVXzZyAVU3000qLgEYegAaPLTeX7XFZTMlK2XMH/Djy3Q3Il
8AYdUB5LqOQTLUYfT6SEu3tFOnADybhi3m65tXR5aCgPZRSYq5+XKTcuD4yMeF6M
H9L1fwzRep5AT3GUVkw90bSj1vW/DM7RN0wcfC2tZ3u59YjOwkj78Hhu2oDy7LP1
N3hq4uX0mH9Emjle9pWfcPzbCYNONNmt1HJmQ6Nunx91P2xP8wKWOnZcIUqxfEDf
ZSQgkb8EXh3BoXugVml9B6qyiqAO2HKRImWMECL3W6r3FF5+6o4po8aVQ3HmIgfZ
nXxRDlvfX/qCLaUf5iyKdv/kj36PZOveyuj7WHYODVNfzGRk9ImH75CoIuu+DRg7
46MTvgG+B9cjf6gwHSR055dHNvBz6sV+8I1pJ2nUhtZHKr+7+XkDxB9SqxmjLG21
kH/j4hQNRKSfkrzIEGEBETq6eOFMd0xEuvVTTvgmUs4LTMK+5qvJf9yAMK9LKthN
yMTsPwqwC/+msbaJEIUtZ4ENDWqIKyKjAb6yOESCykBvtvJcDaQKo4QyuguDEPoI
Or368U4lQxXYE8Kp4cbQvYKQJiudBLwxQ8ZhW3KLcUXxLlbxh0GJljvJLqw3nmpd
PkXY1l+ZQoZhva5ZcoWkIbATo2TQwUWH6Smj46rT/wtj7A7em5Ck7jXzjIcOfIAd
z/G/Iwl04Xns8D8E8CwNzKUpHtQ9vhIiKgE6ZZyYmppScuiuyK9gA0LvleDZHFWP
ol8jqK7LZZ/nuBITqiq0fORHyvykhMShN8SSgcQUxtMkkijAnZHj/O/SlMUUVdtf
aE9pt2dI+vg14UhD/PA/1qCoYejohLHNm5WEcI3uOKP+QGchcCiFDL9noc9g3QlA
LtSv3WERKDnzFpo1UMU2TFBYhk0ad2IuuV5FkHLVeHhkNvwz2WplUv2qaI3e5PHm
7LnSQqvzpDjYop6kXLKxJ3y1keep3RGlogBSHWgsfrsjcxPuUyNeB7c+YDvnDbHk
44heo3LgLNmA4U1LInHef6UVmRQLpGYjhVJ45i6nLOQxHG7ENJt6Rzc96S6ryNSb
OI6F8saHe6X1pSn7/cFvqk8A0peW8kqAm/Vre0ZV+qDpvmPmf5fSv80vRBJZII42
0pxIyQCJphPAHXpr21SA6McBIm1ar4aLG5AuD3WHdCfW0/6nktBMrlhQUEq2qaQU
QIfaH9rZ63je/oPzDFvPaOiKrCaTczjSWDMNLNkFKEO+DgsyP786aA7t2O76zXLX
IzsbnJBcn642NO6pukLCBPdEjfhOefA29LIg3K8hY41wk0N2gktkfzwExXZ6nZGi
zgqDN7h8L6LA44hFtY5AmvzIUBYuysV+E1gTlsapRjUpbmOnMscpxJrzsvr51hLa
B+wQOuDRebnVbOdpbNfS1N/SIDBbrWG0uonIrWu/SXQJAofx9mmWQQgNeX8KNlje
dVpJEuDqnEZBgQp4aAcpHw1hP6cS481DFQNQsc5NuUN97PK0D78bO6MaeL7E0cH2
aEZhFx0hHEgbOdS1K1vflknC4NsJ5BcDuxAwAk7ZrBr2NM9GlP5BgXp+wTajaf8C
k2GfVFZrI5autNeiqwXvBqZGYxQjN0AuXDC8loP3Isfc1P9ROI5o4tMyreIKdTjf
RE8vdryS5yj5DkwsFFMijyQNuX+A7TV8rQXx5yGmxK3/5U/3yM7ZcND+hZnRto/O
L+fh1O770xQxT2lc266F7eR5LF7DNwscHbalusoZQWiYEXHs8MqLLDplW9c0JtOJ
j5+xIRgks05iMrMQpHZpf2a0wslibcrPf5VJjmrFq2TQlHhoOMgLCdlwjvXqiaAg
osNFVN/QL0xIl8oeXTDu95y2Pu3tOGSNx+YEdjluJFXUKKFJoptXeV36M+pYcJH1
rny9bHkODZBqED8+kPKpRYpmg5fc2WNj+Ja53guDVwqsb7VB++gsnifszJsXO3w5
1h7pbQqjecf5p1E1HWcH4TwNsR0E/w2j0/Og13Y1TK5zbMBGZRdcqERaQLKCcp+y
uyjc+bwsSHBJoiOJHgOagZxqQmJHWGu9uiBjh1kWReYogYfzgQM3v1Z7w4Q14iUW
HHSwHwS+KbUlYS0jAKM9k1nw89r+0ciUYHKnFz+/8Vu59+InWGMdo6gGvavonn1c
rmU4ertoYz9G/rcdvdYf6JYeO2NjcczgGyxGFyOtNNR/JOlUWUIr+YCJuj+Fj+f/
DZQ52wLJm2rzuG9oGwZtRNcYUtNchLxcpombY7iI7PR0VZTBBQZw2Py2vJbqOza3
Kvde67bpgeEgMHu3QvMgS37LH+/QEFywLYETUvzI2WasoE2Vm3yQlAcMUfrREbnU
eSpfHnJRs6UMYufA5zvhwg0/tYT2MSnzlrgV7rL88ECNBXoT37YlWrd9q3CYgidZ
6phJDsheMs86R8P9Vri63/cTfy17A9QzF/DXwGyPvmFKSsB7Mkk4jLQhTZ5EWwOr
yFlvJz6lfBdHtmlkZjr2RgaBabsf8Zm1xNygQBwqyGgzTfn8pgG2CeCEDn57voXI
gTS8yhsbl7j7k0PsCyTRYMJfT6LcB72BPc8ROU7+H88qYsp18dyuezNVZ/gsRvXU
GEIg9a6lAkAptn9eaXIIeGvpez3ju4Hgs92NWYL6WVP3Rn0JM3Qt6b5BCnVXymSn
J0fzfio9DoVj8EiJuxdG5FShsPEhsvS78YZc+KsjkmwlpDEWdawW3Xbm9bJM10vB
wu6LvjBy3aFeR8RVb2ZDjZF3Q/lKWlMQoSl1Y4uy5UGBbSSE4ETKI4duFyNZe5DO
xEGbqb+PEJ9wlRLqEzivYv0liMSgekb2O7kAj+fqs5Ytgc4azBLgpao4hv/m7lsw
j7GDxH/rCUZBVONQ8pyfgKV+Qi5cnseCcYB6BARvUDsfNN0R0G99L8VBAHNj1N2M
ZzRaXasECsGbaGA5s7+RZMDv1vSp81Wwr+x+/eXapitglISnPwwBLWBeyv+jokut
c8F6X/nlBBiOJQSeak0a5jVm2EkGJ7l+7YW8IAlUtmv3o6hY4VXMQeDWWX+ioBA+
bVP4tLODbWngANIHSrv/fzr/3FYlFhs9JbZDfMTQgjeEK6iXWIvc0N1PzlvFp0q2
QOoCz45NzXocooUm29GJdlLbuGz/AqSR3N1/XObgx8TXz5Ys0S6Xuhvgl8JuH0Rw
0LYw0lYwTr4ZMwZwYWHTwU7iXSJED6HeuyXBfDg4Uym1xS+xxCLvcFe8b1YTPwSW
BMiepgvEopklc+hhufqSQmkkN5di4BR/+wYfkqhCF/nvP0rUSuw2ZyQ+cCwyTrSM
+eKst4/PLN3hAgQaTYHJcVYPL2nfZisBD9flmEyHzzM3qwH6q/phxL9ZBkvkhgRv
iQ/U3Fy1apFRUMFFRQ9ORPCLHTa7b9c9DsGdU6yrYTjaCmrk7OiESw/lgXRlqTZe
QldLTWUsmENEsrNDUaXPDillKdy8R4XQD9zrFUuUKwv9QCunea04BZc0vr26R0FX
Vnnnv2XOocdLoiUqUmywVQkwogZNc3k0Tc43sgMUiuob/+Q+0QVxxTVt75fi2Wix
36V9GURdKYIoOWAGFqtvWdMWagn7+/SvHWoOCueeQnEfWDZG3wlie5I2f0UbFi9q
eNrZR1ICyZN6yFl61MaTyHxa4VZ8PjBcY+5BaK5GL4ZdWG/4USrSikKPzgYIO+xJ
bpKO6woa5tJ/slEQwPJMG6x5ZtL07Csuogr7CFVlSnUENVbIe0yBTMbbvTYnzkj9
JXTAFCIQc3K83RngtcaAM0sca1zg95zYYInTO0IkMbKcc/eu7BccXO7MhNPL6zUd
XzwC9nVojUhw2HK+vnE1AMumoHoGIx3Hhxkj9HH9U8vLtxyfZJa2VZgbQy+n1rgB
yVMg3fuF8C0OziHIarmZniYF4EQSHOMLARJes6VM8duKkH3G6bws1THEL0H1TrW9
V1ee9lfLyBEQ+IOF8R8zuBsSQCcyh20SPdYOZbfZEW3wfqeeW4kHDQdwSkz7vCcQ
pca7NfWWIpbp02uaa8eXa9KsAb2dypJwnMnP4E918Vvdi+d6iTl/w27GY5QTHk5v
98yX3Z4iPzYL7vagt2bBPctulZzzyI4YcDl2KxS//SvhcQe9aQmtkvGAf3FRqj9N
KUaSoUboMJDOM6W9c5skURtOlwaFLfbB5lWUUrmHY3Ucj61+Fi9j/3+3fq04ZVWK
m+I0kQvpE/7QhRCUr91idnryS6I61XMHX2uf6Sjo56kX+uhgW2yfstHCZ1jzwOF1
Zn2r742f2LCbRuhCqVnf0kAUV3bmy3DwRMbd0O+nDimskfRnw5FT7WS51MJOOKvE
u0KPQwHz/SpCrX26R94WyBLHypqmXzbfqpcZLSv3nZlRdlCowDH2IC50MGBCR74u
y+wRRVnXzBHrbC5QnbyuPkPrjR8gLD5XeZxMJzT7fZKvczJOsJF79rd2Cyeh95Pc
iwn1KbGWANzPXOES7Ae+Sy9yV6t8E2gq4eZ6iFs1nG5vXsRg+5+B39fg/fOPGk9o
moLorN3wJnzwAf/lbuVCTOdLJ9LLxg2c7GgOQ8xSPcvi71ZJLO/mIpvD25heiIbf
CcXazoOFp99WzQHxhCrZSSk7nNO/L0JVnicFpYS4Sel44SVoUJzlu+jj5SX4U7fL
ScFQ9m1L8Eb1SgcUQCfn5mzvN5JejLPTlnP5zUM9TzbrEkK2ZH326VA2UgrZZurn
B0uiiHMBFeRwijE+/Nl3guNP7cFKJ3lCo4vCUkjdj2pghleslQ4HuA8DJAo7zGVn
n97LDr5akKFKtylcLRIBZu3otGjT5G5L6krcD4i48R8kP8+LHJkXmz6Vmz5lX5dH
+V4YFC154q5mU8jaq3SVfBpsuditQQIjP3fGeS4ZMWu1DhXFUrrnVtj4sqAy5YgY
67t0hEjJA5mDuqZ9Et70hlhBF+/jxEvL/ct9AvYcIdk3YY6gisypi6CS1mFUvunc
4sJm8JE4CdDwthUpN4VDAEFiBwbtofUIXoLgeuAuyk57+NpahN8ZmH3QNoLeiUkB
pX/lxSgmGAcDTUjwsED4h63ENsz4c+KXa92RIGaJX+Jg9YjyaFzPpNEMskEeM6Vc
Ron8eyyZ93wODnpL2F/S1TBzMr4LAqi/Uxx1GEOnXuSbzxflx0ChrwHa+3ryOmA8
5mFklL5o1Naoa3xCd76J2NQPegrSowIImLy1nBo+LvfMuIr8bNjYCVMPqoYetlHD
RzfcClS9Hiz/nUEZG/3nFCSDFLqtjyj+9JuO+SOg3N+I5AGdsXWqhhTObpg0ZNJK
Y2RXZOA4IYbTO9fBvG75+JqZSQuzbOXsPmeDXVk43tLfcG5ygh63ObqO0dK2jVLC
ASTxwDNyYEupzEA70SGyab9llPETRiFbeZCjyG6iZuTyh9eV0CzSIMXYWf4lBgu9
NLkkxUOCzBP32K8TXUVmCtDEyKc+2FJWNIyJ+1i1xU49Tk6q21v+JxfQptRPLJtN
eXLMAOQwuGfNkTc/jQweKCkGsIwUXZHpbZ8q+W7pP4IXLpO4Jo/b1VWZ069yYxwg
pT9qWcOgluRmrRXUl8vqqjGN6mNyqA60CcjeN3xstZDmj1LHIcplgjizvJuBxB45
EwuxNnZtUFJM1Tf/GJE1zBz83gHsRqMrF+iYw7Jlpa68DsErB/lEANo/31/oTRWv
IHqrybHBNnpOTay1pM/QsbfcNlyILVAKxQiHeZ/ivPYHt4dgHcsDnuRtJgTCBSq2
DkLQWzCYhQdkfuFDDn79JJhT7X0GAgCh6E3SIIykAlIOvDuAWpL8N1zqQIKJT8gE
5ZTp/BZy9vBO1a4+zMQuqNGsPLiFkGKnQQwPbtxZ0amaAjJWgWkLsFrYMDxhMoVq
Fk2IwabV2LV1QeBDQ2sNYWkdU2ps3QjbFwZqSkiWcI4/4ETPoKuSpVFYBbuOc407
ABJEQ+PLyKSZi+LjFImD4en7EmhuUiI+4Ogj3dXwUMNCbzqbnkPnU283h98Tw5Sy
eSuFDejMHRo0s1I5eDP0uthssAY2SlLcW9eh7rgkJS8bs6yDKujM/vSpV2D1z4BP
gdkeNXiRBCSR/ZG4X+tSBDPDTPUYngp0KkC1UsWMLRm9yEtpSAoCd6oF9m05kVIx
9qRb88mALDwqSmg70NdxXgKNLdgNHBFXQNUdY5Fe/6OcJ/5ZCpS+cLG/hE1dpPPY
IkvlXjDorWx+z/hQ9yuel2bl+tfhpaQLrE21+podrTwGOMPcAcdWZQs6k++U5wmB
R5zF5D4pUcBtu7EszY7+uQTeHhHu9oZdkR9+TILKpWv445UGmz4GBSi/10GM2pgi
e5Pjitk3lnezQcJkAZRoCa3gQr2IiLzVCaAiND+yu9T0WBdH6DG3ur+cAATX02J8
LSQta+YYjTQwpxya3EN2bjGMqOgfhoCQT/RAMZMO6rPl06lfhX1tLz+mLktvMLB1
8YBSRwy5le0Aik3WUYxcn0sdgnAFuJvdzsutqqTcU9EB1PIIwqYF3cK6d2Lb+Tp6
yFJi2Pc34rpWzHx80faM7kA8HjS7Y/1brcsLX6RI7eN6KM2MkvoHvRmUbzxfpLgF
5jl00m5/YnOZxv5BegzWXOqLzcGI87LpP1G2T6ZOE1lzOMntM2DAvNjrU03MYvrC
9AFAecRwD3QB/Ndw6ZtUu8Hj1/ueGXne/ilSmvd4l5hgubxjgakf0xljE06grTtW
zK86ZRWMaLpCjgLuVa2VvKRSKvn+RckdUbmmhO/OIDl49gNVzK5uVDfMbdIm1A4d
Zvtw/WjY0k9xOppPPmYdKwkI8wf7n8niLjB0v0JhW751oSSDW49l86S/O04WDwfL
CC8Y66ZGXQHhgfV0Sfqql8JjMIWG2dVtwD3CneZF/vFuOF68VVv611iJ1TqmTIM/
VoDABnhX1q59Lo9uLIZgg9Z2okkd0QC7MwX/HdC2vvQOzb6rP+/KDZnBSbmkZFJV
YEiknSRNPZabbAENxy/eA65S3Yv7qNFUfj6VBhUlcwef0XHn2uQ+xfGP9r07+cZ8
AR29Ns/lmwqU+0vsa6b6NWezr5B2GnReRW3E7OTP/cO4gs22qCfukF3vsMrfxTp6
AUzm+7k546AqsaoCihlh8oxtICpcH+ZCOIBnX3+MatZzHim6RysBvSdAZiMJbxtY
L6v6QXPv2NYM23nor/RYpKV08odV7PktikWb4eDsLXzZhCJzIwYLJwlpeI68B/IT
5u8c3UPLSUb36NY4gbAugLLxvDUbTg+vKqPVDubnpXnUaFAlOIjrJ+zkkkvWJOXV
pNcwsQsAZXt5Ou3txaw7y4O7jS7FFCrOK9SEqOsc+SaefbAt6f3UmSF7Qm0xf1Kc
CSPoc9Br/QJTloe6JJVtMIKaR0LRFpiDvUfe/9heraxlZxclyzoe+mbbAV5DDAWy
VAgSiCMhjHOD1Dd3IGpvsZyKZeDeoa+fefIg4ubFvEa66umu/kdQyjq9lkGMR6Ur
Po59Qgp/1Zdn+9BUUWIsJMeMglRL7G3Cq1i2DKFHs5Wv0YibpDQVUm0j7ntsOb/R
zPc/IzB9iCPStw0AgFdyPpytbKvwZD2r/Hc6XDFpAEZUl7SgALs4yHx7CMkua7yj
nMTrAjNdIOJdOfah6cCon1X/zkmkXr5Ie/O05lYqO+GTYkYdgTf9J9hmKdidONA7
fV05slFU9enJpI5QdQX+qFWY+LwztOAqc1itW55WGUl0zHC7udLsrkxfatrnYNcG
/APvKZmM9cOTmytMfDQeaWLeNIO4cM2mm9StGLYcIZtWtWKVTFuY3mamJoZnFqbp
r9/KMuJ+csrhrDqIGYepwOaFJQpt4OHb1cdZTb3RWj4cd6Kw9Kiu38jw42yMo/CB
NtjWhxrOTO69uDO2TwKH1CD3bEWonm6VwVkiUrS1bi9A8arKgaTXcnhQy/kCXwuL
+p1EZEMDA4pdoO6MtmUDPvnp460A8RqSGKuFVslDN9SRjM6JVBHJ4Lw2UOM9Anmh
i6LYRBt8G8iwEPnPpfdbgMTzntDLOKn66nQOYVVoHK8G9QKY9LmvoT2WxI2iuwsf
4xaqUSExhc3PaD7PEbda9Ces4JKoMqp6bUDjS1i95ZjFwgw+zfpOej3hGgcXs8Wr
8TrROUWf08Vp6o5nHNI4SPN9+LGq9y6d152G9GVd8dFrHrq3eDUcuzyBXZ/15PlH
UTH4tEzSOL1SAPTx8eImBmBXA1C019/KlocOC5PSlkK2EenWjayu10JgVgiF27GC
x8ODFhc+AjqdKRut8Qvzj2kf2s7O+SDUtZJ5V+xL/fLBIEp4JrqcR5azBub4cEyL
fE5PFnnyYdmz/SOo5QFMp2ZVkYchvfnunmQ8qowjM4Ftl2HJTF8oELLCa7yQ1BTS
eCHh+KbTngylnxsGxIwQ4jgzpcLuAEFeZnv/5vuwJ/z1d0yvP5SdHA3r71F3qTBs
ziT6HOq+3G9293ZR3l4fKYGetwTfFftmDIwfTDAapQVGkc7jYvvPiWVPI+hRK5Yu
vxFKtqRZLb/Xt7FpOgPtapt46OzPziFWR4qLjMwlVaPFSnZDuCw2kEvz3TNwcjJb
o6JPtq1om2QRsw69Np1PByT4a+vRTGJAMwLO69GDsjkg5/WcqBPb17Mm8eonkGmo
UGa7IeWUPZr7EVXEgFJFBHMW1qvlhLRGX/a0LXc6WprSivfVrfepiBrwRycJp4+D
WJBpJkNG89uqxioFTqQn7bQFcw6fjYc9+4V1qxFA3VF9YdtQ23QMdsUF75PvsS9K
2lOk6D/zrVj4VgaG041jS9kbyhVKUWH8KknhCFUrcTHFLPvJ/e6rxjSMObbNkCOQ
JXpHUB69ichsK9iemLE1w6eRmWr7c7v9Xv+roDQcav1ZYXgKSPM5NOWrZCJtVnFc
TM11NokzE356WgUekLS7+TlCqLq6DIqO3wr6k1JOO5DJyOw7zCuBsDcT6/BV+Dwl
Ph+8DiJM0W7u5yPUgRSp/5mNAmUYmjJWtvA2jq18Afw8+jUkasv3OyOoWDMCS64Z
DSjH4fpklD86MStdZaqkR97N/EMtRdNxtx2OktWfCYiDuLx8xXjbUWRV6TLRi3yz
EzllvJ95/uuwSWOkpuq4JOhGugvLwamFZD0f01eFmPzQzOGaGXiB44FuhqAUN1f0
1fwXJ7qkhIMw6CgqklCTO/bqL5ItIovYyDz+gnvVfDF+5F8pXjWtTK5xAbDfXkq2
HqdyHHaWApyy9nBOJZtsEg6KGplOlQ/R56OE+2zlNCpygw/RLfnB0nXI5IeqofBo
Zrd6NUZOHIv12iCP+Neso0mGrzZJklUrOJkcKGf6Z9m0bNgRySfHIH8KkhkXjQ9K
w1hTpWX581ESgmh6UZ0HR0+jD/ZBnoUseMLiVuqBPcCmMzHzyYDJfflXt+Go/n9Z
9YIPB4zcPK/dMoPvp/zcUx7yaiFL1z4n2yg2psM2X0Ga6zGre9k1IuW3eX6NPuHR
AqncfO+FrHcJAqkp1fQ31r5yIq7HGNUwapMiEliyGxEIhC2ZvlSQ/ec8U8vA+msN
Vb0yGchPWASZ81o8d/LtrBPkS26yAezrz5rCSMpPS1FLVrKeLZunf92WLoauC0PQ
lBzfUtQrF1O/bxid1cayQDyVIBxpaLTUcwXUcodIFzsew0Ep4a35g2wI8AsukEdr
HXBz2/CFZB1ACMAhTGBb7v3L9s7tieW0h0HFlO6e2pzmXxn4NUnELIeoZq6mdowr
Ev+PH2P8Rvw852b4JMH5+XLi4lq3LrGWteQjB7L6XiKD5Oc4MHaNpZFMPNFmTn8C
r1huCuJ5l2o+XGNQ0l8CzUTDO1N/caa3j2iJ4oz3WhphFBHKS4Z0sGgtP6xYJ/I2
vqjaLhhkqCdtOGNq+7tMvpIxt5/54XMDnc+DT0KloTgo+OmepGWa+wD3BmNkbBzo
us68jGXFvz+Cdrjbg0GSAMCoIzVQnoaZjuHZNWJYE4UKtIPm4Cu4KouIrf0Lywbd
ysUFZSRI5+SjCLBxP34nEBatdmsvrHE56z78ETDR9yKf/JWkodAxpu4p7pqaoSm8
8HbG/925Cux8fKfOlLcA6HtBPUL4CJjAVyC70UMqEv4h1XhO6TcWRZf+FVX7Q2nA
R4wX/znsVOY1GS/IuspTO8tQjZi1H9Lucny19yP5/jL4k2jw5AmsKHGHE7QjWVwU
aZkj8TXb1HzXzNCeYgarzRu74LakLJ5CJD5Er9Zz7Fg6nNEOplSe8MjqCXU3Vf33
iSek9+FuNWBoVeByCern77dfRBoFs+ISg3wG6sSfH/Gygdv8tqOj0/xTIIP3BHHR
KROXt+pTCOOHBW2cfr6APPa4u2KB5Naenvvk1+gHBSjkqRizDNBn01EcegAE2aMZ
QIJaJsSfq/PCViUoDVXd7UZYFbW0K7VAeIwfXjfliD3yII6uDtQNzlas7ygbP0kv
dZpxPXvNgigSfno2DMiHjuS9Hc9iHzZvxS3TxntGEUq4ednRfdcGswRGsplLiSfu
iZ1HJ1yQT3E4w6NZtHaYHOeYTK1lfw/zZH9vD2XxUzw7HKpiZhK9WMFOtBDQ6+01
S+/DMNUNz8ptizO8xLRieMO1Km2ji0E5KX1P357lL8ASOhY+GAh0l6CLm6BECwt8
FRcOBAEz7sFQyuTiEewct9wGaEq86ooyYnS8HvcQQDfoSwyyqLfyQF1Vkdw10ePs
Hgli098EZPEh4jHvHgF2hf1RjDp7UeovXBxcKPqsOTwNDmnWDy2L2slusXsn9WNJ
ubMttB/XJczsb6R9eiJ0yl7f1gP98J8flagaXld1cnL/SFj/YvZQRVp55dmH3NXC
VrKNjBPk5DFtBhhWryo//nHWTAa66dTjN6qcWIhrGmr+SRwvnyW4Ecfv021yuE46
StKwPTzI55vtek8yGl7WBC6cnp9zg12U3LcfuuFrkjuOTWoctQ1MajZdx19bH8Gs
23atPrhqSCTSBedgQUyAMNVyAnnywipJeWj5+IMzxeJx6oK7YyN4A1YQHYiQprDJ
2BCws55LBS3ZXt2MTPQaaWEJjykGiwnbUQX6QY1RLMLo63Ew3n/h630kwRZn8VaS
ZrwBgk72sSzyo0r1FTbumjsbzKDPfaLC4ll7EJOqtCe5M39LF/y0bYDCFNm8vbko
4uN4eNd45IE5ENYn//PETZbVkNKMmS0Lzms0LZvgUtjrStWriHkhag7FvdnGGFFs
2qg5G0XnXoe/HCnKH8Qdlt7DmIKzMfu6HrjFuLIY8nvDe2yW/6f3DIylQTGhvmBA
9FltEUK6W3rg6hlEBb62yhsXXJCF5i0Cp5otO7uJuTLAKa/1EWXHZHBQMc8JktMt
GpBLqmK+1jQXyeYjsYl6koru7RA5EiLyT/q3i3DAPEecYC6SCtmstwtmWa4qALnA
c5m33/Tbhwof7pKmJqfunvAEQu+1G3CwoUOBF7IhXmwBVsTLvG0Tuq8v7EwOQjYa
cjX9RNWVISjBIShhWj3XLxI0Xf9HM5BqCs3Swa/Gq0tTTqvWwHpt6i5DV7Ix500Y
K7wNS0eyMfMRBOiO6xJ5ZHya5EXMVctotCiPebw7M/xnYfWI6oIIsJVUMmgdFie3
TQprgV+UfqSvhZgQGpVz9AS16Cdu10eThb7pSUJWpeR8KWjeld6naG9ICyo/O1EN
Coh6SrTbHVtqaz3qatyzMxCvbUT46xS7IO/WS9C7jyfE9i9d2BSHoagYo+lx5LcP
fkHWuFLfzRhbsiKJBRCOmkiDUgTnYSvhcs+Pd97z1NCGEj9ATnIjt5L8XXbrpSKU
Rqn218rs3BnQt96EJQZGvZ/rQeoVeVuR5PwKGM9rcpTy8Jd7cRSi53hCgPUQvIRg
BsMgsJCZlbSrY+EcXMXy6w1D5kzw2cJ6kRsbfvUOVwNUtUDUFPo1BctdvGcqpkQe
71py8R/j0rVyxqcTi7ZrOt8+wRTFsUSQRYmeoYmOmgOXEF7JtM50vTS1X6l2aRQs
2yarQWrE4cjopD4BUD31J4I8PcWTTdMk9acCS7Gt2NZUF0c5mT2C6VlI6MBC+SHK
MurUCx7f0opFAamjfJftjGORw38tTmI2SvF7lz7TdUfJLgZpznQAqhsuwUHIMLrl
T/FaqjFp/zsXXJdtUC/na2ksxCwHyTcRSve18/XCRmSgFLLXnJcR/iYAhkiHDYbJ
vfbNN1no0cF2aWFq4IL/8cEbjnvVXQtsP1ECQSMuaCNiOLhGda5vnxvtmEsTDrJs
pRQaFTWE0DgDgKBnT07xHAqRkATtPi0sNZ9GLbHyzBC/fCSnCTT5fQsW6O0ItFuI
Prh9dQP9zINZ3gfMVgQXSzQXMexu4uys/+nbjQyaqlKXYoiyOLga98Z/GzBhmkLM
hTWclN3TKRESmOf37nYexLAMIBwlqz/2KnrE3LqnyYEXKWlYZDYJp7fz0pXdzeU4
NB4cuaArTU46zZEqnzpEwVNZgStW/rcDHizW/V5kyWRvS7aDmr9PwGzzNrvZpCyB
xaS7qSMXR75xbbkL0/gz4CfCKwve+BWijlRpJoTMgwkrXGWkRyheRS0f/FOAEvO6
JS5YlhKqopjZ19hV9ScGD6xPXx6MnJxZY+h2L/Nr/swlGnBR9StHd310EDgqLo7D
+ezHjtaBFCdd8SHkxs60B9cJ+RPHPcPtiDloG3uPCUwunH5y5xzZFBDPx3FQ2iIN
qByCjeNPmPePTF1kWaBY7ifNO3b/4wUzXvOYPJZ4T6g/uiCm5p45O4OcQui1M5rM
vRJvvBlZamfxlx/jdJqh/hCnHhIe/91MUAmMh7NUslBrF99cCNTSCCTF2lP9ifAb
RztvxygXzPaBx51f1fMGD1U0nXt9K1iCqjv8OWgblcLUY23R2SPG1f+lxYCYpB9o
WIKb7SqUI38kWJUjwk3XFnl7rHk9yxm+DD9VKdkG8j9Em0khmGskRQL6lbIqxWaN
LM8HnSsL6nkgSQLcTnTMD5Wa4PtWXKYW4KeNM0M1pF+UcoJ8JEPFNCHVj5nBYBKe
5PxUVgZTU7Xf15U79+qvVT1kgOJ/heDiCXJHyWZDs7oD5Xtk6j+Gd0G7XQwaY3Of
xP9mfjfByCZAAh4QpA/e85FhTeadnKJNHOYd3/gWuoUSL+c+FbFleOfQu21tGCpw
rOmfEnPL7w7TtVE56/uUD+7ja9VYElO5DfeThtbybfc+MAOFk912ZyOZHGsc211L
Usc1XytEGwbK8t/RjlvAFfXNR0p/l0GLvGNfADH8MPedSlSlaVObEPoHgA21cDT4
yTe46IrYgcvT6JkTVHwIeoHy39+ZyyaNCp1x5VlxoosFrDq6U8vBbClOqeLbCbtf
wolqQOt3XRrx6ydTQkjuBVDR+VOjgg8P/kRLifYEKSkDNx7+aqEZAEETGT8nydTG
6/pXUFDRvRVghfZ9r/cbn9Sv0dcF7UsEhhM+82kY3fLdBCndX1ON6l3WdeD2cwPN
kPPehJ0gu4/xmk+yMl5IfQoYQyDc+0uUsTWJ7UF+pDudgJHsPX49muHZzjelaGd+
t6gnjmC6qNK/sFSdl1FQMpxiMj/AtLqvF1bJXQEF8PzjwynT4vRNsz9UNqz2Xsnw
WgFuKzKQQ1pFd/uble2vecdIvnQV0KuebaHBISoIZWof2EQsyuWeYPJzzn06ecWo
izuHSslNe6mYLcC3kn4YZfitZwRLzq8ji1a1a51ng/RIzoRKgNFO8oQ0nQ6OzHmE
YrQVAjdUCRCXdSaxMWQ1cQ3JqT1zHEDBI4hsE0PpmuG6EXDulW1dORFsU17ROGYR
svZqy0jprFG+32+3hjiKoeP/HIKoY0UUpsIsh/GFIY+dRgppq39aPDpy5kg+1I7f
b6eKz4fsn03Ka88fUWKLkZsFGZDs9be/xUy9tr/65aaJXnI5VcnVGuIHEqpOoSmC
Zh5SqzSKMUtmrnxCZJayTUQ77sRJS6GL2a4pGsxpl8tWIuz9UIS/8PE0Q5+z6QH7
nr8a/XX+l0ncr6Yy8YMUIdWJiiPHQ1NMLT5/5gZqDnmqx27A5Drj1r7aYHDTAt4W
PpyKo9jmc5R41i+coT3B2gBs3sfULeYVVhQAO6kuKai9QVYOzTtPFC0OaVyPaFkJ
sQhJcICsuKXCudaqHA80smh76HM57GrpgOXx8Z0bRs41NjD2ERgg4A/A2iGW9KkO
i6t19C0i3XOMMeXMvLSkKj7uEvrNcyFaKwPQr4SlRP8+EWfIDKv2aQ4VAboa4bxf
n/aJWxHf8qFI0OVvNoMEoc3BuY6bPtWcprtsdHnAkA43L8Q7PQjIHzeC9VpNYype
cpXZmCPUC8WUCQe3xnQ8fn4YS3k8oa88JpsaReBkFvV46xRAvYTPYIld2tHYHZMB
x3WLqyzqxt9V9jcjUl2o1JPafMAY2Li4laTT5BBTn/1bsHn8IRrb4PCm0kgMyr0E
cOeYILdwW2u4RQ7RnNsLVoTfuZpvEWkuJCA91kDVkGbspVDjfb7k7ClEq7fs9D+f
6qmoM1HgZtC5+4tVQ9G3Z2vdWSUqcfoycEaIi+RTL8jyRZN6vYYfh8x/LcSdFd4k
YphZYaLs4P+CVekoDobhcJw4houk5pdx9gTUzTYBtBfw68WWWPsJvlR7mbcRJtcD
QUcGgxXp7zOIoV4PgFxeHxa0snGZNK5iQEr2w5q6+9LLEdy2MyndcMFjRtSp1Cr1
wZEjdZlUq0TY38Zk/Bo4YYrQMwXP+YNI+xUs9utzA6j9NmwF6b4if7bWPXTMPXRL
NVXRPGlYngql9odHxYog2ePWevqdDgVgd+34cteP69UTH9PcbJdzW/5Nqqt0SmoN
ozKt0MfTMzegCXuvhlYArESoQRywK/JQXu+bKz/9E9NeicRNe0IHX/HWJzdnKWJQ
oyweXRlIC4apusnA4ympww/ux872ko6Fba4Rxv9J4ZVAKMiHr7wvYSigk54N5onK
9Y0pEARnaEoR8DP7FV186PG4mtLzqRph/RB2OoxKtIKS2PPHfJMsba1dgr+dJmpc
90TMcTMSxm7w+rbkY7krkGqfY18R/mp3DSQgJ5YyDQjj+v//DQzY1l9IcmXL4HKK
0PY1EpxMQX5TlZd/0JyIeiuoBz4dTvXGMlJb4vuSoqLNX1TQvJNjPkgSYzb3NmBh
CB+QmaUx6aejdu4L9jQHFrEe3ghu9EYRjh+RGRCbSTRzQsQJnYB2CBdKOBUG+LUe
n8CzQ2Wf/U3YBYFj/GU/DXHF4MsIpQCPWROcGfMyrCml56Z+W/i/rhgn5NU+LeYh
5m9KSuzOsrGMSt3al/iBVZ7V++8qTZor3xYTmqXNOjXlI/MW1E0Ltuy/QZjj/Sdk
Wo0rPFu45xUShdLibE8jN2jvYEUKAA4o0JY4TPTKR56dzXhPWf+NXR6Ib8CdIyBh
UFl94hiHMjtrzxZ+fU92cmAhCs6+GdzSUP/z+Fh6N5aCukIzFKn/tKfa123hm39g
paPGp8EFz3udBXqHOJnaoL8wXlZXCt4lMOW7kn8NCtl/cZn6KRjJNbRTaDPbF++K
OQFUqBmx5YNZRDDRBYKiRcUmViWqoU970AhxWUaQgcISkDTBWyCXEieqSXUe31sB
cAPeyErdDieHCieuq8NVs64znYCK0eybAaARbzDbsGsXV8Wvz8cBJakypt7zK3EU
JTVqyFb/0Du212sIBOQaf9+N6GlDIh1HHIe7XENZhuyogHnS3ykSbITct1EvgNUI
K2C+gXuPR1EayutydQ8bSXIiOyM+ShSicsRhxXr5SO3ZemalIb67mTKdYecIlabb
Fs4evVKAx9L0oNpREaVI1u320Kmx8GOqf1vf2/bjiEXgO7256Mb1CpJjObDuSab5
2OJxXoTNs6BlAG05OBB0ht2U+mDHACM/SfebES2nlLIrWP4KoXkpwEJqPm/rkHwu
/UfNKG51K6WWr/GOBXt4fVj+fSmy2ElWOTxGXoBowhf+RaJTDSmRJX+5oxtZ1yxS
ndBq8sXEEMMgB9MwIrIbscSv9J5K1PTEDo89RBM/5bHRtDIbxY7MKoG+xfmKdoNq
Oc8aCnnirZg/BO1r4LNrTo6dMgCwMpoCfS3cZzahq4Do8lOdBCeTeQI5oQ83vurz
3LDZSVBdWeShI+4V3zybKsueihBbGQQxpBTf0Bhg+152FbVNiiEuKi3L2Xxo9Ioi
O5WOqwe1INDN2PJTfC8C7tYW/T1mGU21KtmCmskX8qcSzKgT+2/un9y+RqJxIePN
suu3nCYc/m6bVGQ8KEdx4eY1bUMQL1TTnFdszhQXotrPXHK9P5b2PJrDNJYgVH54
6yO3WCMrZD760GwG9DfngeqDyzTJNWG1W7db/An2OFFRsaoWOl3RywpVuHIgl/ZO
DN6aJfRl2/OgTwLmIjewZwexC7ffVfW5KoJRi9jX8HabT61qN++d0EsImqdUS6km
f6VH/muCRiEPV7BNpgtjaynrd7/Dm2ZNUaJWb6Ox30JCW8nVoaCdjZSpN72xYjDV
wnAuo6AUOptcFwExt3LxMvpEyH+HNkXLn+MWRKyrtCm/cYnI45qib/zuOU9mocpE
AL3FwReFMETsmgcbfcqQiyd1keMvI1mF2Gbie2OHtsenE/JWEzHjQl48NIuPGPZf
wwB0McVod6dcqxK7e5J0NWi+6j+SnSHoMozl7G/blfyvW7oEdoEUIFNg19r/XUDc
93JSr7zmijmetC9Z/UW11dbfohBwjU1gV8LtSFstwOTokaXZ2ORLBkufAv3vptE0
ykiehz/mCzXjl/X173VS8z/Zwx18NtE8fxXIHQxD7v0RrFwxtjhZOBa9ekLliy8C
CxbO4Cufcawm48uvL+WO0PKdpP2uxSl3mbgZsga0hVmjSWLtZQ00XBNQCFP+Qi5s
QL/N8HEBp6X5pXlfL1bZm0daKMCU/Z/PivirrV3BFMi1e777wq8xXraTF1NPi9/p
djNZVajMvOz/Q5zTfcKRmKsdm+JI0daaohKOwAsDfJ4Ng/dFPAsnzkpswqjTYJ/E
MWxvWJilG4QktcYOq2P+A+Vdz1paNOiDxe1iO5MgRWFVs1WJv6MFYkevMLiX0nJl
E3HC8Upa2jvkKOamPhuwYxXjmTWRWnjD6W3XfU2oMsuIw1EuzJycq6YObCvdtlM3
cZuhSz07lxyUeAxb0n/VdeefwEuGldkdVGTCRjrME52PCjTlExlcIXV+v4QlPZiQ
Ba2sL+nfN1ft2N9sfw9mhvPk9lAUuC1i+sS5jXgopoQxJA0fOq9FTM5JBC5yUp+J
RrlCekZHiMkqizoomi2vRSfh5bwpnGmpThkJ/iuxHaoH7AbKRKPppgl9wXBh3yq6
WAMgReZDVy2bVUsY8FC9w0WmFKgg431b5YrbT1a3+ZTiFaeaW1cldmJ3trwUBd6e
DJffG14nwXA4nJ9augmDe6pZ+rhYYLloOk9xPOenoTs46MH5652Xgb9mXmaU0CNz
fozO7XdmCAqnjlm7BvectkHMhB+2U3XcIViyLf+psp1BAe2G11N2gq6GrtKbX0Te
HXmgQxSSB0DCyrLzxpXxbjuikF+YXzHss7O5TIpeS5shAFHV8HC+b6FP909+hvLu
LZIJVMNA+EcVqaPUzJjgguv6kGnv32pgN2kS31HI9S5zZwTxHgFJfXe38hniUhN8
9ebb83Ja7r5jxitPsnD0i7LyhPGZVCW0cSsF8Ztvv7/NpKuKC3CDFPEvYFwshC2D
pBtYF8NWj2QgVvzkpMriIU6VEpNyFHH/z6IV0/mlSfVflR3AZvBj+U/T1yyUfQK1
K7GMzISXROVQGJrvnAXMJWGrEyoEfE3nXcNkpqWctMtVaRJ9TZxAirjCfzaHrnNl
n5cXpXYO2N5ud2AYd4UlFq+tXg6iiI8pQFWmMDVoK6n2Wt1I061oCxl259AGq+sY
n3r55ff7wshTUiX/1i8VU0OsF5L1cgA28XuUSKCcq99miarKxfZWHswlu2Q5aTfp
74g6u/QNTgwZ6Z4FyGXOlBdVbfleIa5s0bzXH2SX2fdXObLVs1YkoqLC436Zq2n8
RgSJcoMbAvgzsjP6hfT7fpMk4XlT4cE+YANdwx/tklni1CZ3H3wdAQSJ0ft37F7i
DgrlE2WpRkWYWJQ/bAeTCksEJK3tDqZJJ3wmbgTaZl8w3azjUQx3LKDEiD9y0xLV
ucrN/jHcxI+NKdoQTIWtWvglRCO8NQ8bMBUhRbZjnT5pbxLmJ7I9m+5Z1+HPnBGD
tlK+d4dndtf5g4FZMEhSMZYz8QWA0J4Fm+is+nfekiS/gBrT+Y0puRhzZpRhAVHX
8m5MWCOQjiKxM49j6kwYw+o8VvhAeam+iLkkYuE1tCxjbDsO5QEM/9Shgzc/SM4Y
iXy8dT08GBQrvC2ITp4lVu/3rtIwXKajcUYr5U/9fAkxlWjTZgqTayG7g7PvodfO
6B9BBSlXtc4Aeu5GdyP9RXQ+6U9kx030wygqk6LBHxzfAOS+POxX3qxOPJGQeYyn
qnQEcNXII8xe4UmaFMMXpTpbDZgBm9p4N7GQnSK9AcWzAWenlABPIWqDWbx09rZP
o1CM7RSqA9h4dqAS7AbPCjteOL/6YMT3xqRCM7Az0IqjpoRgYsmAWL9erO8Hr22f
2lMLTiclMXWuIHG5ULae9c1QF4wGMhh/dNZS022IlQjXn1rXvDZyc00vpQlUyOem
aZExfPSTFynHeAJIVPJGP7eutnfXAw0FIlWG0vmUvV45wUUBnlLGrwwoEzCJ3VjP
IIrXVmMGr+olvXx5bkybzmTTVTA1ZXPFURYeImuvuKHfeCzd32kFts6p90V84gMk
B6cYw8Zl+ZtLA0d36Tq1zp1Sp5mjQavAHVvtb3lFRuedxlX/ZTzFnqqjeUyee9xT
o8d2z1TJhAnPEHLs+SS+Upo3Dh1gtm8+XVohb0bhA1Lc9wIIhlkvvHMDkXlP1feg
Y6bxzMk9OD2kOc19tXQS2JSpwoOCw/6lZlhpzPkoV/0DFs0KBJ2App8Xh9cUZQrc
4KYMkXvQzcQ7nBXRpE0rPSbNl22WIQcC9q8viOgrAumtPxKncMSgIR3JuMGQWpdi
R8F7jq67lHFruzONk/u+NpaZW9/pvUtX2VnI81WPm+f1gNYpnHqa4Eimm/h2QF0Q
WANfxjC82ezPXzX0csECkZma6mn8VJqBsycUHOzHad++Rco7yy01Khngx9oJwD6n
cgMF5BAHENPPPJnAH2T0imVOjGW3ItUpjYWo088u8hLwHetoStfswzujPH7idpwB
7YLyothazQEHud0JE/9+WFAMUPGUC7hMrTr9jDpb6U08DhifKX2Yhsxw6olWbmaz
IPLxcTTf28AvwjQYbJeIZpJVLzst0qdUuc4tpW6GTVnsbnnhhPk5icvmcjOYFYHx
Sqj8WXINzAfmswYN5WJR6xLaiwn8xKhnefO5YE6DL/S/5iTcCuru+cCBQiVWiDoa
sjsxFwi4F2VA/HBEOuH41jV49VVgXB+WEtYoRZN6QLIiaUdZH0z2gIu2mCvUXJ48
diHpjSEUD/tfoOsftiMpCuEgYRUbI+5Vwc5fdvSt1M5aurrI0mq37wH9DLLqL7h8
rPmBHXpyPazigWIYN6DaxXtLuBM9RswMAL3/C2KgZUW2vrMbk++Pc49ZOzSVa8zD
KPsXzSLI8V4XYrLeLBsbu/v+kF6tFJWUaC0sVA+SgKu1LwHMxNklwi5kEe0KCxu9
uvuU7r2rW9FAMnPE4bKAqezA8oLYVXgf0Hlz+9oE/filZkH4zToX+wopT4L2RQ3J
tctjRwiogt1hCncf+Q9L9txTqSDW33GcCWjn4uLCHc/w5Uv2/DiaUG3v6NenxxJg
qa1lMaaI/qsxU6/bGMf88TO81ega8da2vOMbhOCNjKgMYGQmedEDAZeQOy8MeUHq
5TzmuW88oKrZg8oqzz7HDWR9TkF4dS39j6rTVytIqi0OQlb/qdt5rcmBU0uaF10x
5MQhBMdMrh9MTz0qDg9yUXbDtUfI6uESvFhW88YnufEUK5E5Vr/fW5DInfDmTRnT
L18SuzPgz+yTl/NsqHySGhMK0YRGQQ5ivufl8yi1ApB7eRMnrowcoI7Vn470yxq5
RhyYfxFfmkPrLyQcjk+Ug/FLo4j+cUfNdyHohELfH1SgaDi7zSIYas8nojTGszWr
1ChKykh373fRteRzGXJnOYZEvz8u7jAfBkAchA35Ht117xCJkY8rXeYSNR3Hnjy8
ev2PzzMyn1V569v9O2PUpQ/UOYpOHXjvl3WTAlhM8WdrGlxWy2I6uWFyC3P3orQS
84+mntg/04MO6n4QRAyeNerpidNWOV1b/k5MVZVGca8yvTvZowC6XjXC/QAuBC3W
gekWLO0mlp502RFkTh9huN97rc26wOAw4qxVtUW1Nm2jcomAeOCbdYT9C6CxTBtA
xRjUpBFy2VgcjLw6usmvs0+4NSyivdfEBRaUjpu60HMTSr4Hd9jIJsXiNLUiB++H
jp0omZN8xOMkZTz8xBviPt+8p6lLwA/BXbKY/EEhu1iqVOxjqIXJI/IOh5OcG0de
9hLuMSrzarVmlLeY9bSTnFKZPuUV4U8tZyCkdfRVBWP5NMl0LUUeoaaAEqdUXKmg
VjVxujN664s9e03V0gFXXyy47FhTiDHseb3VGhRr4vgKbRQ9mEb4FF+AUQTQO603
64jClyXbOURZd//9oR7k95RglG8SIcLW285sVlcoCraLrYbsL3isAdJGm+8ruJfB
PLs+S47U1SjQNU9qSP5b7jn9gRJyIOTGp1KxuxaWEfviAywBkzlcndK/arxynKUG
3vbQhvvaRbsY1/O71E9Xj8gZA48pARyLUKvGnVT51whaXaHcSu0mGpiv1OaGa8gs
f71E8z7eE79zvubSpEsbsWyPIhlrITDkzp+kSn8papAFRHea86oNxDLJEmIxcN9r
pvxpCP7b2wFymLtUhXGy2n/h0MPoT9zCRMulnLIO95uYw3KYwGNCQRT/jj2qHzgj
yPduu5VXVNCxPYGMcUK/H/7ueBfd+IIycsbaDhMSH8bVxwqwfPYOl18+9QX5kFTt
n1j0fTnSdwTEZwWdSsFjeGOhUDZlE2AMS5KM+RAQjHdUUtuIcX8jf800Cf2a0L67
LiCNhBv+dVwW7a6hivCoiGq7g3jU07SwLbn9FU4qq289yS5R8xNl/alslmudVyHI
C+IWh9+ZGO0GbHaNB1+gb+zfUHnl8ZMSnBZ7cm8fas6fAS2L4nqLCvlu+mftIjIb
tLZ3YHsqC2qezhk5V4pVplIACUASD8jdlBCpbScYlPQwkUNmyppc544paauCEYcE
8suCbdi3DRkIdoe9/hFAA7syuJN4XDbibUtrR0jCrA8/WIilV05dtepf34m8R9et
cId0hc3qazqiHtsg5V9I3TzXPSfOoiq1oElaENR+YDlI4X4iSr8x4hQGeLsP1PCi
VWQqLU/qdGSRBx8SWv3BHGFTtD3MzwRdPWMV8N3LnprQ9M+VkHav9qmD9NeTaRG3
mlS3eyccp9O9V5lHOIfOPYm7BwQ0rsRiHzxekjJdva2VRA3Rw/fREeRYxueMnxg5
R3tayPcvbetfwbFCsJ8l2zj/2vBWQUCJ+96mgb+4gZX4vriGEAWrxhn0CeotUwW4
skLGgK7XYvRHsszbct8RdeyjNKadKQMbFkmLKgJAJFe9GmUSFnd9eWJF5BkcoJ4h
zwMgE4s2H4lMHfAPUODAQIT3GL/N7ZWghsmGQJ5FrceAhTndVPVzgIc3EPuyUzdB
7PjBgAmSEgklCB88xCLlv5bIITra0RG8uLTrYc03l919Et+P7+RK8/ZxrlQFnRQd
rnrzYrJL1VwoBn6gKIs85oXdaOl8Gf5TNRzgNsBVDp2cwQnxnrIq066aVqPvhU0E
3ikysisv2vUPt90CnV+QiqEnpZ2Ntv5mSBk7TpsZYriAQUm+LPO72GpK2QFhLL8+
eXTnLVK8Egq1SmZ2egvsl3tWDAfUYv9kwCt9v50JQPMpkMtXwdCRJCt0Mtyes3KH
FFsjPv/hGVWG+0drT9D9ouj9A8umUw349tTaC/m/XXCBXA9Cu64e1wX2suinTMTX
IFM/MYFUeUGhaA2c0yAokALQlkGTWrV7STGcEPAuygaC4v+Z5p96xziY45W84ovz
fISUh+OF0myNf8/5+MQdp3pO8AcN4I+oTrhBCw0DdebMGDtf5lzrYBlih9/+6vYs
h+35K73HfENW1ZUP90JdLgw3bsu8bIqG2Eh2jE4ZvCNaZYWrkqu3VmRD4ib32YTZ
tyE+4wrFQocbIgoJ5+ZOQmTwZc/RlOZ3ooCXEfReV/kzw67s67uOCHcMZyBVUfQp
LSeAngyxfeZhUy3rD6qP6TVigLt0jJJrkn6wUxlMNKqnANQrUVbDq4t1cwjH4JJX
WC0D/eIME6gjiq17F33Eo9R6T2khLiy0STLzCr9vPAQ3JPtYTPProX+wHcM2nd3U
LHclTqarb+U/pnIXPwG513HMcOu5dhTL0FRwzdNL52B8LAv8nnQ42YsAzwwrnSIN
U8nrdJPqZTiHciOinFLuL8+MT6QbAABHXLoal+QO8vCyu67f34yGsMgHEhubY5uD
BSWz6ti4YLg3sruGJ/cdbrB2rrOCpoqNT2UjuVXofYij/EaOO2qdR9hme/X9uiaJ
kkgGvlHpqQmRUpyamBsdNOvFdmT0UpvJVKaDxnrLe2pME9f7HoRrRvfCexx2nLYj
Yhs7gtY/YU772V9cPcpgcm9i8jCMXl2BgG5rtm7i2W1xqCK2684vUD+iOTVs6qWd
Qpc9TAFdUYUH2b6tvJjavFYlpRfL3cdXxMj4WBUbe9ArooxpifCoFO7Mo/PuuxDs
K8qVQObBWgeTMj09lTclEwWQhB5p/FotZFJuMxhNGwxflYAdtyYC5XRk8pgKvOnq
HeVZNFLd4fN0b4TZsw0ze35HnlvTuXj1oc2nMTBJTo2PD1r7//siUGM2j6Wb4dc9
Z/LKBUcBaFiSAtyQCI5KmBnAw4qW7lPNYbe8YCP3fZc6VC2H+YZenVk+cPO4lt1m
+KYmzMigq5xuKjCPg7exFz3XNAOI/YCrleHQTY6t0Rvxm5XRDiUYwKUAH9ZtI6yd
Yb66136BEL2wIMs0jaH6tXjfi/TulN1wCwVo6LQbzb4okTnjxTdAUDU19qgcpHuf
S1CFcS2/iCrcfSu1jfLrDkQJXE3QgE0/CudEcahl6UUXlZopHIY6wL2Kb+eekZ1h
l5skFB/HBxIqVFEegH/tUISnk819zv/A2cmvTflMAKNBRvjYKIgNIR+hlgxuGJaQ
nUsDiDlzR6Ep4oJG60kkIsHYioeRIgnYYb1Krd9Dftur1SdAQHw8ZrDTPAjhbsxU
jZnocmvTtZAWrAL/FzceSjloi/rVVcxVzm/osxPC3edvCtSCrNqE3+KNGRE6QdcI
qf4NyJOIwJ7uO2WtSWJSDZMH3kv0FwZX8YaKV75j8h1MD0AlL3AJdnF+6I7sPjH2
92kWgiC5zGldpONVs2pOzaGoQDXFpLsk68TnjM0zt1pEAeXrw+/wjJ8ycdxLqiyt
Ep2GX/QU3hlgqLg5NsiGgqWV32hqjClpskn//QYP5TjrpSVP9OK8NxXjbaoT2wld
55ePiu4jI5Gb14d7vdBJzLBP7NpHdmFzA0f83YdPAGSFYxa6YIDSQulnx4QswZN7
POwhoHm6qC2kS3koFW8F90JOtztZsgIhvoB0VuKXebbREkO6nSMEHSndhXemwcnS
XbgocqDk+lmgn3FpAiJQAHhEO5/Zjj6aQby1mJqj0k7KOlOlL8R0oDeFSH88iYGN
o42Rpn1d9TzoNp5CSjQwKw1Ssy/iKhvoXD0BijJKZo2I32KEke4oeLliu+PIJyqh
oDCYBsqlxM77CJpF4Fuc4P/1Jjk/e5rBkd49iHGDFvCAAppoMIgxlcuLsINkcIkH
b6Vb2jKVEMO+xvl4r1v7W3rM5PFxGGanrc1f0Ao0PALPDIBsnhiOdG4sC6KcZq2E
UpuXEE0zmG76oAtQiIEhgSNmjGc25ct7FzkCG3fMaYsxfN87yJSOJ6mi8nUWAmRl
k8VPc0lkTVd1qt0otjD4FkTi3l1ZDpdcjpJHkwuNQWEE3NbnQQnhSrForHEpkp5c
a2IEMiFX8zPnlYQzK/C1QGK1lOkkujaXLCqH8UDWSuBkkPWAPDjnLEJMXT3IA6QS
Rb05hYrZdEMgzY9D+IT7rKbMh+LTURyv0oPViDBEVibgJzT4Pm9NomTl7qxdipSD
edC/J5njCTXZdDAM/A9WEQhEJuzcZZGMxqkyN8WDU1hp5LE4X1SrhRu+YFM/OeMR
76v6F1AfQ4G4DQzrtb9cYffQJU0CehVXnF/qQw9GezEbmTB25P9smW+pEFh8LCN4
osq0fEPM/umD5AakutuvgD3zTai8ddHnkhYCGsdXi67ISCGD01a8ev8G7w4mBeMh
FxPnNw2ba/Iw5eNOJFE7xMKCxCLuhL3DwOGAtAvyj6zLzxCe35vmzVTT3Te+bvhD
MYlej31gaC+MAZvhFH9X+i9+XwK5U9jsFzSxtJZNnTTNFFfGU0sYCR29/rxsqWLx
QrWeuxx50NdiKxRFk5T8BmK1N/oKq/jOwz3G+Ln7WhaUjL8LuSuvBiA48TMKRTgZ
6KnZTi9G7+LmBA/lH6CZvgi3HgIsuXY3DuPz1aP7dZZOx+cQpw76SNanDDi+Q7Gx
ai0KcIvucKD1RPFm4MWtb22AixpWjA39P2qvKtQVwFAyDxMUsKCuWfCKCP9kqY2k
vieV6PSWdo2LkQOjlrLUJ2ZpkOwJHQLuhuB/NI4r9IX5067G4fX1wwqgTmFs9DCz
KV+8p/VLiPkKN5C/y8eyUN1fGSq5y+qdQMw+xyG0Dv7tZN2bpHaQ7tnEunVLc2jZ
5/7HuGb+1wq3eyWQlirclhlQt7rnK8HRXQkzqTujh1B5dfVu0+RAPOm+QupIfvhV
30elGuVKW7Q8sBmp3dY/rqin0DWF9G+ASJGhp+IBA5kB8FdbGMuvu5YKmolFUWX0
7Rtzbjg5wRwd+otsw3M+T5tneGueh4lBHdJlikoF9NXz/nNBLB+FSrZR8R80Ef84
uAIiosEYXsgPycIqUPD7XBASnpPej2FYXE6BqvvBZXvdm8+/yfk34HhzdezOI5g0
WXPd2Rw5gf0FlMM5RJnPE05m/FVbHwSaZg7Qn0DqUtjZc1YhnVChFf3H/4lzGJmE
8QL4hpdaNHSai4JaVDIpKOZilNYpKT6Eq1chDlrE+FTLxGQRnGNcbkU0vWhvnl3O
Gy3nJ/eWDDDkGogF0e1mnI3TWdJSAJ//J7P4sK5hgkNPrOrVGYPmiZHW1CnrrqXt
WjbMMUye8FIZnqNSSggfwOXjtQqsWj6dXmzDP2rZZ9N0ceerHqVgVF8jRft0q6gC
oRhSd5icsNqE/lnYXAmGIpEhjtaXdgz6qbz7u4cUOvnU24X6K6EpS1rcrhpwhlJh
bX5+jWwLWaU3JowEiNk9xa2b+5jb+WWVFdmHqW7W7ql9Vr1NRbf3RxPBHc0kEnWe
sutQwi/GeOca/8OWcZM5ILz+/IqJqgnLEU5TGcqghFUFNQEc8l2sw1EPigQllv9k
ezyqoO+HxBx8w4zmoFZ8kenCqp3q7acjc3aYMxhanVC1MvDVvcJiOk2AQug5JhyK
J7oo56Sm6FcBtX1bnVy7oi5ZQnPKBiJZ66pc1OmUstHpa0iyK3J0Ze81zUJjjiic
wo8mnwa3yisVTEW04wcpIUXgEFXE9KS5xuHcRiUS4mw8kGG5AkhISpOCSDVWsmhm
bcs97wKMMTUiIXt6HH6bS0ASUT/s6yySmreAyCAz+dL14B/km+L+jzoumUbkKt82
QY3VvQGVXoNowjjcmpWFndw5TCep4svhHmuchbd1xxSJhjRmaYYZ8YPUKCEaHJcu
AQPXtFvLKO7dZf5qrLkQ5SKufu6r0/uiucJbwDdFy5b4nJaMaSbO1om/iusVzdPW
wni+NNeDgdW9JlsJFhijVg6DBgJyP0qISD6wX/22y+/bqeETI7gZTgJdnvN1jIS4
6o177grdu7KPtMLP27NJQKIhwdpJeEaBq8WUB7RlOU31T0ZfCYeIR96j1jUhgffw
+rFh5qFTIHravv7rw+ecSW1BzyRj3CqmqqXWrTa6BpWQxDzJQDvjV1CjxYWJLdbo
50ZEByyTutwF11XV7HEXgKK+f9xhsDqZpOfuhKWRWqByf8PQOr2G5VzX0sfhxc86
ESR6iMVVXDte3TdRhXJKuHBtfU3bGw8NSUme7BTTtyTaTnt0KXH68fBVK1yckwf0
x4j899KWSBYiY2s1orb3wFai0RnyOLRQUT4oLKF0fXl9L5FYf5Zf2h8s1ntsGFan
Z6sDEIBAiEtPXDxR148DuCTcBAqLXbTvLDivmj95R4uq84bZHJj3XqDI9sK8rFXg
zqIQLWpBW2wJoo3//gPQp1YXsICfaCHWoRk1IFT/sYhEnSAbCyTfUusS7SlczqKC
qR3KmxKUZIb4N3FImoPR1vGaN/7xVIzPW3o1RzCEF6wwKHVd6eQR1ybqEJ6zUw4o
T3eUBbxFSUZd+MkIntWZsBDYhozCAuQpL1ufkv6Aw0EmTnXQNbcctow+ddPlck9z
T7zB+cFOkVyG4ld3WyO7eG6Ptt9IpcFy4/BMZzYZ/FDRXRiq1K3evuHrCqyb9YEn
q+mONaWV1eqdbeIyIKfbH3FmaFZTMwYnvHBMVd9RFUxtgKEypPEIX7Loib2A9VtP
ULX3cbV089/yhjKrpuNICTUJTCo2eoqfRSuPRxtLRJms+ryA8+ASy/OP1QO/6EzT
ojL0gNQxwwgNeDvzhWPA6XJ67MQ7qasK6PyhHkNt3tTPgyo0nf62rQgjUfeiZLiM
DpYyVVbfkS0l2OXrq5k5bWkUx8oxljoPuI8wQDkAQOwvRUkAtFfWvP1XKOYVG6My
r+QgbQb1FEdFQeOfzyXmEm7EmnobE8UyO2cT0T8WxOQ3huQs8t/RnrnUU37QDiJN
xmfMnQD0v0qVvrhgtzT3+P7RzFJt1Gv2gORjiqczMYUzsC2rThYZZ0Ua+m5zxhyb
HJ4hdpxsuiRbsedTyDZNvn7j8da5nDxVc25bvTOm+de5bxmC35HwmyAvhXCmG61b
qrU27oAycwjD1yNY3wmRXOeAfAOW9aN7OowL6yUxuuiKonWi0lUUz1rY5HB5H8hX
Ke7bTU8k80ekrHmyH3wkJKAYoAavzf8CQbLVhSwjjPA1qx7PAnGXXsVpdJfHhv+3
eDSWnTVB7LoNXdzgzgZDphjyXiImBkRT+ZJ3WwImTvpu3XzAJrM9RHq875eluCMX
X91e5S2nlPw5+70wRxPbs6F2sLGfShj+zfMwK5n5+rhnYIVlcIgSsnS4VlAdPHF/
UX1esLdk9CWo6iPz3pV/XSc6vuPFJDVFwK/LwKLumLcJ+n1y2nxVtTXxcbNUz8CC
yZd/ECcCe5R6UySFEgo5/cwRlfk7OP2CQLfyKbpr6WMlDYcuvgx+XN71plxxamF0
xU1ausj0HnaHmPSieJlbEJWMwYeLiAq0ek6KAIHMCZuc9r0jO5GLpFfMM4HEd6HU
wKxfsrKwVWpzRSYHrfvucDoyA7YYAoZZJSj4eIDwyHvD81MfSFVo5RpXjyqemSyo
REKyZoIR30SIhmgcyyxix9CC/KM3fDGky3atWVO/aVuQv56XoErJnJgBGsxFp5QY
erEzn+0c+4T4T9UufmYbbk/SX/mf2lAJsJGuLkcpP/mz+8wqEMbMXOgH9zmhsHbz
lwWZPVpgqZyUeAjvGl9eP/1zrN+O6SHYgdIz2bN9vqTxQl0/KsVZz+wMYMBUjluu
Czw6NTLQlWd3nWqMCYttaHV8tvPrvewz1wEJr3l+NppaQXu85ezITMN1ZVS2IMXw
rz14cUdI/01G6D9JdzjDTJp3h0HrqasHOHjOl5V5yxqUMXxmyjflv13r/QD8yfXZ
q4HvEk/pT6n2H9P1b1acuKUD7Jt6cYTxxCVqycLZXqrZfobxzqKlskOkK8rISkJj
wDz4Q1QGiIrt5UwKslcgRhq9M3EH6O7Jw3bTlq3LpIIYmkMBFVEUiEd9TQGWOxxh
dUZM3wC9AS4nZUkXhFKMs5TSblxUwvF8amIhbE6M3EQnKncdQlhqpJ+ZTdVU0InO
BNVSVc4E6ouaOXpbFOPL0zf3R/PpECmPPyst0O4okJtxvQzJ62dAUa4YMbAIR68F
xsX4Bj/FNi5HGJXTJXg/AbBFB53DC/+iASvivcBVsWJVwLusGoP3UMaCptly1zrW
GLtCSkr3r+o4s5PCY0MIieVAYxnNV1mUeJRUTvq9yZO93ZOdEb3Tq5gzgcLv/tEv
XY/8vtSyjQQYpkSsQG1sLAP0kUWH8VSoEOwosJ+pUT5f2sASmmK1k7QZ8n11m2/O
fCWXzEGPAhtTuREruaRtGRGI27Ou8tTmLmmVZdJ57PxEA1Zy0LrXSWtuTsO8KChf
WTIZxxDNdYYKUBhSib+fy8z6LAHphFj/LMEcubpVCf4gBOqST9mDZ8GzC1yLEVTz
9DfpeMvFnEuCQ8zTQkmLTzRzZM7lJ9EAxkHuvwbkIh1G7WkRzbjt1nBB2xovSJGM
afW0seVltCTsy6mj6XP8PX5s62eKdd7A1uYJ4/JgA/5V2dum0bvt0eDEqguZGIH2
bpQqA+HK/E3zq64g2GWJJy+bgmbjVOvo0Xa3slM8MfVJz48ppG+3tb/AJYlBiNwV
oozf3XaHSem3l5f6uzOV7uKj2Kh28fZ2gZqqVRgbNMzoG25WBaf8ijdxvqBwcHdH
rXLdI2NszHPNfQsMJG7yFZ96Q/hayV1E15h3ydgoFVNDibRip83b+gTnlWPCeeaF
pOcwj3ShekWPGIioE2wqcDxhCf/vvdxmSxvv0KO5ZccvEtEbEz2VQhC8kAsRHl4C
u3NcLzih+0Nxu9sUabMG3192x9ugC7RwGZOp3t58oQSFj9qAuB2elDbdw3RenYI4
UNCn/+6evTYEFbfMiIApKbkpLccTwyvbeRV/ZbBnpPJYnqa70wtsoylhopJujGSd
6sVmwqr8Iei93p9Z2pPy0Ph9IMXBSGuesERVvgz7TDB0CGHonOlWhRmjklsMK8j+
ah0ZwRUOqrC57zuvLmMSmqYefyXCrI2txQJDj6HywBd+vMRsYnULnjVxUOrkRUy9
oAx/4mMIAJUHmM6TyzOk55z5s27WDEsz/g5gmXF/X2KHXaDcqYunz4AylunT3m3m
pmj5gUIfRn5lTK1eenwwXOoJhI9RVdOqgNfZzureuB5gx/AbGVsLu9IYN2mBFx2m
Qg9qFZqVhdzSQCweUq2Ou66eERZoiHi/pf0AtNL1RylLZrrpHVvS5q581A3lPtg+
8jqyMtLiLqlxo6TXBGxagK4etGXNgN+6VWXHlduvXkiL+vUI4iojyX3+5vd19nIW
IT+l9vgDO3sMLZ/ugTmUdRLy8nfTGMmrdOwgbFTowBcnmHKxRl8F37ir5pkDmpjG
LpyYn3nUWAc/l1NNvENQ4uW6QmPLbbgbPSXmhDAMy05yjwD0tqZkVoJqGoTGgjmF
/8O9zrSc3UrskuaSXRgJxojqRPQb63MEpbbALWhyqUl3GhSzr7ivud+JPg1YP4lb
wPut/RxxgY9eoPYmE8pq3u4hCD2P+7isCJxGe85KXus48WzK2gdszxG3HGD1pCTC
2n96GvElMexFk30UdRPciY39zibOLwfql5OCWIPpp5t/I5GZeCQZYpM5VGn//VN+
F1P6ejKtmUWnuxWVz+7OZdXBz/ZlhBdSy2PTOu1DCJuQazcWvifM6a09ZBwFE7R1
yGiVIUxHKtud7XuB41ALae9HebKujAVDIGqmW53r3obn+9OiewOA/e77JRZQz7aS
/yH9Zwy+WgeeCx+edc05giLMRZ5E2TZTdKOR1/KYDp8pBYcGgmOFFsMI4qcHBedG
l9+m3qGdtAp4KzJchYknAhbUiZV3+tN+v+Mop3gjPLbyShPhm77m3zUfJKp9WB6F
C51fLnJlAqxkVk2ZquOKeIU2Dsqgj/mAOVhDvA4MXGpZKn+ygPk9OP9P0ZuGT9sn
XjYcBlPXJlSh1TSgwu64VuRY+8glsX7jpWyMFtz7XThpyOAUWLB58BL3yJZimxhX
l6Cndhb7zPDegbKHYBJEJbygPHP9Ep02Y/GFGzBx5uW/IRmWNu06RapuIQk9RN7W
CW4Jl45wgBCrB6yA1/bEFUcpSXvo6KG1u2MIbKz+Q4OEno6t7gSUmtdEpahAEj0H
R0wSoChCSGmdEJWlauARGEN6aIwGk2KvhblMNfiOvwFAvQMb+bZR+o9z5ITXDWFo
rouRj59h6Kj2ZxvCNdF1gxFUYT0Orfvt0nLGp6HaKhF08i0vq97J/Hf7o+jXn3ql
XXHSFrepBs8Zz6/UEHX9JSJIbezUI1FQgDdvjBL/dbpI4P/Sal9dmWoB6Vngxt0Y
FFbfzh3e/1L/a61puLZdd2Tj/p1vsVpF5PYF4Fn+mgBB4khzUeR/AtyQvdIJZ+WM
tsck7fpOWFnScvIJTLJaJaonBb6zeYko62iAkCIBQm1SsLUgYwQdFV6wm8O6dLE9
zbmTVMwDY6Vky4E3A9zbtExxyRP0KPrKoo5MqR5fvjbNqE+ZVNaedgg5/vbur0Lu
90ZeeFUjqFfc4CA/Yx5MUThzq62GkyGik2I4elD0uh8Oss+1viIWz+6s1ianh0gv
6qZ2puya9Z+woJSKwBxb/FIa8JTKHM/qG8XjCuwRHvFHyxTsNYc4wmEaU6LfYDqr
9S6gZJiXzgf7oT+wZg1U0PNFPzZImIuyDnS94+CdVIKyj0PDqbzJqxKLg2BqVq/I
RsR39RQp9P9kmpd+u/liWnBNmw+uQd5Wfq1eiRj1VbwwARu6+uf5mpgyhZ87vbmg
zpixfdwCqbIWuvhtBVjE2+NhZ9/2xLpVEgvfGCIUnzrPK6pJd1/yx4+KqKkMmIzm
Dp9fYSC3SZoVEpdEdp/TStfy25xbEdN3J0y/kkQVuYYQxr3j5YqNMbUZOfZgDRvo
3wbXFBsuDPs7j9+Ced2lkh+m1Yjfsu1DzMwGfd1U0xcrXgi+/DBjgPc9Rx8GO/es
l7nxRd7GeFGARZdm5RYmzlddCeu0NBpoWi5HdDZuC9idt+mqP6xYoMJS8qWysvF+
oZnGGbkiRROiW+G7J94fdCwUnrkRczBlyGAwFxwKiDnyhDF1SsJ7V+TzmP4KbE6W
jl3D5AdV4Qo63oujyhC+74mraeQRXq0fomzrSROn3GewJyY6nuVyCHzcF6hlXDn0
R/nELr4yivJ0tZXhubs/TRTB9LJOyj19rHtC1AnKBFffCZV1ZyedU03NjgNQTkdJ
b/T22xrE5lRFwTCXZBbpjZ5FJG9bnRi9+Xa8teopHn1Y+66z9lMzedgfb75/zN6O
RMJHQzOTThousRIgCcojE5//Um58yBv5Fp6rW/n/Zs1qQtY6P3avjP22HcKWNKFq
wpRTnld4Y9Tx4ZURabxsg8n9PXLh4KbzZFm/vlRlQhfdSVVWPHPI95mcEX0bbKdS
rYl+hbyUE6yk4eEuh0KpDeuYpcwOi8UwQDSLLMAayC4xnfFvRo8MQmsUJMwKjSVh
d5TIpFyJjt0OcxjF+EANQrL+HGR5OnJ1s5CUjf6YLqa0HkmW5CIo/Zen2EC0cGtW
/eaPVqDkgVozTlJhYufWJkKds7+vDIJ3BerDhd/K/yyG7/aRnwf8ak5YLFNVgoOV
+5w1pi72ajmQFzDckWdRgPL58eHeaJhbmDQwdV1tuJRlMbFeW1dwIDPk3zDmxQNg
raNvl688YS7Xc4MO8J1x+pC7ua+gMdUmraYheMgsv1R6d9+ZpRLrrOeQuUTFJScL
JBpdWKhdXTTfLnmarGfPwcbrnrcV5jT5zeqjNMm+LV2xPdRqTPPeQyYEn8YjU9IS
7t5Bh0NithHsDdexpJYP8ReecleP1z/1mNJYGC5K5h6oIWNy93hDkKxsQaNrVL0+
RftOn927mG7LY1nPay9w0i0Ns8U6fnQFdiNeznBHmaDyVfJtGh3VDgcVdMYH+gTu
Arf+4/urfZbX5sUrczaj5CymJTmSraBs8TND2+HRIdb46yN2Fsq0UMsC5FrLPzTF
Wn4dTzmlL9VDLhKQpWsGuUeQusPGh/YK7FKaHECKEHLIPVd7KQgDM56JVLiSjmS/
cej8fIioxUtUJQtOTmmtvrsM8dH9GV/heI87fIOMVnwG71Ny7bFy8TiPQX/4jIXC
iMZCn3kvp/2+esxJOXvjCFwFMgynx+i/e0hUfGPo07+LXyG74CNGrZdp9uAOdGQK
YuqVFA8ITljOKoneJZmHZo5u2yD/RmgmjU2Tf2/AxkOQOxai+4Oi+YplX8QvldoE
C1FW91gs75m295koS1puhyTqS5OvyFz+w+2qhYg9c7f3aYDsqpsqsIBgzBTGWw35
thB12NSNA7lHsQbJLqNEEm4fekxQ1NPRBMsuV2SpXdhw/JqZ0FJ97QcfaWPEusgK
KSkEl2iSg+Lax+dcZs0FV5KWGrQeARs/RKY3zuVLvjKWXBx4BV927fKVCuzdQ3wW
nfZ7UBIKolb9Xd09jBYBQCO2wOvPzzb5Tu9is1jYqatWoLqTCW/U/Sw4eJm0uWCd
wuPmzJ9NtaiDH8TYRir+3p5F+bpST22vX986SdPenFUT9ezyqStd7oCGxMdLlkCj
i6ZokKp9BTpxc02FDCBQGctR3WOwawGm3AATycU5L3dsbBtwi8wRVbX5BJmmzjeA
SgmLcDZUqx9vf5rrtVwq3ZJXtOOykDCNEElh8PsD++9J+D8LSmm+14tWdrtrFEms
aGbbRv/TuXwFML504XvqSweLBy/fM0iBxb9iNzEfGtt4eJBMDrlYqH02Lncsq8dr
+BX3/Vjxcszs6PhcmQrFye78ash1VpyktbZSm5UuOViG70Hne4zkGvcSE8YMXfyd
tR0j1PzaqBbucgpPpQhuhfkQxkRr+UyxED5mWqdogJQikQpt0AsasuEasZ9+dlI2
q35dP1N7sJJRjsN/rShDrCOg2tXMEwV2bRD7A/Ka2QwtlDwkff0BkHx684CWKKE+
phZBvMLtVCnjBoOAFDzj8xuMcfwul/W6jH7BFLBdMGUZXA1Nld808Ky1QZF9NHKE
ghIJJ9GpUlHbIw+Z27HhwLA1qIHQIGPn80ZyMdJ4ZGwvlQIMZwueZi5kY7Gfva/H
f9mCRH3sMr+T3gU8rsKOynQ5w0D4ELinmNNtWzw/pCzz4mYwjJVed/czJ1oIqHrC
Aqjnu6NJjPbfwPFN5xsk/NsMTCiCLcSj/u3oQHDEsvp2g9UMfBTcVuZSkvrVn+X6
XtQasYTzCicyQAIAR+GtduhHOusy+LmTY9Q/aWHtfUNaA7Fv82g/5gx40XzpFaGf
6LhiGUP3CXC9j8LVec3iyhWLr2XP48VFVDQ2/vG9uQ0w8TG2gf1JnivhYIpAXO+V
SGUYqNznokrDlXHZvF43U8yyCqzogo3EsNs+8X2MrHw6dwcvL9XIdJyR0hA7dtPy
DjscMiSvGpVyRh55ELYEiaTiYuDJxxp2Qv/89UK5jmk7PJ2NDoUzQzzfH9k/d/LY
lHzKhqwDH4QOZDDDF5cjpgxQfRTfreU42WBg4ZwFlR28/HpT+7iHh/uGhXz7GG7M
49yRwiwXroGjhrhBsRmPmVDvwY7gCDzwWP7ncnf6Xawlf6czSpq1a1wBBxTrbSzA
b8zLjTLsevEARGD9PlWN0fIjZj0Q9iOV1ZVSwM1sOZ0RCGhVUYu5IuT9FzGT3gQ2
ArgPnB6/QBXqR4Ojiib9pvo9QQC9fpgBDqa9EFhOy9a2Dsb47qILqAGN2lr2+W5g
BF27sdGTuFMgb2BD3HPUxyYzb/XCintDKgOHlv8hyZmgBfEJOivZrZj/vkWeaKKb
tqMovQy/pB/+3cOaasiCTzUsmigCEdX+pzxE0LbdY/rJxunjX7ysNdtS7Yb96sH8
1Bd6OuogoARWCSPjkhS27317POFoNPdVl6CJojc1PaYSa3uqzG2B1MiMNmJd8xm7
Q1flTAjU0fqU28i1Eyb7ypRx+xsCEdBmzhUhHzvWkfOfE6BejjxmqwijoNl7haWA
CtsTPDxMeq1z5pvQLc92OMmAbrCz5mffbUtSvRvTdfUwsG/ZxxG7Ps2ASEL1IQ6l
N+zCbW9Fn2zy9bdLGF6yhqrKLxZOXHEz6C7DqLutMuIR+TQmtgjZ+qoOfwzxceKE
205tGidDQu1cKvRymaZeRnsk1cY164/cCSsu1IDVTl1bIHlQnVGUlSzo22gukUqK
cf6yAz1g+rPP5P4VHfSFSQEIAnfmTIsVx6NzlxinHmK6lKF213KG7cK8m+MjQULi
SpOU/PLZ+Ugeo7onoAodwK/tB+zj8ZZmez88WHrk7cmWwi6JhxeMa3JdDPkhB6sx
CckVow6QWaHYFVlRrT1EJXLnb+w9sp7/or28z58VFlyp+Wg1HfOyHFUgmDma7MNv
Yk5hJIBPatbRB0plRrhojdrrq9d5RjyCOK6o1nQFDj2pIQzqDHM6BMTZ/85gPOyf
6OknDXB3hJR9a7XkUfVw7YSLYyAgGZO89P4ToUiro5xbGgfza1npEWs20FdSPChi
9u2IIDKiE8w3MXIAU/5pg3Us1exsaM+C9v2VZlVaAZlH8KduPgs1wOmaZPS+ytyX
538unNkc/6aAyPA37GPYsYhB3KLUGPRLp3ow3lGbsTWXw7QwVB9+QvnKlB35zElE
njseSy/YGgpN62fF8Vp41cze0V7vpXmvkqS0cxmv83BALswWyhsOEjNryYKbEln8
3SZ0ok/WXdVuKfPfN+ZKNCkjCjQRNTpdCcTdGX3In60QANTX1hPKuhlpqSCE+jNT
P1WSJP+/PfEPja3JZAI3/eYfNJwh3jKr0XGMBddtX2NhvifbQF5vm5uCbg616vem
dFbxwuVZgfa3m7iVIEmonLVmg3A1uojJxQiwNd/uYnNQJxMIqKMFNIj7dfy5TtVl
kEyFEIQgEAHnLS7UR/+t0fabL3Z58fb5z/ybf8sPkRLSYeA4G6JY6Or5zM+r+HG4
/bYStwc7nTj6ouD4bJQqX6iNg5xgjYXByBE/P6H088YrYFycV7azA7QA8mkvG1TK
Jb2f2QIFgVHetzVaFsQyisGQjjbzRb7duixa0serlkbqpsUNC6RTMtpFQZVpokG/
cC3eH08RhJiAidasXTcbu7N2DqHnLFLPPsAgE7WfoR+2KZfustX9+ih1WcA0TIeT
lv8osR1fucA8yuuVVCkF3jSucUDs8BTb1gnsDcb84adCGP9sEhEggYFlyfyaI944
fBYq2lx2AR+eivyxyU+IE5B9guKP0wSSKjyzqn+oVytax9vZo9daY4afdxyovKjL
36LM9K8EofSY52A81vbeOcosIL3BaxvwgDEahv7D1OlZwddGnXeJgH/YyAD4N85J
hl9ABH0g10duAIA8F+oWO1300WclY9Bb+owzVG0ZeA79L9uRAxrLNSJC6fpbtVmP
ONF+KPamwX9k5aYLCRbzKFbcJPCmgb5HBdqZcp59kY/khVD75R2hPhKleXy0qq3E
aWP72qLgSorZqS4u2VRRkrEig/pHojv9xPdjSK+zesBD/3LAiW+H6t8xazIWyfEz
ZVVoekGC6ahruehH9GCrFLX1BvQPrp1H6WY1Z05wTHxVMrPJfXeEd4W+3qlbXlj2
XZ4cU5L7W+h2JSzt0HmShqPaOiI1Z6sARNupUvkauZdLSYgUyTXxGpeV4RPxA6v8
oI1pqh0gN07lITr/2mMsCManL4dXQDSjOo5L2gBrQ4axIK3Oyd5s8//mCG7FOdWD
ZA7MqVfMzdk998HyGEGjWHci5IaOydDDRahi/BboLjlIY3QgoBjZlGkkWjqS3S5o
017K/t4gCCSsrsVZCb3elNssKQc0rBlJ9SnxZz9N2FPvlAeTkMjo0iYt6CpJieG/
NLxGmrxdDhJDD6GK465FtT47uSI/Scm341nLVwMfiHEQ9fMkLCLwNwFUtcilliWV
h1rlL9r9YnECD/k3rvB+9wQQqoT/drk9Y/iUnrIk64ZSudKlkXA+mdsrSDk4mtsA
ZXEyLjhotVv4a30EOSmDKXUp8n2VIztPh4fI6EL4zQ8TgJEX9eet14XMVe0Sj2pP
VXxVE0SPtvOg14buw+Qg3FQs/xq5U1NmsFyuQ26e5cOUxEQgCwKv3NDZdvqouKpp
QxZpW6vCViXxQZuZHqDyPyWMRBR4HxgX5zENBNVvmf8EYXSEwemLmW/txWFe1GZq
BoXemwJ0wfWicrJrfnmcBnEWkDRgUEFXHfjh6MsMdowuTBd9SrPIJLxjfPES4zQF
dHpeuKZY4eAMdjeeiavMZ1RQoT2jt2JM4XLo0tazTsqA8PdliyiLlJPIWGFVOBS7
NwVX10phCWf0d94JohJlazLeVE/4Fhgwr4NM62mVqba+HbC0e2VfhvzrwulbCzRM
87Xp+WLa/2awZZaWbRjCC4phlx1udQOx0CQhvtQc8HKSozmch3Fsa+WQjY3ZwDy0
Z2DiVcHXUC1SisV2b09AgpDq5jH0bWyVWhCB2cfbsyi5tb8cIVEeWygGCvJBTQwv
zNJmYQv1vLyHaBeRB3DKi2dcDwgrxeLNga2H8g6qZ8caowxvN/nRekVJHzFIgZGH
rqTyQNKSxgru7JEQAxt8p6aZZjsys/qQ1+ebp4RYI9QTtWdQ4Z8Zg9atyM/OHP99
KC1vrYVCwsee5AfgMYkwfWhC9QVN03DwAv1QjJCkRq8HmbAJrWj6q8EaSbjNr6Ql
OSGWrw2jj8N1wmUx9gqRuukBmIFaykzdjF+/6QtUvV2GKToaz7BRBYZNI4QDNZVT
TlCEXcdoD2fekjqnQ9XWuhwK4wfXn+l89YybCV6d8g0QJe9FvLC1buSbaihawnWO
bvmSpn0kElnl6lOpplgsPWKbFTSkd4+9t7WfJzmStFc5CTVgZ8gYLHXmI6GVMcj6
/QHU3E04TrkM9ud7c21bte+pfL97e8dI28MqDX/Ou42qE2kZKQBKYtIxpvO5o/nr
PEL/dA4ZdYO7eyCH9ISQb/PX3C6XKid9GK0aYkHHs0vE/dLHYg3EeI8oewDffGiC
ZMuW3bUL8mudV3AokHkULa9wTDz5RVqkrnLws0ulD739t1FasPJ3VqTYGfrfHcnU
/hdxyGPeK8FN5jv7HZRi/6RRlPE4N6AaCKcswB6SBGwVrlX6T+v+UN+Gf+l0fi89
wRvt3F3273R2JgxwZj3ZjgLF2WIMowbYrlbqBwDCMfsy6KV1lo+72Z/UcDWMNCbf
fFFM6ISg6wY0vhyoyflktFY4AV6cHcifqzcsobqHlyKoXkGg1OEQQQZNN8jUHE/P
6ZClXeSCTopIpmfAp4wLu1FWV20pmwb3X6eIatUnnZctl4knIIWcSEIvTxOIRZl8
N8GcIyyS2Y9IINOUvSm/kMPcbHDD4AECujQyqubZu8pIgy59s4z/LwFCIYp+c5FW
mv15ja2lVvMvGqrN57trqY0VrZGxyYoyD1aGMTWJyOOYl0wjgYSXenIDS0nom5mu
NA8ZEIbduWQPYkWul+37ldhyhPdKNfIQ5oYEZN/h/mUuGDEfvPzLzjhWIzo5XWQd
4hythrU2pVL4m66L+bDdF4Uo/ypQPpODrT3MBXuTutACgjtS+IKKxYQd5Twh0Ewj
ZK9Jzq8JGhG3FRg0L/oXpDs5tA8WmyBq8rqAo5IvK34zjatL6tH0RYD8rKNCnqG6
Wu8PvPjdJp3JzZaSnkleDLe0zKsqwB8dYtMRmqWLa3bpIO8/7AU11gmpoTAFdHej
9Skn1vrjNWVJYC8eHT3XR0QHeLs938cNvG17F5gHLwH2Y7E0l+2tL7BSCIC/blHq
DUR/cgcgAEsgn42aJKeserDL0kFBlKAq0xV05cMF3gGmJdZIkHKPjgKLsFgnqnvL
NHiBLiSe2PA58H2LKmiQ/2tMTB9dOTWS6A/UD3dM8pgzZHZXCTh3JIA/lWD7YVeG
RTJMrtWI9HosRNjAQsk9ZSKDiEV5MB4eI2VLSjLOJPsvx6x3k8rmF4nzoG8rd4Aj
N3R7erbaYnokYxb76ho8tu2GHR3k8/PSBQSZml/Wz1ND/fsraO45lwbq3NJXRFqb
QJq3LH8kx4oYkggvydwXuFz82PgnCUTYAfz7NLp+u1TaOKjI50NsYmcPmZ86V6x1
zwr9IYVKQTGQ08JQH1sj6ktoN3+3QM/t4zvAZRNHKJv8KXA/OqWgPN40FmsjR40i
CKwfGaZ1nAWqLCmaflekHRbc0iijocdxvkGWMWtM6pzXPM9vZ7yAZJ4F6xbP62ZE
UoAgqH2BxMCtNsU+5Ut7TX4KHv2NlLfwRaz9x0E1HSgM5UBe+0CoqCOFMcLkNONP
qfFBugLX7NjMxa8j30jTHhGgHik0n5234efG1t74pMH8IAHBPPA5SR6WXUM/KNhf
+XuLYSlrw1+gtqEEXEd1KoTFazeF8VlchpeklsbTifXJtd+KOwbBXSs0crN34Pix
qbt50R7eo1ddC1HMYAxlxRcxAca/xLHpeNxWdA3OJf5hLfXWk00bpm5H6YJJd0SL
HBfdMqqyXpoy9Tu7tOhc7jQgh5eq9oKcoddbMUlG3qVYAWXN5YgnPnMzy92NxRhv
Hnp8ZVRLlcUPsKoJJ/3Un6I6TnTc/6ulaFNG2zofK/9y7F3VA5L+r8/TNq0weqLm
6l4Qy8Y1a2vSrGslSMoJMkcTYRZwzx/YhdS33IltJ0IRXwQS2OOb+WZiHNStvTBq
KAHwzaZoe/AGMhzeIMPYu0uH2P4k+7LIGB165AlDMhk06cpwqJltfEURQT1OJfV5
llczlZp2nsZ6V5rmINeXo3Y57pQ0QFp6KkK7CWwVMJyIMI2M0Kf9aMQqeo6nECNQ
sYq01pOakLEctDH8mhj79mLjmaxlI3WKBY6lxGymG2TwwcT3j+KFJCg+G5NtZevr
ZXp99kMSRcFvrmutEEzEGzZUdRsM6uu/n9FwjBjQw/KMXEozoCox+lniI4uC+bdo
9rtkvD2qrZQfUDUD8MYzLHvrQtFmaZZ9+RMTvX5WX+RUnXuwiuTVTz3KymvIFAYn
R+hoyBVHzgOaDg/V0m8WNZs4C5eOtKdPaci2+qrtmObBpBpHrXffyBBGVQyc/P1K
8gjONrIcS7lp2r9ogHYVdGhb3D/GDdcy83FUiwgeRSEGrSQyLGOAc7oazwjSJeDm
sofCxu/bMgdzVn2V7WN7OZgaZb149Nq0m2DXVPxorbe0c20N2pa/pANaZY1PyHq5
O1TnYbHmGCelbg4uoxxVJZAO/YYI121+jHERvdIeX6kjHL1fmn43jtzbG+BrAKnI
2lJr6izqwxCx4/u2/dWekuJJTr0mODfd2CrDz0pxoPwIxj3VLqKSk4DU2dmo8om5
hiHyt2urdcJdpdHBD6JgVr7mwePod2TEwcz2EWBgtbJLgTkgKvga0bw7j9rrj2l0
D8HyjMAfNfrPIv4mWfHxwn+8Ghy9xJDLz4d/MtJPaX4tE2cd9Aq3nclfsIW0rcNy
xeFz9SzzkChZ7TALoG1XZBjn0tlg5qZ0i9BPVFfttCsRg2yMOSTXrbvx6p1iu4gp
/43JwsCbZDs59eRs3ZALERtQtLqk52lwg0VxVOI1sDRRmjsqGUg9xo+Su7EnWH1E
62Ykp84msPYWUB3qLaDgEttGrtpFutdAOoPXCAdTb94O4Is9ddidarRUUou7BMP+
kmwcqQPYlnT9EScjAU+iyyTGwiSNlFQ3Dnfqalt5rX5D4qWkjV5w0XFyGnbGWMUM
fHgXnHK0cVVrFasi2S/SMhw4Oklm22oLOZIpDzC8nGS5SdwCscMSIE+MF7QwHzlP
MKpkRzx9/ylgb7Dgpzd6ly6HXiEXFmnfiGMaDehv6peOguooX0BfmVAwLErQRnIw
LJyiY/woEm4K/sClK2dnKKDhMsQPv9MnoSjK/drIgPZ7ehEJtSuAVM/luhKqdxLS
BUmm2sAB8LZdS7lDSlcmh+1CYDkrhZDyuriyzEqdEHYYiFQJGn9hO7T9WcaFBB0V
Er1lBPA10W10wllbOd+xHd3Pqbk0iMODz/IcdUxjnIpXxHrz4kAFvoK+8HG8cXLP
RzsxK4LOyg/pwiYts/e8fx/1P/DPwgDjeyvpV3mKNUTo7NeNNAXp9dPJJ2oIPbi2
v7NpwAAP2OpkNfO4ROhgr/B2EMM7LJRyb+jySIrsK2K8nMpU5w43NhZzSbh5KO5q
6A9gGPqUmZgpvHufMjrXjPS4vPGKRrsB7WPLzPsfmOJ5ouc0Zt9ZK4a0bxWHrCV4
Z0/o/mREfLgrBm+xGnmzlWSNdGJhY4VEgjTMmNv8iapXSzTMY3pyN6HaHExJdO2T
Ok47SJ5sXCF4Mdj7J5f+JD/ZjIgzO7PoRQ7TLvgcWIPznXSXx22QCkMx5RCwzWkt
9aKNZbi2T12O4TK0d/aASrYuctTcctACJXivDZgBwkZyCjnwQ47SeQAVjdt76GQA
RK9SG8uXYDB2Rakhzg1DEkmgt/cXKtmBmn5plTNRXIsml2frXIKJhq24FCbdQN9V
QyRUSl+5FDk798JiUAzjseFAlBpWn/jOWaO7G2BluKJmMFh1kW6LTtKeYdNJGoET
xxOwH874GZF/tWccAjPlhl2nXKvASEcdUgqpLrh7bnYbr1dp04LUa9CfdW49BR7j
9GzRgFvKKUV/kKEwZhLwRNC3szhhh3vhdLSgQAp074AbRrrty8RYLC9cdXPtJgO/
HgKQCefc8dO6imMOQQEI5QAMntYVnXRJdaYEDj2VkcxKHM8AKwIhRpDMiqSJ255Y
UYdS4pbTp7q8+WUbvQxPdxU/UsF0p9w3xmx02HeQJz42OG/5NkxAQdXhN6d274sk
jT9L3GXJ+mfKjkefr6PBMOfrimEQ9ZkZ8EjwQQo+Hc+iq/5RYOAi0T76zRA9C78V
gS5o1g36mNpHTlEPrT5s6rjLxluUfmjCMo6RMZZOw8MF1xsKFpOoAto91Mh3yqHo
2uxb9eu4Z+EAOr2QGBheZeiMvIxvCUN2Q/kR+haRHgVnmFcExhAC8cpDw7FzKYH0
GolpJIDaRjMSIonAswb4s2fbRiDn70yHq7Rf/RaSBxZB0EJALAxEGhTMkSsNlqN1
KIxvzTchEolLoIl2thyYlkgvWXjblCPNsP41CBYRvHl+4kPFv2RcREW+9OjanY8L
OR0rAWwcMKGjQTtBm/dR7BJ9k2Y9ypMItnNMLwLIf7QD8dt/3J+hpHapc9E1UPau
XsgmpBSTbRhzEyyCRcNG09idVBYdzh31zeDU1pXygDewCx3yWhzOdx/TtVU0nG9b
dLjqBHJbSEoNuANKOgJVuqx6UH/5WFhKWDzY+g4/cvyuLmSaoFsm4waRn0/uiK2L
WQ2tjYthskt5m77EiBTzhgFSc5d3p99rCvEtgUyc+hM6ce/bmhDZqVCd4TtZ9Bvw
v8PybJPAX30Xoi/GcOdlIQS7JlgTZpWRY6YgLk+DhGiIkMW6H6nooMv2nKWSWG0r
tiSiI9sArNr0GPxecSUGv+/LyAIhOFwCVxrej7O305Vd0d8qWTmzrhGQpI9/U4jz
1CTomjlGOpR2R1Wpe3GxdB3jgn9iB/1SdojF0pNG+N5C4qOSMHEz+UbYgAW9E7RV
uVP1x5oqI1wbmauRf18styPwsVzKReL0TKGDBX4ODepZY+Qh2keQI9ozvleIh3Dd
gBrnGkOOMEdPeh7qifgNByd4zutFLAFsclo6fKbRIZ+YHoCq7E0prb5SR2ihPU39
WAVjdUO6Vxs2XrL3S4tQhZvuKHP/F+FqAd1IXXgxaVzUc0gsYHSzp8ZDEZYthrR7
jlkWj0ZzupiyWcALja3agPNFX0DAkTrleRRMRMLN5asU8poJ+pWAhkN5AXhHtSIa
tEeRk8uAchdjTBN/UVdCuXYkvAzyuoR4vv4Ja+/ak4Oir+GOxJlPFH5t7NVsK4jj
augHnC1ZPbQ1DeD8MgXdKQcOnyhTe43mNGOvi1blsANPuZX0vnO6kDdNHDmHJuMf
uKK8d1raRPVN5fBNZqXdprTVzOqGmmH97uTqh011uExt2ajypx3cPft0AXDq+sg6
NnSYaiUAUdg0cEe8FwVxyN3Pu1jLSo83ATTMaVFIkSwmklG80rJcB0B0ChYz6E4q
Fv8MNFJ4+ZxWiNTngRkxBxacyOjTieQSX4Aophcb/QBtr8xQrXVGoxDxGhhafdNI
Y0KsGrI2pWPcT/nrZkBysfdzukpmtmlI7ViTxUzn2VZHxxic+Whh9gac4sm9w0ZM
Hzm0AZVX4QOYultRdYlzVYDbuF67xFeN4BfNAwjdQ6GwOZPUJj0G+wQSDGTBA714
cnIGFQkojdnY6QX7XLXRu9fhQj5OJyExtQeIScF9jGPbHUPA8Rv6t1RQXwE1e27m
DxGuqWsP4E8scnUUJHqmuM2Yi/SRYGa6GOr+vW4TQg4duLH9o5xPqFzTeNtZ4MFx
nG5VnKanKWlo9im/OpYPvdj4dXJkBkMHgiLDodvuCvwU4zQ0JgzB/eiKp3fkhvoW
WXR1tBocpRPlxNZig89hrwo6MOLRmtGV9fpqqlg7TdTzev8l2bUMzPptxpZbhNvM
2Ss2xl5BEEY08LRHNLsOh1jM6qjHyz3rZUsO5jy9hE+f/3AE/T21+iSvqyCNx/rE
vkDs7xgWCeskYjACq59C7V39sDmUgeXvJc6WSV08bJC1YHY++ZGxmfYCNnT6VIBu
ZQ0vUvC9l29oeVgrwTEUE3fzqUk37g7Qu/6rFqzqrJkxwU/cm0OndUjPQVOFEQv3
/76ab0VdY92ASw18Gq/2Ct8nqtl7mGAET1wb7fSRmdhgJs/xzCLD4RB8MvcDfm42
kSCL/Mc6G4Na1YDnibj3fBv5pNfoVLD4pni12J0qefKaIed1yNtH106p2WBI+P6Y
Zb9MZBRhx3rzcSjF/SKDwj5rYyU+2bxcBySxskfHD1vxkv1o1PN60jXY78qEtw8I
JJVNWHtpgGstJKYKSQwjlD+B8BrpQI8J7dHf3w++4q8Dd/L7y4apdk7s009Dh3Ws
XaM4kfE56zGS655AFw7lKaaecC29bCWrDG5jumpMcs8UhD8LuJmfBItIrANYSS+M
FK9WnXHGtCYrSM9XhXeklfy+cbQh+0wz2mPdzbBWYjI6CO+payzCTX7paQVza/QR
u8s329GUJmRd8uulbSe/4J28byG0a2hr3n+bAy8lmXLxuYf99CaP/p3QfZsKwG28
BAj7pRfGayK3ifNivlR5UfM1CdA4/g08ArItpS/J1QDBFCCoAIOJ9PSbf4zLDX0w
RWBGDwI+0tvEwZwpS7yQTq3wfMOu34PvoBKwECHG8LHgGFBEzuZDzTRC3pC1dIuT
MlyujkwOImRgneHiD29eFtRbZTF+E8JrTKGKALlvZw8lnhphO62sLIvqkxu3leY/
Md6prEA/8d7TpKe+jxkT3tC8+U2vOcEs5kcevyzTMfRbQfX5cJmuMvh0w5a80xO5
+uJARjfJ2cEo1hAmWtr8+qVel2gn9WOnHQmacbYzM11rNKE8GsSDWlnR95BhCRAN
eXZH+QxFDYZh/goQGS7qqRbj3TawRlQfEEtCrACfPZyvWXDm545rqhaP1g4ed+W5
7/GmxktLUeeyV74fOmxrvvnOJW4i+KvgKJbTtv99FQT7k7VwFKdo9ecsBcCwPk3/
k1CC//2Jrg55RFNYNI4pN2IQpY+WCrGbhnC24cYEGdLfq6bG7Beiku2xDim3yJ9g
zbvEJu6951fOVIfU7ZgujOFnuGpOzio1M5l0hWBdSqsWSSLPrWbXWry1JvFgGLkx
7YlWum+xl1RapsOG5UWevgyUg2T+ygs5HF+P7fYzgQRAmCE8ULcjgrbjMI0ANggF
+bQt6P58iCqxYx9HbkWGHw5krea5SIO/HORvYPP3g0lh7SrDF6GkofWFbU9i420K
7br1JNO2Avj1aXsCbj0y8g3HsZgGdjnuQx/sCm1JbHFLdGDf3AXYumwIKf4wmwoE
Tr2WDpgqhVLJ7ZnC2BLUbVvRQCKZcJNUY+53t2jluxE3tgzKn9tXcFrmnPU6UBs1
08xHfDppORCAToD+FeNkzB7JFGgNI2vRA4hbAsvMXAOEiJ7YlW25N09eX7/fugLc
x0bQEPCTq5HBLitvOMeaYi8rKW9f7HM5dvSZ6Wqv58h7dWblHyyd2hxl7aM/1S+A
Kw1ivU2j01X9m69dWniVGgzS4QyaVQpmxf+ARMAOuskTxbR4zYHG6OZvpozNFlUa
TfYAa1EqhIM81Xi/+x4/SFJFeAMN8aJ077hy/46s3mdB1jqUY2msCvi3zYxHZtjV
Bei1OGeAx+BeJuuUt95wuBN8MztmWZNlVwY+kGT2HtFOlBfOVUAG9Ap763QvrGBK
drrvR4uHqAH1Ex9kI+XoBhjd5CJNTaR5UJlnn+CWUXLqCxgLeLLpGKXcrwkYrjIW
lfAKzzHEIVevjRW/mRTQLiQUNWrMSW0BR8c1KlNcRozNsTFZLvslKIzUFeRHRKHM
Vthg+w45nY1vPYGd9AuD9BZzvByWcWLrp0m+H1KqPlsq6BOCn6P7JqdIs03yXX/7
TSDyPbnvZuGShugylfPxjFMldm50xxVrA3hQ3Rr/+oTJEoQLQlWqwv0KYUk+sPCn
KvQL5Z06OcmZHZqHV/WoDwopDx+gkQQK7gRrQ1zREUq2GHPmQgLHGmSbMzT/rRFl
cOrOSdk7nnIkLb1MTR/thSoAp+57ObQRldMsMSJPA5+Rx3V5OS1P94n28Gb626hS
n/yiXiiQVPJ+XD3qn3jgPn+uJHiYHdN/7lRZAdu37HTvLcBZd7/B8WnplLeFLexB
pUv3jf92RoL/T7/G2tzSB5Ooz2UtkO5sIdvuuHD+5YzQZMghFE3QXAH78kbYRXOy
ZFeCfj36wgJtcOHhJkorQvAsJfvTXBmqATAXZTO42IIqhAPimW8PSwNiiIRbr9vH
o1CFMgFiCipwfWVo81nLxntdWZwcgA7aCEOYxTI6JvKxeK41tw5UxCcnZL8MAf6i
j3rybkJPVlVXfIrAjrrWQqXv0xTJhkOv00tVAJGBoiFnuaYo+Hm6jbuY5dXmDlzX
J4JNziv4qGknrpc8hocvHh7HTIUrinhPX9ZWPDRH64MCTS83wB+tNqyarD9gWl81
U/+p6aNTl4v+KLIEzZ3KmVKR+cbajdAOniJi9NpmxCA6qo8/KE3q+u1qu8c0rZXJ
BFQQoogZzymWR3lAmfVL+MEeB2I71QxKtzBa4q3FIKly33KkSDVU/WX+VU3ATpjO
Is+fuoKok/exbe2BdjTpo+/9Xy8kBh2DwJXjaWWakQcKMmhogucd1n4zGbsql51d
+3iO4dssQPkezI9ZKNRFzTH2IhQr3OB3SLO+NTNPXd5nXER5qzkhRI0EeG2q7VgY
++f+YARK6l2kVZDVL8mjZSAq7ez9FMJEcg1HnpGJNxi3OIadf2t7kyLROQup+feY
4sHcGc3MnZPHFa4lvxQKxYcOu4cWGRemGsWyaNn3fphWB882l3p3C2hJEVEnYCtB
xaUDQMpDByu8hYbz9kwo6cKmvDSVN1l/Tja1ouXosyUniRC5dy3VO7LHnOgebxLv
18Y0IP8eYkiFsJ+FT8+Q9zeWEmVuiJqRw12oryJ9D/j1J95jsat8zwZW7fyWS0Nk
NyhT1knwZ2/veKBENqvfTWYzJwRbNjJuXxb3hX38jRnk2b24Z/YBMCuZG/CuCKEA
ORz3/ToQRqF+mVCy6QXMeAjsRQ9sPcUQ+z+h+SXMonP3U6QwjOWTSYnPRkIoCuHu
ZFJFJnZ/x/zzzANig0j885WIQSzJHqvRN2RTY83LesxVx/7bSdRBB82vpKuUsMDv
1bAuq9QfqX/nhIhS8oWLJM26SlhPa/h9qkoN1uXQ3XMishKZJ7gDxITCaS0rQ3nm
2MBiwRhq2Fajwhe/9XNcoTUX3accHRtonYm2ZvieOk3oQ9U3Y5JpA6wzgIv6jQpq
RWXL9mjc9lgDuQGvA1/GNEKCVYhpzzDQYnrBZHRdOCfbk8Y+EdfnoVrfBkrkC/W/
wA/7lAn/2yyLY1umgBk5cdUWB7S2Pffb5tO4G4uIRwvbXb2UnzQB+KwnByjOyldk
fd+SgSjnVUktAG114ZkjiC/G3h21NYBZU0kv0FjQJ9ymiZN8EsIBdKLrBNj7Nzev
GckyUD1JV3rMJ/9GDhxgZDn+3nsmwNIh4P56k1HJIOexa24KjRVjsESLnLJRID7p
Bhv47We91WnB93TXDDvH428hN3bg520ub643p+MJ/jTS4WeaWGa/PqfEfG9kMBWn
yh33Wlyv/QHtqzMM1RF2rlub9UsA4SbSTrV8vhgvPaSqjXSl4IWw5UyvWJPMuHMR
vXGZXzge465RY4BdRE6fUscfenw/l4FXcFC/vJXOPeMRC5gHUsOjxolXMjCH7dHw
wkW2hxGgePdP0NkckebTbxvOQUwZQayJBuypWH0W0c/DxFF5sj3Xt58n6hNDF/lk
uoPXcX4XNzpTbxOtREKt0ipp1vkHQFcdgQitiGBcZ0NSoi7m2jw5XaX1R2PYgz7Y
obLnmfdzUNxGAl0hgQ2Ps2tpYUD8nnJhGSXXob1Kw/UlSd5g/qaAkZrTDf/Pnr6h
piCMW43u/37diHPgyPQpje0V5w2520K1dBcdHGcLxC+wxXQM4koqDzxFfg0h/xoN
vY0LHlvVpsa5/Glh/B3fBDBN/uJlWWvd/SXlXrnbO9lxU84ZzHfgU/jBXpAldqPJ
lAu+mJheZm+hGylxgyuGuNKyj7A3Njbqo5QTMeqMM5dzdmj7obxkjTyBIoQAUygn
D0fEpNcKFRxvXmcYO6dLjXdtksiY1KN9uANY/d9kIzaezcP8Vwoi/KVD+Uk/6TKa
ZRs27Vmul9Hjzsl+ItcB/FBTXzaRxjUuZs8LZwfTcjpvEYM5Xf1e3nelxPwC4Wst
aV/l3/fhjbrB7UnwTWw+wQP7fcTuqf/LU9SbNEfQWri2BMLD0Oy1jFtbwDp1CDXy
AuiCoYyg/p2mE+0gdTdNI+BKP2mPjUYn0LbukobK0qGnFBQDM3H0vAwe11k+7bDc
H5XLwTkYzvAhdSOhRU+KxLJiwIPcqp3cootb7MPyCrfni3Zf2BJ0R1IXg5WMVBhz
UT1ZImBmBx0eQfsBr79nvuqCWH9T7fWvPYuMRpTILOeAfPAwLERA6lIMPQIDtYiW
SI8nNd3KXiR1mFxI3Goavtyq8qOnHgU0JbPDu/aBUMgl4FLqpJQw6BJSuQi6LVGE
1ongbX1f4WU1iR1jWEp/WsGNpdrzn85X/ulBb+AAXPW6QebLDMCTKIN7Y9CndZvd
Aww9NHrR1B04Z5dOYizZFooIWAooQt0cUTXtfgEpJ32KeRc/CuxEjMXHfknhBYgd
eIkNINM4NlidCKVAvcwYbkvwSk1YgM338tcOg57OsGEqqD6ntWA1x60dpgfF/89u
8PsyveDCZyNk2FnZpWxIVR3voEH8V2/S1RAyNIDChLOZVb0+3BXI7cSAwCbJEaCU
7lmM5S2D5Je+U457a004k7jOBkoOf8rjpsI/yD0eqrgrFJf7nXNqDeiN4n/Z15IF
0z07s1/vvVDd/GijewYeMBI0xhLG8qNyxkFIZDtNArexf+Hof6T4sknEcxr025HD
EZViiyv5We9BL7GtyccQi+DPSg+PtPopKy74B8gR9fpvSyeJfunw/eCPIdEC/Wk4
C3Xeg7AR6XQyCFcCcwZNCgAW3S4yrfKJ05SADmMImxzIy8myBhDeOEkf1tzpAHjm
7NQXDu3xD/MHF0hJmoMWj+PXHdtRTUzksHW5+xNGvrMcc4qdJFLAJsceUaWjMytM
eCi5gfW2vWUlMPuuTvwLvM3LEQeRY0IEOiRwmEeOowSm2fCXEBnwWJKeuNpiyT4N
E36mq/GYzUOhAh4/4vBEq0hIDZKDeXIfkQSRJosdzBPOOi1ekBzhAHvE+9/MsexW
oCP8KRN2QyBYvvmKdLq4UMn6Sm5RfBTQXfm84hF0d6GLvxY0bw16OcYFcp8bMqxi
3iMqlrN+2Xd3nEEkSVYlmSy0C5Mbb3JVHGzRFyxALsXejgMqmODgKXt3OX4Pr5yn
QAJcsFe48+Uq5yBEBJzrUWu2f/+s/RwJHM5Z0rlKAZ9a33kYHk/9M5aX4H4lpedc
bQUp5fEkg7ZOr6GCe1gwrmEo/pUb1tGGTU/hyB2otIejYhLna4u3TwlV91sbyoUQ
/g1wQ9BSkA+aagr72BaKgpBY3utVSDX7ODbgu3Lg3d5E2hHPhVfjeMJk/Nd0M/Rq
1+M6MxxUZ8F7AtSRdgreHBMWUMzPriADnbobGyIYOG692bg1Au2x0TapkJPb/H/p
638JBTDLgiIZ0vC8dJUt9ijQk/eA0Bkb32T7b5WP9v+iDXUnZ8DLEYZACFh3xDo2
1M6YFNsd24q+bM+VffLL7+SHom+X0RSR8c6T1mL4iCfmz9GAyT6e/cHptUdbfObf
ncGPt+Shq/9EBBb71WMoRbo6fLYEKBxv7Cp1AU8eGObgm/uivzERC0/TraLTB7m3
iHlK6TgmI9IotDD0OsgMp+rXXoS90RUPLOVFtzvA+oBcM3kJIiR12HaripXSQIN+
8Ho2llKWmRAncRaqd8Cas0MXZIY0IBb2TEZc920ir+pSwDd+xi0NP3J9Ny5eacxz
0weXKm09svQ10nuSJ9AEDD/ZIBEbHJSfGI8GV1bg7M9XAt8O27XWKDVjg2mxJGRU
lePGFC1yz7gDmLAbck6jRv9t7JHFlZeiTJVz4ksoNJJMlSXioQj62rRGrvA2YD8Q
FdvNzbh5UJbRTJH7E5n/uiMajkPL7V80OvS57lfcYhDY5OUW7NTwdRBFM5fHWOL8
UFJk2/E7hVnjfVGg56WqG582qgbvjKoOOVHwT/yLHeOAHxEgF0/2I13gF4LLlqBu
Hgisk5IL+bFaHOfbsW0Tzkjai5CRociyGz61w/S4KAVh9Nbz286P7OGhwFAXbKS3
3iYbGfDnqjPZqjBMW/lUsU737rIN25Dl5sLwP8azmQouOYxe2IZYI7v+WmgzVsVq
UWhWLuIXc9VUHL/mnJd8142wBOLWrfcYEkHZvBdhyDDwRhhzUOsUymc3/+FKyX+W
SPRW62xTt45faccx1etDU3BZbqcYAWqX65saysBGt3qAh4FxaG3KX3Dy3oh1nYne
1Ff9YFC2onmET14NvsJnMB1JCoiwRq0TDqZnwrQR4pQeQ5XJbEbQ7jWnznphyfqi
IVqIlQPW8JKhhu2tcUtUepLZaAmZkWuUYIx86Ky8kJmtHrRv1M2f+wztsLxusbhn
qTwpG/oY7zwljW5+KU1/dGp7R0gxA54kV6FPNZmXQIirsCEmIN9zNJ5NxwzuMXtJ
F0WK0ZznQhgB0Zcn4AfPn+LaW3p/tox0s3zPRXwzjIEBHCQTEqexkvWMBAABVBln
5OK1jnQb2htpdvhe/QQpeSRN//9UeZ2FE04gwYARDW2sdygtUIYZacxQzSBRI82y
xu4G+FRXapcm2oRsA25XnQUmkKITruA56Y5q87QGrw4qPJ9zKKbBPTUpr3RZwcHc
vcnVdApH0S1m86XDQk4GsOsx4r9KMjnjMkgzSSPUftuPRqwP/p1uM2xfCxvLT31o
3UVsyVbqjZVuPIT/HBhk1LhH1qKSGDAw101ZMEBsCXZ5CsAV39SHp3ZBpb1Rx7lY
FMhGzdhrdvO4cWGSOxc4sKxuDHoFhOcX1KKtQnQwjdI+K/fMDe947Pv5t5ozLeQ7
74FXb2pmnxyifoKiMcsLypWwGAG+3wMP3XYFAHjJceOW2o7JmHDy5FZvPSldXpOZ
BY/NQ5egJgJ+XTd3zEBQ6zyDrGfPzDWk2NRBG5bEYEKmhXh7ktp5o9ppqQ9WdNha
ER6/ghAipniyCBqKfdhC1jH/d9hTRA4ubmR3xXUM7qBxJ5WBk2tE+UKM4nfZUUaY
tOGYy5mblYH1Ap4NrIfl2RRHdzRgTn67MP7BpRHNIPhWi7StDlT81mq4xpum/+bp
tG92wSAUMuAmR/bXu0yxawQYAOBMstB9kzuF/P1Tmy0fue3NgP7yX7vPMa+jcoEs
gJUohPMlv88HfE1FG/FwkRFQLQ1PYghc2xk6PBsywixYL8GMGLAp1c/O03XjY2wf
b13WWjmO56zpRc2o1OXFYfYof/EUmQUHe/+2wi9o/DjX7fMHOOf6QxttSxi9qt1H
XSLZ2kQxF9y6gwz4ilKY3O4kDHun8WmGB+HP0qGsh5NxzXd1iLMda1YNXSHy2FeD
kOwRy9GdMkCGucI/R1hhm4o+XxR3aOeMuIvVSAAax16oYmWUNojqx2R4XlP8Bhbu
XiurhZmJ4TXvSMAqLKYbj+QZ3c8h34A14H0D2tEiOOwuStPbqXkv01svMFxQjSTY
0lpU15G0Ug2fB7Hv7Oz0LCh8hm2UNSI7c+5nyX17x8zjqwv7+6IKfxPOrfQlO7Lc
l/jc7ZTOI5kvqHPodhJ8ksWgRxLXyGAG3copromGcIiPqLdvL9LNcUQ9TwsozoUs
k8XGXmDOIpwH2G3BHcS0/7mZUJvfUbKaOnXtWIBCAYynLNCrd6DFpFJGH2/qPgbn
UYN2GEo4GiOEUhhYZLDbVunxTUOxz0J8bC1Sb3hTDL1XCoydJDUk9goRD9jkTLQc
6ZxRdlXmn0CAbeWZM/bNczVDWeAvRXGeujLx+NOT4xgr37xkwLpDuoc5jqqlVrAN
M1vTHxAdNjA8UvL7ogQUDUAX+EDySeUnER5EUhbRMKyQEfqjB6J2gWG4p6ZuzCHb
hF8tlU4oc85C5Nr78KThZGy/U9l6OQWQ5u/4q62m/O7AV6oWYunzEWCukxax8D9Z
tddaKxJPwEjB2EBiW3Wa0xkjpiYWPqOMpbqCgWVDXlUJ6abc/kQgvuHZ0otiYf0p
jPHEPleInCydmh4OUDIHV+Q9S89xUaVSKBK4RGFUjIhruumbLAhSQ4TrUK10xcop
WkUSk4C+jLAdX5jZGf6dwnsTKZBpNEoSBc6gY+t9cjpq20K7YjI4JxhGMR5ywiMQ
UNzqVEb2kPBPmFzIWZlNIYU5LGzpnrn6UWKBs7okaaV5+ERJmXUgsIsBFJuy3WjS
yD3+SGHo+pEmwVhavYypPsbHc1XXJx7KwX9ykrWufEVHj+5aRgfPEattpGL4Dxpl
gY8zbut5twtwocXY5PretFFFrwAJvTyeW2Vx24zsH6kV3Savc1mP3ywMOyg9e7Um
WK7l9GnHMYXxD9X5Jgl7eKZv6I5dMYvuFlZG08+oo3u8ED6b91OzaCj+jDizOnHN
r2zn4KVGvnTOuEt+u/UcWrGN6KuwvVx155zYL+I1+AYMF4ci6pJ1ZtaTGaJrs/p+
bY1C+4VQTMLBBzvrWbJs2DFNBuSGy3U+UHfDPvVPubJNZXBvzC7Pi0KezYNPUi2s
23I7sMCi2qzIeUT/GLrUFGhUIOQsgPNYC8LKrf2Kdp15zvRUBcX16N45Qf9LQcpP
SEd1DHrdEZKwaxuuMXNFu2DD+66rHK4XKxmWClR2/xBnz9nxtu1tUtjTyGfmj2xN
Ogaq9oydMhaUttThZ5FiZ0VOD7H6XUiPkrnKtfIJZU54QLC+jyd8KJEp9+BprPL3
tHx8V3v++mZA5g0z4ox0xSf8EBG65ZHIkIguwMbZ71eVJ42yxELGUiNyRcQqjvLm
2x6d1NZXI4XX80Vyfqhm6MJ/LJrgTIJZtoBM6B5H9mzyLVDVd3D+eyPnDSD9VvwQ
KGsMBMml1zMQLz7oTi1iOUwfve1ESysGJS2X/foZlTla8kRYt3WBro71K8RMyard
dsf5NHN15WkNDz/frc6DzNSDkUfzMys6LQjBmGiIRaa/wvNilfSk3W+awXNRNRcO
8BKjgSW4CgFn5PsVeAfUXeDV9tgwnNfXFLdZTyDEWIZ2vAsSXtEX6EVId6WZvLUr
3jeWbZ901mCpGWwVVr9gtC5cpFOST8WVEMi1N1A5al5OyS7EGLXiCMm9x58UxF3/
D4PTY2jfjPL1L/tET4RkpuHrYA0dujhZ1F7YHe9tHu1WppuEa33B7Y2nNvwM726b
Z/roIzs8hCuQdTiGNGcTmk1Tbt8RAz78Sm6BvhdZqUF0YPJPVYsZaRb7hGpfsZsm
ZK6aDjIG4tLObur74VJLiT9VldY1XMf7MUuWeyKY7eFt6qVt5RU+f2Omy7bZ6jcd
MDnvl1n74ZwvFmXqn0BI6mHhkwR0Xa4RgCaivYUqI3m203E2GC7ZBo7UAtQjAH7X
H293gFk+8uMtX0yPXkTXpCe9aIRTm/u3bYhP2hBwl4WqG/hVEjpF4a/EPZ3LCTTE
gx73N4ROA+9isspDYPMUP+EqUMJjnOQF1lsoGuUiGydJG03zp/Lhj8WHFRlaOr6X
fy/x161oP3obeGt6mJYqT7hk8mF1lAC2WQxEXkjea+y/tQMrG/YPN7fGuHwXHxuC
gG7bVJzrwMRe8Yaq+pEKhrLRV3l/KwTqCDBUFC3Z9oczh0Vuc66TFj/RXNFjEBYn
na1hK+96qv/dcMEpxaZGkwm/pKjOVgpi25bPjyAqyiUwyJTuYkIjhwI3gZXFhdRV
ndrq1AqMsoiYzRhg5rFf0Jnz3CvaDaj7w29042IYNSsAmqia2zb5jx1RrVY/rpV/
LVgGFV82PH1ZVRKCxFr5uUc1W+/8KjC5EXvlvamd142vFZYeBp9D9hMV7l19+2Nt
BihsuQyEnGcoGt+Eq/iOQVNvaulgCODPuFWH/phh2d068k68alF3tNUd3BjPrSg0
6HaSWe3VtUnOMxywIdhMnLI5MneissEJckdyRw7o1Oj54bupfiRQbKl2SJMiDrOn
uFixa8M0HKiGDQDRyOZ6Oljw3QgiFMdMeg1XxEb03MDmwp+SxwzuLaQMPMh26LIP
/VsG9wDNxJeC0lMG0GNzOrxBN04RkQ0PT/HBQ0IROrUlSVV8THzYY9IjABH8CT9p
q+Rf7dCrpRRNrt0rbLIw781dUbltSB/vk+PPt6iFjVdpLuiQEkSRvvGDe5D3amxc
uEHnpxfEva2yj3V+Fy2BMXwF6N1i2XajbM8VJPjkZeEHxgDpjabQazpSQ/sxH4kt
QjpHFnJd8cmCN3J2izAfH/YVWlpzfauGnkuSXhs6199oW8UKBKX3rtmjnM9gMw8e
QLaSiIb/qDIqh7QG5ACnbZs6WBUPS48rUw0OQrR3CcSKFfPc01Vvtf78x2hXCafk
oaUPwHF5FW/OeMcM0/5ojzJGTsyWdzlVVEZLft3hZXBaN1qTC45Ub87Tx5szq44s
OdBP0u/jzzcfoABenj72VM/huv+iXk3PX/yG1JciZWidveR4xaQknEGYX4BWFrjC
cwXweL51hoxDn/zMeodpTylp5wDrXf1AJ/AYOfaoLmc4L7X8y8wQZ+cThtPTy7Sr
SuDKSsVQjMek7yvHc2bH9a//HXghCuy68i1ufR1ACVfh1DxrQjNjBODqUa5BP+1A
sB7BlDSxPBol35lKgZlopurfU2NLueAsrf1rhUBkTV0fyWQjGTyiNX3U4HqMw1+i
npcOcDWFa04gZau2pdDeFAhMmoPxuWphlL36NFlSmjDuM0EjR26g2KPel0qSi7Xl
W1SYPlD/0lEh9zWIVSs+BKEAmkxSI+nu3XcKMCuSTkezqZXyaCs3C6aPKytorY7/
r/I2/ctym9SEHF/QskLYjv/v9rwQYhqFzItKDS7wEK1dsOCqxPGV6cN0fPbLtCDq
bua95sDksvbQIYZbgK4wX4aaCreNAp9+eBWe9L8wh5NqAutCohJKIQAm1nzOLijH
9/tMtFUiC49gcBQoQpA6M2nYg6kFmIUYAQePAhMkHzhXToJOBj5cp5yoDQzXsSYa
NHtle07qt6J9xY6Q0BAoDbtQ9i+hKj8wNJJ1K7e2n4ck6GsjfZuAYRVAtCzJx0g6
3UZBlJVZFoT//XWk3XmHRunwUbzZMvTJBKNhLXzdbGoD1mcPM4Zzt9QUdnVIgebJ
Heunvg2DCEH37PKF6R7pHJOrPoBdm7TWVRMUHeYjttMLtdwxZpW2Ie6E05VIrzSY
DJGW04gxYehmI4umZORZ9+a47/H1iWkAJVp+hVZgf3cLWahdsCt9GxS6aXM9oudX
0mc6wa0OvGYi6vcmnSG6CG1QEl4w6g+lhpEHvLSziEgiq59BRJ0AuV1+whR9dIeM
yOWv7wg5XL9m/hZe8amp2n52bZCzmemEKVpvUn5lYKViBcHaf2qzK1tMm3BTlRBa
DgglBK7jI5o80nyrwtZiT5U8KXIdPaEa+ZAbTkEENfTOoo7UlJ/vmWub0RR+xjr7
mDkLiGWsoS0tXUTVWfwFF3RRIXGMUpIvnbHZzFT0bkS7UXoTTmrsctO19gzyGa7a
9yUageqAakajHKbSurU5oK6r0f8k7TxxUR12z4Y5dnWo6rudCHTz1zlpG424ZKN/
cst7fHV8MbArStKvg4j9Fp+a7ri9TYSGYwxNex5wDlZZMq1i0pb/vABKAsork8Ra
WXj/Vw/7mEKBv1XiDFk1Kf8oerMuCMVu38R7uHY9TB6jvZZWudBlKVMI9YWgG7iW
4H4jwgCwPxx3KRfH1WXXlqf+EFG+F8X0Jfz4sqxKamqonvw5B6mUV3IwtOvAwkT4
uymqcGzch6kvTi3rb5jO+xomQcgw/NqETTgxRug9LI0DUJ7G8xNOV4nmBeLQIQC8
VigX5M61P9cDLKo1HX60euQxT/yzpIQGquqa8kuETOPwDU7NAUimVvBEOTVesC6y
il/9S8Jsu44x38WdwDGhobrTmk74fohbEUp9mtarIbwIuBcsQ4+PfundP5s+BWeS
0YcOEbsO6YOFd6ueeXdHgif7HAgk5hcj0uzQbT/voQ2V5bxP7hp0Nkk9naY0b0NI
Ev2xn38bSmWgfTZQTsBJgmjRYfZZCWzh53itMf8Im+ptGSiczSHwwiM9JY/zrT7P
gr8FDdr7k8yV2w8+6E1vyfPgGbMuhN8ST/RhQnlMh/XYs9RKZsc9B+JjKdaqD15W
Ki+msZjTJqnNIS32QOnYFpaFxPyAIPKgzoQ/ttYaZ7PTcZqk9/o0VpwwxEZ+UWQV
fdA/d7XJlxxdHVfvh4xh5fgsw6sbFjRd0i2S3x9rMiLghVTmta+lk7WmKNpPhH8l
YNQ5BqBq5PNSC7aE8RVedLc4pi6xUWKvjtrHERXxJwkdAWpoLfnDteKb3SzR15QT
KI5k3oC+/9HpD6WrwNAzTOCzU2ueB6KMGPCMo/FEypDJXYKSEO3EPcEGJgazD71I
JGYxk29IHe9Cjg0kjLwcui+0A7FsPpHOxc6KucAoAf0cHURID2a53ilj8S6E5hDk
/yI5Cs01p34BuGlDGV5BlqYMU2Gye3BQJTjhxt5egeb1TqUW7xCRFCdy1Pzj9Phv
qlSR8/KKUKlkGhHq8jVtlsJXEwI29P8fho6uVUMU7W4DSeZgtnTtgAbbk4a1GoaD
Mju/sSV+6d+AFz23kW/KjG8+6C+8/EfHHqypypPqzCr+woPlo+M3B8kQozU3vynS
j/uZoswo4carvsQB7npy2evbIRNNyWbuGFsn/s3LxrAUnUDlfTjJLFU6Ku3JJo4o
NSMyE430oQLJXlAzS/GYvkjcgZfaR+B0NY+dGDDwpbdAoBGU+f3NHxqwaBIQWNM+
wJqkgZMwGUwEkM84XqQKyA7JkutBBCMl/fSFpwC+0UyJc5pYldVzowpxfHvIUWVk
Lu0LhQF/kw5VS26QhIEoBJeKHAnM43PrjncLmb5utr4EHStXvmAkihP6dKPAmw26
cHQBV/UbE+li4R6LDuc+Nmq4Z1siljECQpn/KOmjyG44wdOCXZ2o6cMR2Mqm1MgP
+IwzYSpnm3hjXp5ZQmkrH1ilgECdsb0OzFqMb/kn73ahd98a7VZRqW/ByOIubifx
0+L5cwWCDQ498NIkjMF8HBdJisun6nVEOWe3aXM3jZ2z7BcJxe6sMYT34vym2oZA
/dzOZxeurRl70Zx/LtUiCdwY1xrCtB9HsCZe5crRS9k5VeDIXVRbTsYBvzqV+pNM
CRQc0MsKT6UZysq3+5ah+0K9sRNE07sBMLeJ+j1SNdDM/NlBJYA3eC1BAjL/ZIkJ
Z7B2MJa+PFygrN1A9fw1zImRjDLfMMunEm/kF+TSwFF1wA9vPi3j46gpV+HHszBX
T3j6wWINbdGu3Zv0vmRJZ4X7ru/fYeiBps/Jw0tob0AEGfCkR9dv1rouRP4152/c
FGfNkdI/mlIfx5rBChG7xrZL7jdi4elNmv+5rhPdnJW9s8oALR2ucVLzrDx1NIdy
qen3aJQiWl8J6UYKJu5YzYPWVUdQ8gzH1HkXg3EtGESrc2+lt55OqLeIgKF2TYbq
DTgo8zIqxIU1eHVe+w57mz9yFNpVqCARfGSe2eZGtHHnzEs5m4ES0d4F1+eYvMIs
/6qz43zcYvKXbAiDp8I8G7zdS6G5/LqHFysqEMWZdQUDLq9nH5pPHuJPNHSQBtTD
SMNYsrX2GlMXKq/GGXRew4KCl9jHFtaJt4twPFN/RiNAmRKK7DBZMZdojmymuWQj
4W53/e3C0HYGCgRwit9pJu+SDfkBCPnZT7hBTdFr87XzdW9slLtk4DxAQ7oNXtXZ
fY/bN+KFBVDj80wJOCh7oU1wksCQJyGUGgQ1mRK+Fe7rciTubB2k720+MVoJw6+b
kjMaW2mqZ0twHGPP/qkdyR6GRQLmmE571tLKYSUBL/wntZy2xaVRFtLGh7vgu1nE
MNXx1AdpSNJSZeCa/UskI/Gpmmfn+GtdTOskqG5PEyQBRbVM0/YtRjEsZyp6a1r6
tT1/0l3SKsAR3Uz8vnICTaXjtqRZ0viFPyGhry+27NJxAAgDLurakBVpjnxokvSa
Sli6gxznOOLuwJXMcdNDZb+QmLhie3YwqujjB5+8S8Y2/axpbhAipZjf8SrnsX5l
WoYnP1HjFGfDklhCPIDQKtPAla6ELfgPdNi07DFfP5aKYJNMG3WhonMPnlX5L+CZ
CGH5n/elBZaCUNgvaAytDEJERpHaY3t0JjXwed371VobJ57NVFFlhUKRCM77xiD1
lG3gADeulhGQhZ5+ut8ee2uCYi5gkjNKcntYeTCHB/KSmk6RtpCHLgnvaD+ug7cy
uDK8T6VmckUxk7ws8vxRADY1/HshQIC2cuY+onnmoYcrk2ar9vcY3yEeGiJep3Ok
dkH6YRgOTtM4on3V8exwY51rQgqmiOppcPblJniXfOCQS5l/ZoxoQkFmbKKVL3sj
q0KYUb/x1uj+qqxXsdcYRzMtEl975nku5s+OR+Bw6ks5M11hEustfCqXTkHcIwLK
ZQXFR0WiHdit915XcS0+J+5Ku3Ul3JgDJ+K2uB1ThKqzsproG2XaAGyfBLefvRIj
q951WBgTTqGZnw0XSlSrTIzGUIEIof+hjH9nZokK3saVFNif1ww2zN/mFi1n4Qwg
UNxSNOs53GJDRZS4IoOzB6+0PAYoLZsOw3QGGEJ6zjP/EivSvf9h64GH1SSt1qOb
F8PdbWguWh3Li7FxxsVVXPdzIgOfZfjuq/rh8T+4Rtc6rtoqyH2doIRgtcb9BICK
VxfEFYvpGs1xb8C1IrSUTEBQCmco98CH3kWFEntEz+QeGmLjV9i5zEDrZ5i0XRIu
nHG7TzSa2c2Po6lVOpn3kQYetrhvkuxdHQDbo+F8e3xO7oZcIG6XgWQpBwhyhp53
HzBiulUpLXbzRu+/YKoIgl+inpNDQy1KHuF2Kx55B0Xyp3OYLGcEZyM5clzc+rhs
u9qo4TOVnuMUn0gNEqo/RTnD+sH6eqsFg79DVg/7eqRZeN29gBzGxsXTEBuoHs+T
lXuoUH0DYB4i7Q4+FhpEh4CyWoSZQWEqxuFCenOdxQSZsVJTYPAJyGP/810BIxhn
+anxWmaALpVAskVrHhwA17jM4Ez8V6JmgJzmzZM1nZok/405MNHvZx+cv8Hip7zp
pDcRi2sX6WdipBkzLMIRehOiDFOEF/Fx2iYJO3NcnbLxLTNQ4KMHLY/1CnirCsXH
ElBiMK03rnZNxgZQcG1gVtAVuOeWA4CiwDi0bykPr2DGJc6jXG/VsPcdAlwWGZ0f
rLX/Xq8bCv+TpxcIy/33tjkxlwKMbqBZ3M0sk5rLpzc2l+Px24wHU8VVYFkN0nxN
kh9WSsBeQQnYq1O7+7QJ1XvQRkgAAFFRR4Bvse0AutgGekFwtKHa05JsQez192Gx
lrSjjacUuk0a0lS693pYKJpzXYKNvX7dj8JWPew4ECE8twHb03XwbMKUl0fnTUSz
x1JbkGlLqj6ZUKIflWqb+1AmkAPt73vE7+88Xwzhl1WC5qAg8qhcmzSQAL8Z3KZv
ApfXKqIsjK4uX4JL+KXCmJ+4+WUQV+lPVnzSIvgUopVBfalrLqgrJljzptPoxps4
u6xPa7qWHTLhpu6RB8UEl/sqdsfgT1XLAvuvm7CQTvy/vhdwPC1zhdMHp3Ch6p+L
4q3LCQ+d6uguqs5kjIhTv0WzhCsKJAOj2GXscoT/i65kkrcSA6le9WDIPH0Yhqe9
AoydNEdUkCDpPgLVh4xa+v4yDZuZAZayoWkXnJUynjlgtVme1MXbN1xC1MtaSojt
CNpZ6rBIh8Gik89BJuJ4wSbIyuo+YlgAuHOLMIM/BVgyjHrYmHg03LDoDLwQeLcm
lZ93RpEddAETKDEOrPIRgdXWl0wtRj/SmTgYVi1/TIVW9mavz+EIvePUCfuB22V/
9pqKbZmyj5e/1MBdKfGMstX7J4HAJtZh0Wh7uK3NN/PoFP/3pkkUPB9gJ9w5eXMf
gpDtaehaaAm1fWglgT5KudTG7B3I7QdOu8VJjDFfV15OLg96ADINCJ1MjMv0Ee7c
qOJchQ8j+UoKS5KGTfw0VihENaddlm3GJBC87ThlOgHuRFiYcEW/+rTH9RkxPudV
lHFnio3iJePzDcj9r7FZtUhN7K9OarSNUpq4IxCpMZlN/Pg0hFqgtK0ylbBx6fAl
gKPIXgr2VKpbMVNqMZqC7BGNS88bsavfKfhlnoJsm2dHyFycQP2hclERVH84psGL
A55Twor23c5OdOs7+C1HJufUHmKeuazvtNt8sSuMDOi1E6HULJ61O/UGZ//I0fk4
qPUQPwGcvV5fnbffr/4BZkY1HVTDButoo9DhhZap5B1gN8leiMp7RTf+4l2ZiXZP
LEevyjOeMYUu3j/GX0Vy09gOnUgRMzjkKE6edZCLTgb8eCvftJJEKtc05VUUPqIw
8aW23v28VEUigvIv0Jaxv9eQIFbpvgfQ49My/RJO3TXIgSRdfNHm3EVWJPNN4Scb
j73YaVmHhNyQhRiU4S/au1Cpi1X9yEBqZBuW1GviOLAT4ezZOJZaVtuaqhNZ4GTv
7d3W0ONsiYV369T3C6AYeR40/4SCeKXm7F+d24qEVjyRhT8xlFVMw0DKHMgqk4Vx
HyTyfOgW4Sa+MJYNfDdUIrW2hWd6hREhBdHEchlVJ4ku6sRUWbVQtnNWytJ4IQIY
8XjBa6gT0LcjeHrvTZq4B01piZ99+U5x8xYX5C7jeUUvq9CMkeWkoj/fgb7v62co
ex/ERTG0Ojz4FzLzfmJOa0UCJRVj+bDbRtX0i0ehVzmxQ16goGKzPlJIoyB4Na8G
Rl3gFaf7Ep1a7ZQR78zgsHPmrV8975sEaD8kgBSNhavWnCRRnod21TlrnXbQJ3sm
mngbNBldlFEnH9s7YXw0C/VxIFWITWJphZ6lW7hnOcuduW8ASyn9QutP3nb5TRq0
cuZW3mUWTKV01vaPo9nr24cW7dZe020wZ7OpKO3eOyiUi0G5KDUE0z1/RcLh28j1
rttrXUtaMc9mJIH2WCEeC7/CWdF7hPQuh8Q+fjUlUkAjtFJBhorEq75xlYseOFyt
ggTb3OJHVHW8Wtzz3oqfZnEUg9RltTLDjjUy4g/EKzVqiJkxX9Ce3g2/4P5oKKQ4
NUv5NMFZHphFxVuEQoi5HGPDI4AMGXFTiS2I91Av/fU29K5k6WziZnXv6wPucO5p
ZaGfkRcgcGzmuPnx4bzkCk9nLy13uBeFgZVXnkvjaWLoYa3e7WptBFoiVjptgAu8
avTp2tUCyMJdAtTOq63No6Zg2Am8JVbAv+zVl3MPfjXCMQu7ZC1PruGp8+tiLkUo
l5M41euVcGmYomNPXDZBGNfrQh4P73mj3VXXfYXjDfcHiNhWEqMub4AE5AV3/MD4
84WvSORkdg3kka0RcUCPBaQx4Y2hWgj266RXH42wA6eHBqyNWvnhbzbN9SpHuZ9j
JxeOewX22H12y+5mgEKPeXPrrTVgmbXHHMoG3Lo/k+ZNqWPZkaV2s/rIo2LhxKAq
+1fBO+PCgzmVTx+iT/FM9aHK286BYrK27sbP2ddMxmZEh/m5WRLvWm9gBWruvE6V
sJWsgPkRLReMhvcQv/fwjnc35FXqtkbBqHSlzLHBCyGcHYE2lreoCsbBpIieGoXj
L7dRmeRuYiLwSNtU/7meC5GLTOI2MnJfnjuYsaj6cQjTFGJZHBxK/ratv9DwCun2
bY7YiqTz2e6rLM9tTYDKW9ceDB7hLd46zNQA+3RHY2Z4/MRRRTWq/hCFB8Og4XTe
3j8zrnWQ11N+HgquUVtCIK48k/x0laKCSwS9BSlFtALgJI3pi1ZHGv1M+p/KZ/LC
4Q+/t+um3Im7Q4fq1C0FpG4JHjaVQq5sS3np6gLcvGraouPSHD/DzdjsnGRhljx+
eYnp4DyjI0J5Obpm9fn1qrhCYZV/AuGneDkXBNJ0z5F0OLXpFR3cnMY2o0sLRd4q
OmUxl/opcbMjGy5hAzKQdvMA7QwWk//TbQFl18ZPs1TJUyN5AuZ+jhd3CYOPNxUX
q46aBACdy6NksZflS7nbwwHLrTr+qa8UeIme7eAd/FJROThDaSuXegN/Ufx9+HMy
jjPm9jbyyDaUBSupS8Q9SL8rfggBORpXZe4qGzBighzErSDW9F7v8w5hsy/F+wAS
yHQE0Wbu3rJXQRpqhs23ImamC9EiZ3Lzivdlc/JQ4Py5QwfDMP0142RyDmzIMaZr
XiU1AZlNC+69mkBwN3//CK/927XXxX5CdwVbTweywjJlLZEKp8NbM0YvFX4GMkjc
G0Zd5mJT4q3wcLr0hpNywlt29g9t9KEXn9kFnOqqxLqaNNlg74GGLd0SNWZWLzYI
BXKvNqprem7xexLLWCnA+4rhHYehR6VS43uLZBojVLH1Gq/Dhx+L/FSJJwHuar2z
eyxyTzTAUm0doZ6zwTxQlBJ9SrFKKGOHOc2Awm2R2PYvnJMRQvi1iQ+OqFUtdwfG
ctO+0NuIeFv7Zgvn9Jadz5oJe7YyvPdVv5lARsWB0hc3OR0O96Hq6qKfLVad5r+V
+z6rpRfPb1wwOfivqk77VROWI1N7ZGh7GczPRpQmxru45UuxTMFZKNuyzlARWxlz
/MonkJzRTBEhqsZllgOForwFoi/nXU1gErCjmC3C2wgbe4QIedYSzVXLt6gu51oh
8t7Bs2Rb9rxpbxfomTg4UzXBCbRgLU418M42b8YNIDSWq3wSYo11WvXnn0QPIRGx
9x2vaB/+gyC6k4kjW9ebN74MLAt5vlcUv45wv0jl7KFVjo29JSYM8idMVPs9GV3B
+ZnAMcxe6TUjKZX9327kRWvRC2XIxtFuzyNGfisya8aStLieod+iloxVauNY5v9h
XuttFGQ4voD6n7UM24itYOdokDm4zg+Chr0pbEbP44nQCg8hovdKN6kKRpoFxyvt
PdzgpHp8/yU/oqE3anlVrTwE3rBlK9tHhDartHAeJbbmvqaAumjPdgVa4L4oOhp3
Y2z6ujSGebnr1sgtOFZOjMCasgVYXWK/N/Z67uiBsvRNItbOa1z4OJpfhcKM7V4T
MGJlLIjy2uCEh3VZx7GQp0rhuAsFEZPizUR7RorETLyVrY0VsOozdMG4dE1PZ14f
y9waK/G/+k0xBYJoNKfZNTNwy67Yw++IB+U+e3lyU6fD68+vAHzqRskKUttpHqFN
M07I49RrRhlnrlZ+M6COdjTbR55KAuuCH6+YLY5bX+TFbYoloCTvWTt8xVmu5rTQ
sSjPlf2BtqL7ASWvncIo1b7clfsXbW1fJl6zpEaLcHHLmb14stPr9lQYngTmHINz
1eo8i98rcRWr0WBOWfeJhN5rzbnh48ob31Ewl0WHVrKm2f0QSdhc4YExfocuyixC
+y8PbfCx6C27PncQXTBP7WMgdYVBouLBMafAXuC4MPdrvamUnpawVUslLs71kgyq
LcgGXcHagT64LpudXgarMQT5k/Y2iZ4bstCdEsdaUppofjSVfXnm7OhFJwcuEbWy
JQY+1UbIW5OPN4Rr+JpN2pusQe2x9lZJMpflJZN+ZLwXAixb8vYYr7rLxdPHsq6p
kwPv4hIwk+uKNQaQK5ZjFoVT/pMLynASBukYA23jlRssXDODQhGPl1r4aDtdAwsv
3Tt0LSwwI7pIyMyzdkxCRXzaVGE0jSaPB38VJZEjPJi6eexD1KKJ6aAVXddOd+fy
i11JC5fd+KnIAfbN4BqOcmZnHB/oDxyk4z98XfUbg9+vrxA6NJJUMDIJqeJR/AeK
zZx6LJiMTbHz8+YuBI4vV9kSfGjtX7vx5F4fEcksXC5FSxfTqBtgKYVkk7IyA7J6
q3+umNG1CcPeVr31r2c+yGsj4ONtPoCj+6kCxnmsYB5n21V03kQ2oHdODVRxbkf5
D1Cl9M2aTOUp6dweNHjcW1gF83OeU9II9fo72pvbSvAsk2lI8k82lnTWIIwM0I7w
41yd0RzYKAyyXqyZKPEo/kl6mAgrmxzpuPlZ9Br/xRD8ILrNA21Y0RxjXVEopgWS
IJw9jeVDDgBhUpyuJWLvcuaP41MO4YiJe5zHAd++G7oIyLEB2cIQceJoXdYS4mjQ
o2OYofEg9G89eydGU23KkL49ftk9urqb8Sl8lMiOSmpH0wNJLRhNA3CvCmoGQhW6
AIO5Dz6Tv5QhLosF06hi0l8e2+NguP+fa/se70Xtma5l2qFM9MDGlitT6srqNsQJ
XD4Rlu6GykFhpWdeJI2WMKNPZVpCHrvZ/GhNxaabe2bRpQeLFE6awsFIvqxpkgdv
NjTAsMQE2v1suv+584fCv+rWxtqxx9SrWog+cDI6IHQ4WnBvNmrPaVInkETm3qF0
Lrte7yPjy0YlTVj0vnseUHjXSjkPXCLZDhtb5UkTKUNQH8bY08Jt/4iQ++DUlPxK
3vZqNszp1FZScmBBFmT/OOW8A5vhxSSc1npkCclzckvl+AyXfu1eV2ylIjgg5GMg
EJsrL2eZKbbV/rkMkvcFJs5J4Ip0/vl5OwqrE1wMLtDBC3hl63AgnAXUd6Vy5IH9
wDUawqw0Lp8gefAh/7XlkVfgIjkhVGy/K6SPj3pwap7s374dVdrKI0dHlNWFWaWC
+Lh5z8SS+Mu3FKiL26ekz4eTKZM2/8XaO/C2r0IWWFdH73q8jmnMZ673EF2F43jk
i4c7Hsao/mc7WEfV7J/djoJwqXiS/B5kjaek/dVMm7WHDG/+winzzLuttU29/UjT
rOEcgFxSe7Z8bkYsb/oYRpK0Vg8SS+6GHFBD6YzpqQ+9ZfSdX5tuC6ig0OAGi9xP
h+auSMt7qQ6kdrhs4X4avv1lJKIa52mRdeZfle1yZps+v/p3cpwYJM9MUMhKtMDN
O/TLxbg1wa7OO9/fQ1k03R/xjD7IF8AsMt5QnVBn8gjpkNijgh5WNkQZN0CTTvfY
88iiriXIcmePWaMpLmenTjq+depYturVBxmGBGzOnvyPnEv/V5kXmlnqtpkxLwBn
WcwEyHDSDG9CLP849javdHenjjcS2zZRoPugfamLTVosL5tMhF4YOZE5Y/NzZmLS
cWzW6arygbX1gQZ0neg35dsnfZrl96HKrmXQtlBSgooReHoKWvpYF77bmRqvBC70
GsI0cIFoYkWox0YR3nCDLaazghrUDobvtwkjTENiehcOX41ddQSQmf8Tbbq5DtY+
CHjTTmQGrfXV8hJbFCZd3bf2XOqSEk7ae1p5ELVjLd0OXoPPZUw48jgGWJAHsDSP
EeNx0L4Bcx7H9LeGVg1m1VIK80oEShRaunfhLMCOey7USlSAe9EJgHQejw3PpJsX
xsdWqHanqlucn1imum6aaaaECWfsu0mRVIOsCVqo5FIWlUO5vQwUuNbYZQMzgn8s
+LtrEMZ03uDe1jBuB65qz1/SakVMT5YSZ1uxOqyAzjkP5ns9CoGfnTrsthomq0Kk
loulBiGHaCbN9ImGH27NqbVyNmtqgyv2ni9rf5AP+WLADMj4QNtFRunBwMAXghMD
3C+p2sROOEsXu5QLVz92+FbpZDMXGxcmQV+OaDdZ7ZsisQ1IR7G9/1iPfasuv/4U
DCx/VyvrDWGhmiXswQYKo2ekO06k53iJVVS4bHskoGBGICcWbTF81VO2PZN+co+F
S+BidJ3Yap341UfhR7WZmKELfgaVKtP8n1McCNpBHQzXoWV4YEYIOb/z+//IEIbg
J8izBOSwbOUlSKZihyzj223UTtQkxlZNrHnUs9S4j1qtm94SOYxXEUEFJH2jvtG7
+ztdXnPKYyvzLPQW1H8zAmxjpXDqpU3j1WS7t0rafJfGpquwi3HXqG++WgZQgxgs
+b8Ld4VxPnC8oaxiwClUaGeA1rTmDfNOnWg4LbRqucGTDBY1TEIfldQ2Xu1tXHME
zPA1Fii5sUxm3lhShDy4MPDOI+U8ltppr6ot1avja1QCbombSpnPL9lDPBUGfl+M
fLjTyePabLXYl/tDYNv6BRDHrZ/tFzzr7i97TtRy4rL3N6eJ2G0xIiqiChRQEeBi
uNRYTdoDKN73Ja8rIFm+pOGl/DNKD6Bl3sDYhQHiotfXI4pewX6i7dArbYjs8/fc
QaEwhbD1EshPoDWy16/0g0jgvbSw9o7h+xr2PvYfK0wDvZRV4eGB7NfQcoBeDLDB
nTIFR9M7X7onQPXyj6sHCagrthiABC+Yb7WJipuO9HCDNMIwkLHE+L4OJzkBunya
PEHdNEl3sdJM3G7MPwwrAmGKlWs3nQvCRG1mr6sqTE1hYT3xgPl5zMbSjcAlf0h0
73DTJWRTWKmxEQBlFBGkFOUHO4vHNx9oKxAixJ7O6h9ryUzSExyj5cU5kiG9gWJL
4Cu+yzJhUYlKVWymavRRJvuViEHnajTV4mmsVLEL3sTKjjLxwKcrvNowTbZUzVVq
TQxc5RhOQw/TEWSNsdI4ZCCGEzGX9P0EOUlweZXzvnunewW+twwFiSEv0DvL7Fug
UHvQPy3Y/Y1zH4xseZgeQfm27WTZDwt6njCzzkE1Ym/BWNOsSig13XMeXRI23fjJ
/ZrGBpty1LBNZZVcxpmSQD53NskK2o5wjbjXpJ6szCz9aLtqhQJj8VvrBMm6KV3b
JBiJt2K0sbVyOi3774FS64tfPGaC+VSIbadEac9OIq93kqktk84I7LZD16/o91iK
m6gGayY/3SI6DLp5bLGBUkLccJReJ2SVjrNMYrRQiJazW+JMWXddgO+6mNTsiErK
ClwfNQnZYgGsMrc1WIVUifK2HtL8w/qOhZhSSFSwNXJBML24+awoIn9jlRlXQ8k3
vhYfyf7LZ/keof1nveZgPer/y86ITN3y0OBQgJXpHgUmK+qB7zZia5M0r/gnz9HJ
p1iH8+KVue6fWou020Y6gyQkBgGn7su2TFAVUEhdr2ifrH1TOIj0B8HkPuoMDb6n
mEUjkQk/wOAUO71f3LNutCkO3zWhq9fZMLgdcEGNjYFa4XXyYayOQ8doaDEp0hUu
dUJaTuX+Kmbiese326tbZ9Bggt4kZ+9+znc0dgPbycyqmvF0Nl0awSMfZLwsrPu6
oRbdpA05UvfsiTEwWJ3K+U4tftiQrhw3y/F0evpb6kv/nczKzhSXlawY1psXnk5E
fq3jkNYUCzSyx5pbeuE2Yw082+tGkjIzQSb2+wTHOBfPFWgrbQ46acU9AByTeprV
Du+c63Y6T8kp5xPS+yDnPH/iqtStHu2HXHkrkT7OqaccUTHqdJd1SRM3iIr2ktUR
1ZQxwVs09yAtsG8fjaC917kZUrJFqbPUE9OBBsJow+UI3wewN+cO4cym2yKVeJlS
JP46RyBXB/vZ23x/VoNOBagAFgQZSr+ZK2ekhKTJrwCP7EKHOgtgQN0kgQZcLcgp
JuXC3MwKLrNgmwyY2iM+NtsTMmLU3JCoxaeFBANuXbalnOpX9zWWZuc0UWgJO1PN
UX+a18NmoTZR/R1xOCQfPLnIG87ks7mvNyZgTa6fsUG2Mnf/nMNORI9lxWllNaA9
GQ6lf03FSs6j6pEH7OxI5ZcH3r0vaDMguMWK1p0p5dzmdeWt8Q4GpLsQquHptyZ2
GKqrdxziXZdNh94pw9gCLTTPf/NizvUsiSVIuCfX93q3an3PnjOZ0Tw/jcfSF3r3
His1u13vyFGsua67fr2EbHuBFeOw260Y1tsmdsTU7UqmH/GYJbPEbQzQYVEjmk6o
hCEjPRx5tZK+DjOcybIL1zydh3mfetD6ziYo15JvuAMiIB+cWBsdpLfonnavuoFl
FjqmLKelLhzkPqaW2bCyyFp8GLzXYwDevUGMIKfyanawZzA1lFllWm/hm9DXNujH
g8PspqHmIv37C2Vn09CO1ik/IMXy1UBFJu6meFUeWeQN9SoetuAwqWv/dJaJbs6h
UGFti7bSm5xBki0nOi6thnpeJ6UxHTP3iLx01fzCRxNtiPEupKnfl7DVdn6u93Ft
JkCW714slDWKsXA2V5w3lOZg3nIdTm1pVyI+K61wJePRUKr+m57f3w+yTweTGOnm
lRIqJE8QdodQPT9cCkKBQLe4i/7vsCSxYX5u4C/oKaHMK/mbPDJAAPVTG/jZEShX
Caq8H4yeSw5uLkaFrLZjoRohMgqqVh63erVu6I2Spy/VtpyNkOlh2qyZGqnsvazs
Z3ggK3kZgpHTkRClgcyc1rKw6lDUFcAjsPuTKjI93CB2okRdtOXeIkckZAMeesdr
7fXAfuySH/d6kPBeV7WmdCmzGmRvrYDHurQ+3toX5NOYT2zZonI+QaFiccGg94S7
sw1eWoo+PVfUH+zB3d+USBO2c9Bta4BNkl11ZHN+qmeOlYCC8Jq9w8xh9hwOvFhg
ybflZu3/buxk2fkZTDOkMSm8XBC1oXLymCJuA1KiuOp9QEN+FuyAqsE9vpink1C2
CNX53lUgWgGORX3zhNh8h1vFDP2gM7eexOgClzv7ybXYORI+9yw60WyKP1jeWDrG
N/bDRefnpRZUB4omUhHNjgsNFEfZYYAWpvuOQKQwh83Yo12PrmSV28WZRSQhFwSP
DWblZe/as/ucqeDLg+lDWtw7hd6jkKAnn3ja4ahfKU/XdQVxUpG4jjDDUjazcB2n
xnscTJRd4NIfvsTrANfb3l+BR+IMHowEOiFfR3NXsYagugkN9dI3tSDn7gmbWelE
v5z5gBKX1x0ckhOcKf9gJfSwCirWc6HCy8el8YjS/iqA9okV9UUbqVY076l0IOuL
ctXQ/qrHvoLsNvhTkJMLYX2ck0pU8lp4B5Fw2kkIRFj8fFzvzlTRgLJk8tCYKJxi
h9qovZjV5/CWLAuqZrV7eSdOrPsYKDkrZGV3LezbdBOfjKgqkEtw5xorbhb0eXf8
4zKb8PCOzU0k1GpoZhYUidlYDOezoaqOJ1E2Zt/Vaonjgaz3SDTeoI4P9GowpF72
yjr2E0+Rs61nfJCme/KQ+dyv72hU6Kiet1rmbMD/gxc1Cu8XoSC/54uhZEv1/w/D
b4HhhqhW6q683AzaSF7bvvGir612GyA3XWV/YuUyU6LSkH3AEOvBP7prJ4OkAp3N
MP+mOvzHSv3TgebdZ7oVAtI+81JMS+JuNwxpIX9B5lJJbTHkNdEqTS2VXdOlORN8
YddMUmW424MXJAm+w0mXTIQ5FoAwi7V4LiLlgem+OuB3bEFH5GiYjVgxpf2mz3Us
DowK+ka0CSFpqVg/WfLvk9FYy6X6hKUeBjCoTxM3nSSNF3hNyZbzQEGzKHeVajSA
mKFlSSgjbBhzsu6WvHux0niIbbMikOv6wgyGaPCtH/z8Ek/z8Atrie9O3xHYafOE
z6a57G39eW4gS2esmx466T8k0y9dDOUq5Vud+UMOReN2PpkJju+82+7aE8H5f+Gf
11OoDyvhv535ZUkEZE0JdtSQINC1C6jYAUcyrGsVtP/vXWH0NB426l33q7bYyt56
hRIvBnPdTCwsd5D5y/15fT8G3cK8dH/KASCbqu7djbcTgZuJohDCnKR16prS2USh
gwTQfp9JvMrrwYHTLjCBI9p7eg+DDrR9SyW+muOH1b873yKu2R89LAgCL4+1yQXm
3X5KbSQhZ7YvDQDM8WcX5VUF/O5lPir+4g9a0yI0OdMfwnBohZQNY5UcGCHK78bm
dswD+IH45Oxv5bvJ2zLv/Y3XPZVAITiBD0Z/6kGzPKyqwGDkRF9va5sjh8tRHU01
lkcNSwz5VA8sjhL4tfOkHMgvr3Pa5XB0myYO1zls9Ztaj76CnsIrlR76Wk5mVRDE
zBTFUUZEspsXgsEWqHTpWeODrs9WDuMwxGFuAtqMC8JjMVE1LF+FxnkVM9zK3hNd
CrfS0xec88TPz1nWkRmbzfkA6rk3XQ4bFmg0RRKIk5mH/HcaY7Ll4Mbk5IQno2G7
fDOlJfrmAYSmCP4i0elFPg==
`protect END_PROTECTED
