`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbS3IdrSo86UcutHE/hqkdGXsQRAbzfvTxxPy43Mz8QbWqA+x9DBSHFwTy3uUYGV
XPCbtvMoNBBUbjbglrtkFysU3fbdcj7+uKDCzhyZKsTVhHpJ0lXkKK6iO+amurrC
zvFoU06/4k9U91lt9YYkW/z+Bw5Rsxga49hXg79sSALHro6X59Ku19P9U9WRo33Q
r5BXOaMFHP6/u2ozSvGeDqzfDMGBK4eiDMOr7aasLR74Adn3ezBNce7avdV+4hLJ
O8kS5IJwAOAezqZKKW31buX5jkek3kAwaUrS49wVws8iy7B/BAJKMkLolNSQuoyl
gYEqNjkh1HO2w2PXLv7X9ssJcwmSnPSJpqwEURbZIt9Y5QA7VHnqIh50GgwUCyLq
+VEwFkG3F6SyiIBt4dORqlMAXeqtoYtiG7AALyquqOiCydBaQT3tEInCxLOEMBeo
EmdZ24xlmy4iD5EFPoGeVnxRNgXQl2w/B9u/9FyhaCV08g/ej0rECgj8/JcTovZl
j7ocbnfVOmMPRx3N64K98AuAkMgZ+z7gDnVdCVW1iRyw9SGBw4w6c4QBULQyB0CS
3dVDzm/YsKBj0SlzD4jY7qyOepDdd2kzJXRl3T8U2fBCyk9zY3azBLhCN7zJBmSs
nIkaHr00Z5aL9n8CJNRVOnk5Qr0pZdzlNVQhkBmJEOuguX/E8WQupmW6P/XXaev9
a3YEFAhLfsqQUBLds2CRgNzhO3JXQ22gI0nrc54a8/fVqv3HsLP7DffvJmoY7u/z
uTLu/lUBWI3QEt6ssH3FkOCcaCVUfZHplGT4BVC0HkangZ0BWcLe+e8JRSNRxiaw
FDdk1UjT2Nu8EkPtvcPIfT5bwXQgj0wxKc8gkxfWxjnURjLAZ7QLNb2IeuK2gTmb
HpzE0wf/5dH+CwtaWEmabDd5RFE3S8W5hRiQhEufa2CJQSyHrCQ7H6cEUJRX2g5V
09TtaooPQ1Kmu48nUm7K8K7cbdCkMMtp9KpAlNL1ukuj6H0pdyviBkeu3w88bK4T
ufmfAostjKF+zfPOcPtTEBUD4ZPyp4TQvKUEfON93R7ng2ClOLw940HRW3WmfM2G
/dbYArzkr0OiRYXGFfBabpIChSzDJNRZ3tz3j0K9X+oYi8qq70SjvVmXd+5oSYPj
J65L8/9vAcGM6RfkixQBgL74qRITkZnnwTU2d9+3d8xmJXTBr8BBc5woBlnRBhgW
NdByzbuuGbtVuhWbqg8tF0yBG2n4o/c5tYe7sC/W+v42eVx7T/lAT9Xev1G0wH0B
0UvagrsLl38HGDz4ZBE1Dz8DuP4RA8FPWlfLxydzTzBPg4DgRODx+C7PkVYZaC4n
gcbB0Xg8+hXozDrxCC9BYXzdUFxyuzFuHtrxHvZUM9VRjf9XQ4zOIeywjZoAMpQe
E/TScz1D2OfZv4eUqE/lnzzFNckhXOtB/if4DbyWLwTG6UTq/cLNLkjTegAK3ndG
SCzcnuANzg/+bZQjDJ01clrY2ozuyzMVnUpy0xSHES2vLBPpV1GEARteEfG6CNSf
GNIe486pOOwT/2SSpLXF4XG5fKz9P2NRQKKHGDyiJCFVqGYiJQOGJGVXeor+vBdY
NnotJLnL2x/07yy2rdKvXqE3OOyngDzY6zDwU+mta8IvYHF8jet0cN6hs6hKq3Q0
IdLyEKO++2Zj3oS8Jhukqw/HHozO8MeTey39lC3jwIYb2fQ76q9YB0uJhaE6F8BW
Ca1rD4tfN4gBPESJbXbY7LM2JcgWzaahm/IloL2kJi9tZTN2lX1e0we4jxexr7gk
`protect END_PROTECTED
