`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kFJJbP8qlIdES+9Xr6Hz+DVIOrJFi8yx1zNI0enurKuyAT883mJmCXTl+X8pCmE5
7glmUTLK2Z/Xh/GRTPiEd3++DTwUCZRaid6+RxQEHqudKuDNP3LI+vWh347Zq2CX
eNd7RlG38O4ayTUllpk1BnIOXnM17NP8c4ockpCuw5DD47NvO/vDwldm6S4pBDm8
yVqn2BOLiL5Yx868ZMD05AKDZNfMTntSXpzVfdcDFS86lBQMa4dpF6vUGv6babfH
23U/1BZ6ocNXs/7m14qqXwx+PyYoS/pdrSYJmVUBqcv3VteNvIVgeVaBBJ6CXlfg
tTAEi1usS1Rxijt1bg8RH+9K8KoyAneGyPT+R43FVKZXj6xDlpz9EzzXGabOEAw4
vUMR3XqeHlVBbVuailAkoAG1HZGkSUfEtQ7fx9LTKuWKdICNkrlEi0FGU9Ewg3/L
rbGWSZRQbfdxz7s+jh9Qtk8IGykoxybeuAtGmH4s6tes9Y345e9IY/BSxQXXUwNx
Z4RAHaQhofgsbLh7fYWDmdZdtAyl1NlCONJ5xSd608fQUJn73IET+KeHLLjgb6vb
AC4diCvXhp5iky6r1/78dFSy8rfJfkMr+0bb6TlQE/K8PQMPvbRDGlMuBXIAvHEs
WPH/40GcZAnHzti7hxkmmUGfgNrNTRwI+JRyec7RQfmJWnw8yVAi/7Z5krdp8yDU
`protect END_PROTECTED
