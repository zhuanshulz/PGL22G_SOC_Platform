`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wuQHuoqAd3rXrh11U6IHLFpWZZqmZGRy0tEQ4hSfho6S+ykvELIbdby9UgyfeMju
OvYOaYuHNhf0L8EejOECSF5m1AGn7EopVbz76cur3Wops2o6Y87c6fm7AzmUgFz4
8/QrDVyxCwc4WuZSnjMqv4yefdxfI2qN2fEobAYwzqj3CStS84LD2GKYXBySXzu4
sakbr2h/7Wi2jkRaQ7w3VzYa1ypBdZrHy2LEiNHsYlrp0wjzI1yKqdecv1Q9wjRd
DAr/UgAcP9AmEoe8TomsOnOUOJjtH2QaIGWJoIZ+bPKdUTZRuTr5Hva2k6JRjLHb
`protect END_PROTECTED
