`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U1WGtzDZMivcOoEjNSXzoHcf3mwhzB2UxglZWCpe7wkMKsBgVQQvbh5vC1ZZ6Ota
WilCx2ce2ic3m+t8rWk2Wp17gu1/hJQTNr/O2OgH15iscwXkJAJaxZABLjjzuNkZ
4OhHPIhzHMXR3hpW4YkG315L5Ywj0RiLbnfoS6sA17aS1O2rB2GN1f1IELfxkuGn
hxEhyw7aYLMv1jbKklnklqBZAYZvYoil6+UM5fNmFExnweOwkBi9ofyA6fOhHYV7
+SZhmcgzfjXCj74io6OPCJbru7IXpl91ukR6Ds8hvcEfJCOxuhV0RfWJc3vuwUFK
9H/5j34SWfPzN/B8s1hS0EDYWAsWefHqwSMzm9/eKp/SbGHo3w4xAEE3aX4xZY2o
jH+Tc8EcIfYEN6nEMIevTUMWVRFsmUM4kNcYCw17xw1SU4cWzGmHVhTLg7EkCNga
+iq0kpsm+8dXWcO2DD9LuYHYCnPGQSmva9uk+EZqc5Es9F9mMmILG5+2CY4PEor4
INkDiPW4W37aURyuOyM8wg==
`protect END_PROTECTED
