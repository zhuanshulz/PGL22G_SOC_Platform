`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnShP33Lqwtqxv6jqFWgOoT1+xxiEsDBJCou8LfXKuDHEtYXCDCUEPciBotyuKqP
PCToFDs3y+Y4T+jJupTtHQln1TERx4OnPeGuD82yBQQ50MILH5hutcQqYgsvSGBU
3BxH1Ngj8mx/ci9iu3v+ouwVK1RLQC3fhohrNvDZlqSAyiBfmY6OH1rQHdTEi/0n
p4nHVw6W8KDQpDRh48rIR/qxNs+RrYO3QeriXzhGkDNeNactcCVAove3wHONCKXw
8+C/m1c7QbXV2lUh8iKfyFJo7i7nJ88ZRBkL/ora6oaBWVMekrwo/7y9q+0Myxua
eryUwLyUeIgwJrmuit4HyHhZgmNQ2CG6bU1hMNpVqExEHygyLMzcEsVpCL7fbETK
byC7ozLNT47ZAScYvBFshwYpxhD9uRoq5J01Z2RLOpdkUYvGJYvXHwRsp91DdGoS
Mwkv7El9BORXHDQ3sjgzxZzgxlYtwDqLY98aRM9TUK0l7oqdGbYGPevnAlAjxHuH
SicFY+nS+61TpWvPs3DbSeNUHWDIH5C5pqovlRWVOpVKODj1LR6SC+CG19apKIll
2B7TreUtdjcr0o2RAHQXoXXwDS1irMtKf3gmKchIYj8vw0qDj8dq3oO66CfIl6cs
Z4C3146sXREZNWU6ApyERWDQsoVI8Jd6iAsgz3BqJN/slDz2nAmxmgGVFUqPMLRv
tDS5yomndcJTJx2BvHB3YutuEiTl8ExkRqO31GD89FY=
`protect END_PROTECTED
