`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQWclyTu+G2wPA2gmSCEX6L5MGoPcH0jFEfwr2Z5WlgpW22/hbjVzUGIkerZ3PfH
g+677OL+zmDe1nJVOBE7p1R0/168CfsNa2sAyW//HyXrnu/4Af8OtjkZSZ8V212O
WrNRLGQzE0bcGh/lNizWH5B/mBifpS0aFMgMH5Jgjn9b4yPNnp/BlVMD9KN7c7BV
LMLq6TZM9UMqI7HsTZ7DVFzYtJCiO4ygbJbYg5tS707NwMkaLXwJpMgsm+M6rX87
IzAMdwqe65SGcGd9sdZjyzI/w/xvf3i2Ut+rNGYNKiNOvu22knabajqukKb/vBn7
EOHV5q1NA8wEQWN5hH6x/BHA9n0WNlFxuIjyXcPKE4eI3Cwomahc0uecTDFq3OvI
JD2fyuaqaY35Fhwub1A/XDO7cb6cXmVIMGreKgA6EAvG43MJ7B2rLr4LXeVtod6C
7yi3b173G4JWVBzR02i5YTO4rcB1TRnTvedXuvMYiPVEINSe+9S3D1gDgmqGOC4z
aIzsZRySYG95ildMvzaqrfIrFXW6F4OzB5JUgRDVaoYkpnSiBBVgyL5KwF1GD7w2
UWQlxmHiphWTu49pkPOCifzandI3n8n8gU98liLADXGxHJZUU9ghRtS9UYTP3lFA
Xbk38p93oa14061B0Vi/HDITazB5sZDAx9o5L+e4ZUo2bPRJEX3kWgC4N08rS0XM
`protect END_PROTECTED
