`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUrkI9MOVsObrQHSnxVmIxhTD5QPoyY2DVd1lzdD7mje56Xq4gRw8wbI1htLpfF0
DXfLLkh2s/3SLMswAGhO9voLWk6MRAb6ACwsi9q5lAkqv/S0s0gfdjTbrrSBJA1M
V/J3VgOvKTQnno4XQPowBbJzK2FfEXlQ3lypLOSk9VHq6BfsITEvMGFiRYUuhmYD
rsBesHNNPU/Lmtkl0PrMmewoiE2vmwyGKzhwLkTcryQplaI/TVA9Nd0smkcIz0ud
H9h2/NQUwgasNcX73nuOgXZpV7QSNWKS+mknwWUjLQtVb/xNn7+0Vhl5ERdT3ZsV
oOvy4MzLYqMSJK2qFlEAlie0rPoSBrUZDvcpIZw170ZA9hll/9VsR2zNc9VJJtRe
KimdAI+F0IGGdH2SICCwnnK7dOG3ssRA3yYWRVoA49o0bLdWsRzcFw5CJHb48013
lhenJVj472Rba6GtR3Rk9rRsS0YJsbLpKMmm02fkEj6fIKebK/qQYY0njvIAU6e4
btxDoqvSq3lWbvo41DqMzj2563pkEEelXKBLBpjhQ2n7Ehcw67+hobH0lKsUbCl5
WmwDR4a7hr0igxne9xGsqti1wQLYsKq/vKGuKel/VqC6XPB5ZiGe+l6RnTvG+iMD
nhKk01l/V2IxDsnYvaqPBoDzKcK+FO+GdT59q6iDMbZ8IKeKi89jxE+k+FrDmq2A
qFBLyjS+yFskMUHIqG/iWbernBr/OOgxXeHy7RNz8EkLHs6HRpT6naLT9HqujICE
i1RmWM9alhyH1so9f7mYLqT73dQj7I8rXttSoAHqaRFuuI5Fstv+dJAHDfM0z8un
+FbbZ1zyYEVuh8RMgkugcJdP3q0jbu5NVgiAhG/v4x65gdpltoda91cZEBxSUeQC
KcSOxAbyDSnJxnQmLDJlxXBuOTJKckPf0Spfv810FAm0QH7H2XzttWb5127oAtON
gqR69T5DlEybnMuxfpSaJNcNLcck6D9RjV+goesMrVQItCkzqyflkNEPUWX5EvnJ
uOTRFjeIJ/BUu/cC5uCzOA8DXTlnF0MSC/UKeY2losamxE+FhbNV/g8HPs1cVM0B
Q9XWKXRKOPPy23FoaknUS4AXjJD5s09pqbQfZSQ38EL28CtxJX23rTVaG8cg8aOG
sKR+udP0tj0IJwPGSWGeUPnEy19nit4RID5uldbK+iI=
`protect END_PROTECTED
