`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X6VTJi6nUQaMUVot/9dAOoa2cnzkljYt8YyJ6wMYTH8LDl4dlN2UGK9JKT1EehsC
mzQ4t0AiFY+BSUcvL8TU3//21uTlpUmpZzFYJ65hUQqBA/EsWXn1yrvlt+BXiuu1
zztcp4m6sNuAukWSNXRX3xfiqIUB+6U6hjIo/7AmHYAlr1ORDBq04bO9HN1EBWnJ
+LnSuOy329rE6wC6+qE+xQDQCsMMBe6NOtwJYDS3Tx5i/sWjDr4BYWzbgwLrZwfk
ByHt71wYpyEv7J6epjj2THKoxljiaGlgVeX2ZK5GFxWIWc7a0l90rc+M5/RoyyDO
Fr5+2Cy81zPAZS+yOdhToHS3oS+pjHElYSIE9p5GxRRMXpTbNbplfumpx0TmRexr
uJqPJAnudV5FO0okxjXRr0HwmVGdJpDhB3LQorPOBOPwvod08yFq5T8hTC96bQ/7
X4GLGS7vAEQ7um2hASiS9OqwbE7e6GJ/L8rVde0xjOGZWmsSS3o2ULe6j5VQqtIk
A7UWh5aZXZ6PvEGOu6kGBlLmdBhrfTVh2NDKk3+0JlAX3C5Cx/dh6d15FoDc93I1
UhqoGr6hzeFlhEacmKELMs2Pe1pDTqFyq+74DZLfhDEMhU9dCt3vp+mCYzn4ee/N
BcPASl7yE68syvVxwvpB3M37kI9SH27W96horxeYzHYYLu+2fX2TwZ9tYzlNdefG
ireqrSa3RTNE7U6Yk1+ybZv3/al0tclMkzKxCJ0Js32ZGeVtY0FjKtLK6rwmYNM5
PGBscqqMTd9kzoBe3JEYT6NCvwuBE/JCFMub3zEbVHd0QWueiiCHOcM1oF7Vrdrk
FLuCYbDc8iJ8M9nqK1m8OQzpf3TI8DHewbLqc8hFm1mjGLq4sbohcHPitsH7S2bN
625qh9GOXAcXOHLgE6ZduBPzMkVWseaZhN0vtII+ar9/Jo8Y2ZCHy+A+PcqWng4j
upKO6OpJfjrCML8HWV7wbrjfYRzxmgDK+/Fgfa1oEGmrCgu9whTXjQl9Oc8ywLQ5
W+khvcFMSfu9AEmQjoxAnJi78kcLiIHzzuNG8X0KmA8AnPuwsQ91DV1eSzkBZbOw
BGl3EIbl7MLhd4myzTMESMlmYSJ9+qzmYPZSjW5EHjEflwvwl6nWhq08RPtJEXy/
mK3+1vdERDvXsEMZdJq1yaNeLTF7RTQZDFTMO67woF2HmGzDgRDdoStrGcUyfFhZ
vJ9eYsxP85bVEBPclU29tHqhsis4yeVzplBJQI5DFIWMCWTcP/KsOD/C4sEeI9uZ
XzvxVIdnKSj4OKY/0JFxPbhnaxNs6yuxQAgLfnb/b260vs/I6pNw75umj/wS858F
zBR6gdaOo82c62eZ2dhyO9n13P00DeNpTwKVRGdHlXmHDIVFWvv0HXkGqPGC6TqI
I3CVjjAkxxcWKcQro/BEuZYeRz+KnfqXM96Y1Gbb59fv849avgIwF7sKU2H4mral
df+fUiY1+0ROaFljVNODnpRxSZ+ivpNv4+8ZirhT6StZy2cf4UcR4n3ABaGco1vS
DEA976qHbY/F9klHJe9Sso6bdGgODzdeuLZVrdWUwV3W+ganYD9DySaShrmNFVmK
216DRI5Ilk+eWjLaI9IUyMWr3xG0GJjK14D1cjtRsX/y8/kq8c3aTyQVdNAEXSIG
3lattVH7AQguUybLk5ofW0D17yPXS7rBb7eFHLZmYuIamVfAB98g91V4s/EvCtpW
22DIVfsMM09Rx2am1Gd6bsCgomddEdM01W+MZoxrA8pRERXjhO/iPdEl5JCVIMXs
nPI2NJymxTkIM86uo3iM1Vp/NJxJ9xQ/JAYIjtd92jMZgh0Tw7QKIiLUyGlaubIR
YwkCzKLcJyT7k1XXhO5dj6q6g0JH4MGZj7enZQ2RKmw4jsRulYrWlwjRC20rOXg+
7KJjkNxchMzRgu3qpnbxgzXmucH2sumrJVXjliRWZqaDuRzFORupLK73UEdzKsgL
G6SbgoA8m1vrC+ah7KEYj+CXaLPo4NeNOv20+OpzTy2TKp8sODGrnIphOMzriXaV
sTiGrVEqEOi9YSeL9Y9saS2SdjlggP2G9/ZQrcPONYGTpYC1wvAFIqlVJH4Xkzg4
SX3w4Ln2WRYuu29NN9/QbLL64MnTOZNLFikyVdZOKtYJyYqtOxHP2lw0Y8g9ZegS
+kCn0KXjBniQrcSzWcKk/hTOvr88tqrp5HTJHFomivrKFZ8RkFCYOKMyHK+ulXBY
yB3f2d0pxt6v/1Thb18vj6tKHfWEvYktNdO6oVHAaRckgiPFA3o+S/jKV/HLOQ5z
gjdv2tik/rvIwP6KGHfgEYhbXDK82JXPSo5QG7W26lE6OUeCbTlcqHdgvMe1R41T
m/2IMZ6oUGQ+YfTpmeCBJvtGufbBfiL7XduQlrOufKuVgnYLFqB4UxYCcMpKBYVl
YmZ+vB0ydxo2dvBf337IUNMDy3EpB3qW6V33Anz5aUT6E9KBTwqwXnrEGIsb7Dkf
`protect END_PROTECTED
