`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lqQY/pC7+HhbcAx1k6yMntEOXvRaZBq/r7D5VtYM/QIt4l0HBOc8WBon3aPJq5Hf
+QvX3bvWtFgCWV3YHvZMN4iUexBp+cIBCNROEkUjO1HTfqSn44qau8yrvLR1DQ4V
0/ZhQ8f3ESHanEdMEBUV7cZixKylu9omu5Ff5m+7Yspf5lnLf5EpCM2gegRndl6l
gewXY2+L7REDVVsaw2J4CYrY3gsUU9xlL+LUtm9NckwbVPgSY0myyfd2fLXu7wme
kGkNWHaYF66epw1cDxql1w/GjVpUH0ibEsFehdXzLSrIkabp0IKpQlqh2Vf4DpD/
5xVJsbU0dd47efBOQVg32SJVqFeuRQTh4uALsGnvW/y6rkh+fXWE+P9w6vAceIEJ
owhlNhpe9SllquKVXn9yAAS1+CdqJ9H5MAdFjewl0KM5SD2VDFmpOXjG6PJwwwrF
L3NRuIKBB5qGOWq1ZeePAH8QmL4bz7/lBZuvIWvKkRlTpJK4ACz2I/YRG2abVSEv
MFGr7oDuXfvjgV6YQYtLuu/dPCY69frdiiQwWg/TFifDht1WpQOTC0vy/jlrRRkg
j3kv4N9PYNEG26j94B966y0E4Q/1PjdgUvtiRSHjnToiZ8FAmXHxiK2O/fw6aTqW
7INDR3W/VR3BNjZYGuMIOQuWxQcYknACO0L74H3tfIIPDynq/ZrkULwSTdl1YzZM
y/Xvpbqqnmh15fr3O36Ty5zyDhVUfo9gbkzFGlCpO9kpVL9+gNHWzBVvALL8R0Qa
J8scIcb0oCP3MbwG8+IiNHoxG5GH0q1o+yJDKpUDgFzBqRHlXNSHvcY/sPsXgMIQ
V/TRAYOv++b22EADTBB2SayBprAgPHa1Oodaxe+tQEN874zcKa4350MhQaOfrDwC
nmEUJlp29Fr3fmhghVhKoV6HiCeOxYwAxiCVUhd3V3UvHHTPYRjxE6NIrfYnfEU1
zM8qhQJ8/xgiB8zhLAwwbQXhTD8vVOyi2JloWLsGUbQUCkxK4Z7qQbSnSERIFnar
sO0tcAwC+AIqNE7en632Lcex6LSwNVsgYLurUeuKoFe1Fot0EvkXF3/DQVWrj+uS
4k3Rwi06Owj1bt1idBixj+dSnzBVGuviGKeQkHRucfnp6TAxuTFZPgDqK8tYLzgu
oINxelvLSpevqEHL8ZIm9DBYsOPdn9kidzfy01+2x1C8lBLC0aZmsVPFFV3vKQYE
fXQTX/aaE1ayI8D/0j10VYU4QKzLabPuBr4dvDxbL14=
`protect END_PROTECTED
