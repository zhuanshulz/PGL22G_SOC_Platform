`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aicdUL2plSz3iOrS5xnfppR2kboJ8q/wXO05FdQQ+pr+qwU85MA6LntEEjaPL6yD
57URFBeEG39kBRvIpW7GhItN5bGmLsf1Vut6usR23YOTrX6Um1a6+8BliG+8KiPN
lpwyMcKesaMv1wbHu15mD3ib0S6MtQ6M+yZJ8uuP5Nu6pcslGNIwwmJIb4YzB/3P
iFnuQDQNUzO7DFZjRvNL+lYEQ58WTY0yMD75q9ONll741Ey7sByRivScTwxRYYxk
IKWhKKc6gwHt/3UwgLnJThXX94Xu+N7KSbskTbcnhS7F3vYr6yxsvaz+L1DRdyP3
+z6LAF9uNzzidXhhPPUobKvDLYgAfMdckFue/n+8hOO/+TsHSzGkLeRp9Uf+/HpV
aUlLiKO/v5Dpc/E6tPIP2rjNQBCr7RgpZVivIyGeAtcoVPPCwFV+GG4PGPVtmlM8
daOX/bj117WFwO/DlukhTAHn4DXjR2SsDJWqNpX7D66m2DKXFSbao8NqDuw7SzWv
rC2de7yqmAlfDovHoTQZL0SsT/WymE1dKvVAGKGmejtckstARQepUhIupXMHVqoL
zF4+WPxjueKKokfksHGQX3ltYrbHIvkCOO3aa2HzF+2p4qmNlzDv/Q5JwaCaIBFg
zOuQ9FzdZIgYVj1LMOavbOFipsAmSUTMvohag+lH7Uvp3AGXGe0c5TtrtvIYZYne
ISeqjICPJ/oab6wJPoPYsGalhA2MZcZ0DKBr8/HbD+y71f8HiX2xHVy+yhMrU3GM
seV0VeY69UD0FWIoyHuZoHWuMANHgrpmjzvGMp7mnkRjjP5x1zbLCyY7t3FVZtg5
rjBVnT/mWCeHv5cI0JAFvH0DWwqhW8S7zADpQXfKUUJ3fzfwpzeBNAN66HNHqptQ
nFd8/yGrDWiJyHkjViL9jymgct0Q+n+p6IUyvrVdRB/HENGI9H4crHveQBYrhTgb
YHtqawnR6+0xC35xe+owVkQEmjmPxV+ZoTaRxmOTfs4Zc3xKCDty5mQ0Ho+C+ebY
laZyGabXvUTyVdvV1IUDHdnAGIUT0vNJwu497iZu/85k3/J7W/N7ztjU99i7Bsif
GJ7W9Abj+/bZ8qg2p9Hl4B8SpL+rbEHt/p/fGDFSwTIYar41igmBO/KkDwG6Sqz8
0XK+hJfm8EALm9ME6oAAs9+K8xyO96ibkIxaoL3K55hPGQ3d5YsKT5g4rLetXFKP
LnAEJVqE9XOiuq9FZpHWOZ1zQzIo5vjNHyTcSvmFjbPUwxihsqOd4PLzS56Plu3m
xc3ihkVgwv7vmLKT0jjXmMti6A3v1dSyIPPFaohfCNp/zQe8RXcUmaDo/dztYZeJ
euSRwHQrHbJHv7ph0JInBW60Q3RiIFT+YqJGhjFuK5M=
`protect END_PROTECTED
