`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AJIoC2+YwEBLkdpmU7NElu0fIfwUQOqE/6dgdIZslGiQQDRXKNV0K7S6J/5cnGjp
kpQHrnDI+/ri9c0KSI3j6xDU+6B8+ZjuJJFxA/HSqZwgdTUvxDWki8iCrKqC0D89
KsOhVeujtHiE3Hu6CA0h+fspZs0LV7JCWJYkHGwJQOUS8bQ7TwXp0mMz8+osWkC9
qO5lG13WEVBR9PoRbG8Ln/3InQ912n6TnwkxaYoRP/yulWMTQHjCTCqVggOJmoMK
/IW+YWRWHbAEm5mHObpsfp4ewo9urFgv16Fy1b3QDqe9J1N8spMxW0Nl8RmEu1d1
rav+pumzZzdngfsA9zpD5AN2Exo+d1BJPICeTFKoHSjUl2YVhmUy8jGAPWfWAkUD
57Bmp/4BqzgLrivEAYTQUDWi5w3ibzEP1JqXtY3+/nXphNFRhn7M6YHHGm3z+KtB
aoE1E2k6LVqUzk0gibMe8s8t3yc7f9SHjRCBBw7KjJYo/qirwcSaxDA3lU0At5SE
x3kHxz8OJsysIjY53KmKvzJOZIZbst//TIUJVggy+bYQKSFOv3/1Ary/D18DxpP8
/Jd602yoMpsKk3smEQ3jXnAoZQjXYdbVehtyjke2QrAPIYIylJzzFkCX8pxYaNWe
aMthVd96F9UBQSzo3oa6eQ+pm2+OMX3X8LZwySHXOUensOaKKLoVJiiTXjcAWmgD
9mda2pPzqqQMHDsbLGUV7PLnT9VRXElZF5lVaQ0zop498ohQpSL9JAULnc6NFzoO
ZBepMT9834ychqmMhBN024IO8Du+O/0uC/IEHWLJMwpurEWeSbTBWC7/mhMCIL8n
HXiZBRADcD+9+Cgh9nvjUx2nRPtEKwsL/AnfRNQV3E3ZEumxMC6VuiSQV2WNK+Dr
h6I1jMqPdmf4pox7tKIctnftsSRIyTG9c4lbz3lrVfs7ZSV1y/e+vFnLRD2RFxrg
7pHBkrP3q1SHUGopbqNH5is7FpVo2v/xXkQ843t+DlOe1wjzmHD7+YcKup5eXeC6
05+N5XgKBmnItT2SfLjr/xAaQEu2+pJLYCU1XW8ohJRjAXzz1esuPn3Myj8ys2/q
7DQKuAaVbPD+b56rLNG36F4yKP8DLCMGiyz0v6ZFXq/xAN6GYWchvKxs0FydNOar
8/ZjZsZ2gWMvTSXuDT261KZqrEhBnO3S9RkDLASOybmhpB5gWiLZo83M+xAdfdtb
szvt/f706KNH+LH6zp62E9iJxf2F0FM4Q1yCHkQuqFKExeQ16ZIU5VJ7vunw1ERf
5AS3/jLUAoMWbhQqJSsJsNzQewSeTGLgZds78+cmTJGNe1GbfA9QV4WQk4NhBFNl
69Xxu+wSfnC3B+0SeP6RwIvHcwkICFuyIX7C6kJl5WHEC4Bcer08E7U0NXsGVAvt
I+lE6v2djCEQUPoezW3qnUiIa6e/jCbj71n32uvNKmQck+nSuQ+fHmEEVnnzJm0c
6QfCjf2lTaD9O5kLWkDpUYBf49Yi7WHO58/8Lea+We8tLVlFCYYqgMx8L6SGBVbO
yX0aTauo/76lgZfLuH5LoovYLFvf/HN++EErlAXv9XLut50uVPp+i5HfRNWqOeym
AodUMbxp1ynq3Rt7K6qSa58ozRTmXELUR64EgW0N6CCtAdp+ukQNUVRSYFrk9iHN
MKgBl0F3BfXeePU2FqxumiVzEwq5Hw2YzBvraF3X57myVitKPstY5nYmB7OGa/77
CxE/zzLcxB98ibPtkqKTCN9ShHewbqqNYBHwOnZ/0BoTKirdnupDH++w6fp2rPTm
9mJMkyWR+bt0VCZ+Da29Sf7B1nSBTFhaX17RoAvKGpsaE1LZFWw0Pvmy5buUqOXz
faAK2ZHBi6uq3pJFqFQ4pik3XXJi2rvK2aHIoLNHAcT4gMpoGib1PPaPa1MWY1KG
qnWU8hYNwN2XencUFR5kE1euHLJa3Ghlzb0jsqDlZ9zGVEZIDl0i8SA1fSRz9/vo
hWJdgGiVJUwuVSxpTTLA+rMG1tRn5KpqY9Ijmz47rDY4K6N2Y4ZFFtvi9VDmT8VQ
RV/kfcNiofMWqHeVbygVDAewdQ6bMg8ovwYVdGIfzm/A/Mvhj6/57Vzjwu2O18Yz
nKi97FtO/eJ5r+fuLPxGJ2d6hO+HyW2YTOUzF+kibHOCF4j0+zVyp6+167qexu3H
Nknxtk+oojKgZppzYIP1l+kJN6fiJOX+Iyb9BtIJ/G2+Drlgyrg3qGkAmZheY5ED
2kQen9WiDFrYcsYWXGJmSeDZoeyLlK4xlf5WWvXUCLUQTObJwZoe3DWCTQmPNOF7
+FPDAHuh4X4Fb2O8mlbWPfO5D7DK7U9+ZNC4dHVGroQ8OEQU/fdET7Ej6G9nWAL+
2+wR+n5XCx+hDkylZtUf0kZKU6SSTuzO86voqEfVmAza2VW2ZJTsxXsxqy1HJSHV
IenLkISFi7YyVb14QGQoFDmxrhW/scKgg6Itaw+mJ85onviQAzfrey+mBAlQCs0o
LO6N+Uifw6IbZURtGoS9Oaz5bjmeGUupB7boFMmsqx1BPEjD1CxikiHSbDeWRLj5
9MT0ehJDbq9t7k90CRZAcRLN8FalhRLlmRf207XNr22LoLIV0VYKjVcjSH+mlStE
SrfgPL4FALqGUXTgtwvkhF5Dcf66yaaJHeeKl2nBzgzVQi7Ywprf1YImmcH0ALwR
yIAnx4b5RL45fTAr2iY/3ieRFhv1DpBIhFUDITzZZujwj4Ndwo0VbRLkWf4ApzB7
Z76WJPEF+9894uTdDJPQOuuklSYRtdVYGbNiu5FLNdQt9cTJyYzX7Bcqmdc7ZB7I
Jq4pI+Ctqi61+FD5S2KIzCvLssoxznPHoqOGj3q6k2WDYgCSb3l2BRHUD/r9KrEc
jGPS9mkyhmn+BKRFF1hWdgaWl37H1tpRGvJArta5A9DagAr+oHkDtNSDNrStn7Ki
mMjFfNm3B6KAnhTFrX/fX4ASEPW6Zbh8mkBG5xZcxwid6fHpKUEQ0c3CnPJl/Ycs
zK79vKhXiEAEfml/y19+3zEcwnJxLcJbTK20BDX4eUqYpZCnu1GQYfqSfwbFH5BW
odNnjFWYISWlBkADBPdeEfuSAU1WzRcVKZIcC9Lq9AA+0fgIPhNkZ//n6v3CPfh3
5428Tl3ZnHNu5ODlgVcc9cxwdh05ir1RI04iGP994kLqKpqNVqPDStDBAOJI4g4I
jVDs7bOWuRPcGggjjILk68Oc16ew4qKOD0y3zh59XkUczLnGRcXSmSbebCYS23qq
h1PQYK89UDPQH4y70m9Al0tdv/B3QK2CC2l0xwrHcpvaXgyzl77rKGFMXteGXsgS
e6A4Xxb6+RW5jz5pTuNKU2lgmBSd4llFmmouQEf8gM8iCnwxebng9F6H9y9G1tB6
hJgvD2xwDEKTopPBrGVfGebSv1VbZjXCH0C8cDH8trrmgBmwSbsxmTIQ78BF2Qpz
64322mv5p4lqLRGjtLIh/b2oXtuzyEbhPh1lAcfhGFxB9m1qhPClcaQ/1U+tSnRC
s2kgkb/Tyk09RjHQgwjUXpQPICQoIE921IQzGWNO0RbCYPAUkFqWmuAdda9HMwkv
gTTKX9TIMsS2eUxEaDfHwaB3DvxXcVFnWCROZscyGYQBH7CsRf9qcVzeI3tvZB9H
22uEStRldVVv+UIQkeCTYCFLXvCFFbiYBG8O5Z3gbgxFXRGaQX++GiurSUBWMtM5
PEhMHlp1jyiufqLRTTOMgfjA4FZzBgVEQl1nbPPW5lagCf9LI7Xy0rPFCaJZJZGK
L+5rlzQNQGUKJ+QVpOtw+eCK9CKF1QnBnGolHBm0Ft5TAFeXp/1CB/SIVBvPz2Ov
O14pCcHj54d1mbYxjWlM+b9t+Nl6mtYmxslfDX3luFSrfgknSpmknf5hkt4yA4qP
rqlekEqFNUtiV6lXdDfkeHSFTdqwGxlL9lTRXVu4sYGnehKrv/NgmbNcEesy2ALK
JCH7axcZe45ymDjsV+cYfA03z5v8NgW9kFPII7RQnnRBJperBLhqUu7O7zmf8D6X
84CJlf3pGrL91ol2mT9ELSyzmziNq0FhsV8JL+OWQIdnAAYE9r+hlGvQUsqNkN3r
v8HYin9bBb/txXPawo3fP0MVsRZ0MnQgs1vHJMB9QQQGYeS3umwex39o2NxnzTie
0xHyBAM21FJnyDIRt3sU0oTWjoaFyUBv9hKV9NAOW6i7vgMYkaQ/kqxJe8SHLqzQ
oTLeOYcz6v9KxGPy4N9D0Ot76YjsS5yRUiV0id720u/xKHI3aFsiG0hz9BQJ6nAc
L7Zw5bLy2pPq453YsI+7J5iHcZ4pQXxd3Zt24bto2WHSu1uDSJocl0BjHspdoln5
wkXveOT9HnZPD9CIXW1hZnZPdT9fTWJQifYkeTBHvrbiY3bnjayeIoQY89Lgs5H0
CamOu1l8yFKXHSpWOByEm8SCGb6HGXeR8MtLcSYHZs0n3IpmCLhUJXFfLoT1edbj
osZOSESu/p6ku1mQOak9V2kbwiS96NI+8UYmX8Cl9gio7vTWSrfzYFv2qJhx/Uor
FkfnoiXZESlt0Qx+ed0BEYiKY8NhJc3KYOEGaxUhSDNkLjxCH9Z0l2tDwDTqk2AG
cSPraCRctDtU12bBZxAele39wqu6UBFRONkW9S81MZyYkxCnP+/7nrSfbr+Undll
oKzHVCZ6TLEVuUxKJN7V2aEO/78s3oyZNCLs5zsDOBcBbCrvBqE7/YUfd+ITbUx0
42pH0FZJfCvee007JratASop9Oigjlxeh02cg9u3j2g4hVptKLvR7XSjrt5C40Tv
MFMu6jCNzyWbmXA9eQHvNnMVD2evkAv5giSgmBWQUqG5vZNtgF8XiddqGYRWw481
9mO8pi1hnAAWiSZwAeLr7iIDOYAzfwZI1HQKG1NuQrC8oS8FEwsRnBFTX0sLiXi2
jkfqqmHbBX5P3Vj5KUF+9KC+p5mX3PBmkifstwSREYP8Px4CRHKtlWa6FqYCQhCD
6BtnyKFK+hlEOXKOUK2G7jmFrTtvomTMdebb2dw0VYADBrLlC6h13S6A5YUV+VuV
buPFmu4C82tonlRSN/mC1rg/KYhvPV6fyIw6A+5T+PmYZv7aLH8KN2eRHPvSdaxn
ixxrCiay8D8f9j58eeA6IDvG+/Hb9ZRg8kgtgm5MLu2ZYVYeOSGCwJre0jSgI2zx
InfpbnO3BDz9x1IzNX7aPavlJikcmcd66qzIY/I5occTBaPmJemFll/ahozpZ43Y
jvKCVC3AI/066Pfx3FUmKYVL5cE9wGrELrQxDRTEqfL3i7/fG8mjlpjihl9O0135
Hso8K6MXiplYLS+O2mX8ZYgHz3xNTVucXKCAzllRSYEAZyauu90hVJcEaGKUVZej
exdlBe6qTGGmmFMBAJInBL9vzsQigg4uZYAVDazB54ZXd89qUshuAj9yP08WP3LK
oTL6Xg9nXqg9xVPaFvuJ6g==
`protect END_PROTECTED
