`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEPOcQuiKulPEU98PorznkMCwlWY/N4JqSbnJg0Ni6duHIYGB62auwWOkFMf1JLR
QEmG8KwgF3LjXnuqLJ5MUFjiQy1TDqc7OxyeM8iufjei2SNkPvvq2bks3bQ08/V0
u3FNxpl/WuiU6dQREBqckBsA4xRbkN1WikTJ9sn7q2VM/JfslBlB1Qi8U+wYXdbE
rccexDgV/IE10R8t9kO+/ADRYr0gPV3a3bmFQXGm1+U4Hah5oBtlIeDghpCnVVqZ
J42/0HFRRlwIXZxTPzQ6r0vo2P1Csr2KeYgB0ANKbvqLLeldV1k6eEX6FyqYtyqb
Tmg9Vy0WUxtMNQT9M35zkjS1PUImsLyU6TkcSjZI0uChHDQ2O4psaoq531qwNn7H
qK8EuZ4KqX8v0RfwnLDhkg==
`protect END_PROTECTED
