`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbDJuunfB0rinbirQz0DEviwo/Hj1Gyq/lRIre8LuOj4Ej8xo4gMGbmZiA0wguxl
ShmVG4DuEmialwZP5hpYb9Q+XEAXRDLeRhJJ+oySa6fVU54Cln5Oabtfm/wFSusK
mzC8yS6uKIlo7tXRZKAiRPjgw+QkEh+xnxGTaPyY6a0YvIRIZ0jpyQHAlcBPKk90
tpMDk4rPIMALxGdBgoffpIUPoou2eOi5L935uE7zHDNIIrGBj08zLUyF5UPVgriR
Tl6Boyx6JHqmP3+WqygcBQrc1JBf2K1O4aYPbIkSYwimS6ri81A804tMze2zJ5Qr
6F0tVUnxLqc1y6n71++GMzrq3N8rNeIeRDGVBMgorpAuDfQ5f80WAw1KhId/2hrx
bBL+maXRFdOr/YgeFohm8nrSStwVL/zOwL/YqUVBUlqaLF/O3B5vXaXAyM6itbYc
v4Lg/aDQhTGxyhiZe4d08kEWkb9n2O0q2MecswVTGJ15zITdvDiwJx2YJjWjyfRw
nbaKeRwnMdNRZlK3UjKJpYXueiOjpzr2zqkrQ2oWM5HMpVQUPi1jyXdAcMfH+qlt
YDqOgMZDeCEYQNWFdvv1ncOvUxyp+1GDpsg42Ko3guhjx8A+n1fE+kk5PGtQYnNW
MjSEYw0U3yiB/ER3lVWpOLyc+VnLVuScrM9n1OPk/BVvDTO4Wv+OfWaWjnO5NjER
d1UGdR+/OaeNpBvzlDyjbz/Gur12od2hhJXPULrqbJX7GGm1cdMCFb5LcZw9+kph
35dcuif2b8DjIsiM10fntJtGVGX2c1YSvOBZCTCKJreez1clQSEYGtOoxqYmLklZ
kfGQ1+pcEyui7M9nMDl9FUhDDBcw6gbzciK1epPiRoW+BQ7sXo3Cg1mA+PAv7fw/
Jzfe7QCg800nS1wRDg8sguaJU7b8w74LBxO80VjLLGH+oAYCrW1BBdyD6BM/xIks
7tFVvkdsJ3gelgG2nyQpHpkLfbQj0OGoAir8aZzmmZ7wilTSI1vNfeCNsuY7LL/x
8qnXbRxwy1vrqguCSTcTWGDW1w18kRrADJWOSkAwlJVhB5lbEOF7EWpOUiQUN0Sm
EmExpijU2rJKz7O10bkcvyyPq+ZXV4knpvOPhhIxZM8bFEwPMUKPnS5eNuhgZGZB
6D58tJOSwQyLDZq5E7Ovcbm74N46Bg7fIKlR9pQRQavgAczzfOckCotHdtBjouWZ
oczAby4m9iUEnyXNw00+b3TvYt2aD6bNEp5lpssFJDJUgUeSG3lNe10bMAGngWSV
nDp5nEPrPuoGFNu//BK9z2dy0d/9VfqKwVs56IZxw7is+FwTWIbJfrPgaQNlWfT/
a/zG6uTcrxVR/Hqlx6RAX19SlhqszSxsOPShNYHk6tLCwF4tRwBBhNtRuRSIkTtB
uKkmZTP/HOpp+5LI1ZePyaKhGt8nFsnb3mH5DWorsOhRvUhfg9O6tru3ZrX53eb3
3CqYY6ZlvVeM1wI6g23EVP8zCHeYdjuBDsZwNT5B0fcF+PexhxgO8gQmv2qcOz/x
tgQhNQRpfe+uUr/uOeUIn/6BsAx4ROw7TixDzdQaz8wHMCnnSPQMfk7v+9Pdnjek
dZDMYafDiDuNeVwdlubfitgWOYLPMt5n77XiO6yXJGkVzDSUUVkmG/JunMDCcs12
TCtDWy9qSbdJomsAqoaeHDr5UqSF0djg8JiCc0JJzpPCM5hv0rTNX+mG93NsNLFe
B8mQMF9wsTy5Y290fh7XNLz0MwLlijn/4rG0514KHa4GeIfiVwxqysBXpU2AMS6N
I/G/te16+F/XcSxr2rXKaQ1Ug2DiampqXHpwjrWPndvQpQ2XDLRcGc10cw/ldL0b
tqyv9EbyJ6zZNkY7VfDHlvgR3ilJDoNJ30dNMSMZUE3JOgV1hE/x/6FbUQB9x4lB
tZLGCwRtENPrAwYy9K06VHhFMoEuywj6nADoloWUT/3M7UrmQitF7fwRluizn1Pp
voGcFGUNNdAgKtcS5+Ad4sRSwV94L84n4MTe7jlFyceOvYJGV1RdgmBy+Ubkkrta
kROL4OXsX6HHRvXx6awDzSNfnloQxkbA+wmE2crKg7yjGNWqXjm/YlfeQGJQU+HO
vPGDWEEkZtXQVTZGFVuqd2GLNCgvGKpkj0veRiSTozVKysS037kIXGycQx2lA1sb
tkA8Sr7tyU4IAaPaV9IKbZZCXNw3+yZSK2+HLFnpE1pIarP4q0sIhzJwCyXpgbSb
rZRNSlbb+ByTYnUbck86EK736q/efnmTDNpN64XoRQCgLcvqFvC2ZCY+1MjDMqkq
jG4OWKtzCXZnPaQPHf7RFNVJI1xwSpIyN1Crt6AOPKkJlzsS2SkMB8YUYQsqpvXZ
Y4AuqLq5Q7xwIQ+hHF9KBAbTwR3Jef4qtVRgMQosKsbCrl6uTfGCVj9aIWH+EoNn
grGuc4e7cEy1Zn977b/KA016eKtaOWm3MSoSanu06BIK3hJ1+bakSBmUplntHwzg
JcxgyPHOmlTjWSzBMtrlRTkHUgr2Luhnoqdck8bcqZu3ne4juVdgLV3MA9v/8vt+
rinHX0ZKFlzarp70RNn5ZOsIZ98vMXL3MgbuCjmABt4+w3JDXRdLwR5a2Gw89+W/
j6Pu/22MKRawhaU6g17tORf0Mczl0mlQarhlYyEUzMS35hGoXLyZ26d9eh9RWL4/
2Z3ghIbKI4TitzyqwJz2qUPi+x7xxmipGKqlZ0u4m6eyFMQngtKawnG/4bIByo4p
PXw3pM0bJhW3EPSXlxyrseWhb7cKlak02VjIIfxzNcfIUlxrT2+oXpFUtDMxdxky
uJebZrw0eJzty+Jv6216ip9Mmr/40H+Q9Jw5+2T2omHu7tyr/HFZhg0h1I/XSSnc
wK8Mx9RNBZ+oMHUWMD3x2V94mYsTErq3F+GNJleMdaq20L/NF/fdRhSFMA9hfboy
`protect END_PROTECTED
