`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XkIkhHVm/q3m7M1QUHqttKl2y7lsdXSNLqL/dP0LLtJz5J6EW4hnwZapQWnPD98k
BgO2aUjILMwRn3BPTjL78/qEIPO6gUxQ+/hFpsSBbj09oQNVizoE7iwu2ExeqhR2
4ZLjq0XESg8enlrf5fz4Gj6zUY5gxjAUOK6ZgY5rTOzntC0bAq5Na2JzNIVIicyi
PMxakqDxOLdgFDTJuowd9JIZ+6pHHDsptee1N7WuDgP9NkuEWhiwc/KwvLSAT9mZ
49aqEjbD035xP9q7fLl8ndFAbDl6Rr2+5MBHZ1geEmmLN2cuXMxW295yzTssw2kv
bJFyA4xYZOeG1HVyBj3KLRdCpDW2lx7MJBMx2MXMSN8lWOXch3k3rDPEb9mOgBrf
YWbj5MTJJia9eNCKzTRb1Q==
`protect END_PROTECTED
