`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djmWl6HmTXUf1FSNmLShG4OBHKWxt+fXSMpUm26zyOIYBiPz7a6qKZEO3Ff2RJ4B
R4uEHCXXtp5x5nYlFXz0p+qDs8EC1DcVGHlNjFjtA+JqEOXlXWfKY+R7jb0D1q29
9XtLCcZWoTas30xqdSWsGHrMXZeOLxAAEUwIMvIfTvM7hhUGRiPY5p8T1MV4336o
mVcm5PMIfh8tpLL8s3qcgFAIDpiUY+mlJZJt13U5EnmUC87OE8Rjvr3GTJhHCIrm
IC9NHZOOGsgakdDJmoZj4epQf77HydaLtY/F1HB+wS10al8lONgo/SVn4s5kGDal
RVFFQ1QiDI41oYScgG1WlEM4ceSSdQz+j0uR3OoJbgyF1tzZOny424kgqagFLjTN
GaUIelIKP9n15q7ASsUOzjPSOPuqbhlDTLB10VWSEw9s8xKH8TzN3Kvy7kTXlOkL
/MwtYAmDPofdv9iZXtvItL8RpsbeembxJozCqpv0WFiiZbzra6ZBXaDoXTraBLBd
qfdJPG8zEuIcaNaQIcEGTAGZIxAD7MCP4Oq1UhYVIBNH4GMVH+Zlm1Ll1lgCpBBL
ftuVprhBIfIoo/kr6lsnYfRrRExO9jLr3mVi9cYMoUo6vdYofqpriSAmjNcU4Heo
fWRw3QWUSOF7XiRi2ixPUpusvePaATwKasN7EqhgmrMRg+q9hZoObsxMdZ1RnUtQ
`protect END_PROTECTED
