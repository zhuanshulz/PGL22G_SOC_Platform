`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XVC02LjV2N/Qz0GEWtPHfyG7VOH8PFgpt0X433n9OtBoo14tSd1yfT3QTWWSnjY
v8t0v5pP6xm0ULfUhirTV3zR/kpvVOdm922JIymySSVFw4BS8I6a1MxZZzt7r5T0
up1C93fGAaw9svDLkaws/NX/T/KhXCW/gOIVIm6ZGn3hI0lmAh9cBlkCKiEjE1vq
nqpOlq4E8K1ziobCxsp7/+9u40NUTTZ3uXQvS5LWpI2RPoLN04j8QsQTsIekK8Ry
IixRDSYRAiwBIyRGLOZrEIgWbHbmsZzZ2MEiUEWKfrUgK1r/tB8kp7N6VX3leI4P
G36nytW++BOYNecwmXTfzX0aFm3OyXoVO6MT8OdFnumbX+TQmI3BgvLVdQhxaES0
j4Lk0mt1nszQ1Pp8CUi1NMUcE2emWW+p6ekT7UCh4PYod9QdH0/hgt+FGQLCWU9L
TaH013YdE1mfZpDJ2IbVKp2+JTY8MQsD6k7kYTRlZh5+6ZeEq5BkrZu6J3qJkJN8
+cacB7i3GowIUDeVcTuUQ2A9rmbCutq8Sj7aG+ns37n7m7G08L4h7vYotU7gA+ex
7Npmnt7Bcl10mhiBcs6POiZIEH1AqmP33lKxXlwdyn9QEe1Ckh0MJ8aB1GM/6v5J
1sUC9h+R3duZchA4VfxxFobFlAcAYst4royLFZDFoaZWd/tgJe/3cDuYyV1GgLhH
kKjxF8cRtR7q0969Xha6Yn61Q99b9IWCK7I/Rw3lRvAYpquNkMzZ5halHzFskFQY
QjIj64wpt3lnhgZWcFoql4derX7QAbHqfx3IBUcCIAsHGV5hhclWyH/xdOQDlgqv
HOkL5XWNW6Tw2DoiPVlcMfblRYXUQzYZfZe1dPjC/yZsO4EQKbkDgHMHv7mFUGoH
F0ykRNX9LUNCJhNz/KOL/haU+wAoUdEzQ5U3FqRbXq5vV9VFpqoaFcVMlq63FJls
XnC+S7ad5TS8uZEFmwDVqUKmjxSM4z7ogeVMLlFndlABQzkOS4Pe67jEBVavSvn5
eeNyJxmWFUJsr/458qUvMpLq+wMFMZxJUiqbPz5hPlWKzYIu1oB0Q50uDd7TuuFa
y19A0cNcTHp2xJEXflhAkm9IJbGUOn45gJk2i2H/WjxoYeAy9ItaHueNdVKwCi3y
OwUu67gknQPH1W8jCeW91zIXETx9asFgBywQfsnDXwwwb66lk52kYmLCoa4KnPiE
yCVlhMVyK5aNyVdAZXHuM7cZ+VbhZ5M8M4ymTHcYFxs4H+76rRiYBH72o/DV2Rp6
I+IKcZ/Z4Qn9kUpCJlpq98wWIrEKwZ4lh6TdUr6UEg/Audjsb0GSBEi15XEiCHbp
7HR+MAmDBzMZ9D0wLarlVLRA915VoEVNX5dsZEUMvBpKZ2yAhri8AIS61xWvutU0
/LSd9Aq5bTpmuQieBEKXViNHi9hrQf5T0weIwQodIcd5wYoglq3q3ebZExotJsHw
EeF1GpsnfBpW+44+O8hv5rCmb4p8ElVj7WOTT1pKJSi9A6zVvCoT4zzBFAl2P3fV
Yq8B009gUG4Ta7ST/W9xNFVQqr/lhMPabtIXNOy/wG09vncNtHXapipoMXh2/PK/
qwK3idXoMdEsA0DyBs+KhJx9ZM81LobAb0gnO3NOTkk3jlm1hMMITsjFwU3fahVc
hR1UnCtkJQVDchaXlZ+dHw2PDcUVxd66w+MzNNzM2aIFBA4dsjrfg0zrAhg11SlG
Va9k/nNgMGUFkqpT32geuurQkajV0dokhVx1HPjcVzv8I/Ain0wyaklbQ+MshDS1
/MA+Cv9NafrPfM92GqhPIEy6hzruZghxyPafHFX/K6ic2hdg0+5a8a0fVMg1OEdN
PPBdpSV4ECGzUEch4Uw/yI1Gi+gCBe4XlMjQ/mrNfT6WnXWiEQswLneFlj4z+Ws0
doGFc9AqLrpwk04ppqaafxlhp041SDBl3n05uwIY0JPeIXw6OcG9b7V9uxRbK8Ap
dA/9nYaZE2BH8fFxGCBHdNjgriTBlgpjrydcM9I6V1ogTIgKSw3UtJ8/g/6HY3Y6
6RrKdi/RvTFreuR/+yEH6QFQx55MvjVjHeG8ltDPRujBnfDUfg03T7aRbANJrekv
DGoNi0kVeyozxyAv/ZoEa5yJ2E/r7gxpfZvO3M/Ri8aZBs0GSF9/ffTtntoBFoPx
WUqOYbmaS3qm58+yTR+G6IF5rvOJU/pbRrPtemqPw+slAIweMEnGp/3jsbxwQICg
HjsZHH7m0VFT38WDwkTNStHw/bI7cFVbLfn6Hy/DwzU370F5Ju9CZPphC6ZpVU+w
LNI/SetZOywdLa2fROdUYZbFYOZHH6wWKtUjXNd2D1zBqk6DtMVaOKDAVVktB+kk
uqZf7NiPtzQA6IA73Oqn1OvdRTtQHUptWol2g5djdRO1caVGKt0YD8JAj6oS+Qpy
NZ94ziKLacd3xhe4h+TGHo46O7v/J4kN6diynkE8lFVY0aWxiomsmQYvhJo2g2he
Ca3RTKB2FD5Z/qoicJ6WzIJUBBvUBICXbjYVUj0a14258cF1bmNwCVLw+1fl61VA
rCTZtfXkTggwm8jnvQ1JSpLqR52DciAHpvB7tp4pqkG8dokaXahm6Nmz2cYMg/SX
agB0pXHxgGKHdOpzXhfoNYJtuHiPSqlYeaNyta16Q7LbthL6Le5/8OYSnX9LHFAm
bVjMSArxxbGN9aAbFW2Wh5HjLcsXKYXHKLtqU1jBtkpd4zRrsmvatA0k+VTFgu5X
Mrc95FiSRPSNtEjYKa3fmtYMAl6yo4n/RoDX8lv80f448gAWtLECtCZyHmFoVxoH
J+qLtwagNb0ko2hImVCrqwILhPsTn1W7whEIyglRdVun8Ss/xyc/PCt8fy/PYNOo
7mnXXeRtdC3oOzIHN/XQnWCKhyQrIGjvieufI5Gn1x0Ve7ubK+0nBQIh+fCR00nv
agKW7noYM9u+Opor71T3/x8eRxpHf8x76+KNsL5RVuSimQaGEBehUTHLsKo0YI0W
hFRo2h0LAyiWMC5nu7KqA9aatK/yGlpsF+v24+rxvtFMez9UeZslnIUFM1bgu03G
3blJ+53itA4N8wYru/JpM554AhziSKqG+/qK24giFAoXHeFmN1rlhdZRBs5DC7QI
1I9dT7CKkYGO4diCwgvacSG30QhAVfRGUMvvoNEBC/pWsnzkz44lccdtG4xJtNAq
5FztLJedQrh/0tR+Ugcp1/gHp73XWU4GIQsQHNlsOvrYJZS/HkqgTYPhvYwWKPP0
fHQ19hD9Nbb2Po+7c3HJAS+1Lakw65ik/9xADzKSS8naSiHDnPkfDbCm/E+oZh6W
m+8scTCCbbuRoc9PgCj3cWK0wyZTaHpXWJDsODTzJYESTzdOPOk6KPkhc9ei7Zsa
0K3KeF8J+3tdqlRHMIJlmv8mNL/oyOHeCmjJoScqJ3PH5aYk/jbSJSXF+Q0QoHg/
8yeUsGlyDAe58V+NnHo+kjX/t5YKcx9e/qTZoU+zmHJKCoKhjyP8loO08Aa6xuZO
GFUmwZzV/EyUvgt7Qga300sfK6yucwi9MkwX4TSzaTVC7wT9/gdbVox8sIL4psUR
++4jvwzCx8SYoIL1Mbzp3q0uZql5jpWzxsihcrQwl3yN6Sv37qRV2/Xn6R1pENWR
AdswawGEOub46OJmrGiM2p2pq2yG51QOm8dBuKvtBit4oo8j3vqLOSWLjz1shJYL
eEM1s2pPcXWf8ikVA2zQuybWpOfY0ias1TI0gwHCoMI7cJxYcINFWHpqOpV0e4t1
EZJ78H+mxRwu3BaDgci9HkiTUyIISuktSzLOqYMTdqq33q24pXiK0qHXSqw34gvX
DB8IwS8ArwVHvRgwO7LJROD3039frIEODPbMbCS2MUDQYl6LYgjLXTAhci7zbqhx
Y+jFtSNbdgLywFBCDcuIEBLXSwvzIxA2gXQj/OJO8BWKy2Wdfday7qoIW0xbuuiU
cluxr2+0gzDjXkhoHX/h31A8k/Z511+w8shNOjngCU/mruyncl5UuGknXbiM+gJ3
mX13kkBaELm6iNIPdYC2iqzEMvMLOi2YMVsx6AnBD0+sy24qh9ClSJE9nrtCFTn0
iqLY81l8IW4lwbWgaZySrumwBTy3sb6ey0PqG7yAP73ArZjX52IXWRhRDelhwu/a
AWdrQ9NmTmRoHR21r2NhH/hRDGzV5OT+N3NkDQsu/gc+88aD8wpCMTjenjGEd7Wj
9/1ypPqurZWQjjk6qnM9gU9eTnNmolCqy8wSJaDvnazevxnJjwaXBh9Zg/wNDF6y
RDMi5BOdYbXScztOrX+Tjr9vouyJk5B3McVAYksAukC0SatC4dBdhSwFxQBx6gAR
Y48ISjmETdlej3WKb1PrnLD6SonHYP8KLIJSgGLersmwGx4gJwr8XKP56hOZ4Pcn
ADggYux8NI0h/64VQDPkQfCQLM47aHGfUcjXQoGyKpei7bRI3CnkhMnGlJHIRlBK
Cn7UhvRDVoxIKZO1se1LHI9vHv4ctAchV27IhhvmN8ehFHL3QjdUn7etsp9nZir2
86hsrUf+YRNA8Lo8OHgkpI27hjFqJQaHBpsV54WIo1VrNyOCH2apNraT3GBTqBx0
fgPeO+VRscJzIzNelvCV1kzkqwTYodk4wbqbgg6ssTTBcRXVGqkaXg8rIvEWynyC
KO/vcG/Vc0DuEE4UO+IhuRYpBToB9CqkwURw0Rzx7LOdkwWCxKjbyuoPaSwtvIIg
gG7O3hzVCmxUwgDdSGI03ZTNrsEmS70N2jFV1Q42ZUJ0BXJqlgN8me1WKQuzezc7
VmWYBnhz66JUu50DuBOys7CH2lNr4uvYYM1xFN+RAuEFd9lFo/vylybGAOwdXeds
+1A9mPGS0BtEfoM9MgpZReLx6L/HY9zgefGzjXYrnrgh+EFvR1jbM9JPPlgrLJsH
IGpz9HzB/qFueP+TIuPbp36vHUNumtNzzsT/+S6QAcIc4kDe93nk1wkpZlusgXoZ
BO0mhHVj1M7VeG6qUqR26Dycrimn5EokdrBvln4Op5jGcUptbyMQhL7lT8LdJ70i
m47WfCEWllMeZlcAi2GTeHbfuUBHvAFESRKb/TkohsROgsWasjZ/z3ggbnf1rKY+
txsKAJK+DsmybsSIbC7jWAMQte7p56kK/fXQ6gyovrDFPXr90zCIS7evCSLVLsVi
TQL446qma1+cVMmiOWKgui5BzN8FuqfmV88INkTJg9xj+U9OxPZvRJHDH7iBSSSM
s1K0RY/KYtzOEHvjiIna4/iEONlTDl1My0fUn7lafuKVkPZYnKbkmlQYtqFBrW0d
ekD2QEkn7nEiX8f2WdbwyOd/x+Lp+4eel3SriQYF4pajSs53PZMsA1Y6SpfvW42S
je9epB71D3yUf4O3kl+O7AH3ZY7soZxz4gKyw+wgGIgX7e08nHxA749VqxLX/iXK
hjVHqB657xCCo/2YEUW2SQ8Biu6U1urQSr7h+KskrEjCyTZyjBY5OqZTSgijGGnz
pMn7C0Aqx1d77XvShKKzgwGXtRoU11axfqKDrcGAg5hc4NKLJ/YbRYYHu0Y8FI83
uQIEb/JVDD4g5mKM+3lpcj6PaS6XaxlfhC7+/oE3VaAIjaroEQtehzinlsiggQLj
04Jy2T30kB7tDOoyQEZWV5M9ptfy9xpu7vrWz6Z1X59sv3wqNBd9jHqi4tZC5baU
jT9oFfEGgrDLF+IbvxPZYYKFASvoPSX7A4sR7lm1nRLNfZCwbkXmng4rJpZgpYWo
MAtD1F5lSkrkYGOsY2WYXxGks6TXzRfUSiiCaQicbltUrvO1yEyIZ7Ku8NPBaQcY
L9iCrjjSld34wdAY1mpbBV8js2m+qNbYfLb+TnVPI/00VBe5u1/cTH75TBR+uaFH
lG8UumxFgQXd+20qI3pgWe+QpABGP6kaNYmUB8ww0Y+2PdHw7R9aBwGAwoWOovgH
lpaUCTjoEdOuimLau3jaRtC+QNU7MbG9E7IA2yt8dxXuLMMn9TsTg0zsEhJhr8xH
gIs0ZZ1wDyahx8VaUykgWQlvj3pEjUzxr0VC/NEXNjhg0AM+zt9GQ+tNQuQh+3BO
wR6Uzdg4GJmd2mbJJsXBZTwCq30fJ/iUXPpMxVVKpMZYcdyaNbfUNJ5VG1NxaOXq
KkNauL3LuqgeCxx9+GjWwNLmL++MQZBVL8PNob0Q90sV+yXEvj9KhnLjf+V3nvBd
Fj4Nr/zk9CRhup7jxi3RzQDD4Cs5AAQkz4Gy06/lm9dtICrkEh48fS9HQkwD8ZzE
qfXj/1j/s9rQVgC3a6NrhDP+tzRam17fh3L4sBFZjug4cCtTpN58ueMLhwxFYrXv
0lWbEVL2gapAOJZgjZ+GcRL4K5NvVks1t5KceeunsCQVXhKgsvr3saA9Z4kfENtL
8JEtz+tVPYp+2KkBt+u625UMjxuuO13hXMZcpHzfT5/OrFwY4RAj8KM/xGPLxW3A
lnzfuhnipghoLbOABP7FVfKsbhMlQfDAKu5BqrEwP7cAVzixmeMh88f1L7Zhz5mH
MI5reyq78sIZHOPheg3XJf3T9CzW42TSrCqP76H5tgkp1v7ydODQ8PyNcwOCU7pL
TKkqFK7ArXL8mDu1xhJ6yaapKYBxGrU+9FKBLWK6n8kC6lkD7GgDqM8A27Pgq727
MdX1S5qoYWWmQMhfAOq3urXCVTHtwpL7cNUuh3ErCIJDC9psPAVvz1DcgVFVbpRZ
EcDzcbwb+L2pn5mHYE1aBf0+uHf0XveXnAJ3QH+clUjrBBpEwos3X2fyM8uWJS9v
wJ3nSf/U9K3AESdTUj+27v7GN1Ols24Qat8u2i0HBZVf4Ge/CDr+/cSXZUzzSAFy
6/RMLIWQhRjb5Ju9FkVK8mcO0Cg6xanzWwgO6biKJo+EbYcWYTc09rT5yPnl0gkL
9VpSWurZTPm66FmyNQTv9lcxsRLNz2c0eS25H9B+f0ty5RSQBk8Mxv9j8gLQ7D71
KO43kVZ26pQxv9VgyyYRSNAwIv9GRzIENmm43ZdFkYY3LQQ2LZwEPvi+FAvL6ktL
9Tr2JeHb9foLJW+Avnpuu0Sizh+4Wrj2RVZXmlujK/zR31A2RstIhvKIDou6SrDm
Ol3Ld37cQBIbFaZO2xWBvpzE+JAXQ4YejbINGBosa663D2rD4CZ6VgBPjCD4egbB
WdHxE94jGCVSZWvBK6PW91p6dRYHbalxB7O0NKTy7u71N+DX5MAZwwod4oNsf6w6
VfvAZhMQIdW1OtGUwnlFnizlxeNfOi1fCTkPndVhEyiK/U5UE0F4oqG0tnU+1EsR
CRqrl8Il6/rSLox5fyMu72gkjfClLGLrEzNo6LgT1wz2iwY9J2Snbi+5TVTG1lsL
n9WFs7rAmXtyJQOn6jhiDaee5Zz5ZLoYmSjbllYOhBM8m22JWc1a+xQNrOKnYHym
Rct0QHQJ+KfBwKG4pKneI5/Ut1GPER3HIoxjI0t2KPKyrun0sCQPQUp3DoasWmFK
53jIsBTQJF2vt0dlajj7DcIYusXoJdTfTB7o/Wcarw+zZYz0cHGTQ5JoxTQ2QaRx
bslbsfIHa30NbCJ06cG59KDHlmtG5P9ql3bo8YaeEG2Ep0ziIiTkriNcrwFjvTSw
3RHKjst0AmzQB8hNp4Nf4EadkKFFIniuthuwOIg7TRfq+IzeQE4//nJbUDsFE/aX
WI/R/fWDo1H5zH+ssqaXgixrmUmC0gn/ADBpdiNI44wWuMvetWk/aAG5NoCruREi
nC+46EVdlRe/YzftfgP0E8CYs0Fbj2fl06n8KtFe8YGmLKcRNWlHINYqoKMuKPnP
eBjxF3yHOy8aKv4r8LjiyBxC0uzFoQkTcrIfZSkAe0P/4js5QJ26ikBi2pvx1IUw
ZzgKWe7mq3pzTYxA16bDS9yuMV3tK/xyiot2LMw59ylwbpWQeJp24N8tkSpYxKGE
jhxqqBlgFgiQxDJ7haVikks7eJ6I6tJ/YjUF9Dwz23xAOABjHJ8stxcVwPwTpsPL
OjO7WRNmCug5Ds4m7ctdTVymRX14Awg49i3DDzjwHGS2dVxLzjwGW2TI4oburULA
0CNVmZvoF1Pwf48nM2x1DZ3tYpSlEJxFNxvQwf4KUMDYibD0aYubo2zwF8/AgPub
CJItI+HpLM1qEv91AvjTamOtXovUTCeo9CjKfSHUID+2JTiz6m8kvHHua2skgKMa
Sl9Gt+g4WM4yZkeaXWFqA7MWl3hmZRaKg20ituf5yYl+4eYhAB0dpDsdG6i57W1l
iZOJkKslaav61ZMhsCet0ivgnyaWcfEUXfOw3qRBsDMNc4X1gTRYGIimTQKFDxjF
JgLpZp0JGnnKdjnXVta7fXRFdRjQ4mpsBDN34t5D1dDppebsEoEpneY0EwhTh45v
9YX2jVgTdURFMyAsaHKHhA1qKS4hSLx21BTVYlzKKT1zmcnd3QPiX1wXU7KtsG75
RALDfI0Kj3tYbZaVtwVgvPItQoPKAhQrxE4jHsEhrAhrgH8+FZ03Pk3CrrSTqX78
p02b6EEMnyomiI4UQVpVvTg2ysWlY9M/FztWL5hmtICE+9c7ZsBbCxyLrOL9y/jV
CSNGtdNhWyKBGy/siDOSdFhzvbKyJviEPZpWzDU5nKb7N5GyUj1e30K0L1mpBYOT
PYRB3c5V8V83byw4eVPOfSYOcnAMezxM3hwIqgR7jNMfYrlPqR4uxmWMZGUx5vu0
bY7kGdsyelqfaL+UBm7ckhJsFlGmNqds4rIEQfhz1NVEJ6oAaDdFwVN2mjgJXeht
/f22TgxKdRuKf75HQW9AlbvfAd3nXKFKuUSFvNMPkzMzwGc0YxfXnPhObtUnYdXH
lTEWR0OEO1UpVnEndziLpiQldWPT9npspsnuiKrWaywtXlSYlTGl6WmeD+kJOt+4
OBprUeRZgYOt2EtEU7+G2qoxU2e9HFE+wEMvgrglMfoKPW0y6n8W4/LgAyC0VliV
bL9fkNVA+TnLR/f5e8gzjvy7MPtAnp3M2uj+BA/lh4Wak8FnI795vwCcqjHrFobo
y0/03/CbUQsKsgWMD/KU2yY4LxuxvVHP5+wscIZCfNdAFb7GRCVlXje38lzEXkE1
uonEO9DXynUndCxEc+zT8/p8JpE858mAOlNDGOGa6cJ+EQgsTjDzXwu79FOEQS1L
liR6FxYfYgwKVlnfiRkMT7s5Ugz35YLaR9DSiO3ldBjhTTe4O1xVEahXKeo0DLyM
zyZ38tG/1JbbXKhLMtQG7/8rFWSsrnSaksZBaQls5uSO2CNLPl4XXbJQ3hI3dIJ2
WmyHVEvhJeI/68dL5HB1SJEvAaOtcAryJjw01UUa0OemoVLNxR6loS+YnFJ0OI/y
f011v1SWciLATF4Gdv584w+04zktkqkBUzHokr0aVL4CmlPgvP1jKp3to/YyzSb2
WDWbu5FMJQwE+NmeB80UH9GKwGmXh3EgRgIos99VTDcrzLU2LMVRu95N3ScN9A7y
T50OYJoVzCYtVzpDaNASRMNKwAFr6OVIuEjDFbCSdYO9BQ+8KoPXWB7pRYdUaOec
zE+0u53S4OSPNZLCbW5JHdnxLGN2dQqaWthJCr2NjndtdlLeGnWPRi/tIIfptsC2
QmZSdvp53lp+qyfVlV4V5e9eLI64NYyAyy1nw5/dN78z8nRxZsf2C+Ded5d50SMK
55bamchMIn5hLkFMt+yEZeOb/7MWAopMKVKqI2AXQyWO0lXvGLGM/SIMtvJLYlTP
xNJ+UMei7kaE2UAHV6xo4ZkZuJr23jpMqA0I/+slUoeLqmekLi7rAiW8KSDOPjNm
EbtKppL11NHgVw1OZGGK4E6biS8XWJxb7en/p0I7tE0StYA5kRUQvJmfW7MMuCQ4
ywLJc1y8H9t1tydoQK3iS6j0ZtWFsRAoGthN4CsvGO1ZqtTHqKZBkhaGu2Vu6UQx
pShrDp+sd/qow5kr2G/0incA0EZweirqFCMlH4yRwIkRPxE3k6liTctCIk45mRyy
0DIdkmsE//GiLKSmn0owFaQG+nEIcbmRICbttpbpT5wdnkFOmWBpFuSmTHtgdvbP
ARSSF6xmn9ZihHDWMXPaR1vNTRaV5iL5wBA+gAt3l+NKn45ddTjGJ7OCXCInOsCK
mpm3LOfNEe2Uz5M4t/eOJ+dme/c7xJVw8QUki8wl8XiFSN8BCKp14AkhjyTNF+L4
gxFJxyNBfg5ErmsszoVV78Lq+JN87ecSwosKHqTQ0zbDtQ5ZiDGysEbAHTvPFXCD
dXMkQyUACaQSk11Fa4z9Yt+4bE3cBvelc1VXr60o7cJcl2EAEeUgxJ8CoXYqPcI8
C+RX0d0JchOdlgj+K8nJTt+4izr+YRsGYywQyVL72eTtJjRVBAE1vqAVcJ3lGTpA
gIw7JFpW7emamxzRp9XQm4amZVSWKWmNOvqKuRaLk6ytDuPPf4dMIY1XWsvTUGeS
KBKCPVEASU3UPT2GeM4n/yF3zkF4Bw6NUSorsa0r2MLk+vutG7Ohgyq+iZGaPbLx
Nh+1Bt0S+Xqsg0nlLirL0pysXbBbLUDNJPnKpkTLkd/tbo0WUiwOrIGL+PXglzgC
LYPTgljwrULGxdYyM0a51NLnMZ0ubQrm59LSSSh10qiLx49+1yaNh1S11laBkXe/
6IsDB/BqzP+yHlf7diDFv5r1QB12DTZggRcaLbN4bpP8SbEvgLkT87LyVa3zgDXm
SDQrKFQ0V2hsQAkHt79w4i65IZDKtEqZQzCIMwTknZlpBy/hl+6TPL7eUO1JeZgy
8Bcgs1r07DrLxRD0ZI93/chcYwGVzCRfRWvj8wdyJPJ7qstYFBHFrqo5ZuamRBG4
G4MyS1U3SvmraFk5dkPUba+gAwBISfRSmeUIt7yA8I/xLo7dmt16OvjN28N922Xe
9mN2L6jxseYA5nt0JMrRXIovH7QjsVqG3KklWbK6edR+8zedfOME3XwDOUpWbpVr
zxrJkmy5FqruHpgQq0CwE5bQSfBSXK81BpsWMooHBIvTYDPqTS0Uzr8JZHa5IFve
1hGqpEqi7xU6SGIw3w+k2AXmfRp+0v6nnPjggipLJnlVufQ9iS2p5A/z4zYupYqz
4rxHooT8UmYoEgLAl+xfbdlNOWRcEPIDhrxR5nnXmG9MHOF4EIPQHgQi2AGcJPnX
VMQFDiHdv8bkkiISlQU3AyExrDjNSjBspuq+MdaGMaUtHLqjWlqdjRoofhI0ukj/
cpwJnursMs+4f4lwfqnj01/t+DRDtmGCLaOi6QEsdWTtQypqv6REMrqixXYmug/t
+j9nXgQh2I3ngC0eFCoIQsTYk4sKcoY5XM8kOQN6mq4I0XZPLbFEc0AKyfhklx8t
9R1n7bwgLPkxadd9XXhdZTOyagi3lZ6PIAps8f265L0B7Dla+KtT2q7IjyKepaPh
w+zlVIFeHQDh73pEiDVe5cdDEiRMKFfHMa9sikQ1LKw+sy5VL2775YP/SCajd0mF
cl7PyqbFuGrAJFt3HvBESKWUpdNyvsDFRRGBO6SE0r6LRjqMUU7wOhnown6F8d/p
R1XCCH0cMz15v7jeVd/fb9oYSD5Sagmxqta7vi+3rr92R6BVn22KPWXst+ujQLa5
Ma1DMkdoRstVKpPOYVKDTntLty02CuYlmK/AuO4gDaSuDS9eD6GOcin3wuXJZOTb
UtY7qi16mlzi1AoeAJszd5mhSfHzrScBCT3irL3rHpZQeRKb246Yz3qqJJ4yHulg
FjT1pt761/CC8IE4NXKP4D96mhW9PYT3GlMNYCfzeei97Rydv5qrOIrwNJQo/BeU
fO3KG/4t1QAcMEornFZMQhIpwDK4fLh5JzLKu1hIoweUIbDTZnNZVc19dVpq+vLc
DFDmoYO4MisPAYZwahrMyoLfgZ4dFEoMkvK/WPwYQirHfI3sQwsOKEnhX2o0Ltlx
zLHry4j2dW4sTiA5mx5u9MEWW/NamCuThT9g35AzlUZaxkTFgbDdqGA7yPDv1m0U
qtrStflycipToXihA2qvAHwYnXDTUy7WJA6lCvq7Z+cg2ytcNzWJnc+LOnnbXaPr
oc5kcc5AsPzKsrIQ8DINtA6YQMw7U4NYGFXtrR7pUQ5+2VGcgvmu5nCcNySxMARt
bN1RYfsCU6bxisgLNNQROoUciY95E14e1L2mb4jeEA6pnwpCj3v22dLb0GfzSNYJ
c4wgmRa7oJm5rfkuAQPJFWXZqkyNoXhNj7wbPD7+V3YMWqlAl7lGIUXqEYzGK3iM
Th95GYi1Brwy1z+xtJWbJ5FliEX85HeLjKnuPnx7EfFAiUEwMtqfA8jn2LPyjOV6
6ztW7GdYKSLO0tL8886XHMEbO/v+wV14RZKZoZAr1vXljS2N+nHUxV95cSmfNlkg
OZ79qIpRilu9N5QwdxsNGQ+0onCat4DumDCBtUwMQZJDjAOr1GkMsF9V4EBn6JcP
nmoYp2tDrdM5cbfcxYw3j9Es9Z9i0Oy24TLdouW6XW6IC3lmYz04sLGlQGZFOI0e
7g5oMJu2Niujs2wub9GoGvxKVH7ooD+yev1aGRhYzJEsbHx+AL69G1c2koni9TxC
M9OFpRSlomkU5pJWjRui6g7OmMh4gW82t0GEsixqp4S6Wduyz0+WSYapwxiw3yI2
ZFH6twMWhgp7RNqDcv5sqKHUOLipSpVxw9TRJUlrwiOfE++FiW/V/GGRbZ5C0iEz
sEW+FXXldQNGKR/kG80sBHEbgTdo93yb2NLHfynbxmplmt7H0FyvSafHHY3+/jOj
a7fmBADc8B2TkINHxFChNOsmi0HP4eRLTcebAKNJYm03c1kXHWB5MG2jLhheFEJd
SqiqXo8ugmApJOFb1mGfx2G6y4YWh86ABOQNSw3e/BD3pVrEyAdLVlhQm0ansHZJ
ShfvSwFz+mw2A52yUMBOqTDy1DbekxPkQOp4bdBaEligxKi/1bUNRipLNMQeVrKN
6NuWGg5/P1Qh6ZmdDxZIK1hA7l5Kn207byf7HLPkdIhXXLQQ0aeXb2i1nhMrmrfz
rBmM29vNoRG2UTIG9cQxe+WDz11w4TDixJ4k6m18DYoCfZZKAasel0GOzr5BC6wu
UCPmTGzxdA02KoK5UylWD4Nrfc9zSNtJwdNvJ/D4Hn06z0NKHUBdPXFlW9mcd8RM
RYm6z11AgyyczHUzXrk0MmTFWEiQX/5DYrBy7CY4urzzajj+HBbygt6dI/9+rRNn
6LaSN9zOgP6YdICeoHRVJwpdkd4Fjuejfr4WdSV8VLJ44+QqZn+mHD4hmFAchiXe
1yiAycoUwJ6yA+uLKS8fcKGge7BBujdINdHns3g3g3bhZ3YWRpzAr7OAk9/yZaSD
XM5Q25b7RI4G4GBxRHB2oWZ9iKA5/YbfcPSrLwVFh7Xh6E2tTDHorSuRz8P8Cr4h
KlHW3h8EEKvumr245BVT5DRQPvhsK7iIN6UQN2X6iX10MJheJHs/Yk/SFWoFX3/r
gRBqHaor/rsKFFMqNzJiEHmoxB2MB0uLT99HwBuIr2sjtxM0C8/elMevCS/HjANm
0wgTfAVD+KKQj27dTOohFuWwoNQYKzwx+W2VgenNSH2/a9fYLYDdDOiKUTznUGcv
VedS/pWzsaS0neubMAg0aX/Q1HdNXI5eeulTUIBAWQ6pd2KECexBUmgGQgd2dN9q
JFs45Hg3g7ZIVZabxG2v8dnI90PGAaj+WDKQxxzVMKKVQwVZpj2FCgZqH0McwisE
v7IWuP7OgLoD98xP+VsOHfXDWcTBbCq9ioJBFZV8d0QJMwRbU8xoj8PvChwgQXw6
4goeYF9w0FGMoc7C0PxrzqZ30VtvzOeVyjk/fno7SP6Sb87v9IewRDpGdy+DXnFi
cQFlxu7c6uq5dYpnhnAVm0dKiCutWJVNR+2pAs2rftApd5tElHbbmLHV2rvlfC2H
m2tDNCJ+vFNXDd8/Elss1mIT+cKuni6T3k1qu9WhJ8VYw+Gk7aQC4fA2POVPFjYO
2QU6uTNCiFi67H28nzRFR0wwpXqMyrEcj/U4QZOspDf1XLVlpHRmK0LmzpvAub/i
ooKI3v4tFFRf8lfv3qPXXBNmYpUGGmz6kHLGGhjHwMeV5971NrE/XDPZD//im5A8
khOAwjvciO3Wkv8GwMtjEX3f2xA4dRRl37ZqqVj2qpM0zw6JShAkbDj8KHyzeccs
w7QIqkmtfjFCpRIdKVfWP//18bUq1tvTZ+Ooc9eelDGMnMURBlytDQ/i+kAqwgve
xyhBXsvbFO6yLi6NqOMgHg9y0c9nettou97mJM/GdYQQAm6B2tZUiR9JSRCeTBjV
Mri5yx4A+u1H9pHm1PMWx3WC9qH2V/b9bpJawadSNrM/rJ0hGaSWwC7onH3MJ6sm
DLcSezpzXELjPOWbHfWCz524+0QhJTg3cMYA9ZOg0X01VNhJTdsxw+ASlq6VPkzg
WhYF9LPFSlpSDenN19SZWxopLE7xyc9uhcWW7kHjASjVUbjWkVw+TsuwodI/q806
1SGFhUePSo7ZdSwjH7ezJbmBkxhqsLU7fJlGm1CTO7ZXrZkk3KAI4jiVfsiaT9u/
wVbu1eWDQe0hEFcM/6IfE1WtswhRibWKnWn0C4PAt2bZ1U1/N/FBu79Kzw8LvTHU
AkitpUTZ0r/R64DAdwB388B5VZThXFwNHBVuy5iiYgFT849nLs1x206OKgl/uRYP
OvGaGRHgjwFzPvMt8nwsOAhVwqkIx2ggDZGU2SUhSYT0N2zibplbZWwDH28VfOXd
zISo8m4gYqhbCAVteuuA27dDXG7CpM8NoEUcX3+PqsFvj9K6/Ot1xY1PoblI+CH9
8MuKk95CEOctyJpgaW5jH4ud/mav8SJBKInXZym9CxS1IJovTWw/8boHWUwtfaFC
Ff9UbEDrsrvEF0kQiX1gF6uw6HQuiXzFixpTeTKxeq7IL0KPOzIbQv9yABCtfdLq
P3u7QAc0g2Zv5sTMB7/YF0o7fxyf+XtG0aAP3QCY3JBdvxovOhd2guvg5fM3nW+r
bvn3hs2Dtvsg4LG+XZbn6wJgnirLsDMF2suVlkUo/cT9RjhHs698kNqbTCmKW3w0
Che43znQd7fMysSrUP0BJ56mVLq2VimLqRY8ElMVHQy2zTFwOjx046TxFOAEzVyd
Mo9X/pQYiFETbaq4+pdnVhG7kYe7rNs9o9LvuM5yk/RISUzBp+0VYoVaZsOj1pnH
rDeMlAcqyq3WYqUhE8DUEEGaqzkihtmT4ld6xm7PnvY9amiEZvs918PWHKwJf7Xe
IEbtM/6gwF3Wcs+LjP5OxXp8/cfFHoVP+8WbL7/EWzq3EflPEA/AIICRAT9TOQE2
5kISjV2MIP7Utu8BjCyzoc7rpEA5Yvt6N3ns+li2Q07Xh7ZA6iq2rK1+xfBeqzGi
xeOmb9gzDlB1tO3Xluy+xTvSLQ2f1V9mZLKqt6BLBn9MApyBo50n/YDWHqXnx2nh
lVF370pTpTK6xwrW8TEYkaWFatA7aA3KskUSIFjzZqLwZJdPZDkm//UBmugY+w6/
vSsDSpBQfNKC46151jNyYHSaoX5CtNAvUWeBMnRC/w8kXIfy45fimcLhwxnfgSwe
7CrikzeGlxZ0ZHqEC2N4j+Iacy0Y5eR4Rt/9zZXJat8y6DHAuaDjMrnuD076/9W7
SqhH2EEdTuQnXcr81ccLu3717dxIjaqUtYWdP6VEX+5x/6vv7IF57idF30vTS9lr
fBRAQwW1joua7T1Yosg8YBay+Og01qRwqCFcrkEg3bBs8Jjn5WUerv8FYMMT8D1m
31wcAWCEEGzuFu0j3jli9/4b1/+w7tSr6xffbwId6e1sPt1foKHJgtK/DeIdGkwU
rkVaCNqQYAf8UDslmC9622QjrYMtEqkzqS+TaUrg05nHoOKSXhyp/u6e5FPlMCZl
KrvlNtcIuzvVS2ah4Lf9DGRs66EGst3cBt6hxKAefe+9s3PKIc/F/nswRPibw3cG
ZueR+CtvW4gO/JkjFgTVcGVIjLHShigjfWKLOsd7ekY61h0NOPWAuK+EINLgKIlL
8nw5iBUAuhKMX4sz44HyGAX+elGNlPwuzyGP8y8+Xj+v7ZciF4RZFrhxTdKy6n5j
Od9Mir7y+ASCLx4UAKYCBFXa6dFvIdTktcDmpA2c/Aj9EcJ+c/54rgkekwIdk/nE
KFgB5t7prxOBkVmJBbxxQ4abbhxtTmOjtItesa5lsrhAmxnoaxrdylFGBg4wB9Jy
3majnx+PssqA2JpGS7vmaO4/VJX+2zjqQBn9qqm/4s/Q1jpOx00eX1sQyKG0pfJS
0iHQx7bq0zQa8z9DM7s1rQAs2vxpy/ebe9/8/er4tNehcQuR4Gwif4Bm8mrrEWRw
tjuWozcObPN3LPZhbh5AqUzalOVpBBsfhFpxuDtOyxjxbDh3VDbYiqf8BoLYMaJi
T1yuptRwkEmanJTtWeMAe4oEVJgQOEuQYQ6EoSAs5R/4otbQomSXr/7ciuSFLfpA
NOrxLqy3X3DVkXImVGOCmd5ADf3v4+fJiEOaaNPZ/7SChFoReLHp97tmray3t/1s
rHwp0XR+PTzkEGkLfCvY3B7c+F/mtew7/XeR9rIZE9WjEfO6NgYp94R1rP/bLuzI
Us/UdTNwx0hf8s3vaNNyc6vsY+Eg2TZmDEsk21fmzDQAokOz6c6RSKoIjB2KRI59
9IPlgtuYP0turveBJ/wV3IsTXLA2BVhcNPGP3P+VHdGLFhT69hEy8EstTlcO5Yt0
5XEqoqi93reH6AG8x/mv8zSTuJ36R/9vIicys2yS7qoog1+UNC9iKmJL+/aPmk7e
8lIRgoQNcdTnVfbLLP8JwWwCr0nclxs9i1GN1vok8/Hsrc3go4VNXj/5QxlMbnlp
lxds2600sxGDYK9lX6D8BdF+XF1s8xH/AsgBR21FilsEI/CCFkMJ4ERdKCNyWPOG
QlVL1sO6b9G4Yu0sfIiLLPZ+8moMlup/iOWyqY7MFRMvYpPj4gSboQGTNB31FTUa
`protect END_PROTECTED
