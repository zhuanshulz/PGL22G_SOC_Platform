`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+GBSza28ehVMsa2KL5T+dXwixXipyJfGJ9B6cMNKOB+xLvPrg74jT0C5kEx0u2rk
oRlZIkJ5ercXoyCMZm9opgj72YfZ9XgHmLDDa1dWDol7TTEgfSPinxDIXNKrqXbG
+PrOIQ7jEp9HNiF6WYRchyUgBJlLQoYWcM7qK5/DBGqBTTiZ0t29l/evGTaj4n8w
Fq/zRKVSjmNku12EbJt1L4sw94uo+vLdIY56Py41a1JKIWC2kHcuNV2vuX897wro
E1oV4v5ZbGkbSDf2nbYSrP87/m0K8cnSLG+5x4lkEmE=
`protect END_PROTECTED
