`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zHSkk4TfzHy8WnpfzjBf+Mb9FZ78iabuBFksgVvhAh/BXh3YUHbd124xYYZAh+RF
/mkZyIwfVRymmSs/grEi65QxRpur9KMzzo+ryoLTi1+NnzjBZ5wwYrBdGN5p9JSy
kUhXCGEx7Ng9v+lxqUBVwJmuATxIj12Pe26tZzqFqszTpA86tyPQQFiLTLI4/Z6f
hexuAOakoRDf4pmfkmkku4xt5vgUJDnfpKmiZZ0WMx9245fIHFH3CHwFFtF7gIo3
EUb9j3ixv7VU+4zoOaNsxrI/rNOITCdxMg/UjuvUSQjd+Dm99UxsbMnMstxtz4af
Uo+LDxrTqbkOHovnV3pXFNsBA/qPvmtDiRpw0jHVIyj7fBa8mwzpTIQOd8wA5Zvg
S4AspvDwTDLuhwdTnWEVnIc2fR8C7X0Omo15SwELkcV1+1mjfEMb640K+g/D9P5e
s6i70Y0bqGh4Mz9iT2Towx58JsC4iZgrr0wOLABKVwEd82eOlbyxIpsD/WJWsRGx
Q1TsoAij/ol73i0FY/SFKNg1nyrASlQTS53aAJ/kGYlg+uZYjP2M8QD3wzZ6+c/M
Oj7PHj9wTr+DPOmIdqk9bCrZIcOk/OV/VUnug9xEUbp9kG35SXUlJxly61oAsQSk
kvXYXaBZTcpKq0i9b+eSozMmvyFc/OAHZCewVHM2e9Dh2d5vKWz/1ThVuHLLu0JF
pove4+e4nqvwI78n9u1jjUgOVhQLdJGOVrdYKDRF/1+CcSzLOaVVqZbPCQCesjDO
TXiitqGjhLA7Ij4xyVEZ7XXSnVF6bCx7poTFG1FfqeCuo4nP69Wx1B5kTNxJgqFg
tSWBhtb51Noeo16LHUvirjQZ+h+AUix1wBdXXX7oh7mpRdmD3jXGPV+xiOdvsWUn
sMOqejXn/0J1R2OGrxh+qOdRL7wL9c4d0BAtwoCQgwAnjp6w1azIMQ5h9kgpuwTp
ABzPuUkKa3Ig7TUs7DeF9pOdpznfE4qK36HbQYLLFHl79ZECZDCZ00SwsANZE6MD
G2tREUdgajoxlPMiWpcIVMoZGGofDt98Dj5TMyfgMWJHrZt2pHqk66AmuP6j/BAy
GHq8NZqtsfdNGInlXdpRvzzNG51894PvcvBj9AAL12eO/1sUiSCRS7IaNSviKRm5
RnHs83fxfxlwCnCCb9IUeNE7DyI9LM/IxYy7UuHmo2f16yha5H/J+gtGDSqZEpgq
yZqTRlThCfMdy0yvaFVIxGX5d6iD0494C2xNWRY081DQLKg/T1fCRKaP6AtvpanR
QTyLcDu9K3dAtROHpS8D96YJWz+xDYvM+xIEhEfQaBXBFH+/56icm4mYcy5Uau/8
lQFqMc+99kbJ01wOWrkxclijKlhYY1DXsbKx6O/NGCzCdO0zYeHSm47IdnKKCTGc
drjLtDDG2AR2uNAd6Mk2vn+drxFfi1LxLfMlCP4AEjSre+q3hbEc/ouK+Ktv+OC5
x4gMTsdyq6S52kNWK8DFnbu8FKsD1gG1uD9KHB+EsllIMzL0uezUVeb97DFW2YjG
A9/XOVUcNdUJD/X0iIplYUI6GJlOKvGGwZ3QhOVIdA5/28d9/7u2B8zvRvegLFno
8aVwb4lHw3uS9TRzOYDwGlY8pJFKeWXmbLc6pTytbnUMa50BoqaJxN6eleM3RlFO
QcEVVmgk7NjhjirH1modoHYwHQGtG+kXRYHWsf4H68onbtE66Je/QZ3PdfhXGvfI
RNQKdup9vDbriKbBnnn/q2mzOJnCOyYlOfBbIJ/hlsSnhQV0POLAXlH98ZzsywAM
ju7J56e4+ve9auylY/o5W7XnYL1vjLxTzOWthxI/65PiqHdWlGcePSwylFeSRy2e
bB1iLGSrq2n0bualqeRTJXi+FTE+/d0Cbh8zLOaADMoV/ay/UnvQhHrmf02Wa7ci
M/ewHgHwDWoyZJ3nS50I6ZszcuTaGMchONgMorgUJpiPiyPJpYr1UX1qvL4OVX0i
qkiZdjIWePiJWbt4k3di04Ip9+L4S6WdPCFH473stHUkVc8Hc4LG1klfcHDmUsJb
LEclKTtSYoiB1B09ZsdQYlYIDXxrYHAxKnt5+oWRuAaNRfMnFsF4F/bvhn6jt0t9
kH7H1CpLQjGzDjzyiwgZMTvZI/2NbXl64zzSbq9uHGs61Zn551/uJQuC2uuXsfRn
869Rri4WClSG8SN4X0Ns9nVWqR1TQOJH9670CcqYVyJfjjheTgnNrJINE8oM4IA2
IPTMw6YEcSoWYO7D0qcJAx25E3P5wJDSax9KknLoSWO9V4HkKor0KVLsRtkR/57m
QlkiCT+Xetb+iOTdczh4/9OF9ZllBVP5E2pv12rUkllO7S+SvVReuikhRXvOL76U
b4L9qwCsE2awkCqo2hossOX2UfljsTpdR8zYpn9SXPMFxUIYm83/lNwOFWpLJoWT
6RbUDV5G8fqd4dX+/M7XHN6VxsdlcOkcTlMZ74NFlasBtDKKk1xYcQVL1Yj03NQh
CTcejwwDZAlchQ+6vqVMIcNu2eRFA6E2WYd1GQQFn8KZPXc1nx4PfBKDf0Q7rk04
GQP9O+aBzPIsF2Iuo7wXI0B3dQ5tzM6krdx3HrWnksDUYj8w3tEz/Glh9csKhWVh
2B24bqpF5v+PQz/xnDVqc+SQp09sh8B9ASWluASYmVo=
`protect END_PROTECTED
