`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q6BIXC7whtHQtgIJ0gy32yGRkq+pjZAFnrVzzlO9afxT5+NPI5p/vIXdBsi/f3Io
OgMcmHShpi17ORp8K0AlyvnThVRB1Cb0KiVn2n4pYgTEr571fLFChTDlezeOwlbM
JZZgFfIF7zQvR/RDI2whd06u96X04jiTd/BO2v0Fngu4zsKv0iBS72iz+ZctyLLS
ybjaaxp3qMnkyDkMKNXoeSH7f+bpguFZ/MXdKl22uIL263Nyu3lhDYwaTDkqkqz8
/4AtTlNNFhuPf1G14dM6MlAMxy1quItQF18jV/72IDViYTLboxjM6htHnQCcduiR
A49oE6f6rkW3t6xX6s/P4AAHj4iIyGxtgQ8IXOXHiX5axM1eJDI47vcQldendj+8
IwnyiEraQgS2wfLl1wYqkw==
`protect END_PROTECTED
