`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YVT5c3YxAgWErQo9IQBWnm6dGRwLcvur7+oDYsWWA4x07XucJqLMxE297i0gXTcX
W9PCplrEjkqcnaF9fyBRp62boPC5XHEXPut4Xc3HfJBiObwAST08YtQltvlakKu/
yHlb1/d0th+oM5p4215MhMgLiapl23OcaSKXewKsGnHfXY3NPmkJKZdUSf1NpaQG
fq2FNt8FO6oBD2+/WfeL/AlC5MZoHPr3x/af2dnjbcGw6wF6T3AYkaGigrc7EniP
uKYkP2CtHIY7aj2jtDkPIFoxa9d7V3iB9wmjfhxJtV7F5iF6Dc3OkNudlL+OmGOt
vjhwKib26d6CJ/HuNE/1fmvPh3iBnKsfatxmPfIhVtKvgbmox8kVhl8u9PGno3Zz
Nm72GasX+ZmMzNRPdk5gLPkBchVYcthvnpMzAbactxIe9aPMyvf3HMX0kf2atkaP
F1Cb0QetyTW/6kHE31uzDHyTGg9iBg+KkkU2a+PIdYBtL3XrXe1JaaSQMWj6nhSv
3tpZSn6BbkQ0zwNdFXVqB2AwWnlqi5Zly/EBnWIXUTNfZxUkli2BzEFJemgIahIc
4HrHYjoIxVukr5nDzVBVIPmLbmhtfYQb9S39gyn7RH0jQWB/AxVYst8siLdgdvfL
gwfotUo9RsRbkH9ibDiPrsfuCHAVdoy9US0z/QuQuNXYPpSn/AHb7g8fKqB4XmC/
abXpRu1qyzIlLy76Bb9XY/E4fw3YUX3jRBH930y39VgIdql/+D0gAVfbJOh1bjMK
TIqml5JklTwzTw191uR/ISBpHOsDDMMAhYGxXUTQ4jjqdMecImVGLVomqIQQuDRH
9cjJj12zDW8fyZnSirTNaOqW/SH6Xnp3GWdamXM/6iunSqPeqZaVIACURluVv1v7
N7VtgSx8i7nz2DZrkU3OEZvShnqr9E3ARcWpv+FQIMU4r7VcpFw2fsRRfw6tbcHV
MmZDCd7gqylXY37V1jwJBZbVdy8VOMjIE77leRoeuH7STIuWT0/dYPAOO0S8b1Rm
Ndh/YzFiiJXZrRslUHTpULnE6Cw4xYSp6TGiznR45XTvDv55dmdpZQaGSp0WvWNL
5idyaF02NVKuoT276hl/aQoRpO37GUuepDOBhbHnUdy4YEJpKAtwHTAfVTaoy4L9
6R39XreW5eRTo/3SHIOqdVywkNlefymkCJ91Lm6iKs5AguSu82JU9vqyl/X6gjUe
F4QH9tCPg0uKlYZnkuBygSBxfpwVBQuMlJDShjN9E5+ugka/4of5Sv0P8mafYkp3
Kp8slTtEuNkkEZntQXqa09mDxDrJC+ztJcTEjxanaRAoe64VYaE7/e8LMLDFu7V3
36c//wPf9VCsazyWRolsFei18f47j+Rcx2x2olpe6vBdnk5HYc1cfsHvfXnpG/qp
KrxjImdZtBAGY2IqskBUfw==
`protect END_PROTECTED
