`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xblqTA6twm4vKvXFVFc6Oxkl8xwcSTGgifWBvlGIM0v1ccBMsVicfoVTybVAWABW
/M3voUnZLrzYifhJd+Hd5zZmg35q+RkF8g7QNroEj7r6jmozwpRYvTkrGQo+iZXl
qrSfcc9velnFsdhy5zO1Po22MVf/HolWbFwjirQX4sgHg1DwXS4OCBx/BRg88Hm2
l1W9O90S4kRp3EFX7rZiMsx5XTuKs/HZvg8qtkFn9HsP7sNDLlX0n/zMn/MwaA7d
s4Ymu3U/TtZNgHcUFM9Ddxs48uvc46EEPwr1N3XBC+DMDADb9kBgGQehIXTxdVoE
WaLWnn5WfkNUj9YT92s/p0jmcnyByJXyj6/mvAWBzqvqFh4XYluym/I9SHrvCkUE
`protect END_PROTECTED
