`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HvrqHZ11dV33cGJjx9XHJcxIESMXZk8Q8xkdmz9cKxRxKjhQ56Bs8z1+/L4Ffg3m
ZpJUSzpj3EZfs23vliNsDn1A1a6Agp4CkdyFmpd9JQ4jhg6j/VRQRGux5XVgKoIi
dC5BKF4P2KGWMHM9lKA9QWVXfuvvJE8dpDQmPuPBEOhyBNaecqLvqs2WuODzEPWp
3YxtL946QDg7MuDPmAAtbxNp8Qc/uQ+sEX7WNbw6vAeZS8TTjGJ+iKOoQ/dNRGHK
9pSlj5+PQudk17hzQMwxBA==
`protect END_PROTECTED
