`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUQ3aCQsPzxp23GVQYn2/WE1gdFyjPfNAnep7Fy79UzjzBJKhopCrieWf3GJB8Ua
2Let3VweGVGb/bLCEAMlTKHSKsJk6PJDvQjN40D0cAeYDqffQ6eASEp0ii6onpe1
sJa1nd/ANOIyaqEnG+yvfHNoO1FfzPaGUueqx0izlEw5gIWEe0KSm8H9gOZSmFL9
b0vmTpK9jf2OfTXSarGGKbxKHueo63D0WBFB5pUqu1mC8+rQ//lKbsCthHcWW13S
rA+YTpzXCnu8Y28F2CBc8mDuUn4X9KoEMRZbCSojeis=
`protect END_PROTECTED
