`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w24jo2jDYHsNIkwPuPIKnwKMrHEDpHn49s4vYGAJY6gr+OqAqxm30P6lAbWP7Mmo
OcDiDRxO2xEjwwUbnEYkS8iLFPD734bMOibZsuTp039lCBdcUjbsMw2TFWI0MCqQ
Cq8T0zipxilIS36hl70+F98mht9SAEXu/dAvGHK0T7fF8ntl/BA/TcqddoJQrNvq
Ttc5BKUA7V7lrP0y438JozmEPTjbJNx82sCIRbWVnqBV6XkDRjXC3qP17V8XYTwR
NZvM4zprI+jKsYUyH+E70zB8r6+PLXtGfU5diDL8FjZoJkhQUdBLPH+lCs+luj/Z
zrbDtUBjzoxYsMhipbulU9HZf1yTJkMGu96TQucPO1W4cHm2jd+ETPqyQXfrvOZu
khcHHwgR99QhEVuTsd2k+Vh1QPRJalcSevCMEYWzui5ICjkBZ7kWkoTCRuxjvI7q
hBX0ymteK8ZzdQ1MoiGG65QKMKWLHawdjzkNbvAGYAW38G1IwQiURvLBWAnlK1Eq
ko43K3p/87uEy6aW8BrGXNFGPAF56S0YCF/CEzlkks0qYFa1a0IFZLaeW9Z+q978
Mwy8rBuDBzs6zdTs4ATBif8Op9R7z1h3TJMjL6WsuJnDR7cfY1DYmVrLsobaLBxZ
iPJSl6QDXr9HNmB1qst2btELh8uVkrh9JZ74EOPEDYI7+vpBn7kcF4TgZyRJyg53
93rpq2e+P5FAYSiQK1U8yP59i/hW+meXNFgTlW2FRvxnZNCSGtSVj8/E1x4L2YTa
EJ6WcQ1ESjP6cJb7q8whRbXg9wzSaEqjSxeclv1XwKMZy4E01LrUfL7IaPjvTEzX
veOScEwjjylYnVU+CWB+8geZhPnY3JQdgUccfpJRV12iYnocdVZI+eYdxa8wi2gO
+kN0kQ2pLp0jSPLkd9EC7haCgkd62paNLquKe1rpD3psSaNpP3bAnO/biFMId80A
Ovt4H2QMqI8ZceK/hicZMvxGAMHbWuOwvc0NMVsI1oRg7fTQC1WCp0q9pUmjg6BL
lCna67XyJin1XK4ZeiU55jqCaUZE5GTu2UnpZTqc0Md+HPrQhF1f5JHeC2t/QxAU
D/T8XhQXlllmBAu8lfbOa+cdx/TxnyW0IyLamjD5I2YGmI9Nf5pwso8y2goTujwo
f++Ufw4u8artADj32FNmfb8pEVO+y+y6djUVQsu+6uez0ZtfYClwiiKvMVHX1KDB
QvRwmUPHTbI+Ze8xlVbh5ecumBUIqZBToJ84taVJsV2QecsEYitfFOE2Tc7ZOZew
kXWuuETg/KH/t/7xlNkJ2PCXtpiOnKdJ5nTP9hxh8UHnKtaYTEBnLDJDNpW/QXBj
Gdspr7JZ55uJVWaXDQv592SxmUhZjEHQS/lrz7KIu3pNVKKKrlVYXcumCQy8VGdr
2FdIQFi3sfbX0cpyfqTswqNwmqWuVxrTOF3YlLb58C5IsNLgy1JlqRLknETeeat5
KR2SSFnOg5zKp0/QAlt7t9WbbwEUKI4fUpq979ZsAAd9LUjnRqGCPOrYhp4fX9SI
jZnnZPiWA+gp7FIubPnlbR1jZ28sIRxJdYjZUuCXrNfx0fMKA3H++lpDDlfYxDlL
Z8xDarb0vr1effJLmqebpNiTCGdHNfyJg4Awyom3j5KfmVTz9axJPZuee81jtldB
qaNRH/e2P9YsdfvHfR8eU3k7MorQGa0KQ9eCBsK/v1UrqjMrLV/LBh19DfdAHSYT
wpaIxhPwX40iPPzDKhCm02Xav1GuPxYHhpGGZK/QM5siK2bWIdiXI1km6e9GGaqe
e0E3P3RbsVtiG26MEMW4gp3w4HMkUTXptbGoyVuynCB8ixW5KzwEfKEcrNDgoVNY
9UctNhVWLZ6ozep8b4aUMv7qhy7hg1KzC6IVi1PyJ9kDufvs+xR62gac8Ly4c9cx
xQ4o4YGyfGa923da3XmDHKshADZwFFrC04tJk26oSz0=
`protect END_PROTECTED
