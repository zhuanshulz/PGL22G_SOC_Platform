`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zF/15tHS72hvmhN3Griqwb78yeX94SZziUf1KF2cFrXAR83TW8ZIIBZF7rSh1oKD
xSMMBdJFs4z2gFwBHv2edifGIZJWKY+dgv1jdu2hcu1Ndqn6uF8nRIzIsb9nHLW8
a36AtmVqibN5VRzQdY7r5zAxMh322ytpSZAahPGNSy4jAmqaYQrXx0XjpSQetSjZ
clroXxDrI1v0itv3RWoHVWT6XMiSCifARwltI9m7GZDEo1pKmAqhl3IgrFNeWV7P
vP6vTn+XLifUC+dbrb99XMsIAGG9ZX/MjOj3aAhpL3k5c3Ia6M/UEEidTBnzN0Yw
DrkaDyZdL5pPGFDwPArKaOv0ajziYywq7wU+AxTI0qdl6caZY6lF5tmi0o2uKN4E
pMo9IF6NOUf0uGxekgNNOmqHAS2qPfXIt2uFC9AO6eeF8k2FxogkdOztm2ISpYKc
ohzXhxGIQ+N5FRxG+vaaukkW7jbK8/impXpTSdUqKVsCHfT8C52Orx+H9NHYsqwq
dAP5AEfXALeXAv+/0KrX6a8dlqxYd5Ua/5ug8/vQKDWd5XoQaktLEC1lMH8YVFQQ
vCJQSTGWHxgHIbw5Nl8jPkE8Us2eQJluDyHK4qSzZGxNnjbld4vXyEMCtbW5Wlm6
8DfjC2t9YOc5hEuF/ekHuYUweILBDomrxd+B68Mx1cDhSh4AVOsWil5f0Qjupfdi
XPefIdQhOI4dXkKszlV3O+yQFK1sgp75jARa4i4lfslFYiDWfJJd3mOg7ZnXZ7wg
jw5qvlL+gP77ieNRO3gHxfY2eB5eOOYFgnf0TmUdyCG1QGkoKeGNCfSbXYJumdQO
Gg8AH/MzYnRf06wahMv/dC8BirlaUKmJNb2T9F3MBjp1ezMHIGEbAUXXhqulgbhj
oZUAYeJPdCOXJpd2bD3pVFnd/TwhVGYjP/gRSmwW9i+HFjFv1mfOo5mYVNIqdFns
CJ6tTiIMtvJkKfTeCOzpRDjGu9DRL2ZIHzLsvAb7+j6jbHC/U9MM2bP2LDnxoPZz
PkLOIcCsIUrLkxywoYOj0VZBvSQ9tpTPKpk+X5h4r8Y9J2xi01GJ+GmeDjpCUklg
f/q27pIic8738yOtjuw4haPHaboTQXgNayatkXcjNg7g2q2e/Xt0B0/GbVFBLYKC
FXWuxUqcvmIhspBKfoO8qaXjM3tgQWW/i3mIsyNzQ71KE6nM4C6+CM9x2PewVTLt
nRVSHdT+tJe9zT63wepJRN5hklVnbkN6RpHJrPc+w21nZBDbOYMphoUy6BeafUtI
ECmQ3EDklbLPcjM8SWqxrz7MC3KtuFfB7tvF1vRmI1M8Vaaqk3TVtR4Ava6Fja3K
wntsDe66RK9eslCwC/B2NJikzWWpGQCUu7D+o75+va1YXuN1cJWbSCTJrPTXF8yv
vZQ+lCAlO7DUAXm7b8Ea1pcFE2vRLokivYjZghWMfVhh+w0PhrIlr22DywqXZp3j
lTibcErjGCrarNG71R0rDuiFZMjV3PnqC/arlIDso5BwLb6CbYFOeO2RsFxIN+Nq
ZWbg3Qz4Xu8FSYyegFNKfmPLYPE75pB5DCGh1eoulS7sxRW7p2z2Ehp0kQnMIrxS
K5phCR1BetNcEI3t4JXHjQqFABY03kpYsCBkxFAUH8NXGPx2wKTq2LvLW0T2QU1K
1fGnONPt5n6t642UjkrD2UbRAGuLFjTjmp2tfiPh19RLqAGdwKR/9SVcGYUu3v+d
bBcqOn3fmA8dqKLoeM7uy5hgo/KixXrBaY8bBs1+LHExWOhX5XFZNcVAhNJ9QI7q
ZxwJoAgQYzrxNt6dIJpAcbAxkYqLNUr80/IyiAif7mP9Jyo0FPj5gWYc+ZKwKpMs
9MIFch1YdTS6UbowENpHBDVJCA3geBeRSgOVEAXUOVhoyaAopKuyDNNLn/Q5gSoS
luQ3Na229zeJJvP6ZXoXORzHZCs1TKAebcUllE98C8Bycf/DmSH9sl0LTeeUdaH/
JkFxNB82KPp0wXO1ODk/q5wUlVfjWWiM2LACzBXVci8xmNX9dtHl/B1fMfRXwoc8
6L4LdiBKsj46HtPUqOkhWUL6v51kn5rK+7tfvaOfuOfOWoWek2H9bBiHfqA01KsQ
FXinp/QyuJTKzIu7R6ipEpxvYSF2L44uY9dTNOFhVb6xAvuYlxL3I7MUaIb1xGlv
TqDGcJqeV/Ms9Bvudu2lBtoGELp05dwgi/EOupJeAqn/QJKShXABUcW6xXRpS2v4
dt3cWcVYoJgEcVrPJUQhd9j2VGKVKvj4wqLQ6mLdvEU5s1dP0CAvNiLzZHH7/QFb
tmRlYEmtpBXITcANsN08lkxTnnztjIgWpSttRLSmteDPT72G2SUperFeZ8xme3Us
kL/od7lpC+lU3F1w8QvUH5H0gKhHGaidlu1XCaAy0Ak0StGmhXHLWpNhvdzWpsUw
yq/FSxoF4Zp9NekTCjF554POLfUqBvnWd3ipk4sy+b7fd8qwNcPrgl1hX4KVQlF9
SUG7+0xD5FrmHn/paEKYF1DvMVevqPU/G3w9E1cKC/e2ODZ+DMVaZ/4o+Pppfo2G
cTR+khofZF3YhlnlTWfGbEiNm4YrAAJjP3KlAKBG+Gkvp1OyqoJ4U4quTCx+zmTE
Oorj/QrJ+HLtmDfOuF2jAmja6foSaezQEnMRGpMpzQFE2M937/5qKxWo4nuvUysZ
lM/dbRQOWrfuBF7mD4O9a3NJQ817zLWdBrGdYmFFzKBMpQ0bVdd4vgy9kKgbPp3C
bynndRy8i95QlUDnljue26Dov5f4acb1xwit08MNknp3Kc7pRchEX4q7DlLPH8D8
BO2jB2a2I61UdxVcYejWLwu1YYCSbNFMsPDttM5YCn8WK3aBmRHNe6bp4XRmNQ6r
iUplZ+OQGjTQmK2FuOopBQD54C9pxcmerO5k0/86aKAErVsV8HhS8D3zB5ADztQQ
mITHCEm0rdj9sYMDnRWO0a9sinU3N6N9XD5fnLV/90ZwQZHBQftmz3HY41UiqNE7
83SQ4mJJfslvZhMZL1uE3pZoL6S+qb7fhqJJg/7d7J9lMylLMCErD0SWzAsSOely
5ur+rFEi07pa+X8KjGleYrQvN+AFWGCXsa2fd7MmSlt3CFITzG97wyT01u6PTHUa
SVxSOONGyj+tVqhiQk7vciGTuRhFD3ROyd1NxBE/4VN7pnYCQHfVqZKIkNGSQYNs
pEuzHmeP5pQe8fj143OpiyzjYEHOYZcHckhL5CMkjgIt/rvD+YqvwVUF6CQ2LuHy
StIWBQGahevJOO9S81paPZ6+Tkq0AzjWs2i1hV6M82zsBXuKXjgtu354SlxEXAGe
7pjF4+Y8Y6T4PWT5CELHO7pGL5G6b7YyIRteUQvpZjjM7ZbG69KQC1shYR/F8tnk
NU1RNZc0A8IMyZPYSDQgcenXpSKUM+6pFrPbm0gs7uPc7np1JQWUpQkpRJ8FmR2I
2pddc1gq7lp8IZ7dxPd06kJaMDk3AQoO/PM8HvtLCENjrELpg2SPx77P7++EhkBY
+4LwPSpAaHLcpp9BGwGIBpppA/q2vTQZaDbvhrZmW3kbnY2RbD3RWQanM50gdOK+
87O0uD1GnYkAJbi8kMSRItVsUbYnIQ+SgOlkAw5aKJ+qmVsasSxAshrBS34Ljzw7
vIg+pH5suPZ+y3LtrZ2GaSsntpVB36UwD2BCkDCy0Cz/+pcOEid9f22Tdms3a9Zg
BhlTVMWnAGaElyeSlPBnKkcibQ+/ZCKJwM67kj06kuEs069q0TSqnR9T25ioGkcC
QtK2uzRqb7Q4tFXcodj4Ki60Q3nVRqTtJNukt6L9710/NDoQAMQOSANvGWZCqMGB
F22thsiUzO/iakJY10jNd2f+GSwN1YTJHFKqFKMn5wZyIIrYerY18L6tCDNzsQwm
a7qMD30vl2bMsEGih4LdEMPGQZbEbBtVEilUUYkmXYeo3xbNSAYPvz4yYK9PaZB1
pH2Dcg6P/5K3BL201EGA5bRYR8UhvcYLT2X8uyeq5DCQmEzqal6qk7+JsH9uyISW
4Cih5+CyZtGZ2hnXgdNZVjNcla6bfzriztoW1vjPSsuM4Yxpz7rHtGy9nTra73v1
NuEybMpqcCBITcoAFTIPd/1LwIuU1fL9EPfrTPTnhVMaL9jMUdcqmriwc+Ee/wru
oTQ4dbEYrKqijNjABit07IeoCLamcQmE2Cu2Tbc8N/bAFryGXZRBrarVqumkE8+3
L1QnYrINEaslecaNopgs/nxvvUOABx3NMjg4uWAmZugWZiZwm10bMfMpO9epcFH/
ze7BWdDjwtMw7LquzTVbPkDUB/VDpfGiGq3C/s7TBvypKCXFhdVis7Zky8zqiBit
VlqwXI865DADVXnADLtTQY/WgQwKXXEQY6hFM87A2FbsPqBHEPdIoGJZkrUz1ONj
UfPCeKIgZlMG2i73ECpIwZrbWUYXsUV8XLzZE8bWEd2E7qK59eSUuiYF33jxWoc4
euOmM7LruLcEUqmdpwrKWPziB1VEoP2yOkOwf7SjTC6wH7mMyYRM6tOolcaM41R1
gKip86j0W+zWnncJMy3tVtHUAAK+NUvql4wr3fAt4k9I0Tm87hcZABXY2Uk3+SDZ
/kstEBSV8VhRWavl+U5tYVCIibmeetgfj9P63sbSNwwiTzZZuWWwNbR/nUZraG0m
QSYoDK/IR1zMZI3JNFrGPtkDfQfsNaVSMLMkpc6+gMiVI24TfxVj6yC4KE4MesET
sxQIPVLjSveOZeZL1a+8hhh/DwCtcoPzQpnI3F0we8ogYLqxZe8cEdK1fyPRbx28
8vRfuo4tTrhOSW4mwBCgKSvbMbRfUH2WFJVoO2rewKmrrqOkhgPOF4KLvS8GQJ7R
KqNoF9vqT3kd+7wTKBiKmAhqWnzeS1SqAJpiOpTM3RA76L+LUtY1Vedb4qzhsRJD
6324sGM8loAq0APpC0IHhNe0FKENRtpuoY0L/3We9dP1bYFf+8UXn8uIwvJu9QpU
MDWpR8Is2svWo5VE6oxAMaYVfUe0oymTZ4lVzh7zO8dNpj80gOw0M731l4glPL5y
Ik360xjZiFsKaviFW/LDfIfXP0tEpM5K2KSeJ2a+6/TTH/6i9kvspdMj1CoiPTai
P1y8AYOY6DlYA/ATwRLLkVi3ekiRKv9BC0ggAdaSgLUKG7xl4CuJGOI/t2CzHb01
+Uara1sUL4cmMYLfnz8M5cAu4AP8hEF8ousXBmnaYkxCnhWVYZyN+XBM/8JRxtXK
f0NsXi8vgltPdxOdLSVcAsU24rw2+KOK7tjJtbQNwrMwpBsEI5GhGQFSiqvfwVyo
ew27nLkGsSSiBwQqC33XfIj3ipmlsuEuWX9es+obR1RsNkVL9JWSWsa+9vYuttb5
EoZfxpQdmPoqFEIujLoKGPDwaMZRvMzNY25SXzXPc1SjfLFI3Y/ynjXSWwPy9f+T
sOvIpdpttv8Ng0QVJZ/y8Q==
`protect END_PROTECTED
