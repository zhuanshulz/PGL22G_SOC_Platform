`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUcQx0mbSycUGWgI0x2zle70Hp6PftIA8Q7V1v7Q+FlGyhKwX5aTQTdVl4W7EHWv
0RmM4t4dmFjW1utzD9zpLNGhy/Ujh+3KwPZMd1rffzYMu8Vm8jU3tM7o5ndWGoEE
jw0HpW6KKSVg9L/eLDgdMn2vgNiziXs8gKhBygP0aET/XaYM5U2gsvE7KTUNqZi7
sP1WTnB8gLz0bbaDBXEGhvWa7bxApmPIdTSNwwNGSbXj0B6LRfCr62n4Xb7PwNk8
ogMtBE8xA1XuGVApVAbD7JGbLIos6GCr4W2DjNjPv/JZIM5diPFjcJhJKFCPt3/u
umqyJ64X0j/5qkBBZ7Gc2G+1nWvPLlI6mf1Xg1Qm8nN+uZ8LT2MXKVkJs6ykw6VW
UpWrx4RcjbJQiwnT1nYsSN09noHd3/zDfjWX4IcBpST4yQOTlpiyV4CLehXgvanb
s3ix3gyXGd+nKqtTnmb3QTVuUxnH/L9oQCF9ctoYQpiQG+lo87mSWpsqUxUDXDB/
eG7KRFbQjgM6ZeiRHYaSjZJQ2DgL8D8sXJ9Bnn/wWpo6LA7Gr4U3gv28F94WMNua
d3e8Vi5WyucWgY83L4YnC9PG+GNWTjPd/Lt0FZPcbHY1YYppueW+R7yJU3x21oot
JdNTzFK0uPCcBd1lb3WK/XzPKJ7WNrtFMEVqIprH+7zapuFpe6G19BH9etKIZJZJ
Pc0ynzAKj5DaEEmn/7PKWUQMXYHHKqjIc39WLiIQUsnxbipFjjwhqXcceauo3vv0
q10Vr7eIjYUyZqht13LSUtP4HJ2NjP0VpHF3blsYi/tWojrvuJomMyOb0udgwGIv
px8Pfy+ZTfVCY2uunVDyM/uWtEMhdeRhoVsVu27f1DInFJE5HBk1pLEvbMfR1kES
V1A+HQpIVkV5UODQEzE0o9cv1VRagd8naRaiz2PtlNdkjRDsRdtQJPs/4XfIEyBq
qDicRIPZqDLFCd/ANgvT7/o9J848f2ndwCQzXllezBWMdepaBkN/1zYkeBVbS8sl
5w34zk6wIQK1e1QzEKwzMyxS4N02Sw19j1YWvJKf9G2jniG3l8t5KcgdoaJrKycY
ISE4sF45SXw6X2XJx3y6uDtPQSMKuhNcVgLIvm/dCk8FjzIHbhoI4oUfPdmLILMA
/YEByu4/dLy7KVu0Isfx6k3EUyXYsHcAnqEPcB22TzIIlMqGUOmlBidltCz1ESfn
937y384AKHTM+LpwCrHHCd03jp9y55K7s05rpX1kzumtN41Gl/F94jqDCSK2U0zy
CHj0YrmqfJlmx3ZQvpcu7k34dn6IfzWv78j+BJ7JJn88zNGdKpKtR8YRlhiJr26O
gqlRf8akTrW/buYMQtDkQVptcLg/CLwbO1B5ANajNHjtuJnLoctXTgYJ7pEzvFwr
GEuBRnQiCjXMilIpodtXst3LmRrXmY18vGNXnWPCRXNYHk+4+byKUwDUgiqPeTbe
0s9PdK9bMIwXs7CNI127xQ==
`protect END_PROTECTED
