`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/ctnHCD3wU/JsQJsOVQyYlWJa3YjxvbK3WKkU5N+rGLQ9d4AfbV6W4bwuzHy6Ws
h+k/e92gIQyABp0xKFz/gUDMZOJ7zQgvs7Yklsjyhxli7Ks7IAbY3FGE8qmSIuhZ
jqSakUwIA52uOa14lxpMSO5cua9bEr+p1XDyWhTnq8Ilnet+7O6GElCSbo2Ics5z
Cr/pB/ZIHeKVOGUiQyWSMjZ1wHwIQASYEricb6lk4+tKhb58jOK/Y2avmgP1RFMD
mxZru64fL58G9BLgrzXNzw==
`protect END_PROTECTED
