`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrwBL/Yn6xr8ZHZh0Ga4RCEKOSnE8hToTJ1HccuusVfniZe0XTuO4212qjre2Zar
nexGBu2QXNIC2/jfL0iK+eXRBV/KwIh2gEg94hSZcGUqSwBj5AhGvySE2IPL5tEz
qAo89xFDjziJzA9gHtga93sroTAU5D625EewW/AghkGfBDh3OYMk1hma2tmFtVee
VWgZ2Qd6oy4gYORt3wU/LhiJtPd8eswrrN2s4O7x6WhOyU48bdUiwg6Uam3CMNkg
Gj4dVN43wkgJrHyEWPtJAw2RgQ9Z3NE9gCXJVawhYlZXyWEi5FkAtQPfjZfbIgf1
+AIu/lh36K25INn1J0k8O0aIyDfXmmJSO9R4nFFU+KXL8tM6OcTlKNz/YzMoCJCp
vbXXoG99Di27NgT4LdJpuqh2AzlIuU1kUbzFg9VNhTjFP9gCgXURZndEwLpYeMAX
CBw7YEgCZlhY9WOoH75o6un6CIPSz0Ah5sBGVUaVBZlgvM9dwsExsKjCpJMFyA+e
Ak5Iap1vkItIZwcgQ5JPb4mr4n3DyJ9rCKLZ79xXZGQQDjnhE0MBTPaLkP+7rawG
Wx+/HFQ36BttUoT4YEPHzEAtCMew2pMlcbhRHYAMik/Zn7C1vMYcy9pKTdYoDUvg
e4a+HDQR6hoSbOsqnXLE1wxs9VX5vYKywcc7riZrUCb103VNLrL4oECuu9AsVePC
LWqDwlncRcKjTUTzJ9CBdj6U49v5zgGv2J90B+AWNRDMbk+EcqLmRm42Fn83CYX4
nc/4poFwLeyqV9l2nuMBAJZ332CBE0XcgKseDYld3DpSnpHSnaFP9mfQOzDpQzcA
D1pUN0D7/7uQvOEw7oR5D+1kP+nfCTFQXkx7h/ckpZIKAvCbfw7GNSJLsgPo+Rrs
hyg7RbmSbeNxcZfW90TZ8XQrPgjtKt3Kwip+O2am0TTirpbjLsH22DYXfQC6wNsB
oXe34J6lXjDr2R0+U3M3SLr0H53p1U4h1q9ALTv6I9idztaz0iH7Mdkr8UT//rNW
nfaYdmPv4rM4iNdRVp4n//t8dgwuTLBKh2FtmTQAH70=
`protect END_PROTECTED
