`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
knw4vOt8aQPOpVN+cmKo3pbG0GeMP2JGeKoQR8nhlaW8TvJ8VXJSWD6CjkDk5ltx
sCMTMPc6Z4/YaIe9KeOpWVsQTjNClWwkL23ndiZmqVSWQzfxwP8kh2RJ2qnbDb+L
Qlifiqs2xGAgExTKP2JgVMXu8Dgke+83jv5+GGKWY3YEMd3GdmDXvRlbEJ9kchIq
kWit0D75uZwJLqqjdyEThwDHb9eT5cDnHJ6C12ngyCPp3quBTDPu/CRLqYge8zeL
C9h/Rev+3WUV3xXBjAZHQweBPdTbuG6JR4MVw+rGCT/yxYVTXufM3V+LEDs43MSb
LvpI6OxHkXMJpSwQEDBSrgBrdusZ1YFEjK4rnEodQ+PnrVgEglw8EoMFm+jh2zYu
z7k7zjgIqDgmiPCZOH7qL+GQ3NuzSnd4iSmJXOKBoy9O1rNMb+OJdoAnGMWz4z/m
FttmtaQhNyA8DRisz7fFqA/joCYi/w3k6vSRhmj1Z1i89pjoGFFF2tT1Yy0hG1Z/
jfFtvBw8uJI5KKrHkr2zKbHDf8e3AoBrlYazp/ffwdaqLvj6M6OPHCMzSbrD3t0g
A2e5zU+4edN5hlb85x053hdvmpmOoiajcTpKRZrMTx+ZNtsz0DtQoNnoCZZybJBg
6lng6aAlju9pHhfZTnemTFXrbWuLDQqnJyHCpQs5uTC7BNzrFi4zzB4ne9NulEJK
nLchY9Lj4eaWyjyD57g+b5T/Br24ZYEd10IdL4MhD42yRD0mlbJerAAvEPvBvTOq
kWPXuiHpgPZ0U8W2W7xSyW/A7jXyfSfIxp8U4SVEiSXkeqXYe7MGIzmbD8oYADWZ
cSubpw6loGusq7XzThteodSDX8OQdXqjxuplC2BSPbtz/adruz7+ZiVT60jbGB7K
EOi6aBWGgznUJpUfUDfjMWQB5FAAxlQbc8190g2pacoBtha6Wy9D1SONwofVGc+1
ErmsmLasAVgbV3CgJ/gwoPNxQjenubrCRsak1sChFrdd87JVmp3KF/fjQQL/8ugg
IYmT2fl8GdBP/TUNWg0Z5EG+IXD3Tkw/y8r16d+hZXCYYr/pEXwqcc+RNLy9hj2h
WVi9z7lwAlDfWjYBCZ7WLv8MSksCuQ0cOg9ReEecu1Cx9RXcYskIyMLU5jDexLKx
4IjbweFOR+fLpkcdgAaxhWgJZExa3A+yJ6hGDqZ47jR0/vXvi2cvi7ejmNC977ks
gIhhZoU91s+KiZ5u56UbHaJhzyJ6IvY96S14YiS/UpBSYQa1oQeUjm9VL2UiIOTt
COKVx77+7q04DwllDvW+Kw==
`protect END_PROTECTED
