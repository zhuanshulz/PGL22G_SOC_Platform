`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lv9ITQplgV+KcuZqQqnps2HEk5KzLKoNsdLPPWJE03JhNXRHumadJhBGRh9C/WkN
6VUefo56Z2GEQtTPDLfOO+J4g+YWMMWe+RFXDkyu7KbItYiko4rcx8uwk1NxY9Y9
JIl/uXvqyDvB52ux9kbbamyuGoxnnwHi5y8SJzub7Q86M0XfwwQ5hY8jte8VU/u2
o84N4QmjA8tezD4PiW+JiUPZGyHlrQ3X6S2XPuThAe7Q3qE1IgE854DcRSI9gK1z
UflZ4CtILxM7JLFf+OlJFPeOJIh4zRGFUZYG51WsGabHVPnYUOPHbWgZhtmzF09z
FQSkB34HlBjkVzcKA+RbIl8zYIGv1AxDnBn7cl8bM8DOUhqEiKMtL6qJvtqXFlUy
Rk4UYejYIXekeK6u4oHfr2bCV1FZXi3iWufM8sSOlNZW93Z3JuxIwf5NiiISp3cF
ZmlmbeXgenkafdIna0C6jjimzyxH45FvDxvSDxtUnmSZ1cXwXkCL+5xK29KJu90Y
zI0Cc5vIiojiuc7ODVYDAwdvQh7pcx8M1kSCmx8kiy53uBSX+KK2kLg2G0aD/EPJ
gg3kPmUoo+27C6FDsB+G7gEPf6UVqRjK0h4YcgRn1nK/GYjGAK76oMmkzYo+ISr9
DeKGwxprLSa+kHNXj6XR8xW7BkVU+/cSDAtEe0Ahb4CHwA1FDqjefBbYF3j4moT5
NvAfMpqo1u50kjJHKoFU5YAd3w32yXQaKTTkb3+e19txFyzd+cI7i1JOSK+gPzdD
b1qQSTMThx5fH1UCHxZ2vcb1UayOy9YSIXYRyhsH/I9ezjOAWYUtLt95P85qls5S
yXgTpKG80oM2OlLrwH7ITVRJIn7cT+SgTgwCaxcWaCJRXXzowlEGoh+BOP3dab/X
BDNm60jCoo+RP9F8Iq2dq4dekjogJcZXXwYj9W478IsAjdvvlg5UuP7vckm3e5lF
sSgWQpOVAl+r0jdr6eLLdhlOG7ddvm/5NCxrh/ZSa0ivBfcLwsNWVDjamIjqYHPH
YgayA5BEfS1SeBVmrGIRGz8zOr5a8mtoWVrJY1L7RLHM/KNiUCrGW3YyQqJk6qd9
38/kMVgSF8Pvua/efvjuwgekENJXD7BjLroAeIQe0JwglNQ6dXNiX3cLucstUi2S
JX0P609bvwAHhwJkidRntHSpLyNE7a8ZCVr6Jtma+q8QBHIEX2R/c3IHyORTeO1k
j9g9NPytRMxM4yi8YXW+F1Qq1Zogw4WB1K01cF/R91Di4ThzvaKN6EyRlpnwyz6i
RSMmFBHc+9EJ9geF1uiefcXqBUjqaYWrDPEyvwrJpUy6IYVV4NREO5CiNq6/PF39
2DgpV387Gr053Dk/860CR7JeA7slbVItFxhUYwe6Q2OZsH7ngE5XCpzE9xhxuDd0
0NLlTIBRgqKeU1a45/4HOs6zWYC0Sa5It30L/HGwRaVsyAD00VUty3K/wywH6cR+
Tjk1KuzW4hj0DpGb5ila5vw7gXhtDR5ykdLsViJNZXLQRRV+EulefbfLNxZyiz0X
hhHQvKqQ5eqmKBVXb+H8jjrZlJRfZGRryCtmtPCWR20BFL4IyZiY9L6yjOk4dK5A
en/3rM/RonXmRVkQRfB9caEpu3v51OIQmdrw7+8OlUov+FC7GGiLP5KmZPVxhyqn
Uj9Bz4NjR32N2Zt/zuV0qX4herJTUI5hozMKqwXWRPyDAcXfxLX60hc6fnym1MOk
u/eD3FWCRMpt7CrtvAGMLjNlkRGqG3/t4X8RDrFJaEtyDy+xto5IgMdBK96SEIh1
uHZBq1JPHG1lYQ6JhHmUgkrC/ZkkHtUK3f9xpDiuDIB2y0OrZayPPhZtHTQcrXWB
ZibnUI6+Ay9tMHlMAHyEPf5XROq1MR1+S4Ldo54yF5iyZ+qeFcW2jk82Ux/N41CJ
FJLl42Lux6rO7Cop8KxKaciKhKMt/tUHXBI5W2IcrlW/OYiYaXWVrUPe/niOPqzC
ZvC++x23gFJE70rg0KDT8OS3vCLOujBmMJsAfc927xszF8MzVPTpVBl7sepUDKxE
eIoXIt0CvGPD2VbjUD863hoPhYICElmLLENJxB0TgnZEH+JmlW3dHDHzkcf4slPD
99Hd/IOLRpDAXdLaZuPpDN/fvLgPAZWVysEt/G/REJrS2REc++UvLerbTSbYf03P
TQm7dPh6neu9ulKn5wOjmtfG9gBcW+rm7CSld8mleRWIyqVjeXtg4NElveOUo9Ud
cBuphkg/GF8qAZwG2FxkjsWa2aKialqc667L4DjYa2coM1hIxObHsGpmYRrwmwuO
5R1A14kBeWGYTx1Trg0fQQA6mHjvmpcc/TXOcnsTRLNHypmE+2EbHKKbycPx6XDl
ModpepVmll7+z8i8wqlgz/tY03/dbMaDxo8zYK8apX+xRCmQ5wSL120m/eIapjO3
95F5Zn3VERvP/PoXtLWulrUjjjbaRmpsPlDkxmjfy71zWY/Pyi6A+t3RL53S+56a
UHbQLMQO/ZTewH+PIKxRnPp5/vQIGnXoNJtZ3GDRykDMPOe/I1a4oD4DVcls72Ol
iIjnivvXhhCmx5bEBHXhCUyR2cXniGKzT2/S8pxZUv8hAoJnWeeGWzMP5h8I3u9m
iurlChidnM3VgQ3uHuKdpRA0aD3cXFKHbRf3kepriAHi7/VwU/4jBT9Vb/+DJLsx
/lSFaAwvXKnIXUs7hgfvlJQXoPxK0JUa8T+LCPP6hAxk6NOTdI3pgtP6Qv46Mc/R
y5dHcZr72YNSbq9Vi4saQRZ6SsQgoP3ldbr7V+0QdNCCc3/eni80ni+XOF46BYg2
iFGS7sSpTLt4F3YmM76zUFBybxtO/CqJWNZhSeMU+vUpdd4xfCGwCxqlCMXYbvNv
4lXtUV58Y06webERt54v0GkYxmaraniCeinNAvXURZUY72AjUUOYGpBGWa8OQZQr
parwt4bg2PdtoQKtU8+CdflZLo55fgxshACsqtPkzziAj9n+h/o03UvZzmxluoMW
I15DDiHmRffPr6yht11nr2L/hwd9ugTQeaMyTLyZWFKpvHSGPsMw4f1bW7AASOnX
DFjmqzcCc07Kf85bvJ2TTUiF1u4ZNAv+lezxVffWkf4g0reGnxQQA0dxOP1nIJSA
59tiVe/QbCzSbmPvloFyrsdioAymapwoTV8Fvm9TXCZrCvAg2+vJpmq7bRPHhDqs
TfgaUSkIH/zBGYez4MbGJZPcZEX4B0XkmaFdEvIXPTxfEU6XLeijbBxKTpXi3MDK
um4upwsSYNGqdnwfxkjADyXGw2T/Cip++ANMlM2l7yNinCD7DHX5UfUgPomZ/x2l
WewnYw7UIgY94MZetjjpovkq7M0JRD8V14t6iswvh87Dv+ZxdLpPyHTQllgvN0mM
6eFyIc4sGgwh1zNy9Fh2siHZshp1/y39+CzYp3w/MlshjKQpGkEQ0PvanNltVTbk
8lL3jbM05b7BLlbQwagTc50Dkca3W1Esrp7RKqXTCm7adBKvFrrm11SRY/5GUmNr
HwDcR2BzW1FEzmZoswZ59A==
`protect END_PROTECTED
