`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6IeRuFjqLSM/qN+5EwetqEMkVOmSSKKt+OlBhR/WQJKf68yszuJCcro+fygu1bt
/l/1Mi4DNZ75i4J2mumaLG9ByGUe1Z7VmDC16IOg4X+2czSr33MNAf5KZRTXDwvF
nhNb/isXseCswAKTyCZ91RMtdQwQBB72Mpm7jxptdGW/J8Tn3HpN02WoZds5I8K/
oe6w0wxcn825QsNlMen1winTslOMeX9NMOWgbsQ9zAKyJTaMucEoVadQbdBOwB5O
U/ebUHbf2YrtRIKKYL3G/NB7CbQqXgQTBk3EVZCRkq3oQyhu1ukK8ptFlNp1dRti
8KcYRDXZsOORkqxKIjHv5TIbIhmb3lz77BMAv3u/SvklfZM0/XQLI0ZyCXF8P/79
iboQNfBXuIsHSDWtwCJe1RH/6RV1RcgXReUb810Ce+o/A5oRuqKNMna+Ug8xx+aP
6PCmLEJWw+TdX2YLSr9MyUPFsifWqioANtq7k5Xa298rLl54nElzhMApBGNbqEn6
9a1ZF27c9+iTKIKYtLbtgLN+n840KivJsCgUyFdi79WWYuhYjMZs0DO3ixTrxm6X
pvWjN3g8dOGo2t84VO1mZ0HrxyykRWkAgiJL79TpI3+Eo5c+JLHuqTSF32NDlEZO
zG5K27ejGv/1kwFfy/A70FdRC8eL/4GVAv3isf7uQ3g9uIBME1/rF1ZdrCxytcpv
FqdHaE2EKQ2k/oDWTkgzX9B+PjBaS63SPsvZnmEaB0NTxAr41II2Jklyfteg72S+
maorSpHWS/7w4hZvlpNQaub8jw/dkjDj+Azec7fQcE4rxLjbp9fCIvnzsXd8qkBQ
4uNZx/CM3S071AZp/4nk4GzRTIiIgAYXKlMeJNCtq0YuH0w8QwJiUaDUalVYAPGA
dqwd6pmVFTDVWChqvuqQUOLUlEsXywppNm3Re+Pc5BsnhCiW0tjl7noJfHmnGCkn
KhpOoRh7zPfXS3ZzADNgdksyz6sMvS5rc9xQea9ahVIc3bPGqC4JeKF20zN7G8Hu
+d3yZzZ3Mw3IM0kk/A65ZUUjYZZKyA92Uw0OkDsHBrXHBuCTeOuO4YyUDPvVG9SB
SA7F2sD3FYW3c9Zj9HtZkaEY50uL01hItUErLE+vkqPASjGuLZO7ch9kX/xN8lnz
w2tmCbXW66VNIFw4xlK1m5R0xP/slrhlgzvvyKcvvCQWmPodzyAgmyX/dCgab/6q
TvYWeMg0U8idKRCkE//V4F3kImRFQ0BMQEOq6sZ327hyG08GCw/wMjUkm6L37RwS
JtszgA4C13R82NUcgttqygriuEDqyAIokAjRpHrlhsFZRwVfMBDcaZ9ZlllOXTvr
gOJGMeffi/t06+I7bb7C3eghgGvNNSpfy/IB16njg4WS6r3EZFP/sADfPAQWBZUy
6b4kcdqeHZOiYD2AT/CSrSbidjLVOiGUc52Fj9CzE6mRYva+e5Vl0EQAwQDJKAi7
WzxpT9C5o9XUAhu87MOO9EYyD9vI/MkNofN74fPeCI8L7q6wE7cvpnuyx0uX7AxO
NP91ROpxd8g3GZoQhsFBoV2w4B7yzf+RqFqvuNbeBeBpCeyKJNKurycefmqWiFsE
yZlN8LxZ4/9AffJskSIMGf58hdpVS4patCGsrbVJs0OLqpU5l6fXNmIw6lXnSue+
tJ7vWl3TBWH77bVBGWFaxc9tXJ1PWYK7A0/vNCr6HmWP1UrCU+3uZ7Vmv/+XKJm5
Y3nIerTMcqNogLW8c2u4MNpaw3JiU+M18eyEWLMkLwbKpQcLUVlYYHsP2AvDNEMb
/ye5becrzRHgt/Xt9FI8bGiEFBAkKxvUPBEwVsojZna/Z+twB9OpQRFgSRvbZzfl
l1XNLhPV8r9Fd+Nc0fWz3zAXyJSozOiP6BhSTGVo2Qg1oHDeGyqeHvbDiv04Uk+2
KV7q6ojBmDAT4BgaQeQPu6Cb6eb8jckIEx5zGq1y9yCcSztYCpeqzoaSobr07sd9
650XV1c93UD/rwtdhynMamxrlTuZkJRgSsbE3ihOs3TEidQeRvF3Lje7ldovKo0W
Kl7GIWgx75ZjeW+WMCgryJRjpUBtFN2nQOR0TodEkyxn/A8wbvF33QWKRBsLpGIM
gHYY49nJh+3jdvi5Qpv+JHsAjc2lrCvIPG7ukjfkMWWkvjrGKtdG4OBOY1b9y8vG
es4+P4oSiCKehF7ie6VFwmvIvdbQSfVddD3RQcl0+WyhcxDjx0+v09ykGUirfnYR
SioGa2XTm7dNjKHWgxOn+aVSQr1rwYRGTMeMhuhh/kFEXRDo3SXkyQgo1lXp3K6Y
VE152gEGboCjshmRR+Vw2AjaBDjElglXuQZFjcx8ZY1mZ3LeUc0jEwzP1Dbk8W+F
knY8oJym5e5YOGxNcgRpzJVwwLmX6MEO6wQvJw4tDl4wZq883IM99Mgs3+WXVK+R
tLiUyOqq0uUWkGkyOzQSGIXjdJdYqz+wvi4kG9m+MKChk6QRI7W3Akaq7gK4PURK
5wOMa490Yo3Diip5TKTxiIYeKqJwOV7GvOXHEKLJ8u3HV+mEYv/3iVa77YzD35zB
ManMGjWcwwP6u5hBmO1UQVllunK62VTKsLsBFOd4nU1WxkVC6kVSp4pRpU45kvu+
LxBaCxjjpwvH3eHn2Dt9aK+u6KCK2c3RYzt3ni9iV4g5RjkaBCd8Ey6ioxhd+Zou
6octD4fgyoXfNJ8VBYEho5l7w3EA/z/I3AUveD+9g/kTyIBNGydQ1V5nbmOJ0XXj
pjlf5QxfVa5bgmUiRrPVrwX0725/Edwfw+brEw4O2ksFkruDxaJHODghG2ExGhf0
QizmYOoM3NVq7thcZleiORh6QkD56ysh91sD+0pXgoYb49KdKObzkM+L4QoQO7LX
9LzoKP49K9pRmAiOsYad5WcReF1mLRjV58YODKaDxiOl7JQ2ilX3T/kPoO9dSWiD
26RzPgxtOF1NhEfIxqNZsOWFl+V+HPRA1k7nbjbMsLwo+XrxD8djhzOO/clkVt7Q
NVPxQlHVDYrwUGLSrhLJIGyOypXZysA4b1y4vye3Qg3OmFbmhVHkPnl3XqPIz5Ix
CgE9CQEOl3mRaTrRD+GTkoKJFRzLp7tIn7HCnY+kRUqITG91sW9dyQdIjX7Gyq3B
P+E8AB4Mpkrj3FQnw1n9VRidAsMQNvqGjtQrH8RGDp391CJJqzhhoxLl/EyvF0zk
X6vFpqRjyBRfm5fmfWhbLvlgXHR6JDG9fuP3dXRtrqaBWUooaWTXsvosWcxZext6
cUweDmcDNgQcgWasw+jUYyzDhTOXHiO8oRCad5Pd34xSAkGBVpwMfU3qnZPooMlW
Sf9Wmhm1evcrnDL0zp6S1gAhJueyvOREXi6toNj4pWuS7vrlcgsfBvgs9N7dS9T0
+xTRfkGWNLKP1HN0MvJ1J+WJJMmsqOwcv59O279nmXVwPoYcKzHJaGNnYt0/dO4U
fOfEmW30ifP7mEaXmZbHM6TJZZRt/fnCZxQIpuI9TQKxlkjl0NB9FmdgxYqgathm
ILo+Sd7T3DcRyZGh4bwPdIS5+uptXidG4EcaeQALhdNQ1AqihysHoNAcjgPQ4ww+
+X/u+1rfvXoK1uT9hCdc+KRVbswyYJnm6k/T6J2YOV3vOYRH5GNx6L8qP5WkFPgY
xh4wpZ2d/GJbk9E4gHaop4B7bSrvEI4pmvuJm7DE1X2rnUAJmjceZWmbXrfqwqv5
n4AAp/Okk5okCve/RJCGeaYOJ318gIzC3pjE216D0S7y9kSYf+EJ2n8r+Ju6RMzx
eUCVigjzbqbkSPGyxbtiAoDrPUYV9IkTtmiHHwTIcUCYGvQ5lZUuVCRunDHRSPh+
+/HTnvYyxY3wX4WKV/qwszhJkInbAxDAWbq8t+2QMvyxRqpwEwRiBvHPnTtLklV0
/Bdf6Gars04Bq73D8tnRXIw7MGRHKGw5uSd4LauArDBSofGptmK9nrRKiCRTxiMr
hbvU7VK9UnM1gLPdpXmtV7RS7LFHLE1SOYVMqmNXKcmTcy61X4H7G1nz7DD8iW+J
XUl36P0+DadXMIAjBLnA3IjkxBnp4TkSaYLAgwB6UNUXDE/stgeQB15OcusYcRxS
8QldcXhHNqSNEtQAhjeOAobq7+GVWDCJneI6U4tWUxNqY1WU26c75NB5KOGaPL77
f5KAaQpBmOlrU0rnGcFC6igRscdA6YXlFSL9/6YTXWYxCYkKtKRXq8l4XSoIPHeg
PcodjM0upZjPXBWM9bIep/IEaSR+degXUSNkvLsgLiDCDrVkCUGGlfRoB+zpDVYp
xre4hcmVVVClHJz7390XdYsU7vAUiolsI+3a+FZf4Z/61ccTjMnMtWreuX6C+CoW
i6EAkEGcZrnuFY27MDAp50ea+nDjEM59OYVRQdlCCFL0w83uT5Mjusp2S5AT5hTo
+h1CQaB+YSMaVmaMy7T5WAjpOegSwPX69Fa+U5fJF05kpuz2QXBIzD+RJb8/JSXM
btEknFbvzHKEz7cN5g4u5tj1gunjFnNYZ03pg6T4c7UrIvFaMrLpMh73sRehSYDc
Dun9+YYK/EN4sASFl6TMMwJZt2ZtUA4wxKQvKSR9T/T+2i24TQHgUXbf/IwUQwNs
YljlahPvKX6cdgVG7jArIUToGkAMCEwB4XWqq7D/G4uaHvC3zt09omZfrQBHmmlI
S6GM1q23HR8yGBdjtpyUiqA3EOzQp0cfR/+bkAdMpRu8UOtZL7xseeQUoKxtDWQk
QA284I/fLoHxkHqAR6a59eld2II7tPFk8VVYXQWFmTVtyep5PaSUXA7hg+fLlEDF
CNkoB3SpzVfEI02WTfb22e6p3sv9qHyEH7d0f14TJNVEHYgBklqL1iiptsmaIKFW
R9Ah2Fjx3XTkbL5wwdDw2A9w79ob6cJpuDUWlOrKjRM6TpdJ3b0h0Yv9ulAEodOA
dvG33X7wfQQaChtd9hKSkaKNKlKPt+zP4tMJUKCBd0eFMlXaDOfPhLvR3SkqWLVl
hoqOFK68Tor6geBNO0RwtLNKTMn1CwXBiNDkLtnJ/SDMmz2L8lMDnup0uRUzNeqY
iZeSBBK1ER7lucCEu6jQ5PmU1iucBJb1LN6qxEyg0z/2h1dzfQPQ5nqsteAHNfCz
BzMEcq/7yxwFs9YlG4YAEPVDTd2xv2hMHOwdfq2ywgu3VQt47evU9z2g3N4LnruM
dZVJHRTOmxTjs0sZogfAyzz5E5lY4C6zzxLM8B4rOrw8JDXDvAubmc6M3nHcjzUY
rpoNqi/i9ERH/P1A+aopZ+0kETwvq2D800x7DJL5+sLHp+f8GtF4fi4XBUKPtZ22
H3+YrDxRqIbNSpAzVWUv4MMBckzVWObbrRGVmPfvJrL0Nk9VO5ua07Kn/JEZL5nu
zdporQIOrGg4Xky75e7iGWEAjczGiRkcO5uzSIr9xNLaYsKYTl7lujoQF5Gqq0oO
dotwJ+sDFfBW8dVPW6nJEuipt2X3M7O667UYXhB4AuBcgLgQjEDKBlyCI1guApYR
qO0jmVsULBqG+DYMmwwUzYtqwI05is7Ym3Qy7WasvVdJc6cc2S26sON5RqnWHeqq
pIR7QRLTUuO4yMQ1ogmtOwDQRzHZl5kpgnvX/iLQaVAZgyhg8uugbNetYzskklOd
fIvpBFPT19rZZFhPG0vIG3vhC/MvmD9ZZWl0IICD2RXmDWZktDdCS6rXbvU3p1qR
fBdtCfRkl+AJnD0r2lfp4grF8yAQuTxxAHMuv3ZICdXMxI9qmleheNtxRNyKFhvN
aekkJwij97QwSq2EQ1sz9B1utjgm5XmQ+E2YcTIjQ1xDGEbaysRkf0WGpzBoGz8c
SOexxsQw44qY326ZEab4QZUCRdxHowQ74szprYGk0Oo3sITyMwNqSr4p/15+ZZPw
IEwd7dFLSiwXnr6HGSwOpjG92CPBZYs3HkU1uAZRNi7emKy8shFF5kHn7V4duCWi
aIxDtN/tS+ae+7QP82LkVOQ9uMvnZsdPnnTOR6WTwMFBsaBporHFi+h2Z9jM0ypR
SBajyNAhA9HE9Z/0UMfbdTx+1oLwxjneRkNiMo9SHd1L+gZ9ZnntgIMU3HWtB4Ay
Hc9QISqj6OInJQXF/ae3K+M/vTQ7UcL1Ck8cW9rUrCU1j+k9o1tSYPIxROM6pedu
33HQPq6Vsgdk9BGupKimPRx7yBa4zR5R7Y/Va3ALVy6mDDlMfW3Qf6QvdvqQs8ZS
4KG6HpZJMWGfj6mIw1OOYF/xaM3w+WQbY+Qg0LuNPCYHGpol2HKamzGD4qlqS+l8
rQJPpESxB+g598pxobDitVbOkGUvouExNRJTUe6Qa5zzOJ00jMqSlbxNAEqdCF3T
Gn5ydzEikZUHZO94JAO3fWvtyDQXjhZB5kZI7C3QNBLQ04W6QjIH3DCKV3ea2eBW
O5PRY5dYCqsUwThlA5ShE/a1fCOzO2SX3p+iqdHnAJxrQZKjVfunUEQ4deN1BVa5
h6PyxtfGXGsIhn0TNbzSsjHWg8r976pYIZs4+VZdywKu8I9lNPx6sjiLYAbgCjl2
ldWOaaswej+FYJSzfQAliRlLsNkECH0L0zNyASP6ghe4pxdz4Qj6FfhvvkTMT+SO
lktMNy422eDwTANpAzDOLskRIk01EClt3OfrJrl6aETP14f7zqPR4XH29khDJwSU
3uljhyVjZO1THyjaty141wAPvCmS+XsxKTGx+r7TKzrMWBUlsG+3rNJaECxCZlnW
Zd+1wTjpz1q1d3SzIS+D2x/nCF29L3+rZqibGGg6pLLRytcXxu6iQALiBXN/p4N4
+hPlspPl5U21eHMvlGrNDkCOsVmTS0Xm8GAZ8pjWVd2d5yofcWY2N+AJVycazZI1
yuDApmYt1Mf8t3inJ09iGoZ9Rgx6la2eSF7aQg4yOUwcJzgR1Y1NQYNCo9rYc4VI
idsUsTSDN63aQQNFh78k3yrLzYLqDqqhtdgK1Yy8bhp632+Vfp1+ibmcs0Dnjj1l
JlRCOEYHShDF9hnM2sJVcwCH+Nepra2KTSfBZby74+xG6U5VFZbiEDkJgKMkpMyv
Hd3/L1uAh/0a/YoX5wq65cBwLbw6lwIiK+WaxQCwp48W9krv64QIxH2MkROKDwT4
LlDUluzFutB/1GncWZW/LjahXTwsXgK9pvY0ELc3sOT3sI7eMaIXvMjBYt4MIlxp
4o5tI8BPfWk6NjBDi6RfgSFJhTTuHzrmJ5Ej17vGExKKxlJG/ukAl8bR5oCOphlP
H+tk/+Rc2UXf/RlBe5Vws4rXg5ggea8lN2IWgj5Si7dSvtgNmggXzC46W+uDPWfE
Moh7dFzh9jsrGLKdCYtMlmgNcC9XREBVJcpQPdUCUOiHM1JLrK0GlWJ0HxutX12A
6fdCUks9aOxrV2uMTmTqhdZoSzRxgYeaK7JDUPrBewb18VZ7j353btfDMJSSVT+S
L+BdIRaIuKn9Ea7v7Lctuv/sDl0K45yC4VRFNWboiMjzmvKOLIy3FFKCF9APr4Un
eHK7PTYgp1JP1b8r4bWvYGCh88/iz63ifFitr7HHNvu2vJcnAk8SGoQTQ1xUFG0/
KTp5B8t0upRV+oljTWpqvf8SiZNH4GO+qJ8CoD4KJPRxW6+Gqyjp2Y/8FrUtFU13
Z8JuJeTxJmjn5xExemU7/OznhRbrzk2oPoUVXeh6tqRjP8PrRfc/awAL4xk9Q5AK
ADWd+TJb8WtrCb8ht92fIctOVR+cIN7X4IAPzmAVpX1ppokHIQFyuvMOctf9FWE4
PqxsGlziQRcei3vdVsTJx2Ni98foDNLCXahC1zDVno/1ugPn7qnygcUl6yXI/BA+
406PatAcm5HXSKh86qeZsDfF0QX/z8oRaGidT7q+OiX9r6sOf7KDhtkSVln58djc
u2UW1w3K2iTuOT5+wamsJlTf32oTzXGHf9aQSn0orv0Th5HfneYBBNjnJYABVcKL
pbKFRKTaOGVfafK4RbWH7O/UQJYC23EIsoLnToJIqQnDD22KiH6nWyc9bDkUgCOx
73TPuJzqOiRIp+/V8r4lMPdlfmfUkyWN/Xj1Wkv+1oCP6xLiDMLJzqCI8B7KbRyn
6Advx3v4/84EFEdXmbJDJbZE0/EbVUT9VsGibchMoU8pArkUshMmTAOJ2NsuVoH3
en07liTeNBFubHNnsYEY1yDpmLgzgdx+QcFsc0j6IxWXMEGOLN6hSqW1i2RlsaiZ
ezuJiQ/jebtSQbhi/jlMXCw8GmJeljjAtBoP5pHN3G/ujBc7zOgUx8JFD8rds7iK
IWRNthxqNEnABpdMdu/Q+ys+5tbH1e1XRkRYrjUGAJfe4Fb11NjGWFOKBByYg+QZ
qEYYgXQ/wSGwRVew9R/sNaK2lsGePLTCJExtY6XiPvuGFBed8DVauiMv6Dl7IueY
j6eRrdKq6fxNgQCKTp9KUQrrcEeDxklsZ7oxGZ+NYZBcvbRCEPrwv9Oqp1JQcwRr
Gs3C0ch15vi4lALbF/qzrvRjlS0fMexs/hrawSggsdMXoc7tB+ACr7n+FtMCkIvK
azCZmxAR+ZI94dVxhbLs0VP0iWNHHv50aX+TJKvgFbmjlmfK3Edl+V2FDmnvsxc+
mRsvEXFg/3mxOJcpn/xn8zaRRJNTT9k9fKCUdVUrYUyyY6U4NN4pR0qqACZbMol4
wY+CdAKlo8C7UWbPSAfsU2h/2xseUAVTeDYtnpHdHPF/+52ssAcZIy6ZhE4Ryh3W
LAMIVPoBG6xNw1N6Lt5PyxoYuZ8TNrBWxYtBrdO0puHCs5HwDY45JXK8Eykw35o7
AWr1ZHi5oBnlZLL+g/5zhOU4NOQId+HPZvyHqedhaMtfNEstosE//c1cVJDPXwNA
lML2S4fwXyo2TMV6NzDgWPm/StzS5WmuFwfkJ1LOnbaK0mS9aKGA3/5dJlk97N0Y
ygcPmHII6aAhwz3D2+lkDgqamwv6N6zJ1aeY1ifrBxVHVYxCytj1A38ThmV2BFLB
QM8kUmft2uVJrYdCv8HTuxG33teOEY8wr7BeN2WoJwki1f+vkqdrDg1ZBlMvi4eW
Waog1kdEs7S+dmH9/YKb5ktiJf1FSUPHkyOvrd7jfOXPior7cvkJpa1ZWFVW+VHg
Z42J3ZmF2uJUVESwTfpF54seK6xbwgAxf8W01rZbuu/NaG3DESv4uC1BpTTmTbOR
izjQmNWmxDobbt2XbhJhrxVb1ZsdZsPcT8FFmKFbw+G+OP78y/EcBJwlCfb01oau
w3BesXH9Cg2nRFDmeo9kOnAlSLqq2W2PIxTLMtkp1a1krnLPDG6Sx6QLNv5sxs8B
8KzjJnvMxCKD3ilxhO2zOzCT4rnYxdYuysCiK04XFt8UXpG6PktEFkYramqv7wmH
VkPTtNrfSvLx/Gb3NQ3kcc0vzT3BBc4aK1SjFKDSQ9+d3fqdvoOvr/ma19+GpJIa
2Hr4UwGGblskIObtDLvye4BB4MclGmJpbaCo1PgR7pf+jEBAaKtmjtuosdVIrfgA
fUGOpiKaSVZ+ztR79MQ+U0rbJ+Uyuoeb3Nm01fNOROr1YrsZU2O0gqO5fxrk2zTl
r/agbEx4XPjAN2Cd5siZpFzVI/CH9aaOw+ApfAyuXLoPwmrKtzottMQSZ3FH3WpG
jVY4khzX+yDvh85kxeu8gtbv6b3uWG//K3t7FoE0qAUwJHnHIEH3+olfZLyMJ/tx
vlmTzKxe+2Dz1CKQ/34b9USmx5Z0w3N8qLGHFFAASPv5RPuXiPpnFRKRzuObhtwu
Wt24UPAD//AYqC/Z244rDuQUGrZ7rALA/AeqqY4FCahTTfHPtHEJXf+qPZZ2euVm
nX1tJHp3wpTj3UlTgCX/16JibUVVOrzVgCYr5Nb02G94zUTvnU+3pWNmlonemnQm
+UlRb9b3kZc1MZflmqhC/aSlvVj72jdVm8XROoFn4N/BXNNIgp2A5d1+yRgX8v1D
KxMXlWVLkFBLdlpnFgnZpU/vH3YCiW1TaRAcxgOvNNlXjFHzq00HcsJBh0q5hsqz
Qe84ZgayRiQ7UfjqPrFasoKcVLkrC1VXcBtyHv05XmDFj9zY1NZjBcQydZ1Cl66o
B/DsrOrZHsQ0k7oSWQHN/J0oCJn9iJOobXJ5DML+DDBljaEKtRPGqExezfRVRlJk
FNtfngcQws5LnuKCy5+Mv8H8xFWn//z15rDpf3Iz9jk5D4J9ypLRFPM1zkYPStSM
qKnTL4t0PjhgEEiYWbuIba/ubb9SMDPHcyZMAtzIjY2c1ewEsmgCRTxoo1wPCT7i
e8//K6vA5P5FjfH0TYC3sOVAaGV059lZ/UuUwxTB92/5zY8+PdNeFAammD+00sAf
/EV26vZT7hyCL/N/2gqAk2PNQ306aUqwOA2C/lV+TzSfurkHsEq2z1GwyeN9Mpg1
L41se54bFEQNuyxdbMEQGT4Gud0p5rhOZbTegAgdLhCoWJI2BwfKxDFILl1q1LDg
nCNNFr0/MuvRpn0Rf4QceyUtnX6HSmE2RHz+qSv3dfsD8ZJZIGObByojSmjW5sxR
dk17qahZ+VPNpWfanWQHRH70UlMpsNOKanvBV+xwFUCBGF2mCJw4mfjMZDT8jff3
yHcWbGxGaJWTWXqebJTFUSbSdXHfIs+loqIBta0H33lEzIcFGhcn5WJUFJLR7lK5
ieuXxqbS/sSoKdW9hZMA70zhoHLT/yrimQdPTtZ3akVbNjl0Dm4DItq7+wWHOxH+
BqVqcyCnOwvSNJ4WWDsPWlsLxis8m7I7RuuZLKkh2/oZAAKro2Qgomx/u6gauJX0
yP7bUNraFy1BiY2t/WnH+2zHdqvcI8mYhKbZnGCkTVKdbnqUfrdpe+j+DOWHCHVR
H5KPtsSTP9uCfrnZvIBjDmA90ASl3LdjPf959jCmw2Jd1FL45XDuhOEm9b0Lq4kl
btR2MDO7peMNLtodyvrnpsjVP0gCz81l4Z67ce0edAEMu1YVx68oN5uve2Oy6AeE
VNz2uHBEn3HVEHlv0q71uDeJ8ojSBsiTxkuDnDv8QErdQJuZwPafuychyYPEfH52
7wQm95ikXp/eiLx4uHGteAU0Ci8/UexGD0YQ9l3UuTjoV7rXbI3FG7AOMu4/up2+
5qA9i1qAPaCPgVN6gQoI3ulfI/EDqhdi/IZE8/H8QcFNv833LenhtPFwV+OyPc5w
L/Vx+3m09j8DHjxxbRZPHBSf6e8R8nU2c1N+ysWfW0Vf7t4Esynep+MS3sn/OEpN
l1i9W1b4V+WuHxkDxKZ9tGIJgOWVdV99HQ67yLy1HOaTAsKjDw0CbO4YzLGzmNTA
f55hoMIsfKVFCXrGWcj9i6wCp8/46+eS9N9ktfvMfj+8uQ1Y2HrOSX1PAbjc2FWV
XfwwDa4CONonz4T5dP5ayw9m5BiuQHX3QPJWaZEkDQSwJ/Udc8UegHi6TUTm03bN
LbSAzB1AmCYCkcKHQiS+RW5LK2sCck+ehaT8UkidTK8W1se1kWH/+gunilMChU2M
we6+wp60N451xm35MZcTbrmlk1qVzhfYECEvupug6k24ql9kUdzymPIdKA8f5r9Q
aoLhLj3l5R5koPi9aDdCZlyy8CjyG6zNCWm98zWzrvOyhPgey/hvk3H4MgGJvI/e
oHISeoYo/JhTVutIulXIe1zSp2t+fU7bmTybfy8ud3E/+S6VYk7Oixc8OJC6GX4i
/0xBbM+WyNzTm0o/O3DEupqjbZw3Ix8kMlijHjO302t04/vLp4Ndk75Fe9dFbFLx
FycrT8uoeL3UkCZjmda7K/j0/tbizzCsygvgbALBp/hC9eegHpYEMyAeAKbm0J8e
tcVU2QXNiXoV1h3EgBTKzxjkL6+p9fv2Iq2kr1ywt/VUUk6yrVf5Of/6KXhyRn6V
j0z/wcXJ/++QF+3/dtM17JLxkKgy44339eZq6gi9M0ptLlOZIb03PHDYP2veIueA
vS/7/48sSZw7VLljT6mIMjZ3Ml2gHjfvZgzJdRUdboZMAjfCkYNofV4MF8SfEUXd
kQTRID+aYs3FRl7og5h++PsE17KjVk41G0eSNMozqshvtKYGxNesjmlTjPKw5Ggv
HNvyckFE3cf1K0JM0u9d5Yr4rn8Mf7gc11sYthEhO9L16GkQ6q7AURUusnyFb713
hI9KNd03KqC/e8+tqP2Y/CITb/Ed8+z6BJbK/1KPjElwNorlHKBUuXdHz7uroEKl
pEw1ar6PsN8TvqAL1taKiRjUDxZrckfuR36FLiAkwNeegyVAPdMtZ3L675KTrlkk
NCPJnFKLdl9O7fNoPD1cJb2lK+/VyANODmEpTC8zJlqD7DYLDfkWb/nZdKrQv0it
pdcP20Byr1XoHI1alxl5RtQ2fnooz7MAjhyUkScUFiA+IfOw8If73+3GzM9cnDCL
j7wCiUS2KMp5kcNJvHo5hCUcFOBCw60NDW4XEkNkzxMZ9Wp1H8ICLrzfp42tS0Un
dyt/YoJgVQVXC/h6XQwqN+wNtwRixMk1O1NUsk4oYlEg2K5OSn53fuQ8/MbCMfs2
8yxKxHZzZa8O4Fy+ejtKqUcNkJRFD7MweMPuX8T2JCDffH8s/1eqasVuEH2MIM38
OKqTJZp9ZD64wKbv7qi7TuO1s72uDUhddZat8XyTx7+LHV1xt3z+sneTGiqPOQIs
fw3NwpQh9vIwfoJxS77YeGPmCN9kMt3iNvykny7Lr+GkrLV3dWC7ygrA58nvEvzL
x+H0IO8fbjQWzOqN9ovH5zW1ULr4r21seegOVZCvDdUebAgDHqapuQYQzhe9tZcQ
WjiPYG1UUNU8oFoDRGCNaXn//H2zPmUK8r1vOoiOaEreW2ATzbi2GovVb7A+xYJZ
L3oX/9ki/wPQ2rzGxgW07wkpIwO+JldnunqEzNeFZ2gqGYZyoYI2IzCt2d/qVou+
52yydvngPXoZR4vSts0p9XgIHGaFxjrn7n1op9OmFDrW1mC1aOb8Na4A4gCmP5Jz
yqJTXKj/v8MjjvMT7REm58jJqfiMEndN99JUQBgs1urtdrRkQhcawwCM24Nw9/9v
gJElNhwlz2uiOBHkaWIw5nnJ8z/NrXiyS14SQAfigtBMeivrRw5KroKBaiSV08E/
DCETK1XuQEPTHEcg8qHlAZVW9NZFSM0DgjPx9Bq6TsnnYpOaaBpdc15bDC1PyTtC
mxsyRmK7z/pE3OBnf13V3QNp0sZoW7pQ1gCY+BSmN6leRWbbHsPK/UtsaV8vHIVb
5VYbKKYvd3nNPO39G8mcaEfx1FDcgcSbAZTu2RELgo6GuWgHKQN6kf5Ns6289Xt0
/+Lp6sT1NC2C3xoz3KcUFKSOGA5oI32381n26iBArFC2AEVR3lGkoATEq9t89c/v
aui+e8tzGXC59/JE2QyPvulJhBfKUiw74RXDWn0B9hk7wBXv8pPmlFaEUPdNRl+e
BO2T89VLxKswiKBASpaiNpPbyPihHkJuaOjV7RdFSPVqaCoC9IvQ+nvEiIHhYxL4
rk9jlOi5qZ7lrFzJRX5fq1U6Y0y4LvIP1lhMYBp3of9UF1Ucv6gKCs22ryBPxRzg
q6P82GJSnYGDz2/k5LzObAbVB7QnEAiVW3NUSf2A+TjDYm2zS6XqBz45lB7wHV0/
QlAIizmwzclq+4ZnLXRIN2MGUq9dzTSBpSz8A/U9nLgk8PKrly4BYSRFA5w4CFvN
dUE190kzJkHVxFoyZILheT0JWAO/xq/MRFNeqEI/zzg2WMqUl2tPzJpVViEBANj8
qZAYW2k/wNY2YwwliQ+72RxYNHZejYYM5CUigcNKKfPNDKmy6oXBUQF95++kWpHA
Bs6N2rWnccxHY+11XWltmW8Jh/Rl9nbK/e/xhV6HmIAEdu9ElYYwnfsxVflVehXE
qbDChl0RF8Cn+6HPyUCFZ41b0sndOIwUBNVsIZhAdT1Qc7JI9dljtPFWj6suPNbx
GHBMEtbQNXPWlauZ6hxnk5Nroj6qyQ+Hcp7ugIRcwYYgx/AeiByBevdyBrq4068R
tcPpXZNdppxK0i2xoBQ+2j3LpHrIVBY3NQywTpBkHJpJLy+0/NHqClHt7OkKSk80
bj8TjDYyRVsSLMasvILaPn87/q8AmCEtnxHbSjJZ1+Ma84/b+SSjhw65nyq0dk2h
ygRmRJGivUAaEc7N1E9mqHI0wcEa3MFpLdt8CGwddakj1B3sk7x6Bg+JuPecfKrQ
5ZDlXISaO4Q47tjg2I4RaepHKD743tQ/uiCgVciqa9VQ035Ykyz73ob9f1VpK9Ye
JN37dT3N6mZPCU4lUrx83Apv/AoNgJzW0kXY7afytbt4PwvHk+EbAIjVQV6iNYGO
1rk5G6gpgLAsm1r6xOb8xOwC6HPYhoxqkKfNN5mkVECBJVXinFO1+YPYnXyCBjpo
JXRkVxiBtUskU2y+tLkd+FEJkw3DWdE2b8TARdz73zs5OteD446pF8oi+9wkSB+C
P3IhcEB7g7T31M9yxaholfJmoLPcL0adeEuZKfYSytsfG10bMii17tweM/X5NlFW
1cVOdp2zHSM/YSQPCHNjPqTl1PBCPnB0kn4GCIr9kk+ld04tALW8F2RPncNNOfX/
PCJ2g/DaOnabcU0PmTj/Dy5EbLuYnLGKzCfBTYjw32Zb1EIOMUwL908qNPEXC0GW
X9aN0XLjZxH2qCK5Z6SD/1qON7wIHBTQI9uULSeV7be00SMTst6n4NkvE14qAWO/
h3GgJgA2tF2i1IT7pZWHLpKFqcNc2kfeHcu4KsOukY4qa5hvXnCkvvwRZBREaZgh
Kxa23+cmMJyDIZRZaMuVtI1M75IzKr3vnJOVp4O352l0wZplcaUxw6zjgQg4DgqY
f8dU+Mwa86NBCzUzJCfJLB6nYkcBS27Mi0yTnEWzszgaZUv1fMEXLpuGNimqLRir
rERTWOi5Wsqm8qPx8Xiwh+ARt18kqWe6+W0EPFCx/g2jUahbHD/i+B2xGR7pErwP
fTJO2ZgTBX36unALgVqZ9+iQNWaU0vgqqepEYsgiJ8f511bDcP/XX6HonNHfQTWH
yPYElQomvXbO6uhcGgwEgqEP0uDfilZacRWN4V1yeK8k8sEMwpI3H9d5+EPT13dU
EdTIqP4AngNzvZFQHk74bvj2eBfXpwQF+kI3gaH/TGB08Ot6PfuKUAZ6jlA24KCX
Sc9/19TOa7zoHGCReEmANhFbvMkqVTWVbrQ4+tGue9j6AVJUvyUKV+spNK7pBqlZ
XWA1pFGqISa/fu4ES6O/a2Z8XM8+/nJlsG1oo2FlOfqNwl2BX+C0slYujdm70agE
Pasw4mFi3DJoAGkj0EA8GfGQdmOKPcXEDPTSeNKuu4h4I1TwG+6QxzxJv0tLvN3i
bz2WIeX/nnh5vOGEUKeBI2LJ5Or8vvrWe6NTtV27u7VBjDZm3TjkJnh7tADB2WQ+
wEdowY8z0d0Ouo/pZOREI9iu7Hop60piIZ8nLNHBSD0nrxYtGpb0YEs/o2ZTyA4B
i47J02YbYqqNPj98rqaOGUN41MHrVrS9KC1i+JCi8QvAxg48T6jmqQ1w6rs15SGY
X2OwdwblOCoXQoIcyeLjoMvjS6M5vep4Tqdvm8JlK/B4F4nT4LOGpTH9oiJBFgQ5
dCyt0IhG/5rOXkc+llq4ZglQCmAdMfeFt++NoujZEMgqquUCQlSICBaqYJIglbj0
mP/BAXSp5M+aOV4r8n8APcAwwG9Zx+6eZYASAOstkT5dh6k2jiGDzKUDxKVfTMln
vcKw/G/7dVp39Gb5HCWT+WWZaeMH3JDm5EEpv3ZL1B6M0UwKb3aZOJhyTP+0hbBm
8iAFoq5sYCFtzJLRyFsuHypiKJXLSdHhcUD1kUM140vZsBw+a6mu5JuzPBRxrmbQ
9Yk7uIuMFqVps5J/E5sOffMxJa0Swl14DaudyHYZqg38V2oJoPz/8Zp2tcO9aJuT
uEQwlk6kdpOgPCtSb8tkQoWlEIfbgxdYoNLgaG4FrttxAT3MP2GhQizLRTCekx3k
pPMjootMPzCdAoBqpxu1ojpOOzPfs/MDcVTzv90AytFYlJj1TwvsSOxqTWQkvit5
jLpDxkPJfNrUcCKK+vNlqkzo4wmPVr6WWvYkXpq+zNayNRi1kKf0o+7fJ3dtvBWQ
zMROhHwGmxk05uCUQsEeXXBwQWKg/kC7NKpaS0beA5E1kMP3KLMaX3fkAnsfvfd8
V+dArle2riR2b0F6pH2QI5nCqj17YNJXUgkds5hcuIt44zsl78Q3cs3fCodTzhTM
Qc68ERM1JSWeRyDjO5+jdo+81fVpwgIRRQKIvjVkw0KGdRWr7I9//CwEABAhF23I
`protect END_PROTECTED
