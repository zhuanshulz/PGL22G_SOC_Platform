`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v3sf/iSlilgzUHB2F5LxAidcqt3ZPCfy0hqzT9kfSaB1EtTEMRLjPZXerKIbUDnI
OGp1+kgCNAKCSI3LOr4RktU0t/7KM/fveyKuccf8O3zOqCKz0jQKfk5romtlkn5c
3doifZi0WkuRmM7hdkBv4G90KGkTJ8odm1jbGSwLgtbNCmCmT0+c5QLw2D1F4ovn
hc/xjB2yoFrNzNH3ayto161OuRSFw/24kPAJ0wo8cQkBexMflTaMjVNWdgcjesn5
pvH0vyoNlm0BB1P+ysl3NaFroa6rARM9IxHsuAjQ6xpS1JWlYAkl4iZhgAej9ELg
JvarOc5BlmWdp3m8GWpehUDMkZ0xhgT0krEqGW5NdGOjCpFhMjyhpBD7FTSuDpuD
B/jHs2BafaZhX9NtnxGHUQ==
`protect END_PROTECTED
