`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ks58Kk4GoOJKuqnoozEQCzZPr0a2+ARSIFlfTH414laxgyze3KAd288PKYhbHfPC
mkSDXikssjytszetrNigFiTgW1wusk03Gi7Pn/+t8UvICm+2dD7sdL7usxHnxHmi
HZSIuycAbvDzZJ+M8kPja0xKm6S2bfiwSblD3XLgDz3J9RZWVx4ve5JgGs0ENgqH
c9OhN2NqQPhBZNPXt7jEHImXQAFltrc3aSsy1g5RoG0Sq3ZJKp5y3/spJ+xmjeHT
RkmLgMZoGkwctAEWxj5kiAtfMxSxpkch2gPnCn9vHEfND494tu8NcMwdZjTMxTuD
kkM8c+P04pTDpw4ZmFR5lST0P5vHJJisTk89kzOjOVAOmUcZB+r2XPuoetsK4ak6
lfCZ1aakEWucALNPXLn4CFXzhJpghHv/AeLWN/bd56wk73ed8XLkwMpsl5zNuj6f
ZADSy9mE6uO7rnpcdS8V1hilqopsNL1N5yRFupTfs+iZpCkSQdUxWZ6kQJ+YJXh4
l9y2ewCIbhTlxT93k94H8Ug916JYNn2SMEQOA/q1WyN4TJBBTyH6o27X+cj3V602
ifuOLVVWFoZBov7ux8PT9U1Wtu9z9Elglg9m2kckbvOPY+7v0h5KWLpB03vE+06l
/typr6/lxLOM/nQW4kYk9C3/q8oRkYZ0XidWPEENPbmRwrjCxSp4ffeZQQdmT6LZ
2ZXAlUaEaiBbVxclBqmIttKG996SnNG6f4n5RUnaLGVLCjXFGfHNJoPQmfnRIdfz
tCHItzpyhotx7+qCY6HoPH/r91BwZpwIvIpaITCp+840505c1xvKSM8HSkAlzFZp
CZyqNm5alE981vi/75lgAvOzXIl0rAtWiqNftcjHbD2ZF1t9rE2c6nQtJJZ4tTPY
f4un2SPjLYyrInofSNz6k8SfnGKObHgjQdKfRxKwUyNxRVSho391swF2yQ48tNR8
2FRPz4tDEx3oOd+sdPBclMyudR2youmLzLduBf3c0ffJHCZAqU+DloyqVuXANywz
eGgrYEHuYs6fCpStGPGN8wJvIpkmyL6u4qIfhm6jUX9r4u+nqultCGe/tvUimFpF
NkB7Ym6qI2GMZnZCJngD1I8KV0ttkQdQIzh8Tf8Qxk9hRMi7ibNq1pLHwP8VLLh4
pYVbTjo+1+AdqB0/5bBfDzbM8YLfndS/0C+0rNeS24oCrxSic6cKyG8qZkDTqVn6
5MCVisCOsDus6H3sfZrdzjnsU+FABfFvh6dfK7Fk59/CFwbIMD1Sm4XARn/Nruh0
U5ONtV8VkEDlw3eXBRP0EFrRWwxjiZ6Ob0rjNDpTLiSUZ4BhdaRt7kn3Tn/1bc+F
LnicqQPE+/f2ANi43dHt4fBqwP6KWZ8o28L87sDB++PMZepamMYNZkH2y/cgN1JB
VD4YI9Or4umfFxFjDhh1wl0bu0Vv3j+U4J5u+sBbSNApbdFw3Gp/pjsMbZ+wnmYH
4AAj/NiwTVx7q/O+K7mXRKtRf9wcd0UiWUcwmgYPNkrku7rtNKqdV8DL06PxFRIY
LqjJ/IJdV13kIA9iD0Gxj6JprXitEiAEFh+X/g+0jrRGM//y2HnGj6terUKSPyDq
Bu291oB4Q5AMpsqV6pot4E14fXh/KZ6AOyIYtvzSw4vwPSjk2/qE7zrIcmN07Svc
yAg/4XP1T359qvfE2/Sj7MTzXoN8rT8oqjGBGV2PvgQ3WPRNI+AE2BG5q8CEoaPj
eI5hag5kEgFqM80LkiPzcGGuoqoKuCQKNvx6FIm2V1GOdrgqtTB19bzIAQSJChox
r1+H5MS10Dq4epY2O93dwbZ772HF//RIVXTaNLvXIEaU+mMpLKxp6wPUuyrmGasA
PWj0p2/Wpzy7aDh+rxQDl4Pf0gASM1S0dJJexKMGuilCxwN8P5f3m/28YBpYC07D
fopyY1NSad1v9hwKBT2mE5qHSzJOrOn7K9oembtMTCrdxR0bnTOdxg8IqJZVXb1Z
aTgAFjYotIQVaev64bQD60KBwhVcAjl0KHXqd+PECGC6j6CJ6/GG6nTL3eILhik2
O62sI9RrIXqZYsbFo96rc3AO06j0SQ6TpEwsiC5GoUFt00s2y5B9WV3UGM7WBar4
kwDzkI45kCknLjtJjmlBkjSVx0aGkD2V78xaCXKM+ADF/cj6VFdavby/dP9tLYn5
znP9j9+kXR2zhFNAVwiI93IDYvywjEGFhbTqnfkxF1smWQKk8yrOcjCa7/mIjF9+
rJtp7sEYGBd8NyaPkYT/dkUzvDEJwyBnMlM2Mt8gr0eBDXTfxKhOBR7Y5Tq2QkP9
eOKOBKjED/+XWESp6NryX79jYm4IzPmuErvczzRkRSf+4n2UIUz3hHfMJ/UWgZX8
s6P9/2AS2Qd+TItYR3C918m296FMOyVBdwdbQGU5rReNbCPEEWxyc+AHlyw2KnfC
vsugxrRivhlRYr+6eNNhNAuiqZaZbJPf9J2s/UxQWpl92fnw5OxJ5VIAeBKJwOqX
Uwf27xvIZYx8BXkLV8e5pIqS1DnntDUnwjETf78lbT1+mGfu1feaXI7SWnP5jK20
y958iGySI+Jkl1iYil6mFqEIEotij0VFteikAs6H9R6IelU8GQeBNFgtqete3LUP
+ujqMo0TsNIMQ+8/c2IoFf7pu96H88ca68nCY77SMT9GOdgJqz4AxK3rvi7iNzg/
o3TK8gjWPaigtgb2NdEeHtTVUYIbO9g5/UcGX2g8Yg12XqW9oU4CLPwCJVre0Hz6
jCyaUR1MeDwId4LJSyHNUsM11UFzamhGEynEn1JyjqaqBwtvz652rSRargJU1qVF
OQod0B5fMhR6Q6a69KgaV0FFoh55AbHzkg2VkAJm9WzGHU2jeiwBphwb9t84F2TM
n/gdQBlXQZSXU2jwwbJBiPG+NRTejIK22bfV5Cweww9v+wCo0mgLIGgB0WOnXHQF
9CSCPN4SHxVsnPE1KVsns3Yv1nOkH3MpOukWIB50i/3h+okD3rws79ht4p4YZYHQ
S92w8M264NeCUQima3kJ0J0QOrqTJOhazyztMx9dGa5kMD8WbjGt4s8m/pOmMlvv
tAxxuneLYvtatx9rskHlROmnFSt8yNhvP2v+9YtMXEwggrSBXpRxmxu3HV8/Dyst
ODInS9qDWAb+lnmiUyTkd1hrv2RI5buyx8CBR95tkjxkfrZYC5Uh2qiwBBT0npkh
DKOEVAKYSxPQ6yVobSbINqp8yinPzIFpgRN4sQFxsKbpJy8ikyYSAL6cNP/gIBW3
9JuIcpxpWBxz4VNXIiSWzfbb1yxdSLiMiLgfTbX0krDmlk97bPWEsSEMq1bjHioi
Pkfpijfc/R2yEjcDRqFIhsTiP8bJxRNEMfvhK3U7dZ0NHahNhuMGyJ6C6EQbytcC
3H8x3N4wn6fExBYKcdf8SFZOXqNzcQ6mbxFCYBOnt3/S/ikBKZGfveQS5HXKNBfD
X9aUE+7SCyBGcRqpwRjl0XPL0ePkNPL2/tFV2Adk76GULDYcWHUeyXeqP9v5hj43
exUDm9u9SwWBOjDl6PBuFH3cr/NrIGx9XduHOVdgBkGbk/VXqSdZKt+AsD2STlzh
IZJ81SpnfyIMbTZjCGWgjZ3GUNp2mmZDQ5cSA8pMWePBfjYnbFmusHJ3ppKq7Adw
0ZatUm0HPAQrCtPfqrEmE4HZeKwkZnB6o6OgxbR6CttNiRSuoFJ9NPcs5nXvNAjH
incqzynoI4DJMCsvCQ2iGaYjTNAt+Zt3JNrIfwasPZJyBoTvdeTYDxs6fd0ESavj
hfe/xbPG/egp4DFnOyoTvObhpaLK12ytbLIMpYmo/PTHCnprZB1Iu0tWAHP6mpzL
fsviNC9SpCI4dIl72np2U2n8CNjedYLKDiKPtb852eOBO2HLmS6zLeYs9VPrI2L/
pXy3jWTrzVX9FZXqQFBk7LTjCYnMbNDqCMxWBA65w4clqPeX6ZKIXOUz1Umh5tCS
l2gNZ1USoDs1kot7n33Z0NO6hvP81x6JzmFTZx4lzPzNhoojbEvvVC3MVjbivfTy
2oQdhaUtcNUDgfpYL3yG5KKk7FnbXA5l43QELmS6bpZkCctwf+nxqnrNgoO+aDB1
5kSLtHxt0608gICtAt+HkxCkf4o35SGDOnEH76ar+fRf6ZQhtmV1lXtU1iRQUiek
GhZOtXY6YR0ymBpq0HuaewTmLno9WHRDJcCBx41tD2bEI+2hEgSTWppFCScSvUg6
XluW6zCpZ1YWETxP2QL41J0Lzd2k1kOsH4oQWl5a3Z6sfdy+AvT6BIWPHD2bvwaZ
3UYs4A3eU7vl2+jcYg/VQkMWzEWR1Gy1kYBPQx1T6w8RsIZ4eBOPpz5unCqGJWnp
NK8vixIHygX8TincFRAGX1VsI5CyDnVe+yDPDx3Sz2ziFjwJ4AMp6JZfJiCQzTF+
BNWElQzMe3v3GAC7oZGhjhH3pV0jsX48qLdzhLs4RY02KJzQfrlYsnfedLqcu3XE
vwWxEab4V6N15HcDfaxhO0MxfINv9TW+KB83FrYyPB7fykCRDbZfnTLtpfZXXgjg
EW5q3Y6LoIvuQ8v88BPFKf1fgf4BaCgJx6qq4CLvhnKqyKfKTPNfATG+NXX0i23y
9+fxLejdxrO6UunpISN/2EigkSurvgxmqFH7+LDDSOxqf925ApqDLvlFtpd5vYq6
Z/Alp0NHYH+BE52EKSVHobjgLxdTY4YOfjdgfVex0vn62W9JIZKSokxhCWqOLdXX
6aR0YY8ZTwuyPIqRD7aqVqY4LU2hNUHCw/Y5NSlLEd1za9hWKgfn6Y+mmlZ6qPMq
BXCYcn6bBkcmcDMKqO3dlcBCw6MgXlW383ZxHU4pzEbkhmyBD32+ONUmQy+4lQ1v
QWXEPZyGx3+N2ucSILhlwDjIBU9Kj6l7EdujuRU8P/GAdvmxFto2x4GScZQ3nHLE
r+BsNvTq6wZ0OIrUn9EB/1YqMElQHG7kuc5U5mouxvFQbljj8HpSMz9f2L6vVPbo
RAqnUvPXPYXcaF0VnOZ/KRcECd983cudF3vn0AplQHI+DrV9XUo/N/Ak7wJVtSt1
YbTZQwmhm+DyyhV+tLPasAjxpbu7119tgdUwMu/vVugHPTJ3RVec77QrH8YlTNDo
vSx21kVbO8u3JFT+Gv2VdjPEkbx1qQxbRyU/WpgA9FrOU1n22nfWv5cf+RetAZhK
cjXKMVTB3rXIj/cjq17lVLDpE7hIJSaLTb9+DGJFwuJvaftl1B246EM5rjPRCAzy
ttJLetqpJy//N+QsVh0Tz69aeNOmGzeA3t2ayVjnEurrdaFvCR+x6khAF+DoqS+J
D8R4TZGdCw9Azp6ykqAsEqtvzXmnuIWTwI6h7/NSxs3D1fOFYiddU94aEAB9ua9p
KoRTQieNpxOZ1Fpn4NYUTeHWopoYFsM1bK9iGM18f0rMHHbFC7InWvphECwOQk32
iSlhFwiAhaWESSCS2P+ZXR5zF/8exw9B3/6zIBMDEH1X8i9NleFmVrl7PKEG/Byf
4pG5/6tbhP21CrMH2GUMmyUu56B2ZB8hyfZJBa2hzjVkC4R1ZZscrxX09kDFrF/x
me3J1TKC5+2CzX5UghVZq+btNlKeQySdO+FNNr6xj/eNzmjH32x7V6jDu0z7+7aJ
rD7YTu5PENM887x8W0iwTUUcqDIH9YssRUj0bpfQS1+K7xVF5l031fX6xXD8/ay7
UBHGZpERuWLq2ScBn5W9Q1igahWEwlVepfxW/MD+728RAwdr/XNFErbrubqVhXIi
GDLlIgYkeUFpPDh3fnM9VtwjjXIACcAFKb5JcSznHnqvg8B62MmHChs6NsCfZfWj
R2BjDY1Xeoy9M8wl5dm06hJMEKYWnzphNPMXXVooGwLLnSgfBa2G9Oa9T+q+i3er
FRXA/xnzWEwJyjuBhv1udsZjQ3Lb739VL2erlN6rPhgnQtWJdQg7utlEMkbtO2Fy
FNP5QyN5q54PeuL/yP7IFkfD8iY3TpA4K+wM0qKON3qMql4sa5BJsI6Iu3I619Vv
hy8+RQl3rjCjGb0NkotbQH8T+sT/Yo/VClAdr4jYWNKk04zEykfsPneu5nUPzNTQ
WGmihfCnozANBhD1FhLY3tpGp5QAeM6x56HoOw/9FRUlPzXYWWTvY7r5Q3Nc058h
90RAT6MBD1yMhtJlHRU9lpx4gk0/Mf9Yw1xxPXIrD28yL9yBRoNV3IYXBTdJSrN7
YAg+QOfUsu5elSL3NJiS/l58YbQkWaSoJgvWVGIWXh/X73sBjpm9V9Lk9QHHURD4
KW0s0kODpaLoIeZqmGEEyUUJJxZnJ8SAsHLyxw81xtd//z+qOPtckRgL4OlM52Tc
a+GJ2cQ0bOx5e2BfDnYlDvawGkwQSArslAzH70pAsEDyQf3jtOUurxTVGpeQlc8x
/LBXhZpdCRE0AYlr/XK8jC0gOjKhgDjKH5G3FBUoykR/5Oz0Ott8WbtO7RryJVxV
WYFdpl0LtMmk6hwdptFVnfeBQFmj2hknFgVQl6hoJN2vUBUSL8p3j1y3azEv9dMI
KLHRJ6BmIGvoNtP4/WZMe1+O/N6HBv24zVCYxYoryY7uBTs2IUdQfnHZaZZKdWyF
IqWvSYJS/QF0xZ4mchamVFh9Uv7Vj4asUJb+1xhZuRKk6YNCBa+UUVf6mx1OB9Kv
a3tNgQmQOhy9Ljz1wMjtrjoZjU6qIAhIZteplXvUOB+bvJR4+vBp4B6846rhXITG
zLdokagQluE1gN9FBBh5Vbr/YXHacB58Disb9aTdh40ANlsctREKpstfy2p194XI
G5T7uLSV94dgiBD0cuJWHzWCIkn5hqvH1/c8xRypPogVPNaAV4c/2Jg0D1BVAxZw
ph46Fq5o6/mAsbuUDWVh8H/pv1HqXY2i6QpS6oPYqupXyjWZCiW9dx99/i7520Gc
5tHsnA3XqtET9VcU0iT72eKSREeY9YEQ958xJddURu7mlKxyxoW1B4lIeLJOnJfb
oMCxP53vImowmC28TrS2OEpS06en6+BoPS+O7F0zU7Kt39otcfeC0QezrUB/RQfQ
quepljUt5qbot4Mb1IqJ94wvQQJZMXogxPae2ZfdpdERGM4YbFL1TFg7HePBWsq3
+hI6V90DJoiCACdTRv5iAV5aNKxWpRAQErEPJ5P1YCmZZWc8GB8G+XNtfLzK2HyD
OwH0BYAfgZ71G9o/DA6VK2wp/68wdY04fSmiop6mATXSXphyRV3wcclhj+Sg4Cv+
CxoVf1NQRJMbTg8g7Njw0pk5RuPFA9eb2N9wxzNtPY2ImFpjBEc/GExs6cnAfqio
sS8cFNwstq1/eVb8XXngye7Biu8ZYpdw3WbxsewR9xPYD2GUbzoItO1Tx7Ab/rAo
uj5aqwB1HxO8Prl4d+C67n9f2ljyw0sDRxzEwxZUgZdtAchBD2shO+RpAEAP4uxT
x9CWtaooC1KQuMsIwLf7woR6YhyQhPp37ipN7dYs/GZek+ZiNW19vzFBei6XcWJa
6y6sB3ouhLPXHqFw7S2luUlCrn0TemRd+VloFZFOXUCalUBX2RQN/4znJ4r7dmEM
+yS4+zNaXxa3Caqats/Va8PwAEwCPxzcWI+aEdZjjjdmkfOgClJlNndtQBzB73IS
L644R4SmxpC9hfc4YiIZq/45h1Lq0JeNFvU5ViffmEMjvcdnz3PJRqlXYkR42YzX
Go7OvmSp7yXqNYD1mbnCAoVh5k2DDVYvoxkdVz1X0IcfCigwARfjvOZIr61WpK4f
f7jOdIcYjGIn0gPJtoBKu+3zvwf8I1kOiyWAhC8+Sg9x1QqDcprikW6Ls1ofBDr0
DhaUDXRH1xTucZBgIboUgZainqWmhE+N232UUCwlFUyidPv8ZwuXPFobQ9lYZpCx
Fzb+L9VxsFbg1/Eeio3i9QtfusPaL3iqE22GlXCA3av+wgyRLuK8kZ+w8zIYbPYC
lM6XpOnqRzU9xubwMftyuMrQKUOGs32WG73LAvj0nQ+nTxPcaEpfVSDt8r6Mqk2J
HblSG7dcIKIioZ055FsX0JUvdiR9JvnS9edkNRq30mgBntCnZMgSesGOmMRwsH3I
6RYMHVRg6Eu6nAowD10aSOqnj07iF7xOFGsoS1PDJayBNPBJnIT3SBOGDNL+jXY7
DWNQi+rVH40lsBV5E9kBqaBr/Gch77ykmaWphQLb5BHGuBKLF1TdZah2902Y/lA1
oaNytNXX+hDGnC3RpXw76tcP23Wb5jWQKNk+yTufwkz+MSJchL8ePpjWT/kyhP6K
osn9haDKL+WKcZvM1aF1L24aZJ2dUGYWQwIOfPDq+6tASLhd3kU+YMq5ECuOMBlW
rhawKIJOyH3GmAWzrV3gOc5rZwfVillf9Puj+XPw41hCDtrDkaqa92HyFX0SeBgA
scs8efT0Gdc3/pXvtXlLgNd61YlcAv6I8/lpM6jjhvb0Q+EfxFUJF+flJvd0Fd9V
+Dn8nvUhTzGmj7sUjI5iIPUluIBOyR7MNIeFecRMr8WuY0BF9y70/vvEecJtcATF
ZK1C7mLA0yO+ljw0PzFqVpOSAe/7Hwjy9pDLYeHnHucxI8wnYUPDUkj3muwtSxtV
vUF2bZppK0Excr74+/yXvl0WLU8RCMMaQ6EPXSCfshrF+SlrtYmMDJmvNaSK0ReS
fNnQBVYfsHPirGwcLVCp931kMGrO6BAx2lkP4xE+7aycgFBWZjgbe5/uviGFZ/dS
ghX3NseQAEVroI9Zs85+wMGBVwXnk5zbugcvKdRWWkrv0ki4jgdIr3KEpMniCnnW
U8gGH49lSd2lbT1qSd8YodOJmHmvw8zVebcqP+5Fixp9KzvcPVG7QOfMaLrGE7r6
U7jJcXlqUhpJQCsKRWqQd8LXTcqeTCGl6sSYkNfi9Z/jwiVR6aqNL/VNBK9w3vaH
tePR0zcKdTdvukAcjtYMkwKA5G5oXMHPVuwkwkdeob3CKNKcq+YiJ71mg8Z67RBY
tQkQS+UX7zotnn+THL+/HUnJyx4dHjJxYTCyEaS8fB7jl69k4IzAvLhiVwNOh0P5
uVQd0WXj66V+k0d4MvHvydKrxdIVQM6GVErCrUxszgvTrsy9Z5crXjFru9yGas5t
pgxZb2hbwl7t2g14fhHf7neDP45M30oSBN3ghxFn8pWLFNUh9l08d+aNmjzi65JX
OHIrXtfZ43kT1THQOh3tZe0CKM+SbI5Gozaum8xAeWgqG5HOoWLKhTW7lux/oDVk
Nm2RS/ZuzhNrHQ1aUci2/MF9bosZsm2/Aa3Anc82WuKD669eAzFHv4xGVo+OJOhI
NO9N1Y5B6Be04m+R/zVNP4EYCijUbmYwd5tb/SYN0Zabq/v9q38XJQQDkMEHNL5u
5jprjT2x+h0O0lm4bVjFpmvBaYuA+FgJJ4bE1fglqb/5zwM0f5M8cLd5CxRRf23r
1g7OSOyzjJhZaev+C5VlSyGF8Aws4ycG2MbANXIWRLnwu0ljrkhCVpD/TO45kCPi
GYNKfWjul87EY9z7dPMyco4HBX4iY1rwFA+WWERR7h18enUrDUOpITVNuIuqIxVX
w4/BFfeweveT+cQrBgDe/HHSHHPWGnfCQKrm3XrJA0txBgzT5jdeN/0kmwWXJLn3
IASZyVMUuzsNoDgFKk9ebf/iodW375bPXkZHbQ0VvaNMl/PpRTC1zpuDfDQcfph7
uvVB8wNiJBwbc+U9MBiwZHeXnloM7JygphxLHo/bZj6I1AIzHrmlZxLjbPv7D8eV
5Fm4g7n6KFrGdGVJRa17VTbVvHdr3WVqTuv/7ABEopJ6BT2tATuB2qAEzNzYJDVT
QtdtoDHqY0r0jCNwKdaBfCG6iQmc5xMiQTWfMYT7XhSZerRIlNFy4er6sqLPIFH/
O7k3aZTYVBllKy/s/s9ORpiYr7UhvNOevmtFFx89T1skxSs58OxAwneL+tr8fowh
wlZhiKzE3oAamign8jfNzblYeWZH2xO04NaAHDrS08HQljOa0YULLCk54GlKFyPj
aVxE2ct+/rc6pzJnngiAakd1exCe91wIaXPCaAD357B2A8AcEPsatmDLv5aBmEen
Jl8fxX7/QHyE6FI7Xe9LLriVkgBvy3bgShKt7oex5wzLZyMGIHBWFoCyhDDZNZWx
ZnVzxIBUNBzcbocLxHVPWoANdufXs4iJVXNerYCCAZYH6A1R34wb5ftNBx9JD8XQ
IcA45nX6y3fjuH+2fukytHEBkuk9hgmq3j/PoiA7edYt7yguJRp8OAZYvD1gnPfO
3NQc8zyo7QYiaQlTXao7plIjP3B1D6meukcqeO6xv7ttwS/4UrXP4H0tvqC2oemp
iA9Uwr1Da9TARmX0GHRNDZIh/Gh3uzVztlic0JDA0+M1IiXlRVcSWkQp73W9sL/u
N7EMp5gSpPoDAw0VT4IXqk1icKe9pjxxkKyHSkC9neFd2G3HxwiqdugQT66+pxIA
RuSGM2kAu6cKUFNMfwtEa+a4hnUkdyo5AAMa7HkI+eUJker0F2KabiitV0ARZRh0
R823XqppLE9IGggMQ+mOSnq8lEsBZ1QpQ7Qc4mUdvmPnLEVIWqX7aofG7TgJPnO/
dcC8/T4m0tlbFyjmMui0gI209v89wC+TCcsdvtmxTLlzliyLf+HEqKZpjaCJzr8s
a3CujKHNQdiUwt5ASeOC/nxcKn6zSk1mWJHePNC+hultqQa7SHgRenWTSASYk5wt
cddlnpjT5E3WOVTwJWVgPQ5qPVcYmVSuYTYJqyXF+7K8AJelTJz7+Zxgov5sPHF0
g5+MzWU51SIuIhDgXMsLM3yFMIsm+zYtw9uHBRmG+QGQq7E7IGmzz2iFn3xfnZa9
tFGBNXY770ddO3tip+pQ77f78z3MX8PgOY9KeV7e6jAE4mzihnlLMvRbwu7rBLM9
EIXZj3mrYYY0GGqJaivPWLaUpfIPyv5PRaEnVw88ziOfWYLvx0sdM31JWKhfMD8I
LgVbp2oc83KdwV0lWtR9sq7jBxDtUg5GJeSAjNOFrwYYM9/wyWJBhnkARFybBPk7
1FjPO8vG+OPR0CJIPS9oloKDqg6SuG9CS8BDZqWH+DdBP7ayVzwVR/MTjCTghoSO
frzGQI/THHHo/LyxwIgYDKKWZ1eU6rNrU1pEnPrGX/COFA82YLmc8UFnLv8+C2DA
P054k1Mi+8xsOq+s7fph40wtqkzwRQ7iR71l2EQlpdEUKNbS0cIrDwVzKzpSNVFQ
/grEOdTC+5pFPV8gdQ+H2LwcaapbEqXHo+YyFPH1ftQHFUmAkuq2c6xyi1r+18Cm
XT+rK1OYDATcjQ/OWlCMfwPR73hVA9rYe1g7AOZ3AdkrTJqf0wxmgAUzLK3y9r1/
hyobRJYe5c2yLOsx+wmd4mZr9W6CLSY7fuIX9JbUcmvfsghQTS/gl7iy90byDU52
1ytBTdw8ZBC8RREdQbXQ9XykyIKAiPCR5/EBAiC0+Q2T0JkPYPziEW86OID6rU9c
XJLtXXdak7YV5ujEsgWmZL1whyUXIVIu8Yv9IjI/tQCOzfssqHV6BV+7KLo0+67W
XE1ie2eONMzucrb3CX1ReecDWR/mdc5Ftnxf9mvyKg70Y8N3EEFbpDUO4rgSjzNK
yyIM7/gps7gxxA5WkVrcbxpwONQf562rVX7V+n72FeVeJUdElB+3xa87YxzNKOQz
7SsNxcDNCv/KHneW4XTkDcMz1BjcSv8FwWWTsfLhW5upr4yH4T7olJ95B9l2B/Es
BAhI4eFle10iCx5+siStmthPTJ2kT2EOpXXGatk9XI4GaKj+HRcVejcj0hc06IVU
lQ+WVWJwxyiFr7b4VEsrl/LwjcsHYIEOUE169DW1fL1D7dM+1zUm09+eVRU4dvR8
LV4OEqXacwWnptlt8k/fKH7VwxYJ72SO9bcuG8mBDEy88IP36KWdUErcVkPKC3I3
qzTczxpL9yaKLakcxUNptzg4TczKLSAE0CohhpUsznAubOTAVMO4TAYMdhngnwzw
KAeAQ3gw0ty0sXJeM9trl7z7ppMQxpc3oSoC77werVY2USlAD2rsaktxBZ36zOx8
iLTkE7pQaSP9doqqKUOiXKiuQI1CABKn3nlbvnIKe+dr88EvdYTHgiYHnKl8Ubjc
xA4EvXODq+NbTbq4oxW5QA7xDTNinn73R4PIfp1ElBRKotSSn85/+Bjot9ZppMdN
z3YvfjZumZMteLOPNwuqhtJqiK+WGuKpatlTnzDa+M8d4McxJBr+JUD68sEcZOt9
NDM1+x0kNb3BjmFRL4emWqlS92COIslcJeJ/SEEurAGeHhCb8Xr1aBhfXau134N8
ycepQhkSE13d2yrQ+XgKOjS+mpgHWOeygqxiLvlhWirKMT93KUPNpaHX83BHHJee
g0yS1XZRxRG9gMQ0esmfHaGjhE5xxfDyhzDggUwcuIYKoOXzouCWfH94g+09j5PY
Ej+oa2Lrmjo7IW8KEeqFeoAzEg9sJIwqfVzWeIFpenjWxmbX4Fedice0h/UowYVv
2pnGhUseGaUwmNcSiTfm5OZTWjQFV++N7pu//GhlKe5V9zON45y/QhSquRZEbZ1f
ie2Lp7JfwbG3lmoz11AFg2s0V20rqnLZvgqq7+oTrM6moyMSN/9l40cx0l5/Kfow
YjttPbPXdXznbo4rJ4rxAp86AKPA4xlXEG6B3Ryhr3p9jE/eUoGoV+M3ATYorn5N
Thz9eRuhsQDMuSBquqZ2rqbSHIMBRwyld235yFQo7jUR4+J/pb+KjzrTfbclHa7J
nSK7F4Bys+2MwbRZ6xIoXl4GyeRrtrCC/c+vFcp3ZRchtV8PNFWpZa1/CnvyKdZU
80PvsRRJCvGEuCKX/Go0InUf3E3KF2HlIc5K4M1q0apfQGMHiEH3lg7CfsX7DCdg
N8jK//EuigQoquusATpLQfq7oKAaomqOd+d1BDXeqrWwaB7WPKtIdvkWZuXY9JYm
flcUDECXeq0vIca6OGphLkbabwuuRBh2t6g1fwvtu/zpUaWcSl3oagOaToQKanh7
VZaQIt2zzDbW3iGbVG6saGUyTugXD9ywOnc0SOLNYA9R/rTGGWBuPPRYZbjiNbv9
cE75Cllkow8tIDVMO28nMg0WzFcuJct7mYDrJJP+1dnZAL3x5WwQvxUfnZfLxNkM
MHuhmbPiQuN6DxbJr2E8+tnle2x2yP/01YUhdnhHP0EQNdmFbIBWFeWEsJJ72IMu
TF0U5nQv1KuDTrpBvxghLvj0egBjUTxmxkZObmoTXOt9PWNsbWHQ5Xeu0KyaMZ3q
bu/DPO6OVH7SfKkfkPgkemGzd4MnTQzUgOKvSP+uwNb3z09ddABsMFtV8dC5u3jJ
aRjrFhUkv7pAToSiNYQloPVFwcavymAJOj5rRt95T7LDuBDvayyi0NU+x5IfPhzu
5bwhFAJ8WenAUkZnqmnQrng4s06d+tg2oJTjxtW9bndaCJlsmHUZlgF06UVaQZhT
HH5JRuSqiIgjL/0lLV1HFl1joG8SHwggWCSXqAdc+zdCq62SWUXvYLlPZx/XOB8x
YYTcwRxXOEdLgC6bw/edDxUx/4SM6KxKpPbjB474S37tymH5/M1DjWnRlQcZtIpy
b2Y5mQriOBRUBZfwQ39Q8O3V+MeLSTTZFQNfvWZlQ5y7HREh/yt+QgPcUcvCKmCK
+EZi8t9SoEzfOpOZIMmieAtfwvirXPnmRzPgSjrzI/Jqm0l513JayESwhsMFFblS
en/wu0vu+qhRxDXJ1sdr383BZFE+MOmCfkzUga0ypVLuTx4ajWNrpM2csUHgu/UG
t2S9ZfVAX0aIkNHMq/RGrhX2BGAfabI0b9rIcNjcjO75kMcr+QnRXzFRtDZ6fFAV
J2wJMIqOEfSeS4hC2l2qzOywaKrmnQgT/m1voV8Rc/0=
`protect END_PROTECTED
