`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkRVHaVlYRu6K2lqI8UgjINIpgmtLA3C14UZq7PBHFoytFYtvHT5lHSjTBLSpO7C
Jlt4/V9GrslklPwjG3ClGltX8M7yqhqhW10aRIzOtzDIchB9/92DYuVL6xLd3xS5
ukCgJsPgpzVs27EEW/12Jmpzni4QClMy7Q4aNejCcv3PqhD1Vh5RjAe4PQHWfCFh
iaJs7qtZE6ymh5RQ1Dabyhk3KXwEGcrQevQZtpIyWvc96NUgZrmsI3U7KM4JHt6z
IkbanDyT8IWRdqIvCSfezSgmtoonjuLDDzEIfLrcmttu6dAM4T7+EWMLfhHy6VSE
/3FWAcnulacCr9s3xZwBYKZBrllQFi9IzaxwwqDcY0MA8UnmDMedfYPkq64IVBBt
iAfm1Egydygfv2Vt7Pc37xZAHBUNs4bWE3/1vr+flC0QQ5v3j7GIi/t5SWUaxr7/
w4SzGAG5oSJisxA29EWYwXdO1AFwh5CCEYjWgmJUH69EddtBIbSItEjd6lo2dcgc
74bIvKRPaFsDh451lZbgbr1on9T3pY+JDtmoBdrN6XxsG2/baGjPfdOL891rFEes
2fFDh3gp4SDubw6WgxyEPTKvtb4tqNPfod2WPv1Zn8jr0YojRjMa+0G9CZo5hXNv
j8/LXNuhpw6JNGrjJDKJGWWNipkANOfS8GsY1mb1JSmz27+jfkDn4/piPhNixqXD
OLmMZX9xnFhXDa1HGlqOUPL3pgiPOwSXas9smo6G6MnjsIXFFrxrXHpnLklpju2f
LH/QqtRcyHshUlyjqpr0FJ2bhwOGrPVxMj9vE6BOq5E2jXI43LGWzC8pJy5bhXVN
ZscS6+P04DnyPK+VwuZLcUT0i8ktaA0s01Mj3PrGXRn/X+jGeffEEey4ej7AD8kf
fXsQZ3mdqJv9p64d0eNkb7cjfJfssGBZlCwKaz11B2MhQNQTPHD5xKvXqU9yIzbF
jKyfVFYxN73hmZEjMZnw9C6bV1tiQhfQN6mozTDbhzVdtHSqdUtLKSo1XmRJnN1E
d2LGRez0P4ipyBgvk+QDyv02ypEgjBMBCDg9kSaITAu6+VHWMg9wYutbvWWylgK7
qU53oMJspjlZIW4gu6peaz/7lvMbXT3GJnID/YAow7LIMY6a3ygc3V2UEJbi6Zu0
X88GrnKT8s7PNuQkoKuebgUzUnsG50XcSzUgdDjamZmZn2qkYBfT227nGIVNC6Kr
zwqe2BmlhxBw5immw/j+QJ6kjSpSFxw5UEQiRQVurhvgIRxTKZ50Ec6iVwlgQos3
kIvKkGHHA1HTHLjsk4CMxJO3prbd+Zi4uKWuJB9p3zlDflf0ZWtCSpq/CTLughwe
UeKXUWFPxR7tStIoxQNxAtDFieq2YJwWrH8uSEfdfygxMYzoaxWPfO/cmvS5Pr89
2pyw65YCHaEwfqwX7p0Bm3aATKI0VGAAoaBeB2Y8jYcLYnEhU0SorSu59exIoYpa
bgIc1NEPFEu2ss+eoCPjJmO3mV2ouPZjH8T24naGn7lYrNfvXVHF8W0FQHEmuV7S
Ieym5zb7ltC6zYjW59HEAbSF4YGAmauDfBrAqenZB0yMLrMTjk2ghaDExj8LwVtb
xYl8G3X579F2qNtofbPglOW8YhmP1PZ+k2X35vVOPeOmaXLQFW63p5MrR9LBe6+R
sayUXzMVTz3e4Nura4j8CRMMpy4cpph45Tw3QSZW8XN9SFi6KyYTgF8nBmAd9iAn
oUnys8jAe9iyKu/liHF2ou16lMMUTgmoorSgTc/9ZWM1drYQKjV9/8v8BZTPaiq5
PEsLs35T7sRjcWZy7phRU+HEcpypZmDQHRNHjlv6DK86fcl60ST2N+872m2/MWw2
JoeuZkVh8PCBlEo1ugerpLo5Sb6vIZJPJ0HkUrqGTfxzXnoJyyISZId9IrYlf67X
UEpnkRW4b3NMxg2ozWQPJtgS5qwIFNvfR+vMBAyGBwYUTGHAe701Z3qeUeChHLQC
RkdDmubqYZjwpMZ6G0VBNB5KwFdeSeypgvqE41r8wpjKgLb3OwaP0Am/6H9648fx
YOjHiKvgbyJANtFy6VjRBUy5OuqVG4kBmgrXuawLW8rWe4qf/SbDlnX1spsjS4SR
jjGAVAQVjjKqjAn+09TOWTTnbTGTrfS9J2rtWWrSRd/ZhWP81mzUryJKxoD4XRwc
oqPqCTO25lhxYbMBjugUsVZb7NnM56gT4UxJiA9l+v4X2DsYG1eNs9nvvkJsVQ9n
YOBc9itXGhuKjiJFpBzCBiQ9YqEy0d1Ke8PkbMOLzvBsDIv5gS8L+mVk8MX75q41
vHF2NaLoGBUJv49KlS+eaGk160Mj242vsfw0jMP5Zo5eLdcuDeehhB8Qsg9eQ4YO
+VCpqVvzMvOsqVPPzn7vSH4TtaESxKvygPQhvUWt3rStO1e389/E+IhfJt5aRjt+
bgUkVsm4td/u99kFZ5rHpxH8nTv9tGzOdfZgdQPgGsTzrtiSn/kWzg1e23XXyT9L
HuO5OxvundXWhi2lW1H7MsZD+OD4MpiFHl76gLNTS8VLZ2jPZdudWXDbTdYzzqx1
iIGax6vOkHFkhyErCv30br3YVhHTEK/x4qR2lVgUXC5r/6faGUUuqwZpryrLHI9n
wTo0gIrOSDgZSMwQp6/uekHQ8zBu0t7Exhc3HifgOUcGaKVAm+Ksf0j7WNn+egAR
ePKEvFNge0w0EmO/clMO5PcOxy5sslxTzC+CtIUrnz9KDpHk1jA1xS1aA0AxhtDD
HNeD3Igv4nNGbMQ8B491SaIE3E1pPz+IgretGnP5yx9D2lv1CydQcEsD/o2d7KjI
dvKMOhRc8qzh3wPPd5o40UL+D7/EWVDYnX96D/P7zqjKD+2RN9UxPICCeqLIv3A9
NFaL1oYGgA1fnmGAsdAmo3dLQySzOJzI2F37navtdnFGcfL0+gtl8kXOgub0kaYn
dJwOEHa/3X+A4ygH2VQidRNpC0CQIOQz6F1181fBVxsDhYycxD1mERSogXg5Qqka
ynyJc21oE7jKo+8aAzSHVzvhZBHl5/EfyZRJkHwNojbPkila3PGXjM44461zr1IQ
kzHyVMjv8r+d4auRZ8yCZIowLL/E8tM1XgsXH2RfZDt99XLMdST3bvvTZGyIX1dG
HjsobbW6bxyRGlJbODREwHcLDp7HM7fMQT5rfJ+St9uYuLf+m4XCsC1X9dxbP89t
LKTqb3lP2NU6KDcE20r2UHuFOcIO80NfiLcqkg6SC3w=
`protect END_PROTECTED
