`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BenLbRxfayYgdGM2PrV9uyh0SKqcgb8dFnS4mP1e0r9MW+VB1SJ7xBRF0+vspK0s
3XoVkHqrrtA8WbEs1Xu/t8P+N3CrR+//ImwjUAUzZXzzcX3b5mAltz42AIg5BWyn
Jh8ARV3NqW6Fu1EtCtDD9aZ7L7+jCvWBRaHrQaf3TDEa2tDqrbkVkoL7CRQBcrKl
6sWgmfCoMZ0RTj9DniZTxCr8P0K5CodCWcR0ddMjnH+oVvpHLdalvz6BD0tQrZeL
`protect END_PROTECTED
