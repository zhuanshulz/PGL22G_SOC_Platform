`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6qVs+f0iGbSjJ0+byMUqnRZOLRlNZERhNVFv6VXKPEJBS1ZolW4e9UnNZbK5eqhX
Mvxv2I2xf4iCHsGLe9INjrnw4B7Wb0qi8ktgiGwutXKgs+nw30BfXzb/U8nWRKud
aaTS19vYK6ERKjuBVuUKKGTYZSMliD+TT9bkZa5d72uJBkYLfIXeqIL+TQPpSK2/
voxgxocARNRhjAAl3w7SHtci6HPV+YL6eTtfZjQJ2FEEPI4s71646OSt/hpYhibg
5Tj+WafwQm/PomyWYi3Ow3lz1Q6AHKlgTvEY6rrje4/fOyNPaBWILgPYhGbrbo0i
FDuGBi0U6JnTiiIVadL9gBzglNu5ynZaJzuaE1V0YkSNpGz2k8fTWUrmMy1haa9/
k43D+DS+0fj2TN+/sT5APdM12OSQlG0h0egrSnmUvqZEE6ADFvhFfPq4PCZao25L
LkPAVnMjw08N0Tc2/NcF5kWzGA0h9WJsym1uW5Z+jU1YKnPmrKidkq1583tYm6H1
wzVeXh6bmFt3eRlBHMr1iqqGO29naFdL2B0zzqg6Q0Whzx8CJFZTdouDn1uoZ15t
QZpyRgVr2DifHGIVzqmwIGaEPdDfWjIwqwk2PtZFIAKOxvI767YgsKS2K3S2bEe8
9LSjbJlw0fHtGc4p4jn81l0hOg146cOxAOa5y6CunrS6a2HlxT7ye81U/omm7l4g
xtYPFNtb9anNzYinyng9tYk+nkRT1GU4PJJ5twa4O/xf9xY7jGRKopSSBimf5ksc
Cu2kssGjuDWNqzeEJHEUnw7MXX2sQbcdNIvcT1QTt8om2c3qnjDcnrepiLwnvV5X
XX+07ENjzDkegBj/DjwNh0XUXKsqIcrSdJKLMrse52SorSCDjx+Xf+w9UKNdh+NX
yWKaeYZ5EdeBcOb3BLwfbcL/NGUgdpyAB1YAkVd6iKLUzDbyzFM6Yj/9zxgwUdfP
p+cs0j6CKr9RxArDneXNBqrOjTTkYFlVDlmNoml408xoqLlPQsCfoAIRDTKgaR5C
ic2LF60d4IrNeal6eCqoXxarCki7SEb95JAz5UgUuyvUuDldFko9BoNjJa46JFJB
PqzzfxMbdhJv5KI32lz9ye6O04v1YESYfH8Ji05EF3ImJFFtpZxI+Sen9tWfWzeY
3VGorcUQNa8LZombKVABo8PboNc57sPuGAt+fG4t6zcxvdfGp1nl5VgtqYMa9y34
7AFX5W08CcdeqeqeXknkK5AjOLTHB6vr4fsfve/SlxuTEeLO6ey/I+I2rOelgo2f
tQsMKHNRugg+EaLmrHB6rRmxylRVrqp7ai5PrYoMQLuA1SVW99PZmKJdrEBb1u49
SH3x+ztqslkxRdZijUd7aK98oruHEzl8qZNvwUHHg5s=
`protect END_PROTECTED
