`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frjKCijoZOMPdKugRkqSsjUvgkm2a93qMR8RpFYNn1TYmbnnlEm+R694pOP/qyLI
EYAErc/EtF4ibKoj1ReHy//ajezQfp+0bXutJn3fhG5XTOk5v7KCocCdW2DBtpAw
qq98MLF5LwjUO702oyyUP9vV72nJkW/g6rRg4xqpZ559muK6FYKek4zjU36U0hJL
FZrjBMnHTWj757biV0NuLXMghffx1L2rEhD64VwvzfdXoo1cqWtMWnA5++lcCSBu
CVjAr3FV2zPtknZbBc3kYHJ8FF26qb6aiJjFXxV+yEWt6cZRnImXFR03eEdPtL6p
JUGkpO0Pko/PwHJiYtQkUJI27x4fcB+8tLtrmUH5ZB3+UkQfcuQGZdPPQLcHx32J
GNHD9D8UETPjWSnq6/6XMOqdNpJcdS+W6wXMuX5EKEwXHTZ+KGliNUnSIkQ9ISuR
KYuxJtCZuiEHkW2gDao35BBuph+NzSddr5x8W9UuDtBUovNaMTV7FORlHiMVIYZI
YEvDiFc4vmRbXilNqeRMkAlXNHxuSyybWQFyP+0G5F2Wi4ak5sWDzT4EZD3FesaU
WgbsPyZH/J4p1oC58ZWnDKxYVQ4+mqMGTaWg5Ksb+wlkmF2bH9gF+qeSg+weNHyp
mWoDgh1iX+chKItb0z6RgzydFp0AXiAG6LQw5z4O+3xJEgufaG0TpafCdA1qpK9A
RkFCmXN9lQeZos1VjkFfsik7WTx/m2qIhhsHCUtwCS+U9fmKg82ETRYW3wujQ2Ov
rM5Qy18VGqvtkjJOhwTVNku0JzzWFV5zWsICqWQmcJYd2B0CBmEiayDdSe2ZTR10
`protect END_PROTECTED
