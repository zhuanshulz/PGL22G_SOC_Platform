`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V6kRr41JK+/xh0vT7tO39b5TmcTtQZcv9f3UyZRp1h7zNZsPrz0ubvIwibn/f4ry
JVr8eLtFKqEJx5McQ7VwqpazpbMQuCJlB/PvCI2fBYqgsV6vqCkyMp6ga9JHt71V
a1BIoPtcfT6f+69f4wR4SfDdvdPaT8fSyrRq4mBLNgt9kpCn8sKBGUsH0qprTDd9
nZlneFokWW1c+8pZzORg0MU3EODO0tzHagCJurIHB2ETEKXd0lw6Lf1fcBQhA8k3
6ePM3DSYri3h6kZk+wygbrRCCl8vxI/wz7JGX0RfUiOple5kV3yzv8QBBzWOXSMs
cxY0aQO7lul2Frajjmn6C9H+rPMc/Q6yS2KQoqXUTPdxiY4omXuEi5nZWxj3XcV8
6/isN3jM8/hyDmwVZxKlUdSdEQWeUn7Nzp2DzldRn9s1SqpitSdVVbY+oU3OZ9pi
xOhGlGf+g2BzhKTxl1ZimwqzlmRcWaqycKD33+UdVk+IHDU60wIq7OlkIo94fQKw
EwtWaFY4IWGsUGU/ww96PvX0MXgyY6SNoPhJZChxRTvruna4w8QazrqB0bg5JrcN
`protect END_PROTECTED
