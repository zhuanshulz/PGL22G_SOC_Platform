`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4KHU2aWFgM71+kPbghHCBno/SqUbSRlGSDdN1KhQfcnALdo6k5ioeCHfIjWC7ucn
6gumcbx5dZPB1/Mjzh/GJZdgDs06iaUiLqvtraf45Jrx+8iLEuWNmARt7078tdgE
0L9Dz2klRndJTSVCCFfgiIDD2OcpDKODz3uVuwouUxBQKGEvl/LXEuLDPC0/b++v
Z/GospRGbe9dQKJpnfrM1WaKmq9Q3hudwt5G7LPoc8KCZXoYPU8wW3SZ+ntpWfw+
reZgj6Q2JWceNKPSzsWGRvEfnMmyiVAv+Tv+kuZJvacF0UU5qqs2NxR6JKw58rtT
N+wXzFcqQGERQp4uMm8DhWviIJjzAno4BK8pPZgg+MHmT6farcRqHCr0p4Dcune4
1oZFGZyDxjWJgDQzLLu35Yt7PDCGrKCx6U+jImAXddcviRuZcJqsnGuZ4P/p4zlX
6jish3rZlL7bsOnPoShBDt2i9dGiXYvA3ipOeL7rjwosU1By/wXlrfkHJg4rJR9t
paFZz1BZFGMLn7QfslrM8A==
`protect END_PROTECTED
