`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JegE6mEbS1Fuw1hPfaZRFcU1tIPMJa0PY3RNnDAHXbLzncRXxFScEdwxq1DbUpcB
d8jJdH+2zADVDZ5Xwc/iAjfWWE5/BEZjA/Pvt2glFynV7mvfFAz7m4FORZ8uxWXH
zv3gkj8MmHHRNqebINCrK9IqEbBd530rfW6DLQviN49r1zqLopWJKeOy+s1Eb8i4
+693vw+J/V4nv7aEhAak/VfFJttI8zwTQhWfuEHFmzNxEO7adAfTyihP6VHzFrqv
4zfF7PHdIrff5L6tMj7e5ZdsY6+LAL1V09OzMknJY9/RjpZrYiqPfZajYW3Adkb5
eLl2fGkZjJ2zQi5++QMwFYXQCx1GPKwDraHOWClDZM6AnN8SbZuVKtok4BzCij2p
0+zHwNekaKbSeobhsMy9W/siR/hr57qQ2TpTT2ks9uzbX2TilC8/p4cYvpjT8s7g
zQa1mngDLIzRJqomGPn8KJJJn3ejAmWbW33tiTUgGtHVDiOTQOznMGPADObWKhXT
r/0ksWxnDg7ZRbg38w6qmpDSnAL5i28nQPWIWyItQjO4zpimvkvDFNLlAJKz/UQH
gzLkCKen8/TD5Z9KMlPf7m5S4ZLg4rCjNEYN7Gnk3A6yIHb3iop5vXGIqZndoOUy
gjrwndluCB8qZ8cqGxZjIsn4FzblURhCzcS7UM2hdanIwH3+/nBqVEABJvFMHuD0
jGyZp+9bm/WoTMe5pN5iwz5BcOa0JEmEgN2XVTHEZ2YF/hllsJFFhOFvX0iT+d68
tGhmu9RPCXaBf8xwiDXMfJtR/SOwVG4eGiebT1TYuHLF5mhIVpjlZusbZXXY9CNc
9TR0Sem0mrxsIRgwpwijlN3EooL22euCJhXCqjckqARcNBR4vni0nbHmih7hAA3a
e2sjnGBymL2tBP1ZFNFGPdpSLFd3AhNryFf5vT9xK3n+5DX1fvcm648foIsa6BT4
qnS18XKSsJzMM+2jriPCApXA1aCOY1hRgPrOl8JAB9bwsB8I97WmnavlhCzNUuWU
o3jeslggfyAGdOWiwUoEaOS+MghPp2B+7ttgrcO9qUUNPnhyNQqAO5rof/Ix9QyT
59wblY9k2Z1faK3egALl0mGaxWKivHqBu+QjZ/ZQf3S5JIbyhu8rVRJ+PRG/VCgB
gx1dZTDCsK4WwFX0w83yHa3KG1TdEVNlJ2o2hkP3cwRevFeK8wB2keNbyntnAiHs
ZLvY7OzGnlTbwR+w19Hj0Zhxzz+x6xt/rqButhUi+Aao7L8DFKvGCYkJHPilY6eM
dNbF/3joj09RuUT1FwJKwXJKsrvWAFB6BWoIzT9NOTJ/1hXithGPslc+3d0wnRM+
pJ8JYVw90OHlsEAvf9P1D5wPw9WxBZ/ySb+n1TV3Ro5SlmCokAV/1TH/iOPmYe3n
6ueNIiMrNvyhdRFhEF7XKBkqOCgIB27CGqF2ekd5+oxurNBMVeKp3JOYn26MhGb/
TdcUiTkDMetAYPnvWuKC82LTQ9PKW5s92D4YjhzxvJ1lbc0pFfY+XyVryeWoK9At
ODLKaSXd4It6Ge7uPyTpR7ammnZG/Z2p1b/xlNaVKTy0r211Ej4/6kXICe8uhhDH
9Tmu0Tvh+ZQXIKvQECTNV5Kfi1v5DD5IEAOYyXX+2scTkXwX9sRB/I+ijYhKjcNw
VTx0p0Ujj95JCX7CaBrNGtulMj9h4r8NuFLnqjoHJ55E7+p1y0KOL7Gt8KFM0Hej
0TfkSj+vx+6PxY/oFW8eJHXfeEzROcMFoFC2lwZK9YelaxTXXZa+DaN7fTmQIdp4
qC9xDJsL07RBO4SVruS1c5PhXjVNDsrdsmPEVqkvQV3GkliTX5Woe9rO7wZokpIJ
taDAC0eq/ExFDPVMGFoB2SgPsiC1WOvQujqFmHjR/ClSesZKas5Bs8GtFzOiBO9E
oKvUi7O+7YwO0l9ZJUtV2cPBzfXaRzQAjBW92UukH2TnmYk22mcFohZp2xYV8dLd
Ca8F14wBfS4DcetNut7Mmme1VHbCzlK/s6GO5XRCoIRllj636MeG0ZYUuJJF3OiG
LLXUkNPMzq1+g2bmsSByfCAgKs1pdCNbo9Bq6IS3pOMYU21Q1+2YxSOnv8ViYEGs
zr4T4FNn2LmPz2g3mWMzDYLCRvTad7rYd1ThmaVh63EcoMcXa2ni9Pfv9IWPuRdd
3N2kJQk3KZ9UdaNYPBoWwLMLaU5KbXJPIuabKq0+GXWeE9BEYC8RVcafFv6D4aCA
twPrfWh1LMd5IjgnDqtvSmZl0pW3HAz6WsnwXAL8cIfbkjwCMWGOSwzfCPqWBD9x
2lYv+8c62cgrketUvEpvTnkBwTC7DbbYPdhZi3MsSUS6U+qnBi+//zy+62t2SH/O
`protect END_PROTECTED
