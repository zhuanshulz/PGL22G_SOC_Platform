`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OF4eLrubzfJrXcJS3gqKf0dGjqDZveMTMow5pzfG/5J53D629PH7QIzMtGxaV7Gz
V1PageaiL6x3uXx1LHl+tU/22ILaOLyZ4c8t2+AQp1c897T/BCe0mvux46MGylDL
CdXdK/bjGm0BwyLVoxHQvvJuJTdGYoxYohtAmKFAdbLsa5FnmOufZsLeCUd54iuS
WyP4tgcsMVg0wnQ9AyDCZtcIEiUiIvmb2/WqaubxnRUaMM1JRdUL4ibB0+vvFELW
S0G5Dwg9IPCRKVAD/yF4lpEGA0RaoySdgfuZoR28iajLM/fPVCHc6i9o462HD9Qk
1PmvNJMH8lZ883tiFdrnWk8FVah5DxVN0UxC6Geif+93exSDHRJzhnNzhCEJCsD5
/EZyX5DU2hCMvKrCaY0qSUNZboKDGfvSrOqP7ZjdDeSlkGXJP44/zAdq0ov26JZc
u4hgH+rOmAcNXu8NbFKrEHL6jGAnZeCWvoxUG3x7LjaTO8ob5NLz1wu2q3oOMTn+
43Rnrc3nu71PUF1aCxlSe47jOjnrHYyusp+anoLNq3ubkcAgTom/8UD6+tiOTf5F
uSvTX/C+yO6NvJsJbBTnZ3fk6XGULqGfdCuidRGrjUc37t8D1XollJ2Pmj8CZKhU
lzgN9WLbhsllTBhtbjEbsTvq1NKy6x5Bqgr4060c5FEls0ZLfnsI9hvWVRVEwNcT
p3Zov7sO31Ihu50c+e6kjFG2QigLMe7q0J0WxY2VZg8VlgaJWjA9/sNlHdMFvHmF
PZo+miOZSipp+02ETs2Ixcuo4Ug9tyDm0y65oXOeRrdMSfpRHq3zXzPtzg7drExG
2hCOBytyAH3M0/PD44tK/wB+V5ThEQeXDuABmzCqkpud2hO/XV08+qzAgkd+XEHt
EnRMwY8vStOGLyE7JGtLte1xKDUFMWMS16tGYZunmLINYI7SGR1h4FWlHhJdkHe2
cEDNThwVXCBdg+ufsJ+Pslg5uCiCE3TRydnB5ACglx26wu5de1/yBI9Y7fny0DJP
3yn5xDpeHHs3Ftfc0MoNvZpwWrDeEA2N3JeYeunJRUO1iv3NCdeVTEjGwlaHt35O
KoEI3cMT1cFNX8rMJ5bWRiNumZANBW74UC5gqkrVE1u9lYIFDBCko6pHxuIErrtX
vPF5SpkjXq8DvJl1TWp4c3SDBrNa5DWjHq2ekoNlbhSehvIRwiMk8HUwUUYV26IH
qKKJXCKn/cZyUvtXOPHzdUkgOq1wlUzLb5+FU76DcEyAVvxTnaqgoWWXF6Ju6qei
Se7ywEFQUH8+tzljhek54DVjegs006AFSL5nZbK0HLkv/Z1mTHAUJlNYH9Y9NFJh
ixLu3oJ2sBLleyKP+LORLIA29ka31HaVhviGvDwXz3xeLuCtYakhmhYnsUFzKFdY
Y4/gvZaehMmEMECc2x8WjkwHa9QbGC75Q7ZfatNhYvf5XvC8THZMSP0xmfXIQ8+I
/XoXRHGN8hj3qZmUpz9hAJHNVN651PPx89G/Cmoqwz9SG9I8YjAO3CvVQ0gKZdBN
iYxYJkXzpcR/DSeyzEhl8TDbUYXK798Ro1gnMtDVzOzaGxbzFwbMlwV7GgAWRBOJ
O6bNEUGSLEinchRJV6gY4V5JP1Y3HO691jXs1n24DjJeOo5AIllsCVCgtkaZMW7O
pNOXtGg3gYQYGu1Se4ztrDq+oy9Ffb/JDAJHM/tk9T4OAR5cMHNodlmgzb82guWy
4BYfU05lcxscOltUAWD0EWG5g4m6VNLds6u2t9Uzr4vVeLsKkK2CKBEITd5LdoPc
ySpAQGyPPsmkKiE48/NwgKPKM4uvqoHHL9KquOHzJWd9jopAE2oQiiNut/JMgAUd
Wm37OwavLK6Tqy2y8qumO6NC4UGGuLt14/DZlJ3XOrK1rzPTvo5zTkPJ+TDr9III
TVq6wJxPVsgZdb8BE3k8T5KcLXP7KzBjoFczD0Ymu7eVCp8H/1v3lQHmutvZcKig
NEeBAVVjmHKC+aG4rf1ZQkG+oGhhfRHap9dycZAh4cAg3PzTtyaKpGvLSNriZDtV
6I+T6abZ67IDu1nV62MTaw==
`protect END_PROTECTED
