`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ct7MPR1hajEOnL33gGvnlPQtJfPOW36Igjkdwz2qtHE/y5dwQCGYvarQYuXz8zJq
YfaHBezh+7Wi/xHvUCqHwEd6TtwVwRwwDL7gftLcnFRrTaRN2jKTT/4ebbDGymR3
lu2j6vQGWWpY96nEXqA4Lcerqr3DkwPv0YRGffzf85kTJH/f1dfMqv4Ytkpjf+2v
YHj2kOJ1bkKcDio09rxXhHYbyLHZ88QKA2OO/jN5xBgllOFxY/VE7+Gjw2/mRoOx
QCDwG3AYXxTYQWNp2s8o33bIpXWj9BEFeeRTBZqJ9vX19FaO4s89H2I+AfiQQenV
lv7IZZ5qsZXGxQRtIXPgqRdlg6WcxvWJHZ7dnnV3cSqZTHS7c7TToPj6KcqCpgaH
Gmk3bTXy1V/3EcZDGrDI2A==
`protect END_PROTECTED
