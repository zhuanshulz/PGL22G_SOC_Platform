`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XLQ4/SkTPJsVaUtK8uEF03OUcahXLYnBQ/5JfBHPAuzKdkgcDzGRR7rZR0d/lfwl
MP/5ZBYBGR531NL3IQLNHhEwhUDpRcnlbJn0XBET5OpM3lsjmIi14/GHjNaA43ow
y1c1ODCMVzMYLJSMBU97MMArB0DLVTk3q7Tmhj/bxpaG3kVuc3Rblz/8vWhbEQko
czKP2C/DM5S3J9somsh9OVp+Ce/jFZ7GX3hSOtmLe8pzW192N9CbW4ygabnfPBAT
qKaOqRy1v2YDLPn07XCsc0G4zO4yfzvYYXSyev9MqCZSUQIQwYLjX8Y6dALJiDpK
kxifMeco3dCYb69iL/g9UV489p1CCvkr/NIWkT834QSujnovjKHP8yWK/HCuQLHC
50BrjlJ/WhoSnL5RzN0kUTd8jExKn5jcWuwPSnBdQVGD76U/xKvdL5lJra/qlBUd
p0kdUP48JjOyYuXFLWymNYhShCxzYXubkqlJpcQr04azGcwJT2vK+4ONr0n3haDI
qfnQQnTgcBvUwkW86B6iIhuVh6V4LBArjVIOhdj6o4sBP9wUMhPdbvwxIK39O7A3
s/XXGoQc1IKYv3VfQ5xs41px0nJISac6u0sRxiRqw4jvEWAhrXQQ+2LA076pDoKc
yPmqL5uL8EtmicRpfXa952O8/2ZgQYfSo+mSjmhHfRuPmg2jZzDrbCoWuXXxhh5f
BXhYnRDIpEYnpdC5j+IkRxgqy++8sHUVgpcrsJhRuH5iIsTU95HRb5LpYeZi9Fr7
kaA2LA6GLZUd/ODxnBB/rKTxfQOX0Exi28e4FVUmsGcMah9LujAChHYy5xkTMe3H
blxfn0nHSigD6HyPfw1D2L4aBd5vKBVTYHswWoPYXV2ahVH1GTB8DH8DvGdHWw70
gC9SWqW0BLLeBJfwoylulTDUEnZoPUhuNG2Mw8GR8x80N3tcvKvImv8+D+H3WO5e
RBfHnkDcmnnPRXRYlhbnL+7ONRfkDNyADdio3/1yfcjn0P2WdHvDHu7DmRI8Dwd0
pId44qIRAlR5wrHACN8oKgFfmI1ovuG+NuXYATmisamqKa/unS7uBC5zuAs3yCtL
B7YihJxhMKvYLFlLdyVEQ/76ARKzrgRTyPtqy4kIqV6ns0dfaOBIEUpvyeFIG1G5
azYVgSM8s3KBqE+QNkUfxooDIf6ff+rMrtv9gNVEhnS7l10TIb88WlveIef+1aue
+rNDRl+qG0QoY5n0GNhrWNtSJzPelSToWILVH1BM6LFZcch+0kyWFdoDON2VlwB9
`protect END_PROTECTED
