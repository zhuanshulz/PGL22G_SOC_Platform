`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/rZjVt23v/5wTVShibYugzJyBT9aUspLlLxjOuA2/Km/2undMkpskA5HdoiUQJt3
RGGavZEwv4kwJowvV2H+d7lojIxLfeBqf3clQAXPiu6eZ26pramRzfVl7wN6uCOG
XPcwWOl+OBe95GYsJN88QAIq8DdGpLemC3y9KAk28nWCGRVH5kWpA7zo02AqMSiZ
MQqiLs0kSCs2wLjVmw+Gq5xAv0HFMX46GnkL2dxTKb/thvbszLcwMGx/EylsyOV5
nIK8DngI9nvKLHqUqcr6/eHoE8YAhdd/VJ1gOvo9whNgxGN5/N6/JVCrf1dXmF2S
YXshNOCl/u7BDpfb362b57WBgmSVx3nJ24BR/4WUDQGF5iEUdhIeW7F2QJ04zm+u
oU8+LJ+Zu6lOk9UeGu5PcTg8Slsa/p1//9JpUwwuZJVw5SLN5ZZ/hGthYkbSKwZU
iWumgqmW9Q97qxzpLbdorIsS+z/B8P/8RbjupnAm97bmDAjROro6TtVo9M7/IQSu
ad12s4/Xc1DCwDgrR/N66IjCf39Iu4cwSxd45dpKAVgT2rHSM06sBnh73oV/J7ED
qQeEQMiz1x6txB3unGVRVVtgRwhoIIx+w3PAxRlkEJZX8B1PmJr5+y5tjx14OYlg
2RizXOJluqiihM8Vw4eAw6MQI6nFTKTbQmbHKKwG7S4=
`protect END_PROTECTED
