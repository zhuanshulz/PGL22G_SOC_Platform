`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHYj8joYvqxMrCK2eDw4fH6NQzt58nP8cfHMqM3fV+OELPFzBLZFfyt816MVBzC3
T64dVKLgrQJlp9EinJTiZLKXJxA69TMNYMdywY0vKAojSbRHlkIXCRnCbcYUE1WG
fPhHJbrNzIm+1rpHUNb7fWiAZbETON9vO/poRR4/HTGE590tK4//jMjAUa6MtV/Z
tzBbxo2RuXRfYR/bBdv1eIRuf4bNYKqmy0SMVCigAaYhoqpoTTOtxBBbe3NRfBeA
1B9NvlFqQlWCTa3gNRusj+/byDiLCVPK++J9xaNK0Nw2oyfz/6BvkfC2YLM4IMqF
iLDdbou2wCfHMbI1UOYFd2HCH9Uw1QJ33fnaUaL21+ENKMgx3FfKIkxRriZ0fPDQ
hI9GodY7gUrOtCXQXHKDHvFWaxrRZ7f9Y3QyMV4v1pESGst9is5jm9ACpQW0qv5B
Rlp4c/6uhJ/KRx9OlN3Ej9XE0ypz24k3dScgua9IPZ56GMXEdvelR02/zkN+Om5U
/uyV6oJh2KdkaOM/lkkzJce92wn1DMmDTLHzFklZP86x3ETvD4SM+WN8KWqJW2vZ
lh0FCO0aEaOwgHw0b2pWf0hoLVrsDW4rQIS3a5XKLSHYDttYYklAvVFIrQszdF4d
kWL4nyP0EJvIOXGPIpspYe0KF7Vnsz8GxXjWTqElPVuOmbZGZ/LCHI02H+pmvAgl
59urkDgWl9x3WpZE2SgRq39WtYV3IMXAI8oUapn7e70Ep4Pu41qmFyla5TIdVB0z
RUxEQ7g8zyFWowr6N1dEY7vzhQq9WdiSyw6CdgQUF57gKvjEi8/We4TOjIB6B0Y5
J77oaIpAs+o/QIoyWBaRfibSNvXxAksBsnhBRb/6DgjstVD7VcKbfZDWRO1Ugo1s
8e53/k7xKK6wNkttfmcw3c5F+OpVp2ai2f3SCd9QfTrbxvC3KM68+gnqNF6qQuw0
znRJYi/mU1Zy5SIm/36VdcoIgFRSMNgXk2jdBB89NdlBEXC+WCD6TlkeYwUZKy+k
0h01flkvkMGLGwG6Yh+tYGeFDPAKGrbPK9CT712S5KOUmCDZjdReDAS6cICkis3r
yWLs/SctyctJj1uADLyx1lXFoNGv4plwHP+XaWU6o72bBAoQMkZrwmMXVIOCSZ84
aX89+OfwwE2FS8L/2qRcPr8pTPgSWlVa7/NIsNqPkbCMGeutsMoH3BBNc4DIrh3d
mc+kv3wJWfgUud++ab4UT9ImamYzJ9oJOsh6/Dypx33zl1rNvGX5pziC73+1ZcNI
PfphbsX8Wu+mCd4VN1uu0bwOCxH/EDREfneUKF/mMXqMc1TnTaFuCEs43bmnodal
bnXSv/uOnmXznEWM2pmuk1T2V5pckLVKAbf0z3lLsNobUkEFDwRFCyyeVdYwkfsF
Q8YooAwlL1kJJFVywQYaIPJRmSrg1FMSl96Jh/86QaLLkCD06PwGEnLus+RnslBk
ES1MnOq+N3GdQBo9/VilkJa1XfHvB/QzDs4s2eTBzI4H2r+YatJXjEc0jAGs3Ny8
4zFsoGxRoudM9QX+cUSRTAxX7HmHYShxfNfwNaoxNN+0ka0gPVQFD5q4AUU4LQe0
/Ixyr+Q6TBa7tVE0P+w7AcUX6LI1XwtCk5ROAm/fvq3DitEXs6jzcLJenL2Q+jSs
hBuJmv1wf8q5DlMPfIqNGHfGcTLvlAU44oDRY7FYVlbq7q6sx7AqHytxwrYYRWl3
fh29+8MOKUKXxVKIdRaRx5awEQz9WqPEtwJM9cryrod6Hf0H9/VHbUBYlnNw1H/B
q18xdsGvwPuORTUU92Fljd0Ahd4bBhCxxXc49PDWjP3n+EUqw+mOEmDszC5IvgQY
01p9XKzMN93BgvwZBzUyDjlfHP+RALLY8ZHLpwYsIrcv3bNQtzP7tEiY92x/FY2n
1X8CdXmJbuN/zfgBLb7Y9RWYT6jV2PNjcH4zMlqv1vTkCWsZzZsH4AkArbjCQ/JK
mWmOya87gVF6XwGjdyXRl2h1hZcj2DfW54b+k4GoIfwlm2IQOyZrD6BDh9150Ytr
`protect END_PROTECTED
