`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7BWBOTZap2p0y83r7oPSTiKatKGz8N3p6gMFI9Rqbr27L+KecDgvvPg9mVrCCS7
/xB9jwL7eoOVwpJk5/DDZeZ28qIBom8FgSIZUa4y4QIszoa1Red0oFmca1mMnG5u
BSXixVqU5ruHhEVmo6OEeF0cU0HGpVrXVt8yMpeUB70G+l/T2iojRBjHZ3dIcvdG
YibXQ0AWBDFZQCBg98ChF1QMwyiydR+wFuQ4i1/hWCnMwG59DzYTmdTIQMYTaEBg
uIAW5ADcmPMlu/GaeZbXu5wzn0X2EYJukaK7XbZtYRqKz/x5fvuCG0Yy4zII3/LB
+3uV/ehQfzsJDdHnwl1lBJUEqC6F3nURWsV7w3tBAdBztPmR7DFbLdm/IoU+Xx3f
9kcSEMRPMu83gCBaaXJ2hJSU16IeW2aAy6gqEFrwG6Q=
`protect END_PROTECTED
