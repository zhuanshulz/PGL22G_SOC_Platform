`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQn/xjDG2qZ4jNC8U7Us4jsysoSQWXv9ASTv23dCmV9Nwgc9BsVA6ZhT2dDgWmZK
BVGyKdrtTcze2RVybGkm4ujUL4LxnRWqijHsHa31d2ux0GzVEDPCv68YN3VMOCVC
jJlWbvKZ8lR8/ajVD7B4zm1ynfVS1K+FyjuAtsi9sAXo32tQfwu02YsFU2+xxwOM
0mfgUC5/F45vggxYOVVVHISnD325ySOa9VyatFk2PXtp/6ptoAsCYEm8UG2Gby1d
0uHgOAm1v0ghRTkVOszCZa0XKrC6GxmNuWEOeYXelyS2fKl/MzXHBKu63vj+/Jyx
n2YNMPv1D+6rwcuxhBG+FnP1kRMuW39Lu6yLNSGDeKtSmZIir+9jF+1xBhuusrTj
+2MljanC29EwXlgd+c1tsY2QY1aX+jTzesCKXpdQ5B98iGvP1cTtopvra5K9ShsV
C1E1+cOLyVwiLFPg6vVoN0bnIstOrnqSkqMNXVqboOMfznTKZENz8Ci+wxH4wyk4
rChXbEAYotvrMADBcaetUr0pRbWcGahRPVKBub6QGby1T8ct7rLrWOACf3TmUsXS
v6rEQkwxW9pBzJ2y7VClgHp50EP+sai64NZMUDtirIRVHlY6wJpPWQK7Am0VElkT
LwLtp4vLHeOqnl7fVKwqXRuH0XOQ7jHOPJvweEy9qwP4JIANYqb8xTuNi6KxFfT0
HT/v2pqebvltCOQqfBZT1ybuvn/omT0+5fi5wV0HwIsPWWFKhxzzUQiV2soMYlDa
FiOhlV4ekYz+e87QP5u82r4o4Sux6DfZHRJYF4HKUZk=
`protect END_PROTECTED
