`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RyvUMFDJ2hFn+mCoO5FklokHe+LASkXPTePh+oirHooTyMbPFAik4rznKxxTslV
hQ51GYvugER/i+xp5MZ895UFgXvIr3MXmpmm4C5tGcy+pUYxeNaW2b4NxrMUwKlC
FxNfZ3SrU5EW6irSCNejyKKg+yLaPpW82U6ooC+nSysXLiSnQn4xz+v/V3LjwE2Z
xSAyj+mYPESIoZSZijQWOSDcr3ZvWkFiyN9VJUGrpxe5e7+AngBdsTP6Hv5qadqA
WmfSyfxcEGpjhE/evXAgfD9/Q1uxKuYlIMqR/2FQNA+YPJVOuHmvbZt4TakydbZn
IEkvO+UNcPwq5ocaSuD5GPD8p60kS0KX9fk02r2CG3UKlm+KiScKytc3fBcz5zC3
iVZ8rBMEpl1YSYsy9StPE6jsLPCu4H4R2lUC9PZGUJflE/SH+uFkDJJudnfEXAXt
BMmjzp4M4P+ZIWlaJClpv2OlQYzCSWu+7AFvKyhRgx0WslTyQ1Xr9Eva9n1yctCw
kaGRKy68aIwWX/A3rBep+e9k1cs0Mg2WstYNcTtNv139fo+mWrIiUhXWzr7rr7sY
jaCP/PYV/gOmt+dthCIEaVXUdnbSUaXHCuwYoaTmU/p+QMr2ZVIXxxGdPErAFF3d
ok2CmhJaDJ+GseqRFdVQ863Us2DjIeara8N/xmOslvXT7cNOeMiLNH3sJW6q+ISo
brRRxw4lJtteu3oEGn9A2OQQ0UGyzY0dVVUCzG7frdC28PZhJcUZpWldPj2Fvhja
UnWjbfqrKgr8RnV/cc/8mofjtUb1XgdLa97ybujeQh89xK5GjQfwGrXytsDTV4Ql
orSpPEKuS5Dxc8exerQM/EAK47hAz+TaXoPjVoGc8hLCQefZlOV0os0AdHD23vm5
QWZeHyU7Hdmygr3xF01VJTTottRzDoggltdxJjxFeLKQ3bhh8JJzD6XPEOkfpI4l
loq7kWp2Fhmg2WBKpGlJIQNASEKFTFEerYkr5nMBpJuDgd5zdRDQVe5GnOg1cdpa
JrojpiHprN0anH65LfwqKvqfdW/anWl/Bdz1epJYq7KGn/66fxOsrPXlC6302Stq
Po+AopVGqYMcYlelSatFF0I4qhhcPHj6SRoZt+G46TajH6zSs1YJOUUSpgvTHvWk
T9qvRvElZtjuYbMm1qChpLX4I/MRKLZZfW90N4NTPi6UMYwzCCEEdjGTNQi1njZX
TCms91TbMAUHX4jV+F8oACoqu1rxqQMcUnaSI0a1HI37cHNyGk+gzse1F0HFTCcS
IuD8pTW8sgUf0RA/SXj0KmQhuPDcH0SbI00YDasrgMpymoYHXlyNm012WqSGvXtp
`protect END_PROTECTED
