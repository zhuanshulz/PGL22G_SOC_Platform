`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xCwapWy3MtxijniM5lkdQAFJu0gDRxbO/nJtVTbM3i3kuyXggALk2wEEroCvXqu5
GLuaIeJxnd2v4x03bnylUSjxjay7JFg0+JzTBAaRnF5Q0HvEKS3dDwrSZr9DuvrG
lLK7S5bOIn7P/GBt+2J3uJ1aaWfafPa/Ys9XNyLBHgf5gHUEPBzh23mjlbKEnlHf
3ctQJjUSrhzazm/yBnv9egyUgegwIAbKBmfERIPueh5ogSd5/mCaAeIgMDF4LHPr
D1C/FJscUUTtRtTNxYkDUXWoWWl1n1j/y+u2Ek2Yn0ooIz3Yq6Fi7oaYmllf5II7
hcuyvvdwaf/YncyfSfUVzbrVjX6FEK/1ZCvl3Ccq24RA8HlwwRcikkeRFStLbuUw
dY5qLWy+rzp76521Y7iJov9ml2LyCMWFWq3iuKUlLl3hvn1d5XJv4fTOf0hNyzYh
crTcX0B9IqZJmanhYz5J4uVdh+R2B+OfAhiOXRakiRyS2N5TuXHXNnfVBN2K80d9
DHZ6nKAS/vFP0DwwhUCVk3DuAP0g7aSS6ToOrgJXF8/pAyE6kwaFccBfiO+AhVyF
0qibVHUmJ9NN9RDQwuF+Rcj20VuAvsvtXXZIwets0m9ysrjP+dgnnkXRx7LfizC2
nnpRJ/zf0bTaH1p1TNEyE3SvkQ37+t5zFx0wi1b5Pk1mQrXu8MzmXy4mYXM052Qk
Ln6vaOxwhPdw6qYAnSjbf0XMzhySa0jCPNK1JG788yhEjPtzLzU1bEh6veh17zON
QUFPL4T7CzMYRJ8zwVpMVj+7dgO1miQUGH4EDjvJV+OFiXqP+iiSyLzciVS9Jx4o
VObBnMHjn090zgE0UQyqibaJRFwYbXwh+1Ovi6fho4S6Ju88l5NBi92W42+RHnam
omR4YPkCVd9CbCnZbvJ0jH+2vCwejQveTvlZTNVN2j7rV6hVRwFr6QGcOSQnoWcc
zt8V05csDNDqicLGISf531l6VBZ74TECfS6qUjt+TT1kzxp8/Ac10l7Tnp+5fUbH
q9jvTKFMHISUBP/1M21lCiWX/i9Po0dD+SAOU4nlsExwB+t7PTlsDfStZsDBqFOz
`protect END_PROTECTED
