`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a8l8Hp1TwR27EcUUrW5YbkzhR/KyQdExob+vWmyxy8ygDRvJB0VXB/AtsZO+e6ko
4VaE7/dSUxktbXMTP+K05aeV2OEYpfDHjEhrf6YtM2Net9Y5xRJxv23KUrbZm+kQ
APVfErg4/O2Zo9E4RW7XCasu86RoaPjwPfkh6Qhn9cYeuDK15w6LT4WSizcr8w3l
SRrn/qBWhyMlJ4t2EeonID73kcRm4sRoZKW2vbbTv6m5qVOsKcv7dMeZIv2tT7zO
6et4lBR9NZy9GQVAl0xGSaa81jKRtZmmtSc9GvhLYx4Hc3/DJ69m/ymQruIjvSzc
TiCAu1LnDCop/j2b+gm6b/mPFFTItWOuHcuStaKzcAYcSpGCKktBTDUH1GM2oohT
yGt6tfLfURxjCX/pXMXEUSEc7u+AlXVKY6tmAiDeH0arWEPrVrPYxn3ligFInb7o
zoTjYyu0PsUPkEpOD3FOJxE02d5t8XChjV1tdtuW9VjIX5EYEKcNrGsDBLURKpBO
OxxC79mt+0sTpNaz5Lb1yJ6nnT0QfiRpE9mI0pb8LB71POa9YEcqlFc2g2lRx8by
Zfg3/SNrz68b+hbbJ5OUF9L1h0KOazc5WDFIr8axxjRVlUSU1wk+Vawz39nedOuO
yTZWKvgz+xrfa5Aaqimtz56JKgCIiwYyYme9CDP1hX2JMAA0TZ+VH901+P3iNB/z
oPqIR4t32zAXLKnz7f7/Tjw5F/eRKzfihNo5LhASWYuB6am1WrukdHxwV7kOIoLg
+ugM+dcg/D2JP7raYmW6gt2j+nfLVR+LV/I2YhBY27nXBk2U/vBs/lwA/lw2aEXJ
6CaL9/z9u7hnVx39kdbOfPsmEgsoyLmaaJu9p8rbRo6kIOUVRYZtsnCG0jcO6Jp3
wlCc3fsR8D7GDeJo1599uwFGYJFCMvDRtCYDkVIpY3rxKvg3OdESbHOMQkYcuRh7
JbPzAmfpyPb9cbGBwEBZi81ghlWgnCXZNVRNMoYjGwR9MLhVDkkvWbWWWBf8TZ+w
sIBaHkUMzal3A2u2LCDndU3AzJ2GlvnXt4BnscJhHPj9qEv5ChdlTtelf3ZM2UK/
7Xflq4uLe8p9Lcs9CHMnJXHgS+6Afz3jart/ZUWC4q2OUIxGsQ0wDph6fyTlRfIr
kFMedK5QMDRkDOTDZHWZ/+vrZMz/BXMtnrKDTkIhqbkXkGq7V2hjmf7fA0kHwY4f
wMPIRoByWnR/83Z/ER8OpVUwCQ5X+KLC1HmXViYt8zyRwVTvL3dUZoUXpQVk8ct8
Wj3L9pZEl69+7t2mVzypznHjs2rMapOitoRVho+H3CavlluAkQfRGC5IEIjZ9TRB
RraYEvxSF9x+Naei0LeYKg==
`protect END_PROTECTED
