`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycmZk5uozik2xbbmZ6VZN6rIaReXquzrHlTpYXO8Opoh2525OrZHap+xb89yBrnm
MZ0XjVWBW0hi5ELv/Q0vc0LMe9zak2YAwSD+5HHfmKu6LZFUZ9QzWp43tKGCnu28
lU6Mg88mAKXoXJx0duL2ZKXNM+h62CovSebtEQHZFIGIC6rt6c1T9fRODxWNcQcH
omVAQFKpD1wlwW3U362kevz3k04/FR7kvVnTk92fzO2UHV1foiPLAyEXhZ9YQQEc
4VV0zDzHq9WWXwuNhNzdEZ0bcFnMPqugc5Z8AMnt3axweW1K8PCvHXHs8/PapgBN
yeU1sC6tRAc3Tk+kH3tXT9FXF27koBFkroF22VVaSDeeOvGORqUbF3/HvY6MTBOg
nHr0A32BYcCiXpf0ZZ8OeQ2zPRXYBN3OZ7ilwvCspBJmXFB3MMIwTpsQ6x3Ktw24
t43HYpkkTfI6gSEtV3KDcJ9UuynqOlEuA/TxuTzf4zPlb5Hx3AMmCsRxQOvkyJ/J
INFvl1wjEgmrhfpd4KSDIkG2qG1gn2vdEasjnd6Kj+nUkV4s6qahYNSg9NSvaZpN
UmzUP/XT5/UrH/vt0QJ7wA8MzsTi47Jj/ywbvuM3lMiAfwaPnspskjFAu85svuvz
E/vSA4h6XtT159Kj3fkgDOwfjbUiQOVpc+eCXp7NfAS0LZ66yjStuMpIdzRI8sX8
yLv3Zy+8Rp8GwsAqVpJ6xQh1ccVIihngdyVVp0CMhiB6M7kw1HIJeoeNe+LS0BYI
q1qv2UmcYrd37ZnfmSOADJCy9wwVZ5KYZUlgPnbnlJ9WO1IqhrPHxnsj7hjm3OoZ
oi2QczmAYj2IgbHRluBUXEPu3/L/Esz6+gYzll1TbjzILTRCiomFlAHktNKNsWJ3
xVc+4Xx1E3ZfQbaZdh/d/uScthWFOcbWKUX4GzkOWjpLi0HTYTi+vPz1O1wGKMxk
fqA7vwgXEr3sM7Dsh5m92cn/+PfQNI95jNBZoJTbPnkm4jXESlh8ArT7mzc3cS5+
vALbUY+Y5ZUPbNQCkpL5ignrA47Qs3rokGzhHAlI/q+kuW6Te3LxaIqOCsPAHcNz
LvjGxtnhNwgx6tffi/ziZ6WprFwhPvt+nc58kKiwnV6alYp9KcdTWwjcHgyIeJZP
1b4HpH1JieXzin3lbVnm4zm5DQJCdEpjxld9/0NFbFWXuZ6eRAvhTZJ3ZOdLDke6
dAeXakjHddEWeDaojUAkLjcCip1rfK2SHNBVI5U8tZaMnzwWPbAbkCoOxaJFdgg2
GpeGL9q7gxDRMDFB/hrf9df8xsoAWkbFjWp1eUnfOQvUAowo00SUzxgZ84ahJyHF
8yp4mU8TsLiqht+SZypAAFgdKSF/oifMcwNHdPUmVy8UhH8OF8kGUJxTriXXC+X3
HrCGBP6+7NTYDnUtzeVOYAftQm0KFrDo2l/TqzmTyGIzK/9kdhjQdv6VHtdBGXiN
YRn+eOewATelRYdpGAb4TupiJr1HCSEciEe/XVj6PHKfruG+oJMCad1marIvngR0
Ej5oDuzdLC/V4T7DYGrFCmdUE4dgw3dZe9U+dKgXTewf0C/7kZAHSmYJm22jGJaP
wj7x0H3Shf0hePCDPrqgle1ATRn35d6ep+Wk2QJoszi1sPsglt6wMdyiTuiGwEMh
c2OG4icO/AJm1VkRZrvrZ0v7udI8PuTp8tz6r7r63eGeozlLA5eGgJu91bjR6umM
D4pP3SLF/3gdteRyubO6hflaaPGcopbYzkd2T1jg/dd4e//YozseunfC0OniNGd0
EQAzAJANNm3a/A3Yxj9CmswjPkwcpk8VF6vfz6c9ny6vtt+fK38tRwGyXgoJy1jr
GTGIQSRz9ntF5yYxzWVuvlI+xJlrNhJFkYyVzx+c3qGwdlficrcaMo9gPA/CHzFn
1DVABc8K+8L4RcFyxJA5Xtp5E8Q9ORF38vBbrmuKAUPfUYElREUsRk0TV4zg4Iak
G2D9d8QlQkBY+rymBVSYp/Sc+GBa6sHAxhDcWvQizLyCzce+oR4E4yROVuGcjxnw
xXjhNxnvtqqVpmzpqeXwj+/M6pk5dwXs4pBelmWQ4nJhM2qGBhrrcM05L9UbSNqH
UKvbQJFy9rFqIKRdRRHbkec3lmXawlbBpbyfsQF1Rfa8NrLhJNvH9jHuolcUSkC7
O39bcJRtCoSXSoAEUasm/bwK1O92v7CaYoHNCtFUXEAdUOeRHWGPjWbf+N4mH4tl
LRdFRklhPkNDWMlUIMrKig==
`protect END_PROTECTED
