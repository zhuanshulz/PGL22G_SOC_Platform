`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sLP0TKheYJgGaHZ4Nz65b+rFaHcYcaRmVo4Oovkh4zLYSU/6ltHjhScLsNmv1SAl
1WBVmeYJ4RDWcfH3XN1/3aOU5NJUQTCiRwN0zX3pTp/yU4gEL6r2IWWqGnHLpiwq
s0Orosgy4KtK9xozqfpMMW3arIdbrf0XslUog1UTgc3hQvpgpFRoIXAgE6fGXcHI
dOwebfwHcD1INAorlzkfhvQxK9QMWISwUpgyfb//BI2Sygmg9FjP4Z4nT54qFQek
Z9Xjpt3lNeuxBg4TgmBaqyCD+FVTrsIJ47JAWjC4MOuI8Yc3cBhNubUZaJW4Budr
VfR2OnWKOGFm9wi8kMKaWXr/StqxNtfOwEJa+GPNfyGI1KnllSzmTLMBNxvZ7ouN
jJFnJYEJYT/HhkeBm/n45sQ3pBjf7PsMJDwwrx2k5Jmq+V1iVVTdopZN9VYRjDgS
CoCeC2Lxm1be6GVqOj/ygxfn/ifT3nJffkkq4XaflK+3fWEbm5YC0aV1i+7H8KRz
0fylDGHI8OumfZsfgYUtZvJsA8SHIpcDqRcO0iLD83QShgMTFFu+1bK5QixxJ4Kd
d0SDkrYv3adLWi9lJRpDe66iAXYbm4KeSoSwhYaYdkKqxKW0EgMS/6a0w+KEr0jH
3FveQ3QeZmTzuk00pIIP8fFD7btyfmF0gTEmtmPTZFj7hdqBrA0dv4EXLrMYvggq
Dw07yI2J880CSMH4h78yJ0eGjhtqtEptioeexbDX1thAM5aMAGcCDU8XjY14kgPd
82HEBD7omEZgs5f2CFAS2utCwRFLxfZxC4Fr4rHurKp6geZB/wRMyaOHudlasNzt
Jt6nBaQm5f8tgR+8QAfIsHVgExBoH7DTQZwJ0BbpGPb8SYnvzir9UEcspn0gn02y
VVwf7oq3qGRj4/mSLAmyYg==
`protect END_PROTECTED
