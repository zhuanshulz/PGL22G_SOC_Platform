`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uiVEf4NjEmxnPr/fv0TrxtjWKuZGkhCylyU5Nl6e3f9j1wUTT0FuCy/sygz71W0s
rHKBzwoGD/qQSK5L7Hy66OwLW2DOaj5rk/mTQN6TyhOeineifFUl8pMkUPZlQyOF
2HQ4npAUlTZ2fHzGTD6+HCkPHTo9F/Z1IHaQbgW5s9sp2gC7cLfyPX4aQbsS6xon
P6XI80HcgVy2Vg+SPSkGxiNBXJIXDfl9unhfJxXx/XPA7m3RNlPPXitEDhEn6xqN
w+Y/qtn3JLbzAD6tO3DTOkKEgz7tKUVxhUwKRoLq93mpuRZdehcHdL27O/3PXJRi
lsW2z2ANEA1B/6O2pcYM2uzAT9wLb51xHpSeGp86DJ4cW5XNT8/wXk7rsRvGM53T
m/znKoWVe820oTHmwqShZUVPtP9x3m3Cv6bwCZvtQnfxk3EdzLKbdcLKult61fio
TjB2+WUCLg3/ncP9Kcw+cAbs+/DiaKG6/iHI9qQVaSGIKV7viQgTJc0gBGtahRnC
rpcI8e1dYs3S4YVpT2GjEJ6Mgiz0IQZElZCNmp66K14TD/K4pWDGAYry+Ibzd28R
nEQ0YnFQ9TxTqp3+bo7LGcWEbwjepPz65GN3D9EO96m2OvapeANHsofZ6o34VFsL
XMhYq3mexg+VfaQuXMcKR725+zHyHtL0TzinOwxIZp/68YnlERIG2kP8x735Dveb
JYEtQ669JtieKON565yttbCJCwOyxtyXnt1jWB3nOB3RyC55UNzNKfo+eTCGQXYs
biWcU+YcixbKQhUSVM/8hXwGWuYwcg+4gZiRKAtW5sDfxUEo/RisB9yPxjyZYVC+
azj9uXeSFDejLOQJVR+IlZZGDcKzTiqjWs4Hy0h0JIdRef4i0FUn1E0rP7D8IB/7
At3gQFVagbwsz52fBAP1CChwiMcywZqWOcxwv2nYT/KWYxKuJHPN4HmvMT7SbyZa
uLGhpTrMOpr56XDzfcOhuirsF72xhkDyTEwcOGY2TbxM6y/7xJh6wqTp/RX1MuUk
HsCYE/UAjCUyCcDCLuU3A7mpOSNNCj+lEPUriDV/GFlHvBpN5ImQ/ICoyDS0iD2U
beJrGELI14Id7u0ukPmDtUxsLfWzyf2wCXhyXpyR2rEK7Eth/7dPfmZgblaOfgRc
hcIygFcxHRCPrrcvLSZ10eQpsvwVYV/f7thT4XjcbUj8PA/8b4hAbntnyt/AwdOV
n28EvPBNeYB1OOxzFYqMbw==
`protect END_PROTECTED
