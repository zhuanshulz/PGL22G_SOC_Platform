`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNA6sDLuPBjbqfDmNtIHCU6etYUI/Nar47uP1VfC4EtF11J6rUzvEwtKp7T9G9I7
7tV0cAG2BY7uNxCeIviWjYOlmEnNV2Lw+tXyvj7jB/3kWsz/dui/Dof9qq1Ncvxw
5jvPAxClLym0ztZ9w/4Fi2c8t5zlITixGYIQeeLjwYw0IyjGlLbySan+hdm6sZu4
JwxWVqMF9StuO+geVvkybvz7G5/l+HA21wui0B4UviH5ruDTipqZPtto9iKbx+6E
CUmSUptn+u+thk80oL5c/9lXK8aePtkJvQuPp2k7+L3KqbGjjWYRHYroLRofJ/Wk
3Pu1dCH2sD52mD1hQjELqcQ0U5M6FXjPTE6EdlxnucvBVRoexpQ0Yr5wMzFR8qQR
Q+W1pAPb9pA6jMKkkSrRRMftP39Ae5UZGvMhLzmWJvTjKGZJdFMkhmPIEM3MRhca
W8TOufY9oQROgwd8FWKLKFsT3KF9vb73r7zYACKFfA9noUGTJgcKoy/PSPzL9+oE
b2UpSPeSpYCuu0RPnGl9ed9GQztarw8rvh3oyGlNIk/RZclHjUo/5kY5Du6ILSBP
mPEDhkfqjRrpo83mOmDF64PETNpwu3fXZpm3fkHAlvL46FMQw9CFD9Crzl9E1/wn
SReqjcWrBxeGXxBXA1Ubc0u/hYbQEjyTIuNaj4zCR/M=
`protect END_PROTECTED
