`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRBjybtdzo35NoyR/41MLhLx7esBPLenJsUOF8MDtiHAwkw9e+4+YAiK1wWj6Gik
JxbtC42MnOfaKWCMuyAesAQkfOa/dkfvC8m+jmGl0DJSRK/nmscLsjSZYhCpza5o
7wfHmucEyt8OSX1gBsHTkP9vSR3ZJ7L1KZ9zLnV1nrhCgb36Pk55b+3Z8GhjJ620
S6H9W5VKSm2jpO9/o9BQLkqToUYneRb4+7mOlgcEQICPrdXBQ6KlKHxaW+rVybTL
bNWse7+SAavXxtIqJeM0Glbow0QS7m86Wj/k/FS2aOjOMrt+P3pIu37c1fj9wsUW
oOlyjyuAVBs3hGJhGRrbqBZq0uK5YZMQRTeo6PEUB3T7VdgpHsiv1SIEkt10ugUg
7/QBFkcT9CeqWlW8nnJnw0+Q7bmT4mymGX2M/r2I1Fc4mmgR9Iq+bYHLPRDEIhb0
w9HqHrf21qUI5ISH3IVq7LhEGWZr1adSZSf356FhGGW4aOevTAz+ZTK8WMtf5nnV
ieiXuPwGwA5Um12rLo9gtLnm/v2zeQdORU3U3ZYpOwxd81FC6Skse/4p5t7OYCQn
IU+0INpvLmMmFzZg4QJ+a702zNAEvkiQb73npg+TZsRM9/Rthx81NmoAGSqU0ieV
bOCOTrqVJHQYfY5io8DJep7ymOfBb5goiTxp4ocfcJluXVtsuyx6Og78ds0DIkcx
tIiXUp//7+yMWO6+YkcIH8BwIAScCvm580Vyu2wO+pXZSvyStvMVlZF7nNhx8XDk
xXNTcyGUo7x1+2uVsbqXQei5OZXbZ8B1IQkDNkL5kADlQrHYdI5U81HQhRrKJxa/
zMK63aGa6cnTauKTzrOANIMWfsTSkCZPJG52VbBfMrmni8eq3o8RlNY8hfP5E10r
Rqt4WPHzer0cDhpr8Klj7Q==
`protect END_PROTECTED
