`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpwsMlb32hZykfUsoS+dL9KDDX5zoxA8eFxtcSv0VFDKKw/m/lDdIAkaRTHROIfJ
NaomSQxLTCAWDWnY+822O1PjMIuNo8yTApxTA8Yi96Y2l1GguauD8C8hFB6iGb3b
2qetszn+RTcpTjQV+yGK6QnCayLRsB7R7w6wqEC/k8yAB0f/cHMMBehGT7reUD9T
EdkVolxfRDOBAPzn/5TqLLwuFZQCSSbWDDgdg7aufmkmOK95o8nJhRroFMha80I/
Z7kidxsv3quyedX9Lgf8ihWKEfjCnJU9b0H0NFbP7EWK+rPhAovPBqhxmYqIElPN
0mOZfAeujObV9lf3Kd3NFQ4kuo9WX3L3C/lBhJyiHHVFdu2hxyG1sOqFMFxR+989
`protect END_PROTECTED
