`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sse2hxEJoHlHjFXy57tnbQPrn/59lcGv22er45EpiD3SFUGEYRCMm5awQ0An6HGx
oHZ6bHzEQJi4sQZnHm4jiPfh7Ki0CCd6q8+tpN1uV14Q7ZcHPA6JmOfl3OpTGxOS
KK1cJp2iYnp+meLEPs4OMMYJ1zGI/psw/t2tRY+j8f4BkIhgfCoHMsQtYlq0YJQt
intFNWKfP4Q0xTeVe0Hctv1ZQbMgtrSwMYWp6P0YLKpYrvvTVN+V7KnKq70IYKz2
Zx29YgZeOxC/0VGozI9IqhMevm/W6OaBwuSsXOY026nOuSG1FT3MAaMGj2/0pRwE
YTkujuj4BTNBgxd5IHUROgxlpM68/jzT5kWQ7B806XJNIUOqU7B3ILJpQajV93Ia
1372SKFSxvRx1/W07hmzRhZI0IcwX6QNP1OEIpscjxy6NZWVOxc0toe8Cor3CGJk
aLZ2t0jB+7OxThHhUuZ7BRUcTXFjsI46u5GeN1bhe4Bm+JLaXrhN+jrujS3y6u77
eu0CB9g7r9rUfcejyUXmeER910znfwrTYcOK7xWGKbQV6y1g6cKvNmlABMnmAgYz
wVIYtpYzF9MKXJ56ZoNfwQM5xdl4KmT74LeQOgIMdTaFhvBVvf34QSPM74zuHqT/
6RxgbTKN4MXVHJVaLfJl2WQetOigJWyeSQUdEzQnnwcS+OfN0lTRoA6zAUVWTF7r
Rs4iDHOJe9t3jMlQJCuQ04Mo6+3tVCNX/O7VcmexocgcxKMC2Wm+TEF9N++GVPfQ
L1N9pB4yx7Hj279DdeLfF/YyEG9dchaFOQ7Qa+lebwe/xaYfy/vjEQxDsPpw1lMQ
iPiCIjKwEn5GuHgWlxFYM0gw874HXHmlR9t9PqmsG8AtnjOS2FhPDAbSZFBl3X0i
zMYJTUYTOQ34qIji8SAkHQ3f4jwncG0IHv7rsyZjZXuB0KjWiryz9EciGkU6ZVj/
aGmCz9XWyhTCERFgGU7d29ykVB/l99hfH9g0K3SROATURbclYrDWalRb1+AJPGOd
P46ULCK2qAF/Sh4enTJsP+RIOnbmyT/BxgFbr04b6YzhBEa8fqVP20Hq4i4/9NVz
SZwMAcwGKoyRi/U3HxiAz80QzckwKNIcuwqOXA01WQvDQGsqrzCYsvLCbxGv0iSj
JhNYcNb8nxeNFgymtj+uU8kYsrmzN+3zvgjRI15x8Kyn7PMsmOgCQji+WwGaL7qf
6cFLxSrR/kW3cXADbR3izs4vfoelB+hqmfY7aGm6cNNiglhKu18uDIUrTQqaHPJe
Rp+MA0ddPe9Sc8hpboIqwIesjWdqJEY7+mLSZU/IGTM/UpBdctrqLcD6EhE4ATjV
bdFqPNDZJvuCoPgWiCf73dKIJMUdz6+e7r6EzACdVCjtXMeKs8TfcaG2NhW4UgLD
R7Zno8GdLXo5eobdd2KW9iO+rh0jcccev0vGudScHxeBrRe+HnzCTt4zb5Qe6fwy
VhrN27CLF39vUsvHv2+f6x4YgamdzuF1JbMXO9+Wyxy9G1PT5iuGT94FubuK6aMt
4dt61+WTTb6hOjuv4xJsCCdI/XOzg3uZ/n8pN2764Os8/i39YtA5U0zObq+739A1
wb9aA65qqXk33Y/6E2em4Alz3bmmRgBQCSxhDy/+uG8MyrDAIOmDvicLfNrFCnPw
8z7u3i6S0Hc23FFaf8GwqVgtaW9253ADhAm3W5ykgJgSzWSIxY2uUBEDlRgkl1BI
Xc3q/O+k4JueSMbFkUBxQQte1+djqTqeBQIseJ5XGS4owOS2R98irdBnVahFWGni
yJMHZV0bOz8dgeGwmiI7iKQ/jqZFVcfdz+cJklndvfK2kOVstZEkHpEczaUz/Rww
F4t1IeCzbZZSZkDglj0BtvPPhJuAMxbv2utIKSss899lcC0kGREg8pVeyR/PBgiY
oHkwxapIQwcfWlktTjnREYzpaFm8uVK+DmnGXgt0QiBqNc5AzvvW3aK+51zR4E0L
QRCJQ+HrJO+46ikQCvI/DiZnALTy5o2T5ZTaEc5QrlXsagWM8uNDh+hL6Mgcop9z
hgluT4Egh/mc3qBV1xYJdhVnj8IsGYvS5HhlKMsuQod/WDHBVDEow0Uw7n01O5me
j2EGljyp3TvG3ipI754ACifGHtCEn6NvNjLwM3m6WCu440gecBvVQP3HXSOEKXjT
CQzoRTAIXRtRz8+TXXaFc0X+ovTnLqYdrc5Ax+JzgzFXoMi7oLEpHO7bmjwhP2M0
fAAKJFxl7+XqgitxnKAtuIWdG5KnZN9O6ONe689NOG1VRd8dNy9xUPL/eUgcHX0a
OaIVqqwXuFeXkyhZFiA/Awhp/driygISQUrIdKl5zNll+9sm4H0EOKWsb0EdNBhM
cLNHyaibEWRpYRQGEgk64GfzsG2LhJo8vH4LmbN/C8OC2dfIMwL79I7KlVOdAehR
1Db+E9aX70nszAzt81yWXnBGEEup470sc8uUMjzzYRggUwYH23s9Qk5mgAFY8w9Y
8cJunTAKudkbHLD3Y9QrtRnfZ6L0vIQB+I0t4qqP0WZsonmQGKg9yccuJoH3RwkO
H0H+70b9bGSGLk8YvdLNuj6kIAAiKtXZH3+M/rLTBerwJJMPGPclcSUzAGJcAWUB
KwxLcAYkwTt2h57p3woJ5zUWTpNkbmOqSx9PzUQ1ewJbyabzFr7GOnL1xkhSoURJ
nYgTqA8EfLF8CVduEW2JX9QjksgTVxpk7/Eh2Nqza0ytSTK6Lq8eQHLwqnPVoRjr
kYAGyl3Lp7U9zMj4mj2kSKSEhlygilwQpaQBJCpHplKH9X/RvZ5YilPZ4xa+7Btn
zjzw0BuEwfHsqTj3qKgVqSd4Hj+x6JHNc8PBuZUD8h63ipPYDDDMJpAZUU17mAr5
ES//oRgmmsBrRyCZD9nf83Teer93rykC4KjtIgyLYl0DyPOUhXYFTnYY88R3wRjI
ba6ogftnMhoPz5Q1Iq++K1BzVwXJhZHlKxzyZ3j3sz4mJPlNlt/7dFnlaLiCaVpx
H9pO68XMMoZrElahI+uoLbz2pyO5idgKCnsYqUus5ZGYprqirAk1+JUB1FE6M3iv
IE5ltFtkdLx6wQT5chUqPrjKLO8ThoRGIgyiR8o0j8V2FvqVTbo71n3C12tiC5oF
S3mTMFwbZxiuBiA4w6xwKO+Pf06qElYVzsTPftADyrE3OWKO2vz3EDytefxUflQz
Eh2GZqhDTJT5aCt0TNGbqcMSLOEsb4NddHNYF9Xt8h1PjZshAVNVQsRbUMR14qVv
AR1eFmKFcpzUpDqvP+DMoE8AecTz89jgmdfrormMG4KCxt0bRPVsyqeWCIEP+YNa
fKFgXmVQl7Mzymbqa+Q3x3bYdbvJEojVegPfDXbC7EKTyfPyz722te4W/z0AsMRV
ChyWiI0FqOe2/tOUVV6ic/z6TInHFoq8p3jI7xqpV8kFgY2jJpgFBiT89YQ3TIMX
XIL4mmolWRgP0B03QclHQipCKORy6b0i0DQqdB/vaXqJyueAchGWAB8bZqiIhtae
Dxu91sctBEzMibqIfWPN81eew6PHN2qEeIIZ/CDXHoVgibdfwLq5oiJqWoHu8HEu
Sc5/AGA2BD4awdmpDJvi64QuIVWzpEOzaTQRgbesGIxt99gIqz7xiInPl+HkE1gT
6fEhxS2gA98BM8YunNPZUElw7xsCd0zoqGBtGh8FHLyV73R3/AjC+bbEk2o8DBnI
dMtBlWUwSrPYnt8ywgUsGO8gbgbbCEyUekgLmjq9SXF+Ib1dUwVd4Jg8QT9p2+fk
1/9Oek05DvIK8EXUzKy1mz6yG99qHYkL0YKV1IoBDQP3qSRJSKYukVuFc48Lpobt
2GkzEXy0NktfYCtIZ6BoDC3lOk5Y8p1Mr/La6hawp+7HO/V/wK8nvSB7zZaT/WI/
+fTAoWAtWjOPznAW3qhBLSSWWvxNGdrLGk7O8woIDXzhIlEzrVDKDU33alAGbeKb
Wtp0oaPF7NJr8cbam6099lDBUtt9Ne4W4GhN8JNxMcWQIoBReqPMGvJVvBO1dxek
8ApYL6CfxzJfvR+sFMmYFgvuxhIrsIjQlOx0UzO032mrUl72wkcJhHb4hVS/Kk3/
T+Wy686YVNccCAF4wyyW1fbYf5ct4qKvrSBPNyUOfFRtZWiVuW1OQ0yqPVIwc3ef
FKzts4qoaHUn8d812CH2CCyXcEtFPqvj5DE2FSbo6Ij1hLapUEMrwz0OsxFs30C3
yewZrY292sGtxDf4kUytlxvtkKOEVrNn4pru+d1VSKZf/LeXXq8XnKWDCMNqW1zC
oe4Z5szumk9Cz31SQiYNfvw/v67LRoHd3vLNMNSQBPhfZQiJcJVcEJlNa7T3BRtm
Kdku5vjYfuCaxwGjBfk8L+O4ehZPPAJtlT011YIHs3U0Mk02vWXiWWPrZ6EFBMyi
59H5YRWn+4VEmsxKqoiczVauSGXX2/4BJhHcozvxRr50sX4z06bFthBPjRQXGg8h
41BCKhQURMBFJTNXkITaWgFbcO/M3k6MVQhqOjv0vGut05YpxfQCKfOk03Eb/2Is
CBzfwyLAJFf2yVS7a8/RVOJqvQJ9r5cuFMfQvS5Kkyed0QfKjCV6X04H++78jWY4
bFwwFjryv/ZcdbRKHW0hN1QCKfHauQRWnMvro+CdLfWZ1KAPy8ok47ABRSjsTAjp
3A4i5ekuhu8qCQV6fgJMWWSxJTplpp5A3JKBSjdsbY8FUL/gGpRG0yx3vb/5daPd
2G7GQQdiLz9/uHzD9XePD0c6ZCwkOUgmt4NLRpkanUybKD+NQ9KygLDPqj1BwqFY
9ishWEZSRa9wHW42AFiiVRwqvXEKH8XbQTFUerlmf1mT1ab9ZiRnzvqShW4rcKlo
6eqjbp1/I8T5zPGV6Eg1Gu8ksPvugM0rYHRA0LEU7G0Syn0xV1BGAVhiuDChqGBH
KelQaPqCAaRluYPKMCApTdj63wFje99+MpbJUn/aOJmJfYZPTbmcMcCrOQJhob7h
+SygHAvgGw2Y20W9kd9Qb7AlZfECGK8JBdBpGxHT7hO/fswPuHjUvgpZkjtaYE7g
RGcduhgvKT7XsT05sOVEbX1SLXbwlUCqukoqgt0WMxbadekBewDpAEV/LVJd8De0
helg197F7IGShw189yM7Za/4AB0x90sXOq+tBR8m3ZJXtqfKHTDqqCqfjI9IkDBu
PK6YRb30Wh0DaBNEqkgQ1ylECXNqfwiwFuBCrZ2Ue4T/ZzJcDvfyaNTqqYT820nC
wWccyZQOVQWQuGnExlH84kKb0n956QbUXqWpVrZbmWz2YIYui6y8Y+JC5tZ5ole0
qjubZIP3bKa4y3HDYjPwCapTnYznY8Zyg31jPfVdPsv41/nSDD2iNRyvaB1QuWuq
sundGoHbvROOdwKKXHICLnt2rxvlJam8WewmesJVD9/gqteTCcn4ZnIjOkEIwsOZ
Yfp9AqB6/bdO9oQ7TGgXfOMlvo1TpMf1a9IaSJTLXWy7eKbD1S5azr9FOyDgVRv2
0jORCb3wGZvgM5pbDQy3330b0DrEFBkTpQi9DsXJxWPREE0QRsQWJgFwZCsPISK3
j7nn9zIaUh35b0vergTPstydvCtpGpICe/kGQ5LELWzlu6zZvgquJ+LC7WS6/AQT
vdeArHSv5NuyCk2b52kEDGBYrJc/KkD3N8JFWRVzd/BvvWBjVnf9u5ivatu036fo
bn4psmXDIERDyr8p0yn74/oOjUTDTf5NV6P5ZCAHspuYtlU6zFtf48NiVCX2Br9K
rnP9GCawJrvhER+fulRQ46SytPa94buDjcfo/U/chizaIXG3f0D5kWZGDn9fPAYa
wcCGEHesmsue2mNNVriN2Xc3xWQdWG6MDtcoAYRWkXO8nXYk6/DP3Y1sRFxS3swC
wVjxEp9VQu7/zcCC9OtJvY3DlKmiiexN3+rj7xp8zmqUgZvWGZwup0BEg0BE1WFT
/vusVpWO8wHmApq7f69vpqfvyg9PmjFTYTxQ4QZW61vIITkwcRdnNE90Oy6+RB1D
NC6sdM0ePl9uRwdGd0BcbQIghxThdIWPzOPrc7XTT8GCtIDDB7ZK6fgtRpZz0plo
qmAFi4fNUYfg904+NcgKPmjdQgV31JIaaxO2sNnxf9qRpAbHNqMpuH/kBfu5WQiV
SoQTbsv7NJ6cpsZidoINQUZK/ZRW1JEnh/6WHTBQ7p35baZJcW9n3NL811bS17a9
j21eHy5yTMe9aLW2wTr7S6BDIVZhIKbx7vOim7ePKHO3gltN23bIUz2C8aYDSbad
9XaJI3eMASIpZ5gnWBULU9xBmvAuHKQuiCuxMzCktIvXFUWbEyQtaU8h7MLsLWEg
ZQQsTd8CD2lTJVrNQHt1FZ5cXt0Z0rqrNt2ttfr7t6GXFuRb7OGNwLUzXZT8ud+y
lQXjBV/+y5B+Fj0HhLCpi2F0wjRQ+ce9vJRcD0bYDeXVLYmkULMd8H+VxbXVeP6Z
0hOPwtRnzwvEkx3HMgfOakzrMP0dru6bVUxkaEN7KWQXfrUfegb8PN8YJiLimeLT
NijFRINtSN/VndVUVvVNRKeYljjYBYOnJxpE5QQpGBtKwfLk8fBw1qI3sFKm33mj
PZ/KIXbBtxJxX2gkyfZjiJA7DmEUCP2eTAwtg5ATpiC2JXFH5haILMUdo+VqmCPz
NJmXR9lDsIs4ZbBr1CnlBJHO/xYQyHb0ToD0+DZN/6bsgeO0NsmaR5nYCHgV7SUo
1T45+o84gCt+6HzJ4FWb8p7TDPwsw/2lgV1Phn8yBbXAfvlA5mIxTLhLayBivtwe
/Ix70TUINkPJB9LJak4G5C2zxJ3cHPU+hACK7ihqtDEIpULirDgrvwYHl5Owbw+f
h+u3tIh4JceVSuw+B8rHypS4f4mdap9uzbcdAXX+cy+HYKuQrnT7WpvoXp+gTvgQ
xhqOnxKUjAgsP5wV73oGrfThLRST4miJlWrVC5GE3rq4DGjx5HZxs7NiDXb04mBV
xrD29pEGqVx+k75uJcRqx7NhXhvSkxYDc8gYCecrFkuyMdfQnAqdtJqCyb3EqhIF
DhCqW0pYSMVWpj9QuqytFtexebdFPvg2nOGUfLLnisnig3gLxAcODxm/KeNHpB0X
pwNJOwVEIbmsYO+vhOCP3IDsdmuTHFAFrd5Z7E3mYtNOrJBxKYLvDUxgsqotFq2Y
MmFvEd6quw3Gkucah/ZCJNe9T/Mfs2oP3NxGgxVQxMQctOggqKQS62KzXd7db9yD
wytY55H2B4gqx1Yn3ogEuCSGGesDiNqL8zIzgVQFf87Rw1W4zn4VPiHvqpPfraGW
ZJf46GDQY9fLEg/psB+BNLy/qojYSG+lTUps6q6XPOHvLrssg/Z9jd/6uHEwqYMu
tKvvgvAscjnyuYKf3D2UI9SK8D8kihKyg0TFTyqMp+HMoQbe044wCzLpE97NdDPr
6CVk7aAWSY6L3zLEwWctLffWu9SXrF2nJTRnoRini3FuqG1TyMf+eoXwN1UBZSI2
x7aqaNizhzJu4E1U7Lq0Kcmd1/3WWT8fPokT+7OHpa/qNDISWLDKu69ktIDehOIf
qfz7vk7KJu+SzDAazHOgO6Q4B08Q4gtJMO3ejZ/qv8IMOon+p7GV9aTJgd35eUBQ
CZsB6jUuSxvAPVWCqralF+EM6HVY56/cXZ0IPXmtaPpiuEw7BvBZn/2QXdNU4RJF
Ep3CakryTrazqvEhX5H0T6YG3eiNb1l6KYKO4ItmZLgidVb/O1LTmZCLMWCTfm5p
UneTj3YzVjn18Rnt/uAyZT5Pg64ju064MP1B+ViObU07/ilvV9CKJxnOi40Rp622
MTNx55aHL60xX+D3tfXOHp/jNA1e2nrevPRQaP1WE4X7Dmh1Ae6T1+S/415FIyKD
wE2hmazUeoiNygS/+Jc+DRfvZAcpfOQ/XsaxjIePc2RKJIjpbRSneD4DRFk5I6M7
jTioKiSJUqIIvYg5090tDHghuv+rBQmHOh2ZUzzGTBkLc4sZLR7mI26I6SmhvW/8
0BF6KpW4lLVIo+LO3O7KeKYK6GwH82y21E4YqPJ0tnq8Ee+L2/Cf5CYw5d5J83Di
zuSRXk5lQTMXUI9sQm4kj4DGpzqDAFDUakDi7uDfcXohJrQNXCyNIpPwgIa3sK3D
+d7befCEPAv0UxhF8QLKbBNfSO8AkjTMi2TutpaK+zgDiExMv5Qmt39pKkyglFI/
tXjEZJLUHv5n0X2kvHYedtpsls3Ggz3jVmU+NlgEkZYNTXFdqFEi98U/PGxYU95m
BFo//uluJZPnBS+vrow+3a+napBX2drD54hqOUU5SwTdENeXsbfcRRfluCpLbVZG
PwaR1V+AGXqqEoshobtT8iVPOJyXKXaHL7wkZaDWcczYOw6Pqe8vCpxvyhfbpo/a
OVJ1GBFFx0ufNcjkBm0VbA7YZtW3GrVeJDx1STWKblzRKmZ+K2LITcJ3/qV5953y
wac9t+AnFjokP0CY0kMwkSHRDGrJLIQGfD4X0zKcmPI1UysO/HzjID/4k7IqF9MP
f3OL6aNgtCgMdpbe29xt5Ffca97FHbd+CGGaWo9IPxWLJQi1/ZFmGPpyRlegXe8b
MZQFb/cIJ/NRgfAj2SoQzk4AjOf+SUKpiEY6DYlAg4ogi/Ol1y3/5kM4dg5i8ajg
qRRjxRAbLX3yxxROeFDmA3FQiTq6w5/WlVGyPBKNbapdfuBvo0j0dU/LRhFy9HQ0
0weAiowkLPiuXKDo8wjEUmCca6pmPQrt4C1Hu0oNVGhOIkkUj2nLtMu9Ev+lnpTB
PXefwB4YVL+J6y88FyAsPmxZZYjtv9jL2sFC8MpsBiRWlbKOZWH4XnlwstXo+7gr
4stzMjI7zdIF4eI33WXdSgRA0qmWbAbmXS97Iv2liYUBSTl9I07k7GuPu7jPA+o7
6vJ5VFhy2Q3jrjUzJ5NiwW+X1t2kEkwyQ5HhSKsQ7JImVl8EDMFxJohzsStic6cw
LmisjkBBXjkNad9jZcM38D6OV7OUj9aS+ByvLsgz+J0aLa6QIlfIYsbibq97UqwF
gQlmodZSD89KYAG8wJ6BkfsjY9fum9XGdyV3vLtJnKrWqy44axKw3rxa15M8YRm/
vNAomFjYLVih2nnF9vUDCfDsPdUHDDRO1J4RlDUlvMToF50WDtAQ3DiuIUU3wI3Z
ugjHNXmuoELoEOKAyJX1HMPqTbJu+Y5u0TKp+RE8gQEyZ+eMrCntsxjkx2K9wpCM
MUbPzKEFLoog67S/sX46qCAppndL4k5KNZjE81AA5dcBdrvZs8pzPW/mY8oxZkC5
YXOfrSDn6W+XVdFCmGS8Vn17QbfMIZSBmz2WJS8Rd7GPdoLm5hHhSKpgB2JvIusS
1nVHAVEX3iLO/JoJV8gWEZ3c1G8RRB/bty0wQPlZKabgyJgy9XHdtSngoMTAOwYr
5kyBtwV3XkUpKeqBoDdE9OEEfY8IwM5EmnFNbpSasJ9klxTqCaFUlcgsbqwU8TIZ
HxYgTOwBSR4vptnpjwM+yGqycxOjtM+T7JAzD6eRR2JcteG3Jogdff/4vKyLsCCe
226YwWBgDJEK/CbrK4HpIp1tGnqbbuxQ1QEyJIzLpl19iK9+GVxzj/7GMwH0NMZz
7liIAwu6K85njzbpqRH1gXGsBzSs2UBhsaTzz+s4CFKdOxDrGKamnlZoBjeTMDN0
W51Whn+KVdzJRNx5PHwOT+YjXrWYwl2rEQ8rX1KzUqiJJ+dYemhrpypyX2zAfZKv
85DXk0+eWiN9BbdK5n9whhAMk5uwbW1dy8aYP1n6fDYhl0h16SaS6c2mJ22+mJ+y
r9iWWbDqwVjx0CVnGXoNjcVGIvif6v+IDFV/DCoZpI/HG9b5CgrYWOKz/cKsQZfQ
wRflFoyQimXqjOITbprZmgH/xqiFeloAAJdOrLPIVTc9+vBCRnNvG2lHvijSiwi6
7e+fyHFZnSlBc6DFtFwqaSP5TBBtQO2+K4aOWiB5JdxSMGXTO+yagU0ZmN9CGRq3
QnONCc9T8ThcSHnA8cC1qGChHoHzi0otDjJPLyZU46/O8i1Oe8Ghhz8hgHQzQQMS
NyWV99dsa+K/ZJ4SHA8CilRzyUYbC/kdiMVADNEN+d1rWSwmqSDmfHldkYGkmgBW
k5FdX4afooVEhGvAF/tg4QWkOB+D76RlLeT6PoRIvUS6fw9o9/e+y5tDvNuGddja
xeQxQ7j9OxbJ8NCfU2K0TA==
`protect END_PROTECTED
