`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0+7n9ANBrNaqlT0JBvHLWSFAsBIs5jNi+E/slI1HSfcVRR54BQLoTMAXiHDOCB2
P8upZ2U5JMc98cQqHFQNPTohCDIqpRTxbCFINF1A+MjhPcIbAuuikpfZQvIIsP+R
dt9tSPXCKQ+Rut5B80+9NSoWkuMYGVikLYrJfxo7aA5e8q2xZsYEUo/dLqmVyzYR
L0+ScH3qhJ+h6xtZHH686EDXMfqqaps9CnXyq2y9Ml75ieCg8Wc+wBVITFfnQojL
4oT9/BZONzkO8IWEjOpJtKLEqXptVcuACwqfGohUiXEkraOVXOf3T9ANmDnoZTLP
B1WVrCN0fJGERoGFRxMeTNtFjJ/ZCIW6xa/1hy+eCnTrW+V07N6c4u1yr+Ka6/dz
QBMBMzj2cAEZCsFPPE7kszss8K8IgXYHFGe0Z/c16/UQXVg//vKRmMxJ93H5ekip
rb4EjQPFpQd5QhjFpsMKSwwegUq2nL4RC8j2Zq3WtsZLjvQSE2rHHtW4xp7V6KKj
rEKLwuWDAmA9kqtR+LXfuAbUHLUzHczHGZ9sSwzSBmGdQs2F5g7xD7+Cpid2SGuK
ztGDq7Urzli8bxzpBcIZzDet6l9e7yl9bjoKW6agYbtZaRRsCn8ZkNQMc3ChwfG1
ftobONDzsX9kFD8ALVFh6/kHssLUypbIQfZ5ZmvV6TqbYsh9U+uhs59QQ6r0zKoR
DxCGikCcxFP1UJoUljPEb5yQytaPAE/X7SABQ4llXgR+HbijMFVIOjaKzJYwZ8lt
qduCjxT3TucJK2PTS+EWVALu5Sc0PEqNc2x49KzKmhko+5Iq5wGkSOonm0skp8xc
chn9TdcLcqZhHhcoPfGXyySq3YqRWTwyUeWjTqdtq/x/09KDaHqz9UN1rkobPBMR
ID/FeBHq/+HBn0Fgcw1MZRM6+ugcanxo/9ZMFRgyunQjzYAGBRj4soRn0K5nUa5C
I2TYgmUfCvIZFoUwXWE11yRGv0LCWJGy+uL6m1XKZF2TppYcnhxKo7FsJM1L5GLb
HRzS6+PFffedb0635eCDl9sLpeyn1e0k0lVM/bgWC40mw44rU9ssLzPyVLbvLNkK
ZR0qQmwth+/0FjSgbUGhxAsGTFTJ7Ye8uGJ9fBj6m/h4u3mj3X/65KG7ghcMKyZG
PvFa2qszlz9b8KGAp850dr5HN6py3xNG5fkeJUPZsUV6BWr43JZtCVPVujVKZZVz
sP5qO+5z15iY7rbKyhfrkcsJdV71GaLPQ96Fmmde6MNIDqPrkXw9r5bS3M6bsYyG
cT6jAB0cAGbQQNxeNa2p43ROHUPL0Md4YTGaGujfJaSerCTqiTeP4LJfozYsxBV4
R57yBeoACOtMg2kz0n1fKSufh24tCUCafuAxDqsj5IoqKtzTCRDUC4tkJbFMmxK2
IrvgxL68pxvqu5IgbgC98N8pQtInPzwiWjpCtI2eBn5nTJSBXokM+V/Bjqy5FoHD
3SFXC0ewe9z6Z25dQ/c6oDRTcd4e+5QYBSVQ/0hZjPONZ3yra6rz4Gk0amR6hY6c
UzxtYT4T3ZIUE1v882rOOZYTXdlac8B054gxwG04c1xJ7TK3TsiOCILHS2sdywZB
jArbfeDh9DUa4bxtfFdFELCv+5cC3Y4nIu7IrQ/gIIQq0LDo1Fmkcbqk1ryyymhz
+tUBUlJ9l/8oMS9B+0d1lsf+OuuJmgwug9cXDREXYmgdjPeqoNj9qRQBab9bNilK
Kpdsz7NGJoPNKEScYZMepfvLSBphA+TfQGMp5+sU7BFf1ynweJZjAOoxVPkWjdn6
SE4090FazO2RPVB8grlyMLjl/CK+Sx38JvZ8Mkg8D9q4aeAZ9o6WbWZFRHginSHz
4quF2KLhaFcE9PNLxOhDSLj1SkNhoN2sG7II3wZy6l06YfCrr7X6HWwnruPyTlhz
I0eh7SvKPcO3v7ybuxW2PYPPerjZM5/mNH6zNNgI1YPBzvET9DaIVhyOE9YVmx2B
99dlG9cb2kQG2Z58KuvP3LxXyfwuIdUcZeNgAo+oZk8WRO/xW4ILZA47YTAOtrEq
zbYoBCOaWcjijWorM5ZZsBg/9+4pavgrQuATP1tdwgoirNzx29d9Nr+Gt5rJdI+V
OHNsiHEIbX/VOMOWeSbgzjAWInazqgagtjWuuoktPN/DfJVk5Rju8GCUTQp/WeGK
C/lBcvhGuhyhRvRoSHcM0CaRZwdgnQDhY0AOHMeGuDBdKYubkyDhQwoE8YBzh/jp
kChaXnAq2M7D2OjtaaIItFltZU8vKtpIRC+eYqHP7pf7N4cZr5sEcszeLZMhBiXp
fWRUKdi4UWAebJDAxxrEVjG9h9mzAz9OziOofW7moES25oPdh5ZWbPgAOP08mXgD
sAhBGeC7mdFYczJkHrccrR7laih7GL7D5JpI1ffloPk5sfFyAueVQ/ilNd3iNu6S
tJW3W6yRDvKM/ZZm+8CukXO3nFWEsIPGu0il9yzLVpxfAjltxxOdYkV4yAxQ7kE7
5RCsamY4fYkRcVodhTmGZNzwFeV5SOKqBEUSZLrru4GeQanP7R0rg2wBhYIXV597
sx6W3K/4g9BmokVaoW9/8n+zPqQIYichMMu/Nt/7f79+dvvdhHqEfkETlKuoHkzc
3M+kiQ9jSsXjKd82M0wFs5ITQJWth3OyYg0tKEu0R/zbKGwEY0KonnoNrgCEDq5S
ugljVF+Z0HZBO5LPy/CIcOy8Qx1X6HapzbI4EZu8PFCdor44pQ4huotgjMMEm7va
j/2yGt5uHdlAdDyMhxXE8+mwqlL9zaf4gtx6yEXArho2SI0Zwu0ybJ8K9TMKQDLq
0qXZv1P32GxTLzTaQQ65LrBWA4xYVRIM+R1Qct+q28X0EbcSzBJiaovPPrT7ciNm
odkOpyVXmH5pavGUA8DlwFAwZu9Lx+2VVfANdI8X2sPYQrWki9lcC5kOis/zRQSW
+H5u+CtVa4osOygLXE0Y9TBpoHJ0U3d3cvEMLU9UIZ+w3MmxKzJbxFEEFxE0LU3Y
xtvxKMuEWcvlcF7gdhLEmFZM6IUcWMoQNQvcUOVL7lDVQDBaRwEKd2BKWwSLb0Zc
QgRiJe9dEj8hyg+1yHib+A==
`protect END_PROTECTED
