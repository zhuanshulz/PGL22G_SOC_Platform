`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3/4M3C4zJMzhkdTkKC0jou5tPZ8FpX2D7BZNqFQD7IcOI3XLRTC2onb9bX097As
pR3lO+/lCM/28pHpwGB3sDFf47KlrDvPFmPPWjKcMbxcuusTkbY6/M3GI5xOuYG9
HSOaS+/i6NWIYRdjO38DitSn6sWiXoZPw2lAAHLBewTQeyZ02xkGimQQicujKkvB
ocUuYPPExsFgEU5GGkA4BSOuj33BsuII9lng0GVdaIi5Cw3llfDLsNOnllS4yVtS
2qqs96Wc+CLS9bBbEGjUaDZ+EDZSrdSlGkCPjosVZS9RbwMTdw+UPdlSWgGTNBWQ
u5cJTolLGk7prJTKtjJignqOZVGXr/Ts1LIJvu/22mbKZ6rY8XjaEFPvTchuFnmn
bs+9AqFIffCG8pz4tYLyKx9AJ0xO1R85oCRv1calya8V2OUv1n7hOvnCM6ht0HvG
A+SNXu3YU0hnP4Os0cBq9+hmqg9HvFusNat8hr50l2tdfC6nngXG9saVQkaM0Pq6
dbwRrqhh3X91+3kEIwp4z62iQZcMANryfhFD3JVl+wSBwIwHa8tCrJ8klP1Uc0QV
cZ14mmEoqtMnnPGhH0LV/NNVPhVFjMMX5RJzHXQjBlUqP3MIJJKfqD8NNFxr5OzO
WaBKO/LOdGkDlk96HHPkuuLIHDmZuNnxLmWm4ybWNDBmRxhUzG2rNvFpGhFxKhi+
DoM8oZuocSSvU/Vv++EeUCoIgTNpTFpLhRm0vgXOgvHLfHkd1w752w+45KkSsUJo
dhDwoGdBdJceagUO5OGIHnBQIJPImTH0i5PhCX7n7TnOa5Fno8hN2k6d7ciUSOqy
rp/yGkGur2HymRGnZ2byAhaZ66jmGoU2+2vfXDNwYl9YVmv2fx85h3DVZDfSD7kp
8PSg6R6GDm5T+/LCveeoIU6WjBtx/XM2qcMn6t+IobZNrrLBWHaT3FdJvlsbwZq2
gja7VFGjP0QHbQa6aHsoWIdOCDkTAvVxOh6+rNQ4gks1sDGsD13Adk8m6CoRiNuN
ah3SGgm11z1qVI7gAJ377CbeWvOEcV9kvpQTZMfeZNmsM7Of9U0wQ0NnlAVd27KE
vQnicMz6nq4CMiSfwmM1Gq7MngGX5gKNuDyZiBqcacgsJKmGUg4oNmLpCUhZw/nm
WuaftgonQoCXB4iSU5kpXQzhHCO6lB7yv/PshMKUKC1179d51qvxEO4R2X2WhTSW
1PPAhz9CcwhBzfI7L9MPO+j6o2rctRuHea67fFjy1XpM2PjUREL3G14oLyaYslAl
jzLCfUkTLw+Utzs7ovZcUyyUSbWPQr8E8A2gNwza9rpUpERoeqIMX+/zZihqDSQb
B1JZx4fMSSj1B68KlRfoWfTtxf/T6z2IJo7xG/4aqZsbCjB5lwuNUfvRjPeb+LXN
b9NZy6DCYc+YKdm/ey8kSHzbWiwcyx5pszkSAnnD2jjcGE5q4pf5GYsUJ2II4SR+
P4XwinRW5JNSKYwqBYwlOueyqIQUUa2rAdbIJ9EqUjbqa7+s+Xax6nScPOj6Q7+V
/1iIj9Yrg7xDjnTMSEGS9/vgnXhxjOqF4fs3RkuARjYvhLTObn0mC99EOwdfjF7o
UFzQMazwz7iQodLqGMQbdd9Q+e4bTic9t7wCc6BKKYEijghNlDlZ/obl8k0bP5QZ
6UOzAQ2G7l8kfgmjhmWQgzhJIcyNBlx1WpZv/TBqS/Ej1lY6DaBdIUsRU4GplC0p
PK/zgJZIqhZsUb07+XcAs4wQyXP1HTxG1V2iF8aKB+w1DFckpZyam7+AwttWZIRw
HI8VcNuP+vtMSHC+0IsE+Vn+MY5jXl9QAzxWp0aGUFDy1568ndS36VNpXzy+oebT
37rRGTTUf+nsZWwsUAW68HV/KLe3XoSWHQRzd7BNIUUbuuMbwjMsR68A4xjdzP3i
ie1sWvNKVSIa9gDWkiTrOrwa4wbsib90PiN/AgHNZYaxEGMfPmxlPAyfL8vT605W
ivSRdjXIw+0Ww0ajl2o7tz4pmLcVKEqrFx40ym/0Tt/c8R0iTsHidOZPCUZwx1bt
9WqErVxEPhkB4Yimf0h2nL8Yo3sUkUPvcU7yIte1jGEbieh6qBcJStxvdjZDFqGA
64HP3JTl/BNCbxULgcGEq/w77Qv97NG/CkuOygyPEFDTSKzX++CiXFE8gSWMlIOr
Y4ydXuqiCAiTgO0rTwtk5EW+AJUY7/tRDLBLn+KfyICOVxqMBwIk4uKyEUw3/Yxm
yN6ygfJ5gbwzI+5DgvMqhNsYmG9w0YmhHAtcaeNALta7dMsFo+zwIOmie2GFg04+
P2ghLLxlohSTIs4+I2ecGg==
`protect END_PROTECTED
