`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dpMFoIMH2qfUaTr6+bUgMuLy8x3Xlp/ZhsUKxahClqCwfDWUbZPjfXOh4eRsCxOK
tOACPPmv9jEWvfONAJp3+WVKF0dcfDhZ87cBudI6iLxSN78TkzIw+sXVKEziaRDZ
A40ySWAtXrNgrQqvPVoOtkZSSifKM4ELKcX+pq3GNqMdf50to4pg8WtA6QPsKBKN
QxBVXOjh7H0r1P4TUBFNOJ8O48iPysHE8Q66GziqgfivSA62rU38omrWcF+ksLPA
d8uoUxqMCJeRaY7+5FIu/zJGSoIBd0ik6niQal0DEaraPuoBxYLpyn2/bozdrt+M
RdYeo36j9jHD6QHwGoYHkQ==
`protect END_PROTECTED
