`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rN5ZWvS0+iekCxQ2kOlOT13WD45nG7sNYHirUbKiGiydKeAK4D/hCAnPJAFVcz4G
nWLlGJ5PSNSEtI8vOurvTXFjUnQs0zGuTAOnGBmCy/jeaaYqVzLC/hFQ9zYoz3r8
Gk7gv8YPBBG6j1m1etEPHw4CrQH6W6AupXEIND/D2ZezmWMcAPlry17POsRhHDmi
w/7yHy7wOJV/lBoglIQjyOPu3Syk+sREyHnQTMzY6I1vBc+wr9wldwAvF1qjqEYr
g2E366xVQf4uhXp7hvAG6r1tPWAjfJUXWbZ0BmnT6K7vnMkPt/5ouehECgmhvpWS
qT2m+vtRtensqnLFrmGTEH/f+ytmgWR9KK3BI8dmnDXlrbhhODJu1tPUSdEpXqMV
a64jUAol++PbqXBLk17oT4UCp2SsVUu/QNipWQq9jw3kFNHkxRpLolX7TXs9mEO/
5lsSXzhtizUs6lp6ycEbaOIUHIuhp3Xso1yX4c0i/os9nwNJvGLSefxemupUawgU
Ys2I0otOn7lsPBUJzdM/jj4t1uEndkqcOT0tFStBXQ8cru45qK4Wb2XKAL2G6qsY
UEtEwPZxWQAn4h+cGz691YSqSSx0+0LkLZB672Wmzzu8IUVAx5lLRGYuhtU9XMOk
mOQeKVX6jFBHGGA7K/LITy2gf8xye+Vig5qphPNUy1kSSVDVnDvrUF015Ly/rpZ3
vZoFijp9mL5Jzb6UwLuQSnbPGiK8FRKCa246XQF/x5U+q5pz0KeUPdwUd6PodERe
FwOv1cggluNPNfYMbr5bIBIwCfcECkkYq9qoZiEVuVw7uV76TFALndz//+YT1mn0
Nopsu++cPCeOG8/uiLKAee9eydDuIKt1R90DZAnhv1431+pAzetSfkRsTAMOExtb
L8QLrsnizjHqdCt71UNYw+DS5RBXKwELh/bBoG7hjea2oxvGrEviKJ+F/iYTD12i
i2/gQaE4N5MFC4GEcMPhzfbBdK4Eu/Fvdp46NL65NLL0IUF399GCLwQ8MPB6rGlb
H7knYJdeMqhBqasySVDyUflw2r+PGggd5IajiQ74/WyAXlmIKJU/+qomx+E9tPQ2
Z5v0tk+lTEDh0adRsfyr90STKzwdtoeP/TixU7gwkr/SwxF8dGcwb+wlRk1w2qcv
j+7kPdYfC+sjOqNflN7Pviwzt7IgElLb3HJ+cni7olLbV5OONCyuNCD9EdS4X+Wn
q3v7MCs6Y1ElOTCOHW3MG8c9lcSxmEAu4L8NwLqGtQamA6MwwGFSKRg0ovtCng9j
HtdG7tYH5qUyvU2R0sbInjoq6NSIYWa8IQsX/vmJadE50aj1/itaJDzmA7Hn2UVW
rWRLtg9zBrIJdO2DifjnvT2jVi2P/JPpcTtrptKhGuN2PdIvvTtLOzn8wHbIfqBD
MSwXQVPBft5zBv7eiwfTpdLFLoaWJ14+7GL2Vpm/sfLAlzscAuEfn+8njMKSQVaW
TplA67Dpofgr2oA0YBgxqE9MBLHLVpaEi9eoSbZVl6Sz0HC/csiB5Y5x36tvvmTS
MyICogG2MT/JkvJSc3XXkmmFXY3v0u6V9m8NwQkgjo90cocYWlF3HJEYSZPOWEMs
MB/ZVqUxZGlz40OZuuSBJBd8E/xvmKgNPaYOQnSkC6z2YEXdrCDV/hbQFdWqXfCU
FY0qsHMRG0gS1bx7UDYDyx9CKfj8O4ku94zKfDUdoD4hvsVbRBGGkI/vD3Sknhhn
Z1I/MCuvEhXbLU6F1W3fQtEnvrhIeMeNH8ZNv6dGE8lrD/wCTHC5owil0sTm/Kv8
VjF0c7VYJDm6bdKYmjxg0dPMszcu/w+uHlrlQT38Fju7/iolml/3gUDDKf7Nk/cR
`protect END_PROTECTED
