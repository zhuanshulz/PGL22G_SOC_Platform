`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BdJr2UDG06VKXYHUrJ7kWORhD6EL0JBMeyn0i6YNff3HM9AeU2FJt8vEvmIWFrtj
5tBYqavZLTALFlGnfPaRzoyfTV5gg85ZA+hvUxT7IhBt3ukOHLuyb3RObTF7MG3x
m41cZTd4ouXhI67x8SshWF9zHDu0d57gFw0uaRpjO3JHMxbG7Uqykwi4/T02tpem
EVj2ecWUWLQ0ZvR5/52/45TLW1TG1N9re/5LWFW8cHM9OXI7YY+Gr+aknffHaNGz
pZig7CNjmz3QUzZLbeDeyxodIsImEl/C93y+EiIfamADRLKQGSE5lWCM8jZbU/oX
Aq/939khvKbR8G+AeviVI7PLTCKoUwPO2X5X3u8Hkt9S9RTkgHwFR379/wSb+J6j
4JO+j4hnb8IrRJ4YvMhC24bruc4GUvTZ/Hwnm9bKRSceVItQ7pl4VMM3jiYqYy7J
jxUOllXmoUTQNFBu7pAytahgRIiqta46CwmF8Uibf/w=
`protect END_PROTECTED
