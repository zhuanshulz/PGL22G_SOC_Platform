`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h0gWh0fwLzaRGVxF/ocmP5l4hJRU1syv/s3RUwKUeozKIkw8H5SZ5SXCWpNE6wcV
UMxy/lWjyeF7RM+VVI9xcntCMs7jOXu+6HxDGQQt+vVVAhDSM4t49G9SH/ucEffL
L1aGYzXl0w2ITpYS1O0kFpfe77SpTcYlkJeeBQ5WlOyeJEm7/YeoGm3xUhCzkvyY
mEcsWj5TalvV6TKYY7fzlMVz6zHrp7wft8BOoXmOqzlrAOxGLHKv6Hh3DpfqGg43
8Qct2urpzzktVLR7l3e1h7G/vRuPd0hx/w+kj0rIbnFxCYBgkTuhdqVbOH2u8L1w
i4483XKBfDzRfOnQeQ0u81G5lvg3sr7wXD2omwG2uDaGaFPa0bjKQ4VqcFzwAZRM
X8nGPW+OudvNd4hUNanCuAUgVtCP7Bf8MIGO71Hn019aym21g/7MLl1j1JcHLcWF
LIxXjRbw1SWGqUvntqpeeAKrA3KgUPQycRIGnNo47/WtNRpzNuB3Tk/BJQ46s8Mf
MxqfBU3Zv8i6LVixyyGz3ANcLrFDl3toQqQCgNPRpeodQ9wq2JFjIumygAQnxSLW
szHgJ0WC2v04EQuU+bQ7SAGkh5vYPm+TlxzbJZqfcMJTgDnvgjrcm7pPEeSjrtYb
ZZoNfZa7krGX9R9lAXR2i/LBmuJ+GwmykenQoP1oXp1/LgL3Zz7y0T36hMbOvaGZ
PosgQaAmHJAtljk+YY7SO1NutABq/UKAS9TIz0gizSNR4fc8DiIatQBzayGJo2ry
EIEk7GPsdULCj8oeSD44P/8NG7Zj+gnvTjihwtuwITcRqsSr1tiHZNKW/Bz28ZVX
`protect END_PROTECTED
