`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7SL+36dSererIlrI31z84LByyJ5kqj3BnS9TfzBPj1oaLyxjwHJQ06ImahFe6/4L
aDmK0gtgCG7ol3Z6VDWvfNEYGGXsZ+QB8nVt2SwmVg0rRILCXTZd0gIZubFHmBHN
TjZq403bb1IhNcmzX+LvcDfNZiKrJtrpGmmb+FzllnNeF1cW9oaR8m5hFTE6jvbz
KhhmD9BHvdmBg/0jh2ZsXaSXdiAwclEal4AhRlj0iGF0tgBXlbJcXdwNJJ/jI5QS
tEcecXyfZHSOab+UufPqX9eu4NAdED9+jf3nOK0dIoagt92gktNvDOIBpmt7gU9a
uD/rCuRtRRBh3GPmv+CxFeV/FmnmSX6Ssm0Eey740fvp8FHkfU+7Vingt8/3T0Kw
OSZIzPDgI2U1JFXmZzm6nBYhFS4bnIOmmArRhczwLqD7k1tMwBdC33AThEcYIKlB
WlnRoklqbsVDyUBzQNflS+z8LySRGVyizmqMILG4D0CVUWrzYog6DI+VRMFZsPXm
NJvnMA/E1jFFD5kk5OM4o69W+6cuA4nWDmOMSWbEADU6QE0+WPQ5Q+Uchzrr1d0O
H8YRqqYhPF43seBiWHEgKSRTcl3GTtSxsHHEnZWHOJnupp1428kigNK60fq0DVqX
wsMtFh4oxgoaZoppd4oWwrxBDNtaehW5ZdeqtjRf6rMkorfPzQnh0IULdxvnnyAs
H4/XtgD6MrOhXm5J8U9ySvuMW+rZvesqVTPXpI3xMA/8IqyXklSrEzOpwMLJf3+j
JllWba3yspfOVc+xmGlMHuRp31fi7Qm5vUtGmZM+s3P7iPQP8rFIu2KJGZEmCfnm
w1a2GrzAbnVP+XDrokjDCakzlpzQDi1EoqViAbiYpTW6siC5mvHTs9+pCV2G8Nd3
V+6+M78utRCsqrnHI5qQqeTmBgDR7wY5rTuw7jzGaRfrGzMwZYYu8GKWy3FBPe+B
jBpqGAKfK+BuKtvezx3OrLzz1tONjfPCUPf6NSOe/B/VaaLWJ5idmGL+owq5BQSH
Qnyea4cyGq6I0EZ1fMKR/U+V3q5mco1cRVXB45K7+/M9QNnCcBGiOCL1DstZTRGt
TkmS02jM/86fV8QH8C0TCR54AIlrY9RZDQYh62XGzYQkkzhpgJuMJhf2Mp4ItAnN
Lw7v26szZv9eurTLWgD1FLtyhJW1o/2NNgbuh4vFr7p7JFPxSfb1YeKDSFz+LcaP
dBOdklFcZpSjbWl46UaL3JQFPmCgyXJiRE92RJS2nOFt7D0Ps/JIySUrdxbKSPsa
esVpTkOgom6FA6VvdaYVXu3upG6plysmBqBxdFnfYowCEW+PJRbVtbGEiLK96l5H
2T/TMTtzyihFJVZ3K2Pjslo4oj4iClx3YZLa7qZOqmxHgNz3RNMbrKyAvHkvdyay
8Bkb9p3jXic3/qXSA9T16iaIWLECJqw7k5xGQntAliPW3CjDNNKG6Hx7kuDM3HGT
sYOPYH6HxHMuDC+u6Yown8movTUKtAxAtcWInp9/HZ754JDXSKCvfBSfKNDksc+4
mDQCSinrE0Di4b5bdvMTXpp5vOZlI/t5olNRlamru8kfOVQh/O5FVRyxc28asKb3
pYUJ6tyAaUaIQkvlcKzfWW3woMzoyGPVe55Cs1oWQPtlhnx57FzPrCj6mkcg6ESr
EInh7sU2juB7xe6cIAlKZsK4gBL87QRQoUfjSTPU8io+uT1gbf/fAKxZxVtbUIJ3
UEKjnCXM6IPO3ip1RtyrffTjnvlHw0dpxjNq3DiYoLQcQchrpzttIe7nuBxYByl6
7Su54H78YVAZa+qqqtL9RbB+atvyedfQZt+EhEBPfkz93BzN0gjmHClwXIH2eELA
mnQ/wsYY54p36VHwHM3IyNVxNjAPF0GTvHvxzUnOMIfThCM03bPsFDTh9742ssVr
u7OpXQJFwX+vrVVN1gqrKIyc7b3h/8vLSeibtCT1vQwrjYYaMxRqwRKsWSjtk9/B
QcWF4731sTj8ZyZY3OMhquojEOxwYRyblDi5YGPaxYn103HMxc+YjidrxV/PyI3Z
DTWvCrJ9qGEZWlQjEs2Kh3ZBVNsejkESIDI8c8sQVXUQFpU1PdLpMLviKLrc3AEi
if5KNA/tuKqN6lf2LsualJn7b4bMdidOezooeWto3par2ySHFzWwcqtD/cf+AdMj
AamWWHCeFKNac8TQIKj22iI72Si1S4UqwA6voB0/E1szArgFH2BtJEHl80b67gv+
UIxs0tvnkboWfr/lWltYHgKiToFYcRyLC5UJss9XQcBJTJvHI2UDNI2xJATFbPFW
M6qH191WyquiWe6dvSaJz3ioyktioeujIFWxqDHIxopGQppDSaZm9a5x7G7gcDH5
JE8EYRBpWq1CRmn+MpleHXrEJ4LIJrqOGcLCw7U/k+uzf+eBSdhoH12/SPYHog/G
uHv8pexu8z20YaPk/+wQveomWDqDR9txMzZNDDmuBAwTnnp5DuCk3hdCP/VY+xON
cEGNbP0/O0VWelTYAZA0MKrn58cni1+Mvkv5X0JX62dEuM8OosM/zQyLJhQ+0El0
cH1d61LokKTW+pYH9Arh6OFo84Q7gj6xn3iIxxoDG89h7ne8g2s6Z3e8tSARww41
MM58OuQZTjs2e+1y4gbLzyJPe6vYhlC7Qj0ykt8c9b4XWf5ZYd34JoZPLkJ6eOav
QO6umd28HXnTAuEsOluaiFXTzYI/3im4HGtTOtlvQkcsVmTqLkv9L4y57pO2eqaS
VW/K04PQGDtePvpMzFtl+CnGAG447v4nNBvYH3MSnQYo0mD1djsmvza3/sRvXpA7
ZH8VeZWldYDubNEb9tCeqvHG6V2eP4Mf33uPsCWG/AOvzLHTFe0teatf9UzSFqkJ
x/RJi4jYI8KnTOoEL81RKBxesymP70XotXSgiLZHlxEKwMAQ9yv+eaIsXDvYG+Ov
VsSyudiln5yATP6DCgI5g4xbtkTzJryEsAazz6XPx4GdRx907SZj1QWhKGtlj5/Y
X51Ek8Bln8F+DdsMZnHL0lQjVBdXpbfrY0OaiXYsBnJqF1b53cAtwN0VbCTyScsy
bsRzNhN+o85OCJ1Zf66qjw==
`protect END_PROTECTED
