`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TyH8vhEyb4ea9d1IWl08fFuJv+11UmJZmfrPxIjQiJ/E+etPUPTxSdoMFzw3PivR
qVKsTJlfJ3w+8egASpBpVHOdeDPsE0o9tOo/HF8EgMqI3DBjFAdG+e7iXftO9I3N
V0Sv8gsVqG93YWI+USKmPEpE+BsK8m7CrZSkqmMZXEnAeV000Wlow6SqCKGpAG9G
54ZeXuyIlNU3TcZ4NMTvPnB0yJQULJzmlrESxw1c6+ywlfQRIdqXWExqdMLP86mG
hp7ma+Yf+CinU4nXKlU+T6E8BfeqVlbn9R0QwK1Y4E5e47pwmvJkcIBfAdN8KHPO
Hh4Rcbx7+lG04/aRKkmgsFwuRfD5Nzn3960tx6pBVm7/16Tcez+Iz46Tqc2iBBUz
8tz/hZQgQ+WAKKZlJm40v6nURDBDYCVmHighbLmr8H4Mye9jQdCANK/f2mdWrOHz
RAej/QlHCU+A1+LzFZrEj4+GzuXt8LBLOGFQb3n/xpsvK0gCOQV1koMznslvYlx2
1SF4A71lAGfPW/LFbzvRE6zgxRxhStKU+MocQVOLGScoEhYQ20PEC/zy1nolaQNH
hf2W9grIr/kugOi+KCMqPGHCLux8u8IR68AXBndlsJEruOmdErNH5iKp0nZBpWBc
PhzH3mIyV6xNVKCyHqLOdJhZXOGccl1xV749+BScjlUibXTDZS9ConrHhk1CyNTu
OnzGnZm4cXnteXCpC328Zbn6yNu9vLFKo14W2pRLWzn4or09fbwH6ZuvKpiEyVsL
S3/PDHKITUo3UkofrSZtD6V9BvVKHmCrCBiVXt7Rm0khqfEsOMes9Exp6b2rrWpu
rvVQ0zJrlm7lb73ZkpC1BOrdsW6m82ps/7FkE9zZl4vDmm++tcJwTT5NxOWj59T/
svHNk5jveBGoUrNXypDcPjh+iYIo0meF7/RLf4Uf/TPbvKOyMLlfmijhPd1nUTG4
1P7vHgZodVubAeyLXAe2wTi9qM6tvdHGrrnQvqFA3QwXBLUiDx2gE9JYctFgrnz1
RTW3qNqMGUVDuay99RIqk4UNcwOvH6AedhAcJK8C41iHsyYtGaP8BKD/slPIDnVB
BtaN/qt8pN6Y07f/RIAlns9WlRJyFVXbeMzB+Qm4zUvCdeZARyEfYEls+PwAf6SG
sOwv4m3w8f5cVbHkAxZBL353qWR9EAbf5f2MNcBvDQXsyOT+isoeN2LU2p6b0Ddu
3SaZ76wsAFR++THwrc/nfyF6pn0dd1bLBcBh/i46U9LquSE+QqYJ6EOFk4qzvqny
0ZEMoVLTHO8NSaXhUmkW/SvBaJRqBDcwWBUE0P97Q67WkuVeQkI20JRhDVIK9K+J
B0W/P0s11unlyoovI+lTz0OX4kMeZ81DahSB7c5oj/6FZl7IxeHw0xIca5/q8GI9
uUKPNZvcrobdqhUX4AopFFOSVHk5n5UywC7FrgMuwl8B43aQinZrhLcwSl2IBd0I
SfJxM4IZghMpU53Zt8NMQtRNuUzNsQq5wYSeTiuS7iP4C8Tkrwzmy+8uB+ygR0bK
VR/on97DhOpY7KCkeCr5n6397jWlMgUXNlt2Umn/c1bqRHyVxdycECTonuEe4thj
E4SzOdHpk3Zj1ZDY0UVxgkfoxfb5x73pFvUmnUlqcFs3X+qlyAhUedFBMpLXNuKt
zW1PXc8zNi5zvh4m6Mj0M0lEpF7PK0M8XN5PqXEGl1Y=
`protect END_PROTECTED
