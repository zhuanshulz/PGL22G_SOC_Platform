`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iTez0m2hvWbv+I/Dtu/xHMsVS9bX5M+M0Wu0I1Qtp3e2ZPB2Idj0ehwXtiQOY8gY
PkS3nA+CI3uwThFkzAvJK2NUPfwX6xX7k+bgvkTBDQsAcPfYNOEsnHOdlFAcEOl4
kFGohzx7rIGcLccxWSAKl3I5quyOwn1DtnRKrkN05cOrpzr4XxVKc0WbrAcRMY81
7wqd6k28Tim+r+U3Dgj4fu2Q4/Fv62aDF/1E/Mv2jQ6SuT3kvdvhKq/vjepJ5Za9
mNQd+7HeYcvbsq8W14wQmNMG9jbBii61kXPBopHpoeqArufJdeQw1g2cPwTRVJZs
uihxD2wBrHQ5nmbDW0MBuqzp3UjOTIxnQDN/8GMFWtVFgNN1fr0+nl+6wmm9ulde
AqJUj8kydIZRT8EJy1c865Coy9iUO4a8FlZGzXaez4m9kG4f/GFTqBZ6X2GAxQbh
sbaKFov5Ndop9xugrmJeuHtUHfaGlgiLA93P9GhTOF+jgLFq99MKfUDfIO9doZaP
7I8BaLGZAHgAGvWHY0zx5xmLuiPXCL77+Q1ziEewxsYTlRSYr98ZZoJ5LpvDHtTQ
PGEkZayegffzHIYo0Yz/UFCBND29UaF1+LRWQq+PLNP3Ez5acBvJRq8r6/NetiEC
eov0U7RUfg2LCOmv0GDOdeG0fQ6M5SFkQ2HrEHr/7dhGRtU1rqBhsajxNQ7dzPcW
1soomG2YZCxLQiBiAOUhCko3EeHu7Z1/2AvJ2c/HCx2DH41bEdVmgCs7h0B71FTu
E+MZpLFg7djGftReIya1+Wh2yAExTFRpCmD0v2t39KlLIt3eWZ8hQSy0UjKKyIU4
LDLoDHa9HbCzyiPSic+sBHeGkR01F5ywa7zdLpAJTAYfbiTDSTTAF/vm9WwAzFFm
skrUIXjMO2xpHi/FD6sWTTZfJaZ6pe3kkKbESdkpCietnfmaaBuJigiRF2dLDnjL
5DRI240vdQvI5do4LouVrLjIHTsHr4S5k89wLJJHwjOFH6VK7JbQnp3ivnL/Pta4
zUWk5zDxi4Qmjq/LPID1iYYkBkWVs4t577+lps7DiUPihm/zQ9rfIfq7a+uPi6Mj
ebl4iuac1LpyBj87goxXVXJ4HPZ19s1R7G+zUBFRKLn0rGQY4aiHNRrh+6yITD80
kzlNW7fDlNCwZVgByP5UYTVFodCvwWpQQ1HeBQyqgJIIOIN8X9ymUw7YnHJ4Oefu
Ms4994eYYaPdd1CMGkA34sM66NAmVaNws85QJjJI6APyhHRcOlAFzE7P3aOaO1Sk
UWBAIiWmpJfU04eK5XFD/Ow9K2O8RSdFkDmA1q0sVSUW3UGvqBb6lftidgdR9Bkt
+eCiHMxCCxvxxSZawvILVtR8VYse4TDJzw1gcy4A6OdLwhg+KbQvt8I5/UukQiMf
fJEFPCRk/Q6coMr615jSB2zDlUR5bbMjrykrzIw8ThcpXyYXl4zf+Tlg0P4Qt7jP
daHj0bav5pSzG6/YtdcP34GBi6LBFDoMFVLoATWYVi+KM3ZHsLOSHQzOLyLu6Dn3
QhmnvyUWFmSg9tLXrLWrKIg0GqCGCeLtf44lWCRHbk1We7wKzueJJv7hmkkQP3lA
Q4JiYTEGCyzvcgXyC7Lm0y2IqNNjGc0pHpmk9xYbDCeKkZxGhv8bR8CBEOy6C4rR
ibtKrrArgwjjujYazyaLouKIsFTYcqOeQEp6CeS82gTEMbkn1s8zOpd7eDZjLMtP
aV7R4+VRobHLlf5bIKCGQ+GKi9pIeodxBncrMcwr3dy99TajGxe0jJCXIoRClFJ8
wxCD4nC5Pa8nUjXV1ufxV7bT6syhHo1L6SWsMcNULUo0KKfEXrpeNW8n8/5ZEg0T
ik2sHJKUiMU+NZ3Twnu+n2WpxIjYpgEcTVSJ9HpYrAW5FYv82ap7IBz/nAy0LxX4
Ppt35+fjUVtAWXfvbqECtGuYnAZ7DtgeAj+Jc2Dl1yRb8uFo/eUXqagZMJU0bQK8
Z1Huipgt4Z8RzWKE0PaRCo6+G8RcumezlV9Qab1dA/FPO0YTiy+TZkL4s7TWh+Lk
sBG7pHGFysI95oC1l5ZIuejSYzsZ1Qc/006guLap3Km3p3zkK+5NdBm5h9wIGfgb
7APjtaKHVwCppEEiCNe8zJxbvJg9a/WsSH6wv7KCojxkQUqSIOHOb3OGADa6quWY
4y3aDN69mXMg8qFSc4nE9SiLLcs2y3ywmqgdBjbDrBGQqcfH9QM0rm9IDzga8hbE
AicaM/pcXb8tNRklYmH4s3Pk2gMN018Q2C33A1RactThfNHZnhwMfrptE6TxWOkM
siOt88nzlLAYw72xezSqV3Mrski0RCOw3yXsr0lX3c5zVR3vCUz/7klE2PUIsxgX
0gu5rHZ9MTbc6YdrW8Dc9GsMaVYkuNmI6XGYkPrUBHz0sSz1VSm0QjFFv93tCqv3
TraBTPMpluZfxFY01lRtGK3ZUMHyFt+8Fls+4+s/ekOq9FCIEKEaefb6DnUrzSnD
zvLjLjCC2lQ1i6QfYkAHi8coAKooGpbiTQDZ/XJwlK61mv0ADR+W9/PI4bFYSNdw
pA4NrMtMDxOPIyML8P1SsNjOTsMnCCF6pK67MjoppwoQ8/wlxCc1XSPeBhllQ2ce
3UbirMlBzmq3oyMN7+DyytVGmrclFG6R2AHsDljVdxrXE7BJbfXGqtUZ72nz/UYO
f00L5QhR6ltvN9YdI6dYs2rnpL45VmX+Oj2OJBZAmzxEc1IPuP1E4+thI5by19gk
/Z4RQToW65X7JIiE1VFKhNTt7qThNJeJshDWm/qIeA5Zt6Yahr6qIlpwYCMGxJKx
hclfxirXoNlFuoU8B1sANsENQFrQQrm1kgZgkBzwmbygKNet/2rDB8rptPIs/3gq
L5lEjy6n+XSxhv81a0zBfsNgGeTN7MtI28XChXvDix8ZQyjxbJda7yHm2ZPpcxZm
f2SvyRz013ChXS2T/Twha0r692Rfo6LR5uhtUns8HnfWC3KTTtw4ABQleku8hvOC
ViELVaNKE0HI/XyRk6YzaMFFpS5zJBTWyRM8TOyWLOqP6mcvhRM23yMI7C2S8go6
YgquENepyp6Cfi1vnZt9lJSMFD0g05MSlsxnJrEMbIYUcrrItKkBv6kv3etkZfMj
Q3Pf7FbRamluW91QyfoJXceC6OSxxG1y+iSxe1AU9bgKHh2HzkcZ9oo/GgVnOFrb
H31XAHca5lLlitnRGuMCCib5ZO/bGYh9kYjAbb5ofhw+KQdLLGsrGdBQ+1yOxQAw
bJno8L+/3rLVTUaN0apSX3AVlT8fCSZrJoR3t0IbCXG6T8xoR/5k0Qys8ObStkn5
uLZ1zWf9eH8oNRKWpRSF6kisw5QwTRNytjP03gG51Cm7NItaTcVOBlXc/1UjZ5pi
Z1oZyRbs8dXg6JNSqdx+YkNDTQK7wL598gnJRCIZS53W37LjhW7UZs4TshNA5iFR
thVxw/Hwqbj5RO8FWGd6W2JChYzo+dWE4vRDwe3PrVo3s8ZvxBX2ZVR9RI6d5EqU
aasre5LvBFvJFydNHnpya4k4bcIHYRHREmAl9zPL+OxH8o4o1jh6YXDLpcI0lROV
CYxwhOJizcRq0tXzQIFutEZ8k+K1MBduIM7Rqlf/C8JKtr+iqUNs/v5eznNYO8DS
maHG++fIZay8qYvx1JraEH0HzPowsv5RcBRZXokgsdPv5X6sxMZdFFXq3JnP56ra
t2+m7oJxn24MgUC5xxTOTxMQyyHrnwNRbI5PN0fjSAtfSpA6hqV9nwbdKhiWyziF
sCc+8F3gOuUjKIh0/pzb3letqOk7NDM8I9Sy31sA9ghaUWdvXY+wPxpLh3ACOTxZ
MkOtO8Lscb7LjOp/cCGKroR709WSruFPkqxvuEvfJkFNGOzniH49QpBEWoio+njg
wS41hhPJ9vYT9egKKBrvvfKkg/GdpWviL+cPGiZ5pibpzqcztSAQzXfbokk4BETr
RyN2+BLSIjCMEkqGdFpJq0RUtw8icUHzdAQStaJ8tWm7E2hhqJMAwQ82EmFw6zOe
tHqv5xW4IdR3qaQYbN9Rqi+BqXr8yaMVnj0kBb+jQTJwx27A4lLJpHWBjYiEO0bB
EOPTX+ahO6EkgmT2QBSSlAk/EGdYXMaTFcBSU9l0G8oUSYGkxPl6HX2m1qkbcZy5
+8nA+osaNXVPu3ufpgDe716xINQ1tn+tifdeaRX3qjI+3ECFduVpVhwxAiHGh0Ul
3XXx4nHDuMheYxgazBnTk84YYQNcitTAm0k+FBPcWyeE8ehx7d9iJXHwmoAlhd71
aTfmk8YxW/ZdR484yY5z6FVN8xoKmew7irNE3nCW8o38V9CVZ2whkkMXuGqv/AB0
HtgaPE3LGJrzDSwWh/4arDB8ixcjNSxpZQYTqkatcXwohuGMX2b0yRa38Fj9RxCS
TiFZC1DGNzkXlGoamKdiPytGg8I370HcONhM8eqX2E3fNCyK6KUKeO8htTrrRURb
30FZ533KvEbjO00zavvF194VeHPeSzK9FEIcB3bCw3UR1SbVu2K9XJaDCJmTNjQK
pnOy0vgyClkTRTkKoaDUXGapgmvC5AuE497zJD7hVfTeOHyaahvt1WVBjnK6Y/MM
N1ASyYPguWC4ReWevJALLi5tKnsPcjRhkMIqmJI3BRXb7kTW0Xb27QGTfOHZcP0U
naxbAGaY5noDxiCiBpFU5vTXbUXRGPWRl0OMGJrZ42G0t2OVnskeDjCnCVXJKQ6M
+sw2B6++wJY5LcmYm2dtzQdwP2SqUX5bWeNba2G8bedAPMkjmcbPZKa5s5oBE9PA
tr2q8clZ6e+YoVCe96DbkmryfTJTm9AsfsWfWJrhdWY45GFsP88PqQcAPvOCcZVq
TgCIEQauT3n3lKiHsrA4Yb/gBXL3pPAW0NBDp0Dm8mpOG2QJMsB8zP9evFeHq03a
f6UxrfPoxfsBC9xPZTz2tbHrwIZFH7SwU/PUcbQ4isxlJvyadH4/ZQHMXL0SPwqc
H2LRcIjF/bM5hAhURiY8PxSifbHsMj6oavSSaGAlm4oMPhDQt9wu7FPnj8AuYodS
SvSBM7ntQxycmpF/o1+9Hwv638NGHeQx/M/cvqiTwQpZB58T9CQPdEvBKR9Lm5Gy
APH4wjY3ctWmPFTP0Etr0NGkILs3xD9a8FJqG7JHPoUCl2FNh/muum5LbL2DsOWe
NamFhCxHU7+pKFW6tiNvlQIUKrCRuLAovh3Jo8AHG8Q6ku11ZzyOvQQ8SLtsZ5ou
dhp/AZG3Fm/q4cm/3+KNaN6IaINQAkGhHAR8bHYDBCKysqDeJLmP15TZtHeBkLZZ
Vm9g5gJRzNVzGV7d7pAv3LcE1d7RY0vGWFIHUj/T63dOxIJDzYrhj5W+juHzp/pf
vqj7p1OMAfnsziZgfzrm7wTsc5zH50ZnjIVtqT68yYtgqLpARVmugiC0yWJAyNxd
qW/vFgd82LV3Cb48dhlBsA==
`protect END_PROTECTED
