`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
79JAZFAGh5qdWsRmvzbzW4S2UL2hZX5ZVNpLr87XT1Z+8DXCROhNMFzf+T48S3Nc
TTKRPJq4wCjXRwOVg8s75VzCPLAVfzAvrq8//GTY/nzrHk2mjRok6e+TPgYsElrW
y6RjSoSwCdvWojnR1YOHuEe7fk7oW27vErzFYOkW8S5MrGZ4W2Z4Vndma0SrieNV
ZDOheNTjX9IN8zEisBh5gRus5CQYzEIalddYHEnwrSZogC3wvwBabXPsDWteJR//
zQ2xkCHGY8D8B295eP480d02evdW+5JKyDRV+zzelbqAhjA3VrLMbMIsFkuNraG2
/TpBEYcUEKYgzfJ/28iu01u6HojTyjVw29JHBxcjYYkxZqO22O8bFXu00v2AdJWl
IjL7fm1MVc3wjs6EjJ+kUrI/aHskdNDtDYlzrKWgAPMxPCahmBxuRZOKRdAbHxoz
TCN4CJ/LR4rzcQnHOmIBFif5HAYQ/GVTXoX5CXKGmvyO7rMEQXFRKJKHjbSZ+2uS
MYv7X1gF4aF4pohBhSTKPetHX8cAinW6L1TFX0vQLDu1WDd+x9Bnt4LK8YB0qm7o
tUcbPxhFqK7qyCBFP5G9CyQnuWamBkO2MXfwirSsF5dRXDdwVUEdsH4zcDXYrGNv
NkMcoi43HA2HdHujW49uQqmWABpOYlXJaofHlyNUJgaWW6aMUf1KlCrcLdiB/tuA
BvMwhNQ6xynNiMi6C7rYxpeHeLuEAAVo14zMkSE1XjGPnYnFeM5sIXGr9pjovoNb
s101mBI8/Ixp/Qss9ynENw==
`protect END_PROTECTED
