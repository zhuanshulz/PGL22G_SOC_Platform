`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNrfoJriIW3l1TA3d5HYpuBs4W1jSHAz6uhI4Y/Eo0xrpHgGxjai9gwKn5rkNOUw
PAEvW0FyTTMsf9+pDGqc/cv3TS4MKNGuK8WEIHCfSE9M32H+3XcGpE010qQDveHy
yfA9sjxc+LaG8B2wZZSxNgvGvTyucALUMKIJ70CWKtqw+4RWr4P4DYWkU99VDn6l
LnZ1qeFUsrefNE/0KxNC7jxDKvrgvwvqh8thHbzGHVWHur/v5giuAGlqfKH9LFq/
EdPS5ABe6dorv1qToMQ+IlQactcyc5/gPHesR3OUARvnObUa9hgR0XaVOt2uGf1t
2aQLnwo/Ixb3K9nV3hR05z76VOmSSfRLHyy/xPr7vTZ58z5IEoTy2NA2at4jueHh
cx0q92yLlIq7pgsI6gh8udrl+/1ElHmXhxF4AdY1MvTcvoYL9lbo2mptcHgAdbs8
+MPeEJRE7a3KNzoxpJ75Id1D3LhyHLioqCYUXhQg/hV0GdS/DQyoBJZkJZ4H6lkU
WsZ8A2cVAI3wcXZ4nhAdlNTNKzbW5XTznx/vxggJLeJmxM2Hxns4z0oeqfCmGSYX
WUBEeMmLa35r4jDJJEqR8+ZCVGO/8jf1H9oDYCaKJ2Pz/UcM58nSCGuW7GmP3O6v
9lLROVqEQF18HwNU2mR4dXvxRLxNHb83BoB3QDsaBAP1f22f6Iw75o74X+iWofkw
/RSLNl9xBx5jbcpzGUMoc2X/ONzSJ05nHS+1gjb5hz1BZbabmB8ZILF0ji4DK2+2
FC5yoTlMoSD71DuXmWtOuyT+KoH9RklPjgJkacHZ63HVdYq16eWV/ZKANMnqf8Ub
TBNuJYLssNlR4WwpXJL7jsf1dYD4VYKrO+0WChZUFXJ4wFld4czK+JNh/yXxVWzQ
EN8Kau4mU2kn+sMNoyifkCEdmnGpa0CdEwCPCKmKUE2QbqFitVKXpI5DxYPoAr5a
NCIgEGWBL5FNiVj9+qLKalimGEzjh0mOIn5OTPS6VX4tP+6b5aY4M6W4A+8rSIZ2
Q7J29lpPXZn3cKc3+z4DLzLSl3uPSgDYrXV1waDgdOkJo80+5uJRienTQAIWNb2H
iBmWxa1Z9dsBWD+mGMbhOQfyBJrKZQ9aI6A4wodobWn1AsV6UcoGnzew0UQ7SlGc
1WcDtkMDQfM4NdrZuDeYtL2dzn3O383x3J3e7ny/FmnbAnP5fJZvqUL0EAg6J3WR
Jn4gcB1IiB5jGel0eDfwCgYk7Jzvmds9gysTq1HRXDMP4k0mXdrh2dBNNNLZtboD
/uHHD1/Eq0bbu5yXGzBss4emynYjcTb2OhdRtFcS96zOTfvCDbAzRnOb39PUpuYc
uRuaRsH6ouAODKyLOBzdb+jSb/pZGOz71INrqo+Hs1Q/zYpfNo3Wax8hoyGRcqjh
wMyoZh/QSu0aDV/cEznXmC7xKQxH29t9zkpTkOjUcHm3Q1Z97pra+Vs63TDaqmg3
nIdxCtjz8A5bZfV0QjsF6jZxJ/F388vP5/zpNtIJIrPtMPIuULbNVVy9Y+Yod8b7
GWELqqbOBgFHw69PPKJdSGkCs24sRKtupjLL0g8C7sYlqqNQbciZzVSbVo/liWgE
Vyf2DdDOVcVN9T6i+pXt3KzOifRtuvnNFECIAuV6+JFYrrX+kpZ4lGiHl/MMtVkL
`protect END_PROTECTED
