`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
acf+bFqQkFE0s3CecZutSS7yuW0z+SxxK0YW6JrB0WGOmhxDo0mMrE9PQLmvtqT7
ResQZocCt11Toii8BhqqRWvKfOISOgoFNQCyuvK55FtHBejxnjIDCXokAiT2uLpV
ybOcwQe3VcCbBCVTyqVTaOa34On9VEqAFgdtENFWmZba2TQ43ktNa41o0e85UWHc
Vd4DF1B5/SNWyFXu5Ik37LcnQ2s5Pb84qk8tMfWA/nPZqBQPUQVPJaXU89rynzCa
fFx8H4+BnB7FE9cRc5NwVWKymWqPR/6lfMRFlFYtqmjm09U6fu8+wKual4mZ9jok
zVOUHTxjZVxnZ78kxPauBpoZ15aQnIsX8NnbwVipuXJgCjBQ4kTGoJPxqrQ92fS/
SNn63oNJhIim64h+Wj0QeEpBDNw9ZtoVsaCYfF9v0rFMUUyx7jIsU+PYtD0i0J1W
9jhk4stdPSZCU/Swo4luHteuLivZ1I8ZLKYwrdmKB/7z4G9t5Nvquxzwkgl2AlW/
Wk6oIBmR9OYrfTPh5QIJwPIUq6tY3XThyiWebGlSykWhn76OYI8uTLJ2b2ucCdmp
uTLgbZnblpddToNAjC2FqYo8/eUh/GO9jF96/7Un+sFPDBAyBzt4bHCCPXavT/WC
/Hi5MGGnr5u8kHq9lx6rerGl0/a+mLsRiMX8IwLmrLSZUs0i9+YcVuPubyQcWqTi
YfCPraaeVJcjFvMZO9V//YbqTVI4fpGTVeFfFc+eUD8j6cr15XaHFPMJdM8mO7sU
zKZYB8Yk/84oI6Q+hCXgeloDGLFXU80MObP4VpJDU0QXlYI8lyjn9rPJz8trBFo5
7OO+QBzaWd7WsKVtTS086mlwak9tzy6Q/B232vqglbwp6oYk6MomVu9XzC4STxuf
mkE9tbENYmx1z/TID0lbhP9yQvvkuQ745BjbVIMFMrBW+mpa4+x5jDUm+NIZhTA0
Btg3v6SURnxB6u46RxfgFY/CmYFP/Bk7Wtw61X//N1rWPoFvwQBykbxaOjE6b22R
QC3gWU04k26AY0vs0CC47jYc2oBDAPJtNyFjfgQK4arGWcu34hqcA/Z0SIqMPUJY
M1sgPmvaY8BqWSFulLfqM4Vp9vBJiEqEL25U0rXFzQ7vnf43wtza2L59Srarexzw
zix7Gyq9zNf7NTvKedvdrsyCS9VyYDO8nDZrozYox+gg+iq7kIZO/7Bp6Vo7RK0T
wXGn65+jb7ajwGlwg77+NqY0HKorUJDF6mUhUyap58uvZTbU6Qnnpq4NfzEinY/B
c6SxJ3PV/k5ncdHf1PUUoG2eZ5W/JWQsqR/YvAUxPDmd+MvTQTPSretNLcT9pnzO
Bv1cFWb2AlMTzNYrBx/oZ4MQ9Xe6xHdS4kKd1Wx9XaVh17GrZzHkFvYZuDRQAUrc
vuXS4AE+rP8FN0eF9cecrB+dAbOUxhNC0AazV5z5pAAQs+YwdkTl/3551zMGDCVX
UETiN3QyC4zJ+IsEnUh5/nRcnDEFllAEvWi0UdEzvBtElPu7sXQMDijHQDPjk/jV
7JIsoBdFVnZGD6/tNkrNTCqNx1b3gbM5U5Sb0zngZ/15+pr7XcWH0N8VKZrxeZMf
Cm473HbLJq+yM4vUponjwpNljrgTuy/E+E4OVl5u45rntFxiGI2YBkysChdhsYXi
yV7z1T16KAXOmPnuwmwpjNV34+mAbskZU1KO8bUi8FWYZit7jsC2pf4ps5jpBONC
2KFZBok5QA3OmKjG1UwRvq6jFF2x/BiD0SfIiK9/nOzMWbEBVbSTHtcUXs4Ajke+
RKcpYR60tN0p6ONz9+4tweqcsUvXfcMRtC+BU4PFgEqUtGSCzrsdZQFj1E4O4ubB
lgapCa22lCSk+yNuLizMDIQutqN7g3dDuzWm5zdJK94Aik35ZAwCQe4O5+fqD8ai
RpXLsG7TF1u9otoGadmN5ydEDBHikXXmCSDOEL/LzVaiWb9tMmhKT8ZK/6uSpgYc
Bymr6jBNaPQgioAmKGbxT/uuvPXxTvptYyaWH/R1jHp4277BW1k5m3h+ulcTqVYl
yqEQHTjmbGLXDDWuKllkGovPLS8IhOuZ3D+bHmfCN6CMaEdf3fV7nkcJGGx7dhIs
8C2iSf5Bg7J6dJqpEt90gXJNHpqff15WDz4mwow69aV3Zo11OG0bg/ygMVZ2oU7d
WjNT0vpWzf7aPBBR4puWbqt5239MOwo95EztCPv8jTxuOchBqaT5nU0hKR/nT7IP
NJS43B4NSVzn3+dwerJkSEfJhkIpp/B0aT0KcYFnoOmBFdIYa+DVa5fXivvOjsmz
N/n/F9Vslno+42Wf5SYWuKXDVIOWif6ZenUIkolw7ysHFckXgC7NfelU6mujCk4n
e4CFvYbigztKV5tuI7s8VayXoeIbwwz8fVK1uYg9v4dbEMENdgeSXeB39GVAF/VM
uGsb7eF0p1VPTSNQr3gj3bes079IE4WWk54AJKcudzm54er06JbLmcFtCMfvnODC
s6Jk5sq0mE5gPVVzesFKs8VfKcTZGX8ucC865t9LYFeSmifeJj5AQlso/bG358NL
a/X8wMGEOObLYw2ge9Nk4v79lmj9zs5AN4Karzx65bKI1LA/HwQQagWbhIS764XH
QYV2m7gp7vV09Zx0OP5Jt/vSNKJGk3LLuH4EOLWxpb0Pi7CEZIybXl8mkYvwPgXo
yQQjsQAFmedS5pYhNVtsuRhvcLlDJN08wod+7AJnvDt/8ZfwEVPMehVWNF8upvZa
kfgKYVumVZn1IaYO1Xdt2e6rhv18CGNOUx7QYblwH2QZSaBwKVVJSM/Cqz5Eef/z
Zy1cZ8LmyN0xnKFaUfNz4ZKo7fB8QeD8GJSNmAHcXPngIPgKpBK3tYG0QUhWs/Jw
YELOlHklKw+iZ3JwT9jaQeBgi56KQDbgmpolUxqvcH6dqPmBd2tkW6TL4DFXwlN1
N4gHKerz+SqtDKNT2259Wb0/GJG+t8JVSuxZwSgYGMxinrxKR3+mnCtDa3W1X25T
xMhPvfQLU5MUOXpDCOi0CW5ju/N6X0thfhzCzSYZymsBEpsqqWXlFawngUAf2ywY
NtIIHRR8PBOKIkbW6MMh/cnUiKPxomz0KvVuu3hzddYkejWWBlA1ljtTRHTttoSy
UkQ9ljnByWadDa/3nVebsoaUjDC+vkwV3OmCTqoULlnx7+FGRatoWBC0a5OQBucw
qLyHieHwF7eK3uuGiIAOhkXI4AgE0c9YBe8zLYszRsAN5U69cpcVqCEb60O+cYLA
RWy+4jDWNdpntXkr8FQ1MDWY486s9tFrmkQjQ/Kjw0xXBLeU+i/IahYmdmuAut7i
1uufTuby387Syi8E8cxYA9chG92K04JfB7+eABoiSXYztJRVYaSIkL9xawLTs9yA
XFsx9CETLigZGhq/fgTmL7XRY7R/TXhi1ALxtn3s5Ptvdx48n/UEYRwval9dEb2b
sOL3sQpZAE44XlTz0iKglhmx5rHXVjgtL9zeb5pUOQdPZ69FohkYXUjo7oFKoErw
LyO9GIEAIVNUweERwFYbVmF5Y3bfJtXhUnQTIjLsoEVYD/6nckZ7EaOj6nK09RmV
y4jpwGWxQG9oy0EO+4pKOw==
`protect END_PROTECTED
