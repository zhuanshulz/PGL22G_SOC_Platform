`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jxOOj4kI6QE/RqjrL4mU89hBAwph0I7j2Xp+FHkgEYTHpIWzkCqckifL+C6PMOCW
Zp9I/DfkMeUpz0oSzLc5n5wDL97kqLHV0Uc1V8ydmpnbZxNefOKCZTFzSjWpu6Qk
dQdMZonX0NjDqFKSd+WE3CuCtPBwtvL6+jYJV8KI8SyRBmzn76T6BZ1oiN1OvTXF
JH/suRxHiLu+xHWTJrnEOHu9C8LBxwvnWGSAqUGpIMeH5w84RiiVfTtEayBzb0QZ
6MGU+S34V0/MbTq2xxjubZwWv7ugkx3PX2JPHUiwyXDe14LdZDSLte0QWo8U4Ssv
mlxTBxlAHuklSNYUrcJU5sQFdapHKet90XjXvbK6oX71KeGuInhVZ8GwbmzRY22l
1VbkaXe1W8dTTmGdyHw0sMtwj7b136aZus8rus0flVQxNDfU96MrxakMJzocEz2I
D1L0Mx4I+v/panQmVhxYJR6Z50p9rbPNnta3nrcqhWEb9GAoqjMDwu72DcT83pty
lCwtsU4hX6G8ChjWSZT8Wya+YSTjNLbVSr8O3JAdjp25f+O4gMWvLQkFUkndEMiH
SixS+guEZiAwqAbyBUE/nJ5ke6BeA00qMpbD9Iv/y188L39MlWKOtOwUO5ppWV4r
EgKKHofvdjyzskPWZ6Ak8wz+cAEKzpLbDJB7iuQ6YLzutA5WlzCsuti+S2x94GN1
Wtj8BSZPJXw7d9n0sAjkzhx+tvfj0sLopH1pKeq2/Rpu6ZNnyjKSpVru1JG0GWAi
0+ws00R37R+2h8pMWITiif8eDNE/7ckN0qHXPfCZsOUfXXDRa5xVntJ9rX5lVtfX
CxL/Zk7Rqa94y/LZymlnhd35vC7kNpJlEhBtkNvSqS4OeJCw9EQSHjR4BtzpOy/s
yjdsC1yjfzicHBrMIG8jNgW9Hgvh9pVNWinlDMQ4icl9I33rOWSDkbNAtNdnDxik
HQ4awqknPSnNYPccJAugjo5cBNF+jmWwUjC2Sj2dYiEAyaKuBUkmCqOIp9zuqJgW
VFYr/7bpBUp075QD5Hhbwi7dDQRJ1z0kpuzpVY2MMhxmEwDw7dKKXeEsqUIEfc5K
K/iouZwXEJKMZFYB4xCUEQia/3mZng+dvBxSyQj5zaLMJSalM8aUeHegB1U3gdZz
0xJlzZDfkxrFeoVULexJajdJpu5RBe3BaIBw9hHuH47JFI8GcdEwzXKYjFuv8YAS
st6ow737gvzRYVOss0eacCFMJjAawXgDIl+thkVG5I4j06e2n4I6+/Wgukp7/kWJ
qkm9elyP6LtIqArby79zxPhR8qTSMYwezrYOQz9C8ZPMaW+y682e5/6DYfRfZWjW
hlckDVQBNYXGQTLaFxwHDZvpeMhL4Ki0+Lx4O+6KwpjaruWpeY7tc0E6Dwp2mo5z
caH8FgP8Viz4UvyRoZlrVMp96vJnRT2gsUkqNiNiQBhcvLl8ADowMLkQ1lSvrO2J
bPFuAJPKF9eEz3p1xpUG7sDsBWGkdPQXr5ph58VCtZzyPC2NWOJAmCekXHTfm62d
IjunLsgEzI8uLfRpdTmRK9ZBcZANOpHFrIraXcAL9l100kp3wfZ7zZSfQJwqWwHM
KH4YgER/9HEvh2Uw+gI8DJwyuivpZOolUWCP6AYtqk29PbKaDl7cI/8iMnduaoCF
QDmS8H2e+fzYHYGLVEDVyo/lCJ6ntR0t4i8+VxWMVZqRrfJDJ5tY18JkqK08UflW
XyYCCiJi6oBAZEkMWCvFyTDyaeVOItXIYktchkA0yMKyCBhtDo2UvRVkT7ikAnFI
gMr7U4NbP4U+sDRiqnkZS7ZRifplyk3itb0Y1ohSwH1FYqzOADD6CXd8l6oM/7s5
IYdxbX07sHWpLFxTZl2tfbeIMg/UpEhlGyu1BNqoqYL0v+t43v7l4duK6XtIqNPU
E8Vmxh279iaAUyggJe4Ou4Ynl628yETqZZsRdxnOuu7rtOYnoP8uGJYeb6zwddyc
SDekU2M6fr2J28D5SjhuTAMKZ6VmU5aEDdx6B+sm7Q1c0UATrBDzN1TrVYBMWHXr
q+XtnXOX6hHMWe0uQbhMKYjSjHlzwhxRe5ELgd+JLBo6jFp5MTLh7e9WmdvM6hLW
rHe0wemQ9Wp6ldNJWoKHkl7aD7zCfmifba1SS4NHBhMhLLV3QCJ8caf9H4bx07W5
uQU6/iDZTudarVnOqBkVFw7WWV30RsmzTJDWfPwd8i4IvDhTTTotWiQdHYc0jcGq
MYuMRub4A0YJxBiy26adFxfw5rQEpm2FfK7k7t0rcIOb3FHF3jwvSRo5mBzkGpPt
5FiT7Q6UD9FF/SUw2ENMHDygpvq7ZvQPZ0QhK62d2vuyl+t6z7LUN0NcwYtv0dYQ
oRqQwTHbePZ6l7hoxKUYGvh7H/b8qMeYiGnBsTJkNbVtjTVqDtpTl0yBdLggO+IL
0HfD82X4/xvRmSjLBkhBlUMiWtPxVPBWpzoPGLG1pn5Xzd8Wrt3Nt9COyiOhnSg8
x7d9afbNQqL2D7xSqSve72aV5kutn5d5VLrlhKcFlsxr9wbFSXTzKoL2QDlsNtoN
jmbnn36VExMKcwftnb2wapiAHliT+2P5qaLbIVRHYZXTfW2d6f6ssamioJMtSnUd
qiRK4JrFsFcw9wkHK7nEYL5QoP1eCnW+JKNEmKAWMArNIshDYopt6LMtZvnW4yOv
WQqBwBRfdvpch+/Oxctgcg==
`protect END_PROTECTED
