`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rQBBlzeIJqEl4mBuuG6nmve3Caufl6VznZkbUL2QjxlN4N/KQGOGtnH3Jnwd1BTI
etGzpG/TjmpUnAbeb67Wfw0DzI8H/kukCLC+eLaV1zV97T5dvdy8KrzBBG63fpwG
o6y16e9Kr5EokllPSzRh8RhshsCjscmI5UDEChbETL4vyMTnDGYdMzcWoKP59Nr7
rLeiEv32d1AMEYFJiNWKbRfIjNoRhuQJBrwS/Jumb7kQ9vysezvleI/OuNLgfNrm
dIn4NbG72q+MpK8g3OMm+2tr8hbBX+eXPwaieEAyLb5xUjJSlyC3XVDzyaUnwgvj
MpyxyPpSmePH6sahiddXURnocvaopoYbQko93TjqnL9fKO8V6QWrrACnrcYMedmo
aMxBMOSMF3dixG2MS+cS8A==
`protect END_PROTECTED
