`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JmrneFM5HrNbk/ZDqGIyJqjIScgAlxkRy9QEADA/zw6WePVpMyaNVsBxmnCHd+ou
bizf864yNnQPvTB0Q8Hh/+oieiWjtJerweUy8xmtvTnGPrx72Oc99fwZe3lsbbrZ
jvGxcwJgp/8vQn3PUFhmiQHuTcfuRugyp9CJUn/gZm8/889T7aI0rlzFgbd+tQjR
qcGWAjrCxwBbObtO+wMdTblEdDD0TVFNB2CTBLHHgQ1queAsVNkUHhlco0C0E/wt
K+/fWFYl0Ment/Zygm3FeVdwTIVr33oIZKoeNh0w+NQc5h0GbX6OPuEvUEb6Uo1I
WeQg8EDYV3p/S+hHncMKWGOdGMq182ErEUJFqnzaCbJgZCzIICxdhaRuh1USx8Sh
llQRVFyRFpr+9uEYTZHE7Fyik56ffPseUu9f595600MtIC+MqOdZxcfHjXqZT2kJ
UeP1R7uW95KVJ5OvQF6Spom27moNn+DhPKIME6I7nO2mbwXtzJC9OlTWlfQGbGQ5
XiPyxCWvqzUnrlmwFKDOn6ki1r+gEuXDmUnp/iTqySdA+tGm51e1BTrEQ/RU6bsX
jpfQOUzXTAJp2b5z3+Td3eah4FBoc18ccgYJ2znbZDHneOi9ovnlxYyQyxQcRiXA
jjfqaXjrnvobMHcvec2G50v/vBHZcAjniOga2HBLT5CG6/wQs6evJ79CdUgojRfu
vDw4QiBEx2d4RnOdvJvJRnElUv2HOrCKykA3LeaPBtWSETUm6N3UebNTesgT4+6f
IE9KeqLjNgERDagR6Z243RDj1MkKJGC2GCL8a34exDhy2p6v0eUZ0CUe3AKEae4j
hGm1PvxfoZrNR+IjBvJutPqez+tFZIn8PKrLkGg0IO3um4Ds3QxLuWsas5sDCzcQ
Gma97IflyvzdicI+24Fy2tpYxTrhwPE+vqEaj4oJtoUE/rzECN9mo7R5lq6dvJaQ
CKZQxGcpMaUP+imYSZkLMhDArJK7livwxJNazlWOrp2MREAInPUARpfA8vzvEwPs
yKxze7PN2uQKXDdzgObOS8YCB5l4a6qSf3aRbmswbMw5qHZRIlK8OfHBJ+92BX+M
VsgkobzX/uRJXYNIQejV8eWFyBuFHL+kdxhLI++JmMClDigHonGLDvHo0KsKuWZb
y+dh8Cz0mkDcQxgnuTUN+yGUYeSaELzw8EOhNVWL5aFfK9eysBgr98fg+EzmKZdM
hl4//stAis9Nvo2vkAPIWYmHk16FNVaFTDuU+J/BGdrmOyCo4SP6aSqLoYjgRT8X
TPbfsjkft/dIFZQg1Gi39vgJx8qfdOI1ld9oDavSv9rA7V1cQuoSa8FCG/xtKgGy
iTHOozmndF8uSJyDiceOXtuUtpYhVw0iwtToAAMQOFfsOkkUQI0Rk28kJQj8MxL9
Nzxf2lX8L7HrluzWTFcdRuRn8ohomWjee/I/4heeG+HrkyzB5r8QXJwwlWheu+Wg
cCijwx/eaaxOD1RH/JUjXhK/MkdFFMRqnvuIi79yAcXb2UfJGM7QAJJour1xO9fg
ZMFY6UQDitbLvsv7cScXyF3uxnh5619ubeI7hVEYLQZD7c8jpwvCpuRZXYzkW03I
uVcv4oroB7UAdHwNyUFRqm8eMT8Lt1BUvBMvPHQMWJQN0+C6p289TUpYpeG1TvGS
wE4kItl8hiWXNf8wbXDun5qnyZJUgzG/F6aFny+9nhFzpv3R5CzczxV+k+xoUHgE
+/gc2o7t+9VgSKkADwZLEGSiJNEsR39un4MmEYqRoE6FovtDvpoKY0sNWoK1wJZG
FJ06icgTaMi09R9ezpQn0SyNQSvXS25vU+tMpppTCz6I817/xiBO75uqykom90cf
91Dl5C+xIs3EcSCVMM3Zn00I3AYe+IR5h4Gn1u05xkHT3nayo7kIcS2od3PUSM24
qq9HoH3vy7321KzUABrzeAE9M3l9/q2wfSKD9aEpSVvfUqjVFTUM47d9+ZtAdIwq
E+xQu7iGGKa3llMVelpaOe8uuw4mVsYpips2TwjVS3FJlwsMx0mI8cQ4W9Xj9b72
i6YsUDuyAVGDnLGmWLs43KDpHB02CxbIi48Xgzrv+3RS1OhZKaE3Z76jFOt1SXM6
EYRxez20sfMmpIOudRmdjv3zgTsq90cB5YXPoHmjpleRXDGAJ41YFx75Jf5Fs998
3PNmR3Fu9dXRMT9LuArJ0mHBpFX2R3iHnNdHxleRsLzfOZrhE82ZRwMTIsz+whE+
IHd65nqi39SNI1HUvQfpwldzl3xtIvmOSVfHaNnj2fH3h/4ShIbv07r+zKYkzX00
SwX9xLWKbitsyq6ARhaGzgszQAug9Kxc4tSVnqjmzuDMc/ikOqRWypyfBVb3u2X7
s39ZaGsNTP3UdUdYqalUBI9IEX5rqXHqBjzkZDHuXAuHd+utgF2ftlA0i6jAcwlc
urIydHVVZwQwJdVVY1flT3XSDCSr7Neu8y+0+32PLboXO4WeoI3nQuL87FVO9aLO
AHdjfF44Ym6RsP7V6KoHZMz35Tz8KMffx7TuZFd00cKaLmXc7n+etqHCRM6z1Obx
IksnfqTxZcnQrV1epY8nqKv95Po+Bm8v7LUDXZfwjL9Z8IVbTy0nYfqJD/tK7WYq
nxvrdM9+36u7nN9xIarMp7XiH7CPxljmfIagUCtL16ssWJOBA1dB43BUIr/8E/OV
EO7O02h3bwep0sEsSXXuyfdaU53/NvAxFaVE1L7bn5jQPArjVWnMHgCgYZiQ7X6W
RW+yXGUsMkB+GKObt0Xm3mikDAY8R/1gB9c4lOAj0YyAxT3MncPDmiaJhQa3/GVL
HxIG5PAgYbPP0xo+ToHVEOqs1B4KOcgaer+8lE5VOP6Q6aWy3+E4+l39CfwEn8hg
xVVjyniBF1XMNerHl8IVC0pesqbk7WDXgq4/gdYjF2umVaDQ/5GrwrzZnaOHJQ5F
4zxepo96rASp9iW9+UCZgYAuG1OOvG9H5yJOQOhu2tdaiuZdQiKUH2hq5XO8msKU
zHU5qE/BXT765tU3aAP3QMRqat3bWgZlxgDgfCr/wrMvux1oX5uRWYgplge47aIE
UnWCScbwVvsKGsUUj4Hi88K3AihKQF8Qu6W+Jnhf1YSkxLHWzqKfagU4Z/2UiMS6
fR7LVoPjeSlZVZsZyygNK/4zHD/gqmqzdI5xNW/IMmtcSa7hSQZ6F1UI/gHJqb8e
gktpxzrmWDDS/ovTno8+lp/Ipe/sQoJPiIpPVG7WvVLnDeua0IQUTRjIA/l/9rC3
eTkaG8oR2dbOGfDXM+mpqmZm16sXEV1n+H3f2HzVwjyJmphjZrZF7LIFZnvL2MTG
oxjL2mWYiuXO9lQevWT+sw0nJ/0KN88YL5opwUuKkhEzhJLsFiPT5awXsMsnMNgq
Rau5/UHYeI2BtoRn3wQiy5Gc28Vcsf3VY/rI+iCzenSAvECto39GJNzafBEK+Vn/
O95d4GligF7O16hj4CKlu5WJ9//HSxaRDiY3RNwhpJoJO8ueJUvQ/xz95XS5/B1K
JsnJkkTX7OxGJcynVTYJ14egYGG/4HOjXiA2dG1hBYBP4loTpO1IgEJfl1tD68nC
g+hLOZRU/RBwbCvf/cWPk5LBMlG7Mmjheho3KLOqRlxrqqXyiX5FFBcRvSUGBka/
xyFahiOzwNhLnhEWEYkgCwT9o50wcCS142oB+STUOZG7dOh9AvlSzTDBb0RNg4E6
HhV85b8lgBE1m2ba7pJoe37n4BhusJPUd70VGR8vqvcHI2J5qprmPo4Fd/4aYs6P
FjIEFR7ro5M6cf/cG+578zQHElHkQo+Rm9VL/JIOxAp4DdGRv5Hfn987dsm2Ybcw
LVXE+lULXdEx/0Fm2Wj2e9ZoM0ccE6p7ddYPMtNMop7tCQWTW2qNwfv4ZcQaiCeD
1KeQvIsDTv1Buofqqn8rmonYAMF7y0EAqaVxti7ZKdW0+c6SLpCUB5hIjW+U1xtd
ECsCw4HYZxPrrs/9RSSIIMsHrhJd5VQPuivDwqFecXIdcK4ZaYKLu7fh2kUdUsIa
06q4pElqV8ceB6+n9cJP5vb51guiHePL+WKynYNVZEc6Bk3Bf8C/KnVmX618l+y6
EAVvvrT00ihCPXnavq0wySozg6tJpZ27o8LYH44Swp+2iCKD2V6Y1kdRzMn1qtyN
Q0Xgf7Xwe2CpNEMsPWk2rBck515AGswMHLslkhWRFqUqExUD0KNR29k41pVwOdhe
vbr1WVF0O0wPRtK5YyJst4jxY/rL8OeBGAC5M+G5H5UaYgiP5+/aHNzkzEXOGW5k
DeZjFfMsVc60noOl8fxa2k5Dh2AoVA81EKDtk2nRPiN104zmGuHGjnb5zWtL0JDg
npHURGNYDwiQgVhH+yo3Gi4y0uQYm1d52z7Eyz7n21RmlcHeCPhg0e166mWJCjft
2aLu5t34fC7sJ8vsMokBrkQZIjkiOu7PE53LeIPJEj/wehzLG09DRD288TcsDSXd
eMIy5aKG1BGfjsUvyXGvnRZIKe6eQvg5q1CK8ieMggJ94Ru6GJlK5jHhg+68yx3x
4cHMVjgwu1KsDREUVNvjIm9Zdo9lc3X9cSOhdcc8T/Eyi9L8KGwFDCw7IHSvX3/c
iaMpyPba1Cp20uQOrdcZcs3jytZDYdRwQBksVCUbg8TP/kHPHo/c+98WkLp+WI55
qjkgWjDfba4dbMDB5dm5gbKatMx5ZqmE+Pst6lPVEqEcvK8VLKKdgQyLXuyxtS7X
+3Z+wwhP0lsteDigjhIiWVoe5B7fo+lK3N9aNhLaBTExZ8PmZeOpCsCbl+X1dVkg
9vWkDy2gL71q/PdqMS5aW+PMu405CDeTAfQWzQMKXCnkg0nWUlsargXAWbB/8ae7
5l0ht7SJYjxCwSmDYBHs3FCxfilMCoaI9PwKSSt4ys1idxZvsu6T36D4p3WTy/dr
YcHPHofuV1z187wiqStjOYjTys5o9LpsyH0GWWL42VvyRzeJ6kJaTKbeRH2LoME1
x5vgTMJMPP3TDPsHaDejiSFQviV0qxXYcMCO1dMvxX0NAlmGj8mp9R/s3Ju0mKP9
ZudV5KibKn8EsERxTbPEupHzGydhoercKXbEPmMXVPcDcsDxeG/h9NXH5RPeerJh
iT0ENI3kj0aLJAf5SyfpUpBTHCUPwgiWliOXuzMmgzVitMMa3ctNqYKrro5/cjIl
a155tKO4kKsmfG6U3Vy82ErSuZiGCxLHmGDZ1LQs86erxBYjRSh8Auqt27VayH6u
DmcNfQ0I1JknA4hitxzoMRe12T1jdgxzK8yc8oEtEO+I7tnAlWDh2UTG9tcuh5W6
+rYywnLJL1VpKJxP3g3c9/ASeXACQd05M2/yipbjGPsI7zPHFbhGl/OZPi2xTB9E
jFYUSar5jufRkKBBKSQzv2fhE2pZPapiRCe7Lp5SWMCe5J9ZnwLTBFqo+AkLp9Ic
A1+0WOW66fbzefmEGKSs3YQflURa19oan44s6DeyhXXecAuv4UCkWyKlNpDwUFYj
8PV9uYUfrNEBI17YYRyowNE328ANjT58RhLe6tCO0Th1rFher2lBQHjMwFM4Psqs
pbXiOa2neOOiOiyZNYnl2QSR44oB+f+qYhGIQyZiu1cGr48LjJBQFJVLHgcK8Hng
gPv6tQJ25HYjpbLArG1nkIn1nSGiiBbxoNoW6RorGeIJHfDn2D+PqH192gaJAY/O
pCljI+XcJvBQTgyVTD9ocpZ9sgDquPJiwBKTmQk8tNZChcvdtYyFyQYfsCv7LQkO
YtZlN4LmeTSYn/SsKHTbYbM4kGTW9z9wEl3Tv4ihIdTp0NgInOEatUGLEmiClAUT
ZlpoLvEtHTeJJma0wytr3nJFDYg4OodRLBgjLisUmo4Cw81QdxAk283jf3yZsZYZ
NLeTw+F0RDIif8pn2fgzJgOwm114YCfmht0BEqVGCw/O1omY98hE2Pv1Z0XrOugS
oWtW1OzRNtbypB/B54rnNeG47nXjZ51P3ULvASq34B2jk9ZKUGBEuhbfyUk7Afue
FHhOJnWS5ux0FqFbjKsbt5oifjWUdzQqgWRUBaqtB+FAH1X0RR1YAxlK4JPiCUyp
Qr0c6svUQOfAMJkQgNXXpFg6oNqZ807FbtnvWdqH+9MMVBC8wUmEL16z4xu5UFm3
ET0/s4F35O5pULL3oATanqGqNpATvw0+WLizhKej14Km+LHQXLUyMSBSJQAmWte1
YsRVQ48OvUIBybB6O1f8OylO2KzcbbeDHc0mNOHm8SkD3FjbWCJZzkbdPBUFGti8
0Mr4Oyc01SdWIl5fJhNtFqS52PyVDUtduQMqCf4+NP2ZPwGV2MvbzX3lW/h5H1nP
Uhc1eKXHAcA2Xr0HJgUYGvd0JPTGVXEiMoLYfRvE3Fhdg0RukBlvd0Bsnbt8UH/H
0qyXxdo66sHtJNHq69ZikaZB42U+LEzVK2fJrLu7R8+jw+uLoyk3TxeHlJu9cniL
Rz1ZzQU13S/Fz1KJnJgdRot9zFhN+Qi/bvbYqKuAGm9V9wxDTnB6v/+Nr3/FtWmW
ObCanEzRtSQXWqgi1f8gIFUj5nHGh8EJoXrEZXM06pjpfAn+CIAX6U3tU8ufvb0L
ks1y8W0AYW36b3MgLH2abiKAFX4BUoF8wMUGZRTtGpAUBC5etvqucZl+3CYFUHI7
1UuiZpw8271pK5ROu+IX6gmfDLeWq3cqG8X83v9HGBW9ckSsUuyNqPjOg+yYtWpk
adpnZModM+7lwRlFota2KiEag5sYwwONw4PUKFjtfL5lf3d/j9LrAK/YK0fKeNcm
7VBwzwR2Xjg8P0Im7TMZRhGSEPzzUVm2656NJne1jhfomuxUkTXy+tMaz9oydj36
2G0YmRsF0PWEr3qlFxyrROo2Kq74I4Wl3mOO2V9vCCaGeGipqqV16FiAE0YvBVmO
6BHXhSGyU9F9jcveEZKMgSEq5sCvfQH9Xrz8VPN7aMZ3Ew3ExlgDHHjHbnUErBd8
ZYA+dPoJpbCB79ieaxMZdYjRRyl3UYiQiPzu7shaUGLNESRY9QKOs6KDCrc6WpsY
Xa6y74D52cx2JN4SVMUh90nRmp5GR6S1t6I87mlti+uUoy+kHYVyVDA9XsTa3DS2
42tmdnyR4Vs4Lt3MatxfzQBJEzRS+lIcNYehg9SXY4FLxsTdYb3mi9CDgJpNyxDP
Tr9sbTAv0rtTa83VV1p1NW8sFHerjuN8XmFOQtxDD494gGt+ooERsNiOdkbATCnb
UVyubG7Vcr2hLsBG/ZkNRNMu99xWnbse5YN/ZcPg2/I51Xzs4LzSIi1sxM7Z2u4a
q45f4+4qqDg0lj6BulknEwRWvW3YN5idsdyqMFCm/+xRcsAHgRecpsJhEsa/b8JV
aKXiMkOV3/HDkiFm+i9Uqa2PuIqyhNHOKALI4QW68cOnenpHPMkTaamvZevVgVl2
pKe6PcUEDZORQIu5hhAzBY3jSSUiXkG4Q3Wpdv8bwnGxCca7Tg4VoN/OVbYnKAe9
C93l18rnqAn/meSrSsBjjEqzuQNqarzH4MliN+2yE3kh2nbt1J4l7UCRJmvP22dn
gG4opPGr+W5qan2ThxRAD1u5igO6J8Z/QpfC0crl7aVxNBqLAb6vSDAV82oddHA6
GzbPoekCCdAMCea1y/bXZfqtN97GzNbxlv5W8QPi8jeVPceRETmg33yvfv0LnhDh
GlGrYSGXyXaMxZc6gziGTXUSH4FY6ld10YeHkrU0QGkx2BsLEuhHftUT0eyT50UT
ArrDYUMhGwDPWHcQ5gkn69PrJNjeikK79yoqBZ1LrlUMbpRB3h7eUNwiWnXpVYSW
zclmu09XFodhOqK3IE2kQD+jfP5IiivVz3FRMV/2nA+SUaCwfvdtmh7OagnBS/aY
yE6HGTdu5LfFfmeCVxNSDRB0ZbmKg2icAqOpdHGFNGVU8SgkxLN0cqdm2eoa2IHb
iJaAjsB2E2sjq7E5IkdAjsVb8Q5pozmBZUgZUQbQWz+ACDLs8cH98JmEQazhfvt3
+TgNBksLdz49UbSwXgp6HbKuBGuyhhv+Bp67SEpOnnkDK4QO5hw/ZWxqyznaiQTO
A2aNY19eYwkwX1ssteMvVW7OqB9l+enSwjAtRSDrbB8QjaRH781BIuJ3k0ziF+vB
k7XF4MpEHstrS0mbC+jE4eRDmWJV5Q0c9Lofg3rBkHL64eA0ZvWKvu9YKFsez8tP
bqJPVsM0pHO19WO32Fh75i1Rbp5Bq2+OR4L+C4yrrEuWpkzzt+JCwyqzsV73sWCe
Ro0gQwhISd+3QBlRk3n8dht1i5MGIretOWPoenu/HlV9NiLLWI0dCGCjBTWUhuW4
DMNfwG3M8VVR9v3DYuk8N28z9Sa+7ZngZpjVkLxlrDVy0W7KH7TPTYMWvuBc2ao7
v41jaO693mG+871S4OqE4qWLPnQZBrVdATxi3CHNnU354kS4r5tW0ObLqi5e6KMb
VctADUTWjsHEcxXW5BgxW8KMdfkqukq6+rjJOIyw+caFwUD83/QHakYX+PPQNE/R
WbVlxdGREq/A4dEmN6BUMUtxDSGnyP8ZPAL13Ru98c8+QQmGwembcjP9tbbHvvQb
ubZkPxQ+TljUMesNg6L4QltjR7EHThFU/QqNg6epGOXdZpKVCTwFHXNOyfxLBxXC
F1HXnrji3b6wKNeFU8xPcMFsaG2evzEE1wkZvoYf7rmnPY6Y8c9b2/9XthuDvNk2
gCev2wMUowGM1k+HbP2fWMhcsUKNdqbZG4FLiaSA6aGg1cUWOH9TnPifRtU3oVQI
8J5vvkRJcRrIufauBJtBAnsBHw22ZZLOOgAw0lvREZu57MQiu4MVbAIo5MxuzSpI
P+3bTOaH1F34IHnWnwMfNdGLUs5Ssl+TIztDwW+SBCUhz6Jppr23toq3KkUxwW/c
7degIqsNG8L//HigcjvbZnpDYsf4C3zwAGy0g3r4HZS0WWN58tTtyvyuXu2Ebs2N
dnoDbDBzVwW21XSTh1Uj94YSWmhmfPx1P96iNCm3mAjHi6XXCKCvorxgLu84nfQA
azaGbAFEn0kM6XdEXZ7QqmB8jrO64qMT8zs6W2S+itKvRHt2SZW7Kh6hS142ADrx
GBv0KWCaodFy3xYVjjOAnaY9+lPic0lQhnzXwnBsneCsTT2Z7+4vSD8aHQWq9ycY
KZ16xuJVEZvr+VqyWcdD/3XGhtKcB1Kdaw1M4VKbjkg34UQGqT77RXam/Ni4jvK3
d0ycJCd0BZCxkcV6sk8ebDhHkxcPJnKIvpYKdY/fLspGIE/1HhFOoJz5zIt8jIuY
zs4Lc6DYwdoBpvQTgkYSn7t8PSWsRH3u/LL1W1z1fRJm1Vt1+VDVjSYAvGg0l+Uk
reXPSIlaUGZI8d1H8BHSYJWXvfBMo/n7K0qWG+il7HUM1djnuNbs7rRoi7HfI7c/
5dH+Ycw+pfgQ11HrG4k0anTleJ3E9QMFbwhJ4L1wqQZ3g1jWUBP2B+TrhIuXxgf6
tSDvb1s+N9jNh7H22FGIBw8JmhL4zF7WrkU5khgKksnrtBIao51kvUmBXCxPpCv3
d75i8e3pKw3yrpYX3TFra05xzgPPJcrX29lSGj/rnmKfjt3DxQlCgdN+Nfgo49Hl
eZQoBB1EfVWkpOrnXD25vrm73MHw8RNd1My61AlYiLJ5TM9GvZI/09SoeS6nao0C
OsGQmC9BKeodTXVohue7+nqUyvyrgDU6JlolCoq/P1kb6wjDZIdiIQhE0yJ3fPcD
GroEs+n213bqZCw9rDyWPNmkhn2g57p+QVBvyDlASSFWqAIX5vT/k7M7lnCliqsh
4IDF+naSj0Yj3R57YlOQI7xQUt3PRCmzkq9wYLyKSoq5Zwc2t82TzElwPRO/qOsK
a5c8l9TThqHvxqik7TEU21NISCp0RRILzY+9sNaGaC5tbgJxy+9PAgAYrAmHSJdT
XmrxLKp6OpIjHkGeZVOdK1HQpOofuhzVyKdgRtyUeO+w74xDSnYDO+O0lr9k3boH
2lyq6kadde4wpJ44DPVOzIe0e1cCijWKi5gCKliHQbPUJ5Tvic+07U20iEEqNHXc
Pvjjyp9EoISjWwWcpebOuwCzvXoZhjOaiNgzhpHZYnK051hC+GUbPq0hphiH07Tt
cVu5ZSM4pukNmiKkWi1vE45Nt67ohOYwq8fXK2pRxt6HWiaWA811F56ocDD8DRHS
0fESB8KLqZTkSdKjNc91zSzr0N7E+8rNA2qj0HRBqhLDgKDGev68XQ8Y+BSIvNQe
5QBomto+0BqoVPCpV7AHUFsYH6zY+YN7xMy+mQynSa8V8U2hfa9u/DKk7zmE+RB0
p/An/FQUUCpVBVrIrKotPqQ0ipjn0N+r6NkM0RRAmtiVbcgHFB5hJCeyKVxfCce8
r8e+kFG2I0elgvESHOuxooaKhORyO+KC9Jg4H6OvDTzTHZ0hoJTiFmkJe7rSOO7m
1cpX4G9BC2Uou5Pad6fDZl6EzUZe1Lrj/iw+N6z/4OvHCdzbY5SbK7y1x7/WJOD+
6AEl+F2gXffA9oYAP1trJ94Y23z8A29kl7t0kNEqn004fGAxqjHp9wLnkvJSJ2AR
t4j8jRDx0n0tq3WTCF0PlwrS2NNMaQ6Y6/gWfv2St6gOpQl9TJVSrmLmcSp+q2gE
bndPl1kY/Tqgy8qGYXo4YOQUMK5yufKHgIPlmvCXTSDp5Uz4LLejACtQ9CRFDLik
VHJiCZ+CyYSAjDHUPMcdppiPFT3hWm56VvBdtB/x4117+2Vp93bsh/3ynqTEMGni
TakeH73Qv+SpPq13jZCFPFiLiQHSOWVX3hXhdDimOXrOYGXrjshOrK1z0aXSr3Ik
T4CVE8BrKdca6fnzHtyMvLbl/7SmCP87J7Uis6ph1//7lpa1d333av6AMbxPUlKs
Q8suAKSUOaMZtMhJAtGyNztVD7FYUaogKS1GyzKRpYLtfll/wcuJB7sA7wJInEGS
T7EsMTHH/3iibIJZ9/z6sTuEHklQnki0hbdbPkLPL/MorFKWKwsSUnXK0LSa+IG5
C5hZs7tGGaZyUTOpFRZZ5HHZ+SVgvIPMdb3rhqXNCuq2WraqcMjqQS/woMrbN4/7
IpCbKq2HM7M5Fy1LGEOIPX0tdOKiDekNPPlLu4CedB9HHZrEors+4uPzUUXYUygC
rnAHK/fTcy/UC6dEjDjfOfmETgs9pKVCHh55znNQO1yXFMZKk60vx0W1ZalgC9q3
ZGdE0soFUDw7Kt4J66yeCTmwMwbEotaiBPi4FYW4kdd7FnYuf1dvfJ92ELzbKPqx
1LYHYJuNMEAcbaEV5ieJin8nv2dWTSoQg8RXfbKfswry4XaPQJlxbgjpyALJjzde
E0rIE4Vl0AM/QHIM9gaVMFI5uzwIJkBr9v1lyJplznTqxIMPSaVRt1mbLuSRrT1p
6UQ0qRBMb/vqMISL9aNnOcgjzQpp7GFDIRbSx3zwY3YPcu0sWPMhf0gyfPX64Gvb
hQwXSUB1nd8OPpbUcsv24iIxiB5HWh9few/loc5C/c+uoUw3lMCxsyUVSBom6c5j
5RbW45mB1BIzo1inR27sNiRpfSAQw/zNR0dQCH1iHOLxkzeRwRK3uhBzMNenZMY8
aJeF5ucVli2WNDPH544CzdHgwV9XxgmVdlWGzEJl/8YlQrLXTJ5xu81GfCSXDeGq
R4eN6hst0bid0x06ZRBwhztCb6/CMI+s/XiZ7BocETnOXrC3vyUtMzm1hCLMlPWB
+L2E+2kaB4Ayk8LpoLVeaTfBUWuJ4g4DTgqm452WAg8yl/cQyQUl6qE6cbWGAKsM
Y98WVJUBnOonlEsfQK+V3tsBIEe29DR1N8eGN58ARCoHupHliE1cuJ2yIbDSzFNI
V9sBMMgJEN1w+yNDN/7JXO05bm5cWfw3Fm8xj+2lg8kUNy7hSMbyg3l6f0engOQK
eThQePU4NjczUhxxVmaqRnvTB1yG8wGAIKcavl8HY3+00gg7Ngckp3RMQl3kC98R
mPPUq612CRsMRNnKXWrCfWE5V9cGkQ7gQB+ffwKJj6vg7HL1O2Uc9cH9/PwUvfwd
8DxDNwG00wwBCffj0Tb6jqsoBNsXMNm34z+YqI3Fn3WoyIbor6EVKuWz8yJmz1Y4
BWCD+GqeJWH2ZdX1CIniTXSAAe36HJ+FwOULsuyEvZw1iEqeyj0Q4+XGe5+q8RB5
nB60DXu7MLl6QdvLSuNwEr0JIOD+dK8lzqev7UDyVF5risLXeQGDwalf2cuLuy+Q
fQqpBFzMEv0j83fXQpYUfk9Ych1xMpysJfThljXTxwUgm1F09IwXoX0kw94YNZH9
tw1SaDag9KHXEWBGJx8vd80M8wUw4Ty2kLJFuLohOUVHm3e/hG82fiP929WtK5o1
PcskiRugbnyiO+JoYaR8Hl7ycVxDCLyde1/yjlzSB9bm6JAsITHFLnYB1CkQYbHZ
JluC7m9cagPDXkAwu8tQsaP3XVeZCpvJjM4ebVBVRQztECM/dPbvyFcmaRo7nHx6
Nq/b8paw4DT1OE2Ly/+eyXPhabT/lc+l4VoxKs006TAnICOja8TDeMzIL51gzeAr
vQegrl+1RZtrB/23m6Ij4TUMEBvIrk5y2ph2bxdO3EXEOPI6+2697RR413yCPYJQ
fYgNOOasGCDoGOFqH/cWF7FSMXwVIukMC3hNU3VQ6ml51x8Ic3B59j9F2UyqaYhI
p2U6ZXUDWGqB2v5zJK8jL3evAv4/bnir2IU5MLwDhmbueMEpzmTUlVqFgLolv6/F
wYhGRc1T9+Y/a8KoN2AottoPfrKxMh6RkoEs0N2SSTXQ+oMWuqdN73qJPRBPkZBf
M1ua4XluBCIEiR+EJnidU8PnbNtGsC0oCbzYjHJK3zwVJ0DYRU/+jtucohxK076K
lcoKlu4LcuYfmBMZZQQGF+xwaUqVs3dYJFhPt2ovH3jIviKA3Nvr1eO8R/CZt7MF
0Ezwx19hw76z68k0AMtOr/FYYFIb9hm05en666t3/RKKvoZmgfhb54giONpEvfhX
6ChPE/qqaFjEFglO3/ltxYUXVIHGKsgqOeB49rESaic41I4EgePNyjJ4VjgZDh27
xlAL8PpGPfZ0yz6doG/vuDP0PxU1X6rXNXsoe8wKVXJ52PimAH2k6Hka2PKwQK98
G1P0JgSvz107vAcYm0h5KWG73EBqxXWdrHhJbEHwrNW/e1QBjRgmvspOvEhPIvmL
gTFLF1qhJ3gA1Coy0mINBVRkgNanhUe0oW/XaU82PJ6veGtIQG4NBldAUEJx3mcx
VtcHYd5JNn6ykeap6PKr3giBE7xkuMgeuTs6LG+sA+QKNgAZKoO8lnZCN8BbhSRS
JSy/oJGx5O6XRQo7mDRJJ/KnLNOyK3tddPWu4DKIN95OeePh5+aGqCGUQaJba+NW
NkpkwBwuvXlQ3/CHadBubTDQfAzcYbvX+fhn37M1+VbZB3Z8ldPm4EZePl3KnjoV
FEkllIp9Y1pu//m12UG3HLXpes7wPAetfrHDYdqbuPBxBZl6UOZALAshTEA3vpGo
lJf9M+U7gUmoZ/Z6dPIpLmNVbbXHUEpOT+5LeKUCJDsft6FLCWfCsLF1YJFERTS6
FRrzbRwU5DQPyhS8I/3800MTA4rAIgq8dHdCRkzIV8O0/dZvBvMS/rqj7o8BgDSt
6qH19Wv/ueNR4GOT4yPnYsztzzbG1wEZ8uwcg3e39yrXw8CbI9+rbtTke6IxE4Zv
VEs+xcBvpBcphz7B64wAq4v3b38Nu+LzM93syZy4kVABDZc3IxWkPjvkizxFqEpD
5BaRX98tC3pPpZTXOA2mG4mqJhuogdwqpcYSlBKvPRpciIweFayS+N3XGE+kWC5i
931s9NOqk1rXnMJkPtSzX3o5T7EwyDAEMN3TPINnH/8=
`protect END_PROTECTED
