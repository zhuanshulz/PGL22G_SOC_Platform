`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uErpXn6WUO12DCcWnAlsTTlgybCI8mgAVcvxVxXZCZ/Tz2VOcH+gX8PbIqTUdeny
rfomr52f8vy2gbPBrfY1qgQiurNyhCOjwS2lYiCTR+gbHTLvV1NnfjyxHZY20Z/i
QjN8HozHOCSr8Vkx1999dXff534TAPGgOOltOsAcCGE7oZ+or4n6ZE2T2OYSO8vD
zXr85ae9/gtYGM5lZxh1whvEcAsemK8bo9+rdjGKRANWQ+wEuKvVfwYazV1Na7Fv
sO2TWdVdGdCkePHX7TjzC7pA0Q1Yunug7sRSUDDwgnK1ALgCaFfmxAXDSBHw8qZw
2J+NmQduRM9OnmNA+FZ2cBH4pC2qGPfnK4FuS5zSFGYSbzS6hJk8ezjudNYC6NxS
zadYej8JOlcQ8RQNnmkD3jG8o5tUXiotXPwLX9Q2YifuKhjYMCxZ0B1j8BOnW01r
GbwuGJp3mKFmNnqdVPF15gJs/jmY4nFfune4G7VtNSrYQFGzhjlYsdbYcSlziJco
kWQkpcp6H7GK/UDvfocGJPm16/tLP/ax2i8ku2X/Ndt1AU3cU2IbseWmg6zBQuR7
p/TLFP2EtaogEuIwfiTERw==
`protect END_PROTECTED
