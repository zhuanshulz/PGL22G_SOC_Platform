`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MUFX6bjkW8Fo67PQlnQ3K4b3hJCyUfoULi+wV2CTjCawLB0kUmJOZ2rlpkYcj/oP
QK4HYIXUWMc2kfG4u0gkjszXtsYD55cwTtV41iPEugVx4LK5d2B2n30cfBRZXc2u
gTzZILAMNu32oRUpm44ErKB8noEKDf6W8NTC3fMHpMHt+v3TITNJu9Y6jH1vUOnw
m1/KYsdx9gBJKfsZic+VABa0IIV9JBGjUlKDqXpeVCpmUYBVXqwSgVbUmYGUWrVI
5XgChbfu8w07Nt7uM/y3DCCFqsMl/9knlEa2nwTiBe+EYq+roq8lJkBGOuIoMbXR
JC9+OlsKZOY9HO5EMHqaajpEFg2KuuuWdr6woRpyFc3TYeBWl5l3Z0PXUoppRuvU
HFbTUClKBtay6la+zcfCA5WXz/2+++QJPiS35DY3vmQQPt5kUWjN2oIBX0YNGej4
RBSw3x41vQndZtU56d66zoVXAX5enVzLHwbzQeN9PllikjL1CE6/VGjEJHNtAQSd
hiaZ4D1R3Muo9R9AG35SImKWY9TBarI2X4IvSrM4UGnIocr1bi4Wusd3fOiw+9Mu
+Ikeda5uYleyqkYmhveLr0POzFoKZj1Qfiz22SLkXlO9SIdMu+MM/ZB+Kf/JxtrC
yqnBNpqcqa86pGqg7SxmNZatKRqYXpMAZ0T8SqpwqHjt1RPGEK3IketLEHEO1/aF
x1sug7KO/CTvB1hrib0iCdln57KMmHf1AjDd8Nw2EFHEnjgXxMcZNHVUyF0/Zysq
XI2/pAgiFMG7NQCLk4g6fpdTUuspbroOBDMHpYIvI9ize3uM/UJ+S86wM3LrayF5
iCh8+TZqBMG8y0Iz49GfPn7ng1C+9GcuAEaVOjUqiEdjwreUx+04JV5pq2LHh0WK
XbZxP5PrYob+Fb7sAlKn2tPk8nfCixt3rHXs+GRA/F3HqRX84nL1oKpfjSHIT1az
l8UqTjw0lh6ao1J9X6Tr+jtAxfDl9G+XTXF4u9CNkB0ChMDC2CYAL1Y+XmLrBdWR
FixSmDSCNKYzp/x79Dm6dh8j5xTGAjInqIphVBk3/11esCoKHrX57+c7xSVzDcLx
7TxWo3FiAA1xzll9LFNmJ7bUzvheP66BJLy8Z+yJlbbncTsuShDTisGODA3+Ua7z
9jhrnHkX+KPCeMP09+ObGB4lFUrFqpsRPMD+pjKGq2Fi+BVuUUkh3b65ZPURXYC2
9fAaF4aCJHmZaFTyK3WEsvRjOu1s0nNVNAeqTrrJYkKWvETgd4iNWoD7z9NZYYu9
p62f3Qt0SC3JRbSOeySY6/1RJVHb/T9R4M/eM9se40z2y0cgo6jhaitrXMDHjzkp
tUiLMP4gLXQDMJxP2mtJc2ntCUk8Iw+nBFFQn6feIcSLYHiNMv7X87m0oDYkUP0K
1y+zZVUHK/et1OQTe1IKeFzz20uaHVoFFq9K+9are3XrFrXHSof2r61JcPEqBz3r
/qutbkD+ez2HX/plDirRoqY3ThYIivRwVM6tZ7fLeDIcPW7r6yUbNo9Pn0aaKIXw
8lHYD8ikVjTMRAsabCcPCfPrY2hj1aVt+jeZ6jH/BsS1zOboaN0YgGVDZvROrCNH
jqzuK+AP7g1HtifZSMYqhvM43rtYeiBa9aI9cxOj7lyZyAS4QdN1hrvNkUT1cDuW
fq0QinFQZVSKMMj+qxWqUM25MRlYlLpNwOXUQobZ8MKIlfK2CDOxPJ9/1nQzl5EX
+N253G7MWUtazqkYWFLNZ76qNfOEfTX5SdUc/cv1BCRUofl57jJ5UH3PyMN8/yak
4l7eh6Hkn10Xifilcc78mL5i7Y0Py4wHUfiVLnlbKNDBPWwVJgXB6O/hHwIP82pm
rtZXw1+aERtXNbXl7OK4xFHn17I5IjKGOAeaD/SjXtEj7WWjvvlNg3pXKt67MQwD
mx6D5IqH3hwD0HO6q9NjeATUwO2VtHme4Qj3ehke5R2+mRZnrIts/30Xi7xos6Rv
i7GcvGwsC4hVCGscfJa/NRq7hOjn8deMpkoAoeJk1hhcsf44ZvCu7rvAgk7WnaxO
A1Jztog9KtzbBWZG60m6s0u51dTiHoKJZNKbQp/2QEdTZUCJWMGbcZV/JTzTdbOF
Geyz3TNPt6M8ez/ZmzZduSECdcdGagDjgiN3pwHp1CxREU++1gU8NGFKpIJzISaP
2IntrfmrXhAKU2iiNiTzIlky0I47X9o1ejEK8HxnakxYUsGuuV6ye4NCeEKX0+FG
RCad/72hWpQS+ae6pkrQ+Ce1nSSpwwk0FYvC/fb2zSsBv9zrJIO4vx5YGPuxPgi9
orYkUdKGo9wSDIi6vbprJMUMs1fF3d1bszne+1E13RmzuWZd9XWs/8wyfxHaa7Uk
/bp2qUIbPyMHNlMUmr1FgnKzJmzB8AeGbNpWwx0GMArLOgxdx7B+dSF7TAuCz8Ht
q9zGIm2p7q4n6+ja/5Rvr4ODaDmu77ekdabkZzPPNuRe84WzGrvwqKh+oC7jtmij
fpd7HPFCkEwMx0Uo/Ou54e/LOFR8fGXEwqwuq1Jw0Ihqac5ijCvNQdCLHALhpWEj
7dU2JEKYwAdNxP32LZqRVJXWoaRKZAjD/xnsNPyn4/93FxRfEWGut8td3ojXXefb
9SprKPdJx6I9uuYs7OYYgVXxz/wAEJYXZVQX8ATf2FH+R4y0MHzHXrxn97ImlgkZ
h/OuswEogUHx/1QYxzVSxcYujlc9AyxezsAMeqD5iwEtWeOHOazFnn5z4maIJDGR
VfIBVM4Y0ntwbafC74HBS2v+h2lZpoMLqQlF8hw3udCyfJGLiwqLCeQ2yrLCvyay
CQ8IikPIBSVM2HwIMFQ8ylDN47FkUmIwmEDuGK8WhhZgrOv++MWNbDrF4gGL7NVS
7Hkm1uE5m0OFcJBxSzGbcpqEjTtkmTui1Nxrj61/VFPEAp9xxyk3LBc94gAxVm4W
Jh1jW3UlQnLyll49f3d5Z4w3LqbmjT54ZSBZ0hqv/hUS6HnMaKj0/UInztrHNXqi
MbaZJKXOkx1d2VVEIIFVPpUvEgW4vFrgcgd1lwU32kYMND1KSliGVFtmI+MdMiGZ
xPrbzLX5UeYPNiljvz7F/Z0/SEM+qfkVaz/6VmPbCM57LCpjEN5z/7axAWeD9eWV
oeqDfAB9GPDkjVNKe+V/NS4np+A9qvieBaOO7240e8OoWO94fby4RHnMuTXGPQkK
/r4LaezdOx42vI9DLmg1SIG7qGsIE5PcmDFyGqSlDv34gIK/RjydOZkvYVztskcx
06JmZOkuUTAQQvbV1CZIAZKCi/4L9jEn4NPYAQLhzpZvvh0xRzs/RaHdELXEdQFy
0mqQQOsQPpFe2Odgm9K8+HnS5IoicGObWWlHfJAizj+HB0ZJg/wfaGZJmnPBFqJW
8Nfp8RytB9WOfF8AGBh4BJi3NZO9h5ScEYmNsXkoJtHKgZHEPb65d4xh8FQ+28lY
s9hX3MmlHBcXfuf8q01nnk4mXnzHpLV+TWyqAIQKRW5lFv7So2RHjB8mDDrq6Qlh
djmLNVVzAOpDIVBHJujWMKrxof9xxj1IrXQrEAozLxqbJd3pbXBsjl0/XmAjRdiq
ztbqzViJc4dKzrxG4lBmnBbU1btLzolSfej+XxFmkCIeeQqRBurkkOhZAbPlnS2V
hn/TKELttUT4+3JcjZi+u8wbWHjqhVIcKekaviPirZ9FpJ58PgiCWH3KBbtGJSTN
BxvPi3tWcFLRrw1EM2ZhYc6pqaxEALiRSoV2/IKNEoxHMW+OjDKwU4zHQt38RCWi
xCGrgs8teflNbWqxblM8v7UatRtAcPfJA+a4zd9/mso=
`protect END_PROTECTED
