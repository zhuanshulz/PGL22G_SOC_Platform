`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAjhrsQly9cYcosJAtIHKckq5h8lOaur3X4iX3qvELNtdw2JTvbw1dS3VbJABqD7
/SNRXSk2xmyhUGRXrFvHHF8JwV5D5P0yhmTlCoZ5iXsA+WKi5ZyvVH35wuUcyUds
1mSDlJvE7thKIqmYuHuOAGkSeozw1wbfy9tyTBA398Rpl6btejs5MjBKPmrh3d6n
d6eaEeX8xZ1dKlTg/uamAq8qny66bDVdaFGFKSqyJSBl4w9SvTihfkJP+kdJ0wrd
lX0FaRilBtiQXI3rNJwV9bHlH8shMa0pEpDNXakt7k1FLcgzBlFacr69MezMtR/l
SoBsHPhipELS5a0PISMt+ds12JrE2i42WQa13gGWvDbiPRNQqFJJjcV3KxFtozQN
JejoKPBV7yD5YoJ3/NwYBbTRdjDKhdZk7xbm8uGYg1vNTooQ96TnXu2NaqAAotHX
KLHB10JuE15Ztyu1iFpmpYIQUWNznnlDrZhStFz1IkgaZsT4d/ZHBdFvey0rzAuj
1psJXJGZ/I9PfXYrg6DHYrYe0+zoxHxoXguztD6fxP6xeqHOBQPXwUpctUH4+Me5
w3xI+W7VUZxLqRoLHh+uOJ8VYsthxqO43EYU8+To9pphr2oVR6AxUe0P2T/0juqA
UlNhko9wmPuxlTqoP8xCxSOeaMoCpbVaY0nPawmTivGMD6C/72yH+7HU6hGubYYS
YuwaRE+xS+PAzaS7lP1vAatR6CnE+bXGryHOC8VFZPiEoyhC0o44zExvfpcMLxl5
oTNBSsHt1P5fYEoQXKybBTJwGqAC0aPiOBreMzWgMX4g+pXHH+ZA8SZ2wlT581ye
ZvSrIACb1DHFteA2j0h7Ew==
`protect END_PROTECTED
