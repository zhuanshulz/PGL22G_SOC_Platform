`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJDZKXoWYaxZNOEqhWxFX1tSBypLNklcFUM5EocstheQ+pcuy0m7RbQb3GQGGs9p
8bWJLwZtvkSpJ8kgLVNo5ufQqhf2JDtT5Ief72KDpbOTaXBhkt6bdmjh4AuWek4K
hyC0pW/BNChXfeOXv/rSFeGGe73Ro4t9f2Vh8AewTf5OkjFZOcSXd3VjLCYe0m77
Gicd5rt0y/uSMKCa4luuVQZ0+fCvsTG2J/WlqHAtzF2M/hh2W0PqLzhNbRHDZdvm
9TpwK510PPonMQOJ77XLhpot9edoUOdv6FEXIcsDjlbFTgn+KniQJEyLebXzxjrp
eag/Upl5cp/4QvGX0WGnr8Wmf2BJioa+PEQj0UNTr2z35Hup8gn50k7yJKe8FfeF
53qf/RzUwQyzE69bxYczKyHV9xCnq1t8n+moFk4yu9qXd4tl2W9BlHGyzeerYuWJ
otn9GzdYtHxfGIEL7TVDbDAX5dPgIDw5XlrxB9sAlTrA47+Xby8BwCtjzzkKGrk3
EpEf0N0xtqEo2liRPv0Ij/XBnAqV3K3O0ijRghir0V3leDTVQzlWIrSm7l1tUFJH
1ubh8AKiR8lfdY+guy70sfKnSwLJTZane+ukqybSp4HS32ANeNqP/T/DseJEenE9
hohVkucn8eWHHqeDwxXqzQ1KeqmelcYMu/Sv5RrTudEbZ83DQ1CgR+LjFJ8EPebN
IVnbOLu3fnjs/GTgN4KKi1O7lXr7+pJRqCI49R4ssnS1S7ONO18QDZ3Ll+L39y+e
iJjiiqYcLYwxPoijiEDB2xvRkUn3goe1oT4I8aR8q9Dfn4+gZJYbmYsVKhbC3aQo
oiY600c4C1+fRAui9gCdvJOn3+kiVZ2fWcSv74Y0C7JA0ETSeHFZWEJG+TxnxHgk
HG/FpOaiMRfe2D1LGH2ZkQsmXG82ahkc1CN4zfpaxJ0bX/1VNfuqx3gmpvFHvlXZ
HI5UQP+WptZaDczcyHvX3ps+EdzwCYneVefWxYyyA51v65bhwyMdXiGD1wFSnJgW
dXBU5BdWBDWmlfl0/aromFkksltonBvYXOrPLinq+HWKaT/NsVUrgUcY/5tdliCA
0V4euKi6Yb7Vs4wSzqi5KFqm2DI5Fw1wFfezrrm1cX2wVPOLdnR2wWGpv5gR6Q87
5rU7P+4GtSNvUrAXbUHrkPDGiyBdQcWctWk1+AvclF3Hp6Zo6WwnmyftoJhOMBDV
ujTHVQPa1oScS5IvFWlTENC/mrPVAK0wyje5PZS6C1xYlZrs8A+W39qe55PPgQxh
FrBgShHRebxfpwEYCvRuj4+3hGGBoKFcW4cjA2WrcSfAvb3me2Cgsg+Rt3ZcWfPR
ste5K54b8LF/+e4dLaM8kvd86k3+A9NTCFFPg61PUPzpcZqlhTz4hX5W0XEoxCZL
rcqnzAX9WQQhKKhSx3jVYzospknqJW/yZlK9RecuDo6DRsH/wqczJR7HS1UBjJGj
e1pldG+c6ktOAn3H5FL55uok5SkpxsthZg4eszvdxPefCN+ZXw5XFhaUm9u6OljM
RKCyN028TRFq7pJLufCBynibRIivv7QdWlmmIbZsgwc92XeFoPP6bnlY9PaSFNnX
q3sVVDI9VqDXbEDqsRMav6IlTTD1OWp4upymKYacut7PN+7SzBqL1iYgT8EcK0Ar
0ip3d5ecmEao3TfSlNvUjEyvAFNQi/yGXLQmcrGxbRNPUvlgBHlOj1diTgzGNa83
cYNeqpdg7RxT9c504oqmy909wajQ6c39TzwJKUHuwhClvTTu7DmvdAyVQrGchS6L
CR1l/22Ifb2CgJruVqAznLlINkMpOt+XIuM+WNReG0l4y1L/4gUq3GX+3JuhIlhF
QwCHcuG8X2jCC2mkOpm21J4oCAIwH5DvHPWHZaLhhNvZ60U9zciBPAR+29/T8Mwh
aX/mZxXRVbunyZ7yvv5nVLPg9kEM+t/2ieaBStXQrfKYlD72FWJsFMDkjbKaF5UG
E5vu5mps5l/A8V35xQfOU7pTX71kQi4tahHfCAp6ChpdsfH1FFGbsvqSBr3b9/WC
Y5/H83a36V/MhQCmhNWTfc3w87fG1u1hP+sAl+zQ0OJncsi1Mb//UiqcX0j3KXM+
rIzCpV6K5SLwZHptK4+zUq3HiuThe7s3h//fQAw3xui+VH2fTZE9sGHHa4eOnFMO
yfKqSfvG+PvNS4qBYbnxLvWhUsha3Jlwuu7NHTr8hgpnZeCKWyp9+rijNZ0ltyFi
nFgRY4VyFLH4BLNGVIYid1Xx4zekvGNFLdTuno3TkaPPWKQIIcMHjq8n+9SPWCja
ReKSYEgEYkZZXPfxpau24H+c4Ua6zj/Vodd2qlUgyjwsD8jbXxOF9D75+2R4sEXs
PuzQ3hZ8+hzlpuzf7XI8331i3uVaH5Q4jzce3tVie4MveYIKnAk6oCqmuKUoCS6y
bjrXgHJhs67BDgXLez4stPkRX24ZylfVkI2G8lwNzS1rKwjikKWpLFxguthWkmeF
Eh+ADg2lpctpbEflpRy2UEwDqyaml1/rB5gesjVxE/zs1IdJb2PLu+LN59O0Nqbt
QY1HGIz/68JIp0YSzrapcqhesCYAqVnqygst3TzICI84SYETtq0PaBIAipGUt3Zm
0Sa4ND/SupFgnk+qrcwbKWuQk1s2oDK6OE+qxKA0vVVLJDNbvEV5qjPki3CbPTt+
vO+Ftm5KShh3kZ/nVF2OIbRIeOyeEhuoCsjeecLeeRt13QW3O2LgmzblWU+4Nn6l
Koa0qnU/UGLlV7TDPMMQffw91kOxsR/XJDURqpze8/15lt4Bl7Jx9FcuPUKejoXw
IApWX+C5W51IKhRrsqbuw5lPY7Avi1YvrrUl5xw6lfGBz1R7w8d1jSZtRPpRUaGM
m1yDbsq+5+sW49rlJxaWZc85WOc/DdrCFPNL4xNuoNhc7UxqU5m0jP335Wa1VmSw
0//HPluc88lBPJsgs7dB2qlAFINM0fhvpkPfDCE/CJjkc8HuPiCu8S+US4/pyKo+
3VD4Dibm4fAlcy9nzq5G2JIt+99JRRsCUOUnDsjrwgYdJnYOCVvdSplVj3FSlhAD
VHgEw+3OMsp4mjbO5gUDLZSVmgdGeCpKD4KFhHCojNEMI12ambWqK9v4uE4OKBtS
bNim3elnJd+8MS9vLh7p5VDDaVleUhgtKCjZpHWrfyHH+tJyvvf0Ckp+TaBKPcnh
sZ6TsbcJ7r2377iimNJxFBysoR9jl23pMufr0Hy5PgtWPHqx/b8HdJZCLFVYzHoi
RHPA7e5YAEoXRb5WxUDCxVi1eaMnDYnKp3Uxpi8TGbpyuE0rYbq8TjP9b+Aesxgd
dfz6NeTAIy9WYfolyi97LFcFujDlcRw5FDfUvrA1EjTE/lhUazQrmcIPYgdnxoZV
Aw7nAe7cwK6NUW8CDqEIIWvwb4IU09su3vEX5/EGvNS7MKCNzQu0CJtX6u+SOROr
VUUjn8mHG/h99ADXFCuXP3yXD4fM6WC4pSzJnNFSmFsyQSFgprqUsjidUEP7VGpu
Fp+FHmlHJyMt8eGauSXXEVuxn7HFjHtVTP7To8LWe5w3sQv4uNo03h2uWBGlyt8V
mUOIEklUvGSSVzghXig5LAYbOm9bWwE67jZH/MFGt5RcM4V2bFSE/WIs3UzUGHSr
B8FR5RsTyn2YaNCh/UGUlDF1CmdcRh4HXZklxWBisQdpO/KbYKP5TTaLNSazVI7J
vhF7qAcBWjlhA8k1cOEXvN9gyslSZI+CYL5Ogc3Mi1HfUSTcU583Dx9Qp2c5V2rg
kAX0opN+H5MhwMA49MQjdubm9KRddzNZQ+aXma5fUU6oE+Am0GTrh+d35B//n30W
gMLth3lETwAcxe95OM9P9IryuL1XNs8CkRphFWd7i7YIC0ZY78ExjtrAfNmjOKsq
ZTApCphbN04avCn9vE/GwD2QCa/IdIe5GqhJoQ2umPsf3QcMqCPoiASOeNLCaLpu
OFC6Aran0NgFTUWwoZbTa9/4ms/OgHpJBC9dIvOTjoXPYxg/qaeVrSZ21yLWZfyB
KbqHBVr8H7SDOkl25yTTpRI3iLezESHhB7zq2qqZ0fOYylF3X6BFKeGXeiRZvtGT
NfIlPyoTCmTaToF3sRCHps6oPskQWTb7AQIOmkWtog5vmKLBPsiKXQHff5ELbelL
XrROXCBDtg5/1R4tIfK8Wib+m8M/6s+3PtQvQLX/8TEUkqSBI2JRLb8tIch2Ed6G
MBLRc9jzL+mM3MlCOuyIphBdzNG5P18KMzoNPaAGstv0NMYwpdA/UvGBG/bpibM4
bINcnsi32w4cHJM3F6V9yhkqPnXKglLXEs4kKGLPvp8ZXHwtI7B4W6ZHOr7Fcb6F
zUVAVVYgcVMmVKuxPVr0npE7H7clLePhrFyU7cYmerNSizBcpE6D3HkLoj+Vgxxt
mjMUPuvWoVdMXkeb83eDqRTD1gRkUJF88qvBSnoThQYaShwfp3yIoBG3Z697iWYj
wnMecdN01oIx6WuBgQTNiOW4YLHOIwFwLTwfeIAke9OHj5cy1woYM8nqJ+sXew5Z
WM1mKqJwBziSqdB9Ash3NkLc5G6hsngys3WOtIUtGwJHu1o5gdcpLqjxF/hW8WA4
cBb/NOawl+QSDtio3M+Ce+JcNnSRD2elmENCtFLugj7/+rENGEQncH411+iW4M2V
489Ri6798OSGQA9OXuLRkwVwhP5V6bgkJMsXX71hEQu49bdU2qRVdQmJAWzXdvDH
edlA6NhgH8gHLPmMNokJk0pP/W+tiTpAB0deFxlWCNiykUSbAmWGTOX5SOyJKbq9
ggxNE6NHn4yMKCzeLHqkHnUEnOTK87SMJ5sjWkSLvYoUN1uhpNo1m5wGcE36qLIQ
wIIMNZvy4oehMYg19qrIbcA/46Ltc8isvPujt/mql22DDTtBei/1rklph8fEsZHC
y+wOZYFr8+AJGb2jjeD8RgGw+QOK1aUY9kZhP5zxYIeet2LI0WMktHekD2H05bnL
teNiRVdW/92k+RPvcAaZ1OMFzaI8IHGoL7XXpS/QIW7fK9QtwirMpEdCU9fzz+2U
V803sHIOyNY4z1rgUFr24B1LeXIEZbWsG9BX9JKFb7JMQiw5bm3fmNcECmw0vosr
zvlAtrSlx9xWg0pixLkab+Epz0oTZCxLlZeT2GoGf39QgRmSXTk8evQlk+zlDYri
CPr1+rCSCcw6G4++iFk95965p5KOssCx2iDDObRvFj7eTwmDIEsEaLlHwBRMWWnx
l63jSDNkIdlwj2g/tBx2TUexOzetBj8K4S71btK7QqbxHIB2c4yN8s5pWtlVt++6
z8sE2FGTNr66vOJrFjL/5dnpMjZScWTUO2DhXLfHI8EIkCDTfT3kwf5yCpi+O0fQ
ss1U5Z+SeKUdkcqBMECqw54u0vaZBoZawYHxMXWYzdx9L0K/W8QrNlSzmg7FJL1p
Fmg+afPXSCvM8Ev0zi9uGKZ5ALM5ddvFuBMD6zOcCpVU+/bTzDbHSe2cyQrmASAQ
HTYsgSlUED5NUO4fK83Nd3XOpLNw2qkyusvBbpjUpB+mBbi0Dr+XihNi83S8cRWJ
36AuAHdhMp9GHBIaldFyxRptl+48TLeoMK6jxikaUZsXnGcKtulXia+1rUh8TdVq
7AkzHGRAIvdwS2r6GrJDd4aOfJ8GAyUghNHwnzU6eLYuQ5toTrh5YwBMVXUxHD9V
W2NN5F0y2r5nsL1uuVtc5y7IqTdyU3atppuhrx3jU9ypw5JPsV+HOAtHsnjI2qL8
qcuTHKtjQcnQi+IfDQcZoyaR1auVAYhbmdNucxD7a/cYaEGYWoLrgKtpMZ71USRi
QGpomLxeO16cTPCiOm0vKE6mmpQDT/RNAYXO+hxW+ZITYJ+EV1ckNgxBzGUmOmkc
T7OCrsFgy/vqGGo9hnuPyHI3NwjO3oYYg0ItMJlr4ck=
`protect END_PROTECTED
