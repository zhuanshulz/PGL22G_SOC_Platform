`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Mqtm1xxLEwzTK4ugkhswWGs/aNzST0xrIDrTec8+JyBF6/Tc/bw4DZzgGNTH/zc
sC+dlcWJKE8qka7fmqYF2s4b4Ot7m04wkR0Tp0AxJ2fIM0BTQmQKVd+vW8rfsSB6
RczCcad/qlwGqGtj8cMpoN5+FL2WdCqj8/0+Wvn1MdNkj9bMV9Wvgx1BGDYEUfHQ
RjydZ/kzTiUpfMSGcXGIAB6ukUsbwhylESQCf3C0eaqCAj8PAZLHu+EhGSYA7UcZ
s9Dd6LP0Why4uRYX41uA8dxMmx1f1z7q/MAXuetWLm2GPId3Z7s1Xjwf7pxDl5gW
7mBpurGdPtp5V4HdWj32nWsEG1nlWUyBDDBjgmilMwR8u8Cjf/+ZhbkX4PwOZtLb
bOAchE19RxiO8tvzRTtaz2nsbOlZS51dKVAen+1LNLepyrMQnF/fUk3RfL8ARBPM
HtUSOixDUk9w51C7gotOmPgDx9WzdX+jC9O9Pk762xiSEXOOi45jzhMKPLaqEBj7
cC3vj5HtzLJvMx4fT9jyTQAV1PbIQyzKS9tJ7BF5CcV04t2iBzqVj8gfClbri5la
/EIP+c87IT5DaVLMwgk72sgKz/l8+FyU0TjO52jWKCNO7/y2hZx7VXmsj+cnhQtW
gxyJrMuMY/incv7u80h2gWA2XqZKBRxuSzmMffkW7b+nHVOv+bZcbBFGNQMqcCkq
/6b4AEEUCsxmhjn1qQ+2iaqNKFKkHE+305WLyVC+mMPu2DbJn9gfCdr0x1Gssqv4
qpy5eLSCa0zQgESBd+tcSrrXEgxCLdsrhp8licoU0Jw5OBK84SFFAdDwN1VnZ3I5
w37ynwkoJDj7mdcHDDOeGdeQJ2PRCA0CJQC++Wd1435gLNaRcSk4VNW+Bae+2XmO
uOZTzsn+8lwsjoqXzVLntw504049yY0KWSHKhZOi/S8xhCXahYx2c9DSb2Y69BdL
rZ4EQ1i++I+rP/Oe3BOA3miT7GX3DEVOMsl9bDn6PUl9R+VIfCTOrcQI6lzvr2P1
yMFdYFRG6ULkgtFnl7fd//dlbMuohG2apFK69A5dxcyac3EJWIhl/pjiEUE4bgWN
JgamkjwhpheYEtl9btPX39nkaGlOsowjaCJTlU+5GCLomKw+R4px2HBiVlUbBWyX
UA9eSjZrR/iFAHTrEG7nEKPrUTCNEQpAVX3wDz5WKGFzn/sXj2OAC/rdwf+4uTrO
0UJIGYYRgtzt9EJ2w+wsBrUNqbdsYOomxcos3gy/iUPVFgJG894xVg0152hatAb0
zXwUID8VSckuBfNMGZDWrjWD1M+Tj+MlqukUAhjYisevhIQZFnqkaF/jDkdzPQ+X
MqlLL+P6sv1Folcg1Rkqk1vOhoMskENp6SPzQ63Vkqy8a1wV1LO2yxFg73SsxnkJ
D1q2F15d12N0SFHAW5gkt4rFix45HEN9itojNST9FBD4ongWHZlPI8CvYNx+p1C9
a1Ugw7Z4JfnwyXguLCKLxJNvi56zBPVe4lZegetZIuKs6g7/wdTZD5DFBJbPodG6
LA3lYmfqtdYlJZSOR8fZ6pwuqEXsLedJdCVRczgX4q51tVMPZmywHhPNXA5AkQGD
SRnPULeBDmh5z+ozeXxIsUl+fpEt3ZOO0/kAXYs6SEgvn9/wc4yowkFTS59wGny0
VrZaNgO3g9Hle8JOyQ+WHlbk3gUJTjRDAsr44F16u/UHLJBlMeI7P4NskP5xy+kb
qJUN7a6azszP7gBGlOBIWuFKhfTaHeBljbQZJCInValNnhhtbkeqd+gQ+XEB8N9p
Yh/Pr6zeK/XS8SwtlIdVJKFImClR/kAaJ+D0BrNkxVAvsWTYcyXqfh3n9eGntGzs
bBQ/N7clUoTqJcoHrkC2yMCRLOiouKMeqDBpUfsZOaUAk/8h0CIoxwCmTeX0kpQB
LfrK3FOIbv28+HPIPPaaOc5cymmO5OYL7LK3WMJqIvleiD3JlbShQm5LsKLuh7n2
bEGhiBPT4gP2WTLiEP5SOh/EdGF/H1tOAwA2vZBrx82et7911g1znM5fQMKQ6S9f
TWUDU2S0b+Xk/2J6M7GHNCJGu1JfixjwcWggQ7hJy4ZoPBf7s406wcSamFL6vmp/
oD/EbcV3kc7tGLK/TJ+GLPyVprgTu2lyUQMB9fYme6ygk1bE4EXTvcwbT3wiA1lD
OcW23U6PcvIGR9kY52B2DXveo2inrRU30nsWrysAjZLkt9lQLoQDt0auBfMzaMGg
QLjd7NSxMN1j2a8VSPPNSEPmU0bDhxLvbF8xxnMxSCSgGvmJQZFmCfNhtVDmByzQ
fN/CQAQwntsDWEF0Y50OB6tMYmGqsh2654f44o6hJn8lfQI0OYwI4yu6HuGA05pF
LyF/zR1gyg7XYZMQM68N4jlR+oBjSNmSqlAdXdzQKvDyM2hmGfijdHehqQYLVDDj
sQj0dZXaUlS3Hv1ZktCmknNVm0jL5n37u40sFSUfs7NGnzIlUnusv9OQruZo9P9i
vCBqa0+5ly7Q6sxhe6M6/E/llc5t+nYNlvATNH0qMKVEdLKZHbB7Kz8TaYsn6e05
lAuYoHn64V+f6idYVHRhYxk29lNc/YJb9D24UY1VPiGTj5d2jt0Cr8wo0OY5XftW
tS91IF6pgM7ZrHGtyjfdhmXS9VYKyGT0kAJVyYLSYlMlFXmt2K1cCimUqYWTLRRk
HXfqQGCyUaUyclYk5iXMyLdkOQqpdL5rvR0e/qyP0tzvCYZGK/TgXn0j+qh82dmT
yF0SWgrLKvIc8ya+ywCOtQ==
`protect END_PROTECTED
