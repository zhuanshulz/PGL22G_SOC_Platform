`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXr0mPrDoaViZuluaMDI5HtGQwfxoSETGjalq4gKRt9GxDDDhXL94UoYMWfrEC8k
3BmS0mPYYV/FFE2x5GIOEY2mWOQUEBiFRgq+s6dVEGb7c8pR52fQa507hnBaLP0M
wcntgmg12+rQ9cJo0QFFwryrl9jRivDDcSwpmXqQtfj0LhtaATBwED3APrMZZ5u0
CofolN6903zsOCyMxqjFHzaSyE5D/FtbzSTfkmaZuslCZGE331vhPsLAzX6WTU8/
mZE4bMS65fRC8DUIL0/PmHceBKEiaq+f0tOp38OzWOxz2cCV8yf25r6qFyB1kohY
GDVWkyVd40RN/YbnKW8fLvhyuk+9aKBgISUwO1+5T/9hXxDBrYyFSEXTWSsFiarS
hNFcBAODu4s54+EFtfO7yoIgZWJdHfzJZfPpUlMRta0+HQmuFijVQMlLL8C1hz2M
S1uR5R6Blm0BH2xqLNAi9LUKLZEVdSr8m1a/TT7v+qL7+6JGP9QYZlaq1DdttfbY
VzSv5gqJpBP+wP3G6u0NcASUPb0jUQfRmJ1XubQ2hDEgLkQT/HqJAQpWgyfB7AVX
ibdEaxKl6Ms/vjpBDWR6Fv2Z6oxMuyFBaGTcLlpUcO3xPs0FhWPHFQiwzez/fPA6
fFt6PAtpCz79/6FDKX8wwAl+HX6gnFlPNqdAqmXAGhS7WvIQVOnt9eDLrRMst827
HssAxcFqvscAX8LZeFXRWV4/ky6gu1P7X/XpBEOIns4h5LRjA4xP96Hnqupy4ViV
uEGoUhZL+iIlFXAgQakt92lg7B8uRzelAABlVBZ5lqPW+56bpPbm4VbtGLncjdRF
nNyDLKiLwP9h/NqTqjCCIXWbkwGnaJ7pNfd9Z+C97sgPE6VECSeqKF0CShkh/d4l
yBTaRLrbBRgBcKGr/VePXM9ca0mPsNStNS2wM8Jz2PdwTZqqHNL3eAn52Q5mv8uX
veaMrmPOeREpXxJPNb5vdvq0mza1PKmn03t2eHx6qHPjgX7TT7J86MO+02th3YeU
UigNbile/5qNPUJNnPSEtK1KDKvtwSq4Yl/kXpbpKyN+Lej33UGQmNtAh6yspmA0
W6rmO1OoEKwFgETR6eeup1YDfMUNkqwxuytqEtRRSSrnxtUpSPD8QgBX0mq5Iuai
Xfg47W+3tWnuh0pkEEeCLUjPKxjh3C29YLAq0PAfQZ3vjSGpvLnJqF434868MYen
9CXFK+vCFVWFTR/4cDO2WIyZcGupjb6hdBGefbQ4oq33N9RgppJsOidv5jM6mkIW
wH8OBvBWuBS50Hv6B2dunXUiHWgXhhYfSAEIN0sX5Gx2g2ziTGthtCDqmF0ussjB
pCRPq6DxHKl674mclrDyOY0gjzKHzeHQLnIs+l35QkGfipGZnL9sITErGQgr6ozS
sEQm9rIwmDFlE6nLfHwnyeBkFEIlt75UL765PVCU/LpVGsVKIU0xc7ljXBLLnt9V
Irp1xxA9oKDf1e9LN0JHAlLU+7FEfL0mPD5B3LCoLYzSKzFQ2C1g/dsT+lURLrjc
U8AsVa8T9aJ5vkG4W87de2OPiLbbQxyCdLsGBXCDEUc7CP10ib5LqCUy0PeINpL5
2Uu/+okNK9+IhwiXDpQNcGr2kmJJXw2LkRi9MrMDrE93CB0n3O3JOEOoCj/YfGu7
bH6CLljYyaElUc+HM97z1+p4cj719YXzgu0ZmKh5IXwoG1mj63iRYlF/1vPxOoWc
artsVPyD9EVhIRU5smezDQcTI2gPkkfWtEKTWKdd52708fgWdqQdmxGVTeXNP4NY
6fzH5hWfVe+Xc778xChyAlfZGeL8aK3YR+slybqetvnG26FWaWmkML4gG+8gG+Zq
Sh6Ydori0xhAHlW4xLR0x4o41YnRKbG0WI3vNL2gjGQgjIRtFaYGSW7EsbytbzYl
G7F03mFrd/yhNWDtQiz4zbzuYEpHOjjOry2Dp71KLe2hsQO5VVp3B0qdWHD2iJb9
oBUs5PW5pxNKw8MpG3eJD6V/7dIXZF18alUq0JN1k8GSaIgzfKLdv3gmCc4bKRRT
Hl87O6oZaCyUcpGy46nDdtviBRd0f5vFwW0ZKVLm8t+eVEm80Z+1j2FRryflyPXR
b0yMn/JttECZd+u3ey4ptKFvwhgQuB+ZmAPx9VyleOiBz58w0EhMp0xAUq5syL53
/lwAWlW8+a1DprcMOw/El2RRZUhc2ae9NUN9Lze//5ajb/wynaEAWCXbuPTe3I87
KvV9yOyZwZDRoL6VPPV7UHVKz/6S+aU5KZIslZHJ2VuVn8kAK0jaEJBZaAESt7Ue
B/rEAeJDnZU1Q4AjkMhkcU/Hjkef+hQ13XOpp2Q9qFgnSel2y4CSBfjqRpzY/UOA
eFrUGgooJICDCHSHsgpkbYBHACCKRlrMUjUbWuXZ6o6s+fN10AnxMuC7Od4ATyxz
+GMZUk58zTu/YYtD2p/SxYhZ2cPXsNbsd7pwsDVcXVd+ht2ffJiaqfS7/wEEuJEa
FCka2xTScgtzV7pD8utb4BwpGagOxPNJ3WY+F7XqtTAadRD+kUSMUE06uqGt5O7z
PJ8VG5Ow/gjlf3sbs5f823ltOkD4UM3sJo279bybQt4DBQVZdTZadmC/thwqv5cT
uME4hQYZb/cg7h9Pn/eZUDUXaNOWWELqfCUad6yxPqvAESoo3tt54h+rFG95Cr/f
RW+zhto7SpQysJ92QOzrRlYNv4k/eOeww+60Uys8F3GH3A1DqpmMzMZlIRzTYhds
Yxfftgk7s5icYMzHmecOQylqYOew4ujZlbUCV5o1lFHoiaX4M4MET0LHSG280TZ0
wfQEJ3UCew2L9fa/RcbwYSxdz2gaOMnWwAwHe+KA70pK1TetmlLCchHW2lQvemo/
P3+8/SkV6hgRVkz6rEcKLAuTeAs8doAgfNFfjM03A9l9/IgNboRHKqdb9K8ancN2
D0+QtDkKVAUFMqu5ksCtUW35oElRFoAkS3+VL9sdq5V+Wv57H4qgleV8kMGBR7iG
moLE/y8KkZ+jJnQIGqiAJVVU6leHfAeldAsFB1DUl7LoxsjbnJq1R1pqecs4IMTl
m99+YwQ00JrufJvKA0269njtVS0BKDptheqI63COfjP7m8pReqIn/fYl45CJ3ZvC
b2tsfX0+v5PhPfpoyXbs2goO8EN4irgTX6v9OQZlMMjqolq0cnj8JkyTGfUnHmNj
eAw+qOIIDxF1Bqj6Xxgo8YrhUKI1cAUkCm4BJNlHCgW9lHdagqWe1g/StdO9C7I+
vzdnmPT44YtOjg1QKMWHcoivOh+SQoeRL1ItbVvXjTq0iKH/P6U17OjMbspZczSG
W75/Ew+YReOzG+NVxw3zw3eRliyWFLurNenlQQiMKW06OqnWLTDzVB0vO0HBF3to
BGPlba1WvWqmfDAJ1bql3cHxCl17pR7lIaxfWcQulAHseVkMflxaBlLZoavAciTE
pRgdNqMdRh2TcrH7/c/y95U424luOH9Bu3xdwT/9iGvEoeH7ZxPAY/a8wSPx1uB7
fYSxCfHefp7yqC+V934cFlS4xS+Yom46kIMn7oiQj5alXPtEFhbfD9iVZf7iUM7n
Si5RxnSFgvhqKNWJ1d1LuGCU2uF3oh1H4i2QpuHKKpZTj7oycPnsa4Ry2tKjilDX
LIrs150CQkc1lzX8JvQB8DrB8UUfdwOBSV1gHdAXtVZ5+P5YTuDcqmiBK4aHrorp
e07vWzi4LhVqdgQfHRaInW4X4o4Wp7M1Jwxt8sB9NL7rybl/LBKIEGVCaS8AHzbq
i5WtYon4LEl5b9aR6J0Yc+amujKWtD47NZiqR70r/rSeAI07wWrhL4Sp9eFrq0bA
CnV2JEs1ykY4vdIj0nwwbL+JhmB0vEhLYQYTgRaakxLN5RbjqvcDXRZSPVFRMRNv
iGpaXbPTE8Zklwj1JoDsscyL3dpy1An840CHDA9hrKZKziZMIImavKHHzfETuUYk
+c2YFnIuavI3W1XpJ6JfpHoL1/A7usePpAJuGZlOPt9AzYbe7Z8oVY97u1MS/NBM
3ExsLP9PiaM3c0bVtJzCJu30E1T+bSlhfY1a1+0nWrk=
`protect END_PROTECTED
