`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJfq3+hjsaNrC0PoFmS327B2tMAeZC0kO2Qi0dGPtfh39J9idBiTPnnsLSEA0YUP
OI3qXyntEk4ZGCE97LsK7SB8NsswpRBpC7WNoSlfL6JGaJdG0yed9GzyImZapbRM
lHNf1vaahIlu6hpKnfdFj4ViSLmVtYB3DYB+yMY2dVQAl/5xoqdGhWP2mAhbckKp
74v0AnE3S1mnJHRuuCNtCdeb5z+N/PyVoXJKVtb7O3nCF7oesEt2f3L71K7Arrs5
1htl50Odbhv/ZrhJ2goHpuAP999mfj+Vu3TCJp7H82cUCGqqmqr+Q9MO9czm7jVd
Ob4QcKy2dpOHIVnEtGITR1mDnC/W43KP3DtI9HDNtvkzI41s2NtfgR9kYTV/3b5O
E0wiTa+K8K7Xx/C2rUyEW8bAkUKMp/hybh+IvOQpZMKLDZKd2pvxP9zCaKa0pvIh
/Zll8MvE1Sh7DWkmsKJLnces30HixL3z1n2V3RMA2I+XE65Cd7STXugDQOmJoud2
vfFlWCu9Tq1mBERJjURfbRyw2ctZYRlalPLIdzWppoJQ78g9vowKweBev2qSFcAM
M+HBaEacNV9yz6byCWtmDmQQpfpsyDlOcXykfXO+FqcL7UH/qnXxAd260xYrFHZp
U4k8QSVQbDolDX/cYrrmeNU98gWCVLlSM3PV8ed9Yecfrh8/nHBkx4B4knvw6VzI
XzPg/9jqM6zzkqXr6TbLaLCsKyrPPGRThT7kG8vEEz6XO8BuUm+yL6/QyfzsUoT2
QVutZM+/plmXpPHkDSr21YsUm2WnfHXuk3RxzWe53bO9cFlQsLvgS+Qh+bq67O3A
STjf8W4a4g83aMBjyWuMwUU2Wg74GWKFG6eB3EjWoV8voemkJ9zg+nDFD/YW1u22
2Gtu92rD43buvhtHThk9tOOE5TUcV4LiYW6JlQ+CiWwKx2GIi5s4GDIIdjNC1uGT
yYYDGZaTdbB/52t4YeP0j9/09TRyguDgGPxYkV3jSC2qy2NdbuzMl3hcj2X7ePQp
pMKxqE4E0bxN+7Nz2rrI2S6PSf0YXZJGmi/davD2CD2cK177B9wuCDCNfJv17QG9
UwLMgGnxhYqaQDBf9EslS95LuLfEgHl69sGHrVD3sySBRerc6wdixfhSyIBCv2FK
pjPn7eJS7DVv3hWHIAskH06+1pclLR/CgMLGrIq4VToHMCMeyoqSJ/yw5cgaQLM9
3zzW4N5gZ4PK5u03ZScHkU+Bd8ARIiEaQpQrg14s+y+yo70fk1ELzqa4qX0PitV8
8H5RPQk3jl3cWhk51yCzmGLED9C/COAfOAKJVZc1YplJDmQk7J+7URMpvr96Ayyp
ynTlW+a8EqRLOonVsHB5jETwJqVOzHO4yD00bQd+Rg4McxZKqw3fDqnrXbRwsKF5
B9uEyYcYqLbvUXRHXwGdPfNCF3dIvK21wunbIX00gGuDnLqQpLvBf4WJAZw/oKuk
4zD2OXi+OGnxpRfDGYCJpklgH2v9Cu9oVOHKWRhqf4dsG2hhh8NpQm+QFNZMKxx4
/WSy8wy2g28icwnMCsPEB08kbV1iQb+JECBfGpgYCjUkZ16FI09c3zzu7bP7nnXK
yiDxbV3ZjugBAW8sZokL8bxXdahfX336LaE2a46FxagKJffm/3ItfWc2TTXHxwOe
B2G7rHnVV4e17VcqCifSOIiBjP0bFnpLdaXmjZHWnEasq0w7SEUc18BhCI5QRRwJ
hjo/60yuAl3tMcmlwrPg8g==
`protect END_PROTECTED
