`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFD6ny8P35tngq/QxGL52+Ll1ubo40RXTGydBCkfUtAQLjiO/LB73f1BJgoixqlr
eihKwVacHNpWLEMDhZgHdOpN2hc5EJhANrYm+iEiv3NzZXw4L3AjSNNxAGnd+Lbd
BK2bny+Y/wEtjvIrnPaxt1NFC+c93coSl3idlUAUSUYUDEhi3x8Bn3anizzo4g65
fwqrbgleBgd2iyyi2FeSVO26Xn9h5Zhv0zfhiAXiUgLivXWuXA9HyisX+B1FwN2J
eC3Z/vsntbrbRNl2ZR2/ILPB9o/CtiSSXzUP2JbpafEaX35EUiCIqc4UrE/c3a3d
OQgPIHwcP+0k7JPWLvvMjg==
`protect END_PROTECTED
