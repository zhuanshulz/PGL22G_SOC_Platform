`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/S0bqRiReGkGa6SUC0P8KibEdx5MwS+QUfjvkzt3mTOQ45LVlGtP17gI6SoAmaN
4q1ePrwdkcSWe2PdOBy/fqmdvMT6XuWXqGT3Fe/NgS/74L/vuDNbzJLvsv644vX1
XAyw7EOQ0NZRuFGQhuLHkcwHtK58lfSgLONQvaIQJxRo6pFOBjdVMWlRWOH+uuqw
IHGXey3Uqqc0fJn33ya8jmvNI5C+iRQl/uhclQDNRS4qZDr9aJvzS5pl75kjP0mY
NEDOaWe7J7q/uj2biUL4+Ox/PFdxBituuMUGxiAzXDDTLHLK99ceWQB7ptODCBZu
qxhGm61S7LK9sZcz68tKB7yRT1z/Go1TJF8oXJU0UIyrMzsJVC44wjlr0oiXZWX8
3RciIq/qYRKZY9zezvc2cVrE6IeoZpnfqQT2QupkXHLxEPUYhgqOCshJ8x3Arj5C
uN7kVI0RUcUUE2xvFBkXomd8cY7uvNExBKiGtbrfCrGFfvaWHdDXn6109IewuPPU
VUqa5dRj828s4wqe9KKJDlULgzckwaXGc+87Zg/FfyfMHe2xqlKMbepb6Q3Prp1s
`protect END_PROTECTED
