`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzcSArCGwcuFpDVE10XRK/J46jHeZ58v2Cgt7YA5q7BYTYYsGAhWihK7Y1p1pyKV
swBU0vBJ9taiKrGdbfGMs/RHFm+TiQqJiBT+HhSnfu2HuCjBpSYgRAHYXto1On8Q
tvHhHrHZpGsfmb5SYAge6V5bHpRbEc03zx2aug7KN0pRIExsaw9ZbkEtSNfM43Zi
TBxhl+3p8GfuusM0gzWKWm0FESL9P7mtdchcALIe6JSidTHl09Vip2Kc/7OeUjW1
qRrERcaIo57dYFFBhEj831hEoFEKT0g19p3CKLyHmjTMuTNjBh8VSWOPpLZI5AnR
gLYt/0pH4LRJmJQI9Zs2wrTyvoJ9Rpr0/+wTUtMNJ30E4B48pe5PaiTSek7gwU9o
laCtPlLFIGet7zEd9VsxQS+DtSpjVIatCjc2VIrbd5ZUoSv0AoEaKmGrOB9mL/nu
nws+AckCpgRI4hDlaL9BOPIhEPjUcfrWEy8gR8WuND4K0R74Rm03d/bmOd9H+YbU
KcjwBPkVTAJttYumMsANSTmrWUi2JxhJmckDmXUVrUYv3vaYBn2tCbNRyFPHz2sX
pPxz5LVTjhAYVqNya0EiiXJ8BY6dhaYvuSWc2Xa0NHepJX4iYqGG97NQbiCK4/1p
tOGUa6tPIMHjGd7sOi8COg==
`protect END_PROTECTED
