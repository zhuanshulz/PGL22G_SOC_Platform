`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
brqLF35C+C2+ihNy5BU7xRNlogF29ooZWbACX70bXOcZOu4NNWM2hBhAV9L9WPxe
G7/mu4d6BahdGczW1redmaTA1VhJ1LfdQ1MmYKQle4Xn5xGMCjKfUCzefoi/jLpo
gcSaBEDHDgQB1/zbupm9qSPz2TRxe/or6ebTEJ5CdxESXp0UD4lXuE72qI+q6PQY
reuo+OT+imVmhIwsZtesc3EzLjXraM+nOE2o0Dt4TOIkLzTA8ppR9FOiQf8sMI/W
na5qytnYrzkV1V33IvN80b/JOMWO8gSgSJtI05gCLGZwccjPA72rDmVEylEaKxPd
Pd7/6UyRqX6QsMt23rsHzUx7ZfnmhWJFUYwMFVzV9nRmDU6RFAbf9JEUkKT7EFuA
QGD6Z6fZH/6UpSLi/fLn0T5new6x6plIWKGlFeLYnD+uDPIpAMxDu/YyB7TZfZkn
4ebnIr1WqMHkSPqjrRj1mCnmxjFSjW0vKv2odXeknHYNGGDeR/1yXtJrg6JfhKks
xzHpBq3UlLjuDtX6JA2A+Xan5OG6spHSQf25TcShWI67z0VgD15ox7u+Ggze0B1R
QIYuT2obEo6jgp5zqOO4pw==
`protect END_PROTECTED
