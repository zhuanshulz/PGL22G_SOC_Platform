`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZT7+LIAeSpD3c06rfWeUBktIolMMgSANlBZQWuQmdTlTYaDGmznBvYcYWquGmnf8
cLqVU0/m6OBbAd7L1shclo1piy8I63VRn8ZbuLnM8Yl5oRBH/6A8zPZ2PjbHW9eQ
3gx8O5FA1BJCxet0/MfoXr9vnSShhXOCccMokCOHIDk1CSc9MZo3DQSSUcGkpBlt
8LIqYfWakEci4o4sQBwqFhuEOLlijXpbrqooz93N7Zc7WciXG4tdNg3e0Zs8k1rc
tETvfVX3qQaTpz7oA45V0j19yy1pVsw8Sg53NRE3OsAbaFc7dL+ZpWQ0a4oYX/YI
+qdP66uLChyHi6F/qE/XfHgygk4HwEq4azTiCCgV130YsoNyl8KL7MNxpD5OAgjo
BC5k1EkAr8US0d3XsGr4K/b5MryJyl51DU7v9odT37qlEkEiCqn4uxSfQ703I+Mq
qvG4fLihHXFh4cidW17+Rvlwm069+vFXG1nxR7atK1iuEqTW1WmgzgTYsE7Y9AUo
wNNMFh1iWoZ/eQJkoZNpui69jdj9TCiHR3r7Srq3/DIuqODb3bCpQXRRoDOBOvo5
B6oyujVTRknjphpM41yuskk+7mZ3tPlnTZ/0vchfp5BNVp2uHKHe5sq95GmfCaYX
X5L5Ez6DW9GQwNv2YvFSKwM1XFHQhfH4z+4ydogEee0vuQgkvfqcI3nRv0BQq5Ss
YDpwUYqaRbuB7kXdpYXoMjEru+cPiYavByp7/OQN59mWSrunT1rB7bGBQtS1ZmZT
6c5MYbdWXeoYMZiUcrP9Y+Gi5Tt+nAwEVuE9Z8vOQCbdBOqX8Fk/ViqYJwtpG/OU
R2tEca16tTNMwbJsrZzRSSXYxkjuiJUd+jZ7CL31n4W/HzoMMAQDS1u9mfAuD1/I
Wfkv7jGg63DZV+xQ8dUJ4d7jpa7/TUsrJz2boonOeOksKLfqQ426s50bBhItP8QK
IAEw4c17znRrAKyVpHbkqsLh6h0d9XljiIlFNW+NQd7LsLcmspX+SBtFeDDUuKoq
emPG0BPMGsB+dRkLeRfTEQwCh7SEbQN+6fxUwyTeKHzliTLCOvHOAGpiS8Kuoi36
zNXmWQ+TrJkvAOIv5qyXqMkA+RnrYVfTroe5ekB2njqEfSKtOBsIglpUo1w0gO/V
eTSyvMMBWE2/RpotoEuxvLcODOmGbyeb9wdoSNaVtz0MhZr96EhcjZqwGHr3fJhA
NggqqrrsphT4XqSUBK/pJM9pnBpYS/O4+qcLb5v7XrVA4FmOtKCZ2FIZJLb1PCSG
7qDqIabgDKMvIbm+B8wkDyKDSJ+81VSLUQIRafC7pTiZUjQtIQv1QT3fFkS0f1Fc
Be4A8D6xwpwf+JqcnAf/69VDsFhg6Skpn9cLKctP455/ulzcF1n/lGvo/IrpqMfQ
Gmw3F9/eQ+SdVb2xdTifns2u9zKWjjy7Ndae6JosjZdnaxIncEsidD8W1sp/QfSs
1L2g87DSOs4embXNqi4u0YpE8CZcHnv6b++XraPmd/UiRUGl+E+zZFfd5ooHvK3L
C4gJRe3zQzR0y6hykfLZSF7bckIJrIRuFiqNBYPBtvINLbXrnyQRMlBfOqQtVIwv
CCW3LJ/+gLEPKYK0sAUXs8l7A0bO0OU9OfAeigvVy8VNOegFjqlWEo3A2b2QLfAY
Lo+r7sDCoxwz4Y51zR5rwrBdqUU0+V+Kc5tveHriYT+zPMixwjd/ZJ9RuEzJqZJy
9sePj/pY5+A+qM+ULrACT74LSk8VfgkDlq4SvJqLduB9UTwPTpWPF1EpWCzZFsG2
6qbTFkcpWHS2OJdOA7rHYesVUR2JgR8l4PvWU71aWpMHYm5hKegYAnwHq2obEkB1
5pmDJasU2g0IECfPYGVI/JK+6VqYe6VJVOOuzu/uFJSnEE8BWfD9iVskehPFgcZM
OB6LorEF8By+BChKLpE2SDPkywPE7NoaZlzkAH/sdT05Ha0dG297DgR4h+cHFdk+
iNHd8OSBCCs8puJIXUszFVhpN1PkBe8BrQ3awEa81bs4HiAs5Q3nrcNDXGPDZhN0
/FNPBxnyfmNirIwK4B3wfsSgtYNe44yPAXKMeHKuM24I1tisGhyv/Hxgw+/pi4pT
yi7qn4V0iRMKkdB3SzJ5/GaueTU2a6XodexFC+y52xLqUJABvqgHiDxUZmXh3ha6
qVcXWUloySVOTh/yO+NW7B7xacLSR69sEdiTWJFNsIWynPxP+OvP3lQuQDPV8nrR
NZLSbKYRHUrOEIo4mwRQf4zwG1ba0rJMzZ+j2KbMzDLS9PA13KwVWEljXzikNDhI
X8P82gaQzMd3LZGMfbe/lXnSkqCph/PrJo1nEWS9Wt/m2Li6CP4sFgQA0VyuTGW8
7Q6N5VRGZkC09bhqJaVkCWGNJBACR3d2k8IRxK2+W4vyxzEEFvDrs9HfbynNtFaX
hAtHi//0HfmfTPx+JHCGwa/Un+9coQuTuWKALrxMsCgVlcsgLUFirOUfboCEZCXT
OCKOJqlxW361JSsqsX4By9NrgHn4/Xyoom9TfRVCGvLOTXXhm4Q5zOBn0uUff6Ao
c7v2n1gwkvhxOqFOt3C7eMpROJy1Q2LsCvZaphHahJhhqWj51eC9qHepIIuKYdLO
4zoNmhM9cS0HF7RclJ3x1EePQE3hd5TJtFqbPqj5xlUR8GPI8w6Sn9XRRkosfd+b
wMGyeGbLp0lXOLHiKi9WTK0C/5MOpHijkRPP7aEHEsHFbXghliGsTW7p8+vU8ANh
QTG8orS/c1hd7+nslVE2CjMnNmL2MYmB1wNkZA4FQGRmlbu82oVA6M7onW1sEQq/
PDwclQ+7G6gwxWg+i3xl9tpAYs1FGPLwg9kgDH/HrRKkXx+XQ08/YdJoQdIb8nB6
cRnFVJNmiEMGl/CsSnyXFdGwC9MkfIzqF9Mum1cypbZv8QmyIRYEgp7l2noxFXgt
l6ErevAPFhm5d1s5Icspkfe6Zl63KUBdtRtA0XGbmpMc6wf9OP990TN/OT+zo4D5
vUx8RZczrfv+lT5lS2RvEerhgMepSj1F0kbCyfdY25mD1mTNdpIh2y4+N0CB/q/p
CSzs3TevHNYrBOVoCXOPQHiCXIoQsAnw3qv4/ACzBrpap+JUTw95HdDdDacwNztj
KMMOgPurNwIc1qamkHlTQxxK0v0K7WGw/kIhVWmfum+tXQqYAEKAwqsRSEKyD918
eTm5QaBtpb5zMQddohEhUzOBiQteXRmE+vtprnfpo6NxQqKKjhiChFcnP3zatQAV
b036/4lvr/m0hLHoWVeZXm9MYKIVf7DlKPk9d2VLwWQBkzEx343PFZzpxzd+EjpS
Yajx5Ozub6+s0twmwcFs1JiV+DGtJfyfpYPauQzUuCvPEze+nWAob2geCvBPelgB
qNIWq3zlNcsc++iXZ91vDGMyHYSweEFhJ2IW2qmyzZRDxcnPfqQpGB5kcTArHZq1
XiT+uDSEAmb5Jl3tNO//wPziQwwA+FH+cAq+lYPdsEequBzjI9pvKajOvTRC30mS
ABWF5alySA9P/LCwA+QNkSM+UMfKBiKEh4EB5T+uEMwXlPpJijvynKoYTfe8Fflp
veF2ZhF7Ib71Ays7TmfL+hWVY0zk3KEx24yucaLchSxLRqf0iCKPWhETDn/f3kHv
0MirzA0fi6NBpzb5Km/P3icliLcHL8ranBWT0ywAm7vlMc38llkEwDXKRsaIvglR
BZ3G/mhcm2O+j162VB38BuuFmHDK+GbHpel6I3yQCp82ADZMBTaUPw8xB6+G9npX
nidath/gOIcx/9nY6+q3STN3hruwjtaFmTHXfzvMokzsdC1f4/aZiRkIP5K/APAJ
oGGNJuOVoOtqGfrlbSPy36G8YqrllIle+44p8/YVjbfDBuTxDSqZzvjeDJxmgaUz
8ppWj4Fqzhs07GI1/ZtLjNCGqBONrIbYuX/dvFNiLbUbnrUaI+/n5SXYNuupxcAA
V4R+NTpPRauLGGB9IQtFaFKdRcKp+eBkRnHnIWOjLhwGdtWx4844EuibhX73/lwD
Cz4KUBEodqJgR7slFa+qLkLNYeTRmwTRzC6x91Mb/5srnUUyyF/1VnEVYEdsz6AB
zU437DZilpZYXGThR5xqJyIFWxDPgQewMnfzWearLGzpKCUptC2eV6E61xqKafLR
mwbm8dow3UPpg2y/acCRXpcZ8niLXw2DN1qAMAF61KZoxkE48sH/Gevf+DDVIO7H
Cx00Onp3RwyiiWVZaSGVYmnryGgLVIArdSqJiz5C/IcFb9Pf+MGB1n5GcJyc0Lmn
PGiv4g6jAe0oEPdDNeZnJ4ry4uMMX6psqbKrNF9vrXOoI4yKWtNIWV8CnKChrLoA
aGKL7c0UnzQ+ORNZEtppxirfF2r5uZ5ScPV0Qet7CFfNfm6hOIF4pYc1TX4ZUfMv
gjsyu/Gk+yq+5WdRNHuP7yHkdnS+qAo1J1/smFygzHjQbMavVZJZRHz5ypMOQ5Z3
IxdrUZwVzFScjMiVtKEu+7eR3SRmz7UYzSQ0cnp2Sa4=
`protect END_PROTECTED
