`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TyFS5jNoc0xPal3aCY8ol+OsM2At4Zvzm6FxzujvBY8LXWTrKaEvvaoB8zb+82YU
oArvVtA+mjEeDat04ZQORJkzmgCdQfYZYmyAT4Ik4+sldP8SiZ8MB2hvc3sGqgOA
CHAIccCiwQmXuRRiaaOmj9VmIfiK7CKJckUR0H/01f14PJu/+kbdgGpuMrPSQXY6
dieEhPE7IMQrYSyd8+HB3yDatYyc7ZHgSoQJtYrFg0mQBtG+TB/CMy+H4BG4cawG
0Z3XyQPLfH4Y36jZFvCyskhU6EiFbHzXyYPz4Nt6fo1BUg9OkcqV1BoUGYySg5rl
OmHFt5rDF6F+ezwosbjEr5TUqDyWzKhk9doyFmn+kShwd030b9p9BTdzzZjC8DXY
gK7ZgekVPMUz45BcgrCJOAgryDKLBJ/+u611vjaamxZfM6jxu1Hbfob9uRcAC3Nv
edCdUw56eVP2ZymCqCL5ietB5TNnX5oha6riUtdvKsVDrrCao45xR7n0hxaf57aL
OQSthXF6bSIxqFN9/ez6b8fw2SqXGFKjh5PxWKOAfpieu0M9A8E8gudchvrSQabs
raeVE/Y+fdORN6aotvcmH2CzAljM1bIpI7ACG0Rp60mWcN0b5B4KfVEA69PHTJru
dof6mgYhRHqWfcJLfmw8nSwYXbpv4xUVhgZh//uUcaYA9dlZBPoLrTFt/aba1ON6
486EEGbXIRq3d37Idr64mEMp+NBQRioC0bITYlQI7A/xh/QZp1U4npXqMqqpWwA5
aQsi/yoj9hpHt4ihomficDmXHMessNTlurIRx0cBcsurS7pLlLa08NnYjyCxU5UY
tX+T2pgf104m/pY9ynu5S6avJSloFkyRAEDbC8bGMVaQ8xJH/auR90dhKPSUmz8Z
oubmXkcS4xZ0wkWYmUdtnRBnunByrmaKTatEepO0JNVGVofoWGq0u/MFarNNBEyv
zBsFSp95TTPOM0XWUsmEZGMTzpABEWviAyRpkEajqOOSmdxD4wNaHmIt1JcET5ao
2MQ3GpwIrW+YY8w77bEsA0Gxx9fizjo/jRQi0UkjU9Vpfdb5sMuNwqJxnvx9s81r
0Ec+p3ndwexSUfvSzWHMKXmkVByW3LdYK06eelix4GNihrScFzvlR2kFrmxCqUe/
FP/F4TzM2lN+D11bRQS40Fd909+fIbglFjRqUtaEsWsKwlizQZz+QzJ12Gx7+uOj
//MvEAT8lBxKDuJgNk1dg/nF0FxAs6Gg9q6G/kBjPuRR22WlOKslt7/9xH/wHT0w
2J9S2a79Wtn8tzhwvrI5qlqgVNf8y2KIHsjGyqxlufFTOzJbZTZgq4cK1s2gOcdH
JikrPpLb8KAeActmY3aCOZlpALY9vbuGS9oXFBLRpmQ/FajJBcmvFRlZkpcDHVJr
ua1TpRFDAPk+9LdvOga4BiOOJ2dsc0riq4v+X2jE/SYabV1r3C5HQakTE2sKk8am
dabT2N+Ri4htz4NMs1fE0B1VTqM95TsRG3rJYJdUev6kZQQCfgGMYWuatlOvEBSA
G5jtFs0wBL9QDNaNWLuNstjOcOyn1f4cQeYBgvJntNSnHcqTwnfOmeuiMpkdPBy+
JPaVzu0ruhDd2j5z6k5AszLV3FdNHqiwWQ8nz36mJwDtjhLjGlTUWLDlPN6IQmPL
kgDej/9m/GV6xCM6Qn5nAloMeWSityh2eUnPtNK4z8s8ye1IcNahBULAOdgKDDQJ
L6xNakiPGu+Tfk1szfl1zRBNq2QE5iNKsmUavCTk47q9POfAblhR5yjxYLOrxYFk
vfLAVKLKI5yVJFUpdMFXBf5ZtJTOJjObPeeSkU1mlBlqukY+dLpdKqmWSg3qhWOd
CQWWN012Y5r4NKpsNsxs8Y7gM2pf6cy7j5nY2mTAOD+t+XprdjJifXt6BATiLlqZ
Lw7+ImEgODJEg01pDrIasNfSlQmEWk5r1iEvXzxW430bMooB9ELuZtooynP7NRio
ND56WFMUUbea58nZMERqhHdyWIOO+94Em+y4XXNGV0QA2rQ3VU0soI+qTbWJXbul
57W/0kS9wVRlbf7GtxaL2PhzCiM7Nc9R3Gclkv4fEVl1xtZ0abwKBq2Ctp9Komda
L31sjBhrEJxaECimWyUR3JHM30GTT9OcBSyRJ7/Pnm/6kcWtV1ZrlSZSwRSrvond
WldWzzY60pH/XFhfbjZfVVn8mQ+ZwKqcBRgRbeggRSjsVburjDi1mhX7noBCiHly
99DQnyYFewDULc73gsgbeTTdodHaa9NjCwE4h/tYev04mMeyG4U95qMsv/Du/A1w
vpEmPWx8SfLOG9nwe6c+lnZBGTtZ+jIhhbP34IibZctiDa8eF7wbCopZJsLhPXD6
FGz2E+s0TOhPS6/hv5o5gsSMmHFv1AYKp1znr8TAe1yPiDZBg6kTJf7loe6l20YS
kCFMJQwgHDLcRKElCD0tBwFypyttti1KE2oP0SyqZpkYMT0Ly3tsGn0vEUiPTnFk
7QldcWulfUM26PPYf7T2kwJDuD8ezsnTRiy7RnYoghjVB/j8SKV8rKpf/s2Cnowz
ub1L5mjIWvgVb5yPRjzBswBFdTREAXS//HEQvZn+qtHTVawnXlF6Kj5NNumI1Csi
EeJE25n6hIxw2RVVyDuvXgPXMZyzmab+HgN221L4Z9JPuo8BWPFekJ5vYeKXDcUw
RxVXUQVEfnChQvdrPHvW2kl8ETjF1QZtW6TFQY2UdU8+pyG0oL3l694nYq0evkFl
D+clb9YNmyv/V9qwRSfVflJUMdEi8d0Byys1Fqqn82qBmCv9LEo5nQFe4V8MVgS4
SnPOjU22rE7JuD9dxTP6RnsLYTH6AdrAY3LaFD94HqVWT8+6oXuTGIZrswKHveSu
jvUoQVVK9b70yHHFSSWtDpgLo0zWBQ3Y7AvCjaNDNRIJ+x/B5U3aFdDlTR0WGXHN
KKf5zhwwnrzhCWfEI9MlWzfsd6yL7kcdNtDINcgHXf40FrMTfLBsCGuf+6XfuCbk
OKlv0gtd5wpPgzLzgp+IphvXVzrBEsg+IRpS1SuTeau0JfnA53oBkJghlSXkK2xu
61KlUhuQEQRzwMNKj98/TMhlWcuvVGuops+6dh2ylYPNtlxK5Djr91CLaazruIO+
DFAf+E7hpGFpykKbJA7M7CYyT2Fv/+0tVxZLuyZdIbsJy2osbFkHuNuJCR6MlH0q
5gaSyyEk3lNlmjVZAvH9HXpm2g3+DK64wl3tVA602G2F0U3zqZXydhlslwE/vmVo
1Bg+eUmZAv+az/wwJbHXu2HM6bzj7ZhXTUf/th9U8T4eAkbK3ZzeV18doHMsEGrJ
m11JU6JlbUbcGBjBBDP+WgoHN4J+k2mTZJv/9vjzIrsSXrVH3q4mKgsyxD0frEDn
d7QR4+27UqEEIPr++YuPQxw84F/kgX+v3v6bbnizxDuUdzSLHQ2QVeG2tX3rVdxp
Sq4OrHb8n8tP/+fVx9FCC9SutFrIiSBcaqHMbWs2tqgdA8u6jf7Dhe17E/VV4wk5
04F+YXKxaUckM7UO12QqfccTZ2cbXBbsBI0CCDPlrnd1zyyYbneqplTbpIEZ+MCU
SpwtFnfskIe/hVaBoWS3SKGxT0w9hZbyrLerKspWb0pry6AIQn3oLNrBZsx17RBm
LuHes3+PjDWefCkqtBv0Vy3Qt5OPrYFoVhQ+HnnT6QwNicPRfE5AdxmUq69dHdnb
O1OHZLAhhOizEcDeZSKNBe0Em3VhLl2eaozgo1Nmw/1bkledolyRWk2uExcULoiU
j9AUzDdSO+Ov8Oipsqxu78GBcP6u6AL5Abqow87REMcxT+BsD1cqVdvHSZw/eA0w
tjkIId6NNzpRnoPxVWqnkjoPnQ7Z+nytDOqcm0HpJgaFaFmGIBCabMPiYe/5zPle
EV0LAczqd07c5TNd1TFSxvz+QQVjNtcKAIDgSlscFaXw6QDlff0D/IvmII6ZyOUO
lz/CXPRPyHD3AgxlfVpGE3Mex00KyhIhxWUPMbgNz6cbCZgyRthsuppQHHF3a+O9
s+Zakexn64XTcPgZZXAip35LUffeVb4nuUsq+DxqVIYnF606MbRM94Q8JNZ1afcx
rTLHtHdMYYF2w0sH67JgXjtTco4dLVb/f8huG/VnHB5odofYR7sNmWmScIci1ra3
4CwQdbIJ3RP3Jj3VYbATb2lfpnHyVD7QliGHWrIk2Br3DRZcSqntzAV9oS+xLded
sLw1GzgRNh8TEaTPjmlnC6ZLGoSGHhOPemqiA9Ot8XroFHOZeTgx9iYoLhpXxqxS
r3fXaHlj0ewH2tFIynmfVzMy6suj+tW144AQ8aV3tiXJaTxQ0H0OvsLamzjhmR7X
P4wdVVLmMMQf+V/nOKaLo7bEQE2fMKp5HjKig6Tia3H5ERilXwhph8JuCenimb1t
Skjrqh83RdYoLrxM+D8n+eKTdc3U60OWT+qSHUkfsn6bKSooVuidE6NQOSO04l6C
0Y4mmSsKXpyRiq2cTB6L19j3lfJNKSWxclJskwSpx115E02djYX5nstTVL1b1NWK
KbYWMYrKG5FiJFdu1akn3qtVRmhdVdAxsWs4odkCyQENIPrwBQQ5UvOuJYGDiUlc
vYzSJyvCq4iYeq2X8dvk0ISo3aOeGt3ayW0DDoJ8mNf3Ymjla5KnN4S/53LnXxCG
4A6yfE2dy5Iqr5m3MReignG0VlSuO4QaD7L62TchPkCkqWXjKWH44zqToDNsAyOW
7JeIee9PE+fjcww5flADmEoJSQG1EJWwyqH/gSvAtRivKZW64n6M3ararfaIHBej
rLXtOrJ8LXrqVfJrOEDw6LtXbFtzjK5pulsb7Lp7RnGnVuNsIv71E2GDUPtC+YWq
RQ1q/tJOLnbResH8iSMsx28owaICL0lcyfORZutkP5WvUUa3g1gcxHhjaZhzV45N
W/f6NOraiMPJyGdDdqOx89sRSg4Huc8dr/07y0jhmjfRD1efm3fmm8SQ1pLuT/WV
rgwbdFQLqPpvXnCNX+SWDl0FbNmcG5GWDLhRfkgY4coFkWolXiQZR03yWQxJI/sw
P7KHIQfo0eby6YLFBIkjEKAk3TGXcwNHq73kbQb7JGod6t/hGP/VztsQiexONGmw
ExGQZx0YJ4qXHOe7+d4HD3fVU+//UC27Jz3qQX+eRKaxNfetKXbKO98eUh1LPWIY
pqpl4+G4PeI5e3+ci+KSR1l3mjBqjYijjvc3pfNb6dGpkVt5i97nlJIAt6OlLTyE
eACgogt/SAFoPc2lfLWjejZdL86VBLsNRwYvk6c76ulrEWYoncNLGcuCjOIn2mg1
xku8OA5o9ZJ/qQPL1ElGxJFYS56Teo1hkjbV7PjG+CHRaR2QbOHvFc3xt1nIT2rS
Cbgi9jPBW5cUJVUma1R809h+bxyEWrmeioWgsqCyCjRuAOZzlB6Vu1JGnYpaXBQh
Q7960+/SgQCMPfry297fMnajqylrM9pB+NY6eHnFUHBvwfiluMJsjYO/78rci9t9
Jc+bOhBOzVP5OhDXYinLBxhEPzRSrNn2AXbUZr0WTFQwCsl2aC3fxGKGHAXXVD+/
Su8sXOOegYe4tGHjiJqVPpSCsQYxl2m5BNM857ikTivKdTtU6vwxmUetXyE2GAf+
ubuS6q4mutNWRYCSTrfwYxsKRsYrrhJ2SkXX80nrMXmXtCG49F+DI0O0M0RmodXA
q6iRPl5cG1AN9KTnF5hWzo/5le1pLcv+3n/gXbV9WgsKx5O3u4zcgW+5l13FPvOU
asWpcPEGs91pgeiSMyVnH2m5swDI6XgKdpMdgACk37bw/vCbug2I3BghidfdDRwA
m1YqCEX6aANsxn5ZDemkP2tPbDlK3c123l5bPkgY+fBhBVzTaAl8z5sYcjOGIlue
wYPIaGMHV3lV4ILdNwy6gFCp7DiWyRUJdqB+ZAd7TjAadJxbeFcVcZtQsWRH1IoF
+kjDiIATjDtuatF1wZMMs+GSEjfQNu3/MZCrcirIjXdSysxtkoq3ZWs0uvNDKi7/
g/zmqBHBIa6b7Jd40z2aVVetcb7q3eggXOYGYM/ExZYcOqULoJsYTPQwHVOX8a8D
EuZNnLC5pxHGwNBh8gPJLxkGs8MBubSYcegF+yPgB5Y5PTUYOJjdGgsakz9BPar/
fVL0zZqR3hFPa6uJD5XXyqTRyShsmzzKWBJWgbbfqC7AJN2Bm/92tXvcDnUX/Wwh
9Dcxrsm0FTH+1DA/gLWjR9qSVbwbWtNK+ipAMJLzlpOWD3+HXfGhPkd/kx9u2mUY
1AJ1GOGacB5FV2YyxV8+BDkv4gqe7fdT2t56c+xRgSZs/livzMqW9uW8ng3uDU/P
G6eO/psyCQmiHEitOwq4+sMt2v5G6Z54ghglgKoXc/WNHMtpClW7ZHzN2ZM6AEBN
rijdppMwMM8VogzUdrPbwK4yfNffTaapRCUNZa6xzQ3q+byL5S+oXFDas8x8H3SM
TnIeHmkIHPYhEtgTa8evfawnAiioKMs8CWrwAQcgYUgAQb8n+dhJ/lW8ZYrCiyYl
qsBaJBjxOshuiJ7fNYsXqWxVk+Y9XLE216Gbx0YPHYP3Y/rciNCCSQpqrKb/JSUs
ezfEUzAXM/eoZrchI/JEnH68deVXuyPmGLOSpUMRZbcNY2fXI7jmxsbNmilV2ds2
fc7gcx+Yt1bDgWIG9sj0m+qDQmCS0Ljzx32S2AEJJCqh0ztE4x4oMo4hRfuN/RRa
+CPaBYmyY4wzO6s7l21N3sQI2FGk7VqHY5/MrkHrTjSeQdfPgltQXxc6RQh/Y9AC
kiUb2Lv4juFgTxgLwfQCspwbcSmFdI9VhhL8OPqfQSgToIFb0bqiEnIQ6Ofr8i+p
kArYhxpfrulKyamfH+DHJknLz2Ht/XvHQYVeb6zkeD5AAzzdIvkh4QO7pcDJzKbh
uZGo5rRCdkUFzQ7uoYUqh6PcUSWT/lJWdJvryqBVgR1n79cYvGFqxk+2Drof29W9
iYVAgvV/Es2ucgvJsfz4tBtFTfFtm+XuAHTz9oCtD1+0s/cpulLb/n+hGGX0ZoyG
KMTb+xbJaiEOSV1mAGWFIQbipzFF1RDJb1l1Z6DRm66qGthIAH+nxdZUY24eYiFK
gIFHTKqyi7SlLnb4wRi0pxDhaGqk7Cw6FMCohhbdDZTtP5IfUIdG0v4syQlzPcQi
f4xr1DyWXHErRExsT83PlD0DVMRL4B4byJlF4ft9EGpDKqnL5VqmcvlB/nWKi8Jt
bz9fppFllTvXK4AVV+8s9qbirvWTyNtdeHKycU3gRZHci+NP/xYjEx5otx011XZV
R5clKx4fnDtSyZmVsWm2P4JVC1mH+UR6thp6+wyj7f38JEHtUo+GLZP2IguuDQiq
+0uUSyuwR4TMbkqfQkKv88cUQVy6btSdHX/WRAIWBrbd/5ENzCbTDVSyZ/nfdPV7
7YWAw0fBKjPPZpcLpidOrfOV/bK5y5getKoziC9OolHNN+MvYwj+vWis3CwgHSqy
VZc0SLBj3ycQsyMJEOdcmqsNYXHkt2A11LQM89gGSeT7LPJxI3Gfkusl0WvE7BvK
FIV49m0Jw9NvibrHdc3v12Rjlf2WuDO5JtdZYEXhBRPQ3tye+RYYY4DD0OqWb/Mv
M8GmCMR+p/zm5dXEtIE+2qHK8l+sRG7kC12Qpjd3bhd8+3opfR6PsfUR8j9MSDEr
QpHJKdz4T3Uwcqn6dBzIj+taUu3vA8qx1JIb2dhvEFiWU5GduuDuySdh8wx7odCR
K3jzNjJsWz7OYLBHDK7gRLY41F0Pus5hyxJM+iPaZVJ+5mhQXfIydF9sbOxZU0Am
QEUxAuuEY+XAc/SSpFVU4xzyMjvjVUf9hfjDWKJb8uV131KfehKPDhMk8pnBZRaS
CdWKuHExjeWktukrGiv11pFKS7n0MI9Vp3QhGSQ9H49lA/Fq5VzyGkxeSQifk1xB
FKpmcnjxH37h2oqQBML+ONvVRiLJXRveQOYL4ZvMB/yTQDQYrPSO8xYp6BzV9b5b
7bFXuL16u6rAnK8OSzSW6t5m7hkWMAD7mEh61B9mqNEPw5FaU/REakJ6EX+UMXDr
osdim0IpcHTNZHurVkDn6p/DMeAYawhTYpIfspA9UHZW/qyuC5o5pOz7C2sojVbN
pUGEs2dKN/RsrRNSfMeFhkhuH3W1f73bcBDaWtM6FcX/yzQy8swWKSyFnzRIFhkW
Ig7kBBcIWK9KsxJeQMp7mJtcfaXteLyH8iy3kPdwyQ0/SDWJvBY5ryd86oKUi5zv
0P/nU/zFCSbhMbOb+kUvLdT53bfN1IKbYsQx2UdAN0NLZLN9lBgCIX0POj2StWfi
gLdI3ylwh0+s+075YsSvrOPHLNk6wG0SibJK5kS6W+jXUxmfP6kPyocj0n+wXFoN
QCn1zICrvzelmPyR+IjGLeHjxpNMYzyPTWj4SfvNSUJcUzI8J9qBrg05FcyM731x
pbdb+/gutZqVPp8g61whKybc8sX1cQKeB1yg9Zw9kK7gqUIdWBdVV/mf8fxlsFeF
z7AQdo5iqjievAVGurKpuYmPf2EsmcQTzkz5cVaNYxsQlV0X7I1H9vUsNahAD80c
LzBbJdeyeuvXWgcpXyuVPvrHoJwubyd9l7BMKvSJjv0RKceFCKFBXaGMb+R1BTIp
5hHl+LvS8NpBGDz2tGTCBWfBDV+zSq46KAQaTPDtj1kUaH/wTrlSSyzDxsSIQw6N
7dbH77NLAC9809V4xx7/ERdPGphxrGwmpzbg5BwqPKJYIFoFM4pM8RZiMtc3Z+iP
OdSVTRvqhVgdzIbg5ZEFjObmWx5eNpEWOB91ENOMxoMwTzw6Kd0Iwj0ylyVD1nD9
+89O6vJqcS03bmMy1VH/VIdWl31yGRaBJeswD6ShXsVX08GogNs2xVIIm32puKBt
ItzEXCsZt3+vKtqdgESv5WcxKKSDfpB2JnNzqoDl1EiZlmtJWKgJ5KHtz0o08a/q
Z1uYECN3fERRsIEiVDcT5/Yu7Y24ukidRAuGlnVbeUeJTD98oNTltCW/KXbZEJfK
f3SWnoOPdcTmAi4zTFAEVjm8RVIYv51UucodGkpm4ZumLLgTxw81WLAoPSBxIiSF
7QQFeIqi/SJxbV9dBwT8t/JkLTHot5+gTCpGx1XgV6JBTXfhVX5q3oVNvOdnDw0p
uaZDfF1KZ/fbRoOc/sMaLm0imL9YfGhnEyp5IGPO8xryEZfPUFvCfUzLF3n6wjcp
9poecFzpfPdwU2H1euV0ZJM4oTKqMBB9RjY0yHPQwUV7Iau1NHmCcj+lcZ+x8shA
qBLw7GnMhGNE3cGg83+d1+Vp/EBueiCh/t8fvm9nv9aVeOGytv+y1Txq6bBK6tl8
5/T9Xf/2TSwaTfAhkEurw1RHBpQfjrbsG1t3UzhLuGHN2N91GrGWdH6LDC8dvCvX
JUawRQj1GJQfj41Q7EcsH2tCOkB0OwW8gqUYL0nJ+rYFed8lsb0+VaboeAVb1bN4
pk2Dc7A46s/rlVFFf6HPzTqUcrAuTEXJr911sbGkfDpU4B/kCMj8n/jgL83PA7QK
pU1peVrFatBrv6qDJkdcfDS1TsJrRb03AYAoPm4sjsr+2JQQzLtX9UZuKIPxiO9g
H/gZo5G7ZeVPz4mbMmgLFJbsXjn93KcXUJ1hFgp96BkEEm8GEloLKterpnbdF4Po
zGxPjpGGy04n7V48BZ6BCK+UJARYuOEUVs+bMR1J5whaJwdax9CpEmg7wtsjZZzG
GkU9Di+aQGI3PDwXT4MlNZnlW75KEtJSL9ferBVDiQiBTiuq0CtJHWMsFbyELWgg
i6CDZM9hC5kUMvCfq9o3BBQHDVj1MOXTPUwDYi8R5QgkMKhsS6+X6O57uKxWH2LG
TLsQBy8W3gdoBXoZL5/4b4neLwFsk53FsLGD1L7A0pjXGZbirOezN5GFUReV6A3t
54wsPI52O8HTKDANnX1t11UJxZyUOW/VGbBZ1R0s5GeWr1fZDjvqqyygC7NT3Tn5
QqluCkj5qw1/SNr07q/VMpr5ZqjNJMLALgScL6l5VnTBBBqGMeowUEMG6TuOvEwp
iv36FSASV2KbAzr32y/O1LPJoe583e+3L84DJ4aRi1H4mXLXDQleF3NastBA5cOf
ENKwpTP2xAzGsahqGB5wEmJJ+YMLjLFtcOyf9Y7JwPT/8LlWvtttfv7v+nqvkEI8
nzr/jJ81Uk4O70KF388LtCMrt30/Pj6BD7qS5WDE+rAUKy76nR45DRvRf2XBcTx7
OGXQr68jRjdhLzRYOIPMUfJf5Av9L2Qv4djObdK4lSsRMGH0D/O/fvAgeT7oP/dY
fMwh/8Tq/XP1+SK1OZrmsWE8acw96CFgETk0lugCU75Pwt/kOw/rI21ukXSmxsFS
+CQVyEx4P0goF4XDSdIa//Mus2sKClMAWOihO2DZvvuLqzO7hkvI62UYAu9J+AvW
GlhBU+gWEQ1bQjxQA+WkdUcWFQXTI/qPr1+FKdGAyFwXbX4/CPQLieT30vdxMV9u
cFqNyHFv5YrLwT0reQZtFhs8rQTxyKclZhcvd8iRFrjHxm8cR1iz29z22sOfLmWo
I//JlLhPi4EUyVANjAyOdGm1A6VW9EIT52Xv+KaApDh73BHQIuaD8a1s8Jhi/KtY
sJDdWuSJbkTWjUafikNYnCbw8/eCbE6AWQnVKcPbKd8VoGcK1bHPSFRd6gzKFtEh
+nEjVJTwksGPZ2IZdVLPqeXpa3FtYaD3d24H4FZkZCS1fNq0btvOjE5ixpnMjmKa
dbTJNFyKhrWXHPoR6Fw9gUVrTIVBrBrFQzm/4Yupq49Blkdzg6TqEJQfADIoUCW9
DRFnpqm6NQEoC891Ermm7ZNnbU6n0owq1SGe8YP793pmQctXTCnqMuSc6ZMMo7Rz
l+2ve8MPpANqAZUQZ13Hb6tx+ufM+A+xP3q0juN3r6oIxsxAyMSX5EenSDiFqNxX
XfalVWMMPbB6eQrKxR/UZUr4VzK7Yic33GjfE3e9VApb5RKzy8UrSrfYb7/tSJA+
0V87Byup2w/Pf15eNIpmolfiRT8AIHxPuMnCvgV17vZXnGC9IzkpEwXlUN2jxl3D
P6EZ6/iBVHTEmtZnnkSGHwTCUSEo83zPXDLHs6tS06o=
`protect END_PROTECTED
