`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IOauUHcc03shQbK/reqpp4GP6q6yU4gWHMDLoZUhDBcUPhsztQmzNNrjb3ZjvHtI
fq2oJgzXotOdNJw7hxJZTOeCIyRBbOz8xnoGSEkvW8bNR3L5uqyk1PLqLwvXGlm+
/KGb80oW1nJkv02R7X/qimw1L0pgGLwsZI+OfyMQGZgVJAP4JYJOq+ZEOt79a7dP
oaLr1CuRnEcravWIonxUNFKlYbIs/Z0fs3Nl7rw7Fn4lA64UjuD5A//xsAw58X69
/JC64fXKcJaxBEEKNjCW6Ap0nAE9IEiriPCKnKtB/L3HVWc9YE5MVlA8yWaDsUnM
y5W3Plw2swVHvRK17kZ39xTimOtY0Alhztr0vRuEaj3QvmNbI4DAD2LNxb18ZhL6
cOVkfEn9FBMhCJKL4CPw8ckCsFiKYx6VQ1YE/QjA2PRGFJ6Ih80UBtWyHXGxX1v8
JyfUxiQJGswYzGZy3ECdyhkDN9aKAgQTVWdfgq6EQzEEQOOf5DJblouN/f0gqN1I
sNcMndjnAzVsy8Qlm+rBvl74/GhKLa7H/HnCKtZ9tb1yPNLZLQQqN2wcRlh8GS2I
z943naIjcUmMkAcK8h3IvEMpvKtTv/L3+BKCj/BD/vz3CfOE88gFIO01cqYkOiwP
hCHBx3sOJu+yYCAA6ss9DjKAofGg8HGHw20UjamzmpNBCFGXTHOhJrEniBIShVHl
6Hz38B+RJUay4NX0Q2dIP4/i1AtL/ZoowUGKImxANxQXOtHHaTyejYlNh5I9DEJT
/+Jg6/GHkqm7QjZMUhEeAnnqmtTWjlX9ma/dr5dqnGSXWJ4p+X1+8B5RHMQ1+apr
DBYPSlaLoLfc6RweEyX/BufUrSCzGxLhYnl/IpEMGOwDlqg0n+PTCyNxozVjyvbj
xOIKeu5k5wquFZqMShVtkadt7xGLE3YIuKC3Thu+FnTzMiXIWBFUDE2+ELFwkG5T
YWJ9KC4+7+TZq2D+niZSGsELC2LXR7IP19ngZqkh3l7KE5FcxSh01iNSYqFtBqBk
5DWSwOow4eKqoKbQU24+PYBJzwRPT6cXs9yFUOzeqlZI2NfaOJAavTI0OpnKNFS0
wevvRm2R/ahbyU9cLcFs1lT7zqAPwYBE11+cWo0mYeLnt3ohf2cA2LO02OCfOAwZ
JPDIs0DnOu13Tke8twxz68fniaDja+JLJ8gYP5LMEbG3uC089ETd2YsQqIQvcI/B
HSFhIJFLZpnBfINgvbE+FzRiElNv9VZCGegJ57xbsolYiPAHEFi9mtCF2OX2K/XN
UZO+QbazQb0SLO5S1xVCVChvB7bENVJzj4+b/pQ1L2CW2QygLpCYxGMH+WX0IVA2
Zd0kYtSBKHavVv2ccZzTLBWRhI745uftUP5a/f8p0VFSJqGYoBIfCtmCMkn8kk8v
a1vC2G9VRxnCSp9yTOc+3GReoe91II0GlEZt9rZpf/SgQdNv37j1dClcwB7HBhX1
4cnQzde5pYypRnc5NWwlNp2yODsqTiaPfBM6ru9XTbLFZHbbIvTWJtABpEeZKdoo
Iw+NjsnTZeNSOTp6oHfhMsh1hnBhf9CffEhgQ91sLv85xb9BN4cbVvWUc/FmNwZA
72dWVczSQquXqQDhnUADOcOqrpao8+uBBDGlt6utgpFI83whjW4Vgd/RgzhDOuO0
S4LxbydaYqf7FUQROOk3Pjh6HFo7NCAQceSV1h9BoKptTlnvSvLLJikXY+vtRxT+
jkfYOY35JGISg4OuAPg+nwRGIbwc5QfQ4qm62EUuJ0DwQoYPcrmJ86AzKSSSo3EB
Wwyxa5qnYJ13nGYkLcGzsvkD+aQiaHeoVJkrWZB25QR1g6FASRrVgMtoTRt3DrAu
CWkCN5wlMvm3WVr9JOcqlc+7SoHSYWGZnisc/qk7zaZhZXMDhpkVD3pOZqgShZPa
3Hq/Bc9LEBkrjJ+ywtf4iWP8q77tHQzKiU0JPfvhM//dvsmnL4xz/+8Y5ekxDp0G
0nZHzX9KnFORVxGsQ5gu4YG+PNv1+tpUxLd6rpwmY3NOQFGVsdK5kBTi1L4NXteI
i8DG1UM9KPGUhpyz09B4Aj0PKplRo8EcOEXs9KBuKlg1n2dIzNf9/sjU6yNthP+F
fDRDhLZhbxOoQ+QujpFkGcf6BdmsOVUkUJOKfHfdKqWBQNx6DmzItYjt9aM+/kLZ
9/xyZpQ2Lp5hW+Fd7t/Tc+AeJYITkYJRTHeN/QvEsrvG7U8wXtXuY/7Ns6kJG8VP
agbcnom7+rUcdVvwMjTA+wx+Gl8q6h5TR5w8kDXAFSO2X6NtUWcCdYd9UJMcsLtG
5Au4zipzx3T4mpa8Yg3MC/maFtcCVoK7IgMwVjjiM/NvcMtnlOgIny1gkjVIcCq7
U3fKF9DKplOiCJm5DunApaFFEtSpMhD9nKkxrT+7yuw83iQDpbeKRsxhq+aM2//s
2q7vWjCvY8mZsjhSjOmqf5jBAbpCaZjZUtn07P2R+36Va/P+wu2F2U8MTbKWfLas
y4uxUPmGJ8nXNqDrJNwFOFmUqXPLD4T61dIM7FqzdAULPDLr6cme05Qsb8JyCwPX
9S3SnpZRAR0otovj6ig7S2fIGdZKAORdVz1agb+JiqL/XxwfH5gOlRyWlbxlebIY
PHEAWspfodPgphTJ4Q6uYkZvhPUJaojqBScATckLWtoZnLNVHldWy3Drl1GqQEop
xDi9oWAPt23nAHuFEAD/iw/lKpc+uWfZP/G7b37iMfaATuNn76F3MI44okQTQ/3r
JKpSECgj3mNzF47sqDJxS2yPLyhQLWAeyFg1AD1heJRq16ZmvcjefFzlXNAOLxpF
d8FqMKqlUfAh0A6STMrgo3guRmmKIvjf3eoGVyfHTvYdYskUav+7I/+GyMJCDzTh
jieqwoUlmR1XQrP80jDtf6q1QLVZ7PIXht79UiZRVfZWHgXynS9WbIIkl8uhOku6
/RcueWW+KHtFZnNG6qGDzxRhI07K4N68jhOspTkZrWiqPtnerYxju0tAv1Com9ky
ipfEKGlOp/nvutEttF8SuRWjOYfv5N6HIu3YXqp6URZk96T6qDmzGgxLBKAEhEnt
8YzAUEgXJ8eVlQMrknI6Qhs7/LAbPeB4PHUoDFCZHmesz1YGQdr32+htA4E+14h/
j9JT3sUrs+gmbrvvLPRrs8RDeCtLi5+qe2aZZFXwIEnTq4xokErQUGidlUbG8G3p
O5RC4qcCbnTZxA2ioIffxjLzjekZATMiaaZiQWVUogOGO/1AKAuC+6GFF5Pbuh6M
9wSVA1rCVmqXOcgyNflUZxRYvqqGOADL0ymqd6i+XQgbUhxgkYYykET1BQV9RgnF
3siCNWPeK7APm4VxCrlxHvjU/D82da/5EKQ6Asnx6eG4/0fLHXzMv/v85n6e+OXc
lf1z/Bc48umDYm6THR4ZdnQLdB2FFuHVih2c4ptM0dRqVEycTuhu6y7UCHqk8zIR
ZM7tpMnsywdCkWHETVDv1QxcQZTT3JfFiBGuZrRJo1CR/wu/JYtmRUD98ZrrVFVw
g7Uspj1o+Tf63J+C8LIy13TuNpiKLxAZBpOQ6ARGj94id6jY5FWIzDZgMRWyhR9G
VbKfMpOBz1IzxeCm6WVi7JBoxZyFysFdK/aqXoBHvz65lAG0BIlOjiYSCW+lGjX5
DETK8tkgyfeLSAVaaREYljUZX6UhKDO2zCScaJyb052eEQwEvt/Pk+8fdw20T742
n4Je7YALAf9N5jxOxZmFgG0hxVDlkpOG0t1wV+JXI26ljkuC918J/bOmWI1xgVY/
SojsCMUtjApLfdpT94bXwNAOopKoETf6Ucx1n8dyxgp6lm5MxhpKEy9k4NWWiQwp
cPHi1vddx7fQ4RGuZGftaxmyzxJ5xK1GZcvyBHRVGc6VmUzWPD8MAJ66cqPGMcmd
EAc99NjdfBamGu+T5i0WS9sjtCCIz7bD7iRB/ZmRUj1jL9xBwWHRLFn5oOuXlNIW
peWMb3H4OTqjbKS8z3gFmbKg+xAxuQ+b5aRJ5O5vVmJECu43azxLJ3JrL1ld3vTW
24WnsZ0YhM2Y0OccplTD3w==
`protect END_PROTECTED
