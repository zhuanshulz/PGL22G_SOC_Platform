`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
33ATFK14uwFNMXM/q/P+/eSXREyVm4p3jHtf+vhokeBjK/7K2ATW52MiGSnJV98h
LkDTPA75smEP0lDo1wLzFWZCwdq/Em1/5F5Emw2rJa9r8zz40Nem2BBDTBxRtdWb
LnXnLfTIXGo7s+TDxagip3H+sUqpV1knQXrfSpWp+HsgX1Xxnv4PoUFhMzQ3xnr+
o2iNg8LQtfyGZmn54We2crYptoOAH6JUEXwArckumz/wOFjbZ1evIPCRK6V6h6Vw
isfjR5ECW5Kx9omuwsz+FHB/sZD1yPlPQ8i+CM39A2M4h5eUZ10/TRhTLTDd3LFN
vnc6ZB7biqqt9IOBgomkXkRqYv+rNywzGNgYD6oUX8cqVfYwDBXhyLPJmX1lOrY2
HDdUQgHfFQbM0Lz4vOtyW8ZVfNbFoQjV3Vbiv6hJvqfOmeoiOKzJfa3PoTPqkafk
G7IdpnMdN/FbcjS2izWlqnrKHxnsOniTd3KM74DmB6KqLHcKC3r6JOtMpQHfJy/1
TVkZ8Qf3a28b4bMpE22U4VHqFtDY59KmM7rZeuqgm2RdGcMVpkT+bzuJUFQKAg15
3C5imsDP650hHfF8KpIXYixGf0PdYthZzJH2ygwcXH9o+YXG8BBC2ukd1FqYATip
OO/fQBsLY61ndJkj0xvYft8C8dz5AufKfSiKBQ+qIoBcd4eXgZVlihGpYSs/OjIT
m5Ze4FqsWoE21W79et8rH2uIbaDyy8NOP84AGSbLArwO1xOP196dihZ8zXOV5Fti
AM8wg4scJuBLAjpQwhmfMHbXaWLOmJaKwFj3QSfvbSi1aYng3sQpuWwKTVkGJKNs
lnUbtyS96KEIRJiw3pd+dA==
`protect END_PROTECTED
