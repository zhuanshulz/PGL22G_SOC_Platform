`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A30yRUGiuiNnjtZUcvlHcaRdeyAbwE2IVp+QZMmtc3IH8juGad8tF9PlmPlfw0Ci
wzLwOfC0h9WKIPbZ0QywmMkkSUMk0iB83LmyeD4uzBOlEPm08IVyIFdVhrfhg8Uv
tlST2T204ZoC+TgZJ7RRMSuyahCfWsOzNkl6T2N3kDGLsSvV9ZSD1nZUFMITM1eS
SLJDmsdhWvy+WL7L/Sr3xFFUXnF4bVNORra/mXrZAAft+UjUvlSXoSpetMTHOE02
f09ezWkO3vZi/g/m9gArXPO9z19l3BjTpBq0hq5Cg4TRQAGAQJUugIsZ6UdZeeQX
XrA8X4J6Gz/3iUvDpcoBvCyjLX6s2QqmucX+oNHlcsGSI/kZqZLrAqz8v77sTDGd
Tn7JA/r8aOnqg7lzovAgNfC3NYp1vnpGTGs704kkuTdSR0kFszOY15ifae/gG3s7
PuP+SD7y7jrU/IzF+kXypS0bIDh9WfHooBuZCkLvoMmBu/ryR0yJ+XAyhfRfS3w1
I7Pq5kVBrcAmj6l/B2bLrym0xdcBjQU8/J9EIfsla3NoKrlC84bJpAIDM3pqNym2
WzXepdPZK5MoI7sF2fbZda05Er5xJFlHPEtGD/2ikcmd05gsXhhegcpJbm4lV+gy
HIelapSk2+D0EWQgEZ2hFpaNwliF1ayq1SY8GXbjcfEn+t/jEdGE/9SI6BI6zstp
CrMxFPgHizSf2nTM3Yylu9F+l9drJwP9K6d+jfOJddrjPKFk37nMANp4W4QN/bVT
7qQ9NagzUD1iXVOv8BuV5rvp+MUM80MJRFZOc1F6eLjXfGCYdCDye1Fkbex6l5YI
Qh0Ka27nLB799Xx37LuhjFfBaHnfuSZHy2DE0yMkLmiTK+31fkyELKZn8GulmFSG
lTWDdAbyDvepkn96wCl9tYDiacuN9on7MIjqXYmAhrrp5lbS6QpEPz1ZVQK7+OyA
wDQv3b87TTIButiWSOzDl4wyZTPm0ievNsYw0hD32cS/BI+mp0Z6BbfdE1Lyl7dG
xdqIvVBfajDngBtUom45i6PV5M6L1K2hexGbfss8ySoZbFn12Ljre5QPWjjGN7H1
TyL0WyM9D8PPlUlUOqj1pn7ggR2mVcK8Z4mmhPlYmHY=
`protect END_PROTECTED
