`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QsVGruGMq4NM39XsyBKzHc6FZYCcfu8cX915ctITfk1IhoFHzbuRumwL4wUu8H2K
lQEIzpNAKHRbWwwYRfxBw2te5I9q8wmMvYJSQ99x3mhGHAHVzUWIdNeWsnyuGnAd
AgIU2pTOJlo5Vwig43two95GLcezFZNNfEv3KHROrZRsyg8B93wt8NjvIsluuJ2N
ZLnCVbHeCEos39rpOUQE6wRhqlf3RUVfIuXUG6p9AW/XE5cD3z1wMAA5bB6gNegA
XaWwXMcBGn8ZPFrURKi047OHkeqRjY8emS/KKuZhaJ3hjq1e6x1ZN66gE3aqdNzm
r4EQwFMiNlqGyd+8bwpxHqTy5nrVKCo4eSzNi61Nd3y/KXAkoZJ8OU4Rb1u3aCWh
HxxI8Z23UlPqGUyVhuQ1ZKS3dIZRTf9mvrRm0juP6/i2UnRdVd1BlCxFQjKi3m7Q
BRFIP6i1BUaHR6ZNTyQBy6JAAZ7n7UnGpXzJHPqNK1aLgWgOrq76hvSNrh2F05qa
FOk8NMTo6yfWr58Qplv8zxK1acR+tVFQlMJ+JiLOyQO1NmzRFc1MO8AbchInQjoN
E1Ohvbz6AfRBlWfXuMei7t9sYrEyzeyysOob4PJkrO1CpfeM9EiqzZ89y568bWfq
dJcJQb+Tu9TTUqIm9rhlOXljJeKcTqWYuD51xmjzyTjMVuVJ2a4zqbE4ctwl/b+i
D57/54pEij0qL8hDLyrkG6zuc4Z86fTIMyYkupvvU8bXMB0c64ZepiBe+P4jR0yD
+t5/PLoqj/E6U4BikuW31dAwq3hs6syqerCxM5nYTIQqfgVf1WRmmP6vubOq0VSV
0Ms6N6aMVR7noyYOey24zf/OSYX82Nh///gZHwQZ3rEgMDuBZOELmLEEnOIWAURK
Kr9XzI0OXtJPEoJC8pG7wtp97+QGxE6PBbhtCowcA961SHVdCCWks9hQVE43QdO+
9/HH2pDJy5v91lnsI4c/cienUi8UXZY6N32zsBG/PoaTHr0u1V8Jk+e/Od2SITrZ
FLCBWJ2ryJw1MtqfB6OFhy5RE0JpPfQlqzs2q1hXH40z32URLAO9udw9tGqEfiSq
e64o6mdizgfAfyjof2LJ233kxwNomNKMdPpUxFXA8hEYav/sAcRrEOpZzUlj77ZC
YrCrwhBc1dxFukac8TTv7fZZj3I3uv48Vs01AnZn+/o=
`protect END_PROTECTED
