`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d19WQ1AvyFmKw6RHbn4Fc237BYKLKJtzS+vtz9D60qFO2qGuolNo++vbjjAryhQt
NWOyOf7dfAZKgW6/2BSIvJVfEyhi0etd35aDmoZ+wGdkyr7oT6QiBKihHHYBYmME
yD47Usp5GFygh6JcJuYm/IFELs/CNw6yuT9eeGfLZR+y9NBMe9m0zqU39AejaaE7
wkmMhdlROZMaROSTscjxQxpnM3OMSWl2AJ3EuB1cZ2AaO7+IOZT4UxlpK5S4QBbj
lE+hgjUEgIox+TlzvxdNJwhH64DOsOxDOYG4cWdAQgc973ZO/qWUqHTEPoOA4WTI
agoYhbo74KNbGkx8V3tkfx12xeaDN3BDNriO2GxU8Uh87BHADXIp+fdU+9vp6w+M
Y53YAFnObYd3xO7ceRFz8sot9RTKlE/m4Uoi/Lw6Me9XzOLWHR9kMnvdHJMHFKWG
jYla+JJPZAY9s5i4hMu53RpxowMcIc0lBy1iQSrxniZdfkFPuqz9kE0hSCyf4fHo
me1YqVEYD9+K+j/6v8sufG7FkwuQLRv9YvJpWcJaUTG+cCV6LZMhuERqEL1HukB7
cc7d0oALHMYPygQIOBsak1a8nXeZCTPrK6ArluMrOWLJlLp+w1UIjpzGANFolhz7
et8jLGICmJeFHvHo6mL0Q2glP78TRYnjDiyvTuhKxCm0K/+hp/b4HWlacVEesGfn
PI4JIERzbb7TzQGFWkP54kmSR3KVGF/5A8snOdCdlrFYpX3AjeIIZ3E/poNKyIk5
3WPtiMB4mldQt1u2kozaKZmSHSePHhDWr9aSll4qwCQJMJaU7KPSldCx/yOe7YgF
Lnx037YbKuAcDVG1OVSc248DgibKWZ2joSlDOiQK7PDRLSVHrfnypvg6gxu4isF6
`protect END_PROTECTED
