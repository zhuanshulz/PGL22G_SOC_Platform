`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMDDJCKDpmFxt6YQVW7wK+YmOvOErrgMV29ASOCgot06Ke5XnyDQFFmYlr4oF8Yo
1ehRn+9Oa7FvUZGM1wMTnex+kO4DeDl4hSHs0QF1Obp1gA5TX0MdPBmM3YIyV+hO
DU2F/qQs5r1hBLJfuXVFOQlEkd9dwlNw21KfdBqpguzM/oW3fEuu0WZ84KX3/QAC
+P5ZfV8KArYGYe7N9BPnF3pTsUZ+YD/npmcS9pQvfjfbPiE91b9CaUVv48Vl1got
MqgjgetNcpcghhf2kH3XK0M4Z2TVglHSaw2fiD1RW+bmi902w4H1O6v8HbbLoOU/
MiTi0s59biWLOgK1Btat5l0oiw+r60ptODuvClshV2hPyNSEPoLo0j4uleaAT7v8
kchWPgdy5EZadLKZXvtxeWDiD7WpsuFKw+cZ/d81cD1braO+3e6iZznpbMvo+npa
CLvsJkNBUIK+dqMqPIiN9Not1FLsqSSGGfwJKyPw6RAfZ3kBledJFTodef2LyaJe
`protect END_PROTECTED
