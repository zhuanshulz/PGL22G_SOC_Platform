`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZlPNnfG5s74/qvbiZnZJVWomLQE50HYh1qA/zSF4f7eHGN9tsZQw0CP//fStRLYX
KkF5xQsy5JEFGv6LODE+KOMp6ru3cwRzhPyMMEKJnWIgur4pf1wiDqsVJhFXU8vt
Y1DRlLwbSb53Wr6G5b2zsgbsZxSNyTeZJGMHCip8Ude+KqvrYUC94LlAAdBsoDi/
RsOJAEw19ymOdhCezM26vYGHRTMi3E9TfhW9/L35DwI01WqL9W4rluPPUYKbUf5K
BzYM+AGWTIP2JlVbhW9MSWHzHwJe2FbyJnLG0SSa4wELVrH7KgrAucak7jFbH35S
L3S3qafZOSifRT4uLBPSi5lrwBhE447ehZ/euKb+/bssxCvlqcm110orNaORZcbU
3U0LlMLcPFtAXDDjo9cwmXBG8nKJzPSb24uXcDReQf09JDKLWK7ICclg72uCFHcA
pL58KLBN5M84DBHpFiGLXw+25lx3oamgLX2m+Ey6Nvi3xGq1yOLOsjLL27+zJ/li
z+UGQhGoCfxebl1hKaXwGOwmq37HGseryv22fZ7zYqfSBa7yx8mzIpLbyqoriUn7
AV5Ga7FZdI+eAge+PjITnAOU8lHrkc1nOQdGHbT/GMDsCaI/YOFLVoVRwq+sw+JI
X7vo8+4GARcyESoEXZJZpAp/4OnALI19Y8ERRdHZULgVCt7weN1PExNM6PAUwTEP
7Et/7SjgPM/pEcd8jy72TnzLYLtO7rYrAi8EIPRQy7dvMiM04NJvb0dLc4jlaBbn
pmHdcOT4QxJpky/Kg2C9uapGPwnpTJJKuDPjS7WQpLkk2z0Q3JXMBOj2IkYMhXuC
L3YIPYW2VOru6OQ0H2vQTsJK95rdEUQoPWw8SgcvtaLN6HzTMgzmT+1P9CRAmbYp
HZrQfIQlKKQms4Tp7Sw8RHmInnwzMQuuw7nhCSSMp90cB/UE2gCG9YsWgIO3qH06
MEN2OuAehPQXoUK1L68uloaCd2q4yEoXW5QtgiMTBBQ8zA0QGQvR+pglKR2YqSPT
QfbS+hxyfeks4TIXjiLFaTZ+jLddDi5JRwPcxEhPRPzhcOVDIVp5rZxiAit4Kg5Y
PUk5hLlJ34LApUEl6TKDj11sYjUZQ1SDe2GN0dm2Mef+Q3pa1yZ/it41wvDemwqi
sWQTX4s+BRYle0muBNGwATPrITadFUWtbtDNzZrXFV+ZfxWmIbxKuAwdQ1GEm/5y
o7EYvgygDUPm5wt6RhRnu15iZuxYCCjdDNWXlciSVPkrsyrP0mHUgeqPH9IxDxJH
xAFDP2P2aM5UwlkUDR7qLKnFP44H9d0mxeDHm8p5c6/89M3+Bog0FLotq29bxNbM
x7QdNkqGfsiGg67EX1gb6A==
`protect END_PROTECTED
