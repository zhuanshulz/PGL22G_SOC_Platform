`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OGe86H5a1O0k1+gCExc488PL4TFY3u0eEfhvav55cLNozgIoeb2Dwo/a7UPsjD/Z
0DWgn1hbt4wWAyYFV3C9PUDdCJpJiHzOow89Z6XS9W5OJfrOOFczuHUbWJ328eFJ
UbTV+bLOynHRszC+tAZtkawE//Vz9JsY8AWhxKXr4pdPjcAwVhR+Vl/2cdj13IIA
RF1zW4aOo6Iz96OKw7bOLaJtKXY6kXG0FNY6EFpmc7Bc46HZj+Az3uzG9aVc0NIy
1e5VEJmqcyyWIA1DnGIkkjDxx4DBL9gfTd43YntfAlo9/8ze8u/ARz/OLtr+vIZr
5ikd/Uqn0n2DEf90KW0UCiuNg8C4pYmerq3eaqBRYKckJEBx/lgCpIz/NCWRJoRg
Yk2IEycPtyATbW/v0k+kGDWhrhp3JHrQcADUuueUsHem1uSxUTq6AbJLjNuZk8GB
9aeoUocTivIsiHLNmzhx/Ak8WW80a7yhuPZXVNofbYAkHkFpA9LOcvcWcy3c0bRa
sWL7FpgvTxRPcR4JRpaHsoukZMMazUZFd9sJQMP5ATj6FmnqE9O+EC9C7grAyJMB
y+9fYgkgeh/kMY1L8fZajd2tnp8pzDAtzQ3093iDiQRKuHL0742jOR9eqPIPcHqA
Iwx8uCsJ+lB+JDUwwozIW2uLBsNwmiGsPuokUFZBQNVMUzTiPIgk/o07ih4UfPFg
g2eZNuMkI/WvvSFH+0csWf4jHyxbSVdlq02Z4GnIeDB7ZHiiY0eayWP7jY94iQAL
ClXVoLj7Vwwg25Wxp0uJJ7kCiQ+x9/AaAHQV/F5udAh7Jhei0IYt5pF449IuhJ+7
hLUWzrmwVmpNYlHHIadRUTkLWdvV0eAuIi3jI67xXdWAEMn3ROfUrzz/Tv4yzcuM
jnxWtbo7pxNJ3dxXrV7uj8hn6N0RyhrfQ6Zau98oeIczgcy0dWpl3mZmP1SyWYpM
UI/Rub69YDOVyMbTuneS2Z5hNWcii0RQBrQ3P28cRpjdolA6DtCntCgOEbcDhyyd
`protect END_PROTECTED
