`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P/eLOocPQkX4mrEKkzqCJgbg4JHsSrxDTwagh8noAST+2fDTd/aUEdA8e9lzAeiO
iolcmFccV6bMNjQ5lpPpmO7uW72yR/+JXR7NUZqycJS7IEhS4QUN6qMwDCkNFfZ/
MZ97wUfoyMMypvHollETf4nOOi++HQwLgkQOZnB5CUBSZeJfDsJ7GcvUtinOep79
1qED0OqwFnKckOKTUykWWGiXCmUXQ2seXEu18VPZ3//V6t0BS56vIjifXWrR7JWT
ehPUqMrmR2GRuxbZNc+hgf4lfF8eV5hwV+bObStmFs7lt3/fTxpIJPOLP3TjM7WC
M8UWPQiBE90OhZ51eQB1Q+DmORrMy22MEBLAK1xp/S6eRFcF3lGUX+yAyVtApOvh
rd4nk1xlQkGbzPREYvMEhaudC46IKweRkXY3LOV76t/gb0Ia4AaxfwJm/taYcABj
PQZDCkJUBanzj8iL8/mC28aDjVYmcQQ2ZNboIpJRf2j7Td9aYRoy4udZii670bQs
pKCjhY/2fekVJ0tHVV7ukk1/61s27CJRhokZza/2Q37S0rSDC4A0p1LcxMGCB80a
rQ4UTihlmWuvQQN3BdvwxX3YV81QGZjBI4riFoSF7CJBs2vi2n/duu8ym/2aTEex
aHvlPBYwi27yKvdxsM3KJ4YPSWSityn7Pttzax7ZChiqsMMkdgYH9P9F1yYb4d/e
q3Bo8XFt+arNjOWygOvsHYoMFeukFGdRyiVhIge3EpLUWk72LLmTo34e7KwsU76N
9Mryvp1Vv0n1tYRdOXF/iQs9cxkksNhL9IUgCkx3NCcxYgoVclbC08MXRWiRUoz6
3IRQo0o2b/WksHXCG0f3RCAJ8KmLunfsYGJlAPjwDAiEboibTY6j1FyFktkrI1ep
aNGl4+QabIDIRfD7cgo8E4UoubxTs/BgziUVYjpH6df+q8Bc7Qw6sPRfR0hnMxPR
sBLB5rfgHIjbAcXUqwPOpurVpoyqS+++VTrHPkkdFajpxaU387JaW2KLCpM7Qwa2
rpQlJesSHrYF6odO0yBZvZ3Cv0sv11wspPs4r0zE0MhcUqibVJ9NvmdFrG3zQitb
hnl5BH9H0lQEOXluOXezaxbG0m+lsW5POhuJRbkahXoRc5FQi6PuOL+R59nkAKON
T0w/ycFTQaVNOwzUKkRCnKwson3NXqZ8RHiglS3vxzPn+kb8PNeskSote2tSNbyO
/zZhsQzjyp6C3s24ohu4fvYTa9vRMKjG66uJdmwk6SkVzrzqjsySy+CUwJWNRQ+4
/YB6pS/bfogD4JfnQ2nO9cRm4mHawjVinEJNSqKWhJlI1u84TI81zC4IeGm+R5Ep
TbhNCM6KxP8lS+UuaWaZl7GyKWbxoNAwlgJhGq8DdG1YwiTjweNBdBhiwLHxfRrU
wzKLXr9J6hhA1R1oOEpt775ie8i0Z45yzJJprYQELieqWzQx6gdfBxpFENeDRvuf
MAkQzrUiVb7aZ+04mnPasUTqcF2zhmbXQSpSOVptfwq6SjMHsjz2ahTMnt/r80RJ
KLxMCzjBiNv3Zdf8Dr4UKhzcHLEoluM/KtGW1UPqmP9XPgde6TaOoGi0Cae3HUTC
iWcZn2tUwgEUOr1OfzP56uml4itbz3aA4W3x3h+eTdIAX/W+CtZMSb4H9siE1EG/
0He+QTefedC1dDdoEchL23TarXbwJDKnaFccEpn2l/fEpz/iubBGXJUzK34XbPtL
0tzrGrPvkFcYOq/19YNrLQnPqJIS8QQ3s+Gyb10VaUpod8knRroC8zlJizTQR032
OH2ZpFq8LQDftglNPX+4i6SLgfAyuRMl8/fkEoXLh06F0ZmXSnrHXco/8zw5I0i9
RljDAhS4datGMXAeNdcoJQyDGtH8/OqhXYjnJQbKO6Ba6hgNutQUa2hb6rz62GR2
6gPoFMQsH/c1+kMAc3l6UOJjmbCEeVxjvp4UwVuQkXanHaReoRXrpqRqtuGnrZNp
vOWiwX+vksC6wxe5DC4dLolb3f8lJLiNK6Lb06Cf463SMAcpDmq5BNzZnH2Kw8CS
kcQCR9RSbdxkul4DjprwK31txuwHgd6btC5FNeA/G2339idUTRK9WqPbT3QTcnpw
rdqxnv6C77d7Eh15ODEm0vUUOoFBA3ovYaw5N6impnL1/QmliWnMHa7lcGz+Clg2
mV+Zwd+zEXrhig5uMy8SxQ0nWQcl5VYjDc8+Wv+FIV7DQW7GlaNYwnHYs4ZYeAQa
f5RMR7YDSLdSebU+Ht8801a4GIa+wMbvjyIqrY7AEWOPrzvbnRetZat6Ofy2Qkmr
Db3GWMDdq7jl0eZEnnRQVBgfXz5lwfBMkEM9hvi5r0Ic/uxayqxeWth5YX4Jy67D
1DMP9jiUQc9RMgZXGRZc/nTHXVMBtY8wgz23brzKaDNdoCQq6PGiqeWs7DjIXxty
5QfjsegMJIX48Lo70nCCHdXpqR5MAMug99TwjPPzU7aI9UNwGibfxQRqrYGHXCoA
L0f+FNWRCtZ3nXp05AuoZNmkk1qu2OVx4ONPVQjLksPW7NqyqpMD7pnNdiPATgvO
AQVxre7y9JJt7PpHachwL2RXVbBrdpcUX1srmDK8VQeb6W3adsKbhV5cf9/MLYu5
8/eXJ+GqpV1MGhflUUc20Q0VlH4meep+osm2u24rL7utsTEoH2HEGzvmYvhFbTbt
2Co+bcX4yGzW9lMJr3rf8ktqI2pBlg23VhX8oBHxuHcTB72ntP0Ay7EE8BWbr7AZ
zw3dEE/qpiitM3at2OoXZI7lUbI+HUFDJjucba6Cwux8uY5/nVnjm0ULn8cDVHQL
/bOA+0n2j83aOu9bIiE/EdEhgs112VN5cUOI6BO8Wi54RA+htWNMIG5OVrDdzkE1
WjIBFytnoWUabtGq4OsourRwflZlu1reGVls/UMq7V+s7tRd5Mc5wgqAch9TCx8r
8E30iQ7zSgd5+Q0UqQbPE+7t2B7dQLXUgyXN+nSax8+RByRckbzsmtdoW7eUZ1rJ
CroK2Cht+VMiaVDXLy5KEuhupoGrx3rzEy6S9ZAsAsT4/0ZM/kzSelPmHOkdyG73
L8Opld2Wh2aR9VAr1HfcQg==
`protect END_PROTECTED
