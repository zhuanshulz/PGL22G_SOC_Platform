`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dL/EFocvW5V4ehKKYSCwa2EbIr6/YQycyqdakLP2Xy4fSnsOIPW/3f+Om0MXDXrV
gcba98QNJeR1Gb8jaOGlwU8aRjo300/7z9u3+qTrki/xBYBE5fF92NJVSEdQT+Ys
b52q+ZCtmkvxATh6IvUO97pAnXQ6bmxHTj14ofIGdIVocHIQuDN5CrljNJ/cDtBE
ebUfarTd2Z3n5J2k4QwbU9QHewF9DiJowwTLm1mOX4f0dQr4HXaRY+KbISkMWvnj
QzIodJlvVcie/5QyZNfiH5W59yWkD9SgluvNe8LQkEH/+AG1gDFkCdsYaVmd0xzb
q6BtIMY3jIBq/76YHuGr3rLabYT69JVF87rqtBmuujIQOv7TC94VsTKswYUvh7XP
PSfoU9ukeYIecJR4t8QzfWoPieZ1WRRXX0wCbjqppllDjTi78jkyHVsuXAiVMncj
RJtmX+EqfpXlrNZ1MmmxZdpWJRtvtiR0EA8jQUFDmd9UI57rOBDv0k9FYAUmhWyR
7WyrBEIjxGwm9+jms3MCPMAi8Cakpj0r6V9uYpIUmVpTmtkLX4/NSdzyON6ILEi1
3oglv5KJcQnYAXu1H3PXrIjYn/PHp6onKCeY4cZ8804R9/dMDczB+kToHeY8Zch+
r8SJF09jCnYCogTrawd3hmBIrNB7tCGRQWW0m2N0eJ22cKFUW88jQBtnuYC+KOJG
zEh8DofbtnI2qUgfLKH7iKjadWUftp3TLTyKJM4L/pSoOWM7iR55e0WigBWl42Je
js6ZVCtPWfiaj0NjaKtBqrDS3GF6CaJmjzDgfkDo4ZS5H6Aw3J1WNJzYR0Q2Keai
DLQFQXFicpLgGJcq3RMgknCmhCOyKLoQhy2X1DAykihmJU0262R4E3gZrNFCdoEt
rAXe3O5SqPLUO0RgSzmjag==
`protect END_PROTECTED
