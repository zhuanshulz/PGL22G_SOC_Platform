`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3lphPZ3EeCCKyQ3diGs3kKPJ6HsoTxxQNWlZ51FfNnCruT9jYc90lqXPRKKcfSL
Lyw5lQ/I4bSRRUDpilKMtfBV1Ku8PLmbLzw7LifJS9RXrWy/5UfMPPX+KaKYXO7Z
Ei4ucswD51Muc6R8t+Gh32qcn0RzWpoOZ+Bj6q4ScORBc1ZQV4YlcrOHS6F5dKEG
6yPmeMnS4imxFgRabe9KODVy6w0aOds+229l6qAad06Rpn+F5lD9fJJe9th1Zssx
P6xpm36Hxc6qhS8zMYFwmlDJksP00tlAGE2ksRcmmo4f+oSQwRd041bMqALVhSDJ
aKOuQLrEV0qu058OK5uI2eJuC6SP2neB7LmXPuoZ0x+dq4SWPIXAmoFxBZAVp4CV
hmpBWeyvZj9nBw2nL2oMJ2RmLRc6ItKHVmtTMeJMO+/xfVz+3iOndXQTiTT5gLzF
kb4AhzIL+w9CSg6Se8GoPhACmee+V1U4QFosM8M6ojYBWSCVVvIIp8fBIJFxn8eD
/qbHA83s3PgFBUataujyN+8bBA+iihyPH67/Dt3t8Iwi5N++XQa4CodgQERA7TfU
bfuNOIlF9UjVHD6FvUnZ6Cz6JWMGVoR38mVcMR7ji7iiGllx+KK0610+zyZ9lUVP
5g0UQlk0rZw/Wt2KhUeOBVUSugad6Kyp2ma/uBEyVrCmXGKmtUmJTcirawfPYATm
vYdSxY67bWBuq1lqmEM1rHhvdVqUI+IIrvdLN49zwfGWGqyGSsNG9LhsSkwbjXcR
xV0+BbyO4rg4xVLRSgMrUw8QmAtW4yo+FWcClY3EZxi6GTbSHkYU/Ez/HTsDEpOj
OIuzPEM7LBt/Zgn3Wwe8mg+gi2Bz9ze828HwcQUBI2o=
`protect END_PROTECTED
