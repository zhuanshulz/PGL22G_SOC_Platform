`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NTphDPvU/kDligVaXp56pER46a+uMf9o6zRr7NWp8AHPk7/EgE6JPYckl39VIO2n
q8X/xkF5XfkT71kabZeyjX9dXZ6WNwJAbcyGmL37kdJx6dap5GuD4KO0E0V4zKYY
Zo3vhGHY3lTpT9zroXDQOv2xoonHt79GyEK6rmcFwznw4mJQ8rnEvWw0p2zWEAOV
aTVoyDmW5og8bnLVG7Oz3LoSD/K1WhWe5Ibd5VqL6v2M+xmbdJ2Y1SIs3M9/U0J8
3T3OC8sNkeJjug+oVG/ON7fIByY03IMzKeufHfoAy4GLc4gejxyOMT4H6BWGNU2M
nK0t8v/HpjHNirsfIB7DCeXCzlapRaFUoLZEOYqT85yRVoGcSgrEwI+RYMLpOkdt
XIsAd98iCzEWKNqtGY6+0CBGOs9QOPy3OYl55xmHDHuIpbkR4Q2pM5yqEojHnsdm
qYXTeENb+e5o4k8oOQbJDAqjVECH2tKWWP0m+45UoHJ0vQsOBU3sLSkcSlBsMstQ
/HvR2kbnKiwftaLeg8VgOnfPj1xlgQI7s61TCpMr53NReoPnN0zDqEl/B3I/uRHs
W070j5BX+WmH+2LvqG5IeIiMs476Aps/uZN60ciL/ePkwDk63VFI5z4AuskK/Jb0
9G2C7bEjsHIdIIAdI/mX+1Yf7f5HgjvebJ7ZcZeF2NpY2Yil8fq+SFD+CF3FksrM
EnJwlHVoDqtt4AOk2RjsQMT/K6tDKrIm9LMSB48V8HnAkKBmw3D31rEmaruAlSmz
Llx7VbueDyw1iMChfBxtu0XlpKC087+j4wXfOn4uxOvf/LDLJw5J1l7vOr3bwmOR
qsGnscluFXR2LA931BKYoy9D2TJQmwbIqK6atviCDcrpFB3lpzTnhDL7SQPVDR31
UDFgQnuiKCGniGBn6ytCBuhn/QP6nNWvmFXgAhgg758/XEICh5Xn9ToWQIH+UmIi
KrmoY7CI/eQIyDpwnDSJu7ZIGu8cJsQZmFpPffRtX1a/02QZvlJxn6rLbx+Ykaoz
GG4LQIFskq7tuPBSCn+hhh/J/mpGH0N3J0p501wWNDFJ4EW3+0CQQUCG5o1loEvn
0r6g4p77wKhJb/luEqmn+TvnCcHT04a3Ghqn09yq86j1vnaQBfu4gciGObXU5tFf
0TJDO0O9W2FEzBIIVOZgDmZxb9l+CY/AFUOylZKKwAgYrVnHJ3vfjDh932aeKse4
YEhG7LkTfDyB/0BHt5p3rysYx7xvM+TXOoawoVIKCrc8PtjO7xbNXNBoiS26mNJm
ALf5/0amRRQ/rfl58o3QzKG9mwA+90ssJfDFX7num6ts9RJqHFnhI2AXvDh/wi1x
eO714Nsv1j16GfTJDttC3OENJD4GEVAslZVZwzRaDtbUwj/esXh0tZ7B/eJVbiGM
GvHSyU+RHikFwfFcRC4+/35akg0nkCPUCniEtBtxq8xff5Ic96akVzHAPRNDs/4n
NQB3qJ57Ll9ow1dQkr7L7tr9Rvs1oT5VlPoZ21Xb1cTbNwZVk9HQCr5F541icYG6
p1nb9ONgRHUiL6fVC4RD75Tk/n0NVZbXLpKWUF6pTAfsfRLLP2jVq6pyetOZrbPe
ilcgiUkOPBKUV6WwPGuw91J57qV9Rw79CamI8S+0zIBENGo8ZDzAOnOvuZhnHQ+O
2/47zc5AGLi68Cemdcj34ZoUAK35H8m0DqtcEzLFr1vM97SVDOCkehLNF/kwqFEg
OAZ5cJ4eekXUE8dRjzKP1yEx9xTwzIF+FKOyE8xqxDyQXh+Pq23L8onmK30b8vwL
bER+H1aUiyS13LSKYjzD4aRZvt8/n1ByOnZZiKert1uMdLVazF34yXosnFhcGDcj
c2JZjHcaQxsXOfUsTbX4YKook/+v2LZ4z/KwpTETAVo4ixNgJjDUyhQcvMB7CZ+J
NHelhsTqbvhAZRcRWJpARU6Fh6cHpthcgnG/j8L3TWsbOg1Gw6Mmb+4mWJiJ752f
NkXwGW6QlN+tHu0aPKZ7Z5+FHSmGv4UJoOC4r9Lcw2uXrW6kmDYvnpbSQHRh65ZM
AVMzDFnz5/ZikHbKQpHaRuNO4KLfeLlgitJH3cbsnExA5qYdn5qf0QzOfgi1ST/R
DidxAEUcrO0SpVLGJ8685SLjrjC6U1V+Qgj7RhMTw8vV4ibSQ1WtU3E1jo1rFNvj
TSEKWTMAq0fKVe0zX3GXjS2krC7/GmqfYEZRbQBq5+JEdZ2E+g8QX0cXhg00yVhG
HNUh2dyf4sKAcplOxUnhvvTXWmZ3Lj1Qmoow9wLdr8mi7LvSQK3s3cT6QgdAubA8
lhaX9cJi238E3cGcenXrGYVhxmgp54DM1oar4tBYcup9QOslLsKIBpK1Y0IUdiUg
riqQV4W4RRn36e5T9CIlrYFPSeyDKKJwnLsrBYFVDd4EvCqUR5atkPyI3PmuBAJa
5OO4dm6IfSUmH3mYCQzPZO9wOldYOhlds29T0YPnzbtESe6+ctZhE5eyvJ/qa3ZC
augnbJTUaBvLjBiMQpfe9HNNjfLxXN/lWnhCpPK1+ORyzJzgITBWzJof324xix9X
xH8p/ZHMLK+XmH2J/28eTOENGqB5mr0v23drJRQpwjRtJIscjpRkvCONJQDN1eux
bO3qis2fTXXOycyRYgSzbjY3kYrT0teVU62QMNRZxTu9AiCynRU4gL1/yKHuYbHz
GlGrKCrt7h5/Zq7AoFVUiR2tBmCiANwDMGBciAT1j0WXw1yrXFsEnAuDkYAiXr4K
vxSD17MN2k+TKQVu0a/lhjayecUc17ASrCuQbPHYGeyOp9xkNhwVy+EWN5Rm8RvF
PM3mkLTkTh2icnTvXREJsrgCR7AJr/44bW2ywoYDG3sNDrB77eBheBc/vSjUcFFU
ODokAaCV+foXeG5KPKW2mLd/poeo/BtKQ/pcQN1wxqjUFexkU6IoOuDaVPmSnEYO
P/Ms+RDVnQ8qBMs7gf0urSCZtCBntrnwfCSAkwQy83SjjCgMbWwsaaNbREo5l53L
s/3O+GJhV1+6WMYc5lkOyiEF8KaR9xdflxZD0VkPoZzP1CqEHOvX49OR10/E8ERC
BsztrbfoEbDOCZssf3EIn+AV3A73YqRxxEjws9tVDPD77/3Mop8ajU8eBQV5YLOs
2g9L35jFslWw/wKbb88a9HNTe1tTk8uCXgXxa4Za9RFITqZkXfuzUbZyEVDBVBnm
DVwm9Qu6VliFlXPk9SRwS8epVTdc/zXPv/5Of+RvQDyp3cefJALbtdHQPwzrft5t
KbrkGpfQiJDQkWoSABnp8nMwe4amwdnVQuvflahbEM5ugVRBsRWXBqZfQHsl5K74
Q2cHQCfxg1+5VrAndU0HbDgq5Ky0ix7S6HrAf/HYl8A+JZZ+uEjxeq+qMwZnQ541
WlfYVJ3J91h698NgjhoLfQ0K+Z9PSO4Xxt2BzWvbyRI1BHmNNg0KJyPVbYh7zM0Q
KEaQaqDAIexL6bcIWzPSPgShO8x63jqr2IWmdUMIap13KrGE4ZBUogC2HROb6lHv
ik8xctjwoYLLtoW76lCQOG9Fv0i5PcJAVOOmHUy4KDGeSIVODuMgUpTCACAQNWXr
9eNamTMciv6zfVwZbjc3Jbl4Zr+PUt4iDEv14+E5OqX4YE4x996EJ/7Fdr2+3TGW
hRS4KDNtteocKXA19091QQIwQE2mkyNdiVzBOLPuYohJ+HM3dSqBHPd+gxKRyh4M
KkztWBFNYw4lIywxPXZGrUxQqlJrtnVonEPMZsBcBdCRPXPS41ek+M7/dSjFZet4
JsXiVFF0A3EopicuEaMP1QZaG8EEsoTSDGyTNXjKM2bS7nX6ben6XLEe1ccgme+x
9RIkJdK93A48L4lbRYoJa6lprdHZ/VTec4A0+JiOgsVUdaI5XZaMFHEfXBjD7eP9
dzCobT3wyvwY5y2efyc57KRqZSf4+vjP7eOrAzmalpu3eZiF6/XA4VdTVoE0AYao
wOVwmXCjK1Jc27vC1V4YMcD5BC4/AyDrueYXqab+0hU/yAt8Bm50v7rHglnkQbRx
ZD/eLQBNz7buYUs+PuYafaxxPdpMjcM6KYxkIYT6kT2kERnaRKD8hgOnCKmpZqhD
4NYpWKLE0pnAwQ/1/1cAW154KnP89GY8USnvbJ4F7VtZFc46FntQEKLtSzRkLHek
jcLXXS0r3zsrND8wBPtmpBwFGkLwv9pnfq+CX9uI/IogJHGpLGUTjDRvT1wgKsSD
vdYGRDhPrGNXrXsTeQTX8SUGa1NHCverRj8IMrHmSP6qN3cxhYN5QdLCER/DNrgA
tjYQHVLBeJjZAaDJTII21vqLxvkq/e1oMQBpjEteNr0NDZH2IKgBFGqlK/nrsQlJ
4v1ABOKlfgZRZk9oNieu3OTrLJ/ySeunevKieKqMhaCyDMDIIsSkygpTuDI/WbKH
w4fu2z83LmHnGCOUH+PAgAjAt+v0UrnuJrASngJDMo7fT1E3RTL1AHS84mcuKLOC
MfzPpsJOZGzOjFUInGsSNlANqYAmtHCX6dhXI2Lz/jMZfl67/SY4oq776/VI2Asn
kUfPRkr9fzEHJf6ZDDeDfK0fSy6PkhcTGb8RiiHZGSXgfQ2iMiSxon7yx9z8KA9v
2HfT/DpBdOlJvEKEjxTxxYOV6Tw3a5yEEZINmtKxnOM4DWa+R2xjIUlzcxLEu+nm
yVkFQoaCfRvfYZCmOx2BFpMWXb+UGsPSWlR4bb+YHzPZK6QI4WCFsGXOnb5DIGyO
e2ZMMFZTSeXyHEjHxuBjNsWcT/NnhxX1xTvvtk81GkNMQfkm1k0UYwABNxFNiMp3
pOmOvHJXv+W7fq0n1pOHN40d0hyBgcrmYp/h9rhduAZgGxCYp8xUWsZjIMkAbflX
fg9UPD9KAZYI7JfCe3ZiKSk9nFLCGz3n+HcTz097H0GDCrvCEkZLVClU9b4jja4S
//kUSyaIN62LI312lNqY0UJn9ZTJibNLsbAty8MxLOJ/CgEgYBOTr8o4qBsdzz7k
G4CuSKukvfMRpft4DCcfX7KTEoa6UFq7GAsfvdSqYKtfERqryD6NuNIvgbkSacMe
0OfqgqswRos5VS3Ul0/yXYC9chLeSk5w/dl2xyyItxZiH0TdsFwG2IWiHwoIBORJ
5ACuhqFN5A5X8nXlEqb9U6S/nsjDb8+PFlh9cWmH8bgYU4tN201bfaKnLzPn5XYl
Sr+8BBDW2+HpnbI3QK0FY8LronHkygVKz99q5pwmmgACxjbIWrAlGUlzc4tIEr7b
P11VJBGb7SNoRJxH5CU3YpXa5zxuSEZPZtRcxsjarVBBj6ZRpBbELxMqyIOhNShe
ey7Xw7p3lmaO3arOrWzuByMJmPcqE8iRHuWZHhgga7g2GDHlliaFZ9jMUXupdCAT
oQJipzXlEcum3sZii5X2Zhab+HyYn9b0N2d5EdC98ivoH9c9zc8tkSWPdNtzrrI9
hVpMn/y48RlINFDWt6LQSRe+izGhN3LWvfRAMJE4hx7LKiE6AURFflMvHMxRFSlZ
gEJbQn8QMF1R9lpV6GZoUvgk05bKqU0hN0vEKHdJ+PukW0xJmz/Y0xRQdHi8hk/I
7wUyZb76R7hErAnLVX2PvL7Gd0PeeU2h1BDUGBtQOUhm+xy/9ePJcp9OdhhNMvrV
y4uAiFDGo56E2yfLx87u/MpGMfkyFAwnavvjLR7gHke/+Dp5Lb63Ll6Lw2ecATEE
H/I5LamC2ODhx3haZY78o5gzM7d3etRhgk5EeVPQ5HBl6nUat6f5Ggcv3xSNivWb
/nVxNTq2Qozo8xCgEuFML3gOUlVwYfqVJXoeR7PvrmPPdZOVblWtUHdZf63FbuIy
+XN0ERyMGbSXxnXizostq2HLOjpwQ+Jhz/7W4S4Pa7+dXhXCdz4c+h8D+/3q1A7N
wBQ+3tYcBCECxKwgTW5AdCbC85U4IVCB5MWhko5btLXlLD//XhfjuTh68d5eqwT7
MUs0FeSSQwgjRjT+fmshZjX0BYSuvl/stScIZMM0dvmEBMKJRi1lwaUgRggkyz9o
kSuUEVlJYcluJrM8rMlxHGXMRFDx8lS18A7e1oBGWAFWkgxtcfI0uOyRD0JOEWt3
/n76Ks35A33u6BKYvPCr52JzSS8K68KJCJ9J0h3Gz57uDYGV0XCo1+bTYGyo5e/Z
2w3wmiCLVESwDjYFLTO9PLWArJ5tDSxFt3VC4VfaohPLAi2a2u8LF4zV18kFUTZu
dM7zgBSPigV0SWADGC686T4gkkj12jz6Jt0NpuGNTz5OMJxNHJD0tSyRqzuC6lt6
UfTKwp9l+PzjHn85S6pGbnM17cDrcituvk317G2rmYD2G1RUbERYZfwD2mvxgXGY
bkK92ZKshNvdtjNimdfDvm0p4PN8j6/V5ChOpG/7tAbYFok5fAvIs8omD9iVB9fs
h0IPkeXogKSKrUoIcP4NxzrSdrrrDyKPP+yQus1A7K9PcQesaLij3q9iZqKSDjPx
oEpubAL6FPfsmD6oPeZwtu//NEZoIm9ZsmxB005b+yCbdtl6nNwbu8JDz9G8xC/x
SQz5NgrsON7c5d89gRQeue4GWX0DDOJoxLB9ilrgtVYkUvSbzo3O6iQ1pm+sqDum
AkXR5juPmQZ6/Srs3d37j1p4uTolI4l6PkNIAQSMvkzjC50ATdGd5f6KyIIqOcnz
DpBhdT8JJpCJiwbCfZMq9qfwRTBqhgGmBrrhcBD70gyvo+KfXDwn2h3V7CLz3Ddj
KpiQwawKjWuuhV+7G7cEUvEJokigXVQQkD9hgUgRm0AJt4InkceUG7Za34J4Zq0w
TV3HFS1t57FtzQ2hl54aOSNSXiKkiqTiRkgOo+520I7k2PlgfwN60lnZui0YWCsU
lhjvUBaVwTKkXaeaarzn7KF+msLc0I2xYBTWdApHNHJ3NsGdlxA6LZRyNcooy97A
RejNW2EEXKNmNlk2zM1FzuqWds7RQlcI8+5dHQUaL+mOFDfPw+enwS6bvoUttW/E
xcUC1rctHN0USTynj6RmrCfYSWijXvoq9wtmH0HleJEMQKPcoNeN6bRtx18SheYO
tj1krrg19Y0HpEnrX9id6OArQO02q9sVLpM06W+ZcyBZi5GF2s8AAa6aXf0tx9I1
2aslfkk9nVNnRh3sZfAtD8FxOCYcvSBU0Tit0MA6k9oKIvXXpi21WKC4sKLdOrTx
xwcvVaHSroFVpaH0vT2C1Qb++9fSo4BOZRdJrbgh84CHDUlY3WfHHyGKsnGs0oiE
v4gig+PoeZ6DYIRBNlLX9UiMaKNHl05bW94odMaLlFFxawr3sfnqcVTNlnPdS84C
dRAROhTvktVDHJpPbtJ9Jy7uG1FrQ+b83YpWS2uZtPIc1ZiKxXj9Xj1IlEbwMK9v
oWrgVC1t81pdfiZILNq+LfjN1JhgcuORM2HzyEz0PGhDZS9HnEOFFqjfWIlDddpY
6oHuRkeFWaDaR5pyykv7VDDAs6gr7rRFPqgCDIOib5o5/I1K5r1eolPmG2DYwQvt
IDT28wHy5Km6Ls+r+zpihji4DIz98gUe1k1usmUZMr3DpyHW3tmm0iFRS4nrqm6f
0hUhNg1I0VgVDc4R/CBQTrXhoSvZrPdgpaC3xLBW2OrkhrDl9q1bRQWCbp6fygSg
kjKD2Cl923YjBFmnPdl6K2fjP0Zg1KHnaNrJORtBHMrlWNTDQwUd6Zd4gRPW7LHI
kOdnvDcAOTuGwxbaw6MpPTjxw7JMSxlU9jHjEjEowopEyVxVi4cUosAspB93HYG6
BnJnCBvTEWmnmvZj0MKm/p5VYz8nVHLwo5slf0zgVoSgkNeN0bkUlbNO0JsCTRzu
QPvMFEOfAYUnb1F3rSgrlGxMUxfETkIJZWG2hu6zFVpsVV+wTxoTTxQCL4bWKJ50
VQ+5GWSv4uzb/FVtH2DD65VEICt4/iRZm+5z+j6O5HcydOHnv/fFi4XQQ0Oxkaad
hGYACwmhGusITx08/cf3/zqjUDe2G3is6E/+AjWWk0E6DzL8KgUCFwmO19yM4L/h
iSpAjfqMAuhic71FA608k0tXZRnoXy9c7f5bECaTN5nP+x3OW51qKPYIMnNfMfvX
Ww1nc8dXjubq+nlMs9h585SHu0jST9ZCcKVrocmFbXSR7LBGCvnzMPkelp/S7RRQ
tqEjS3d4lUQSqAV/J2ZAtzYrKeq5uNoG3PZ1Y91T7ihrasgNjDbkMarktJIcUvGe
pQOeKeeeDVRm+L/Xjo0E47S9CTW/ppndkI4CMWbcFLT63iQZMPT+rgfz4oBRYoJI
OoWIy/x4+y+oTdB1h1ShhKHEjtYQqd+FFl7y3u3eeqTAFZLD+0XMzq1hqcVzALOx
fzos4kG4OQtuNpHVFpYyGwUmAcWlDNc/dCv8SArC5ZyuNyZhV5RQqrAImwqXxzgo
o4mFR9l6IvGK16rRViIHn/Nrly+TRH0HX+cRk9kyd5vmPggP3tM7qjaTXyeuXDgw
DlZ9Jr6/cw/pJGerfMD0ImDEsOiHLr9YK6QwLLZM3yddKCgOD4AQlACG9kWcGJk/
Zk44JOh4SnRHOZUekOp3DLTREPajgPfwL0wWqAuHBxU=
`protect END_PROTECTED
