`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGEXITrNnw5ZS7OuuEeLh6IhfgTQsjncXPRngZZ/vho6GT1mMy1qptPl/iy18+IQ
+cQCPV/6KLTLvhOZa1AOjIsJTju7qCL9/k2bpcvbNWjc5hbsWr+jKJaIiJZ7RSJc
cYqewsx2OQHqg4BwdZuWSWZOz+B4FuIIaVDlrwmkHm7PBmLvzA6IXREiObMgbVjg
mee3v87utQ4D73FEWQMg95lliucSigeqZsECFKE0DhMbeMouZ56OFZz4GQtNGZ/2
O+Oo/1jerePo1LLWQCgAXCEX9dZ48noxIlsGMshE7eQyz4KEphZYJdTSI28isU/h
tEwp0cupUGYVgE9tY9SCYZJoS+Xa9eQr88BcD0ecGVe6qJ/KeouNyzi4KgId06x7
Xuoa0wz3gxBa/bwGLfjx3XbJzZnC6Uf7WtBy3HesWAw6kX7ZBs9M8YaY2v8/yjDa
cMB1Vnq9D5+rMrMrHuGebo3wv2oQpzTYC7VOOtx01cMj/3lNBnZv2/JEcxn7Prv2
JGlJrMksO154nXmY7S/qHMX7C4dahDGyjxBqq3EH4aXjlRtSj0RQpEc5pMZUdkZ3
Z/6Jxd8G9Zq2yPQ2Gb0d7nsq0Xn87XKPvAoyqDcr7tsd/wN5xVNxragrIrp6mF4o
joZu0TDDSDNA+lZu40vNr/1++cpH9r744vod4XK+93E+kI8IzcKpCKkLbplg+yGE
jhgZ2CErZnIjdHKvqejGuKwCKHCbJlIt8uuHddaB2WJ/gxPGFz6xMbDF3E2a2ZFB
d0voD4tyJ5y1ZEScY2kgFS4ggomJHjAK/s7RdyJ2UFS7IkRNSiU+a5zISB/7T0We
PTElPUlLqMO6bszIG7L6aPdNIxR+q4dzyQ9+4r+K3l9cj8qQDaQzDzIjPJf3kCpO
dfAGnCHU/DFUW6eg9zjBE/OeSCX71GkDaeTojU2HF9k=
`protect END_PROTECTED
