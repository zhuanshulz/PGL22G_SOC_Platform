`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bj4UeWt7rDPCuYcU8SQQi0jQTpVLBJU3LMM1M8pVAtX5cAbxySxWlNT9xNyyaTdy
PDhCoDD7oxaNWC6u3ShZ40LctuPN4V6y9L/eYrWw3oYXaiQUK5UJLreo6nU7cl2N
hx8EAKJfJYAsAwIi9Jz34UOQ07HWiwdQcXUQeEyGaLufoGec8hvRpRjGFzQOd4+j
+laqc+nNVbX9/dg6sMuuKQoRfHG0ud8+BxQaDRgk967zYh3szefUnxUnB38VwhHp
jwikJB9vi/A53+FGxBy5f2pBFKW0YGJphGuO5jOhrLTVXILL1Pgn1X2lrXpHvhUj
txgQ69fB2nmKohLNsGwI5ag8i34ySnlxiTDeN7qu1Q5K0UuEhnZpT+I+9Fxjt6M/
XxrC7G4wPy2Gb+/u11bD1z++W1w04FaVePOWp+7Qd307qS2tV8sEpcpu550wlW5Y
neZpar1TrvuuPytAtYl6bAD5hcAK8gEh5FE8vxwuoErzXnPd6qaglxiuoACE06Q4
2k+WtEVMJIyNqCNirHvsesg/8dgbzUrjI7CBZw3I7+0xUN0hO3KR3QDwYSuClVdL
OJN7HQi9T/FdGGKBst3BPE5xQimRjaqxtdlK1Lactfy0OXOrg4jTowa5v2nDR3iX
eB+MWA2AKTd7wbFFjXQmV5Q1qTt/skzh/IGBAljTtSX1aRujJToOcYM/obR4kupI
gfCJOfXUEViZ/ODoI5eKJtbe2wG6rpTLpZ9bakbQNQyf5Y8zX5yXIRSErjeQ8Mgu
ZYF80ANbEyIVh4mAp12OiA2T+4T5o2R7VLAutbG4dPllVGCDo+/2jfSfWe1ExCw7
ptH5JHK368ZG70JgneLRgMMrJc1UnUKtSU8545xwH1ztiN7yRVbLJFitmHemtUXC
vjsnkcwmz6fMoIdi48DwBA6wunvBwgnmgMAr28FlydHB8RAc+SyKt0sToTlCqoRi
9BheqWumolFQ8sPYIUoYuXuttQNQwLgHELkjr+SvBGkVLeyZ2deQboWvo8TiyoQ6
gczs6SqTGBFUl3lzVzZJJdD0hdYSBbZUJBqBN3p1C/LCTaFvUl8zm6vQw9tj4LbK
2T9G8xPwPlZZMNTo7AG8QrKoBkiBEUTRlULLGAXIufurCVCcEI9AsePuzgiABqOE
AN//wZcdU4L+weQg7yma954+mmMzMQ5m3v0f3Bjd9I5QdKC1TgIcuWXE5aBFKaj0
0SZpMg4pv5mwQWnOP81Az2bWPIbRIO7L3gjYN6Hn95i/vRxBf3dKckLv0hfkI+Kz
zo6nocUuMt9jr52qOPPEOcMmlJR8MfIsIuAiYBm7nGK77L6znx3E1Fgei3z9F3Zc
pNJa+jBWDqnG0x5ViYGdph9HkVBdBkeVd1B/Hq3Cz+1GVP98tL1ANF4mzLQTtKso
yjhvxenSSSqPhLYSQ+qKTpucbL17fJDl1LMQg4xlJUsHWA854zD2Dm9d3TOWE8ex
g/pIkgvdEnlQQVlb7SvVFSR/6DPF2YwHC4KbCgA0PIrmmgQqcL0mW0WPFBhvt/5u
z7fdKkhdhqLz6FzurCnT80QK8hYE38t4oA4J2IDv8L/89m+Ffcqswzq5V1CLnRXA
TYTlGiea4P0QTyxL7H+O+zlJueEm9QkAoKTe5M79xFQJO9Eajzj7nmjYp/kAevDR
F/Tl1BK8jlrm/FoComX6GNbwj1XCevEjT9per3fRKy0=
`protect END_PROTECTED
