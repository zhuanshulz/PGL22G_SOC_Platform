`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WD/0xDj1AG4ayx77zy3QHDUcp5KChQH30emEhAvFvWns+G6tND6N2gLC0QigYGaH
Xw8ZYVewOAE+QrzXdoq10sIug5v7MxTvzpSlmPpTOcal5x0d8tphw13ie1ROYMOi
H7KEuoSkOiIukdc+Dar041kTh++9fw16bc1MsQkFpunSroqtQVwYa8uAdmad3Cvg
cXDjBueJB89BprD2j91Vu74X7lSBCCgY8I/oaLxR0z78MjSxBQ0CgemK/i/UAy4b
yNfhx/FoDxPNwC3Y1w6t2RRbQuhZvvZ+EZjzGHYW+ftIy4xmE/TUEIanNp8V0ebM
dF/cXxniplUkAn/yUO7I2STw5/HS0fFGRFEvh6P1xboGQnycofGPwosxC6CBi7xX
vwc4/7FYKtcfPC4a8bTR3DJZXQk0y61F3TFr6kHdG1pP/wSREPnL61Lc7p2m6upw
521qUfv4aoyfEY5a5bhO838c+lvo+JQ3daHlaDkS3ENyNS/Mk4pUvFDsCnAk14yc
JWAj1L8OXw/8bzhwgJG/qeIFxIe9W5ztN4hKEV0ysvC0G4yRwAjg9Pnl1pVUjFj5
5V/n0E6YM2FKRGHm8wbmqp1to+nyiJYgLP8KzHQ2SNAdlPTIP4rgDW3fvB15GvXA
EpTCEuPEqGdnsQrrJQNcSJ+Fta0nRh5SQHWirad0Gq+0zp4CbXdBGQMO2DB0kCXy
lnUy7T7ZAe5H3YZ9bJWmidvMKRYSwF1+Uu7xVfEEZLKrMGad98FixuROVzPhnFFF
MzEIGZTfWRRws8/Onr9l2aFbBJsWcoX0U8//vCKl2qZCFeGRCMs4kanGARYBu/bU
7hZq1k41e3NFfdl1MILeTv8iC6GvydLvLWd3rQbU53TWxJBgMoNCbwYDnpJtN+VQ
pdILXHrcgJDeiNPwDqMf/RWCDEnjtUmCukh4S9tJh56pBwTNmZ++kafWEs6ZWHJJ
4tbgcUHJYSWRwCAkLe1Sd3qf/KaN9WKzTpFxTL4oI5gUnt7ohphM7uUdrdZQOayL
q30lBjugoEMDB8EHQdrFEJyC/i5/TMhNuO081B2kxNy5IjUz0QJ44HeUoGyRKKBv
bJ0/MRZzXuOGqdBNA10YF7SWqJJ2Rv2BYyAtAmoopQEri4Fxq/IkqEf5Bz74V2au
GipTe65BR2ul4bUDEpW7xQyUpULJpeh+CReK/Flc7YDDXvXhf8nD8FALOCk7Mz1a
2kQ1+1f/6NpE/i4Bj53CJ9dQIQjsbJOXERIS2vpTGeg=
`protect END_PROTECTED
