`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9G0Ib70iiuheY8/8DCLfdUOt4BxHQCVX4ixQz2uIOfa40a34wClQMUL6HrM6Sj8F
hSY/sEVpMaWv99GBbqK+kjQxYDNjYEYG9IohqpfZ/v5agWsPMDuuXeAOwQy6vw3f
yRdmYe3wKvIi0XOc7vkRDJbYyT9CzWwOrB6v/zs8InIQY23+r8JnxORPCMkS4N8o
vxhsp69BG4h2XuZajxgDdulRsuHCB3POqnG1oznLFU3va/2KfKIQrLUpoVi2WdBb
HC9L2hwFPIq0cl3h2dJSermyF7NWjtWSbFE4/S4axbYcXvpktdrEWbOgArWff+7c
/8slqYg/VOChwSvxwgifFfiQf3+H5WktNt7bi1jbzkkKClxODPbCjhTKiBIt0P+6
BUlWG2i/5izAQBFsoTnegSxnmlM69XrILGLUMAG61AmUs0aC3buYz5jCGzpEmT4q
EeEc/faR4GF3neLDfO3Z74FFoPWQk7zpRMPUgRUGLBImIglXnBpRIL65UT2E4YqE
m91JFjJUeqXq/MTfQ//F7u0QinMxonkKhYG2hEy4F9vxmkQmx1HgYBDhIk5cm8sx
0x5QUlufRc36fsnuSPBYSvsZWZ3NG139SAZ4u0emOAbP7yCwfr1Gk5tiwh62Cn2w
swYsuDg9DhEiz1T0el2Hpe/sOvT7uQ3Xc6vIGzcZ/Uf9Jx1PP0FR524XHYxw5jMv
XHzUeeuYQAL3/P58PpE1TqIOWjatb/flP6jj260teGVh4k7e/6d6PlJ7Yzkj7XD/
5iUSRoDhFzs/+74GtAibejXOt1/Bs4mp5R+WsQ+hdow6HOxHOxRrxeTFzds5LX2n
6kp0lXPRF68kCwAfuYcXU35ssCVlY7OANnS6c2yupwNHVcMRPrEUYm8yBJQQY7VT
ctOg9MiT5Doa7xexcNGoXAgkLd96/L5D77fW4SfMar8wbCGn6FWS7Pax9t8SjIxP
tfSpErd8oKg5565mDqD2OOBXytV4OyLRsiafd6ksT2+5Rsui++4U/RYID8o6+T0x
dK2GsGrmi01VPh5Dvkf5MIirhuieCeQTmQmqgTogTuLKAdlBO/3CuqvaVqwcQCKP
omxsPCeAjMcfC69k6EnB+47CMfnkf7TyyqErlia0M7ETM845ObWQ3iCijw4zrwKi
pUMhFom/6QAgZwygwnHu3pCcYWl9IRiJc8Ojyrp8f+56LY9HnRvtZlvXDdmwz4n/
o1zPzKv2WO6A4YuAsxmrfGVCmCAVJANbjyIKlkvZDdKoLcDOt76iYsHEHh1IIJMP
ozA2pI6jHXKYm6r/4F8wgz5uWmcm6DZt/psVHyjTK3877m2q2LeBKT168roqg5wd
ZB0b5ZYlhHEqa49MUA8EQZOTmYYBOu33HKpfV+D5USNYH0pLK/+FzpotNgcFIjIY
3EXqoUMocxpfIuJai5fkjEfxtygetmeAFpxnkX4dLv75Tbo3UdvAlTgVjiw1GHUH
Fj8VvAYDn/xUxdHzUyoiAFxX7oXMFhFiPUfhS+EiPtY=
`protect END_PROTECTED
