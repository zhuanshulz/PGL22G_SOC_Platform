`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glsREDf2l9VIPPw8ed601PTtYnIQoLDakL4ku3tRMh1hDiDDwM0USGsHjMI8X6FV
i+32f4WanoRwm18cDsXIQQEMFbzR5VRP50sELNfvMtmZGykZl0Uhbe/B8HVQtvWf
50hRHy3gdx++fybjxwxzULqbrGnbTrZWg62GYajitPyZ/TCzsKqkzCNd7M/kZyK3
skFyokIIu8I9CfsT4hI+1KAl3I6sncpraCfP8ytrU4nH+HUE8Oehii3HqQr8HQJy
C9dxa9guHv64nQxk5RwhIaBqikqtK/AxXlHr8/HjmeWEV6FVwxzg1bUE3NiuaBVT
MVnd986IiRn/dIhSj1tEZQ7kWW128/kTUspTq4+O5GG9TgIaezIuqUTvGrsdtodt
zhHlhUNpEWouPX5MyirigcCUB/LDZz4XRPjxrk8yyPL94o+rRB8yUpZqu/sMoAjK
svA+mnDY85DFb44vUkeSvGar0J92YNjJoE6uuMh68gMQy1cYa7TxoakfIzsONJKy
Ch1q234/Svq+TBlouk8ulh9BNbNFLFfJz/3ZBHqdydIZXwy/bPCxmaaVlMZbpMoK
nCLwBgLx4GWFkv5YMd56L5y0tMWo5xwTS92WL7/HHXztOyBW1USVMRAvg4TMeXju
fm8nrNdQ/DN/eowVDu73KSTlzcDoOQv/Da10uSShNBQQz50rvTc8SX8sV4HMMkeu
sZemnRBOVWGYn6gNoyCg1wA3+lVILgq4/AXf8dXaUGRrQf49cH89VOjSuGf2XxkO
3rTWnCSTqaH7PkgMRnXhmFnwg2ix/1ICUpxF+xFx5hrH8YRHsBy5p87KNSodr11J
nZgUCPJQXXZbtCE0BgJMSKjV3HtJS1Zke0p037OVluUBSpjzLl+vuTsJ2jk5+dcN
syjhPQDeQVax+7THQB1h/5+T7hZhEvmfemk2IgKuTgxbJxG46as20D2m44hJFR1R
pmQ+yXltuFlqOF1454zqv/EU91IWiH2lw2I3ZD/AR9XFpIf2QaNn/DMHK+VVjp9J
P1ougjUQSDBQxs2DqKSAmTDpJ/OaYHXLVItFc7n8JkO81O2r4byDinsbKrnQKYMo
ouxYZuTy7R3mCb2qQLGDUe8DnPN3QMzGo8Z4IIO8hzuOPE/HacumLXbU2hXzivhh
x0UZ3icKjOM1doIMCnBdNwF6KjvJm0TW+YYWQGi1DEedl2PKv8mmuFV+0wjXiMYy
zIg2wB+aQQOR2+8auE8iByGQpQywdZZIntVMV6GWGQuOlLDLFwW0YId0uvUrsBJe
BpYD+9MmtP5WISVYJ3q0OmKWja/pkkQWiKBP0GRwhweNRBSn8oigd3OMfYeaFSSg
vVMW75cF3RyxoGoggHfW/5ZTmlnUI+ziR1YA7JdHLO5PDm3EWsVaxPgDoop2yi/x
X672ylOSZuIBmJiylYofi6tss0W9Yrggtcw158Dfv9hG3mrDXsS0b8DiaqFfLsBa
gFGVJ5eJEnJQAaNe5gSa4I69i1s09i6KM79pMympZU6F+04o3YrND5UEAutPnNAh
H9EM+fmsJuVAU1PNjkfoi+o6myfL/2v59UMqhU+uUSvxxWeAOb8QjG8VxETvKR0W
H1atEw+omFhT/b/jqcXSMB4eo4N9G1Z57sS/5N0kb1s+K655L4DanNYNPHBQZGEs
NHxPIlbRqMbkQY3AWi94571TMiE5QnLAPjrS42J55j6XzODIYHYXy8dVfRrINBjz
ET1lGEuEpgXe1pdMGL4Q7mZEALfcY75XvyT8lsNMzZsCHmAHFLzKgeRLPNWF18cG
OE0EieIkNfSvGGT5IXtL0rZpCF+bJ9Z1/SFYmsW3FdXdRDcxq2IZx/oJDgEkva8t
graNdrDF2qzF4mhSb5TK+fy7ZoyRwBRz5IwteyzNHhhiktsYhZuoaQ9jwQWywSjI
0Z1Kt8qrj/28rSPMMVYVtM06ICexDh54eqXj0NNNe0aeBYvbhW9OxzR/wT6/khbK
dXauCuRbsqg7WnNq5UtgVfl13fN778Q5dGCLw/HgePbhmjfV7UsW3BUNE18Qd3AM
lUDwIXXqGySG6+xz0EXyPP34OHnUthBHd6VBFIuiaNUCTwHArnvLNP9f1Sbtp47u
cGfmZY7pvCsZRqi+regeb8hT8MSjLYQUKMnYHJ2oa/zzw506tgPOVp5bNyu83LlW
0B63vd/StTYkhvsQQknGU6T1BTfszD9vuBEQoEQV++cNEWfF7ShjBmnToN/S/Kxe
37OZzmAiAlpax26xSJJNTxaVgPiAmuIkfg7VvVL+2GZTjI8ir8+NJ7OHaKSLfqJA
vIeyJkKXunG54v1ElfWml9OzkyQDClriFN4qotYM/5RiBwW9Stl777nChUNiucZL
csbqZLQ61+5Ba33Zm0iJ228WTyeOxSZKREUjKHwNtEi7K98TJFUEOG4vj4HcpIHo
2LASXbp+ejbyy+UFkgVObG8NBWqmJQ2qa7Qleywu3VSnd2Rb8vPCYEFXQc8k6v9U
a4oMUh1RlD9h+HzDMPaAadTPR9XG/CEzl6yypYkGAKOmVEGhocoZlVAy2/ek4bUs
5trlqcdua5OWqziYaLFE+1ZLoaMx3ppMVD3u5FiM0gl1aZ1nFx/EdHsxjUhhjUyj
teoN0rEI00EskEmDyqtnjI5GbLpep3BftUBFeTX4z4yNKt4tT9HeFq4L1ikGofIu
`protect END_PROTECTED
