`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRfI35/QF+99FLQzo27OK9U42eYooXCG47TgtHMLGBOjX3pm+7F/LdsBKeKBz4Z1
8GYVvh1PO0HTjC4gb8c91KNBKXcm6HkzPfYBr2N4lhd1RrUs8jINeINUuYJuxBJ2
l2NF+AtK5+Qqr2aPhvoQBBk3nvCVaDyCtP8uzjU7g+rzwi5y+PD7XPzflPzwbhA4
7/y1rq6Y8pCr3P4UmtVsBSssFeQBHqKxJcN6dyMRvgcQFwOR0j5hDCFG9V/bohx9
kMyewsGnnggdId0WuapMbAYFOr8OEOGNzY2F7YVh53eCRGfgQUnGJcqcfgqkF0MA
6kPFumzroUjTVwhrq52YlPRKZupXlJzYqolxbLg55UyJrurBPq9TKT8wJhOgr596
5jp6yJ/4YXEt45ThOhh213ifsDPhV8qMzkuyfomXDKqhlqXWsE3nSGHh1vGkOzOA
QjvRMaMf7iopdhma+g8a5lLTSRyD5DfLRIv6FcotARgIy/91OYvnpkPQ3BA3jKdi
/wY2b9Zh2ILSnDY9fNAENUS4BuYIcoV53Ruysb8k9kkUC5ZNhIu/eYvhHB3Ovank
prXP+x4F9Lpw/tVbWJ/XaQLQm8/PRK/qA7JRc/CxRcI7pa3PshZ6N87TVKV1mF+z
633MnXX6Cn9n9NPIcknq52ppGB30uEmH3iIND/CIwaxzIfNNhUM7Z8jOCSbPBtdc
lubgWLfhaCmAkr9GxKK0mf0ia47mEM2lSlnIasvOP8dMDwU856D1Y+ZkzbVpVAlP
/EKuOlz38uWNQCuoBMbkJW7nqpXIwKYlgrbs4iPqR0v6EWFHEmVjXujLPAhlhrE+
la8ET65MRx2TkSnmcPWeOAQs63epMXcczv98nMQrdKLwFFAcVIdUgLaQ6rOJh635
`protect END_PROTECTED
