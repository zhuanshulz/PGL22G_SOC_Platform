`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
634LOe0N6ZsQlfAWkN3xclmTZ6Ohri+4IsfIfWZ/lrh883DSvzbwt/+a7WJQQbfE
F/fkvBQpk/g+QydUnSBJFKDHkG1xv4nNIDKnxSDBI9QjHkBisVLOtQoifE0EnwbF
6BC48/CgO8EfLh3XHMmsQSjCEoomnFCFmgBmxKlX7Ws710foe009xlFknulAjaYz
pgGcVFNYS7T7zozhPwnnVBBJaVvyrUN3Q97lD79VWXnewwCNy3YlWlfFsG2gNzK6
YREfexREnLxuxC337hN7rxOGMzO+44/RXFw10YKG0vvcg6ue1mM+fy56LGk8o5s+
ZuqI1zTeH6PyIjzT31GiEXIiCKcMMK5xS4Q6rVFQi1lkIkxOb0WEiYCgRfyj2X7j
sKLpEbXefGx2sjueC6ce/V9yd4DoJ9lLHHIvambu28r0TjEw0XA2nUu5FiXF0xHc
/gIapUch0mjUI8QI9PhoPvJiKFgtqOKLhl84bz6BO38BGaADDh4OYQ9lql5b0gNq
3PgCMNtSMbMVtk7B6SP6BrWcWg/N4PyOVM1mxwa+2yn3ae2yuupklx9YJll+HXxO
kZ63gdvUf/8lefMbxtkvjv/5mMG1iEscPhQiT8Rameww0QCNY6JbQGsbw9W0XKtr
oYMNe3tfIJnYgjz1iAxept1bVD5b0jc/0bOs75HZHmFQi/6RfxRQPzMGCPb4/x80
Tuh/Gsc+bSPAJ5YxHrUAnijblWPPuodX4Q0GFxiJyPXlW0D1kH0qZo10HtzM2iic
xN44Kn0LHBEAh+AfjtgUTN6cx91GVGv2sXkP626fLsa96ILy78dNSCCSHCFCmwn1
tyxuQwGUh5XpRIgi2Jn1aY7EfwjS8Em/bUNx9KeGyr9BvFEoW1rgXlnAXhQuVt4e
vryhyLGq3Dwvekth2RVHWmko0n5tMnH+pBTNpws+62itxv7KONhJQoNIwegksV64
VxUWcqnh7h0ndSqxXJIVYBfCr+Rn1d3hFk0nHEdObNsoooX9gwCeKFG9if4q+uP7
xXHYMg4Vg7uBSlwutWmLLzrqtRDAX6TIgNV5IyLaSWelIWrRbnf25qzfZlYklZp/
ZqsyGoyxOwMKgDSvBmODpr/jsFwwbA/K+U2/lW6qBjMqWDn78LFIdfWZrEsGesEI
FxB5sa3rVbboDXz4i3I10Os9VpPao8LtYdfUCAKzha0=
`protect END_PROTECTED
