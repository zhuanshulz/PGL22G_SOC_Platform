`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ldlh87T5nL/eypMTV6Mcen2EJls0QvwslBp178pzQk7QdL0nu6kwYGzdtyuEaAf
BygJCgD2+LY1+QnfVYGmUVDsm7jbdGiJNQwhSEhsdk/1+RqajqhJVFCBsRljZY2l
MNJ6IcypcUQlBiAdQtenPG+W1HIdzGfpNIVsaiAfUaKZMIZijVqvcQSpY3z1jb6X
WYAOE/RlkHxryMy/gWKiEBlSyx4raSftUgK+UAzZu+7EBjhPhgM3M/4YdecBrdwq
hEaUJqIQsYC9dCXyMS9EWj4/HzmnMtYnrzMB7CmYaGAwuG9GxcbHi9zJkHdACQL+
F05Aqd9Ui4RaUTVuQE/Z66SAUNLOUz0WQPxyX+yCoN0JcmgJTPiTVSDqQcho4kR9
A/Khsq8UWsCcTUH4/rUPZ70g8LH+islMhaNrhIHt3dEL/NZ7QkEa4Xz3fbAntIrB
0c8MZ+EAAAIyrFEJMzo1RAsA/eKfmlregf9G92tRcE1Bbn7PXMs0/IgiYy08YQPb
2TXzhyqwXFBdq9AeIJ6i8lrK20m/E5ApQX7LPrjsdQ5YF18LonsHnkdzPKwn0PqH
z0jhY47jzQ3LwcVsCxh0tk6JH7oYuGlrRcPQ2zpQModa+SVtSa832hiPUC7vlvZq
EqOEN5ImMJCdvJhGL2AFLAfqs5Nlygd2BuHjyLrD9O5Smi+ZNMtn34Zqh+ElsrxT
EHWEI7aC4OJMjO6FHVnkpT1ihXQJcO35+6C26rNwBnCwB8BVYH/7wNI00yRQf4hB
`protect END_PROTECTED
