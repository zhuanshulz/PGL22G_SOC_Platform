`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ySoj/xk4LutonMPyNGlRVPgRbBC3iBbzh2b7xp43v7UEqXTvnZxG8+fzoHZoofQ0
c5xERk1lgqo8KueQ7nQawM26m4kuCdfenI0/JDZyzTN6Gc6xVK/PELksaJKGIRoM
q8QFXKwHKL6rpMUtogP4j7M6qKI4dsqjSB1LpvcUE+Jt8EEUR0nnhsWimtDYtaYJ
iVFnXPwlDX+NbzBxJHxU6PheVuvlvrHSS083wzE/rSvRe40IQEn7aByM95QPhFA2
27YFOP5qFwfMCjqW4tWwFu8Knzfhif1wSM2dFrhFyRm0uHG19BYVcMG81Llkl568
mQ9jOCJ6PfRodB4Len5jS084GfWoENa9WnaI0VjXmsnU/jz9FZOM+hhw7FKRTgta
88J3+bc8HCLND5hK+eceW5eT6euQW1KyZguPaJVCJbVynogxLakaQS8tryJYmBM+
04ELFS9wImJO/bDRVNhZDJjZY8E/Wm5xT3HA1AAmg8WFugdyj50LyjZlFDA6W6s8
NnFoqwveLc7JZqsrZwRfW3X+dwRgoCX7kS/GxzufR6Bn6kUPN7S+TPKfxCx3mV+Z
z4c39pKtUEt4mVRemptKvUidiSEZWIVSibokNZL1EXx/WrxbdulUaRhB7iumRbQ2
kawnr5Wr1tuCimjYtp4QeNHWOYDdByVwbcIcThexVGOmeDMhqnL0uhsGL1hiJLkI
G3qFHNRllux9cWJYnEc9R1WcOBzk/8rbwYztL1vjwltmrYLl5gkcRPDZnCaGXs+1
HbaNuBaMUubwFY5AB7/uiVpMSu0Wwlzy33y5ifrL43BJRKvq1J/RqN0S3+SsyWkp
FRZ6LbMvGnsb0upp915DLh1GjhvNRYXygM9FsH0uFbXxigzHZVJ238uP0MF7Q6yY
UcrHuY8tgxrcQZW9u15O2XlCrGYk6PGjaZPTNYydbtYVo3wzLcX1BOoVtYszCk59
syOzxXPSiOjted0++foeEA/flUtG6SbPbR03NidxWM3nU3Je+Ilz7uNcaR1T04IL
33CUXqsYRjQAvC4FH5NMkqhmFszlsc/gy3xhpCueeoSPrzF5V1LtgckiiJnAf0jr
AZebUBU/lOb7PwXuVkT04jrH97fV8AQIIbGHNB16WR7hP+nnGKDRBVuti7ItdhUA
YWi22b9kY0a/Wt7liZXC+UE7XKDwH4YcOVJernQC14GXqCVaOpVt3Y0ALhhPRcTI
M81HTrzZ0gVTrYCSW5TYlGW72U6DH/SaBeD4OBLodW2JRR7lTepXD5m7J4zRyKeA
tRPXajoJ4R9TbVJnzYg1A4/CFQxBR8k6ZEScvpg4GHRy0MvG10jDe4oiGGmKhs5W
ziFgymg2lOV6BezU3yh8C7L0uWIMLOTbanNQWIEQvNhvy3dKIlWnhovu1vYhZSaM
Y3heghNzeSbgiD/aziz/2RqklJhgdhZn/mxyFWECOe9Vvze7A/tqbwtTDpjOyCFq
uxSzdrf3YDtUlvMhkxVa6DcNjzeEDY5MDfI1TGeZepaV960XwmdtQ8eGXf2hsAxa
QHDJwesdfWjA3bHd59c+QZ7SFOVJSTZAusFqouxaT0QiO3wU/pq+vkgjLG47qocu
zbJbStLJSULmgpgD3W6FvMxvU6DE5R2FRbrVfz0qKIujFzRrTxWMxVKahpkayrqu
CrJUwOs1TMrw3xT0J5TS6d1yYGb+v7oFZNT0vOuTw9cMeG/ZpKFonfar3ltRdWC6
rLhfMZW7w0S5KTNhaBGYmZdfxQm0mpZY6leYqu+Ui0VESivrVDrytDgfxs/t2Ja7
yAFoTN4uLRsp1+ChHoFf/Y74b5YAY1RLh+QB2SLd4Ag6gxz/4xpYtcyDMwiRhZ++
F5sfHHrZKNDNq8VDkkl/fm0mBmu11458ugTxNKQg0nveSlkQ2/YGBsyVfdVQ4SBZ
2lo7rURmgsONp98wT73KZemnMUc6G02gq69mBCVrqvUvTpDxAW2JDdyfxLBa4Bxs
sdHKEmpZCp+H/Y8qQJ48cCTxGq6yhgKVZHb+nAwwbjjyu6NtkHqEeik4ug9sOw05
INaGixTDCD1cISXcO4h3A7o9bKn1rZyQTALS2iAASWhz+HJhgoSMIx5VGLWolvT1
rTxv96yD6RniUxv963+paBqs+TvvH4piV1YulxoqNo72doDJU1mN4xVKYdM8C5Ld
gya1R4kQrZQg6KyZGEjwN6t1fNVx0I50gRYAfuBgjaix6blT8dcjBb/Bt8lwdhO3
FyaD0ixO/jgVMgZx0pKjPPeaZo0fH0Hao2kwc9pJYb+Uc0Iaft3WhkNYXCG7AH1W
QPyQBkSyyGQTW0icBNwMt+HF7Ds/XdCfPtEo6byL6QTTRi9Avi2+kNzB/XBDI4W3
s7Sx25UJdbP/E4TitI8/PXHR26LmO3XpLg1JPyk7KKvBVhpthlOsUYqIQ3oiSCyI
i3we1Tvrg48KYZZ0+KYZ6XV6ylyPWElhGk+Xx4yb/XdYTdCTQ8xQMzbwqrHvRVIk
nbLhamyJxSSxfpiokScgww5MxeF4frPfxyRm7+fCMIb4Z7GoaMuWmCmYENSboJMG
SJJSnAK+3apr+TF55WL8MUvM5moLqpJoh8TXnxYgjhlgSIrtV2rCDAalSQy7jt39
RwqLSco/ihCuYfjkyu+A/SJVD6t16vw8PBhcieHrdx0zTuOQygNPLDcrMYUu3AFo
tA/UHpfVDHs8MLaV/Z3GB36tAAtUS+bYHENQI2sW5+XR1LymP/XiUO4p/l0alAfA
4UXqtyIH+oIYVMhxXjLM9OVNZ39XiGudu2T2F/bbjcuQE8fKUr60Cnxf1TFY7qA8
8Z5FfxlR5jKfg/+lFl+IeusPGQCDDi/9t+R2Jx9EBxZLM1IT/LZLVUeqIpmtEaaO
VSGTew1zDQW1HmmmzcKmnKWNY7XUq3C3cew7l+5fQPU6UPlkvOTNK2tLSOsyjiAx
3G7EXPt9oOJXZwWmzuMgI8upW5rdCx9n13COF1Oj6VnJ5TcRpWOTHXuRpPNgLPeG
jw/lbbMUSI4z+zftUQP/xRo44QB/xwXxTdlI1fvWN4i7+dLTI1TdW4oTp3HpTQ0C
sfpdLNDYo/vVuQskKWdbQqAR/6fVqjSrlkM/0CC64qD4b5aWjPsv7cXCyJbMPmbM
zrCC86epBjkKYmK3ekyMxAIqvGiyt50P+/E2p0knSwqX3UXtAu+/6KE6wCUq39r3
/QNGNpPX9+1E8CecsgCTvSUt9Z1CBKdQOaEi0U3A6FVrWEh00zwsrg9q5D+/xJvR
nQKflAOeRPAp8dsSe60nbEd+n9zhUIrfjHl1+uqEMX172jgVSCOvnduPzFfrlwCf
Hz6u3w/oA3PC1z5WK5LOzKgOFy9CBpwouSAm0vEe5MsT3sYevos/j3w0aAPfxmuq
7GQ4O3YeKM91ygmrrld1LhnICWGXgetNZWr7wm5K0w/I73M9HqU2zy6YeXIz3dDX
ZUcniQ1WckTHzC5/joiNYR9xfPEVrNMALxBmUNyDLZZ5xBPS/Hk6tHkSpcKzNOvR
YE4jfKZ1Zztg1n9ceNVJSqFI+kIbtzMFw3OXen7DfhF9yt4hsA2INFd6F+cQs1k1
cuPz1ID7spPF8ghmoIzKzwRfZf3gnDKzFubkFX2dus/R2sR5LzjChyjKjZX/scXB
Esy4V5bxtjfqyIXvy03BOCPT6QNrxhwgKZkvoe4oix/74OzBXRU4VH4kcbTDc3Kk
nSrGWJY88JR6cPLOKYD9sCbptpRRwPof2TQcF4mt6xDSWTBRAffb7fcD3Vt+EwBg
gM7uLOyim35D6cuVUEi7S1e/F8Ydwtsupf94LfLyp1+g9TYaydBrU4mBE/bEh9Ko
h7EcEqgmytE83qr12pzqfcR+6Qkcx+yJIi3/FjPDnsvVdQIa7kghMtAdUFK/BDNS
c8jizylbBMd6Plx15yKhb0wAXW/Jz/igZ2Ywsh1AwsqoPLc0XQk9mFKHqeGG4iOn
c1B/MVoH1c5adn49qyvcIaSScYBkXwFe9xq9aO7MBqPEILh4SyGIl4ZyG3MpGDUb
jowhRCvzXnVsaWSmj5/pCnW8amIpoZEj4FWYjNgozPg=
`protect END_PROTECTED
