`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRkdyiTm5ui8MQF1VjvnuunCEj/U4u94Fr5hAmapiBgwOgJv8AvgIa/Rrosh8gwR
fX6FZSVfO+TXKcRLGy/qk3nYYwkMmqEEf3RJweKkTOns4XlACqWvYn7MkMAnVWpE
rMmlGrm+jt6rr8lp/6QGwaLcDoMDH5YpfI+l9Ruj/MiQ5T9gBdU5d1NRk+apU3e6
MxBlCVUzCeLVSwgie3JiKf4Om4HVH9p+rX+uy/YNoe7aCszvKkfTwOChfj/VeHby
rdXoMfuiUiA1IitRqavIKTcF+pO/p82VIQ0GZcuN8++/G+xKV6kTSNBJbpRDwwG3
KjtSXYl1eq7gttTdAO+Jzg==
`protect END_PROTECTED
