`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1FhJwJhdLZmGoMG2v8zk1sU3KjvnEaQNAxtmNJRtZqTpcU/A9MTc0NkRpgbhTrzC
vQ9LrD87vp9DUfqYnkSKjQwIlW8RYjp9iGOdfBIMGrX13vvxjIeMNxD7O9umq6jz
WjP+AzjFxIgyLnjUUKs4t2HFfA0/Fz+vCCKyorfYdsyEnJAw/bcWgJ5IaQL43ejq
zbCVj4M3jBZwSI0J4lpByCQFBiUte1zqwUJ6WLTA4ABlvPO+Came3DH+KrbuMqEr
e5T8yPP7PxoKm/ZFQRjKgMUYSvfYQs27R/gl5Y/UeqOpw16eqM5OuEDWvRJZ3s0j
Va2ZOfpnQVuMp336ckoVym/klY0wb6ptUAwFviWWobDfMECCLicv+xJsDoIywivO
AwXWfRqMOOEJ3+gDTqwzZg==
`protect END_PROTECTED
