`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1RQHYelTv2G8PIFpRAmAIooD5fb/000Sufymhe996RHipK1vX6BBBZlZ87+Ell4
Fl8i0c8djLHW3ztskFRz/eV6PvZZURGkZKL7mQpuFfnGr8bnOnbkUgeawRyd+aBV
VFhfyo0UmMzAM3fJmGlb68zVPPzVwYFUDpCkDLjy46ywW9BYKRZq37foe5c/wONS
OR+vSjKaXEYQyusEqxqZC55LBUrUKpdvox2BG+OLoT8lt41bwb9ilibT1mEGz9Z1
0hnY37XnY8bAzYRkbdGKsQri3s2JWfZfVAbwvUEkYbNkAPV8ZHF9RVzaz4hoWp0S
Ud0D/HTFvA0qZW1hqYOqA5UkSvmnsSnTIaL3nmyNLNRCQxpEkwFDFflovMt+MBU6
a5+ny2uTk62s9UQpUL+FUEfHclwO4LOhCYV06eXQHb0=
`protect END_PROTECTED
