`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OAaFpQkZqcYwWc/3rertP+EKhyoEdNvo6JUZgKdqVFtl3xR9qFyYzAGOyI2YrRx
pKocYmkj/lsvJzpU6PU/xE/beKKrMAAEaslBv0+0h9VQtrw1inyepYYZmX37ON3D
1WfVr6V+vxcztwSN0vdpAA2E3tOEQdJ3Sz+omqr+tDn30XrR9e7C3sbZcqThRw3q
KNbtIqeJK04wHhxJv9+R+JA/Ddbp9A1bhuZxBsoarphd7GIVrTkK3OLf91YR26cT
om7We4Vt3zcyktde0EItw9lMv1OI36IES4yYZYaS8D5NMWDceXrmqT0/w+RVaZzG
d2IX6392LnoBO/J/gH5JsbEZ5Ukd79mynSrO0Pb60Dcz0lF7NS9K1d66aTu+yVIB
z/HHwqXVXXHuD5H8fHdabRETGhzIjfEzEeMUujQdBW3YDYjWIFRFm6H+8Em6kp4m
env9U9JRkoGXUMpVqDwXMr2mHzCmfFnuqv45LfLLMVEjdMjGhqyF08q6zUQhaj5k
cPN/rRXx9oXIx8fi2Pak8DWqzK3WjqTZwAYFmsWU/5FLd9Wr2nyB8hQ+3ufgiR4H
2hposShRB8m8edXrJA9Jp3/BA/gCzf/J9gCxUIPZGhkPKlPFxTkWM/S79AmoMBaE
mPlc4Pk02XaBzAY8/r5QF1XNRJ+XDI5eguHfa1xqxjTOM2D78lJgGcL5mswxnjsh
eW55SfIE0qnW3yRccODdeu19FtzLuvzA8cs/jNi5ZhCgMOeovxM8fP3Pi+7KhJur
oidZmlCFDJ/l8e8/cCRc1fU1YvK8px9oXiDzEK7k3gLmgtIGYP8oa0Tq9hFgbrVQ
emOmdpR8r3uAazncI7b4fIcPJuVmRHZjKP0V/vHvgbzYMLlm81nW7QwW27xZrQ2M
XZsrpXl7rlMWgAd88eeW5VKrpEqOTjUnyBQ+5UloCg/5Sl7OJkfEXjRYcPTZyOkY
r4Yb5tjJ3BYhDphmC5IvOIcvj9QHcc1c42ltomJCkmc0vkd+5NtU3kv1H/JiOMoa
fx9jJeivgm7mQSamqBnBgv3RuPNlCFUzgGMtiT/Btb8P8gj/weLqBAH/FfnrU0qs
MutoiSRfiFJzWBbjjjM7EdFazJ1oXCUoKN2b1DKjKTw5WEdXEuTx65GVGyWypif5
Eojt8ymUjRkszOFaXaM8lmCknJh02bJ+21f1yEj+GMh3+UIV/bL/8IIu71L0jg9g
fuIvhp0F1i/+jiRLYTu1jV4nLBCWfDOrM5HM+AGBVmY/w5mKJfYNwQvFPMP8v7LG
BPDaW8aq50cxH2Gh9I3zJ1f9jk7nGHWycy3hz2CaLo1IJMciD5GPRd/iuZTTPcQU
WdBWyZl3Ph6TBwXoO8MM4S5eWJjytxgPS71Xy3K8t09JJWk7z0WCPOEXcRL3ftf5
N8DSaUaYl0Vkr016rT2V6SMRD1zm75g8h9mlxb7gwws1eTeOx9TphX3wNUTDv/PK
sLus4/wYLP3nNXCVNdjsGCMoWQYIjfb4DEfaQerdqzHOBHaeow3HkbWAIXfHkSEM
uY8ouOlaQptAHh8UVSmjV+8rQsZu7CAeNAO5iSVhoYB30gZcsAQ87rGGJSBLHXEn
CAnrgCImGI9H96IsgX5MHUsTxM5fyUOU54KaoLpC8kBUxMw2MOgFEkqe6ydoCWuz
NNmk208kJ8cUNdChmP3Wf++INKiOUw1z7I8nvOsb+rH/9tNPP72irtyc/vppcX7D
phoD2/hr2wwuiQ8tjYUZBjsSc+3SpXYv/Ytbr9cB/LZxi/EF6GztVuN8ml6EnyL4
LWUviRsSiT0lTidAaPNSP1tnYqef4ShuJrCZNNQQpKy4O4CXJq88ukEii0X7ZFfd
urtKsEUL5vW08pximMcQLCD4cN4kh4ay/CnMYmVLZF4wLuXGaVF4c6IOQfwWdzpV
gtDVzCLFB0pDUpGoLVDzCouIE3jm9b+BRqgxoyp3FQVeUoCfr/YC/ALbdSnpyzp4
2S5Dqk8JBDn1MaA7dpmfPPiw4+22w5bkO3GdzcyfZm15QIVdvGV0zsZFmYjoFaHD
Ri2HqHlHAF+/+bMG2b/wKFjlo0Rgi8Qo8/UkSZ4WmJ8=
`protect END_PROTECTED
