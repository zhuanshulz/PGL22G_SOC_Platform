`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hMozEfIlvhlVyCurSW7DtOF/RkDj52sHba4C67Aow6ZpbaBQf3WqYxIIWJKXl5qP
DH/jnnEboWmP3ejkO02DjJTBXn7kz0rPECHF6LY0A+fm76XSVm/ntN3dBOlwu5Jt
MdVaX0ErLmhtSfz5czNjjnw6FAqDLo/npLBPx7kXIAkvuJ3US0FNPK+qkC23Igkg
LYjoEmyp7aa2KJtgD3dgA72XDrwdJigqaPgHzxlj3C54g4GF1upmElY+tdC4MlGy
YrcHKyjEK4BBZeDSD77ujHkdwcHbyFScwBolZGHiastE5vs4/sBKm5ryvE+Jvuln
xixsCBphC2G1qkR34opcJk0D7buP475NR6SWggNhUb0nn9m6Nhgc4r63jhr7nCX3
lUJGBuBnXNdeCHhX8R+Rz/f1fp1pCsmPXqJEQKTu5vQWS/c71+faV4IAcCbh4B8c
9t/+Vz3CyPT49b7s0PYLcVtzQ7ygdfnRT63L6viPEnyOo985HTcRqlXbYbelMbSQ
Y9vxo/c1pE6f2IsF1jHl20KWSn5Yn12uudDq0VHCbEAWRWin+LlF62G5MifnQjE3
2pTKEQqUQN6e6BDJ6hzKU0Fu69zlhXT0EffwVcJUv90sj2K/FkPXrugSCoOBGsDi
5rN+ko/iQn2+grxF9gKg/YCQ0J/FWfOG0rNn6Bk1s0E6kZQMOQYjhumizpxrrlzw
dytRLZu9Md5DPvfanW8w2P+k/71/cH9TVWgtQ2PR1pvWRrfECjTZTwSKfykMXfAA
gDzcLqyFf2rbS+pBzWzRcuZgA8jAlujGKP1OtjBmMC8JtW+NjfWHJXKObKhwsHAs
wGvD5lwMhPcfvchXWFobrsJKCiZi3z8vY4IIUQY1V9zgnGul8T2F+ss25IUhctpa
wDJ2rdbldSnBru8yQCPqVPFUrwWFdB65gtEySf2qNmTQkmhSDVDKA8PRpNqvuzo4
2cybKSuaU07mROD1Pw1Epl1KCcu86X8pwdUh5tssLvvX2glN/kaNRAFUF+9PrmTN
CYW53Qh5Mli4wQw2nzWVqt4T1FTSTukxOcPoTUSYJOgUxC02B/sZRnSPnyrFNYmC
BEj+oHPGPEflHuirVQax7w==
`protect END_PROTECTED
