`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJd2eIeG5AqLJUGySujct0Jj5IOdiDX3AjR5/MlyfbN9kmfe6VYYgRpCnqKvEHQB
mkbN4+2MvjsAGAEokjhRbt/R/VFcgqaXHZ1VLuCbZYtWvEBkI7NJL+KSHZmcE8aO
H8mgTN/HHqkPtpzGXJdMEPo2sD40wwUnO1Wi/oQW/iv9TxcMwYz9mV4rX1wpKkH+
14LjApSoauVRSEfgLclqoM0GascrgaDKo4iRmxlOOaAzfA+9ZRCEEbAmNyMXJwwX
dPHSyb7s838ZOTA7BIBAKR3g2+BxBbd3oB/oGtgP/TPD8ShNijD5q0C2jhTS4Y+v
NR7X52acJsVRlUhRaet5RFao1zVKB4wZKGRGlTpTHU+cZCyvSgoVEuTeTnuWeLi8
m3MMZLII55XJX9YCl+FjYQJpvvi7ERLw46CDsDpStgx1/Rv7t0WTua6+yBp43wH5
ChjMV60M5LfbXq4VhBsIqbyXT9VbaULQJTAdLCgavqTC3/2BDXWwwlomXGIQhLXR
r3qfJbOSeW6HPH9DrNfeXBHrE1H2V0/0MRAGOZ3S6nLfrx4u7XTItjfsCH2sUe0e
7YQ/Bp3/vqnNroG/mTQknmiEU3W1a5CIlZYaSwZOwv6WiCq3e2NefRHruTezlOgc
GyfOEsABXPC9AMOo1ZrPNnNYgCEyFTYsxMhJ50LmNid95w/Eo+PNVH64Ve9tpeMQ
vA3eH8z6QX9OZ1DmB5d9X8eW1Nt7OSY8WrGgp69MvrgwBZFO+9S/ZkFPZnpvPt8x
N0UCPWvo3cVYxWVapgkZdy/6hre8HBiKCJQ3MquUTzpP7OJrRxcy+fPfESmnbx1i
hVf4xktvxdWq/VTUeQyn5hwDfC+1K8MiPTaSx/++a6EEpZQJmOGLK1gWX+uXRfTm
nK/njvpLLUgC3Om3Eh5YGkp2xQSPa9ZYBaaykN9CLEYIkAr9Nb01mVShuf/pqGE7
6NyjJ6F0TjC9Yi5iBUxPZOPpUrxEBXqmYh+rm1KGeShTovBELlKxA6n/fTd8aj49
aJgrZnijY3qWFPqud9EY4n6RSjvQcRwOkkic0gLmy/NtnAM3LsWoeYyT7AsNrK75
GQWVVW+7sSLGUrCwWFvdqoe7JoJNVYbhmPRKwJhmFWGsWHh9cgqvijJIrNq6AuVj
TqJi2xWWqx2oC/pd0Hf19ohwD30+eNb2j/MDTWPLhVr/xvuJJsQJT+KRWJ20uH5X
5/JYScsYZQ0bhfsOnKSxe4zhmUFKkSLmbihSZJGRh9w2YHQZkb2WY3H8gpIrHGsn
BmBdtpgWDJulh4maDXQJSmQHYqkz2v/qrv3t3Hyf7kBslHSkNkKRom+yRM0JRwxp
XeWIl6Cp/SA0wkrZAiTG6fzX2eidVZ2QEGmCLaXcwmRxqJ8/Cvmmm6m6BghvAGmF
KHoSGplfo4Q5LqWQTICpigu/0iLDvi7ahl+pXTdGJXKf9nRca0fRK414UBbWTwba
1Fb0Ea3bYJP9MQ1IOg8KObq1a+BDLM3VfI5K5Tbt0J4KC747tsm0y9FCmOWBkdEm
hfIUscr4MR2XXhUs7XaH+sk+gL2AMNZMQIoJBoba598pU/JV0K+5ckqeQ+hkS9l8
uwqir52uh255onZLu2Ngl+NDlg1qhJbFwVeYqy9lYLt9OlEGHhCqDBh4CtXndca8
B2Os/gkYrR3I5DzxCQdClxnAAtbrcxq5/JMrobYUn3uUThcfPsBIwYsxox3vfkDR
xYJvbGtR2PPdBHCWmesmUfdHRsuUFzboEf9LPVfb9rw/7vYsGfeVI+2g6usa+nai
hvAGImIlM8g60G6ap00ehSmj1c8UN0PGEW5TG4xNDzimUQwi63/UikZHCfP7w9t6
Y9VQWC2JsJfzrHBA8O7eHDJscDeGM5+th4+UebJs6nSvpgnHos7UELDHybAvvDIa
7krvEBi2jARudKyi8hIgHqYRRK0emQYdVS327RpgDZ1mVkgtbvfgEbj+CDwI3zHJ
OxTAlJlbb++uGUv+wDv0r8Wfe0+qmjISvu3WeYs3CLHO1sIQDsCFcTgVSqFY9nP9
3PPDyH2BlhZuVggxdLu1Tt4bbpqqaHkcEPSbnZtptzQ272VhI/Jp//BfH75wIjBh
qxl3piDR1iWrMeN7jWlUUMgZrZ1WBCBlvcizeu2R2tH24afX0omrJQDx1cyDoT7n
G81T33qJv47rUqvLX8AtcE4gUooJUhrlVIP11nG/agJ4qCCAdgWz0+vPKfnsNJir
wKICCamQy6rUsakY4Rrz19eYowJ1AvAJVYFS9VxJlL9o00TBSqtORUnM/WCpXMsQ
eVDoo9ShnZVZZyXoMIolYhhJj6NF2l68mTQcaNieHOFQtuoG4SzBPO3H0zLVVaw+
frLGvrBQzykaEc4fc+mUYxPV4zQygmCi989K/VW+V859slHLVKj6TtrCWAe1GTYd
69TJwP4m8IV4OLivy3S5k16TK/MMWD96Pxh1Y8SnkFDXA0MXhX15kW5C26y3uinl
ZnwkCjVNAQaLRDrX1ZE0KfhrJd50GfDsxWX4x02R2oA69hpbydD1b7LigVQzdV2G
ChsI6d9NoPid83oXRrjfePz0zYiiERvUPBsX1BWBa/ST7fDflapqegYeJmeQTXH3
bs+7vzqnnoYPYCE7kJHakkKbpRc2YmbIlHtMBugxoEEOhhCji2bzfoSBApgA83MH
UCCo6WSpchPq1uswsqdXn7iO949S/TXzsLI1L6pmPAUXdm6l1FN+5rifoKYOYVtg
SN0OsVdYXpBxoPIlALW0H48mqYRG8nF5QlolVJ3jkBliyIvlX6uKonP8FEV4cCJz
CiKZgg2Lh3BQpdKLYP2QTmNi5hthjNmJcfFtiQEOnM9fZ3Ssk/GKZ02BIywclqNr
Nh3YDcWixAp3EqxgOKbhQl/Lh0JB2hHCduvefqCYiucm1/ne4uzgn3gxVRd91cc8
kxG8/ZDra+mOz4XJjtUWNfV13mpT6QX7auuDh4Rc3Z4aXsAWYqdhWPUuyX8pVN9C
BGCcm4HPUMrs+sWd5JRGCd/51r8L960y+6pOgJxpPH2nJsafptkM+CEIpdP78m2D
nR98cRJ/YeBzcOE5lzOs+Zb7BDCzPmY5Um3czLhYdZSc69FjlylKkvPD85q+Ip8k
dDK8cF4mqObvAQ+sIPjF8uVIe6n2sgUx9Kt/4E19rJ3Lat0hKt3DMnQvAhPqwDAy
dM0gV4UTyR2159PsQZ9l+/0AoCqvTDk6mDgZEvNoGob5hSa0ewMiCU6np9GfEsT5
ZOdJNMr6l1QGH/vmwF6yQlaGeSmqcIfzpPzba70nmmCspjcStvwDhjgibxgw53a8
TPKTg39n+8c1k/ShTpWcnNHD2L2sybrR/VMUeGnHoAAmbQyWbT0lQ/4rq8wWsPbK
qd7sXUTn24Vju2P6Rv02kKO2Ceq46MYnz6otcA9/CWvQfC8/3O3rt5Tgfu2RDsxN
oOpUIhGZRKMep5co4N5uX9i3Nfy0f1pj5MQNlRibuDcwW2XUsVLzQAGcZZfnr8xD
CXVJrS4xK0Z5ZXnKlqMhrSFLHveO2eTtgkThJEd2tnpO/WXRDaECsAn5ijCLDh0d
Zk/y17DIXczV6rwYLclqEs0f7E31fWJJsPvCHN+zS3E6qJBVPF3Mct0HBHD0hPCU
gsYq1skxJ2LHb24v2TJIFQRd2PsmKG3j6h38DM7NACUsFrXEVX8vpWVHBJvBQNtw
1cWA9GaiKm43ITmcQOMMxUZLcsHnQU6UHz5dBj5mt4LUrgn6x/JvWbeQWgtieivc
HrG8vDyxQ7DqsBdGOS0Vvet2OY+bXL02666FSCuE2ACkj2BONKMzxDFNK5QT8YK7
uJxSexdl0Va+BeXGXVGgUY9qgImfDx3a9cYIy1iLlWpqiKumrLJ670juPI6shtYQ
LTaKSkLOWCXR2+BSh8nxshyFiCu9DnCN1esiEbAcKVNS3qnyZxQENpUbPdFeoFU5
XIJnhOaza7k8N/6YXHh1hI4R8tssSrQ7iU2nHALLkq2+gYMPSnhlqMmrUT4xGN2b
Wy0wfWFtYaS2sO8+Nu1AmO1ov0E/OqeAHLtvv3WfRX1yRWXa8enTiiamGuB0egu2
XboxmP5GRp+xaFWrCBuGmdgpw4V3qgyL2gUbeaOKYxnIk3rrjwV/isJJlBwSaG3l
ITs9Yu7lzE1+ZR+K5thzZijEN+p8tmCHkCeiyNDvuY1On1VdAMn6ve8jquLAuLyD
4d4cL3qx5w4+Ei27XVt+8kWmTjvY3NbY4/11w5l5yjCyG7ziKSZfIqr2xv3zCmIU
nswKDOPLyoygJx6Y8G394W1SVOAYXN7b6mR1Di+wpL3P6qR4q8I1vwWM9ri7Nw5U
`protect END_PROTECTED
