`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4sIrZu3L2J9gS65+QCuXtgvC/vCUM1rokAsdCWRpuIYU5BnHoFILdypt7YhqXYA
TUmyN+QLz1Fr3mvqYR3vAlipcFDKVUhUf3cTjwtHN2G6XDggLEbnRfS+AeWzCthh
URW/jUAbM55PnZ2CyRfdQLKsxB5QRqRcX/G+gVAjopX/I1z5WnYR7U/bZ1zP/WiZ
LKKITkv1lMuR5MNlDGgRbOlhajDu/y4T7N64ovrBS6kfmFZG8WH+a7w9I/EHDbnw
B/vtGpdetgt3+PVepjzDuG7UkheckcXFc+TzMgPFDWPYtXqVtaazwL/AoXfS37XA
W2CeueoLh+OiNmdUyL4ojmUknoHqmp68VARylIpstjp2l8Im1qPbX0CtOS/B7F4/
dvh2X3ukILQWETJ9xoB+d1ZGZ3t58N8iEHAW0IvagPEfZgHNninuFrxwUQTkxJrD
GuspsLmF6c34145EvL/+2wDjT5uwIypdv9FwLHneDPiHxkLKIn2pmq5PcOrDwo7X
hb4ISS1gK6rEx8N5dT6WKTRfs2PMEI5f0xmAGYBwupE/e2CcV9sTjo45OhTM2gXO
EracjCce+T7t7Eu5S5gp8D7Px/06wklJ7xxFgl41OGUWctdJqdd4alyZoDYAQXlx
IH31euLmyvxnfcZMfudoK2Gq/+y1IRy1zPuwwk1lPOi8uDamnOTmKO5qn8x/oux2
`protect END_PROTECTED
