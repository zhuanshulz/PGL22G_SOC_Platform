`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAHApak1H+ZkkqsbvEssAhPcdrJ2xSUH/SqeznfJaWnPUI1j6Rrb3daO3UuhIgVN
Vw69zGgB1DkfUYo5gTQYSJDyHhtCdRob4qWzjXLqRji4nUjeCDbHsYGzaCZMd+4+
wCLFQuwZG94ESRifHaiDvl/T8mc8pL/ThWRUsnbht+vFeRXklAPmywesAST9YJWe
+NhRXpFTIBidtsN0/VZSMOX23Nv7bRNIT4Ls9F4IJ3CUBSbgDgXeofi8GYCjgt43
x34yKFWYCgycDgXuRYq1XIbz4N3ADFQzKo8zCNhhhcBg5h9t2riD2NEyaNSqy3A6
EOMDZivXLOvJAbEUHfGcJn/P9em0+VPFpyqSiDuMxWEyD9/d47qPyRs/LuXcNmeu
n7VYLznfR8pNDULut9w2k0SW3e2Pq8yQmW6umdeEmoCYqb8af67bqQ3I8W6CA2XM
CSLndQ0oAtQNSwgl3vcAHvt2DI98G6MJZ8F+viVDTwEoLy7AiRv1GzRQ3VS43CVr
Kq2ZWMZp3fLB+JeB38ZOulXIFT4XOqOEeed0xvhmMkCXc1cpUZvakcZik1/FG1de
rtWG0h0eKLVJRgJmr+IF1OslZ0hPf4cWbDO6rLeqm/UFkxKfr+Qwl+vm4yjuEDCx
wpxBxGz/RiwGvuZtBQMOXK0Dy01Wa8eirA+LZyZsTQkkO3Y+5ez6e0/o0XfvWefl
ShPBBALCEKB3teKpIRpqoSbSdRvw05m3JI0pzWeutGYij0j1IyZWdIpTRmWss2m6
iFTkO2S6YLhs6VTbhWXCG7h5CZKKs27jNebQiaELJnnhArBuFDJH1BlrA2FaWVYs
EAq/O90U4kxTcFZF5zrrZyWbR5pnXox5UDdIJkt3OBoWiy7z/YBwvFDca3lFG3hB
YPqjy5No6u1pAb5jSMrfZpfxCY1Cxi3+eSs33qm/dJRXyAiEdSkXR4juA9edVFsn
xwLThCU4Tsy2Funku6egfDeiAnFS/7er5bmi/UkZXOa3PZOU8NnatT6TRhDjptvF
eArnsIBk5ho54FETPQfQHkmHQk/VR4cqzXJb16uQ95TpeOJsbwZlD3OVuJqfj9VK
nFSFhM7AztWSQL1spKwFqWqh8HeoZsPmVe5meD3RWIA=
`protect END_PROTECTED
