`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdOKukuiK7IzEcRPpsi3wOaBRONDxv46S2FDHNVbHpfpqtQTXxOWlN6EBCJQwz+Z
J6a4k+T576PEmRIUI9TJ3ES4g4WRjhqiIooDtAgi5QZvR43CiGibic4Ua1i6iMXI
aI4rZ40VUPQ8XRGN9427+dCDlnuQWmnrLVuvEzoF6346MQKZOiq39lyBdhdy1//h
HSEUfMNRIVnNscotrrX+q6LfllQTLoeyBnS3mKvPhuw+kgyW31xpNV9dCKVft7r5
f7fLFMBgckhj4Qvx7yLEoaI4pGjpeztDrUkhYEbKXqczs/8lRQTrHyVOi+BsNJBX
HCFAvVVdcvTiVN/MMHeFwZgbUI93yZ9ajrRG71O3R4ooTQI2kvPTuCgmOOyQt8p4
d4buANx5r5KQurbnbZzGBXxr92rRUItg7P8Hq3m0vQn2d+uOflWrii3EeAYANZZU
65VMMfG3Uu7ugSfpTD05I5JGpRXCUjEEs8c7+RXijmKIll+jYmi2N1yBHrEz8uGh
0xTxY0DzGi6y1RwAqWMt3w6uWjwH0TtnE4PHjmTJn1TfAh8joAObrJyZWDrhbB1p
kCVl7G8HtiVxuS4lOhxMWg==
`protect END_PROTECTED
