`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0iN+9MM5fof2KjDjgHKpJJwEYkQA3VFWUwDP42+iK/QZ6daiVNagPePQ9B7PIzpo
0A5ogGkfyxQscZLlIHlQaqfa1OTPi6fjI1bt4j51obB57Q/WvSyuRQA8ehQ27AKY
vx1GMfDdFQBbe3o6ijwPTAQOaaGBAghgBlP6gHh2RRy+vd2nwqQt2g/ndWVPn9+Y
Le9KnDCujORW8oRZtEdW7JXXAAwVWksZUQqo47ivroJihlog8KzshwfS281FkBK+
jN+eNl8khT5N3uyrsndGWFpqawwOTWwAztj99BL7lUmVIVQCei1+GoXdfpOY/mkB
HCdN4t419gsqGzXQgg7euWImOcngKRniSNJmB6e3eSLyeyxDXITzMxVSeaEcH1wC
DJcQGATXGkDcQn0QZ/+jLWFtB/elNKcesLTY2Syz/XA8anUM1aK1FRdgMeAwPgoY
7wjkOo1kNQ993amHGVhRymwG6sS2o+t2teUvFuvu4eMKREqXCw5gA1gCAVa2XvJA
/RQYdtRkG6N4oMfJUNI6CINTKQ3hBsy2ynSpE/PDLvQI0Rp/KQcDyI0BgTKziNdA
mmhXlRz6DEhHwfgBvJMlR++9kj2enk81i6wtqdKHJ+SndHEaYF1YYYe0IHHGe4OE
i6Y/Ab1LT8usdkwsHB2opJlsv0Yf5NyfR2+2aEA0CcjBPED5LkwoxiAKnHDeB/+8
L2F9nqcSLn/hn2UR8c3IvLPDp8B7ciKio7l7/oiP1Iv7FMqTP6Kwpi15kdR0FKMH
jjUi81JXL5buUf/aoC8LaoOZBOkcdPRK75HPSbCsw3oHHQPGVFoCMwlo5dadLg/1
YBsUGfnW4EyZvWjp7WEKDg==
`protect END_PROTECTED
