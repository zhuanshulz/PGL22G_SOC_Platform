`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vvg34b8ax0ywjdi/TFjUGpjEB//CLfaxeGCHLsb7Tw1anz/ZzgNPhkyJRxW1jODm
ZbcROLvAlfdrNDA35LhKEeB60pWPd+/jc8AGn+rBLsZBGEVmMnkv22K7YSDyFrYb
52mq2pzJQjmtI1cwEvZwio2cwtKXfU8VTOeio3/8RttPOjLDmwwYnbFzX4ls/Cus
i9TbejfrM7UKf9jHKg8TZ606/ZCOcmCO8s/cCvTyC5mwPyLBjT7kACPUBdj59owx
NGm8xvRZF3k39bTC7zqO1GMdndAbEB0904OltwpOqxqfgxvmZA8b/ijs2sQpkulP
Qkzm79vHWKi1D/pFrqPjoUShZLBtPeRNpN8hyCmc0Oy1gFtsHqCYHzP4CkP3HNkM
`protect END_PROTECTED
