`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Or7kRHs0VNC0d1iIL2DquPTR9nzoFow1MK9chhnTrIi4JiqSLod+ELtcb2X8iIaR
423fU5t0jdZM7u71lvpFjaahtf5zlT0GtUBFsIcNPD6NnS7/CJrurBJU0NGJ4pIc
o+G2pe8LQHAr/bVwZJRNEl2JKQzTGpsQUmRf6MoYJXbNtV6KP3Na0SNYTs+gqsP9
F2X2D4v5xDV34r3qz7gNLrwNhRnVDGJdfYOrRKdPH6ghIRNuBuRvLYpQ2y3QLn7x
nt4Aip8w2QmsnNS0QrhnrMo7l3E6zRw5VlDTCFH3dIeyP2wgZ60VDaBQBpOW4jr8
Btlp8nYW/aITLLL9FKxzvQZafOt6hPr7xBMb7WSB4E2YX3GzBmFjcO/rH/9bHbQK
HdybPsMHShKotjO3GUyYLinRYviwR83moXnSXXUwApOMajol5NdTFoYgLZNTBMsA
9gP8pu/vQ7+Po7utvWgfbEt0gZd6xpgepr3K2t69XvnvVHrhWzgqDuODquqao1iF
0jEtHoh0sqVX1kzpMdgHEuKE48wXEyKtqaQY3zrSdMvFRcMg5cx/9Q0avTUhkwrd
Y+ffgpyyrWU2v+7GuMWf71Bh35mUn6K5WdOYNr658tMqL8d91D0eSIvDi2RNbvND
nR2Ke0tjM/1Z1NlLwoI5J4oTi8tzYKTBFS0Ygsdu5nyhdbL3l/couckNFC/TV85P
amnUgdwGX3I2D+Xh5GVomJ5GM5VKbyp3mG6DcJlJYxUAqTg4+3ultPZ5wER2d30w
32UuJYyAkOmAq1XHPp8IZiUwO41A+ZfvE7/Jx7okB5Su2MVBzVZE+w4DmKpcFkRE
V4A/jvk6wrfD85UtQezJqZv5nYtWM4yIsoy0FKLN5SjVa6akDnmVsKly3MUCH+ro
vvWE/4vh4waauDCkJv1oNT7pxab26G8sh4QF4h9vc6ipxJocteAemnvGJuVXpqEt
oSAVzpF5Pb0dks9vBiUmu+YJkkJa5qXPodui7nfFm5WzcoW/2aRBquX0toHwMbuX
qaaoTuA70YKiR7Tj1y6vW2I3HDI0EfiXSwP8BbK+ks7RhFSYCOigKEOMgKW9s5Sh
dv8B99SyuUl2YH+ZZi0Z2M8C2qm2tx7zUT+ZqbL7YibAaO1TUKmuvxvmXN3Cw+dr
m/aoReRUHdrQN5HCMB/cTmxsfOP+/h+NKcOID+BNIde8yBDsAPlDMmcFHvsLlvpe
UrCifwT1Qr4CnKmXNXhozVBHf1Cmt26yzEcuwnLzuGbBFplm/WmULLcmPZmf2S4B
DUX23KpsJMIDNH3ncUi7gTA7IgR8jkdr9aDDnVIcW6qvwT8hd3NVk0z9bwSnQSNC
xiVzfQUt44ebw7eOhuow4I38TaXnBHvt3CHpCY20oTEGwBX1tQOpd42DUvXaizJM
VlesLuD39V+RQS96/6WJcneqN/TvzhhSmyVHWQLiGj4J8uQ+ZraUJOEfKTAosPV9
pDYKAPttDBBBO6Mxjm4nUiWX74IcYpjf9p/0v3XkUKs=
`protect END_PROTECTED
