`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lg660rGLfIwRMaVGub/Tn04VzGpIOpOR8xu0NcpDnL3C2dwPrL/XAZNaxhMLbQXl
ZyrbMHcnX17/3n/ugPyY3Ch0RZvD/LWBT4dICAj2hicnWMzep6lJckL2qpYO1WGw
Vu9McR5oD8qEKVinmmSF0NcVwD2ER3O/01wT+YAs3TRacbBW3ZwDn3cfdFuInJFH
v8uWgGVXmKMyqt7KUFZTHBKf0DHO/ve8pMFMk553eNsVaxrRBHKiPab78rnL84Ht
yBGTNhq62LMoCjjFUxflyuRNhYXlNi+n9h9oiET8YQvIDCeob94n14oOCVGtI+tF
EFomhgmlas+H+9rTe4qLbrUo+pfV8xYvMw1w7E5I0z1EwkdTprXzp0/tkx/Au8pL
lJ0DAgvEZtLRp76MOptXTImXKsAuuTBF4gZpU64HqpQJpAsnH80l+LGrPjPxNAU8
SDY1flGmAmQSXGGTgUUQHQ==
`protect END_PROTECTED
