`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n4R+6eNzvjwqaFwGFAVNUjWc6wT8KVIZZp1aLgQLtenho8MwHqvmJlAK3HrHPdVy
AzWiQKXHeehJdZPOtU8pWHbSF+y5bZAWMYlL87de0tM8mfBMB+gpuKhOT9KDnVIh
WIC2fNLBB8r+2FCxnRWuIdGnjb0qI1LaktIaOQmY/x0OZUxwBrbh78gVWskehHl1
3LnO3sE+qS5LmbLeJgMXAXxTZ5gTc3nawX5QyxbNc/5AfMgpijB39GZ1HTbC1zpl
R991SI1OvcK8zJd5aJo6BHabFpIiRa95InDaEJWC84GnymDKBS9w9CnW9TGrE5tT
SmXXglFJZ3nNL+JbsqmbvIo3KeAXxcdsRjb8vRNY1KvMODzBATEuNEWkT6dQ0/0d
VVRcESsuuMfQzxIWwnrgDNi9MHnl9SchbzevZDitbsCZBsQ5XCxsc7i3tuv1ZKui
s03GGpJqWUfQ0bMxo2CCSQ0HB1AKXGtwmPiKL30JMDhSXUD3rWJtDHRpxwTd6Nb5
dw19bQ2A0RjPRCbIO67mY6baYIs5SRq7xjLmYQEDPrcXSlXcSmIjTnDXnYjYUoEt
Bk75IwittDVZWyHygrZrBLdi9wVkwgJyE1SsZBDBsPd1ami9/KQNlxfR9s6H5mAF
5r8ZuGUFfTQyELwdL/ZWepJLowl9J4p1jkFDOkd2tYSRYRyLzgecWC9CVKFBa0zQ
uxUGie2Lf0vI4m83mwu7C/MkogRIXqRbAfAI5BzeaQr4b0tCTbZxaM+3+aczGv4X
`protect END_PROTECTED
