`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NA6zOxlipHfNyAuw+B3b8ico8DTFk62bIG1NjV6OIx1Zrjp5yVhmpF+TMgY7TDl/
h4upMyQk1rO09W9V5VmrKayicJ7PkSTwwOI82dpJ88wEZG8/t/1vbrXF7iGW3LlE
1NL7NXSjTeKZ5ff09cw5K97BaxsrLu407e4QA4RXbyEK6AUdeMb5yjlzrJa3bnvI
S765uRe+08CjuVk2cgut10i4fbJq5FuYW+7pQexxLzHi3ZNIHqMxiGZXTeSGRacy
U0Qgx5iU0Q9VGqTf3oJs40AviEdMgOiivQg0tPUUkTg9d1ruhSyKGQ8EUtOUMCRY
vRiHnSl0K4R82K7zWyAkk4Mm2CnOEogEXhd720pH68LurG6Ux9P5dOmRZA1EMLZ0
6adxnJGrQLAT0aWAPydlss7wdCASvEEtYU5NboyqfVK516ahfod8AGvooCPATQ5t
trCGI5/aa9N8SJs0n1sqGyoQfgKiucayCQTDrPYK4i2BNLKtR6f27JuT0vAo8+UV
3iMGIni/huLomtt2Q2qnSvqGV9+DrFM2bcSTlNX5V+lMeMoknuuSnSi9WV/hNncm
Q9bqRqHzUOsFS020j47iCLwguOodNTbazMmxTDqAK0veyD2yQpxTrlfTzzrLZGCD
jfktuBWql/obBTFdt1yShLQ6itspEMiziy6o2FF+J0/YRZN5SCkPaUGcCC1rLpCE
lDLemZ52skfId6jM6W5tdxbctn8cnQROlUoOMml0K3oVt78mJ8DjAsF77uz00YU5
r2lZnTlcCBGsfn2fD7Fofep36MMmnqnv/ntBOX+Vbm9b2l3aahgEx5e7IzenMDlF
AbP66o6Dq0yHVzqaPp28Cd86VFbbPdVKdNd/uwVAaqnE2dqkxyAC5tEPDOTK/rKd
W5ma2ovtf/mbnRzpkQpNvnlW9CGc6WBs8kym5VIAsvOLVRbcvrYp62l/piw/UjIO
JOCt4I8vck2oD0xU5p1ZOFCcfuYPUbyOHPidp7244qSPuqJt1wxp3+FevnppAGnY
3Q/FYX7eWPce7D0tJ13xacc9yQabsLxEvNZEQh6/ZBWJdc0Jku/4NDnEY4XSSsuC
y5LKJbb0EqZ2fDL4iWsKSrzAS7ME/yzv1mloXvvz4im+OyokEdBdfRnKwpS0g+CB
xiXRJxSNJ74HJ1QlDj1dqmHOm1hmsqVYiqsPDb5mDpC90P6uFiDLZP5Jh6y25TLe
Uk6ZDhlwYyVY18BB7nD+4g8jMMQsxX1UoYJovwV5Xz88lJqER5MkwFurJsJbRpR7
EkxJW9p0Px6P4A9yq9uQ/G/5nOLmnFuJ/pidg2rlqNlxcbkaZA2mqATpI5WbrbB5
ve1WvJIoYjUiWeggxpT1UFGbe6EPCzbuPziv3Ac79PE7hCVfpoOK94HX95huuRvM
pgFcxb472qdCcyzGj/8u4sjnLIG6N7XJNEhk0YkVo2jmMtnNj3F/Q6r1j4BE5WwI
/gNIIIGxyueQrJI1LqzUvE77MfLAm+Fln+Au9Ggcu1eLh0w53oUK5iXm4CpbGmSG
/t7JHGxWlE+Shc3T7WJd2oDXfP4W6j3btoFS4J9i49cP5ZJGkztE/sGJAUk4YSmL
sZYfO4OV64IzrVfpOC160dkFT33pUhnZ0XnR+fTu/BFfx6NmrcqqVjrVUGJpOYrB
52wE1/VkV5jIoeLMK7qHKlqjFe924QywpKfVN+8AZ+edLzBSIpRk9Up263IDQRoP
oRw2Zr4PZqPF+2bMYIUTRVpHXZ1OA0Vo2Ox2kGET9NpA83kcavMiSQVhtiDUMJqD
DbZfTUdQ0DyLqrK81izknCWkCehU6ukUl6E/LnIYlRaV2WlV2QFzmNe6ZFJVvvKH
bEi5ks94ZGqYzfaaAewu/jchw1vNLUZdMRSJVchneBuNfTlli/DEGrm70VWVoX2p
r8gy0DhQ4i1mSmU6RQqxTKuMneZpJ0gVx8BjoFpsY4nrvHfJUQjHnJX3nquF8f5D
i+VMnffRMZtb0jws8FU5Pr8c2IF02S6ICPXDwITCSpQEIkNYtTC3aWA35uq0cl+t
cw0VKOTVCPltOhC5yv03mx/MQq/ZHdwBS7taTS7MAwlBsOTZ4VPL+LT0pTQdPH1h
Aw+f8Q4xKYjawIy47XkFVAD1Epq1D7PGNqWWmPIjWiqo8tQXFp3Nkbf5WJ/x9aqO
0bHG8E+Uz4rMRDe/2SQtC7MrpgcMyGkP8XmA8tM+XSwYRY5gShuQUxs2U7Vlo/IQ
RA3HgeWYVWjLtXSvCuX19tvFclEmUpuhXPH+sKL5wu7qNdT9dVHjkzvPC+uxzLH5
kueov99NKAcvFIHNIpQsSQeg9wKxGLraz0SdPeR83HSIrqGo2cjMN0aOhwPw6EG5
zfuPQQ70crK6nQwX6oIoFHS6yEdSH/mAC2s7wpay5ruQAjVXLYKfo7l3y6yAS9e8
yt+RWWISIvDrrr0zXkbddp9k/e+X+G9yEDKHjuWwwXi7xlCx53uoOhx83yXjOfVU
MwHcmn8ZfdfHM9tKDVAAl5c+NBkFa1ZRlS8Vuy8VdD4P3c1PJ+ra6QhEqTGU8jiD
RePsp4SNmAOiaHt420loYAk9Z+PFPbkgrr8o+Yi5YLaRCIDzPANujXfFpfa54FPG
+MoFDRCQUanrznzgNRahr9YVeNk4ew/NfzbyXvLK5Yl03cHqKt1+DEELFmpXe3sN
+ubdmerVOewoyPDqJlsWoixKKQqrbqucIn4XTbgc8NlhWpoh2inSfnxSXfi5PIen
L8CmVOT4aV7x1ceECUGynGXNlrA/v718PyKCNihEtP2Uejq8u2xwUvD+kOkDhj+m
PgNtbqjborobUDUuFns2MsF0RiuoJYppJRwbR+3Ahq36t4wNSuf7TUF9Celv1PAo
mosjSjr2Jfst5R9J/bamDUiZXugUJzlsdXegnQPSneUmBKX2DTxT6Tml7Z0LtJ88
MxaMrvIoThY2PdAd83LGV51ug5ZXfDJ50hglfIFE/Hza+jhylsC9NEOKsImwcBDF
1xyvZyAwIvhI96j0IJady3oHJq1zdmCW4K799OG1xyul67vcBNGlyichu+81P4v2
T1Ta1qZDArSyl+X7O1z7f6F2aRaWngpSuANCbN19G3S+m8hbWa+GnDETXTXz+RwL
Th2Tly2TVXudCgpaTo3t1fbG9ru9vAKLwQsFExj4RXz5QXkVXdeUIVLqF66UJB/+
OYk3yYRnSQDPDMeVGdlFMjktFJyhNPR6WZUPW377EQGykHW93rn0b45XvDBP7xgb
N1vbBPqrPqN3aiouNF/X7LWxATsCOkqngm6Dvao7u/ffuLeZl6iFlzxVC9gpiRyn
94/g5MTJz+TV7tgbnyMdTHTMQRzGLb2G0Avaz1TF4qvBygBNuTJrfySGC9a7/8VR
yAG3qBXpsAb1e9VvD+npwiYuTcxKYfFrF3LwQZhrle4JfR1jOjQsoV7snKTCuJJI
+esev7NvpqDJjhiDt2kv6KXFLfRxZNO7ZRwzgjB7sqSHB+/K8vLlBzdhv9nQTBua
hivfLaEnaqVXvknv4/vl0CGlu1G39bJ0pGMRLIug8QVEOkTcXMWNKVdSyR+y6sqr
FRxV6MWtcyZMiyIETvbTnA==
`protect END_PROTECTED
