`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r445BymMxquDYHCvNzlZsXmVEBDtGXiHem2F0wSBZkUzir+lW7GMbvsmHZE3ZdbG
5/hvjLvU7JalnLorvoHQZ/5mOpCDBp8y/2eWZM22IZq1GwDY/DpninK074WG04Iv
3f7Gmulro14iOKuhgZpJvSgCYeikMCZ73lUKKum+2yhlsCmuFgXuBiAN5K7srZBZ
XMdDaFQeYNNaOF4qwPAwRe0531pot7KN7x41ooK0FzpCkRzicAt32GABiRoFcfdE
7RnaFGobvGlT/GU0SQ30y6h0LTl6yNwp4BbjGvCJs1XN3icXOwAoAaafXFLVcLGc
+yWcjSZrAK72CH8sZ5M3TCIEKGt3vO/KN1yq5jK6ZlRhz5LmBh3CA6/OZ6cSbhW2
8d4L4ptVDGTGQ7UYilbU0P1unbhjSFiAH5hZoFW83Lb7I8wz5ztm6p1G3+vwGZc8
C8y+UTXfDlcuAMuPo3FZReX18Q88QoKiKyEohqQnoC/aHwHsdKfvzow9GZOU8L8d
w9u7C5+4FUZ6vTSjHivdtIR4VpvoDC4ub5mBeCWS6V0JOMXeZ8m98kVXKn76HCnt
qjAO1fBMnjBOntkNjlkT0g==
`protect END_PROTECTED
