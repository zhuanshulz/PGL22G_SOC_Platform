`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNxQ7Rz7hoK3+PKNknyaKp2+Jy0UHIyooQC/qh4nWxszfaG1h07xnfXIHc7uP+f1
MJHVT25IT9OmdTHDZ/rMTH0WXx403938ETvtzPYqToC+KKQEJ/ufkSGnWfiJOS6X
p4EES7Gg3o7QvdaV91PTR1uH7Zf4SC6fCGqpZGqEUOgAGXMiO6LKQrz+VnZp6c8U
OeRsW45glihwx+gwUGTp+/Ibn/8ijZYfXIJKIVh7YCv3X3wtB2aKMrCDsZ1kkzV6
ebTe84NnGKVvo4FlwUL9q+Ext506ak5KaC60SfYrW6nRUaFxV6GAVHmfvCwSG9Pa
4IB2O171PIC0w42xGtn9gGdLwm0xlPdMYHSWtvxycR5vSv9TqQ+LqVTgPtgAb6jc
oAC8GuXPzSW93Vy+rWLxKSU7ZmajwlMJlKujzqQR25lXfTrmLNKkXK9T9MuGJImA
VZ3SAfRXXCfl+m2ufuM+inAonk198PiTqPQT3SKuv3R+X+g0PCyjMv3umNBnytIB
uzfsdb5rJxmMvxYUB3yKw2ftNvq4kqu21WR2Da5iyx1aNWi6RuB/idt6Mo2Aomdz
XWzd/sFzUvr7rlUvO2WhME7VLOgWRyC0W7N8HT/B1tMJbqX3AV30iAMcXoQH2/36
HXkBnTMUfnLf0BnmxHOVwQTBPueJPz9x2+ghaB91nioYAHgqpyv9FMdZe4tQFVHY
6JxZXw0tbS5WhZXXLTENSbwZmw3CNh2GluL70CXEeuK8nOgkPkeoeT/HZzzQsT4y
kOzLYPOMP1aCFflaj7nV1wb7yfu1vos/Q7snYYil7w1OfPTKkE1S/rOhH+W0K5HK
TL6stbU/osGbzSPKU4zfI4pLEKha4z31B7u6l2YexGff9ufuZUT31eis0umVB0yt
ts77xg1GIjEdOYReOs4D3s5r5qp0ymrKWjiF1txKUSXqGED/0yG/tPqLh2nsHLdo
6wSismdGquuYvOd5LrBQBo1vUgSzU7dU6SnESqho5WvwwD1CzctnVkf/FRUaZmZA
fF0e7DY/FbYhlnbrrIOdVEUFL/GJpg3nbCXzOslik5w=
`protect END_PROTECTED
