`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/XdNMKDRbKFFVFN9TtH/AKcZ/wZRgBb0CaOHwWdqsfq3Mnu+fxkZKMVwTL10+gAG
InfpZa4Ri/jIqWptVlQKV13FPdAH/KMvQ/jgbU9NkzpQi86BnNmAMugVpZg7rZCl
Shfmpy6HHzNofXdjPBLwhnu6cuQo6ObMLmFTL0BUZrtUyzlyX9R+9/5A3VuDfvrF
7JezukrNSEuCT/cRlTvqh0XfgMCUID2MHQCd5cH4swbigFrkSeAgxR8hrT85cD4V
sgjoip/p+TaDB19cuO/pzrJ0Aq1DUk0xjftj1RuXoWQxlGjpImKzNHhTpYWhcOFY
BTvHeSKE5GfsM73sjHSqXZqyzcqgMN6JTEUZaaS4uzyxmjgmC4v4GLtwGibSS+TF
wvywroKwGinVOAzR9ZQVfXtxZMjwCIjGsxs5eNwuqpbvzUxEgi66By0B3rCnkzPJ
sl6ANxxphbfK9S+IKacUBTeEVpNCLlYMIEYlRIuAx1qBczGZlIIsMCFtF24Opf6G
eJYSrQT85depDHUax5QHeHgn/rMu9Xp4BkjY0jZNYoJHp71Crlq++L/P1kHAAsz7
JehZIflbCVHsK8nY0ZrUTZ08tH/jNOaN0csNr4WwOOFCXLAdxwr2hLl8P2u0Kp/0
SH1VGnHHJvVZiBYpuvugkn+EZ1+S8tHn2zIs3m2DXPGJMju4XY4Bg9vfVeSrR5tg
VUXKQiQm/dir8eF9UfB09C21d/93+T20gFteWffltNMGoWx2dn4bDtygSp6ToQ6q
MmQa+iGCmwJMOasB4OfGIrkGPD9C5H7qZ4RN1pr20gR5yAVr9aYeLVqzyYEGUBt3
3uI03BJiAvYNyl6rDgQbQ3wuDlPDdbo5U38HhGCLSWz5g7+7FXWeDDOn6Fsuhpx6
6w25YeOFXwoDP930jMAVez3dHWpJWyqQrJJhWsO3B/jplwUP61sE5OQO1a2QZH7I
yFuTRZDxl7YUH73hKEBtJ09v7tM8KwXKHpOZA+p0ZtoZx0HygU9N+NagW5YfRvdZ
46Zaq4QJ5b0KRDIbnhKrzP2ZqChxRo6g0kPctrBkV2/a0n5Cgwo3xDwhp3TE6sth
nI/6myZ2yB4OUNGGD2GhhtEQdjonmDb9gkvQsoXJRpSM6Oq7tmdvHeAJgaCyzne5
yBaxb/L8R5llazxiIXziGx02hkRMI3Ub/xeH8iZAO+7y9nX/GkKclT4bVwYk9UpE
n+lgpHmE3BjarsDtQyAgDQ1Y+41hOwVOiuhO7q7bGouzBQxLZGQcFwvMj7E7AYLx
6kxqJBH4uo8DJlLV46/zZU2yVpC4GBvAwkgLejiy2RpZMrMaWrPPwBsh3GmCGDb/
SHMy2LrguJFvUQ3zwZicSkGsSr3gq71eafCKYO35UeX6aogfoYThQKluvgoOD62i
gm/72AN7zzy7rKo6k/Opa0wy6RNKu5csMwXjrqlaOIdzlnaX5o0eKywZsTlOK8/p
bud1Eva6erfkVVkcvM3cSaWSKvIITgJf1FdwR0eAJUbEZmDJ5rlGrfNEuLd4QR2f
ktst0kBuNThMaTYQNnbnu1FOHcY2a0GhgNi/nq8ofrYEcPqP/jEgNkFChzFrsEIm
j8D1cNmyWT2VQYMiqgaZ7SJvlRPBsrgGmdDTE96ZX4H7yQGCgGjAM8JFh/ZIqDSG
6r/e7xJLkTM5U4sFhVrK8cpEDIfHMa3BeiUzkG9/sUm+ESRvh7haix+EH4qEKPBq
H9mUHYsO6kQN3v94SRrLXY7sRA3Y7Rj5ohZiCYgwWVVCzHEkiyp62qGuwzPp5KpJ
nWV8ZbxnHi6nru9CUgvvUvck5TrrqbKa18AU8Rvgcnu2dOojQluTSGfBXHUtatjL
EwzvOIfo9RPFD953eFEshg1SzlbGTNAc39+zclBBxlAgRxDbWkSLB9LISFtEIh28
NeA9xVAtuxwzwu96BTWYjsFwd3DjoHpStUr3wN6cCibVnmVpi/uyDVeR0EJ3Yil1
PWQjYi0ceRWuFaW6KDjiXGjtQm4bGb1qi7j9rFOj6RIgefZn/Cb0Kuc5Bpf4tBHA
x2ICm+zR/BzS+yC1qJZACqpb4/kKrwFq67sl5s+mQOaK2eLeGiGDyJbOW9WA8cN+
RRhHHeBugRpPmGkB3sN0dMkzzCr3dOyfQIsR9/zBZVg1/HyANzVT8xWTYtCuqDTL
SP/yWYipjdwLjjmWq0wDD2HKyaYsHy/ZSsBse1DJNiuBgKbucY7Yo43KrjtQP0yn
Hm0A5HflSVKtm4HYH/KvSX6LXR//lQwEa/V6lAUMCFJFbuBdom6sEtQMA93P0f+6
sXDoeukvBrEvRx6/H9SiXV6BeiJxD3YT1XVTIUd/WyLefXETGZThsbXTSMVvOZOx
TisUNiOW7mY7MxL67xg8oiFD0QcSN2oAsxU53zc7ZWO9XvoFCNmdY/uxQG6In415
pfuP/Er5oac1tAf5SrMArvnyZiR6lRlZjtAW9UC3QPISiXoyVOiV8xsLXskn51Hb
lYNUGP0mwyFirfqUrT8NpzYZzhYA8da6b9Lj1RbZbJVFsu3VhyM6dVG6RwUIdStn
ImUcM4P/mWu4rVa3fDl2D5A8BkY+x4f0sub0EqjW+h1JM5F7eB13koDcnnDPJ2io
vDKGk+EVFqIdAxNzBgY2GQjBPPHYrU/CCx4Q6OKkXe+7eJlNUJma9/H19CD5Jysc
J4xbMgjthZZepUccjb+FtmwLWW6bKiv6u6AOIsawA5hWbu/F4abq66f+5Mfzb5c0
Z3r4P6sAFK5i+jfbNINiWLg4hltCOEAxQEZ9gHwZUgW5YAU8dZjl53+RlCLmcp+z
y/lKJbWFiROCuO7Jm7JaeuCwt1Gq71WAsLrkDGYiJ/nVmukSTv820IfBhajibF2V
YDS9m+6RB+lTiYds5GkdL+rrE56ekCZulfU6ZGssZKK11KuZ+joPXqSRieAZA3+i
e5gfK5B+DoP1pmD1WlzN5VaQnLK9XXaXDLik53/V0EgsoLZ8vAaOUH00ZSXPhYyN
OJ56Ddu4babSM1bB9wXJgwboT/La0fRA3G60DMEbzUnH2NaYKGw0gVwPKNuert8w
IccsEf/v0jL6aiQx0pWddklQPIaIKxTlnqFidivvrkGIpOBYtU5bImLIHn/prVtT
Vh7Q+4TD2VzLAUHSesrx7PhXXywgYnbtyFuXQJPVlXxGHY2JNuUYunS+DwqmVUjo
5vEu7vwLJIbPTsc+G/9LI+QqUpi+Jk7ugqKg5lYJqec2I4yYyTIahCmjXXwArwIy
QyUlh0KUAu5/ZRyrZwVgh+0BCxxF1Qxhk66FaFczNXBPaK7O9c/ZQ6WxDHD0/aHK
KYvxxkwGSVi+Vtb6G3ZG0/AqR/9r8zHnQBMN6LIvHAl1TfhOllJGUUqDM0CqSZ4K
Hd1sW6Jn1XLrYF/R2FYzEehF931C062dv4edBG6h2oTdGcgs0ir0mlbEidN1ol5T
FzNvbBmLZpiiLHAWDaV4f+zkaQg1SNDzhjnA/DyBbjhlyCgRfspN7LtKrgkCqPeu
4CVplkiLoSK3T3mVb2roaGHxKE1Nfo0Esn5ApNTAaKn+OvLr0EhrLwtrvoR0K9lC
0IBkloTaxUsPmMMICrptIDzCSL9UZvz2ShOerlOeMVNDN4TzkMloSNaJyHa2IFyn
dAAAfpoJozKv0HfejBuBBGoqrkC1/pxItXb14D+fpGyyDf25+E0SZ7ORXz/qlv3z
06RQ2wi9Z6PjqYGGdp/lg1sjmWyOvCzAowo+eYq0F/j+g0fiSOJdUPOjpJNIi6Mw
E+rFsh8xY8CZXIAk3K21dWy7KhWLYs4IeBRdptrGLp8boMXXGkBCt8QsFkYG3jOC
EoIAbXxtyE7p0Mgxdi6b199C890cqikd1+qFJC/yk7+BXsZdKlQ8ilb3Sb1T0FI2
P9+CuXWJbvnk/AU4+OOFwcdluw5T+gTMpqEBupBIoMBmdfh0vTu64rgx8Bbwe8lK
t8t+sJGUqqYZHOyru5rzazQexWWTZQNfPsN1GeF+o4Uls0qoY00WPw0OvkszjCby
nkeQF+G1OG/4zqDlPKRL4/AVuyGIgKr43hiX+uTZlTsxsm/KlE+Lg2sqSKpwc+Pz
i7Z2XerFBAY+ul/gqqd+P4LTCxih9Dmc9MVLUmA/QIy+vSyBehQeGj1qd4uFmw9A
pRFGX4qagC2yUskFmpWIvMElmSzEzWDF59Ttv6artRdo2e2GS9b77sWZ0lsR9rpP
5lIc1yPc85tREVnJUb29wRAfMlNhqqJt3BMAf0GZBlepd0Ecoufd2dSiw3N8Ds/p
8JzRFAftKJfhdosczn7uSQVS+9eEfzMU3csdqQdk6olh2tUS7tmHHa4A6ImHiVYz
aMHBSN4PCYsYnshzYESYiHv524ZFueOq7wuLoCxI/2mqoMS9n9RNJ/IiD93MPCJr
k/8Td+KoEFr6hdBQ7ERrZv2171uqbvEP06ZolpFkNcLQfvvj61ASzNQJ2fV6QNYJ
tc5otoTW/ROQhOxu6F12aADmax2RBmfjfG66BBKOQGY5pRjiJp0N9LKuuSBm/3bK
WlcRPNkVYEZF+xS4hvg4zqBnCI3gU+VE2lFZ/2yVKt4Z0hlqEbiobBdFHxvnqVUO
zf3AWl6nFua6w6OztRTXVYeK04qCat7lF3cOkzoCirzEDjL72XRBxs2CvahcDlRW
WprwQ45EHa6qw/WEOHaUERXmRoHu1Pv6jVgwEwOwXZFcgWDrNoiLJTK9Bs9RRf+g
z6nXmpUS0G2p6bKuEWD7hLC4brUWgEvSTEzd1CmVRGFxkv6SkD668dXbGbdpseWD
hWlWmYNK4zARaroXX4WHmbvxeFq1M4PvaXCWds6AJCPygRowvGShqKm+BzQxQ+/H
1DarMuUm4Ybt5HzFZX22L17qxB6pwROAqLLiwpHGTyqKGBIdwtPFEDdE5y2zlCda
RPFgoU3qwaJHuaKrIahQfyXn49DPkTcf6nqDRWiOlHFxOpPzsBUeXvz6/PxvZvWe
y35TOxRixc/ra6E+EnKDFNlq9mTp0z/ytkh8Q8z+MnYKmNlgnw4goGk5RyorrVM/
gLi6CLzo9To/ckJjg7f7wsHpKd4iW+qU6TiyV6sV/0epkoo3mJCRBAQO8ssxWjQS
QqSN6yaSTHRbGwkqMZ7x8Ap913ShkiWFYbWE9ZfZuCzPTkrwWpx69zjLP+pYOY5h
73qAn9su45v338x+oYuB+y458MSIf9vvu/Ie+DKqaDmX4FgVkvFLJtHbDank/FEU
YGgVhf62W8FoS0+oNs3KQ7WCPqXGtoS1AL4qhF2LtMMS8KCmrfcs3xzgPzILCfeC
oLD0JZ5KoFJS5IrnJDDGEfcDZ796DTwcpXF9MpqrD13aDpEVTj/B8w00VFTtB8ni
pdObhMGaXfBGR/BlsVbRiPK0mXKQvVBcW2lNtrteZuC1l8TcQN/T6y+N9sPn7t3T
ZF4FggyRQFpF9BFvkNNy/9eP2WEFXp4SUNF4hIbYlfDUNsh6FqEXTOTARUArx8RV
4YawOjwNJVDXfqY5Sws8+gg+3UW+qWUH3Ilan5Ut2XIiYndAUdhoPfE6g1ZUbbXT
z26QnGxmOovk2tF1aEGwHPRVBR3z+pZpA914GCKinIiL203sYAyzuYjKekz0QD9H
hhs4phFqUG2xoh17heXy+PciyqyZP2kCOCT1UYYX+0FPFYPaW6EzsyC0++2t2FSO
oKkP4ku8zsr26VS0EQovNObimGfq4pUjhIKKJ+iHmPkieuNozmR4Wwqle/62LZ8W
aQEdjRofHb91/4wn9YwiDBsQDc9zeSDHsXnCg2UuAYTUkuEzmwLFqr6SZakrWiMU
JeVTyDJofs6nBiMhdoNOWzxUnKC5rlruhW+IFQk3+0ySDGXpXT7CFQn/3YdtZ7D4
uYivtLVRyxVAcT9R2T+7vAd26FOpQ8185rO6u9CXEbziDyKnmcGLASOuwVWSKmiU
qerEoGmKhaS5NFj3g9LObJKnSN0r//7HdvReZb8m1WLj/x3nje1Xr9SWMs17qgjV
iwrO+aBxfAPqxqBXxvteyXAEQMdAcoEXBkIKQmOXwg1RMQdcUPXVRPwGZxcnd7IW
Tpn3uJMRIoio5ySWDYMw/som4pj4yacDymt6bxyZrDzTEGLPKyZZL+9L6d6UJxEn
BDxgtX3KQpKQ4tkl75KHHZuHUt7aZPJJ+APAUC/16dkNhf2jfrRk9bMnhU/dFOov
cb8yBy+UDGwIPQKn4ZwINchoOmHR2/TI+min82adAWfk72+Quco/BsDTS1saR4Wj
0RAFTwigiZTznalN+jih78YKNudhUuPfB8K0nTOn612ddfbE1R+bWB7cg/xsDib7
JgSPoJkte42m3JId7cIrOlVEd9RQyxrn8PqBYFB+zw0wIA0iTtk0UzkRdzOlIRme
OkuompHOVHjhsGk9Le+isaIQiOdo8otQSbNGFy5kdp9EFBy81R73dugbQxzyHKdl
NYhJF7S2iXw+L9oGWHi5jOqgolmeLaRaYOJ71uHe0zrWIJTBpzwxSo3hkPz5zLw8
/MG8SRD7XnXFj127EjHosUpumQONdbcoFRyMc+KK4sA7HGImfwqRfRjWygR34oCb
gJ8EOn8S7RmaZPhX06suLpZIZEVZIUwom1/Zon3Z63UbQfVPAn5fZTGm8AYRWS9T
6pdP02V77nZhJGX+Jmh//UNxDuCr2F4Jp479QvAuWk3UtO2PLiDYtXrx0K2INcK5
WksCa5VLVklur6I4R96+XVqHxvgQJZvwfpT3UPcPurAq6Fl7mqAPvGlDu9OYbCcy
/FcbDhWpamE4x6h4S8cFahMAm3hWUbdOD52zVrnryfvmFgX4zOartIOsOx6Zk2YP
2sVhHarcxgVPMFKIKW24KZHECNPYUZ5HtPTGnJ7FEWDO9e3qvg8w0HwvItlH8Iot
jhwg60bU/Z2TQ5Zp5nXZERUH1nOXvmIlO/vNoMnHVnceKOh2Gbq4oF8OwVvbDhsI
0CUqC1l3SHKsErPaazXMP6r0DXiSAPKQalWm4g1/7ssQi04reXC7MnKIKO4XaEXi
1002bM5WhekwGrWDbwiy/PJ2NFz+lr94+1IUcvs3xRzDy+SAkH9etv6yBKn/8Gcj
ty/hsVfmsvJRG4i9F9UOnCr2s4ekvwd2E9GAHA4lzihNNYujR4494ly7uVtO4VPH
eUlLTbUNGFD/Ev+IKj6ikuo0o3GKzQ+qkA3IZjQbWHfUR7jbiuJcOawyyVWZwxJa
Q3iy6JjXfmXFcNwJirOV4fn5CniYXTkgvESfBaw9taDcVq7baPJLyxuIVLtYIBAo
nku4gULCmwi5Q3w1F7aRpsXUleh6hVU8MwcZfZ1Tbsr2dN5IgpnRs6RrBmRXZIke
G0SnwDi7XwfVAkdbrrdiijk6+afOohNhJz4SYiQu+zh+Je9CFGa5JwTwPFIuOin6
t56G+CcVLxl6Jeu9h3E48eoW/J/WMsLFrrQxYtV9VuE8Kpx6aPSvgSrd/PT+RvkS
8tvU6hoXYomqHgy17p8EKXmEkB4njQJkth/XcvR2TwNIJpZ8ewZHIf/abX/1S2Xf
N3Mm4TYSlIeCyn1e0CZ7M4Zda3/6pd5HUNtMHjo/P+//XYpJvaWW7GA9gk+Bof1V
`protect END_PROTECTED
