`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FRp3ea0lmYhIrJ6V5WJ1gy7qFzWFu0izvwQUjPVO1BMhrlp66icktrDbuuk4ZuPh
7UNFipKzJXQ6JjdcStus6PsbkVoyU7UIpGXtNk9Dj2MK3NtxFN7EM7fBLSbDLxdM
e62O+C14VjnnMk7eLSIKLIqu3eVz+lPv4M2rz3hVbsgqbiq14kt3C2uVIe2lC3xD
Rd/yz3TcAI+hEj+39kYnFeohaA6o3hZkCdu4zyA0zNRgsErOpDhvNFE/Dm/BJ33y
u5KOrO9Out8GRMgD4v2qtUbDWjaovpJqAeHTgmqwkM2kq8vC9TTqZ8qrT7mGqPVQ
KG2EbgZYqXToI70Wj4TG2wTZB2VLxXLjoK+/A1Wl9OqWOCI2AADi6gFKuKQYEnnZ
uYGPFgbqCi96gurnUv/CZaeidmXq9sC9dGIU7ogsJCHUioU8AkLgNhdJPgwalXq3
OOnxG/t7YnN0U4PNzHYbKq9VrvGmyrOSMiIs8VP8XfuzLxdHwDNj3+wz9kDaXGZs
qO9LxZ872q2u2AdhIMfJBSzM7ZBCvIEefFoDqmPJF4xznfRuTBvl3UIKkimZyC8O
/12jRg56RmvfQFD6gBqsZjdTBHr6n8IBUqOZt5INzCL/0FfgOotjzfd4crKOmF+T
+cemFGt5RLbuY7JpviHEtl7JPEd7sjVWg1S81mOevoSvCs0bb4aRuCv/yHAkvwMq
48gOJ76G/3Wm1fhEBcLHrwODFeWoNCKgwJxU6sOuW7C/4r2Hvh0iEbRlEvfQqog5
orRx49g4mjOOgdpb+fgPP+k15XJjWzGTxeM7da2QSx+PQSzeKMK8xdqpT9F4gddo
VVxC/AEiqjEhlm/Ljr8DgnFOGdCBkXlu8Z1tfBx4uAAbtBLmlhzSfCeYt6/YIOp0
6LGiegxn3xTkT6WA4cxs3iZ/NDd/TomrZ0MTc69R3vi7coLwqJ9tycUHi+9dTYo5
u3zlqZ2qKwHpHCNfCTRhznTuanuVs29b1kFf52GdoRxAmp3rKGTpQNGFhmDeJzP3
t3dZWSkMVfJJxex4BDITrxUMHWKecYYhn94qkhLBxZj9wxcyL7kuuC1WY8arV+uA
3qjjhS0WpKAaT4UYuVc9MA0KAVJVzrzTAWgp76IakyBovav2sLGKtr8gU2tQhGTm
O08NtelCrKMZbtzkrjvngLUrigsmIi4y5QXKMd1rydB9/jCOl5TfmpuckmQM88r3
8Bumft7gP38//rLt0+0fAwZ5wRrhiRMu5Tqya0JE3t7go5ygUeCCFECusfX0LHRn
WztzWPGS/Zk3q2K9ks9+a+2O28UD3SkXSWUBecX9zXHu+SxN/3RWBJm3BUkbrMLB
QXbAPWzwiWMtU+dnYeQiouSv/Yt0c6wGYO5/XUD1fwrKid1eiuf2epG52lH58K2D
EF/GHsb9I/y8rboxcebnBr9VjISVYmb4d8dExgtIeUdAHK+913o+JMo1Bwxg0qU9
`protect END_PROTECTED
