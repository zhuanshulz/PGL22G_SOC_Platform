`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uzXfUSEodmvg7l1yJCDnjpwDnTHFbPKr+CrXqYJ3UpCv63PrA7FoCvzbDn6Jtlqc
Tnwd/vuVHNjgN78VwTyTbQy+YWEh9ka+9uXGGofoxNGGnx5YA6YSwgafWpFUzLzP
/HeoINncf1r88isNKa1G0gTkOK8NOtvlAKaNARVPi+ynGONsz2uiW88E4NplDmh2
2uSyi+cktq2Wl8aDPkdbaGX7DWjcyVGlADl/7GpqfbXd4RWKmwAxetpuBVM9CKhH
x6pu2OeBDdPWxHGvkQcBOGc4HSBddvLXFYDtNvkUDqWq5pt17A9VrFpwokOR4qG6
4XC+dsiOBJvqApZ8CakasBQPEeIzZIZmx5TN0Jcg3SIz0HdkVJjCFtm3vtKp6o39
ih3JmtbRGG0aaCGWuSa6QgPFt7I4/qiF6807YpCAPDiUKjxgg9aXjXLrEgG7rQh3
HJ1NnSsvTlaWQr8BCTr5En431L95QNFy+1RP2DbGCXoAxFlXElPRzRXo1Y8xihq0
bJ1GtDePMAQNIwXtEsAb5YTjUVtphf4WN4bC2HafIVJoNKtgHObkmxi/W+LGRuW9
Noid2oPzWLlI5L5ZF5BM9pywx1V6t/LvjCUHGmIUGyI=
`protect END_PROTECTED
