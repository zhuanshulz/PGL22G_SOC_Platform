`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TseQRf501/gBNZsH+d6rK+Lv+DmU7znhbfv8w+JRlhtyLPEjoYSJJvhDKWipSiGk
k5nwAxCMqkOgxnDnAbPywl5Hz7SxvZ33lVBXVtYNdUg1Bi+9M8jrVnpmHlc9Wbgq
l9adQqLcaOlEwXJ9L0aFnK0pWI9JBR/YOCoLf1k7H+ZgtSyFTXxa59KJjavqrp1y
u5wdN2bj9g62Pi77ZtbcY6UrVedBc5Tkapy+kG/j50XcNVSstb1DyoqJBH9inAxY
xeZHXpz9LzgKd4yJjX9s4Mibzxduk3gpD0nI6DBz0EvDZkh8KwXmYTWbD8nzzuMR
lhz37qQ1G9VYv2uZ3fOKzF2nU9aETuM16pVWM087F6myTHR+g+VLARipvXLN5yw1
xri0WhaexSeebtT3OPUw5wtNJE/c5w0jPsIDvsRNFIczPg9pGajq+2so3gmHvBi4
FqV4uccZLW/ofFQJbwTvSWHt565IARS8bYtTz2azR1uFZ3HvJ6iyZbOZMc8Tmjxx
W8EfjhXaStzj1OrSJmlrx9Sdf8+JNWx6EOJUFAy6bLROeYFwvzrNnto+NHVg1iiI
5KHqdcAxkFcpTqQG230GZCeFgsGQ6nwa/0W/y0yDcgZhZty6uCdtRogMT5iT7QSh
ncBvlSSzLDdZimRPvLidmm4CL+TLVybMdlHGQmFt/r9y/kjQ9o2Mqs/9oSfWTc9C
`protect END_PROTECTED
