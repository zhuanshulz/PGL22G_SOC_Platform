`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FAs+Ch0Xa7Q6t7XnXbc+yHH/MCvbJ0iaTwr/cTrumN/pxdyU9cxBfjAE5QKgV0kt
vtkIprzjq6NuIIaVa5IAxDby5hC1YmhqEMlKwLLiGjkkFLqa/YIQvy30ivcqu2qC
DR0ZxLt2n8uQZnl/TxcPj/bdXQxi6UGEx5+XoBOlj6d2YSpeJ8nnRg3PidvSHYdP
h7ZaAVJevRKkraTYLEx2Ff8o0G8X6k1ayGy6eSGaZIkU0Tneah+XMDWEbXRePJwZ
DEItw+fFXFHbDzJHC2olCcQajfO6SkIbhR4yFZnNMpNBkIwM5iA4lKUdIhKSGRLS
wNoUh6LLHcE9Vxa43mVdCkl7zBd8peqz5tIoPE1lPdB4H4ppycjzIglGPMwnhVZk
lPCixZKJyWUXXbHKeYJ9gqiiCfZbFc6jh3Q6ZdPgQnB7a91D2RYMrBX7hI+UaVsD
TXxlQR/yReOmhLBPzXljWMyiiOvo5xI6oq1WLG804S+7ut1OvgOWCJdqEGwT3fj7
UF11uH2+rgx9YFX5iBRuH+VyiMFDT5ioes7y2q69vKcQKqV1IpvVfh8dFduhRBr1
WyWayJOdO9SMOG90plapqYYw10fTZY+uyS2Us8GU5saRqhpulS204Jk/cEJ6SKTR
ekrUVxCXH2muxubZSbvm6mqA8qaV4sM8K3LJqysHHnipLPrxMjrlmneFE4sHdxMl
wx5gO/N6Z20r6TJkGqJkaMQn2xZXXoM/0VxAAWI0MQt/LtIvneXtUT5r9UAHvfN0
DSUZHTyGLxWEfyjysr0xcEITtVvkyEIonG6wa+CqAsQEIq+4pPpp5uElJlfLXA/z
l8+yqASsLBcuYZ0+M6omGTEKi99iQZsO+5V0kCymoBHZ45KP3XdfWkbSAxSSm376
27eoqjigOa41Uiv/I4h8bjX2Bu9Q21dwg0NUBSsFA8aGXINIZ6IvWoh6CCv7D1J9
RJ9A9ypyB8YHOSip+Pr6/XpEj2NfZHBgzbXrMfP3TcXB75viKTqfzwqrjyTpxxax
HL6f37vSgdjkc+a2m8N1oB/kQFm74wjtnJ84S8Xm8XVy/OahA/sFN4PCvjHuWAd2
vHwTMp/6PWboOklAIM2VK4rCSpgIP2kcKk/cOqoaKkFfq5e6ZsazH9ivKNLv0MSs
`protect END_PROTECTED
