`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRh1OaF+B4v2Q3QO/rHLSxiJ+c/W0TrOn/RwCmzOK/bBR1lg9KULqhuHkIFJqfkG
XPCgivHcCxQGrQj2RlgU6yIUvrOd4fBsDQr4/HcONMu88ergcWSqueIui9wtSut/
kJ2fxcFIf0rzIxHjpgNBdZQI6kWx2KKB3OOKUeYyI8pYbFHFpOr1+jR0T5LNgqcP
QhbA9FQaKu9VhoANEQdv4pLNFx1hhael+i1/McfkYcfKxKSeCtaLmoEDbFtKz0ak
sGcmz92WBMkBXJxyq+UTXuqDV2RQ9EQwCFqZ9e2I+IPH6heqFZ7UZq3SRghDLGvr
fLVjvQDdonoH+r8u8SV75d5/2pYiHfRspRPN9VHVIM3Wpay5nduqZO4ZKpedqyo8
Z67F9kEj6bHRTqJLCnzqpIOl/N2cc1S4RQ7ZOYvsfP96oZSeJEUOITIpDhVP1r3p
TWEBbdmm9ajkE5/oMdxbpFLtUCWOpZhvR3YcOTw+NbwaN07ZLuhSuU6CcExeyFYq
C76X3MidRHwGgSNTfW+uJRI2IspJAJL3Gi4K6wzQrN8l1a7PYimxSuc9Q4FogYeo
745jR4je86ghWvOrlw5rj5YTVI4JRAvbRsr0uYFMKl5njbDimrwffPwlBSP7BZY+
Z7sqzi4xzIZwKmmys4OPQjNelNBsPiWapNLLRP76qeTR4pf0Fw6opP0lcOeVD3m9
LiilwmMRc4EsP4rLd3KXHNIGhDXSGX/mkRlAkIvRoOkcNiBKE4Gl92K2F7rhuVxj
uhKBQ5FZ0lAu/QP8VGDeWe9BlBO2D0Jg/WtMAtY2oC+sLSZMPr8ZTDuXSUMNYVqY
MRCDcruQ09JdgPkyMD+r0WU7BbOciwRS9LkQvsSIpBE5rcJrJu97Yl1K/cq6wDyr
kBvPSpdtdglPrDyhGMLq4UVWEeNT/Thmey6kiXWKbqVe8g2uuBzgSV2rjwKeboFy
HxsIzoqA2b/NygoWZDEY5Apu+2DwYgHQ3JD4DTCnxl7kTDKLE/VdET7R4WMcYb5Q
DVLHvmpJcYQ0NgXF73uklE5nG7ezjnu4bWH/QJ7lRl7ZZeE8pOdYx1z1AQG5bdJ2
7TSs+nWG+a/+/A/aN6+Bp2iMz1w7UbZG/VYoZ/pLZEDFWZU3S7t1LiLXLWAHLO1F
Nc3S4MIb0TdWXoQ66j/spItGDa4HgfIG+wCocD3lW7Zm/vcLMSYJ1imnw/FIEO2f
tV9xKwIOhlhDtSr8LHmkVRT8KEuD1EaQfUhn2Px5v98SDIxrM/Y1GrcSistMi3Gm
sJsB96xG9X6dpS7txCTM/FW2B7riJEZdtCtZJkKQofvMGvduOVEW0sY+o17+BAaZ
qwvWYc9CQkgW5ayrPa2BekEDJTUgQ8Ho7zqI1a0a+BS4jKL3FndH1lu8sMDKkvR8
Yc3c0fd/ZC69jId2bfWDZIMa6UdPzmE5we2ON+is+AVyqibyipFJJzQWSEMrVceB
mqvOicWbyXo8TfCK2ZM7qRIYDEjQZz08aRaKzUjzw/LtgJgNtdtOlLSA2MWWu8k9
KWPnW4o/T4dvfzoPp0Fs7t07AVp4xDF80XRLYJWYydRDuSakpCOuQ9lIflQ1+CiU
Ep+fEfe863aDrAVhrNqaUHBziX7499UfLAs+DOw+YEkkUMkJyANDGkNNElIGz4JC
WkQ3xr1sqn3X27wYoBMUSuWXzP/SWudJTnQ5sdr2jDjj2QSZz/+iv5PukYbHfYWW
qlb0sLDkHbDT5DTf9T05wMlSRzFdfjdtUZGdsEpK+7bTSd1i8BYUrKvaSWNeyzqR
ny3RcSag5wBxV/TCZDm98fUoEon1OKGCARtGNCXsFOwvGABZiytPzBlZSIbC2KiF
WAIt30SEcLDIakIXTpiTvdez5lnFrweWjBjAXCcST6uT80qwtRNhsvv1c46zgiUv
Y2yxDTarRRRptlwx8T3Mnn7G7r1faWGAsS/V0yYBOqTPGeEQ1iCLMOi9LxQO6Mw8
JpAdOhYGmzCmH0c1cn6NI4P/pS9J/8PhjzKwkVpvTaUJDt4dT3cy2zlLn+cgHctu
F4GadwGV1t1WAABQ7dcqSJRSHZbWoe2IZ0BDFSKvU+GH4JkNpLwVDz7diS4Butwp
PYpPXhai6w2pBqG8GxQe3GT1yxm8g/1k02ode+JhdtuhFDTQjN78I84xfQQzNKQj
mjwM1ngkJhUM4KnU9jNOCDsHlboeRerGHwyYmr7SbHpWApHdIhtDmGjPqvicJ30e
d/drU9il9yymLvH6nTmAojgz7PCY0fBvPb56wSbboF2G7BFyzqUNapU4kX9xy0i5
eFmsyMje2vWmZX8xz9rTlMp2sDtz4z7aqrFtd+/vf4RSIS9fzzTfeWXgMeZLyeZe
T5Yj20W3WErt6EYUbsiXIKLB0Z7Tw/nHMKtlf4NqaHeZUSF/i0SNCdF0r5MfPy/m
xRsfILwMHT6oci86mqH96zuV5IcwvSbD6agHVHsQtEH6w1aonErPQgw2HAh01raq
rP1t3jL1rdE9+LSLMJr8HC8G3AeZII1E8VSKRQ8oP1NAm+5keYoQQe2Gyr0ZmK/z
6CdbOwkLR3NyejPedsTDDy8izqt0U/hpkjIWQx2LDof65DFsSTYIBwAvTVlP7RKe
7iyebCqDSPh3b820rTbxcZ8091yhJJXXoqeskVMs7O0MB056jABlsXzwkTAnHCnI
NG9RBqiYZADGEiVDLNSzqIYcgJfZr6q54H1z/PWBQyGNnQxHIRT5JWOz6KFeCDSj
5JBTMIqQ62JR46yLBXk74CgJa6wmPoYL4zYvt8iE3A65e52ccR87JNp/xguJ+ENw
/VTrvPJyJIMP2VqYzgNyt/oFyg3HqgrMGt0tLHGvHUXIjqk38v2j3uDvWMQJnuVH
a7AyoAPUx88UrTErlO4PoI+v19Yh7fyj45oY++3VcwkoUX+ITdkpzkPFStoLLRT3
p66V7dbT6HJsPH2/Mw/JjTGdJ/S2WKWihRS1/6JeDywFqHFRuZDCfoIPTCrYRCKK
Z/jEPYRFWbFa9/S2G0j0+egpGY0RjAVtng0vuLhmkw22rnHvd5dLGcRenoEZSeAg
+Yc5zIgZrP0YCwlY+szx5hjbwDlTCRxKXg0SKi2XoDjiv8WEnCiRmsReZBSkngGc
WN6ik146QZl59f5tzvM1DIhp33sAc8iXQPebb4iGnyHHi0SuKvkqQ00DbIiPBHxA
M+aCOecg6FP5LoIcBGxa1sN9dcE2xm+lDYIRX0qgE5uLOKluDATlmWD40Fnna+6X
iGedjGQyobSJAymqsadbo4usq0oiUeqwAhnBlUIJhOEiYkfQ2gnijMZYFNZH2Q7u
2fmtuv6StI/tWd9PLRiERUJY30K3sbwfupsEQBvGdjIPb2fenbfKrKStbuBSMgpf
LfVwD3zz9zQfLiFYLVHx73wNk+3MvvJ3zqZrSQ8daf0dm6TuVFqxqPYPIxfFxWpX
7bshEyqmYpVZqbdkxL2MJMIgehfwt3fk+8LXBpF0tntf8EbS4aZK6cqjPORqju6h
tBbRU9d4WPKwsr8vSsgfcUnCf40geQzjxkKqPfcezu1MXRc0kgHWkVv8VrY9Rck7
5rtNZJJ12KsmJmDXs8FtPoB67LjDPTyE8nSVER3W/+Ae9MwCkBuGvkiQsFTw0YIc
Vzb5F0wEUVseDeuruFqsBwA5l3tiTJcRa7DbTGDD8YwHxDnreYhj3sLg2TjQ2Q5e
+t2EVeR45BK89tGtP9g3p9h9ZMueuJYQZukEH1JI2aGJNTmhfdiJMXnmWVoT64qo
VtGvARSNCt95+HHa5VWJWClHsSBfCjEfANo0qbiwueSR8tY4QeL7cOLwt+Jc2W17
Gd68IAdTLv+lrGC45MXsaNExoyxgtEDU08IT7dBtJGQa+eb8ACXScweHReZ0dQWn
THf0WTfCUyaOgGyC/TQ7feIihW6rrGTg6LwgcY7SIsmEKn6BIC/O5YxuokjuML/q
vvHSkz/8460GaDSZq5bKZxA3r6hLci9y54NB0b7vwlkOSTxy4b0rU5It7Pw70KyI
vD1HhB4kPxfNSmHig4hG4oeMMgBa8jNuJElMhqr+iNI3Fo/3u23bTZMPN3ewEfjM
2F5omVXigEASxYPcmbeAuk9/ai4IHhsX24aqJHBx3xg22Z+9Gzj0wtS7QD1+GX/W
O1g6WIJcYyMo7OieEGJ6wDVPrVhzyJRcYlRKZROn7IB6BoaWdhA7oW0BvPmu1kwy
faGCBxAoM4evXdtUsPWY+UUuJp+koU4XoVzGSF5wcvGcyKnUJ0ov/KRFeHP7AC4C
QQkS7Nrr4ZNQh2iO7g/p3BR/zkh0+adss+huGljt1n/1MZTx42bRk4qbOGBpNC4e
v3T81BxEAO017tAtLxS67srn7ceog5bPw9hQIMpU139qtiKVWvjyDhMRnNBnQGlW
CAYGu7bjNg5/gfbCJIads/Dcx/1JfCSU4gpykbO0erb31LYiqEf5Mr4gATb/gnHK
ZqvN1KMZLvuexHV7RtKdjF5KbzeRrL4s+dMB8FHLH2+brxaodgmVBbawt+cMu+we
bR2V4zsyeanh/s3krrlXCrDRys7WjEkyOEfPUqAhSWxNoWtft8sh59qC2yV98csW
3bzgyhbroVl2nmyTGcjc0ec9GeLzqzuBqq9GPxG9Ykjj/J7P+xTnyOLqrI3hTwZj
sX99R1HtxwVwO1sfzg2gvF8kq0/tJBsFZDigkEJymR2CJxf30//ZF85uzicA6yup
iHnge/ujOBfpxJQo59OkVD+OsMmJk5Rdhrfp4GLR7y2Cshpmpo8Z08dT+yiD+tG2
bg3xjy94KuVlGbGFUeB1VgdyNzyJFGHDRTd4BysnYmHiVWyZTQDva6pgBHcqE8nP
j2VNE/KRx7tISBScP1uagFZ5r7FBQB5fQ5QJWGm5wwr49PX8WjaxH/MJTsIwA7hL
YdEK52Jw3kIy51FNZVD75qJeMtMhBphjDRp3LKyq9upKKLJNZtID0SrvXw1oaAUK
2ofuvdZiYrKh6J+V84SVJO14+3JHBtlKkwPyP2KhaWf3R6DrhXKZwRSHw2BMxuhT
MQb1DtIyV0KNXc+xG1Q3fXOa7cideXCAz3RdfNqSs/FT0KbdywSHsuVpjXQRWqf5
+09tDZnSQ8N48K3gtgSUq3JGylNE7EIYLgfEJKqacgqLMxh75IktxAp2We0gvt5n
eJHDYJkt5MNlr9AkniEdzyBcVvLGbxFHvhmdZsCSaRNxwyoTaWA1+lFaAX0VQF8z
1LhqioAwvbEc1AQkZLkgxYqnFtvGGdMPAgaDSvNRA8TTdc2C7g+hQ+SB5k8O+2qV
b0DuYLz/GfLmV67HjtIx+RGZzM+Yh8gAnh11Qka8xUe/zDnG9uMVoPFNp9j1oIoV
JsCpWxo7JNzgVb8+XNgu6KiPDm+RIx3yIgy+jgaucmBMV3QFixFZvohiWcbfns3h
mi4Gl3K+tk7bmdJ1eAGcKYALa+N7xemBbNRReKWfh1VVPb5CotQ1GKwlhMjxXQZw
HFDRWu1puEEr5wc4e8ZTs6EtVvMKnfjWjIYP1WArwha6IHHkE0WM4miWnUG+FoMB
Y4FzbwwO6/h8hovaBYBvc/6m4V5QXWFoPWM98wDzH0ei5ITkHzOUK3knkddy6Zza
LFjSbVLMB7XCTCddhkm/4ezn7lNcjT5LreEjBYaQbK2zgvYlSE2+C8egLoIHslR+
5lWjn6vcSvY+08zVcYtww/8eTzpzSmg3kDTDB+RqRQSdjp8z40jD/rdSOU91UVPL
r4wEHlvqk+gb1WBtsghwB8uNkTCWHnmeHMHGu8P1wYWOLfcJoQ3t7KIMPHe2XORE
d/c3qr0YXLP3XGiNmfr8v3kSxKZBai0zksWIzSi5h9hZvKHzulmLQGK2jgQWG1MH
sVcahUfpatlVVpwcmQ+DiCcyb6Wd+giQqwAp5kMcngHdGkQBLNGtQOy525gDBhHr
hdCOkhkC+5LTd6+Qpa56yExD+k1pnKhtlrvFzv4mRUDEfaTRoWNOgbHS21ms1XF1
VFah/lG9n/VrKPh3xDUZmhTFUKnNKc3mbHGP/JsdLYpjNXv5nCsLesEEg6nI79fW
LZzyCblfxO9VmIV5qdLPUYkSzI/zrvTyL1+MRnNt+BNlLUFbek6JKa2P/2LrkSAH
1lNzbK8FyICLL2G9SwoGlcARl0xPcsCiv5eKk0kRh67N4/Ys309PT6YgZKPbPA1a
Cu5Vry0Qzc+cj2lRkYnCvE4Ye8MsulbuK8Qg9g3z97HHxXDRjosGD5NeRST3Q3dm
DOBnUiVNpy+ZEVwR2rsl9/OHBj2A5VRlzPN2mta/giUbm+9o+uBg2TnYjHQU8EYg
CbX0QX4fp0eZOo0qJZqyUHNiwmy2b9We0m9GJQuWsy2jD3xEAaDXAUFquoDiIh2M
+turGq9LLrvHwY7wWkglgM4s7JhiBrEe6bk3fT0+HEUvMl7WJhcnYSHSPM4mjvA2
OOLcvWuOhZ5M9hJk2sO82mEz4cwYwxJCaQAWer7ITI3n3TlXndwGSuJ/E+T9AM5D
uQ52369/Ls4Lodn1MLSw8Pgel6zVB38PH63IeRlJl4gzImzYNcNwsYLRUIVLyji6
oIlSWHIMQjVgoJnC13vanK2ErARxk6gpuk7MCybIWRcD5vIu+lxHCDc2V+v0HU0b
cYV2PVXRUyc5v+/W4w5UasNy9UlEXv2ovGJz6s7pO2L0tk8QS1NGi2BFxP3zbdOo
+yDaEm2YplBOndYqZ/IOTxGN9XcZ6cSr8/5w5qCLE60nhEJIze8aNlwZm3CBfprk
jr4792EsXn5rjbfy17qs3SbI1O1h1kyGwadtafXyI675P6RRh7onx/Vem2oG3F7h
DoUSJ2Exm00tKvYX5BJMMGvy3yov71og9GBw/TPrCfdbczh1aRq7y3ykp5Ox3wub
MT8TclwhD8gCva2q2A78LNdjM3hAZSWiMSNEpaRaRbylsZB9R16b8TPAua+4C/S9
jeYKL/smye56Hm+96ZiAWaNNnzVG8lGxE0r41tNEwIxEcv/zWGv81byij/zM+LIF
zj3zeFs11cCYeJbIjyRpDLq7BkavHFT4WfUH7s/X0N19YBazJAztz2zqYIavyniB
NcwORyzG9Q2vL2U10IvSOZ9dz1tUs5a3W7+TUGLLlil9kwPsFoXhZdbyMrHqizMo
mbb5Ulq7K4aYgYlQ+eI5TQGx2PoNygDJaXkk4Dvv0p4OR7JldvZj+l9cJpaACF5m
//A5o+++1n1luVH/5+wvtx3uPehDkvL4aIs5czg55czC29i491KryGIld29QvQcX
f7wWIR6kxyCXoMdV52jKvA6WDe2vkEFIegEYkfpDuJvzuVCy5yhw8a4ELA+TeW/Y
wFFCTG4c57WHROLGeg2lZeU++vyk+BVPds9TbIO8qSePIgDrq36dY5TByCGJ8EWA
9r4X91QK3ene+XIuVz2hY644EDFEsFz7S6q+8BJfTXwBlDmL7bbHHXl29E5ADcRL
tMCVIgY1apTQg71HfjkUw2UUgCvZO6kMKDZWJKq2uO3hAID8a7fGIv/1ltF5aFTb
uVJF0+loNQEpT4KeYkug9T/dJt1z9A9YGjAnX66wBUwoWJqo1s8Lx4pJLfKEJiW8
xtv9k5RDwRKWnePmZw49V4VVLe11f/jGwDmQmYHMovgAWJoDkExkwe/Gq6Sy8TnB
cJguoHX9pQSslqY4mLMei5z8bZQPhiGhDhvRSkFeiHQnFYm4ygtGHUUTSG/fnVWj
rItce8YRWm19UwhQMw0eEjukmaQ4MXusHqyUI9O0N69kM9XREWjwpp0tjrZ7PfCE
2cp8LM6v2NnQYOQs4s6GAKNEye3VFlEGSdbhdqad1wSMrdyA001kX3a2bHv5RSv6
8BXj7K19wl0V26jAIUbfPJx0+eYExnAM54v7Cn8poX2IUks3ZC4uOXEaodZ6rvYG
HL6PJeY/20YO6P3MF30pOcYJD5dbEkm6LeCZYfZf51ENRREsIQaMLyMUzWmxGq0x
vFt8G8kh2jLBr3DFdZuvTyIgo37b0ZvCg+BTNAUSFzVhGoqOJQFt7zxZS+PmE1oC
qqMKRy2pqiHlSvZjwNhYRA5w/JmEYzGTPwXtPr+qcwJI2CUeiSyCPtST+LoAN7av
7SKy7N2UFQPJIJWrTMbjpESHKdsunHTl0hawPq6G/zT6j/YgfyBb1kh6+IA/RB9P
S+7G3kYgP3avSZE1yJyIVvflzzWcGevR/h+1Nj1FRkqk3giGPhnESCA5XGjjfnsM
F4ixkmvrbW7+YOA/rC9WD617oCaVRqY4sEMUSRfINdPC7F78+lA+C6fktQReyN8S
KIN/FIAIffqSTkTFMmhiOrKqIkia7jpEZxuvzJSOthU=
`protect END_PROTECTED
