`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAjFsU86ki9DHtO+bWLmOAYaGdbGF2cM/xeJzYfzpaVi86aIZL2cTTHm82kfEn4z
cCquSop+KSV+lBXbbzXd7vtiySEUxj6j6e2klzw/bUuyfURXn6LOBHj3p3BX7axQ
xEarhzthHx2QOGK98nMYQ0Jy05thOym6p4gyLvWcAvlZQxEoU7FIiuyWUV9GSDL8
NFRQWA77IfJ/iuc+8BhKQR4wNKapYC1M83+6FkiBUNQcKhDiO8AsCKpzSE0TRIO2
b7XOSiTrD8TtExO54W3TcIIHY8vfN6icXR2oi/rCJR4TuUIifh/RPaAsNtp0OJNc
KIVRN2Vf+z6eT57U0XqWWDqyh5dsfs4s9GDsTzW447SxxZiEHJ8iqz9Ma6fvObIW
5qK9v3wiAyFdadCTVmh8AsPl1LiEXiKgLO5YT/BaK0PMaIF72EOVf6rffauUCtxk
oAzK+vozLPSO+tlC2ShDntC5CjkEY+RtYt5/XrY4C0P/Xl4iRdS3fJp/NSJMssF7
akAhT7kUzIoKaKnJJXKF4XpOJpdUcU2N4U7P3TgzOPdFj8PJg0HfklVG9v1SqlBQ
ZBcUajqyplq6vcy39SWAmcDCsfyu4I0haAgM7auZgq3+iFMnAWWlwAschd2FFK2R
ldo5aSg5yXunwUgNAzKpX45HO/5kxwaepTR2T1hG1o9pEodm/UBf/iexEkluc+yx
l9DUbncvrDWPdAfqmjPg2sZh5/HghWNezBnCg/uQc62yrdt448hWrNeazGbZLHlc
HIM0CRL4F5JghROdIL1NM78Tf8prUBMRjDWTXcA3gL1Izbxom7x2E90dBseenc6B
fTxw5f+56Y4gLWfbMCioMftmBJSMJ75rQw16XoLTp6LYdsskuHh6bKSTDpZqXJIm
zTrB/J99dS865tDvRJMehHIQz7M4t4q+B2+gv4y+S0mUwzl4Qs3ofzzBijljKIYB
prhwuz6N3UImSbcL9JnTxS4Wvc9L3UGembWXxGTz8c8fXd36WCAi1/IzRiiV80/n
JzhNS7TEv3afB1T9qKrkYWPLyDZrZyni553QQhM7d3YWgJzFP5T9vdLEa00Sj0Zd
8Buyg1uKLdRHv2+qvwI0VLwPxEc4a8wfLEOxdB4OD/TroEivd+C/GwW9OhbhzZIo
p773KM/tPTSDlvmKAaaDCykECWGlAA/LUbJMRcwhLEXMo6cNw73hFgXo71CnP0it
8sG4/mvhxAOYKl+i9lEsj02/tDsIvyD+9L3v12lpcA1LkU/PzyyKmqQw6glNHs0I
gaJ342Q+2HDEehLT4T/oxU45WMLXd7MCo7eSngYJojkFW8MrGC+tOxfRZvvu3asr
AR2HayZTSyCtinlIrGHh5nYC9bEUkMgpZl9WjcASoKGjpPlU1tNAPip0fXVglmVo
SyZfhTLZQT/FNkN2Ii8BlQMaE3fuXNkXIY4w1v6G4sxQKM8u5vwsa4ALF0Z3Q6Ej
6U5HulI7r6+tUOIXZVH6YebJhpmAIQkNkuhmB+ZuvvOLQf8594dKbKbCn2pJL50W
L0IqPv5IiD22s7/V+4Ax/3TNLE1RPqWKVrQWMWxQJv9ANfJc3Dv+4navq54TG+Cx
ngHJAzm8bWRdVFRf+YU8/tSJp+asbrgML1+QSydrKuVWg8MAjqJIBsToi0gb71L3
JEEuYTe6tt2K9KkV4mjLjYz85Ip9dzcW08BLt/cvUJGFrU3uBoWBHJsDbyysN5na
5AW1QehhUtdNYtk+VbQLtOo/f+Hn9ry0oTPILTej0mojss/NXTmkQOUzuGXpT3QS
RoWOawd/aFChGm3g4Xamjxp/zKkpF0gsUvIxrAkZKVPA8/WysArnVQmxCtW3tiW+
F9c7CDzjuGmL6yxneQhmeq3O/poz4pyHm2a4ehNXs1VVVn+9J0nnsb7zItqELKuu
hUiNBMUxBbib1Ksw0m3bQh+ZXqq6mUta8kpBz6eP501U/CT8ZCfWyA1Yv/DJlZkV
Kw/PX1CyZG+lNRUyOcYsDxzB/V/1OkpBFZKgb+D9v5ur+mbBjmcZKTSauzQ1O+vh
44Sd5bHIMk+Wq/lpuNz+y2HhZdkFcnc9WtVnQ9GC6ig7r15oTcUQNXjErGTg0Woa
ULmsdM9TIB0DeIIZdmrj5qzZCTaDKDEWAQ9mW4Nmaaep85S4go4WKKWH8hKCPBPZ
rr9LwNKFezuePj6fJgHuMDsH32uogmDDJ/pIRhyKk268Gxi2/7wXJinrvgLe0Fyn
9ZcURAWSaLM6GUGBg9MKNqal6tp+9E17HDJ2R9mxe2uNjiUvXF8+poe1Whx7yksU
pKbYQXxKjuih7fqZpCUlaXmOtaJ6aZ/DNKFLBQSk+5ARrNZOPo7UXIF6P60fSX8f
XD6L5ZOIdyDyG7CRjinUUBy/5N+p4pyWAVRcRp31sSzutSYbk23QbDGMRFh5dBen
PjVklzRqY00w3zVxYs7R8sTQ0eALEWSVIFL0dnqF/KW2lHdktpSVxE7k4IcZLbFa
keEUAPB0qTvxX31JA541tybnyGPkrEzNy4fDWeBy2EOmuH0fI7+CLswgRowLhVbO
5SOcmBoTH/acWm8fAK6PC9kYgcO0VRSqpnBwK6c2mK5zHT/DpBeRLhm0AhxZpKlA
9Bgd5luN61DRHtAnefffHBLUf7AVqpZKJeUc1HaA1/MUPrmU5up3GF5+eRQwi/SX
TK8rAqj2xTSv8rDgeQu4/Svsny68r7v8ywtDb5ORTbW6GmgdbdI6VXAC1D4ReRfH
7mz1gNL9uR7m8vuLcmHye6cK1oaDhJb5qqGHf8nMWjFhu/fioMQQlh22dW6XOlQJ
GfnBMMmqHl1xGFLQscyxZvc1zDGK1EvOhNii22FsrEL828xCjJBEQZ/IhvKNVPaa
sPMePrAVoS73fsr9Vr4P36EAnuCrznBJkb5iwpnX7WHOp9JUqCVquUDOCfBPQ79y
pnipO/O5CMgqztnXbXyohVfw7OF0EVUk/E1YDQqkkeu5LrObAtV+2FUOFeeuwp+o
PpgQnLUS8vULzbMyZ78Vc1Ey5RwlUCkE25MUShTG1RHoHzqw1A1+3+JLSnngzq47
RXxkBHCTA2n0ziIp7vvKnLrlqyVBzwR3d7H7yyfa62yoe+tB9oBOqrhVcVSY9qvC
nXdUGlwpyBzf8fVcAgdSJL2/jLKkKIkvwF/mkJaF9zrIMLOIjljvcu8huYsoaRRv
MT18/IIls4bZzPNMJQvSip7Ih1utJWO5I9wRcvuohAGjGI9H26aFPZgejP/dZlJ4
yjPWa0O+1MHJtDllNQx+MA9KmgkxKkrNm9nd5Sl0T9f+ucuUo5glHEJcl1JRmGUW
TX+eaZ7PrvPH1/uxneveFoZVjBAguNnBv47AjCOzoXRLcBdHxdZ8D+W/vfKOwqdC
7t56cOvhf6Fj6PFiUMrRCTL2pFaRiM4WpCBktxYdiJ/41Q9V+Q0MOVrzijyLMVRc
uFWGJopWZrYpQy2NT0CUej9IZimqleWe4sqqiQAqHN9of6TyRL0Z9fNOCvnm7Pf1
UGd7uZSrFLW8r1MQAAi3HhEfHcZ1dMmQmbjuIF5Au4QWfHOVMHziI+Jwis2pF4I8
KcyCSbfXNB/7cNyK/lgM85nCHxn1WZBIOJEzWYOC7w+gZOMOB+Qv+dBqi1oaOwsq
OgJEMtKPCdKWkD66vbo6AWa2nwq3JMAbnXVajEOdq/dzifqD2UQroAU/Ok0u4afm
GtHR/RbTzWZs1vwFSv4YoXESsMHCcTnEgl1rvQphl0d2SuQR2g8ji0FTDq3yPLBt
rkLT94zOOQoRkxnDG4UuMnCLH3wnFu/9l5AGhpHMNemkQWn67T8XHlk7FPmBJj5h
uIPDMPO1Ea8eJlvEf4kMW+yLcNepb2Zevb1dT7JAo1PI1a8LLxUwTxdG9PhFlZ3L
cOrycFHksL5K30BBy5dn3dMGnZjx5GkdNZN3EqqvE4CodUfSy/bPXLGCL7TFnrw3
dpn/T9TREnAYvK8r6JNca+qmlSd3AeNkAWBW0glsnKrBdTO3ThlscH3gVlRyQ5kp
xUA07A3bg0f97owCr3k5wvDklCmnDs2ypIjG/NSQNHa1tHYR0jpY0cIReHgDQ8Rf
xp7Hb3sZTPhhUTlwe1RjWsLevw8bTaK3DuYyf8jXCax3TF9b5ZCPEpu4hIKR8Y6a
KzpC7MvhcRD5oDO4EKd7RKU6bTvJv7mAp6K3/j9DyQLb6mIreexyfF/4LyIaDl0X
L+EEl3Z0xl+yZZX7OQ9asoRo8nZ1XEwWea3olt/KIo3FBu8YQX91OfGpk2BrVj75
iCMoVBzOyWLK6PM4sVJRublb/nz68ic/DZ+yxrvZo0B12CdAL4y8/GUOTPx/PbwT
bVKEAJoVHQmmEEZ7yRTIfu07JAY9x6MaRV7qmReF2pblBpbC1/oUaquyFvdiazaf
pBFlWdnJbiZ7E1ZqSo68OPgOLW9m+QVWP/86zuu+XeZ0PzbxZFDXdYzNDul/ufN7
FiOInGnbeZ13tCd2nj/pQD6nmpL9oqloWLQZYPbxZYkTRjF71fKLqoHgdq1ZLSWm
RlWqEtczllt0Kv3dZsv8iPrhhlJ/uGY6h61SApCYoJG2otMSp1bo7ny+A0czC6IS
drDuaS1F7ln7s/k0oJa53EvkeL3IUbZiIvm1y5LuvDee3+dz+R0liwYBazbmkRwt
ry7Z8HNlp2s/yVBxdhhYlBDO/8wdvHf5/HRUmD4WLViXwFuNc4Z1fC2JJ9QZ/Uof
XRRu/74cZ8FG37scmWA8BN5gwly01JskNRhwLKYXjZxPeGqNefoasTOC8kPg1Q0G
JYLv5ru2vLbm60ueSaMVKKQtaxvTOLHvM0pQZF7SSgXIHGyOe2Q+aRJ64jb2Q7ZA
yxL+hGRPlcRw9yNUFgM39pQ+RokD0FyCDbOszu/CGIppFLcJm79dOR2zfHpida4u
A6reyBB6u7+j7PHzf7/xMNDHN3gBVlcnOVyx2TZCzlJJN+AdHd5nE0LKhWoCnzd8
/X40dtA99FwBuNC9jy6DHa/YWR6iAJLk4gqh5e3UO4WYfZdOS0/hCZbM93U8AW6E
TECwSgrTb/t5xZO+w7YZ95BBtlnM+FAYVRsNGOJw3Gs6I40chbSY82R3t6FZr4EG
GIKibQTVWAosZGm69d48hXpunorrJqL+y0TW2Kk9ESi6u81T2d2dSCC4REUDkPSi
8TZDO8IlzYMiZ6yTboLXFtjVvacmYQRNRv/AdMZhPu/mKmO0IqEOq7LpCJCYZyVm
GRXZuAikGPxkZ2x8hg6jJgtBvLePK7gXS/LOWQuWlbrqXNPwBZ1aQSrGfNToziPf
7lvIsn2zbCInST3z6zBYFPf2aUqxXk6dtnGkcBLnxe4SQQ1dElJtyw8/FFfWRE1K
+o7jWBGtsGp0IXiR4IcmAfYUfL/cs0VNYALZH0r+nxChcX/FgUASPzFpj0zzJCCe
sU3C2AHcgin0VXPsKHwCRM6IiOyMb3nlW0hpt5s1yhps8ki67PNRQ45Pukk44KN4
bzCFo9VuORc7A5+Y98kpTs+LshDlzbz13l0Upw+CybdDoboe08Bv7P4XEd1Ub+pP
EMej0HyYC6HxCqeY8eNFeHTg77F3C7iUYSWm5yrRxQUZHV2nuhHK39KXRZ45a3cq
YOZ7D8nbGjgxhazJHWgwjMfi38yPJV83OuYP1kXYF+pIdOajY8t2CSlW9F1QCZNv
qlDAL9iy7Amp2EFAOwrX2k158z3CqrFA6mR0BcR13NVe2eBu66a6cmTmYk6nn4eC
lsyLIBlXT1SnnMWVFJRzQN1djAtdde24PSihZDbBdXrVIXTIXSJy4tuLsJsUQDp+
WPH9c+dbctH8T3yGGL90WaRP/ZmAbF9p+YyKsY6/UWlCzHZrTje8isIz0j5uFaL0
nx7pO/KSk+XvrmgDaG8nVGb6i/CPGxpa4wnjqMNZHJWh3Lk3b3uwiKN7m+tpsuTk
AZ2Uh1l83+rvCLw5opYLjhyvb3jAhBqmkYyQ8LEXOmfSk9tXjPlKYeVru3CCYuR0
7DnNPH+sPATE1t4xlyAagfWONR+jLvsefSW98yQ1NnXeZyB1AdS/0yLTN979h01Q
hu4rKAEpcTjMv+zOB8XyQQS+22EeVo3S9M5Y5OqK7pVCwfGjfVEb1AHIaa/rv2eT
yKl4h/gfx7t7yrKTptZnhsjnGqxef6mjI5H+FYi0NKTCorQyrq4WMfrbPffbRSBy
o2qjVY4UkL5jUk6nePE2bmQP8HZ4rVJ71/2qJH8IYNXAGJBX+1bkBE4ZGobV20w+
x4wICpmKL0lBSR/lyvxeSRQXO2oZsaHAl1hqLCRDPWIG9F4fPTALeCXjgSfJlxiQ
vgPUlOEy9pDah1oufyPrp/N2l6RCew7tje/vLNSS+Cso9F6bcrg1wplX5ez72+TG
Ipk6ViZRAuhkehYmQlccP14DWoQUjtaybYULeEp2tw/Yh68/Mc9zJsyeMu9PYaRG
kr2FunDLw5it97eq5a/YDVIyODjLei3O74F8FrhAfQLXnCkXhp7dRg2jYEt2Gl9Q
K+3ep/vYYCxcSP116Wo4vyrjDXdaOl9U6zXsYEh+nIB6MSTtEaJVh6DLa4FD4geb
vIrnBd5y4RxD8WBxSMzo35tC7OEtxQYjfGrOiSb8xScF0NZtI80oTvs/owfZHotI
CJsSah9Q2G0WGAY+WSLw5XvR6QaqRV0z/FpWQzHB6/BmdicmweOv9Syg7UdCVSdj
TY4d4Mz6mPDBjNTOgCQbtKQHGCO6bzJgcERxUyUFjzP6KNWpkMhWp5PqFj8U4BzB
PR0NY2/Q4Gjy9U//YrttG43OkIcZgeYYt/K/EC4hYPm5r4OosaAXGpUlhRYputBe
B/tRWv9YD4wVKJW3GUyeUJn4ME0okc6k70NKioaS1mezL2FS8zL4IrTr2O5XOIQz
bHsGTj1lk3ThYHfiHGfoXzl4l7eJqsEBRED4DRXN9M31xsBa4bST41PpX1nofaR4
+BM5y4DYusoiV97Ch3bL6Zom3/ipAw2xIKe1CRuoEG0SxqUZ/evAHBGTUIVJNRZk
Z8Hk18RFHAXoa6cpJ/VU3Y2aFJlNg7l/tr20g2PRisRDfSkGhTLqdbKaw2ho3RNr
G/Mf0hb5JvZw7UbXUI4DQ305JlgVqXaSFEjD2z3Wo4ikgCZ7IgSaSRHcg8NTSlxd
910XGUDC3NHB3gs1NQbaqvFz01tHKep81GigQbQ6xYJrm3QpkqZMKYXvjAOHGCHQ
rgNeMwTurSPjsVM/1K2z6sMgQPfq7/v/bIy8pFyF9/tpESn3vIQqLrU9lN9yfUxY
NY7dfIWhO0cCGgSseQrX9TivFuE4mAYq8XS7Uq5MApgS5VK3c5vFDl5vUlje21kf
COCQcanVcEZNWN/kBnghgAnGhiPY2Vs6b1dId7RycWckaVmr5LB9KZzhMNWsanXn
EWx7AopL09mDQFy0AxAYduY79XfuCZKc6v/m/BCi+2sXYmBaw+yicO67lfpGboBv
/nV+N67V6bp+ADXvV7vtRoFj8cRgpr4RUL4vBWnZWURH6/IyGp/q6sKy8L6J7ETM
PmlrfsH0Pumhx0V2hlvhAtrGNf2W9HUn41nUEOsBfXnxt2nZEgX+kAsH7Ms9si/S
w5LaGumP52mcHvKiOU0ms7wJQFhiIhaeTFQ0Jxiv0wdpeqFC4xje64WBzjoScIj6
klLdUPS6iFTzDUu2JyMFngW4h+EDb3CG9bDnwRBxTIwP3VhcSBCHUqd15S6qU2qh
rEtVV8c7rQuJNj1U6HcItHqnjqpmQozrKjDUHfRKx+kwR77KIb/zFELf4u5HO0wO
ffxbEeHITihDX2eLgMNAIGo79168ullEMnzOx69tmJJrz/DEitskXN2Bc7AozOGQ
6fP1+zccs/K5oHk4tDlMV7i9NXUdHcGwVB4ri0kTIQoOzkazdSSLW9Vxbf70GqXm
oeKMsr7ZZXm2wgeEuUm25/g+b6UToNvx7/IAU5bOc7xFLq/d//vUeb/HtTvEgjMF
430MhCu7FDiOLKIV93mAuP5S3TE+ZGEy0eOj+/cbmOnc+7W7zZ/w8/1isv8K/Xo8
xA7MF7HtGsB+0Gvw7/mrm0Uc00WIN/n0nmUiMjRPH4vFw7qWXlPfnTPsqFCsoVuQ
BoGu/HSnrjAuGiTGoSYho2CJ4L8dOvXQuAstIsrbT18Jn7c6u1m94rmOzNlXwBx+
4HzYmjIlCL2mXrKNcbiOB+n9RsPeek9jl4jkXXvK5Dfu606tDyu19RMp4Poa0RaO
FWPGvwZlLpYFyMCPsHzjzheUk1n+Hlso2ScQChpQfC7GENuBuVCIz/dr1UpyD9+m
rrEBZ3VPDD5eX6yeWPeJxdx3lS4Pmn9pNmP+RAjtvz13ujWGowG4amzSA0MqMuYi
EsLjd2Mx8zA1ZWDE4luARjz0+nf8Lth+Pjo9QTnPy+5mOKiHDDGt4Qyn323N+GFe
oe3aOAYXK3LaPSM7EQhKmy/OEizEluUNK0bfLxoCP8TCOr9wDpdJNwSbiYtHuzJ0
EeqtNNjdhaCxGId7I3qL722sd/6VEH6tNw1Iak9+o1tgVa4G5t6JzSk47oSNRDGB
OvblFg+Su1lgFF7GrpEASFKBkxVH43HqNGCm7/5vly6tYcgEJRg/OQqwy6Ja2WJt
o3GEjyORaEflzUp4J/4HXSArWTDgB52Nb3dkMLPQlltjA0N84RpkEKdhn4p1VquD
NqmlRRu73cFLxuK+0C2YtSZwczYTL9mL+wpO/vuiBfh6uH/T0B1TTKuRvgBt47by
0PNK32uZ0TcPsa/c7qtjOFvpCvNcIO84tIXQ5k9g0ePZXt7WN+2tysncqCZktTOQ
6JHy+1GFa6M8j8QJem2EElWYYQfyDlhXEpetqkxB+F3WmQ0eHX0vA9cvndgz8bUT
I5K75Zczl0ocBeUR+0h+H/0rb4OaYHNJ+fVgGBDlpFlqGVhpByBWynIHx/PrP2zY
Vri26enUgasAzL+4HEnnUzMT39Ux/VZ7MZK/qWiA5mZvU92HaP+Z8gQUIOWpY2u7
H1HlZu35qUtrFXVTGN6HfzgvPqKSI+a8fr3Tjtxd2RSMuSemnkzyCj66wk7lk9rg
NrCNZhuJZzidTTAuBdWAekPLVNmhWjFormC8pgnO38l4YIIEwY06ehYTCfrhd9GL
nehjz5Vx4VKJSKGLMsnks0s65OHtTju39PLvgFOl8X0sxCU05wXFxO6nLxYTB2DJ
HYLbH5oc+tV1TcRPVM4ShF1o+yjoGD0fUo4GoBsf+aXdhZKSu4MsCt0qwuHODMkf
Jx1s8AjizR2UyfEkQHHPL2mp7HqlhdBUr3E9OUhXWikkLTu6hnvasXCAsoe2ppfb
pn8zKB76QJDZodQqYedKBxLD1aafSB2STXpYm8kMRtCP7fG3PYGJODFecErIdyJA
OUzyPATqeZXUqeffH02I0hlxBytCTP6fVt+25QOY1sTY0jcMz3kp3dVo68jTid7j
wYQ/6pn+yx3L2clmcB+MkgYzn+J3FYY4SEj/a8lhAGqVvpUZXCMmrFmEDvqh3rR3
/URMZwgqreULLLFxjFhnO8wuFJ9fCGRNVkOIjrINPrnQj912uHvmqv6o/GBfeQkj
1/WAQnrb+vJaJoDdFLFEIv02e49e+4017nxht8fFH81GKfvh99zhLNs5T69mFvng
MR6Z8RqIXMf9qgLBudw+tOY+ngZQOGavJ9n533oxdvonOWEEqftLoHSU0gCxoSC8
p/9Wxi+OTWj26mkDmxnBtsyBSmZLQkEFK4n5p60Yn+1oZmZwaE1f5zWd37ruDHG4
YFb95734xqXe293rGab8h5mSVWZw+OJMSpk0DCJSKBwhSGymbFvihB5JuYwmNTQn
QguvYGMCykqYVj00wXKlmz/HU3ts8md10bLGjdUeB99vwUjQLxulac/W/dJXzVJR
bwc7+GdMUYPaoeM5dV2flpBu7nr7QbaGX3WEBx/9IhljXHlSedBPq0Y/inSyaHEv
pA6ghkkXCnh+7/WEKrIWSe/ASRM14+pf+JaqX7v1WqCvdLiu6Ni5HKXjabUafaf+
xMJQmc0g7B2NCc8rbWvv651EcsfPibAarw78SMiKrkkpneSAyI2BqAMMmf2TzPsj
ODfhR0gA7yGqmRCNDTq7SUnzw278m9jdBosozHIdWSzfib4UcO0mXuPoy8Qe8gM6
H1PHMQ9MP89MnxHR8jObDN5GBNE14B6JZsnuyRAe8GvMztAWjYqxLPxhun8vT9/m
PBGZ/nUKta/ZocjyIU7rn/Cty8pRcvXAA/ZRmCU4AoOUgpwMkaoPIELItbYE2Bd7
8+R7KWxUAdbBUOySasSeBFufyjIbDRUd/J00PkEZak09b3FvEdNFTYsTmki889Cx
RH4/oO1I7k7ec2KVS772U3QA/JIDQAjRzNYxfw9Y+PuwE5a1jLiicRcHZXzRzpzc
h9DoaXjraqcWYGAQ2gVIw7exof2AD7lPkIo+XQXlxSC7GQ4IdkEi9nPXx1dtdTcN
PIqRD4tmwXacIEklWkVt1dT1hh8F2Xqb6cjKOdyJha6cSO8hC4WKskRDULnqFqqc
+K5+w+9eVvJaROARUA3yEZ0JxA/j7T6jLj46ib0AzFGutKRlkL1UW82dFngM8rDp
QOHFsZ4vGV6j3ZY/1Qm9oE5e8xBnxJPOGHR1oxinC6+G/rXDYEhqETOaMlw3l9Sj
P83MjHrhxFIBgPawtETky7S9Sk8Ei2tGBoZCqvop8QQqb+jLuaFnUatPsi/fxBc3
oToPwD0WSse9MmI8t2H9f0NzX/Son5O7HBYgFG1DI5nkuvSRW4H4X7QaJ6uE360c
gssc/1fWyMUeC8Kb9xVvWES7CgDx6eBRjE/c65H691TXiKxgPbbE4rHGn/Bv3Br7
PvlYUFzPeCQULdEsJIpljSkjCZSuB8IbV7b172Nr/Y3Gi6CsJCgjZrRWGEy8rCNz
M4dlfW6EIH3P+T+DuEh5ZnRquOHkLDbda78rAyc0yfq2d4sZHdlKsbA6XdQLphTZ
Itv5T9/ETiTKYS4/TXYYM/SkynPvm3JJQu15UXE2hmmRBPGed28UlyfWQ4u92edH
TcCs4fCPVf2/KEZDkK7dpUW23YxIq9ss8aLtt4H/R71XMXEJupnzR7CSCXRGR/09
SPhSjm/2/6zEvd85s6K050/JXCtyovbYSfRkk/MNPR4QKLUahh0p1HtZlGzEXKS8
MwOdyqUAqluyAYdA1TWnAW5Kb97nsT4zZyoR5ykP9zlULnYNnKC5AbuEgDWVJUhc
r0cwSYHKjVQM5/a3mWJTHjV4Zoojag8aFDBjRNqlMAtGch9yZo/OAXimjwBD0EoB
yXf4l/EBYIJkEaKVnwohJS5rSU8x5E09rYchVYdSZ58524xkluL+RH/kAooDwWH+
VsgqpdFXf9P132Rx1Eei1g2Xh/iKWzvbEVJXOW8lJin+81hpSExwWccazHLHWI6C
gnYDaVQB7grBd4gdHYeLuHdb5XMCeo8zSJpM23i1W8V6QWnbEnVAZsQ26pDzbYJ8
9vhkEpvafIsKumdpVkOJU8ZAg6k3gye4V9K/VRoZxchybxE5z/oqqgmq/kXlMEBK
mSNTxZRn2I/oo5NFPXq2sj9WrwEqADmbs53Cb+8BElgHQ6/UO8REdY0UdQgzIHSm
DgaYGPzV9Y2L09NzPY4Flpu6TInWOI+Si7ZFCvANZ9WlzqM2AifbwnDEXeeENBSS
JiFdm/Sj3qdnwDEkkT4EbuwpsjVx71y0KDk/acccnpgC2QL8QsRT/nHv+A4Ckx7V
iFFEDM7bgRuhm0g4hhHjDw1H7hLd5lGCGyu5bq0pawLCm9pDidtQ71ZDP/tMfTKf
TKoQWuv/ixFdp+QkNRYsz2XB2/wseB38Z8yUe+uuRv1PqDG5NL1REGOubRcW0Ry/
QAxiupWOfXiRBu3OSYYq5XLL64T0Y0Rnm07V3hAYO1wFdxZps4bZqr8zzLj/5K9O
uSPk0+WvAjwRg6y6LXFejteepMJ0C/4CvGEH4blD5tj4ZSbu4idGscJ1yv7q9GZm
X2F4+oiDZNYLn1vKVE3TmW33TIrdrHXJuk40moOCRpiimzjag5DYYZD6iVNNldxP
uEJNczE8+SuN7rR5mY45C98wEyDDEmS89nepq9V28WrsHD9JATZyv0nUQ+hcQ6a0
N0DPIcFWD3I8LHX+xWcnZGriIz0zmhGhMWwTE3WKeAJhJVKCS6RJtO1gerW//vxc
TBMqE6LYgRyQfvui6a/agcVs0qoTk5gwa+ocddTfTVJ6wThw/QZD7IcFRlXTrSib
9syt0RleKNF5Zrp9LKK21euxw8oHR/MYyUOGsypO5WI1WNSc+C3Tb+dGkSRCmkST
XYuJfQInAZYnMZL7Xxm1Gt+MFZI+iiZEZ7o6xawbh6YiAMIXj92ZJ5IPfhMxnnND
M+LPcv2pLZZDuwUD61azT4nO4CAdPiXVsTMhFXF8lUkT7AtqaZASYs6ZRhFO9Ypr
Rqp7ibTsZCRUqh9bK5E5YOFcGdWEMiX4+uxAITGKV4HgrvsETdDIVLQbYjP1BsIk
Y7G7c9PyTIHM7lyRetef8NUjWUqxfkqrfAOGL+cKidg9h3qHc6fx0gNlj+G6FGC4
say0RoUkAtPxULjQPo0RpvFnBYWxWUCZvVvjULw8RQXwsxzcZuwRbdHcHzEuHlDt
7TUyVHHpnEgpN2qM2hBG3vFoaqbMnM1HRZ1ESP7vfQcy41CQpvakQb4a4a1RAbCq
4oCn4p+uvaU8gNrLauY9wzNpbjIaqRG5T4nTwmkTzOg/jpFqYiWwa340jgRmyrfu
tAxMKmpX/ACcbhJPNkbTLpOXRIUXkYC58RF6kxBz0zd3rYqb+LkTl3czDYMp6E2J
VSbzugNHlDv/2UWr2RxNZoL1MI8BMgpWxqh5lCYbZ6OfzqnkCPJ4DuUzR43uI67L
pov+KjrnN9oVPI8qPl5wLqyUrHF3c0/xh9kh7iYk60Un/t7CgTp3NgflHN54wMd9
Rt3PG2sMJPWu8ATNRM7WoWari4+oPPtikr5LC4G7gknjT1YPFUpbPU4DQuheVP9X
jdqEz6nikDjZc79jaFPohWGubzhaLN1nAPCG67HplJmD+7Yu792julpZ+O70xLY3
YXRUNXmxErE5SzZjqgGtdoJQ/7ZataAXnY48iItJOT7GeVhyM7Je9GtztEbSKkw5
gi6KKAoVWPG90L0zgGINBbRzR+LZnjkQru+sszXh1yAxmKo6tLaNh7pvMcvoythO
aiFRNdsuWUZGpY2x0/rDFf5ghb9vZM2t+IBuABoVuQmPdeVYBc8j4z/2qCoB82rh
2nc1L2UzQr44MaVkKluBGVyNQaieIxVckgGIZKlMzdL58AAFIyI8LB8k9FYxVhuZ
baxEpPFgTVZinwHn3sZ6XyqZ/VRU69zI/RMYq0J26iV5c2PKJjdMlXNTWy2aGmVK
gs17t03YNsTb4D18MgsOHh+i9LwIKNQvsEgopXLFCZUYkFbXlZ+Vx2WHgBj7/dWM
ILe04RXu6MIwwxHlaUCQXJYug17kouYhkY69Sxm5tr1gJ5MIz9+pUA9crAF2nHHi
eyszPR4Ktoo9beECioIbogK3bwyLKztSmvsv+dipwXkFcFb/pZGL1HvwrsaAxnmI
YR/o4K2p76ebQ0sgKM2egOUuhPdS21pnPDw5BU4cRir7/LXsgeVq0PX65zsPKctJ
PJBoYVTm5Ot4FNLgTsdLLxY0CTglHWAQ4W+dNC0HLuMgXoJXO+MsQOGRmbi7lZOq
IgTYfd+fZbK0xzUP8mpyUBrrKppsgm6MJ5kMgGIeNcuNtK9jGubZZaYAgrwfR6B5
fW0ZFKgKCjPSkygDQIZ2WDvrXODtEp/1y+uGzNU5939Jhq4KeET/qQIApkkVC2kd
2JkgtfA3mGNJ5OPqPSHLUp1rFvjeOovpYt9P2JnKRVN0hwb4xDoXwlqwohnoDEw9
MTmZlEn1KWiNhrqDyDyETGij2STYSSPzFrTcL8SGaH8IA7UF1xKXcgQEP6WzDIJC
sTjjnjd5fK3VvHGRB1Gv2EZvwxxD9WKMBdQ/suTdcHhGj3iDQGtZgYByYG4B5ay3
5NhRp2mWXqhayYQdJ2pAyWiGSj90sIzCKjxYJvi0tHFYjIsquJExDxLgpUF2B3ow
0DCVGopuYeygRpdfTNHtSTlzoEug24Cp+FScpHphiWqH2mR3emwgbUJuKVtta0DM
xKGSjJ0LTdi8iuChoUq7R1eO4pGpLJ5dAfCt14WLxY2lWa/KaDWTwoCjD+PvPLyP
qKaJryL5DehlFOFC9mEYLioinQm1VH4MbFpPTcIp0kwPMW51cEA9+gBuufeXaX9A
D4joyzCXQljDzU0JK+JlJDAbV6re9bLzDIgnnrGkZYhMvoeRcspDsmibAl8xnkZi
92MEld52iJ/NStsYqz/vbZM6Vx44Up/pDNJ0ETEmzAv1ifuHprkYvrot6H9tW2bq
DLH3XRTtj4DJBtN/mxQP6FOVPlFGpG6llfNT3c9tpmfJP/C4lH27VDYZxLEz/rC6
cPP4fy131W5reZ1DmQRQkyip562DpskOgpiuk8A4PHN6s9BF6R8GqOZAFn2R9kqX
1/6VX7a5eMPKsihEE016EVjm2J/529DOJyT7xEOuMDPNEfuaticNH4EuEKo1JwYj
lIsbiz3ojc1/YEj45f3jLulFlxP1i07O8LVOtYSLk7IXVwcih3YZ9NX9vV75fFoi
NybHsYksauT/NaJGHu9AxYdpKBP0YUo7ThbKjDLzKv0uBNQBSRt3EEpY6er5c/ND
T/5BB7yG3Gsd0wDT3iZLeHyx7VPMi7FxQD4ZMayX9NCExIiPr3vMuG2G8J0d5AKq
WxJ34HUJPd8Rop6SRkGyKVsJV8w2b0E/UR9O8tScibHxpXP/PHvz3kahrmJkwWOr
obe5TGXtHmRY2YERA6YUHcyK1QVgAxDEIYePHYmkCta3hkJizPmK3r7R8LAHJtOm
6XHQ0BOWeDj0n5HAnAOzwIa63oJkTD/M/NuGc0Wvj44PlASo0VBOtefvLIH+r0kw
9QbWZ10pY4cx/iiUt4BwJmEWQl0RV96LrCYAHCAIVoZKoSi1dM9RQ3kZ1CqGhvNO
shtvGsnQV4BLpGWOG70hMHMKc3uHWO0mwKMQe46H03TgTWhO7fGX8FUcHxqvCaFu
HSEnbIVqWvXY5cSZm+DlMMaEwGgNibcs2KHufy/JCijwX7tGUdFXxkmwwrMpYfAa
Nlcq17KHV6CjL8A+0FLX4iAxgYiQWWxGuaVOhm6CObnbIx8wgT2AzT8oDhnaYVTr
5e3Sly5cT1h/lbOuziBvS6HRA6mO7wtFO5UDinDtRQ6TO444CP2XVffl7cKveeNI
Re0DgKP+tUQSZ3XH1PMgpJ/ZuQaA0obhq5bXeWGXGBUDb/MQki5jwFm0ihrXXTXV
Yertn9qp7gFQjilRExtCK0PKherer7WJgThIPXNcnOvSW9rSlNAXUOhmcMmV9i6R
rwrmMNvQKqdXnZa77BK0B2ueuqIL/TQTmiHBiYxr4PtOEGap1IlMaKqo4rJka/of
GVh9vfFMrlS0QfbU1gyRWiB45nfCyrGqcmElaHXtIhufzxYUPciEK2xniANG9C0/
i/79awGK8jDMtN4agTSANMhG1Ck4g599ktXwHMpgA1y530i5FzxJDhzCN7IAKiRa
WQOTbG+og62Uqc1C7ldYydb1DH2Ck0Ykixj3ItBdz4N/GnqY8ZWssu6o/bnIHKXO
MtHsG7iBzo8gUKfDRyklIePl8V1tHof/cS/y204lu+g4lMEcy0ccSx9IZAAVsq7u
3d3tHx757//1HfxgUkWWDR+bS+2hrIXXnvY8g/FFQzHPTK5riG7VjteHywezEby3
Mdpv6xbXxN/I8ocMNur5fRWAoPaS0YwyMoyIYS8f4wY6ap/4c+7GaCIVGoxM0FLi
NzvtfJtDvfrfpiXQ35rFr3E4sMomcSh+GenuaNMMkFJGEQ0UWQXsWD0ahg6XVErf
L4IB3psfFBS1C7olU6mTLsXy1F9V3be94RY3b93tUzwKWrf4kcwkdMc75J5VkOYf
5ptU7G2slHaSMMirhFOQWSE3aZAA5vK4QiXST5NgbnOt1Gre8QUsEKevLqK3itUw
e6BCXwv3cDKxwF43qmRjpc4Rxh9m0SpGRBI2yQFgekQu04y/UULOt1VfdkFqX3qE
45vvHeZMitSgMvE1695OG7WNktpUD6cRk7ivrsLak6Df7j3g3nTSKdHnDuATo89l
OeR3Sm3Js4cZ8sZq5Zji5LrVvh5NafH4HGegid8PrcrgD71Bgj5wPSvrz3zknZ9f
vxIAkLMsW8IY58ehOcecK5/Det/OIPAaJK1Hw+CXfR3L+0xlMnlch9XI32U9y8PA
q3Ku9SuP/eAQ1wrbgg180NY/p5Y7/+7NaIkNfFEfrX3dmwhtvcJI3r8i63+OH5Yn
byqzEQwZFISIezelpOt33usAFmtO8YuHF2DXJS2OYcGiSURDNSCGgL/wBXM92u9I
S6tzXfBPS08zqi+eDImjyfwshKP4g/2zFMOLwvRNumS5d0RjGlRAaKe9spU7oK9h
KDHKw9pR7G9ulxEgAL6BgDnxYnjq2L/J289wHr2GIust2tjlitYrgdTPLthXGhC9
srw//kyM5G+77A2vXrrnAmcRxeAuW6CZf9UZArqDX2sJw0YHgzGnd4Ip+9duTL+1
g7aHd81NP8CB4Jr1ILBT3+fIf7fBqaKD9yK7lSfEDmUaqh3sl52I40xdMGiJwdz6
18IqT1OXOt5M9BYGnoWC4EhdqjrBmpkef0Qg76pECQObQ4zuzsLFojoksyALtcqs
QaZJPKO7wf+9UzWfyLerxMyQpUdLx35A/ELt2ntHRt7HrSYldgEfUPr95s+ujKLA
KvYApbuxiVPxCogQToIyijg2Gui60ZQ6ktTd/dnFhL+ccq0R8jfu/Bn+bxSvG/jf
X3gPgBYne4NYn3ZFb+guAvwViHvsSRRgHfJjMKdRYVZbclpgfLW0UNcC7RZzWyEy
y2dGy2+/q+y/MaO7aRoaxCEnC8s8bkWWvd1//79Dv36k2CGGE+Lypr+SBI7WIHl6
+Twyk73siw1E84QgkFIhj2UDTr3sIZOe9WcywqjUnYNLkRBwvgbZXS8KsHMBDtbv
Lz/zybz21+yn3cLflbQe67ChtgifvuUoC9lPs31OKbRB76Lrhb8TbD9h2sBWCr6n
AhkfZX2mksnL2QqEprav8caas/8Dykx/TD3eqwgd5rxBwbRGRyso/O+lFOsxK4vV
ZXNCQQLk9EY5motBMogdeflAdg0iL2B5zHaUtzB5CJg7Fk8ZrtzMeE/GETj3I9py
/s0elBYX2mjnVrP1c1yJdk5165QxVRro9qjpYGzBOnUaaXVEF3MsvaTmoaxPnziW
z2Cbik6ngQZaU+h390UuD/YYRjdRmCe5ElXDHxjkUfQyypCrbAnVvsmvXUZ1eA9O
aOann9fsK+DhKEi/mJNINI2lMKL7uARE+s88vqG/oqL9wTDfppPPu4csT99jK5UD
e5TSO6G4w5Owo/fIZbMUpptpuC+snrfsfoYwyyrZlzTYZ9jFafgA8Y/0l7p7V53s
qoF0gkMT8dO492ksz4puKsRqbcQwDHHJlP+Azrc5RaftpIpjE8amAMaAKa37eFK5
fulIJyYE0BwKGwC5V6j0WacGQgar3j5kqAoiZHqG+m17haENVD6jkOCL78cKZwVM
rlvBtQt7W7dn8xdYUu//5JU+ZFEGh1NHVEoOtQNXEjK51MEWDOyUdJlLnXCITDNt
Dqj5T63gziKXY11ugCs7qf2o5VP0Bb89pTPlUrrPHw0P9tMvMbLnIaN0UAUTfWsB
tZtcOiLTHHKjXCNyldOi/By0qLlAA0J3jhPjqwP4737ZzM62c6SfEwo+FvdShxn6
KEiWpt98zhatDRcSDuC3H5rUINwyJZLxyGcKVsp5N0f+EdQhsx/gnjNc9h4RcvGu
leB2qkkeHJDDXq1gcBW1MRms5XOaY7Tsya0esFyH6HkRM7djMUgjENSELlUCa9M7
+YTLGef/YKBsAuIzFg07JF0gpSPPbw0j/69zkZj1Dz4S5HXx0FXRIW84pUc5VoA3
4tQiaBOjRI2npScfUakC05IbRYZblfU7unIbK0/RmDBMVk8SojkGg+T5vihsx8wi
lyeV5mtuR5sP3/loMFpKWZb3lPSW3GHF/H1z1wVFM0vB1RgjDb5MCgW85qoSLu6W
SqirBQERLqbktKIkgpkl/QeEhW4u69tr5nDqw/Vq4hjrVV8o8uJOLtTz1cEuEW4h
xV6nFh8ezWa6WvV4hK1/FV3RDpl3m+SWnph32eXwW7xsFtVYNKRvFA1Zymx+Ebx0
GWtYZNRJ3FWb1L5NygGfNyDyh4IfR41+z9wQIets1QMLSXs2XMYeCbJ62L0ktg/z
5jlTiTgQ63+uSvx3dDVdmJlKoyI4NaGVrBTuG2BzZqYylYRl2bjhPkG/UPg9SayN
SFNX+92ydl7qBGqkgGmGVbg6IgtmY86V2TEvox2udOYgTL88Qng0kgkaDtAdrQWk
9XFtxkYC+MdMtW8SXE3v5r2sURUjiURKXaGFPuxRU7wqleT9mjzRgcadgJDnFlqt
WtYXIo/sWVc3dN1QSIQkAKfbCV9/h57J9vVVH8EJwbyNIT5Tf9KhvW1qbMZ+NZ3x
I3Vl4X+YR6aG/fQaINIoNeGjQijzZi8izfAJ42+cP6iIEuaiKyGMUWJBCICOij3B
MkKLScH4QgRFoj34lh2q69w4wVMCkqaF9SMOOZSeCLNpZSVAi5d9K6wVYl1OIFLT
/4I9pXyRNWMnS5vcX5K5KmA493D+Hmyzl+ibrje86xHUTELypEUmETbJiqWIvswJ
iOfBcXd4RwI2Vzji3SFn+4Blzcp4S6DBuw89wOFVzser53fcVKY+PEb+vsKuaN0A
ukD4WM1LbQ5j0LHOsmu2SbwTCCiIzOhr7SvMyeqnrqzG0iq2LOl36XHHf4Kg1Zsr
oFqcWnCjoPTzQlUt+UQyCtYgrE6Nftk1pnpvf9IOAGK9ofGUlC1mevi7QXiB1gf6
/tcPs7BiYJJBXcBSfFRENSn58lbqXfCY4NPdb1WtbzvJ5ubxa5/1avZCNH4vGBIs
MF0zdFA0N1ho36HoYJ7oWv5FN48rtFkkucJCeXwIMxStPy1OtKAcTrs2H2WoTL64
HvWyvpZ9dRHtzhHy02AfeacfC1fwbycMEposVi5HKaEhmzCebj8HT/TZ9YBx0K2b
obRZfmzwA0M5V1mNso7OpUeee0DIw/g5RQPX3wvFfaACzFsTPUq2SRbyfWIBy9TY
6HflDo6ERaD1k8WvZbYwuyXV6KeXBQP8QNtKf9CtDLBsKyC6IHfCyK4dJk0n80M1
YRgjCRhLks2oVf+juXnDTFFgcTDjnn3OQJcUSbeNekWOb5W+5KICGKfdyLwvXU+i
MMVslUaTddKN7zqwrky4JVIiK4RQlYSoD2JTHdNTxnNojheW9MIxbncwLzz2PUxn
F3yOtdMBjpUpugZ7bmJnmA0m5mnSbla6r/oAJh3EEF/dfYnFCIZanX/XpqlZo9Lu
oyWjkQhjsWN7zMBmKbpr9ZQamVRmCc74l6sRRTiJIALvlnkz5RxK2BAlYSteIkVx
OB6uxfEfw1qD6uTQUe8fN3R28TPXwA2CtMkX4+qM5G3FhH2K0fDiEHglsAUCy1sp
EdzN9gPIj7mw9D2QSM92ZAnt5zXe37SioAd3PSLUliV+q+PasxgrkcJrfW1Q2wFX
a4smnq1JlgMh7DAFZRowgV4XuefW16PYpHXbCBkG5jxJ+yF/IIIW5qOzaTmOCVlv
Zar/vTdjcGc5BatJG6Mw4CGZRJmkvJ8PLzQTCK/LtvvU6RHi3hsVVu/AdlhusA81
Jqi2m3YHKZ9AOrnl3jUmv6wslNsrb3eAOVPPxFGg6J8E+aqBoMO/rs46GeU24+rC
XYH6p8yaQ1jzr0ERhrh6vOE5h2L/JN3Qr6vYCF4ux4VuXNamuRK8DcgAgjrV3JXt
kw37nBTcUtdAB3quO3mqYw9xxn3QviQ0boVzhJp/bQ/fwtTNDhRojvjbrlbSid5N
3v0QMeOUYTTBPtcNR/qkHqThv+NjGIigV8RmBuzsOf7xmzvd/6E9zKjJ1wM9x76y
+O+PLTEyFpFl8Z/5o+M6wM4rOeolbqNwyeK/OHLyFTL5Z8g2OAraYdtgzBm4eRsB
M9tSv9sdttZUZeMqzYD8P2jNPxu1HzuISvaRmQi9javfmcDw3CPRUDVLw7OJ63dC
1VFRoldfbGTAJnr5Q07AywNSNyktGwOkZ7tJna1EjS4uc8k8EV7B8hd3mZ3Av5Vm
rIrW8F4cBw966SKFzcBffhUIfP5cI5jo4cAtyTPWfFErDkTx1sUyC+nsFbDYmGCY
S28mDGYCynr/ie4Lx2UI9RATZKygNnJVko+ZDL5HsnGuQYvly6pc/f8j3j0X5NT2
tdlbELK9DBBN5O7TK3mLhyOVNQBYQ/QkoMPWWFwdkOjpX2IFWO1TxpfEqzSuYJNM
bNTcAUelz+Sve00H9tWpgq9CFD3HcjeStuw3ERNM4WXTfMt+WBrc++Q6+mCxqQqO
+NwHhJ1+dpPSV7NzeqO13qRAVubTppTbkU6GUTJhpY7iLDdhlHEuh9HWkxgalVTX
1GoE8mrIiltuXyo67elpgZOiJrR0L802drHyS5LdEr3T4Pb+mkjImEZmWkEmM4fr
/pcw+lyx3TR4sjSvGQWgcbbMaM8BIucY+Orz9q8yaqAu3RrozqoFQZdVVNu+f1zj
GaUAl6mzOI7/o/b23nDQRazh9WrcKOi+kTGzRx1TqUmhJ8ocvCWEz1gpLCS1bGEa
KKgaqr9YeOLQPkaFCe0CFY6rhXVgx/FKmE+2ye0P70O65qDB/gEMSD2GNuyq0zZ2
L5FjZZ8zBgktjGnM1fa5btxUJuseQuubjGlv1aggHBErAdDiGhQNg+UkAlWeAZ09
+XS2bUnCVx01nwDJ/W2aUsTXIqQxz1h8rURFEcRiCR76i+qDt4JCr9uC0ia2YJEa
Whxr3uP7grnZN4xWrawoZsnlf3DPXGe5bk8WxViyjhB49fNFSBo5rq7dzz6SybP6
u2jn7i0ebLkOY3TTvvdu7B2mejqNSQ23hnccczs/rQWYOQGVrFg5+VvYS741p3wJ
gkhYWFl7waS/gGQPHpx+7UBYVn9+ZnO6+74ncONLO5eSdyH7VHvTSsCR1NmBBY6J
1Qe4lqvujw6wS96d3aAs3UABzwfmif2xuTkxdK/jkNZ44TMPf0oZns6EAAuuM4UX
mp+n0HDHypblAOaF0lnEeLl7K+eaMmjI6A97jHfbeP4rmUrxSv2KB/7/nNlWFJUj
9/Nj7Z0KiI6pivPbQXw7tu7o7xy8+30HhQ+EVysD0vUjpZBbhqiRU8KR9URoJlcX
b+PFUCc89/6aEDt9WFy8oWLyt6NkkBNYVDnMsqRaiZi1A5AMbEJ9GR54Jp3KFxI4
cs+J0hDVvGScI/X0Xr4jSdDkpazcdcNCcGgT2ZGZN0vrav6bz1sFPZbg5IKv9emx
sCCK0I/u6oH8FTR6v8Yn6ZiREPV0lkdE7PYv0SRDhqqyAtVpP8mjQqw9dlvkYD82
kSAD7qD9zMbNpI18iMHdbrqmCQte00Mj5L8qJfXMzhBSFIB+rQ5rSOtzSoiEbLJN
g+jASs0inwqD28oSosOPnGmuiIf8EP/quTQnAr74P2y7RrIOrRiQCeqsCuVL5rw6
ulutY4MUTM87BjANQfky/KRUx4REMf/mC5e0OhKYUebKyBawJUFh6fEVaJZMODNi
/CBNnkLFe5rN8IliH8yidcJBrqHLwcmQZbpsq0uqM3Ic7qwgPHt8XJijq2mIhED2
pOhcFrzuDWu+ct4f7RgazmgBmIJw7kJEVV5GoUdcCByRfd6FvOjJdqpRbuh6Ev1G
zG/SJIdko/yam+MkY3S9txxLd0pNL7uvEjkntoElKYstM2yww8o2z5Qphc8dHrbU
CWQ/2G0PYRRydBL7gRXQWlSOksbzav9dyECN1BwDfyxOticLGt/mO/Lduod51f90
bWgniyeJ29Dpy6zwDwyc9C4l2w/WZtPVA0CJe/YqxvFpmddfJYfX/A1MGYP3ba8j
zrMlTXv14qCO37KHfpB8ZdzPUM1VrgGnNQqjrw64ehNYzqk6CLqtwtpq4ePqBGUX
kCxNpow7/rG2rKG5TbGkuDx27kf5wVeeKjEDM7pjKO36XhkRmpefmaJfNwRtQ2M5
AUgLNmNz+9n+vEJhE/zptJLQzB9egb3U8kHgCLhhYa6MF5L81fkxtrWl2OgkBi6a
nly8LOnQfQNi7PNhjPoNrYD6R5cFRYWdSKgfDHZnHilDDFsL69cZAlVqLxHp6eQK
9cObUs5DoRWb5D8sl+9p8zG4gml/h9MSCV1BrX84oNtk7G8XSzx9v3CfdPGAjrOd
S+3Biqo5ITqlvDeOisUsbsC/LONdGHHvr/cJSjZWhcFZhi2PJ55X2pOt/oomyzwM
DlzRsqUCmi8g/+uFz5/5VHhkKsSUmVrHNAWUYcP000X9RmkSd4apiNVmHJ1MR5FF
WEC4yo5Xx7eSmEwsCoNP0B4p36XiX09D18vDUllSz36vHkcI3t2qHgC15dqymeDy
DAj3cN1ynXKLSkW9qYVbRtZCUAb3uYL0wJaFpS0Qhc1VRPfJzFQKhmuhJF2bMb1W
ZjHoYKfKnpRJX/FfaS6hNqr8r//Vt1By4lYcavVFZaEpC1fR0/EYUjUkHvCqJ0cd
9NJu5g0JB7Suv/7ez30CzOQmU9JMpC4bnQO2xqYpa9nh5GsyR+ApSIKQk3crnYM9
UScDJMlHC1kU9LMIHKlb/WS2bUEMKZmainXkR3K9mbNgDXFgk18ZXHoIrSYXKYdb
xa1FVqy/dIVpxozCay9QCX9Nt4p4WXf60/uNOeyyRHwks0f0Qh2xcs6K3xrGEL5G
Qz215ZjPuZfPnFtOd9rofTED5Kl+gWSdcKMmBvmovFTrf5tkFHbkauAixG5HLP3L
JqoJHIesxYH0XTyzIc63UZzHBNZfP+iHjV+gUkuGkCvH3B/h5bZ77wa5yl7hx+nQ
eQkuJPrzL28dux7NzqimKm5cNuce/qCyWoAIzUlMT2aBKAoYPB/Ne5eVinik3XkJ
5dzRmVHiq47c8lBqJ0UnGyEyOkw/UoNh3M14P5D0jgZ844lt7OAouodHNGDJJRIK
/bXiuZ7oCrIA2gZgBsRkEbgV+Z5+NtjGbaHhFCxkyNgmxu9BLNOdJmKXwR2WGk2c
pvyt4Vm7+nIjr8E2ddlwgqnverekgpJYS/e9cK0ToX9Bk7BcN0lly1zGav/ti/ZA
IQ90e8r7RprOciO4nfvEFRw7pPVxNLWmDuhWGuaDmXRvyzWQkTdAjIWKOPnq2BKI
QLgE9ONaSMO2fpRm8r4Cnu7MBOMXPokywyi+xQ0TlbRPDXttYhIDaBm+TAogB7/R
67YF0RQDd0fOjTPQ/Xx4+wRUt286uU9Uv++S+jIdMMgFPA9jqFxo5IAXmqlo4/Mm
lBGSN7FzwAthu7tIJJmwuOCQhoK8Ax0Dt+g61NkimpWjMMTSMaIM442h63TrHxse
KOaWAOq7/uTQSpq2MD91s5xSogorRB9ZRsQsvRSrpc+6ru6tc6Go5E6F8gl++3Hb
dEBWYT4AzpMSmvmTMRoFHWtlEhnTNv8BrZ6XprwYpF+SwOzwgfY0j/qMVr46hiMX
QGlVWb0g5L07/nxQcfb/ts4RUd36HhSMrlX7e9S7sBmdr4qzvrQrbJDiKpZonLGU
jryor0HxWVE++ho6ChA9nhecQvwME8EVLbgncbjtl6QladgX8CUDb2n3d4p++9SD
4KCzCL0ar9+PCrghXFe9RIneLdTvqdzvNFWpwnC95VuMgqV86ylgTAu4bQWVtfIU
G7uTvd4x2NZKaJC9z6gOFiOJBSmzwrcFTKorW4FQxiYTWVSbqeZKthMDRHpYNeid
l2Py6O0n+PUDmhILk3cqRHs9cPz3LIDE2gC91BeWTDP8ulh9TD1nR8Ig5gXX0ieE
rkBOBTQxHr7pDeVKOdGm18Fy5HltS9XDTLJg7JlgE9PCTeH3qV7hxKAQ48nktYAO
XiigWygMhsS0RDHJQm5SVJUcbcz/M8+fb59sEW8qlmi1cRbiZSRp/e/nnWgKU7/R
F5iT8FdfXl4LK6c54p/zcS/vM5b+zbeZ04JAFbJ9z3nOQgXSoL/NFnvdqySvUdEs
YWSslQg3ErgXO+5kYWTgNLCD4YLBW2MWfTs0y4DHWr99Wu2NXpQzktjMlc1xPEM5
WbZcd7w0d/3w8BqeY7w4ZspklDvGBBZDwlhzkvtlHXu5sNuNzDKasuh9GGzRoamK
wFFk1OldDnnP9vyEaFlb31cJ49IOA2NL8V/nz2ymOMHD2DyWB0+UnB6ZLsvYOZwa
sQi1CW8J3oJWQw2KmD4kcbATECr/GvJ4yEyHIyDLhrmVa8k52ak3Hi9lpn61cv/Z
XNvB4ERczURGZ2JZIW8VySzG0L+tPYEa//DuredZxNyivfOhbIHDwJa2EbLBAD2t
i4y5F0HP6pX7RkOr5VRxjSYXugi4yxbJe7pDUdRJnVIM+yqad9/D8jJaXQb3iIIi
DPu0lyAFGRD87fLsrX482VdYnoiuvuYDRscFSJ8oaqBuaG9p5zJgNetP1Yx0dg7w
PnTKclYTCZJaZetPmh8VlzK+QQcUqfF1Rn9h9iby4UFMEu8D5ttI+aZWZx9Kvmit
1unf8QVC7Ce+4H1M8CYRQOcJ9K14KgWx8VuCm09hCnTc2iQ95JtjI+aS7CWOib4J
VUjAwhWe4ym5kzsbuQii4v0o/0sFVsh+1iEj0bMVFp89CdKC3X7QgplpyvTa+Ij8
GiWuRygoNxZvTVDyOV/W9KNA696nZ2XxxiXCRtmO4lsgF1JzRq/uwix4UJvZCohM
hy+WXIsQ3qRBItTH3oXoh8+MsYJeRJetdwHDD6eNcR5BYZXMgj5G4t3i5AdeHXnY
fM48xGwLiP76Wqczk/HIo/6YU6Gc2cj491n9J780kY7YLqPRofmeCnmElvwkxZW1
ofWWBuSqpvRFvo9imwopR66RnHnqiuJgV3WO10PC1EUzq+eHJZC6Fd9+IHDK5BTl
YH9x9Noi7quwGv5hRM1lXBnVOU26+LkQOIBOrSVmUzt4JUql/z1oBb6I+3Xsivpx
0uJ+fdN6qtU+v90/2p+qbSZYxqLaRZocnHzD+si2O4aH7fkah/VhDwe/0lXn6O4M
6IDjDqU0mB7AEza6yGl0EYamqBmg6ymv/qCDT6iU0VqU4h+ED4UB0AwbbThD5TOr
sVt/WQx74iLeQdWMz+vUZAFLRpq6MKP+UbEyCT7d4pTqgVprkm7SvGG8DChXWEnV
OjDKn0ivQJirvtP54YJ4TppbAocogZRx+4QNXQS/vif3egxGLbw4M4atGNoxqwan
rA9+S5QzRIqqGhDGQq1SjRov0zfiKzGNL6v3zit+sPq8SrFCQgqhaIm/NluxB1MY
TMGIy4j0yjFbOzEXkkHliqr1uYptE2otF3puW9emMbm8CMaEwfW5l1gP8DI8RpKD
v+gsZwra3sxotbvqhc4gdz6to16KWY2Xb254HeS4q2mL342LVAxQLHtqtxKfZGLO
EfdrxchTGYI4GnoAO4Ev3L+LNBSlAcZYEGQlJvBOT5Du5nvmMSRiir76WWRBLZms
Vd4+el0YET43sp4zHrlcNMtRZ7m9NYLjjkVv9waErQvUBdoCyOill/GpO6m9C2TT
4FwCt1HR+Y3gnNmZRSvlnUhk7lDh7KjmNcrZ1lTeDUjWM91EfyBvi7OyEQW4OcoI
4Qy1VMBC69rXMvSGeSbEv3dCLfm2alOT3rZarDGg7EtrMzrpUGCwVesRov7+eOPA
Rk3aCRXU/5eWOSutEMDONdHFEOKx9l1TYpH5N68RRjg5MaJEkhTjorr7T0VCG1z7
wImh3MoiGeP7SOcLpORBVHO0VuiegGXZuvvwx/n907+Ow/1FNzgobAqnuvscvAH+
KujV/lzmNwPpsYRROFk7C5GbS7+MsvhJT3tzsaPAaHdBLmLymmYAEvabnOhFip2D
KCkbgu2eEUmsNYRb0ebHeN+JPsWSNc0yHxrw+vD/LQn8z02LWWeZXeeVhcLEwF9I
KWWfuSEwA1RrZvF1n3kWTOnxGdoLaq9V6dvMSzHQII094KZ6tGVm7i18l91So1Ih
qmObE4Zl0XaxDe2jmAjJDJyn/Hs+RcYzC0OgT6Uig+JXc59vKl5Bb5ofxwx1kFKb
2e5w8jsIhPggHvRELsUcTyI/PU5YeFV1t4DtsBQwht/y9HhNIQyqnqR6Y8HNLoXf
kPDk/JGQeqGXtGq2qdNqVOlMhNulqrya3yuUIhtynKTHwjcB7WPOKNkpIxltnx9X
zpkBDQgRLHdN+Vze5hjbVKIdqdw6i8lxMYKbIJjAYm8bGWTgsD9hhN5FxvH5dzCA
PqySMCfAchuy+FtFty2yrHWSIGTREir4odWTvsMN7wxzqErGlv21qzGHySxd4hWn
ZLEGsx/emD70DFc9MtSOXe9TjXR1ZxZOE5dcTBuB19PUUNwGFOrIdRQQEQEcAI/m
3UxhnRO1TrTF9OG2RKhCp5TVgPUmr1e/sa/IS2/1j7FXTOKSD0BOPFbzJchP0Q/g
A7CA6sjAjJVk7iyxnlc0pcRjMQPxduBecuQH3L501cbPYiEEpkI6HR54to0sbAxL
35BplWOl5bjxLmA2FIVrdFkhz9wg3JW8BICpO+5WgKAaQ79FAyTtNVvTlse705lz
deM0dLCWyUo6I7xyqk66vgauM3SfOHd59LEofjDrR5PncimvLF81JkTpROu3KuNW
SSq/C7ojVIy6neK7TsWJPyFQoyvE28/Omf6DT8UGHGIi02ISpC8/dyP7dqEN+UEI
MxrbDyQiXjKp/zKl4b4wtteyeXRTw63j4xDzbOoBx1hhdd8vjVHd3meY6jkZiVpj
IICA4JUd9gei5HHOSShya62GScht1ZnWe8dqJP7idpkVRmAJrsN7eD0n9qo4Q8tT
p8HeKeKohGy89mz/znMM31HQp+7xW2PJ1exOiyniN7OARxEbaus/EpgCfo7Or0d2
fneI6JWAVSWqpMLih7yOkeCGzjX5Tvxqb8hWNgaLfDGfJrWO7wR2PJo7beAsj6Gz
zi0sD2TWlfEwUP0QwEgfbtfFDoQFXfGJZgjt0KN+m7YLdCsecWSX8kiIXRfArrdu
DLRqKX+Ore2f/ySPzUntyaCAWZlbwLr75HES5xHaYrkd+YM2Yg+JhRA+uki5vHcZ
ogQzdBWP/HqO0JvrdoaHQar6JcBa8iuKWQFwUma/oeZYcxecl75q8jxrPWsl7HWR
b1/1z6bzkFPPbiZ5nj+LIlE56wsJ06QjgeBK9J8KGOGEJlqwmAUg7Q8HfUvMGK8P
VKOS8CMkPlFDRA33Rjm2ssanJC0WlcpqMnCyI0rMTGd5zbiopf8Z8s/i4fK1fHcK
255wzSTLWPVyhjq1Vxbm5WulBLrQg5+wwvJOmdSTJQaQsREgBF0qhj1xZfi4TK+G
hP38ITZgdCaG2zBbuqPm6cMySu9TpeawDVyls9IBUQZ71qXhiMtvPmwhEPKOaOFV
tGXaKKmU8nfS0LrTPc03Tcz30APg4uGLDkB3kgt7gyMP2zdn1X/cN4iLUXgkMXc6
j321avKtv3wYf5lQ+LcxOeORmFMt3wmI8NIj3glJ3sbld0fwJOyPQuFdOPHO9uvr
MwH0+7J6RWkNk6SXI8L6wyR6W8sK3+Rm+qLuPu5l52H8iNrPzAM1IFDvRQ1a4DTf
A18ckU3qMRedkFFRFCQL9w3gznP9xXG1MNUx47IuJto5+ijj15YUr+yl77s3Fd1m
6alp+ZxBAEyOvTwGfAek8LgOpBEOhO3BX2+xtl5XkI5Ycuax5RTFB+CIJ9Lwa2dH
l/gttrwaziKkCEJ2qUX6eEEL+Gne4SMTNjMo5YxK56dvxzpSUjQnUVcPWpg3EdMU
yLK7ql5Pyw/Uyc41U/BOAdDvitEAp1tn/jfP8m8UTpv9mc4iMj6G/G02a8/6LFmf
ZFhXKq2bekpRoHRHfyDg3dQOs8cn+upn9PjVVd2E1Axi6pS1bUskn5g1hyR7XfOo
/FoBEzl5ul1SV4MoBQrMQY14zwvbEjCEFuVZ0sSRtuVh1M7YWXrq7Z3K4yi+Q4lU
YN9296UyUWK4f9BlWgD0jk92RyXkqY/DWfz5ei5x0/rRgsHRLTZDu4YXzBugdGPY
TdbGVP5oU5AKg2R+InjWijYZLMwwcPIPW+39G0KiQHQHGLAhd1O/ogVZho7j/9bC
zcZr6tC2WidOEDSJqgwHILNt/AkPyrK6Kkr+r/2+Xxb88VDC+HxWl419JbpnNydL
mfjoIjypOWDmZHOEGxtykDI4tv53AWgxBXmFxVYvWRdw6O2W7q51HX3WL8j5kU9A
T16GMJCEUpsZf3HeUyksGPiO/F6sH/jRokxMu/BhobJ7o6lX4G81IXb//7Hys441
du+QIPE6qLL9VlQXYZp8jE/XJFUAAI5WzHI2QufZcWwPwsik0hFiezj+tXuIteb8
g+ugEtWqtSvFOspR4HMJk7eV85BxeY4u8qIfcoVXMXFxxdisjYmaO83eIN6QiqGw
0yNn/AKjtUtJDTXwlIua1FbhqreEWVYIIuULw7UbcclUpVJTraGbDz9s/RJEs2uQ
Jfc4wrGd+oeAYGncUdlJsdZBmUYKZbmzv9+ReMnybktvOSSCGtvErYIopGJ87FxZ
SsK9chgDMffIbf0ReNfYX/xnxnYvvj7gT0FmOYE9Ia98ymRNjtnNZ6Ku79ujGP4y
XQMCuwvEp8hyGkxUka0aNDkfTSvpJ7Y/v3BjwaLp9fimlJIp1oP1jvR1qvWsXF+M
Vx1Nl8uwgNKRPEIj3fLNzUFaHJSeW+Sl03q8MSkq42q9Ofe+kRo/GcP2Or4C+jDS
CrlHIuvq8z4mIy4mUYbXhDc2BRKBJNOpqaPr5ume6r+wBekuYI3iAh/22q9FnxFh
3mGNs9jBtToCggcOSSYNM0k1Mq+EqVsR4BNEov2VzDIlBG6KFbx6VG0da8fd41EU
dLMZIFhF9FHz7V4OOylRZ9+E4rZ1EQkgF508II43Uap3MUbY6c5mch3jM7HwLjDU
CR4orx+HGXiYNkCDNzeGW0EJDl1K8StOa84AE9K3J4UQ+SmClutM4ORLk9uF+/gx
MX1l1ABqeAK12ah5fsr5c3goUVpUKb0YlPfVesW0I/iNTqyw00ol4oNSWyeGmk11
RxZ4vZhcegaCnUGaN1Qn4Z0tNINH6sL4IN9EGyrYGc+AfTBFHjplq23DSQY1fo42
CEsvy530RxwAeSn6SCr1V4XuEnyCNhfB/cSYS3Ad8PJZH43fN0LaXgU1rtxv9zs/
Idzrf8nKkTg4jUtrOhvcHRJNeA1KiorkFonVJBW4YI28GGS1RDZR26AyDV3PB/Oq
ug52/C9rpePuRLK+1amlbnjIxdsTFehKvSV+tLWSlr2jOUIyDcVyhHV4aKYeHXXV
GmkgzBCONm6xNaj+m/8GXj0m0rNOYs28gHT+xZ+IQiZOZQwV8uCPkklfGrA+tXLc
I5+SuYL3WO18Crr+gYpe96ACR7HS+q8+exEYlAMBG7/m1dElXEbCj5ttdclJ1zDf
qH+8RSDnvq3E8aQ0GDwTZ5ifwD4m32KwXgK1JvKkjsbEp4286Tzz6kxln8BUJ3XW
hgKW/iW0Fy74zKskILm1cIlYgX1SBMM+ANYrR6kg9+pS4EUyM/jAES1W/dHShjGb
7swe1fcP2QLUpA3buy5WiIFr16lH5D9wCE7o27kZiVospjrwxfVKv9nWo1b2b3iN
GtTGXnEnJrfE+eGEFY72tuDU5vkSaGgBdspNB/XTSbh8DL5XUINcOIIdf7zQF8VW
ZQ86Bq2jbWJjXabels65x3e1Djz9WWi3bNXbXPJLdIZztVcU3KhJ1cceIq57N5Ed
QwyH7tyL06pq/FaNyPyYStmylVSqifXJ3n/WYv5jQpOFBPHN7EngocJHut3BgcGv
jAB666kYa98ulJYO0GcPKUNT6ufOiMWnlFcJxtE3qffxzqloxDoLqqkUPi9mMOB0
hdNOy8/cmwiBPffZIkRsRl0qYrJcei5QAWwSTVuQQ+k5jkhdFoGhvqtJznd+x5pR
+4XokltzFVdzFx+9lmSImlmMhCkNJ6Dsk2enwDLpxvEXUtKLz9lnmmdgEYZN5kbw
mhCzrKPgZMnMnbTpZAde+LhuC1D+8sgfcNvPhj6NI93hTe9PPx4Ii+C50nLBg19v
+Z8F5IVBfvmdAXGVfMUVQe+xiw20FNTDI5pXI7Ska9+6atKcBQn9MPtjB05lzWFb
VwBADzgtS75hMAofLokO9spQ25irXANgsq6ZTGrB0eidOKWNAlcwCBn/5aB4sZYO
rjpZIoEaXlqBlmT/DmS2+JalhZNxl8vOQtGK+0DA8c6oVjHbooUCBDg2EjAmqj80
PwjQgRazn9lRNB7a3feYXjoZXSfkJqNDAKezCr2/gcWogFtWNcKD3rUywM8EnXJG
jPL4igPspSvmAPt41fuWiLksCuMOxbjK+lnlTvmZc/CVhWBJRPohxquJbatzxPve
iPE/1d56XsJtd9OdXlhsxke0g9KdrqcEaUW1jwRDtIJEBN73KrK9wMJ5wMuFwo4X
+2KqiFplXvgoYH9S4zKTps+ePRLs1zl7yfTjf2MtGEK1yq4CvzN0DH5R9XBBe/PO
ADbKSWYKHn/Z9n7pZAtCE4Aeb9y5M3PEULG92JWEVdtYPvB0SBwRKAOcWgFuuPG/
FIpkxQT18phwF8aABAHjQOTnaHViHYWmVvPs1uc+yJkpiLCTh5lpi+Jf9ZGG63OO
Han8r1NLgz8iD+j6oDRxuMmhO+J9Mm+5mwxWdAyKHECdzd3qbvNv9i+Asa4fIYWV
rZPGvUmj+xh2PwKBb/rc31vs84Cf8gdxikrjnuHnN1W9lxilJHkxK05wyE+YnFlL
4mUX7VROwxGbW0QH+CeC6fefSo6kwuw0c6xMorYY+WitpFOEhkcx8R1vHVydQzN0
gsFc6h3nf73i2mi4Mg768W3SkmBIQTtuOazSH565q1NO1VlkVfiFfDBil2AcYrpF
CNDrxFFmUs0/IaIZJqtyfCHFyynFxw0KNellHTiHQU3kY788LAJQadsyoI96dGFJ
/MLNrf9T0EuLBTd20zwK1IGlwcecFCOM1ahDZq3Vjd1VvxU2GyhRf72gS/D5eRzI
w6t3V1twQ/b7sspBS3nOy0J33zlLUHQ+WpILXvJ2U6p9uWtDO/AcBHzz5Pl8rkwh
nJsBYlAHN+mCmMrbLGqlgWsStB1x1wwz61UUw6WuXZ41BXUJjrwDm7bwvhreMEGQ
joBgCNOc5oRHiT9Sb6DduwWQzuG01CEWT8Cq8SG0B8uBKmNqHrhVqMoVZTrH3dOo
z81DFxDNgNniJGiv/RlwJvtixUb//qH6v+vKTp7wI3TyOmZMf5DR6TaMuk+fJx3V
rASwd4Jk7MO9iT/5Svz6J6lo1TDiBVUfGORk6BXLjExW5FSptEMgENLGWrMzdKun
MUCbVVW85GGzBNfleDzxv11Upkh+BYoqTRpYUUYdFa+YHAVGGcZglhRjBrIx5VAu
v2htfYq+ZfWgcJGxYetZNCKKtQ01znP6aJLlKm1+B0xtCUDfCwtxLeZyu+WnBRiQ
PI1eagTN5I25ka1CZ9sC8kVLUHBpAPVIMJ3V83ew5x1x1+d7VVNIsiGm+cjeDELs
/Nw8o+r+/k4LNQwkIN5oCUZB7So89/QDauLoweG1FxudP4XqTfaMbZzYV35I7gbG
aGiOVeaQq2ImCYh+V0/LibWQtaNYp18dtounFsfZNC9qhRhsTQwtgbmq6+jvwNzf
es1QTz9guUxxUKomzMOtseYVPcrAM8fMYUKFMRmx0cIVNfIQzz2d8Dy9y6ur2Eif
0TgqKmNwFhFPeASlvLVAH9IyXNIU29jz5daL8FgqI42dxZ9E9Zq9nB1YkjWWNhju
rDFm1nkBjmPyXghabi78bsYU5cF6DvyWHdWmwZ9oE8tB8EX1P00n0E4fViI2RjuE
HP5drXyGKiPPT692doHgf7ca2KzLtuufNSfyuSWXw70SaApqQ4vgcpshvqdDhFPK
kBdBefnWGXUtKkSn9lxaTK9u3qm1cKp2qKWLfFOaFZ5quOth+RlEJWp2DICGSdPG
YVkgWa7dfHPHUvw5jK37jMQzhL/OgEog2Sw2aYo7vJ5F4vCZykn19291NSP8qYAE
iTTPxciGZCNGYcbUeVhuynQYu1e1nMXV/qZgnsIFeUzY03H9v4RCjKg/B0/bIh0h
nMg4rnznMa8Gj7b+93Zde5dtcvAz4sHmlxbGJXSW8sTcIj4m6aHlJf58vFZG9aBI
Hqw8dPVzmiBWUsmyhKmZZMFwnDR7VvyKMNd4WIw1SgaCRiOEFErSu/S29ca0oeQN
RTavSaGz2mAef0raImsJhAu+xlwjoqa3ema7Ga6Zoa3IXU7LpAQCMr8BmChv9deU
4r8hFRNUAs+Mx/ItgZqS2uDjl37CRmG/oHUSSIRPEgsayQMnHggUKpdHXMAsSoUo
B0IyUeO7JMqXJH4rX3Vy4ErurpiPyzqZLb83MuUbaLZmCUhpEVikukVnSV/1iOmS
ZmpaJ7PWtiLV6ufiUluFUtvEhIvtZIjWHFngux2jW5MYcbibdF4sk7BClKoP39Lr
tPZ8godFUBPvk4DQVAyOqzm1uc4Sei9VVpvXP/OuxQjU520q+F9vEjdAlgCr1YNA
Do53BQfXmZ6qQzSj2DuhhxxHcc9q2US8HZrnMg3noi0gHgds/IetrmE/akiJ/KMi
fVrh+Pn1AxlnfZhXANORkttSKP+gFCcN1bP7dyXeqnce5NXxYVgCseaM3TCm3Jqs
46nu2TWI5mg1ckYgQUTHUydbkh6FB3UyNQJjZEpnW+Xpe24HjBDSpSGbx+YKN9Xr
0+mYuxTpqwPzz1DPKu7O9JdJp9n4K/oEjfOVJ7/AT3s7xPZUNveXZFrKpo3BSwsF
fnqeOx32AINKjsxBIbmx2zgQ0MgqJQn071IF8yEfTgJUfskg593lxOYG6twVqfrX
eEvneAC33btKYYMb6JkOQoQZ0UM6egsW7R/1znH/dCcVhAF2fHNXUXRoHKBhPrTg
d+mVjochGvEWrvSnUauAQDMApa4LQpWlJDY7uV+GZmggoNgoy/wI54MDnxNiPPJU
8zW2/QVsTM4dAMaMzck+QJshVwI0pASU9pY3jqlUxnulQKCj4BWQn3nfFGcOKXxI
vAnyFdcOwIyCoWsIPzdE1hqums7FsEPVQ6CLvdM+PaMZ6P4/F26QtFo35edYbyWl
TNdxCkyhPC0LR7m0/+kx09oz6BWuv7uZn2+EO2gEx1elSsfnYzPX4FgKFLERMT7d
sD7FSeqpHaC4r4sgQCTn5Zm5qnUWsD8yHSQ/Rhe667tcwSZOfJOruSven5lJTg3n
ghidmYvJKhPwYPqSGim+4my13qZQLdJoOsyY0TiLnaydLzOwVKdHEAKpZhsbe9CC
IUe5LoUCiAuPuTny1POpKdbSjGYj8lH3jwvmahbx9T43G9tf/BkRF+dZB3I1QqkI
WLt2Fb/iNpbYJpo47MBW9nVHBoS1jxGQJT4h1dsGX9+TEUXXSWNuK0NCoMcnGzUd
7Z8TwU1tyRzxijAXZPCECi5yc5I/fIrLENZRE8y+IXmtwvz5QZK+uk8xeyhDZbm8
jGfDDtnhdqhiYqIPh0TOvFI+WY4nie6VB9Xe3OgT/3a6BjfSaBr+4U6NIaRhyBHz
ZaE9iHqEITglvZQmRsjtMzaCSDcygk6fMyCRfNzBOHwvtLWnm5QabzZslkiwNSAC
II4Y2VfAvcYZgQn0OflCFFRt3bD3gJ/I5uNeDiu87MRMfHUDfjqQZPrTzyzfSUku
upseZ1WI7kvIGn2PtCJzjCKb/s6wDDF+lDrsY2jVuAx9xEukNq054P+1Z1czFlWT
m4Awz9HP1q86kRSM4TlwjWYrExuGia/jcN1RsIjhs7SqpV1ASy9cf97lxFyRa4Qn
/LyAYrT27lO+/kNMs8UHCdqUHVtPM2o0VgRr0kbh3xPwNaldny3z7ATkd2ujF7JA
9IjaYCR4LnFXzCr2Kc2qfpdZsp9OMNP0As1TdKT1ho9UONb21utq/jK8bld7s7Q8
MPaAfk2gZdbhkSZNEt6u/Mpgfzg2psg+0M2Sl8/MtBX67d3MDlP6c/iXHXGfynvS
py3VGMGHtAG+XgCd2D+DHrA5l4xlgJ+j7/eiLfCCpnq7HBJ3GFYwPLd3g/giKAVo
BfrKipJodOZHfLfX0rsZS0/qI5GG95kgCi3iru1wHX3E/i+67mhui39rz2peT9oo
3cyL1kzhbp8YD5bG7NOXnoKb3vruBhM63yL7DjUtZ5MuqfU5+SugTsXTn5nQY2cU
dPWyvIdacSlF0Cu40A1wAkWLp3OJXOKEQtd/MgaLLvC+dq+eoHoofWGlvIXgZjnZ
H6SdKOyXo9hCWrgysY6PrI2YFuBrZFoa17ble/GoE7IJ0EeTHcMfRgx3+Z59+fdc
chgbS9PQ3RssSuwTkZZEFyfIoQWeO2NbgCGc5fsbud82DVBH1JD8NzEpEbFkH4zK
aHNi+82iU7WETDEzZi+yWRf7dpMDdqbC6yiWpufXpcGkFiUmc5hwrDMGl79dhvuR
NAMnJEmG2r8aLZKBtN6+2Bv0emAPrX08eLrgRjMNrmrOTn5RTBggrz+Sp5eWRd16
G+0q7VQly8/WRJIsyTFKkLmeO1kUR40Q1O6rjhloeOnYB8pA4fRElilQijOlbi49
tKQGUQwLLkb2EsMIpqJIQkJPzxAf/8s8zvWgctvVcQn+GTX1FKsRg7hdTZIIXqU6
OJex+nflx7Kxe1QxiU8cmmlscSFe8OkexxE8Dncbzo0117e3CTjX84bpK2JV7GLE
xLLjvmL9W+1crodl7bTxcVY9oZkrWKserHJwix4EBvlsEgLnLKhObw/zHqHzjTjo
cbWnUqbUj9wHHG7zS259nh/XnXanA2tneBaHLi5d1rwQ+9zUPGxokWZ7+gkhcOUG
Q5kwZsYqHYg+ZMdhOCdQwXsj/thwWan6CMUdPH17PbbT5eQTFtuAboEZbw51wwCz
gOYoxE9cLnrm1WcFVA6mj8N9xHknCxLfhiSVCvQXdxSkwbU+lr1+WRtFi/DnU0WA
EC3zP+BFtBq7+pNahNv41H9VPyCR0+oRmoCeXqQwGDWtothI933zJMd/RuTTLriY
Ko0f6To4mC+2XK1QT7KZaeH2er7cVKw+EJO48rs37tANnpszyJjUzetRYld3m33m
A3bhl9kSMmU5cThGd2VhKO1hezZ2gMcayosQ2ZV8Nl7qkDuFv6bq9xmrhJc63Mj6
o4A+j1xw3DkE33Of7AC20tRHcQ/h7RKqplXcjwcg1wQxDBZS0jd5dXeqmJpPZZDk
MTr8Ezuexwi4xSF/lwSDm6Y9TrYgItFgnJOgNNaczHI4s7Hov672/RiaNHgE20lF
o9wrjn/maN071+VVcDT1KixyIcN/g0vBmCgmJYd5o9YOiNTFlayXqvYkomsdlipO
cY1OVMRReBafSk7iyngI2FwvdTUn21JDGeFHKdMmQS3VFAulGC+tf5MblyY4L+Is
cRP+8JnAMPVH/ZJKczd+H3f+Hbpz0HmrcFmaBeJkO66mVxUj+q50rbjjUmwe5Yia
umZI4leazh28eKHNCoFNUkX74l0/hprkT72n6+u+zi1Lc1W5JIKSDhRUpoj11Bdi
RzVZUC9FVEb0CGvqSLLbUWbCb9KR0xjaiPB1x2vsR3tnTJAYNbj+0/smXAiIz91f
QyCI+JDonl4F0cSQMR2kIMsp9N6TwmSR9+i1Q0hM1TDOP1LjSw6R5ol73i+kysNC
jFQ3pucNBaOLeZuHcIXDL59PZsNfWDIEQhdssOxlfWbTZZFfhy9Ib1tq3EX1OFtJ
Uumy11v77gA+OOr7o4KqoIhDKrAF+gyqNhkMofMH3mOPHhrXGOdeOmN0Qv5sIBVN
6DEz/1JTrFhKe6Z1bp8PpVKwunJAQycMgFHPQwAO5uuLdrLmihaFmhKRI1kJvIju
4A+9oHOWoHpEgErC6xSqS5U5WaXmdnCtNvSyaBxtdNqYPbyDHLtV5gHBKYTJmQIi
TaQMgJPXz2eX9j5pv39CxpI6X9X6mVEmMokpL8Creq8sz3WJtLM56V8bA/1cjqaO
/8xNA7oFhFy2oDCfk2YPXWRrogr3EH3slzMTuQNjR/cxWdhQ9NMK4I56FZzaB3Tw
VIn5M1ifBpOisot7yYwaGWYP6Fum0s9DqWH3Iu1OR3lCWq0j4BpMV2GN1n6B781P
LVqgW3ambSnLhxk0O2+G2j3wJ5Flfy2C3P2ytTKQmz8zI4bC8MDriIzSRrAW2q4/
DRxaY9D89gM5C62LVxXkdZefDgcNq889ibjDpjaR1fL33QjnmeahlGNgP1KaksnA
W6AmpldQ9rIGgtTlQoQedcPs5KC0UxLCVdV2CpKy5pJA4T2aRQrkN/NBF9l1WnW3
7MaZtIjJ01mToe4Azc1S97F472c1kL6DJzD/Rt54aXeWLsxFpSatMwr2V5a4RbZJ
5z1DYZ5RUAtlNdWI5b7bvkQ7/x2zhsfRGPUC00dpbbxE2gwB3QcyPukba+dYTx2g
ftearPCYqhEO5smvtZKvXEDALZ8lszjRVDRXvvbUdYQiPn4epfXRuvnH3ZB8kpKO
vu4Qq+mUINDx9CN1z0Ije7bBeWQqrEs3Ohb5VCmu1CO0ZsjqgdrEfYoZnJfPX1hn
Y9ewseRov8F/0100cPbj/WiNXOxi7S0eQnn5ZU2AYOwu2mR2Tb1TAfXYgsbl8vyC
Q6FRWWYR9E1XOiW79HltdpjbWYXplNbiIktkYIIsyC1QI2x95TG4mmI69f6qymus
Dx1gXx3J8KoP1EFh9IvuinqCjzmpl2cxo+L9PhNKCkpuJC+l8l2CLsxQIV5rmQeA
nd07hzvuTQxvSnxDCbMVrKXN/8WVEHjkQWWPbBEWNGetRgTuNLpgwRb+HSWH6nW+
aKavpHAP/ELMrokEZv0fe7E82+Us6Y7jS9MSqRUXW7qJE0qoT5A/ot3TimYLVlli
Zfux7CCadB57ropWqwXYDtlJKOPmrpmpzkRm549NiFEKFi7OAVd9uDy7NOYdcEwJ
nz+rP5BdQJWHyetfWRPZf+Ey2onToIOSRnpvAbnS833+MuSWfUq1l6bfQnUipczI
IenVCes0jtVgz064dmX/7tkuw6b3RsVUKF4ytvXfibJQhzH5VeZj7u5MYWHaZRii
SapDiAZi3BUTcUedPNefJSZVT1tYB1z2dyqtPi/C3w0FYe7VbtpniDWh6a9mEM3L
Uv8cKIO0C9kchZm+v4pYM4qA3gqP3Jo+08ZhDNndBt/vDZKsWmPHiy3G87ZD3Ftt
zW0RcD5qxRPALelcQS4Lal0d9IuTif6babGegGCQa3BjvwANDNBUfU1CXRA4PsOQ
5rRW61TqK7eKbAR4i55zPmC/LDkizOTisFuArsO8QGRQM+0cs4lY5olWfpXAhFi/
MhpfPNPiQsyQHT/0G5KkwgV/z6n1Shk/kP2ZP3EHhu0NfR1H+ti1jrQBfdQxo6NN
KQXEC2lXr48LMXokxKkBfilySVhSdr3jAKayb8L4IuAMc7pe5RKJrGwN1WTed4EJ
lrqwWiFyWMGWOXKdA9ZTmIwpd2kW1aGL9yyOlq9wHZBtIBbh0jmRJs6OfCwlC3ab
NaXupc1bAuZZFCX8QqSbWuvERcxNxGmz/5jUKud7U+v4LzeAw7ebrXlMNCwPW3tQ
IyK3anAN24Lk98xtHjnN4VItJQKRk8GdlFu6HmrozTkhyB2QWzRtsaWcymqmZYZO
SsutRUGeZethnTUazgyd3r93HonQ5aNeWgZg5URuWYSRSSVgSiWSSmoiNIYoZMY9
1r3ZYjq4+PBQ+prgRFk/xwwjLPgIgIeJiNiMr9Y5Hhb9xJnrzHoy4+iJO/czLc5U
Qk6Ef0cBlthUejoHK4eSmYxuWaorV8HlyZNBhkpGdnXEqf8GFrIQvrXFnZ0b8gmH
nG58U3ubT2XhoQ5ToZseHCM9zpQKrGdnS6hPj7JaPFuHuvYMhdQNDAwQtJgsQ5kW
SRoBWnXS/SJHVLfaS5YumHBFEEjfgUE+9Zajpn0ugRpvufCUs6hsZ13iHQYZ+u/L
umqg17CeXnBgyEmGFedx1Os7wy36Syx8aqCJtrhrBSO0e7wVxWJf/sTn2B3uYeSq
FV496A6MpMvbWfpdoM8erwEwzKaKmtOwWOs2SYTjRJYqk2Hn23C1bEiYi/AEUCOL
rs5b0sasOodmfU0678TF9AIMYTpktsgI/tC7M6RBaBoaempMBptofEdNlADZmCt8
iW2pnlNtxCXv/DSWqymRDUDSqaxxf271JQExLSzo/tbcid64P6qI8GOHUtHIkGZQ
r5JXHH7ZHoZaAP+/iYEV5SMkUeQ1g7+rAFuCmZrfwZ25J/+klypuXSOfAGQXAHB0
UL5hJGGsCG6WmjrmKaqkKrGbpc+bKTBmllOYCH1vasO1wPzfNcvIYhoyZyKm4ZRR
Z1GicrB2EXC/hLSciR0eqos+AGk5Z4PjHEjRtHpPS5KzNfjFhLbrzfPDYyVCgTfN
lus6uvo+lo/JRzQzoBQgM/edWQmK9t4iu01OxDXgKUINChGEHwlWVMiMnLaixruu
YJUTCozB7Z8XY9JCp479ZCtTmhw35mu9kQPn6ZFf48/BUBqHRoqI3sNfH9FjgPZ1
lzia3idkNxGdimfRAFlDMCvJ3dpmJkPH5i+yQPNvaIer+hr5YZGJE13vzXILXDDw
n/UChyymEZj6Obg2k6YVS8E5OPAyrjUdy0YOQ3HqLhLlZGa3k6zyMSWUKav5vfeg
1EerN/V9Xd1QnmPdmK9EqQLX9DBA9/cu20TgpPyJQKp4UZgaKmWH5fV3dJpwaZgf
CWHT7AOXq+4qdcsipn08obg9nY4XbXntLdeViClDYehUp3uZ14czmwCVgVR++A5p
gTh4huxBi1z/1tIFhpsmvHZ8VKRHfBGWGuW1NZWiIyzfN/EpMOl3Oj8F9TvjgKpO
cbASZJGpBzg1V/JGGfmR9G3LUqvBBx1W6mc0ttzWO+dV+TYT9dI/Zy4x7yWwpoyY
I1Lq7VgWExUolvM5FpzAljHINtbElsMAktmsc4cbnalEyjBhwHJsqcpYB3boCz3y
wVlJi4Sbh5QT9W0gVKEYB7mn34BnOwZVUjyXtynZzGxDdzE/JkqzI/qLVSmpGuat
vB7++GFb1RYHP2BYf9FCY93X82IZswj2ENIQmECjaM2jiBgYAeazQD8LTzMmrko6
obpu0n/WKeWD3zgHA6vlxIcUMSIIHVVNu+1h5XbFJCxmd8gRG6xc6/ZppVhBBLV9
t3WAhAHq7iOiq+VFjjTG+m/6T2xRB6m/h9IRwSzgJcgShNYZ6cc/PLKpB+XdkG6e
CGYl6ApNsV4jBHLxBr0nUlDXw/xWhZCJcoHvNOrUGD2N5bcqiBKkzpC2/i3WwvQg
kR/4SCWOOllpidOGOWyeYk+N8NN6Ge3I5EKf1NK0Xels6VjAkw2ubcREx5qEno6w
U7vAdpyoVXBVamBplXVDNDTHvvxdtohH+dbOcjyxMjaWh+TyYPKliFv/GQBgxtLr
ZlmFqdq1OvY2HJ0zYjyMNGnhlj0sfDPnUgoztfmWdeH9wqZF2Ltr+ig1Ws2W1UhE
sMp0q2P2qiJL3uIDj8/W3inpLs1ZUFfnSNsczAxPpr/OzYu7wSMfXWWwlam3yf/3
fyo/EWcy+KoTJzpTjNj2EXTDeruluZ0VmPZGPm5TYVQIGVDpdwTHLal911FmwD4w
Y3yuNBHH4tWruEZP3OLA3yUBl2cb7BJ+qFRHn1fU7Qmpf6U/hFZKkaqBuGhJndl/
+gCkKWmKF+pUaTy1lUvJcRSITkitUm4Y0sffmZ/drxTfKA8itlTIcwUsyXPRTCUX
VBKxa9h09BzWvXyqSiNuDjXhi6OdRTl+K32UJ2JSWApPPFbigtoTp1qXtQKD10WD
J8hWIYDV5l9I0VbLTx6TFEgHAFiFqnpkxumAkPGbSxSTC20uLxWozPp58OQK1G9p
01zoZVaCdxr3fyaGlBVQl8MpfWNHRSSnXl5d/bug6d+63sWuA1sh9uVRlWEJTekp
LC9OgNttiQidpMAwxE24F8Qi7coTl7U9v/xDhIgChiTXiTi2+6iUKsO1XKLvKuoJ
3/Av5bmckh7xbXE8JVg8auaDgnOxO8YC2iNS+xuXHtOfxDfdrhM+R+1Ib0fgy0zp
W9WLelIdSPWzh4vwaTVVURH4XaCJBhZVXmpAF5TUeMcasLaFwWHZzMsue74NyMm/
qwDSK62mAzFvh3CMbd3lyn8wmPf+ujCZ3GMNb5KDtBPeKzrSdGOOi/BisjsIzhgd
prGwUqEfhjWfaGD2BMgRKdc4StgL+UItAi9MOXOfCqVwwx1HEzEZuL4b4D+jVds5
VaYDDAehWBcjNawzGyBaQp24+InrmUBp88XQi7ayYUY49NJOdITtTzEzsH83HPIS
lMTsDBuT3uNJCQKPeBAPmUMGXycxEW6dQK8DkwVVqLH4DEbZY0vjSU7qlEKK4WfP
jKScqE/31HFyIxkZ2MyQmwy/AOfTf30+VTnF7sWdDFysJvRCJDo4TjLk7baLHNFp
omyV/Jew3z2Yil15jzH+lXbd5AylRXApvjHayMMt2ouXGbLQ6XQH4hr7ufCc/nyf
jga3oetPV3CqsjmX8uIjZa8PJuvwt27snO8t8La9v9vQE5wPoEcPqHWumK4+qXXp
vRncIXVdfm+C+xbikiJZ1G3XzGVtj0lb/HaPv02/HRbV81dK3/sYa7gErUkcpjsb
BqA5c7Cim1QPSqnWjVWTeLPXQZyBwaHOLlocup6HZkBmWLI9/V7ZYD1SmJhUHkif
iq3mm6kEZQyKWQux3qGay4W6u60POuzPpRbcfzyyHxqQupkvbheu8QfrhR58PuKO
+0GKE8Kek3kM7PAu2GdJUOx8c49YDv3L7Jx3SCYgRCCACs0UH6OvaPJBrb/UwzqH
VFXaXaMi+rM1IicV1x+rTgK8vCvYtRlaqeHU9wlDpYPGwhf61tApODD6OEqnnr+I
l2FFW8HIsmh99FAvlkU199mKbH6n6DBXRiLhoA6Whiih0B1AujH99yJAgQWhGQo9
1srz+z5kbnPBpioYEh/Uax0n+t7yqq9vwtVBraAm+Zz1nasK8zQ0MY1fAumbOUz+
WkEM2+zsZLD9DJF9rB6Uo1PDJQKaqxqbyqIrW8setwKBo2H2jwcWhClSPhCGWNKh
8940pvtaz5K3pv1N+luW0FXV10IoBk5vDyYQQ8W+kQhPB4SJsnSiuE6pE/HcHFfF
9jP8TrMoSw6/b9PjXoKcGfNgZ7T9oepwn6X23JPD4t4tTZ7EcQ6uM8L3FodJ1q96
olfn6iEQXJOk3baWGDIXu/VDiOR7dKZL/r+qd03ChwPM9Wd0a7afYD8aMBMaOax1
jq6gdpA8F3hpAzr/VVxdBj5ZMCkTqgQjX+piH8UX6MLwPEOKLQvWVfq8axgYzQne
9QHQKR0vXBr7XvIJT2iaBE6wbEzHfzvN8h/VV2ya4EOAHEeCna7gVGsYNnLBvz6j
0XQhmt49+Mk8tqCPIW0q28oqajFkzjiwp3FEj0Ita4zzefOq6sXfUL3jGEUV+toK
/EUtw4gH8YcNWF8eiPJwhSuLcWk0trO371LlB6/YUykIZ3LNAfKcWhJ51ulISWGI
EcY6ZKffRIH87gMW6gyRs7U3B/uvjIYqQzxF5VRyIGaOdtoZlRNB8UjcOtTZwrG3
TFhs2SqBtig0D8hvGiCEnhYU/f58MwVB3AMTQODvTMmMBUONE01h/16xN5KnztJg
doN/K8JGz2MZsMQ0W1ZcNFk7m2bcn9JYFMtlPZlZCdjrfKr8iy99vW4HzryWRXuE
qxvGNw2DirUQQG1XAfs9suXynpINxCNo/W718LBRQ8LJyiQ1R51jNw/ZVGkEG6Ux
yTKuk2AebFvhxe/29/L0QZbM8EsjWcd7YE2uWVLNm/VE9JKr8DnWrTKpXVJZ8BnC
2V11Ga184wkK68/cmA6AfyyP2Tu5tvqSX3bO4Y5CGuExhjptnyPMjkCyQpjcMvCr
I6RyX7NhYWe5x0hzmOcUku3iaSQAx7HNaXteprpbd/pjZONonGUAbX8ibHF3ZGgM
wVVWazSikxGaRb6zJkP7rADGaCjY300iHfTAtaAGGwAKPl4Yz7po3D5oYhxmUQ9y
rpfGKI2g8c+5hqa8i7TqQXXiyzkigRnIjkE2xXA0iL+nnvKaBHYHmHXQM6xW0zR7
Qdb8QDwFlsGMsrQyYlbTdNvNbwFsaO10l1u4QNGh/R48GRDGXorNBoFX9MYSNl+2
l8jQljGzqI72BsrRDJttVmk66L+WDoYu9vz7kXIgyzhZDo/T22bUobRaVd6ktfwe
J/GXfNLX+p/9cmfrxsdGLca3Ml5uhLTUgfd9MyfZDeSuyyXR/pdkBeI/TdMwg36j
Oj/Z5unfjs7sK6qjUYrOQ9J9e8v18zNLRo+RMlZx3x47TAxuTabDFecNdex55uL7
KPgOZhBEgYlTiwzsnPwr0oALoiKeRwv8AoQgvflo15QgqTh6xs5P0FGUkuBdLe0G
HaTEywXgaLUho6j9hdhA4LZxSSDG72lqSIwMNYveLciY8wC4XAtzNnz744//VTF2
4d7O82wS5EPwasgI/GcNF3eWerjoyrjOFaT2skp/xDQ1CwTy4iEIWf5X4cx8M63t
hhiAP5eOOt5skxgwrnoYEB7fpIp8rngxjdvY3RDoFZ6VKSv75n0cNYbuF1CiSwxW
LfCavll/tV0VL7wV6jgNhVcO0PeTm1s1542RSDCIsNemWQffZ/YyVNH/3bUB57EN
G49XRmd8ErxZc4+8AOPcx2rUQrjmkHJ/Gk6F8Q2Q+6LII8SNbd+v/6RPQwuHSHqU
dxrPgcq1z2souQ3Cy/kbnAkshhMVDIUHWaT3uoMoyN82oyeepTlRKN+Y5VlneoY/
3h6XZ7B+Za1YLwTMYzJA3YNGdxWHpH5aHqIt6x7r1igPrJjpRB6CdMoHfWxJ5S6z
G7TQ2FUTLjzkcOmdR0HNg6vNcJtqp7Lm3v+IJ6fwk4DJ7T1PZV/QM8e2k21P3eeu
KznYQFBg8oH1n+xoXmbJBTiJHG7jS0LtLVV7p0bJ+fiwI5JzaRgYSd8/LrEPAGle
3XriHik3pIydv+/J1N5g5CEgDV6oyKKZeyPVKGdNih3gYpDPq9bY6cmOC9KCSLNL
7QLGgRvwmbTeLGjj8uRi2a314KZYwpo0pt+35/OHsMxEuAdeu3M0NG/fr66rnwcq
swpUj5RWBf3gZ4URj1qVy7vxEwE+c8opyXovnELDQjjhypdTDAWdUHDOYWWfPI7D
G4pk83OSJGBFsECHNVP9K5zHyszdfJjB6BNNUL332RFKmGqlHXz9gQns5MztOBUo
mPWDzMs6yk7uNY913mY2CHXh+vqOxNvuLU8Tdw+YxRJ3I9eegwHH1MbW2DTHGmm4
iYdor9HTpbXSvx4GVU5nZo2IJvCmYw31NdWYuDtwPDhCTgTCap5Wq8THvo3LPmud
Yl5xAaj5mmO5Ja6vL6jrSBMXnIVo0dBkZcjWZqZV2njuYxFlUyDrnzT9r9vHuSLN
/sgBSU82QugqXYw0OiqduX6d9v+jgwy4KY9OTDN2WBA+KrgkhQHKA6ubyVslCeqA
0GYLZiCfU+1Wb5Sfi+XdWnUVwPQKnklKkooqGg3RSYZNGzt4+HSW87jgPKbB3+wP
bLhgZLGW+s4nhreYlX/B5x1Xfzj3QvwovsThtpDNPc3/HM3PCRWv4V3+GmIZNlRj
BQMPYMz/gQD0S7o6RRHHJ5NPQkRAeHkjkyymeKtwszZXXoqd8u2EE9mUo+Sl+JRd
ZdzagugDedwwcitlA/RgwD8fPnHZGlvYOcSktu2GurK7cRfW+Gy0jZwvbCeQiVVa
35qGresAfGRye+xZwa31BHLtrJJh8vkD21H7n7IdYoQNFpvG2u0xygBeGNjm9/bu
76oXXgaP4ciQNVHOnVQfc+msq5QZjw4m1w1MJtoPWpUc3SAUpOlWP95ZqG4PWqIn
5sPSyQpUAdTNJSpeFmX6PpHFB40y6RvewAdbip1P06D5cRxD5AKvnKVT7QWgTHTT
GzI0izT5u5aLeh4mLrTR6APe0UruFrXI7qwMnA4d4GJQasdWVdtVYuzNpp1w+P8X
+RPv9AMl9I8DY1gZtArqA1MHNdbzxFH8Yt9RskAOVyS28QPNMsHq7oXttFLD70VZ
Vh4E9JZ8e8FAQ1eMIrX1qpAvqaSk87+UNNENUHD34lbDPo4YjW2MtQbL3Zw1z2XT
eY8rFTG8jmYg67Jfdz8DXeWDnS8yfrQBKev9QjtYNwQUzcWB14D6VsxiBCSBAN9s
MkCNz0GUhIj+/HieLC3z53KfFF9hAws8aIJGiku/qkxCV1dTcZa5Olx654tFabPH
GDmjqBOuoBGC4xCndivZLkoIn8pMSwcWZtDtT9qDMEtZTG2eiP5PwnGP+rR/ZC1N
XoiopxdYwBP/ZIfCt+y3GIuPIzDnqKAQXmiC4cQEChnAujDCjMFwhXi1vuz3QHkd
IfqOrKQ2f0Dw1MkFNWozN28mRpBuBZH2VgzKWMVWfoTwOr7qhGppPzw5hjifsPCW
OhJYg5mP8idg+CUWJ6PEBtDgIo4I/VvQXWj0NHnXyCy5EMR3u/5zleTcMnpONLgy
Mj2rO2fzTGwAIz4ilTXpAcHZpZVh4cTwWboJfHjFicDsHVR+m/YKa2oj0hv/0+av
Hzy4gLEf6hUHFTTG4R94qYCtHYvSIBGNDM5NCH7E1xilJZz83uNMyTfxI07ujuzO
/JlffgqKa9k9eRFPqM+9xE0HRV+9sfb8FqVB8LvzPQbARCR6WuBG+6CpPRoDvEqn
rYhrWNrQWI7hSg2wUEEMxK9KaowHxCuNZ7cfppHO1FVzxPo3CbeW102/o4FqNlBv
plIZ5tW/7w4GTnYxVKgl2PWlhLo8vAd76WIoLS9d0rONkyp0Z19zuRbjpkum1IVU
NYn0FpmOWOfHgqkI+It4M9ccYLQWba7+HtRRa9ki5ksB1QeXfer97yQPAWofuDCT
FQSdsgb5R2K8fBYDEWDWghHvZ/GHs3nnJH6ORmjLCBlH8keHIpIVQ/XcqPa/i/sn
UpO/WiNRTmbP4zofM5xBuH3ytRVMoP722OMDD01Im8uw96FjKCp4ncHDiSJs3OOV
OVaUJpQPJf2DjyvPx9EGOgyTriiV48gRNmNHmrKlYEUX+PfFs1w0fc8dl/HNAbdJ
wFsWCwLPtCc8ParVd1ywjmm9Sj27V/Rup86n9/p6+ch2afdg70WH8F46AFsNaPIm
oFLKgxjq+XPJOIUcw/sOAgj0v2shwJw+opIjnw2NiBlBle1ceD6+GGpTITSVPBEa
BSTlRJ0WqGNu5NtxLqR10HB/5AxPyCwIcDRTTn6v4iBWV1K9e9xbJEMIcMLxr+Mg
mCSSKCS+rifz2w2q6FQtuZ/m209ZBM+BtaUfFXObzuR1BOgHtQHQ7mR/HyU2NJNk
Fg5CArQS40HD20APxdMwTVP0xphUt6N73sG31yLmgBlkbyABj4z7K03lTUYMsShu
P4wap91YcGAiaOLm1DOTOBepsF13h+lxFIH1GVI7demVbkceBGdxFOW8I4b4kHtc
244YG3zzk3+kttpPl178uLaU/0LLUHCIjsjCbEGhfC9PQtzZQVs2puDzn9PXSBPu
3FMnbHDbE8ilfrdYL3nRbsMqs0WkcNG/rYM6Vz4FpQ+YPjARkWRwhhcpobBOu48n
O+m/bxRklVleE3DXxay3EnkQHhzFsMbFigGuYA3RzA41VActvL4hSfTAXZhbMZ7I
hnqRuxAVdq4tcZixiTm3BojKqVctf/++rTdyr1jMQknNSEUDYac3Ifh7jz67PfQj
dFpVOPiMFEnWHm9LMnJk65axNUN0tHz57y2u/uchw1eZGT82cXAMFgaovuZonkKI
HZdOEBTOOdy+ljsk3hKownhCrbWJTrz0mp4e0KARau0ewftf/KP2NfKaIGz1cNhm
e8tmsdpkL3XVMON3FMeCSGF+SMUfgY4TewzIotcepkLETp17x1OKdOicjEBuomMA
wuyELjuOSSBIwqQJ/QYHjKAtOndcYAMw07jo8g9B8P+cgGt933oMUUEJrLQIkC5C
g+4nqSH724KuQyS9/Nj66mpqQIhoJLfde7czhK9brRgAMux4XAAhD2BgHtKDmXrj
HNMx9PAHmwGTxq2F70HWYUKf1BWBo4WXtxZPHlVy5tmB29wa+JJLl5JTfz/vPa23
51KfsnfoZaJkfLuWVJe2Z/05FRDIWqeqquzpZBXtnXQ3GK7QIHLBnBuhEeo4CtuB
bqN4gO+HE2Cb74uxyeq/SKiwB6B/dDbLgcMWdtqKZB3lNZXWUU1RG/HXNMfwJvdc
N/fLrK04jIcN2SEYB9g2z5DmcFCldK3hIRy0Kfa9iEZW9Gk35c2BxHfsLd4n91Av
ViUgEofAd3X96nX2IjArhy3daPupNK/lfMRy/sgtR+bgKZ8YgApzstWVClkC6Glo
yjRu30ZCG2FhUcyVzX3kI9jeHzOnrdRe2xGMRT8PZwhaho+FLk+DNGTAZH/5nlMN
PgU3zhEqjnhPA/NaSYzuyEjYviaEH3ivPyKAuK8Har6UvosChO1E9OsWjhjqotXb
mHY/OP7THcrWgUnq8I4qWA+EZdmMy5PC9safzVMasUgVsRQbHFKzTp224Xse1VvS
pSanohxv/Db//3ZcmTOlV2dW9Yob/j1ePE0e08KTjpQRcNXDPfldxgriOBbFsVvK
pTFzGonV9ojSfmMscdZT9F3cDtkX8xa8MJQu39vvStoYkKl4xM8T9eHeSyHdqEP5
IYjxUmazA14ZJmEpxkQ3WjQep9iF7BycqbCVx8VDbSTdL4fQhHx4aHz6JU/fZhE/
/HgevtRHAkrOIVnOU9tPcWakYHx9kVhNdOw2AATO9nZLpu8sf4MWrGdhoRM4Ie+h
uWIlza4xwGlhW5flWIuTv9ejGSiFYIgc2tvltE3y7/X94HoKiQN6E3U2gD6f2lap
eoO93o1m2V0ODgwFL9MA9uMqsOIvEShdcUcfgNNtdrJ7taX3JWoOICgXpY2IbKKg
T7trhMBR3AgQVEDMS1/yTpvoDBGUwk9cXSfFNX9oQ7upZPfCOcCHJXK5BacPPtjN
41iR56WYdVNaexDf5dj4D8qgC1JrBc/t/l75Fjcmh830CbVZdQUevxMPD8WLRcQS
QPdArUHaBDj/hXNprBnLgHkuMXud1ye1hI6BpQ+YTx9GGg27MhV0uQWoG0fbMkT/
OlXONr2uyWjDCFINr1xftdcJPhsMOxrZPHrulrVOn+mTxMrMbD1grcsYx/IKS+FU
RCqNC70yXqfbm/cpPGxyFvaruKQ1+SHqMFCGwtxBpqBv4+pjMMlbKTcgGdGq+FkP
q8luPtNyv6aJvYfSwGdbYBVlWlHG1s9GlcrxtPTrUL2BgzhyTI5IjBLcRCQ5QGcD
6+IYsfTp5bts2tNapXMobpacatzEyqRr+/HgSedDgd370JVsu4QWWn9vj5vYuIXo
Ct1mjOGTXB4F8FCmiEIuXJWii8cXJ//dp2R0uP6rcRTDhqd7n91q/ik9KYkovw1G
tz1GmuBwcCdkQm87C4jwvmGZ2zd3TDECjShhKFMAgK1nB5fLbeLi2hCqA/epFeza
fYXBWgLTB5BOeL3jetagsF8gXMnJCvvgc8QiC6vvSqH3T1IqI11NqdHgULqfhtXy
h+7Pt6mROWqdBYd7PpZdk/VfvXiPzQLeAUXyD15mnMQN5BOYIPTDKLZ59eYt+tGP
0SA9OoOvaYAR8V7LKYY15tgPeKvDk7Afp4wCtpGXYRfn4CvBLXTHF4ptSvZlfavp
0lUJcv+sAE1zzZzD0plQDd3RGo23fj+EQNo9oub7AoApoyf1WeJMYPJskFJeTUdu
ivOK5GGhgDPyexkr+6cDYrOYPv2XPk8UEEoLAO/sG1Gb0kvsloi+RgMSG7nwSR0h
Gtht0TMH+gKR/DZ8WGNiD4T2TmVWFRLGQKn3crvje4hveHfVKo4cZ3W5U8RdgFkQ
O2e1Zy6itJi2A3U5fZ8AprzE+8ROdkkNA2RMBCv1MzKrgOgTfQVHLJlNweAcj0gh
9G4dPLQ8tM6wiiWlUrmxGq5SA27pw27n/iPnV8Txj1o6if8SJug4G1x7EAA7pHNp
BZeodVy2315I0VqG9lZS3EFfiFVMMXdmwB8Jgp7hsHPRPg27hPPKsPZ6dWYsJKFb
LPN1fADVdQtnNDH9gfwxDmb3rkWLQRlSiTxuO/caEVOg2vFYbAutreny4f85RwQt
1RJd2OrCSwlBMbCdypp8kvr6KpKozGMb67xhhQCmOu2gIgga8dVtoa/rJDAvqQmt
PLlp0Md2GBGVQqI0eO5A0292mRubGKu24XPO/pUfhGQVj3jhoq5AV01MZiv1zxmR
AtZkIB4jXMFpI4d3C0txbD4XGhcjDrlT6Qq9NhOkxfcMTIcyxExo8wHNf8mDPWGF
V0+bFj1ooZ6a1mYJrrWCJK8NcuVxYDhcK+Nb+sI+1UZQGrnsaCyU0YIcY74otkXX
8OqxNZ3RoqB54oy/knB/902jwVdObmG7mQu+OlJIeh3dZaW3+z8kvfi81KJF2G7/
sDPcr/YM4Dsmt6tmzsDP5pnh+2a6vlpOmqiaHNH52afdMNGQkwEAm8iFmS3K+Aur
E0Ztlo8RTW/42Kw5YZ3jb33LEk05x/WKSvf8E+b4RAY4y1tSEOt8yw3XtRlJ7OJR
0/1Nq+soDyIpc4qFvqlcNOPBai+Ui5xGVI41JlHUDeDD4QXX29ExbcxqOZWFYPRV
sid+/r3Ctosqq6dIeuouZmvGvgTx7AUw+A2s9P334j0EyeIdX9DHM3oizcywMQZn
n0dm5AkhyAIhal7CDssb6pAQAhzC6b5N33mPDwXrT21WdoDrF+ZqAnMVRzOqC7r/
fp+TL5p0aO8J7jGErb0sfhqVch7qlcDmgLNKW1WIua6WcuhLRBbu+nrEFIYwEUmm
ml9jODAmc6QKtvwkMKlmO61LU6oltKMBQZGm9ORhTvgM1ZIf42Y4Wz1YVg87p1CC
5TFtYgDzm8kFPmq5lk6/e7nyJwOFB6Jel5ZNPgo1F4XhkULs98eV4UGzBNVM5bHM
3b33OR9iwjPhZszugVPjMw6sYV6BoWHnqIEBg0JiwHkmWJkY7iYx6vbOkPltT2yC
F7N4aRZAO8r0LoWvjybGJac15zmIC7OC3BCjEw4Oac6BrH6MqoI57MzO8ZeGXU+6
43NEO0uMEifFpqKGudAldnw7bCndaoxIZaoUYlaZhUI29rTLZ8aar62WuujZyudb
XnUBiJrJYFgo5GpZ0whxJLD+BhvFcdkz4OQ/8Hia35NI6tbEw/JcJ8l0yPInUHOn
Od5nz+0hJrNyCkEsSLK9zRqcohOnuU8VzF45dXzIGqpypNWfK/ddG3yJi4P0NrdW
Rq1fotX9jTBlsxQdvB08QxUy02ovyF/g4fgY35p6x/QOUBzHfAPLGMruT/+B/hnK
GOSRsK7zmKNTKy/rI7NHEPnXZBVg9qG7P4BdLv7OVYYMUirs/mjmVb1GwkQbPbOz
m0EtyGPYLmGFXmmhag2f+mhCgSyF0PRllD6WEnral3IlpjNV5gQ/fvZ+fParkcs2
xExEu0gBdPiRfHnlrjZT1Gi+bi/1whh7Q9vpBCHOprreLOdZ4j7jM51Ooir19drN
GOwJeOtqL9zIgAwm2EF/FamOpkjObjVD23eEiyRVVW/5EwrvaXR8c5f12t8b/c6l
O+NsSk9o6QVZP6ffQrDLPqv92jCveYVDRmaRtYF9RxHnx5yYs3Ci9E7WqZIEw9U4
DoPtTDOrXzX+db4kMvFftkN+WhufDQlkR5i3guAp7uXxU3neVqx44U02Yb9+qJOZ
AoKDRxGiPekjfeygAfjAicocPBD/48HEONYDbY0lxA11ekIPe6WZFfmC2hdKXOHu
lvuA1QQT/YNKn9ru256WVtIXk8K4J3sfwfEQn7pFg0pRWwbw1mwf/a66fXOmI4es
z3Hp02joM320gYMPv4IDEfLh53TgDmPHZ7cMEGcxLbiHaMyDuN0b555cI3Ev6pdQ
e3vLooFgQFtfI7ZfNrotE2htPuFLgAHpcfux/LXXwAv+Vin4Dy34CJz00INDTgPS
MXYTLhOjw+eTFxFzw84SBQg8q9jD+JcwLiS1C332CU5sXdW0UHD0eClSw5e4PSqm
96wpCpYt2IxzgXSEtL5ipDG//yUVjBCSgt0Y6HGK2gBlysFDTm7qsWsAz+Qx8Th0
mpkoVyHYeZwJ7wdnUM1+YiYLRxRU7UFbItZ0Pl1/X4r15MXDSq81CxF5nLTnFv/a
SwMGx92Y29eP2tLMzIi1IUEMVLRnbitIHcm0eb5/t4+kSW2rrYGWMYC8GpTbAx/g
nm7Oz5gjRTbq95QcAWA/qlF5P27+0/hBg5bfyyu8o140VlMPyiav63KyHIX6vkRM
02SlPaAMXty0+MujSUWCxyIG66XUmUvAGuCW4nbfOQijpJO5B/tGAKGh+5r2M91T
xcmudAndBOlVru3fg8pKauxTsGkNOxkM4JsxScol8hncVH3E2Weeu8qFV+8jU2+i
gnOvPeeGh4xmmjU6A/6ppq2G+dhgXr9vc7jbhLleBUOiIhlX6zf9jQi5dxQRzXYt
4uES+Gm4zYWEFzI35oKUsgiTCI3rj7sKIAbCaJAYWzkeEo/UDJs4XaeH1V8gZp+c
nhxVwtdIdJ8WizKgNgA0TEOZc4aEj3PDVdcH6QjMn2BfJnUXgVKDyuzNeaJDvqRc
or9PQaRUiR6dosqVngt7DSUxIWA+YJf+/KAIGIBHvcbYQ4GVs+cj/C5rdNg/13rW
2xKHyWTsYGfu/G6OCgeS0RAiHRQJNVH2jC0bztyQKBgGg2rS0+T0UeRc9TppX7q8
Y2Woeg7D1zT9ZntVXCglG2M6LFOg7/BQCcWOYebPUJ8AswYcxWj+vGw6wWOWvCVN
pY4AvjwCopd3B8On7o2RVPQqioRxkZ32iC53wXlDbwmSd36qlhF0FNDVOkA/kXIY
Vw9Alk52C8+z6FYRCzPnxBngKtVLB1HYksZAvTuMobX6Bqd0e/kN5019VpTDBUiK
aL/1jpDhZ/UWFkSMTve1nDsWMDCM4lxBZtE3/ASg0ejkVOueuYKC0zmyuH+RQTQj
+su1DzejvLIJboJkrTzPJlLls+z/s5AItmtpujd+KfwgZdPtV7/dYXnk7BLK4xgn
sH7sYufoUGf3Z0x9XAkZUH0taQArp7hbPP/Budeu00lEKu9t522F7MHmxnbjUtn/
69yGSKszX8OFUstjFRFV9BzokSdGfTU40CH1+LoS3K3r7VRVMKt1+oiGHqrg7uO6
ry97UJ0xKtUgY0Um/IjyTRnzLPQEz6IszjH4x63hjACCghlaGZGb4ke9vjZfzWH1
O0PVBHuamOQSrHhp3tMK/F3MqLy2lgg9GDHQj+51Vf0F83gDu3k8Qp3/VW9qvJ26
kkcBEIZxRxknVxZF9r8SuZTrCmi+7AM82lBxwtzPKqQjVZiDRZWXt2PXh+DXYnuq
z1rss74pVznP712xs43+7TtsJJHN693bW+FxQcHnkMsLpMvmcRtBrnvfDLrYbl+z
qIB+F9Dy5dwGbyFI1vfjNT0RzE3HL/KHSplRELjOXYGeHm5rWIofNN3gqVJnOC7n
78XC4GhyroZXWGzVTGJnr3nEBGgIowa8GYa7hR+VUxUvW/5j2cxV+e0LEQVq0yeM
z0zl/zL7PDO8n/cMBy8c0zP/TU6UKRKqJqz9319NJHmWCPwu6ERH4YmyfMIBtG/h
S8bNygrHpnYxrJ8dpsjTSFv+OSMdDPZvsha1lEX8by3TZxn0vA/Pq48+AY3zMBNK
To4ISFUwP2EC18AFdJAQ5NFtBVw5oE2kJBvkPLrOfr7j3c++8tQ+p3/KXqtixtvM
Fg2yTchnD2rbwc8HrlVdzCzh3a2ZXAa/SR8moGdrthy5E0lZ/9RoFC9o2PiCkxu2
s0XF+ehJhIZm02mHTMdFTHcFE4ikKusdYwO5rH2DfJYcyr6HfrlYAGt6HvgnOw/7
FsgMp2NuNo4o/MXLVRZXFY6sWkzQr4P+Xz7QxaB4qAe0SE6sk2v8aX678nW7XJ/5
mbo6TQj3+EAa0tlGWKQitcqdB/cr4x52YGnNQzU0uBkGeQmjNLZuXmJPqtqBCvkr
wMvm0Ve3q7pdsVrM4OXCtE8zc7tOL4sSw8a44aNKNBPzgKy4AeSncMKJjSdXCZoU
HSXp+mvr+JY1cl7FLc5z+8OrnGUbAk8hAWuBZQAGGgLG5Ws95GhXnNyM0cnB60ti
rGSzTHVmv41Oy4XUjFXlbW5iuXFFvLQTbISIIixZbjTBHagqwJxZBLxg4dq/Xk6l
2AeZOn1nJ8gtebXnCqoRWrMfQ5rrt8FQ9CWL8h5x6xj+GQm5B1pPV3JUzBYbEWC8
tq74OlkUk29YNHFKkkPsNFX2DvSMPDev+wjMVNlaSjXwOnp4IjsJnhRezesOpJsg
Rq5lThiFIe0FbcEPygdGtf5cvYo2hYSvekQJ9LORtHs9dTGmwP3n/f+TkN9FMaxX
6xbm6cCfYAjoELPwws7mCh7JyJNpSi5x9jLFOseXPiromJ32d6qijbonDuPQQt1S
oVmGCaoUqqc+a7RdYSxWyLbTO5blEQTVmZOIuEqTs/sHd4YJBUuGQwEtSGbTrkO0
ETwcSUvnRBpGZJ9/qY+5/SnBCerBclWtUdyDEUdhzsyCQq/vHCUO6q2VeOYvesRK
NdVoOG5WrbJ60EJZAX4J4qQYvU/bREsVuNx8+c2Aana250ywSMlYHbfW7N1IgiHE
WC9YK31CQwGpJipRf93/VCxDD829n5F7gkZRvJu+aLcaq0SDp9dteR8YY2AAYjsg
cewWdBdHbAOYboQn5fJr/JK4RdcSU3jEazIIihU6vdstPb7Lx56dVEdByYKOn6vb
nZ9k3u1CSy6pERnsub1WXEGmu6mxot2Xo/BypV8MsB4RVZn9z6Xs2qZ7zeOMvOYb
AMBBMB3QXeDlglFlHKkjE1IzgB3olUzYe7wfyhDwxuYziZ0epGpQPL7Y7Ndr0Fuf
rYSg4he0PgltpBjmf2yecehCB52/JO5Wg4Lj2HlsBoS+F1DlWfYWGITr8THuARX7
5N9UOOVvigyv+L5UyGU9eHVsVN/rKBH7x/HjPzNwOkLadOBbgMGghIYI9xwmltly
xUvRrzdCr78ilIdfqrxo6iWp6E49E/8RPYMZ4RXZnHsx/UFdU2c4BKsSfRiwEMyH
kkbwoehUoeBZUQIfGS+fItStAtQ7LjPZUYo0sEERTzAXCkY0Jd4p+1EXWL6niytU
9Mj5lTKP34B8tmthK0j1Nhkmn6gkKPsYHL+2lbZYEpjtgojqGXryBl0dCMi5wGgF
P19A8qYGbAvX4PqX2odcqcmfQ1ZEAjGQoNoNNDNKXuwH7TSeMy6kf9/OPxjZ1agb
2ftOW9CQByIlskusyEXuHsvUitTj5NpYrtEr59OAqvn0pVRJhRfJc0FV9BvNt4iJ
XyNjDTw8UDM+UF//Rs4E6zADhf3yg4eMiYFpNFbm4AsyU/PgRZQ30htoHnWknlxs
0guLXFYu5Rp42irnbNiHNSaYO7W8mOHcE0JzS1XSXUQFwxm/Db7xHihTOx6As6q5
2P/joIi5vUa4MkQfMSunwLD95yd4YMAi7dnM+H/Xhvf2c/qaVDUSRZhkMEIPssOC
ihJAqqN8rSRKimZrW9GLgAZmuDeGOVAPmvZQd1nh0heqDQ/TBv9MoK1tU1nNULw9
2bmKkw4qkoWvlQ2wvFeVI2ND2op4EjYtr6SqGvcLetyaXb7xYCJR9u/rfTwTCDSI
4AsEAyvq4nfFeAKZ36VKcoc+khyCM+dpOVucylt8xoemns9pf5hVWhVupoNs9ZR/
8zakRPvLYMvuNKuVRuJLGV0DwIkQe3sZ6OOcJwq77tuwMYQyA3Y7QeMgRK0wq99D
3f50panfOCSLjb2fxhc6Hr0eAn3mM8x/KtBQtyHWiU41PghowJXH53Nfc3TWdgVy
AuDTujNE+lIPIAop6tit4mjH7YSnezLHISZJWWcCrDICBF0atsiIfSVvUWwdWh2Q
pVxM/kaSvLL5SB03PAUZdQrHaaPmOZIfnzTzpleZFAoY/Wk27Dt85GxGm5gZKcFX
kPGv8ZkqPERn1CXpSSgvkICBeMxCxK74G+YHPLQ30nKqFixE5XiTsmSEkxWo69Ii
I6+EjdI0djMKM5VTAKi3+K5I8qFsf34g9qM/8vax+lD5UbiqGxQQQ5aKdXG1Em5l
YV3O9pWRcmNgSlyJ0nikta6Um6RLuW4npZ+2CBhQXPE33rVqrTVPvdvsgbkX0qtU
jjPvVDcW/xwWXVdA3ssc2sSgwsQfUW4pM1BeZp4NvObwjBmLmlTfAAaJN9VVqejO
fjJ6fCcZ+1lgqM51J7ovtqwsgO5RmThupWs/KyRdeUVBdv1AVmWfa4WpPoo0ktlU
+ahKM6yf5XkOkbaytCi4081j2+w/EcJuqXNyhwtBg1ObZInPXZuPFpKstAsQE5KH
BS/GQG07sQPneECj5ogwjy/eqy+HnJftAisscCKiVLtBcIUqTb5KBAluTH2nr14y
1EPzdrc9kvBmwn0iJWumTDv5yCcBfROCxNnfRHbwTTr4Ww+4xdNRvWNfdVH/+G/x
3BMdWtvwREc7LcQkQ8TfkTVz/SdZOX+hqaPY6H2Vm5X0s+i596SVpHRxudwnQ3jD
X7uave8S0ygognk2jcNBQnkNM8j5vIYXrtewVzVBmO9co84FJ+b9M1wlmdcrERcm
j3SwJmSCe6I7Mp1lZPRA8IbXjkMqiojo97Bn06xaXcAZAudeNG9HU+7T3nMsmHL7
Frk3Z+04LLFwUkac+3ddNGvQcECMHZ1tiaFx1DCSe1HqmqEA6+lzKwA2I7aTpQaZ
+3+xlF8ejI7xlmrFr8KUyJs0+hSu99Z94m/fSSTwhSvr0dPefPhEpc5PoDiCv2KQ
3Vo8wqQy2jPIhRSIwvi2WcST+Hds9tOV2AAWl3beEwkTYrsouLQfMipai86aXxwK
uQ/GiLUAYEJqxlQgk/qfCwQIfxeDRhfhI42fyvCOFHXvxw2l/kzbNk7pTKz9NY8K
o15Su7tNLqWwNRLVVjRCmsI+ePC8DAp1lWnKzKRxpNGcxRC+H/k/GIqVwvj6qpu+
TGTx4UVX6rXa1x8EjkSrVmx/SZM0K2djB/s/XIOR+hvbSTWGKAd2GId4Lq3VqWRL
IrCv3vwsVCLYxAznNBnyJub4gNr5d0LffSHus39o8q8hIN4tupHYk04gAkBI4pue
/DVQK+/2MV10gjvIYo+BqdW1lsW5DBGkFMNEEkwMGj32QdNXYlYACvU2zrMkyLJk
jrWW6TlFyhKb4cxPKSXt48teY0D97ae0A+a0BvvWNbBM0m/0LLVoF4mfR1pdXb8T
hS7CYBFcDLpdu7YqZ8DyhuHVshLjHHrdoAxb5IKYHV2OUsj3SXDN0jMtU39ZpO9l
xgS9xpkvkd+H6Fjqwz07LWlx9WX9ffHSSoKpXpocA7fP/eXfwwIyY5LIMW3Rc70Q
S8U6xeP/5n4Tva8ZYvjqu66CkVcGjxdO5C5fefJ3E1Qdz+k386RoIh4ITzZnzyWk
wbWUQ4Y7uE48RWUD8YiPz1exeM5giq/uKkJtUPhDxu6DQHngYrttOlAgtXMXjS1m
vXWyQLG/4+8nSS7qMTbAiK7ioNe5ssc1vi7cRWCQDGodXAdVtBDuXfVJLNkP6ULK
tlzPOXnvRhSjHVnnVTuzoauvXPcWXjW2VkqZrALcoQDcphEHh2X8ARfSgvKcg07k
33pfDmJT3eEj9SU7Aud4QNyDfaHfEvMP28m24I5orxAsg1uMFxoJYZggOkNTk0cw
ieb4fFW/lnt+mThJ+ipsme3vgp5N+g7x9MeYeKkmfUoXIQkVUJGqnhBOmaPGmeKQ
k4UHK4BqiIA81iYiRUfllgigmysKYEQIOUR1mXMPKuM4A0Tg+boRk5uUP0SiHbP+
ElVv5hdrXy1bio2G2/9RfK55c/xYHtEYbet38c+LCBRO1Zodpqj0MnzhikDEKl6n
XgjkV6iA+sLWeGfOd9p1j/acsvfFpM+lChB6SvS7p5iMiqkn8o1TCB5vdQdjQQkN
HdZ3BOchoFVW4++Rc4q938eA2dn7OriVd3UROMeCK1PurTBXSu2GLxMMk8KVT5Cw
MKXQwGuF4sRfDy6gf2BNYJuWPSl7L9NFXsmQzefN+xSkNU/9SKvE4bsf3N0cn/Sr
+2FZ6HxG4mXQS0bcQWP6FQzUs7kmqQWb4F4hhPU5Ixh7MbEQkrsFlK9LiyTxNAiP
YPf9wva5y5MqrMKsE5bep8dmkN57O0xRy+gc36DDFz+5sGCRnEj9axVLVTjA37Yx
rNFr3PftEOY/j98OmekeeKU8ibATmRVQHhtwYrkt2l2Sm8unl/Rzzk6P+0ieL53u
RjkveuL8w0BsLsQ//ZpqWO+E4jfwJ17zi3OSLv0lwy9SngCNkgFFQmt2xDr/69Wz
+bnf5LiE7wITn2ibv13YknrZpbvcJ9upGPYepBGkP+KdGKUKiMbZYnKvuNB2hDNy
tJSwkRaJhfiRxPcOawzdJklaYB8zFxa8+baSjelV8VM6kqP4jILl6UR48/6lKLkX
0XpwS/DzbbKN1EgxuPW3mdqZu113cm2+k157aWIL4Vfh6lJL5d7V/powpLGJBaLF
BCuNOTnVeafxkGVDgiXqJNN5WyUm21dsoWUCyN0fnn6pzufO4erE5Smr/bMLFqsr
5f6YDJvbBb3aJjyA+qWcfGvwsoALrLdaHg1JnPW7C4T8znMobYVzRvED1nATq1gk
dTLm6EHHo+0JnlYE0trIRkxheExI38N8RWvu0+G+edKT4ogPEJHoVRX2n+/0HMF2
Om+vpSuTlkgCVYTqZmaOM2YcOsrckdHPmFJF+qwPVaIWZeR2TZ/smb9H5Ew0jzon
iiXeE6ByHkmHNOUI6X8jpxQewRDQvJxY46xG2JtY8Q1QGBk2JXmDVsFc3pxUfTP5
8SJ2i5ppDgijI+cF/GbjRZ0Wy4xQW6xiXVV0NgBLn8fIfkrmACi0uvk94SIHL60N
qkcbNsTP3x9Y9LIeyMCadJtSiyxPo9D60HlVmnpe+47JMF+sW4dDC2KJnmWJmYrp
OAzYcMwc2ebhfNyo/E5C/T2b+v03mAmfkwMNTV4k1RUDYMD42/yIeA3ZkIx7hYCt
8I5wU6Njd730Ctys96qRqNfM6nBea3CHAxo/dNSAqC+mDBQy0OuynEEqXReRihh3
eQKLafduFqR74HuAXtdhXh2BB1FjY5+peHxdQ0z98e1zTxl9OUVpdgQQ49mO6E6c
nCojcoA0FAHU6R/1HOxgLlmHd5pfjmeyZOAhwvin7cXA/ySddsHUv0Ssvp+PFQxo
D0XzvTzQtn25xek49xzlsMBQyfwruW2TO6h5osuv4P8GToAUCXxtZDxfiOk6JT/Y
/GL11NUucVdTZcB8aaz2r6bpVR3gsG+llIjCZW5lyrD5HLNAZkzUjyla+uG7hHjK
Kw5jjMT0kr4CNSfYVC5OoNp4h7zikkqzcFbOr0C9wuPJeO25aYpmkbEV3utjXGBk
G+iuH1MzUnlHTl3HZoI6AIxIz+VNhi7Ga6rc5ZThRjrqhrlkPA0DMi9/qUejCTsz
JMhyA4bt/ccfYbHoSx0cBjOYgKIwo9DPt6B2lpHqaoe7oSiiLkj9WJ8sjD4OpF5y
lZoECneEX0h0Q6fUOvAbQQaBeK105LEEWx6NuCf/G+lMw5Ug5bF/NQ4hLK0gdjIe
0OHlrgxL2RtGQTl/zxZ9Zm1KW1RaQYFYpfB1ggymjWl/yHcUCTWh5V25vDpsj0dZ
18P5mfEMclfJhDlcFqidcdG/CVxSZmgxHTq5VxUW6GnQpxsqJrxBqtyqVAmh6DEe
F91rFq2dh0jIQTtKghoDAFtakF4K3rwuHIVA5sV3wuwzCMR8EJFPFKaeXvlHuSqO
DTJnrVe3MTiDdbZVF7CRLuC7oiwMFRpTCD6g4Qy6tJzUTA3S9D5/Zw0dS7zR/dkl
tMisP8XGgqYX4NIa5rhk2Q5PzfeKGfV7l2FUDgjVnvahNrnt3gb39zOfysr2+NRF
3pdTUb0t8Cs3LM3bcRpBkHn+ravcTsUmC57I1EbXdsrU4cNeST2PXjLIdAsuDRai
RUR857RWHNSWZclYXEOsN8lEFjqRXHYvOhWIDwTZXyM29Qx9P66iYvrMe2FLtkx2
AoDo0BSI3sWm4YEa2H++dPkrRCDI8QH/ZjKiR1IRb3y6TLR1dkxCcv/+EhCM9A/s
T8ADqp6xVumorYjHpN7jVdhpkObr59F/MxXuto3zBNPkJb6mhCC6VaNZ1Rjzbbmf
JuQ6KToVLUek/iCOYbP8GjnaUZS1vS5wjwRDQ/I7waBniSCTQjL6RNxah5Zf5FL7
041DmwkeQTTJ9/RVqC8Xh84xWjkRkUyePgFqdRyxrb7bD3uMxug1NOud044Ijsdl
72/ZLMmbQs3OBL7WFmvv1EXJUBnZF5jbZQOdNrbhDK4LB3TJKxeBvZrjPgqiUmfJ
YCxXysv0D0KzOKNf7HIfnT8gIkQ/2PwywxfMhktqr2HrI19zNo+lK7tdXLU+hAOm
gz/m6wQUXb8cTxk30Xn+/dw7PDAOZaj6naBAUHcE+IxwR0+ldf9LsH5Y09MaiocH
W06wdueLjH31llxlZLnUV4tr++qAT9kdHBfBXS+BB0U1bcHsYr5ln25Ppv3LmvYr
VPu2hjXZXdOY4oBJt9hfR/5ZzbbijO2W6FdqidwqyQ3YSfAQoI69gfVSaDiHZgk8
XzHVM6nsWE9vhaZ1MhHvDbhj7aBsprt687wwAhlLBcx1935/7KreaVJez0U5lXa4
zp6jd3twXBHHEcyJG4LRCdmun3gpU0Oi4X1BqGUxv8Di1LxZIj3EFhRc+/M6ph/P
8CGkbNSWiaUIrVDl/QeIttPG/x8boT4v/mEFXYfraUvGPWfjacykiI3jRpE4zhT6
675VnKB2ZvRhpcGSLYc/Kuapg0hihDDzMWJ7FiOK4ZbOTHp9KuZSrtwN7wvx0neo
zQsk/kN5G2YJHH15QULB/hBIfMBm3en0PGQA1Z9qUztihk4Y8SVdwc2U5mtBUoHZ
1sF/5uD1KAIeh+ne923UuYrYymVXig0M2q7/rAiKqcMM04+aFqmZmY3mI4mb8AR5
+NKun4IyW9HGo1xIz+MWSO+S5fkNtqkEk9qyS6cGQDaqum+CKXyaPNW5ckTfgX1j
1qxWNy5+MkpHyQgBl0V1NmlHTWAJpEXVJ4gBs3skeWHbzl85KaJcrs61hmu3oSVI
uXXkoKHm7D6TKAl4TsCK8oJYWJ1m9OELgwNKXkD1AqPiJrOM8YJB/VZxvmZKAOIZ
0UzHgabRacklyXuGWKQ3pwiI7cvJ55zQQRcwf0b6ID/pSLdYsRW19xUB7SW/ICUu
x0f1omxOdMfS+zPCh2/qawYgBlPPZ/Zy0AnMZfsU04nI2ytHNspBAu3StZ0kaHow
C8lZEg7uLulKNa1QmiR1jWWSGRSzkwEggSKiKk2/fQv093yDYyiC41YcLTUG58Rj
5ajEtiVwBga608nWibLCmmTd4t6ZI9ympH9CnpNqjq6Z8E6mtAEne5xULUpe0WdT
gbs3UXkILgUAv8x+nYkssdW2wEpTR/S4a29dGE6XLqSa40FuF+uOBLLbd5ALfqbN
GA4Ytzc/zAJ2OPId4HoCHNBiC4pSNOX6J+8Xjr4aq9CaIK4ESi58qydO4ZkPDtp3
a+38yER/86BnO0oFAVDZjcRp0cvqd6Z0/ySIgmC9l30+sgkgkAqgbre1vkO5IDFf
U9fbgudKetrK8sKC4Oh8xLpl8iQGDxYu9JRii2/INfMJ6mLBd5TosKIU+n0c9KsY
Ddq617ufJ+KfuyD/oVvmutPaQv8DAtXWAnjY185U0RE4hGa+3ToNnYY1hqkU+KX9
9z3XLcrrXWA2n9Y5M3XEM6xuzGOe91vMD3gNKXEjZrf73zvN6OKM8Wp1LWkwRFMu
hKgzbmIZmKB4W5+PGext3i//HP0nkyn6Z4HU/lQxR9m4gZOWrQoesfMGAfekXEnB
FOTCNdhAa4equ2CZXULCaVj8croIhhvg2+WAX/+YxjKVJRzrdaVXwnFMn91xdpJj
0CEkfD7cqoqT7DMCOAuSGc4lC80AkKh/Itjur0s0MsU8B+bUYEFQeEoGBLPk1pJi
8K4FmmE8drSTUm64TEU45jZLX1D2+CB1lKNxYRLcfeaRtVl/YlMav2uxAmefOnEj
pX11JJgdVi4cHoiGqJxAiGMAGwog1gxtUlbcAS0G93F9WJ0l8BfWXxP2uqST41A2
kXOXzZYUbQzm5+KCRgzVtK4G7s9aDyg6SMteI0OgVbFO/6FffIyeF13UT9xBGwiG
ThdXHLMrOb5PU2BCFuVSSV/YYXC0nu/htorCy6niCIGGJGDujL4D6IEQsIEW7oYn
1cynbkpQKwLmC3k+92G30R32PR7L30ahgwRcn+y3Xei9STaeqqW2SkaMtwfN61Bt
2Fd3zfuj0BK1560AJaiFw9AXSiKk974G9yMcXsb3UC1o97QU5CVKZbsmmMxLI73T
jkK2VLUSw3yG53iMib2+YBT7BwrLDkB9IdJn7vwBDZggDopCGMimeBgogPPpGMp5
hqT5aIsO6qlpbB+H2uUaBlsM1eExTVRXODKanBCss0uontdfw0EHuFtwtGri2I9o
Uf8sHtLrPCYrq1284mQHXH0ppCsqQ34vul31QcwFNIiY2E3pw9qfuz5PXEiOYWTm
IM2ZOr2wpvDoa1NJ55CvrZfUSAb432D+lVl5sS3xIPJuWxhhbok/ICcdzdercLFR
ZL6tj7qXVDu9VMZFLLtT40q9TJPkVtVX+D5Sp0okvzcDNwB8MLB7oGxwB72qysaK
dUEqbgmVSil4ZaqTcRTCf1gOV6A2ca5vlkjGSjQ+7TcUlBTMTPnNEBjcCPKeFExi
I3FO4HiSD1XQ1hIWkb/7lIrwtvKtz7LklyKmYqtljtR4lk2aRG/Tz8gwYCbNfoLS
N+06AltMvebRbaVFiFdZUP4/YikdYIjMq7U6liZk1bCthHx8c2FBNldsvMgwqyKp
TaBf73TiB3HuVKSF1ANLezG6pbkKGSF8pqznV8jnxGeV1g0YGRZQDHIPwy5TATMA
BItP4yH8JTGXb1KE2PXXx9ZEq0TiOoLFL+oQkiGItEM/8U7WDP8q9La69fXHMwpU
F+lTya4ey0YErL3F5EbvHBtRp70xX7rdq8dwKxy6yvfBBfKl4LgqiB0fDsvIvMeo
oeCLCTPJAe2iWhLiObgIPK3BVy4siIrvqHXF3n95U3osS1JYc0Y4fQKNHyCjxKOT
f6YsQPUlIGDHWW6HL27F+SEVUntVZ/FiFpS+Z0NM/81L+Wj+FU8jqMeev2Vk8qZC
Cj2/BriYZOoWrNsb1uJh854cCDmBEGVhAC0JiNDOwyU7DWEN1BUhIGWGJA7UekNX
6oR/q9coibHOhF77JcVP/97WBytUWPGhhSJyCy6uY+O8Wt6vJ1C9NEgu/SEkxvnB
BQWqSUorvPztmjN0ugoS+7fAkY7y6MUF77R9nMDdc+pTLZYf63MVq2KFOOZJGMoJ
h7EVKaBy/rszeI2lvbw9QNZdR9/mQvjfFr8Cx2ou2PywgTaK2ICxO6tzg8DkmZdm
aapDs6bCLNrq76CQKzUB4sOwyXA33DtTEkoxp/Xuk5/83zycGkRUZmLjUxaWEYPE
yz+EK3LSF3s1NX8Omz8vTlwBlTHtyU+JQIqQa7dgA5axuFAY1zeDOjj0klJs2IFA
H6XhZnyvsH8nUBzCi1o482Mx+ibaB1PfriQNgVrJX+YOahQd4ZW1nhwIOhUFp8yK
regKhl46hr9GE6mY8rXmR5ThDn6zlGz7ms513fjCxjPQ6v8pkyI5wDeHarhgQG8f
MhdOLePADLERnRiUMKvt4x4+ktXWy1qkCIGli152F7o0oBmJP7j8WAcdY4knACxl
pxoZerbUPLiYI1tF+HlEcUIHj5crlPozM6GdY4DO3JB9VReYc3CZIgf3S3wZGFRI
21UJ+TK4AC6sr0EZNQ0q3LZZNIHF9ZLLb8vFDYVOeOkaFWiGMo2HvQUimkuz2yh2
YAKsVnKO6fpZeDhYyrKE0d8jf5Tz9RQ5j5lfwLBfyA2gl5iG9U/EwRzRps985hl1
Y3Bz27iUj7kG5BoEb0SqumcA5YEgJ67Wmws7nsRrIKZcDlRe7im7cAABnXCXmfEy
3F0OuBtKOvtSp97+h1aDindUtlruSb78ODUGzDa9o5DJCnTuEV0ogD6KTuDi0lz8
A9yLo5QNoN4R2Snm6n6jE6dEkavfsBVr/wDrPB7O08bvPtG2i0TKGxL3fhBzFsDv
pHVHhwKinld0DsILD5BqPA4TBfqoHJ7GqoK6EAtJhDVc74/LpLzQLIymbSKUTQ1w
rZlrQvg9Hz2CRk8x/zCB08ajUgHegntyBRULr8lRb08uqVuzijXfmxutdqM3EyVz
HgEvTugKLzJeczcUwd+Aey7HmllNYiwQ7UFp3JUoXJjXQewRPafgk2iSgr0MYoxP
UncfEQ+2WGDNGtS0Jn3n5mJ4EatJiXM0GtxPtq39oZofXcDgLJ+bdecvnCTOYOLq
2ZVS+ilESg99pqmcHUV83IrImS6EppT8uLRG1tib/tZVaHXDEdWWF/C88zi/Y3sO
Z1CYR4Al6uaJbjX0eMz8GOW/ZCC8C9jJFb4TftPWJvjIiabgp4H1Epw3zbN+ECT6
LxtAi/45+G9iyHnXmKYl0DbuwXmsMpVpZ/7haKX8P1It1H1dr6i9O9XQMZOCHM85
EzeytzqLQAWnehIZgdaOl6DSFLfk9P+PuJUN4ggLrbfz4XEAfielvobRLp0cy0/S
8nryrsbbkO2mZensIQNk1bLOogL0ocvGpxq2O5ezanj4Iie492fOfhAEMByFOMW0
dGfux0ZENPs5Et330usnR0r5s9xN5Kw6B4U736W91e1LSOpWn3PzHVQAegYtxcwO
BU59ailDNqAhq3SgICg6nhFfCj8hhRuVtCKINf2ypOdOXKdlwIlQhQnBvP4ZkImB
wt+VZ6VF0kr5escHOz6Kz5059VUZx/3Dfll2K2ers3PPbc56LIAo2JzL3tKgNAFD
4PAgkAen7VlUEt8DJzwNq3Hk9KuCG08hye5eUz4Ff6qsW8AeBTIXATnQXdpQKd1t
BqZn23++eIu+MR3zXrD8SvB3ieMf/Fmkg1jkPhLtavS3O767dHLFN5xmElfhllWa
dTh9LeoSZweLS6Y4M1v/g0PrkHSbE81pFycR6E9HDSw0tT6E97WXPdBZ2l66pISm
cfy1zU3NnaKJdSJDH/WitxYzJFlgDvtWNqTU8hvbuAD+G19y9K1CgiH149/BJt+C
qn/o4/bPkJiEUyt4qRbAD/++gn5oQsn5K3cicS9BJxNdvpD/mcryui3Tb1BlEJoy
Khb6ZF1Ghg+1xVjk5w7rmtgwS9jQXmsysX9QaI42Vm0xtKxBGdeDzz6ngnwxRBZK
FT6OxaCOBgpz6Urm51TBNXYP5DzVv3i+cTYT5r8yewbILGS5jYi/hiziyKKrv+ps
fo4aZEZG0Pjtmp6nDZ3A6UridVwUMzI7wNu2s+ZZ4lH2Ah+4IP8QDti2gBrObZ+9
5wzewS0nPRUDXZLKfmGmc+iiNkogX8yLaO0YcrWKFl+4JEoawqMSvIBnVxkdQGYG
WgfTvk86jeeyMwkFzEtpn8z3pgUkYKd/pevtDY0kQxnnjNwxSnds90PgCW8sduKe
Uezr0EVnMam52iIF/tKz2YubltAV62opZ+7HG+Dz9Ybz74hSNp7EcwKBkrQ3uHM3
o1R0Hajly5MU/QlOmJQO5gljHAo0a+/F7Hs7D3YVL9QTaerdR39ER/JymhcLzm2/
vLaexfDZZAQjaHALWeBAuuDEhzWnSIbrPJtqKbeWRGBw5486J43HuBYt2ZLjWjMt
pcEuNmGPbIVqYsOkTJ+iamzrCph2axLv/XVCrwEn6d6j+fQjuWC+lFFlAVIZjx4S
C1Umr9bsEV0EQ/vcQZKC4hQ6/GYG4o217y6L5Kf43T4UG4DGeien7D4xZzgPaxdi
diSXvs2pY3eSxWV68Hug2ppi60NdTy82W7fOrfFV6VThQguQ1sqiiZaU9fTz+geG
vXV95FtBxTp83HMmkR6+pYPwUqQdidiVC03EknBqTs7pLiCNGYqCRPM8a5FnzcbD
6Cm9a44CzhlypCBDo1Ca3FVPILDL1GXS6UyVXQX9eKQHxIYTLk70kGISl+Juw5Ci
MlvWu9pRnJOMCMrxompllwfrLGzMGgvIFgmx6tqKEwKTUBBBVJLJgIkGSa5hR0IF
c/KjGa6FVym9uWEH3pL1TDQFLjEieTh8rPOzH1AK6Amcnp1Tk78lGixV64l3EI3x
RT+4Tjl2QtWVLgStM0HsT2maORxr6FfUcwGzhPBr8RYAw0IJNlghNIivISdDm7F+
Ag/NQpwnMU0/JNdz9tqe2eLR9QY4MXbkG2d8Nex3fEgTfSrkXuCz4LxlbFO+l8p3
DQoUZqlumVyametEdZanw96uKQE+QdQz5nVwUVCgGc4t+dB62HzVVD5hmZCN11Wa
Aq75M8cNeArqvutKgdSTUskm20qlWFFNFYhxpNzLmQxvbaW6Acv4mP18ls58zTdv
cQLtUHqgt9NCncFkLkB7ufd65B+y2RR/LYhUyJGJ+pwDdfBefu7RWQ/OCCQ8oKou
23sc9aMMklq2tzhQsks7cIqPKZrjh3wX8jWjxF5Z1MNqZyY4osxCwic+HAasfMrw
S2Rm9Mhz1Uo6DD4ZVD+lFOjiJlh6oWNGz2J1YrcCopTzr6FTNyPPv+8KoGwOlAfB
DS3EReFek07JukahF4Hpna1b9WEW07nBn5V1GrqxcjGxz7/NVQecvCIdeCb9pjZQ
IkwExnzvN878uYdWHibSnLIZt+oiyALPxxvwxheMRcvz6OxfwUgCb3RhfwEdHATc
OnqPeglX0o4CD+bfaZSk5FRvrHpIW/sk8Aa8Dvjdo7qnSijk788RC9Vac7ciP0p4
8mjSAfoyv+iVL0GiqsQcdhGM3fZvF+B3SF9VD7VOFYkeTmii6FgDaySyX6h1wTKh
slx5AVISMXN1937ingHb9mnh1+F7Aj5xY+jCt7fvUNpUhhdoSDbpKuMx+bg8KqC5
D8xhIdpE82D9DTLdB8x4ZBR5rKU3zdeI3PtC1+UcHxSos7Va+lyz/apqiLgs0N5D
o+CalYa5KE+VUDK784jnDbRGzbUHLOikeey7hZ5hJ6Lg8FpouQnknaqiPe55/Ge8
slBGNFriEjzFSd4vRK4t9X2ceIIQ7t4N3bXvq8T+biBnd780noccKJ/ukDADVnwT
KobQTEqM0Hq4o0STmcRwtr7vXOg4+Mym3SELSQPsVE2xokXDc1WI6s5gn10CPa8n
tlkRTYmWf0qqceQGlPhwn9WbFG1cLoj+Ek2xlZDuHGIOQtLnHrUB26OvhjHH1LuB
JN6HkZFh0KqxuPcq+o57qApwIdv3IPQB0LMSljGnC+3UXuyJnjIooZfgiIKd+tI3
f5SjWO6XhptKP7DIvcD61kh+/H6W7HYUHZZ1P9rcmYjxyI0rzConripXUGbgHpGG
AkEn1UYRy3maXQ8iyb5vD11s5f2QhvaZgV59GSfJ6U8uf8TuVthvX520UIms50z6
4clFZh7VlBAR0roBaBfT0NoM/bpqHEtR8X3YsOAqBvbWnuWynZ48ywFgYWnRhCxi
0U4vImv3dWNOj8NhR4QDT4kjIXC53BXkNvsURe4s+10hOhhxA3kgm+tqlL8oDUEg
OV0EbhyCF5Ho1spRNa8T8nxaeq1bqelpoi3B4gBWJoHQj7SbUkG1t8lJZGFq49Lx
lphVSyN1AB+3MxlH1dO5jvZrND2pcE+vWYc346K7IxCXzdGFELhDeXXn308XwyWE
K4gt5YRIh/H3sg5lzefu3dQp61ticlJ0xx0Izlun6e7o08v0DINnoB+Zqk0K3NZb
w7t+UmbEUFCd5XSvRateDPsAj2sj4uQSyMHdpeo7c0IthEpMQVzgWK0UPzcKFnWl
VUOBmhU30AXhOs82eXb578RMT3KMVD0XNJmdmLM3dQ8BtMdwgJ52L0LEOXNVLe1F
qXI5YEUTe1LbgBSXkakvZz9KbdwC6PsbM/8gbkHVlKTjYt4JWF3ICQaauvj5svU2
hSfEaHlRCSjpqorcGydGcwgta/fSpAcGXBjejBAAoOmkvFtLTDWMEaEpJxmlgQ7k
bA0SEP7HRyXdUwbp/EBsXe/cbcAfC+wXSgDZ4mzuPJWPWMlInlsRI+iA8rIXxgyb
XtVNXEKYUwSp4faTWcRSBgOtMeYhjpaS8ce0YroEseOaniDaKMI7p7otfxJqkW7F
Us8c0eRyoSgcEuXGDxoR88hCwknV0rtWu2K7fMNwH/ssPT6qiySkEp+VBrmmfu3P
sd1vVADAw5uFv7+1Xjaxj7bBTv3le8St3aEvdRBKUG82WDnn/uoc7pNl0cCV+dJl
FsjH3mjTch4qrXDqSwOryEK0FEdnntyYgxcnRongtQ2v+1TJ+h37vxP35ldwVY2V
U5wy/J2h8eUVSjoQHVDAXyKI5T1VoWPBRnBsSxQtOQc5iADJdV7uKt4KHiSdHlm8
SateUwa/WPrfbhbmpqHNDgMsEXcvXbzVQhfH0akHzkL+PkJ9f1dnHrbby5wshWyM
CFk5E70X1ORwj5EDQzbXM8pb6U/6m2LyVzAWknfrAjiPU+jeRS1rWm3XEktk6Csg
faJpfU2urXpmSg7qSJIH+4XFCn9pLcyw4gx3gMPOe2+ka85h3fpj3XwGNy/caCSQ
P4/jjU5jgBQ/xQ6/fMFWMDLFY5eXNRPMWL4EpFwIo5taz9Qj4No00S6NtuLYGZLj
qlnRvxzc9DQs0wxjrhIQOzdAQW3WsacmykpvPflNmatfwUBRCiQx6W5jqs2QA13K
cWdsbxU+AWe65BCypjEmn45HicSCHdbyLk1CXe2acGE7tM5X63ssM4agfLIT52dI
bbFQ7bfbYGg8aycYVXsTb6t6/ieZSHzv9DbsK+mDiDvib5mHc69Bcs7tFhws/eBL
+6ok6knx48M+nzFm+fV19ytCStP6jjRyP4se6sMcfut0SXF40lc7UEM/bmdDhp+W
i67oQrBsVnSIILqGpFn6G5xkAHjdjf55uyxGuMPL60Q0ZrNTZU8DGgBjOa8f1ZmO
3736Yz/NtqSFf4x1zjHSnXdRTwiE9RI2X1G4dQsCP3TXM9pSHsLiK+KyV6i/FlLr
86j2AdRI4ptDna4NaujC5KcbX76wEIq4oXzTma8Yd1aSNaRDWH7DEyDyZ1iPAbei
mrQp9KF/mxQcGntV1Uj/+Nv9iRpQj6C2IBPfis+2APbeWsSsQJxTzhx91fV+kbfN
8DbPa+5Ll9bN6DQlWKHs+Z32y7jEf4jbDw2NF/yZt9dN6TpFrXdIW/sOwFgPDwFR
tTR9TAije59bFjmw9vY0aSW3hVRI/KXKanOM3mgr8GOfNHcIN7T6Ys84OFO90BE2
pEq5RZrWTFPmLSlvsQSRRkXEORP5ALowGE3+X+r7NymMrSWTNUmuNUmv6CL5QBQp
M7Um2oBwziQYFgon4gGkBE7hlusjx01mt3hUnj2e4ofo9vlo6ZblgXfslqFflMzO
iuB2u6s2lmCQjfLiMEK6kCoVKZWTiZi96RbuGKUENqkzTML3WJbHvacVEWx8SMdd
0R2uH6ujRYwCxbSkdbi1RmWSqfmujP+/QKq7bMiVpT9MSWfrNYhd3IJe+484+SRy
O8f95JPMYv1TwM138KVhACZDnjw4MJzBjGIzKbtsaYZnkk7pOThi2O8Ls4Jdrb2Y
9SdbIRYAJGSiXHcBlMWm+gRjkQWbI7Nyn0rENriNI6L/J8cvMctOD7FpzG5bjO9v
8ZOLmqxZYFc38rceWK+VCSZ8xXdT7yMwieP6Z//8gnXcbvfeLSJqFS5AaxcKT/2U
QPebKXj6mS5l9wcP9SVsHUMX1duge6voKjtWRWN3ed7o1sKdrcTtSe6Gu0tMMWQN
PbnZX3a3Vmjc3B5M0crrJ9/P+C98X5xt3l6e5oN7yDHeWPG9dkSel5VcJrsM37iz
J24a/IOPmYJ9yLMNCJTBCY6RFXi1b5VNy1RwRfNbYcr7/6XJTalnlxUps4tSSycu
U/ShYh5gVh1d+Dwvt1UWu6QUWmZ3DiWuqwnyJeYX4pu88LzdvQU6znTs9NEhfBrv
L7mDJNzQefXILZ7Vz+QjmsfwiPU94SlR7u5vG5gD8mIswpYgrT41I+fFYGhWC3vB
Vwemm8A4zxicmlvW02DXgGM5NpLOQieK8mZMaA74+RCOzXOJ8ZXnvExBZJZTEVl+
fHlRZDFRfTIMjBJLizTDDATqo7OW56GmJTMTeEnCJqiNMwLVDTjcy939A/zp/hU6
ri53eRhpsW9XbD4yEXsb6CukWLFi9nT7OiowlsK7mjqQU8jLl8aBCxo9RYMHhuI+
0dgBniRyD/wle012YXmbDQ2Qwv1bz+mik5FBm47E2J/V9SmUzApQ2YEyjKbuaWYE
c5UL8F63clrIct5oJIalGKezFnv7Jp5CVmwaY5Q3aLOR8oCH25ABkRNY24BfI8e8
csTGhKzxK5NBpQWGw8+525iZzmtoIOnhvg5YSBcOjG/imuaU2a2DvHFFN5gsRIdw
qpTkYGh0yl5JxugIGITvlX9p9wxBu9lRas+jczrmD4lx1YzMplo6Y2QeRjSKTE9O
hUyJr+alhqqKKTWRR0wvMASePWQOyuSB/dEAIr4uu3euUin7bkcwGW69yhkYI0MO
dWvYOsBhszSzn3WJNsRR7wr4ECrGAAi2o9sLCCDIgoP8tyETTf0KSNunuLSo4TMG
jqpiGxc+UCQO1lG2UPH9YCcRTlDDYsfGOjq/nzvG507/dblZ3IWcbmFpTEm117ts
e3yAvR2gOL+k5VOvT82QxOgi+zDkI67UwY0rpmLBnKyTGatuLwkYn8NvBURLxJPW
L4VeoBKfTCwoRWvbhDybz9vQ090l5DjumeOtNap0sOdn6SLs2BdbQ1mwHPyrxiOO
NUmqf/FLpUX8wBUft2Jadd7vOpoQfWDfvJGKNDjxjAKBtEQWgcg90q/NRqcPebsJ
dgtUyJgSr3B/jkb90PWd9REB/QdTo/kkt+UvP/YdibI0zdkUy1L9DDzB8lf5v/5F
iej+42EybjZGGcDpEtl95ueTL7vhgnUZKGWBGByjK6y/TXMSH4o9uchZhNkZeL2j
oTjJJr7D97FOtJYoBGnFiyh9KKvHc/WLs/lSWWdHvPGCOMjW7HI1iiiTyIHzUzUR
Otk2ipN5Ix1DRnh+59af9Kw0I+HPRSkR+1sepdOKoEsAXa0oVxl8lNR2LfqhGUyg
nLAKdyjoX430DTEyAufHPSB1NauVwlmlc07btAHnwzdcQF3Zhtiub1Ex+Pj5Dwzx
rjNitR46zbs9+udwjBiCr7QFgVIZGs5NKdw2VnepaYFgliqXGE3x74V6yMTP85nV
C2DdvkTf8rbMvVtLbSzcv9icx9OyKBMqedXTivj2UHAsw08JKR168jn1Ehjw86c6
BhncsIr8wmTvs4IQYGDGAGF/mj1ZcvzcHdLSxpqb399PIxYxI7TKxhd1zTglarZQ
H3W7R9wCcjP1wJ9dfLOSXqqpmujlMesFq4JoJcURfFS0tX5QMYu5940D+MHL+eXA
YQdyzlRBiXPrm0rveaf5J2pFSEKfGEN6ii0uSnuaCcfIwC3LTHNZ+Gsmhd0AADLY
Kx2BRBnxemNVoyO6vVoLQXiryAImnohPBkgdcI3WNZ9RGqWMyxqWqjgauBNKuZWj
l4659EyqzUZy5adAbjLhg4udi0DBQWVuaddd7g7/Aw9AD0j6hy9/xwoXaheUFGfx
+ZvUGEa/NvIsvZCAsSI+ia2E+LddPQbJKA/srX1kn06Wf3Q+kW6z1FV1JwIkfB71
8OXFgNM3GRjkuoNPrZjOmk4YyK30GaSLUcriHEpH/e+3gAdoPNaTkztfoayRoO4D
AjrLNXn76Wy9Jme8qWWR5CZeCfaPUYoaANgbchqfvj6fywt9u49qnVnBq0WJG3KD
RaWAbhjAvxY/WAq4VzUGYltDUc0ciVrW38arE7ueuY5ZVO/8iFIRn26PnLt1Wboo
JqMdTv6CCr8hQ6qzB54KnclbBTaUTAwMqOQ0TgFYUcq/TB9WhR8SqTJyTWQfuQOe
FXerXbYokPORQMTc3Gisla2R3c4gMO17ib/ch6DK7cdJhlpnIxWlyQhu0jEkJAiO
D8iw5/SfQi8S3o+ntqiidfWO59HSOOv1P3xyBfkg5VmWF/f6HuCdmKRJrAhgXzDZ
BYWKlgBFj8FG+LNMP9M5x43+fSnsKdqy6pXwOanqeiEY1IzXrrGdT7VqkvonZE1L
CT8bockANTkTfvBBKYtooXW3IuwT6lurB5f1OERg+s3AFB8mnMKn07sqbuFS2zrs
ACIsBeOoVUkiCZGYbwIt1gmwy38tv/prh2O0mScPsRgp0H+SDL2VSXXNGY/j1VQN
tps0nsptV35Gp6vm8wHrHzphuSP0Em65ZxTsZvg8Q7yCX5zWKSaVtjxWNHwIfvZd
K1UbFOipEREs8VGyVy+b/+ewVlY+kJexjVjtFMwuc7g8Hbn0bCQhNjth+tlnucIA
h1ggK9ENfHtwUylZlx75bDa+VlGD8i3oIh0ArwquhlyLLLIQ/aiTIjRkpZBvhhz/
AVUbijdpXvnbPuOYkOIg4WZs0toVxImtxqz6T1DJU9q83qkJrTV1/wOgj7GyTXN3
jjbI4qxTyno+wkb/GHeg+r5Yx7oIyzOxQtyc9nNppuCKtDRlRmZ+JS+hpwYw6hGE
dg+j3AV+s/WRbW4+CYmUNQpX9Of+VS7LQ+390vuO/ci+EUv6Dz85fOUjQUZPi0TZ
QIWtPtE8ruL/WxuHnjTkuuGRVjmokDWysF1nYeUtFNAM4IhTxWqM0G3ySvgVGYju
G80i5QHI9QOP1qNoiHm593C6rQ8OP3fGpmClXYBM5P7PudwZyzmYfm5sAbnvcunI
E2C6ofen2uVhVfPYcZ/7bJadXT6rqx1poYH9osnb4N8jHe4AKHw8pe5CfSlLZWbI
p64DArcjQq5JZ3bd3aWAc7l0eH6rZwKuZ8SnSVvIz51WVUkwT4bBnigvsDDZ0GgH
9jqKREQ2Qp6lnySDqxhbqiSrMrnyLPxndu6Yy7PaY2pdn9W0W2iPDnsE38OVjljs
enhO2i0Jm4OnX5D1ibf/7ffsgVW3RhQKEwiUv+4RtfQTaRakrLb/m8OFt2mNUgr6
nznK9KtFkPyoAXtWd4THC1BsedmdAtG+idWKQJJb3HzBIWFu88XZ8N56qoljZ/Ge
p/D+vwa9sVFDiHFnmOj4ZqOgIxPK2YFUmHc+/JX2sjGQFBCKf9ZD+rgWl0XuqowS
pIoYbPxbDd7oK+0BvinC3flqfqiMu47JDzazPXy93ez6d2Uc7jmo7kzxMXIImKM0
KaR3JpybqfYqRF8dIS9zAYV0EXOgn8QU/hmaBeug2aak/T7N9WnTW67ofX5f2bfB
nhfSobc+CC1VivIL7gBOfMoUMYAeHCTUtRYANVohI/Ebvea8YNGxsuP8OWlchyTc
Tegm2ZB6Evetpq0bxl3atOQFFsdrTc0CBMB9/OjwEVMTTmDLEId2V15g+amTaaZv
M+ajUy9/y4rpCOukFtytXWduD3BLYTPhbHCpYfZ6kA/OYeDLxPgD9KwRZIV0mq7r
GQ4bXfwKDL8BvyuGR8VYqGtoP3s/va9hyhgCGhiTqclshYq5pAuhOKvT24aLcfFj
DY0LzEPXiIccX2nBLYdD29QARz5wo5aOtWrLvtoWU/3Z5ePoKvmUgVQFCakkrwbG
842LTcX/tQB7HYOoNXJXpPmQMRPJnkjgQLsPXl1OVKhDg0+8UiNYFVPx33Ev8raY
pNhMngoaIZ+YltzJncek/OuiU+fxSuDQ65Qyp++nty2XK7tNax4Byw032o0d91BC
ZzTfpRyvZVgbjfhOce2gHyYYrik8HEmODW4umHWxLfrQPDZ2PeL6Am0MSGVdG7P/
n6Dt4ixkFMqe3MBm6Yl8V2NqWV5R5onMOa5ZzqXixBQWydg2AHxuIgKwmeeMo89W
YExEFp8kL6CdBJ/T5THOqGvPBSv+HOt8tTNkgCcDgGeleftGXShFMRyDBliwEimY
ojS1q8ON7EGBxXuUyxKL/W910gaaBFEctmYUpMawGCC0ImrVjb9eNtSFEH40P+sE
1giLIXZD0qEcrgNRT2tkasWNgUzMjRHVqE0Cih4QH+gRPCQ7jgWFLP/AuZLuO54J
ntZ3cx/9uiE4DDLHxAf0gSeb7t/c0fc+BxT/WEEuH8BtgZsjQDVwiS4MRrtPR3g4
99U5VcXZXMAE4eIh7+xFBA2Y65pw7KpqbKGN2n+L210ZCohDxkPWZzrm+MW0GqCa
UrzQ66Q7KoYIDCwFWBO61YuWNTQ4KFQwCqmzlftPo5DRjPtaFyBelMtskvbZONZT
RmXfh8v0Dk//EP9cs+F0LmKFf0Nn0wc5BnFRxKYiQqAp2vijr/cMjTHHyilg2OyS
Jc2yqDydA9YRmF9b0rj19PsjjiF2kWLruuCiZt2Iu/MKj4aJZXSjxKnCnGaSNq/r
fwKqXssb++r+XDJEhQHFYzI4TtgdKqEw05clWLKjXpWCeZBIAxDb0sQc3WUzWEiA
ZYeXdnjbpSSaHaSDLklDGlMv8yb5Q0YhZGgf8kcE0Zz80VEtvx05xKDaYOUyv3Cg
21GJJgi5vo1l0xr/0Kv7SGXy/viZXQNAKh8ng0QqKUPQL6Wm1hyqJHr5G9aknE3j
ZcnKCXacvVZfrbaUqKN/sNhnK/KAZ/OIhjvwGRBvxU26S7DXKqlCK+PH+uBf9ahL
GOMnsRlf5iyiIJ5bTGypZvb/9P0ut4ZCmiEPLfy97ysReFbySL/BMRw2HhxpBQ2m
arlUA+m9mxQxi9CvV5f5i4VfJ1ww7DmVOcqOgTQvz8WgZS8E4zKMVsFWrfwU2lQW
IsCVE0re05fdQVbkV2NAIrfx3p73aujCzpEHpUIQDmkiP1AG1VA+FefJjSNLVkAC
othqVWQjqgIlUGM/5ZwyvOXWImHwigN54Yxw2XiyDu3CqRpPasUSZgzia74y0ND0
+IAoeNvnc+Vf+dykk1O+HUpXpsAyHAQ8OSy4eGeDuBNKJRrIHZMaf34F6U3bKGI2
MHLjoRRTGTMZ8v0TWZSIZJ6d1YY/u0uWCDtsuqwX9LU8ONiTVKNoLbbZ6AXoYaEs
Gxx7KcWjXswH6SatovyVLhvGTZH7n6IF/IuH3RdFJV9+qZAyfKnuQwjMUrm11XyA
NSSDmD8NFx8Ei9BouoAogjtZOUONUuI1yZnXFjAUt2ZhYFwLTB2IQD1vA4zLC7Hy
OU2cIINvF/lTVwdAPMdyyq3uPjDdrtKVHmtNIOglvMSO8Ew9Iwx+PLRW/CZ0qX1b
l09FXLuYLHX1AmyVTozDDsxS1IQWo49+i8Fep8wmomtwCEGuEMwECs3T78LL6YCi
vhjyybnkmYyQIBGpAVBaJNwXVP8zzbV9iruuMu296CA/4Plqm7uEnYfqVqvLNSdW
/icp5jVz5XZr6Jsw+OfGmhhWFeNyTRujrNCqjW0SixV4QqO5UCnX/DgckRkw31Vv
cTkAy9u6jYsXLMEC5o3bQ2yvHCberCrjyCCIagzeVoo11gDTtblusx+b8QDcROiV
riITs0lzBcQFJteQYKJSwF5m55SmwgXUdz3n6eD/4ElbuPKuwkMdSs3J5RYqol2V
pDBKxso1y+Cb6Qc6wQzTvA3QRAqho33SMkqvkG1btvKY3fz+j70ZQrDNCs9lvg1G
vnIiIMaI3UkIDk3gSI7JEcGOiciSQlIH0VlqASd2Mwy/tIhvtgVIywDcJtdTkdmD
mZ4K2AyCttwFsRQzdMraBfYxbtrpG+brCHVf5aj4ZT5VbiYeFvud9blgwP9jaam4
l6j8a8GaFM0dgq/fC3gx7TMG1oWe5gEcBhWwKO6V/7KrNKgiF5ycVrMX6adap+9f
xMsMcAzgMifjU4fFnUNuAmwI3bqSHhuyFJzXCUH0A0qz60N4xqnrMpJuc92zET97
vtw8ozjqgaVR/eF8SAUa63xpUmQ0H2Wo+eulxFIm9n6AeqP50rEaiV+sn+Qjv22y
RU456PctISV01hqrITojFxFzb55l86Q0rnDKq3iNFR/wLphT8qRRV7lxRsJWDeCe
SdzBn0wozrR8rxPNcaEcag0bKVHf7xdSRvXMHHhkZSlK+GeHEJzP029u3mLJClud
nOKKy+JTikX1ghUSgjB5lO5hrsT6Z78XtyyK34y/BY1QZMKIPv5cfKbPkgdA4cdP
wUP4Rqs9Vle0xPHN/a2rj4MWO/C4a79ugbVH3d9Wxo38A1pkFT72O5J+I8FA2Koj
aGIfuSIgzYpGqP2JFCoqKCWugs5/Mey/ZE0C9tNhXdDg3hBhOgfwQ2uSLT83AECS
aZPzqzRWW0kNnbgqTMgc3bSEj4WVXrDByvM1Ut0zyXKBCuwsyx07ltsghECC99Tz
B2bhtT/cmImNWlLznEx1s+Cp2Vsc8E+wEsW6FkijJPKfFnsHGEUsoXraS30yCLbh
giT1MU05JpIms0HIG8BEwngGAeKidUKVBaAfum9euLwpAPJMjIDcAxRC9XyIVn8y
NiUxFNxm5kl3IyAyxUgpj0OOwzdbuDUNcoxruB0Hw+OWB/2lfYKFDTTJncLJYhbw
CaS6qelczl5dF80a01Vx3x3INTdQrrsQ0bjLUlumKxZ3foEit/PFGS0ZkR0JqjNx
fmt/7GmJANPQFnpIkKredaPhat+NcYsRNtxNC6LBrwarCQnoxRVWXq3ghh0E03/g
9yl+/GZvU2hPABcaCUdfmhEGZZIhWjtsfWsPhKexprxQEcU4KIfhxmAzBI0bcqeK
9wTgSrIND48zyrig0Iw6+7ytHb0FTOPVCGE6hshrv8gihv5juMQui9RQHKj1erJG
/rGftlJ1MWr70cQojJfPvVsB97DXmwSfP86Yrv+TyGucfj7/NUr0cAIMNTgLhLFE
W359+tBFTcB+dWVNOmSNtCI/xima1fRiUPq5av59bMsdFG965Tq4ucqG+j3csnfz
gdTxVDmt8pjfIT6YaM6BJk7DssBsJQSqEktIhX7S8XGE8acWs0lK8+UDkhxni78w
6YpVIpARXjce9aCyZWzOTv7DqxMRYYraGkp4bOxSoBSw42wVXeC37g1qY7IcMbWR
HXkvV3wLZBZcsdEO7z4hTInTWzscLY+1eQM6TgYYMp1dxtsW021abRkBe/jfPJKs
PhytPwmg20R/S7yIepJacc/HIVJl81d9A7xWR+FDHZcAfAhELLDzRUjmPVqrq/Mm
JFSGgrny+tyNziyKCYeK6usdbEEmQAQ95obkLXRehZQEv3CITUEF624shuivFxY+
7XJ+z6osdj6r4YbjBIZ9fSrQXjC1QbVHSYmTQi2ALCzP9mUDuZSTado+yS2lQevb
mG/0Q6ryaCnb91wtgbdnfOpLWXUSM1JOu9JF+81LLQzK3NJLuali6s6tbWyF+IpQ
s+fD7bt8ghrKA/PsKgUne08ZME3YKnzlSGx1qorFniaXftq50yoql2Czs8GeSV8W
xnGl6aDFqkqtTAiA8NPHKugn+QGakIpNOIdzHEnDlc5HLEIQaRYsPBvAL8BFoiPr
sw9tEJYwI3cXvxt5gP2TyxUFDAvqZFfBjii6frrvsjCQfcMEo/co8cW7u6fzGoF1
RGU8Y/0LjWEqeUm79mraRtbXyScIQpaDLJLsLE4F9NJXsjYLWfx2CC438RJT3m1F
XuHsxisFbIxcY/WX99G0A1W7o9a/Ew9wa8hy3TKVdsrH5mwp8FAtCcBL0LEU9EcW
Zc3frxp9oVq84CkYSq2E+zXFfSFfOktl2pCPsshwzwOxryuj7a47SrgdHeEpm8ZE
Y0ZrDOl+Nb1qNDm9FsxJItHFJ+TJFjRCYTrCC+mJm2nNTxCKsDcMPuO3x+Y8evlq
eHciiWkJx6NF44JmyPwmppOfRqaAMxlK+/kFQhJAfctisknUnM3sLA/5eJ2UbngU
L8a8tA68WfrQrC3roxV4WtXghFwhbw5A1dx6VetzJUtdpJtAfApEv1WUshs+4Ehn
OxdMBQpRgTtYCgBAwkJ6tqjx4jEqvcblXY3VZRsKf8Pl/T2QXid21Z4TKNvS3Ef9
wFOcLx76mVYGReI8TofmU1crqDk92dBoV/+Fps3y0txRUhWaaS1gWSzy4YgyI0Sm
4kPXdWhPpPUJ7OhpFqVWww0lGOt2JTFqGLpc7ygxywRblL/2mLKb5TtAzlTX7DNK
1kFdd0+PoB0d1shuTr78o71GRDGvOXJZnWoSkAJ8Ks39CJrEUPUktLtmYvyIQ6+4
niaKjipgWezPHJhDeFalQWn9YfR0gXxUdi/f96bGDGjMPbqQnt5K48bFdrqZ8Vw0
mDf44Wr+JhaWGTkWPF5DleWqah4aPQlriakpeURJQ5Ufl8ZBy7yaAgC4nDuOcWMn
aai8PTaJWia08GTzj7citMrYBSKI0LecuRVC1iN0l+/NEiiWajuYJQejC2SplB8I
Ej8qrqGWouTZ4IgiQKplUSOEVQ/EpSN8L72jJNPC40WSU0FyJRsWm0oTQT7wVjew
7raa2X+2XAk6NH02KyswjvM5MFmYSgxD3CwUXUjwPIuI/NxrUzk/U/TYqf21wygI
rD/dY3FtpV6LLqu7+WFOq/94s0M2/KkQN+JmI9RVa800xK8aWd8yKqvLQzxbDz8A
hzq8L9fRgIWY6zEo2AbUI7dDEBAyuqCFFP3SmDfOkk8eOjV7GGQw9zGOJ/eeuoHf
DgPzPLlAVzC4E87x34vHuSY0i3occHA/JKSu/3cCAwIL2Jftj+1fN8XOww0TkuEk
TFxKixE+XZprd1m3zYVJpWztDNNcwVmFRWpSs7ggvP5Wwn9sd9ZSrlQOiXofHLrK
uQg2wQcngKQK53RAOAZLMx4OttoRAM8MA8H/STxbHWLu0E3z+OVCVvNgevOLg17v
BkpOeFSvzf/r9BhKCGJPnlyjkhVFJVVe31YZ1WuIoBeAjyJZ7tnocy1W97ECE3Tr
237sOT/+IuyR4PbPyWnPg2QN4J+P8SF5uOnlk70SS4RZjkd5BxzDvXMt2U+nhNez
MnCL/LLqI3dLmMa6uJWrokC9IXcXqFArkgevAQVOht2iD0W2HC68e5GMGfmJQOHG
ARUcpf4fTOpxDVBX9NVhnZwkWcvcgQF0WJ/S9+aFxzQzmYzd46FLtzevEiRuH66z
SQS/Cdx4/3TzM550bi3KGdIkpP5juw9+Zr5Gc7BxqBqwXB+um0y/Bwec8eQgv481
kRm9/klFVV2kfijfus7nxJM0hrWi9w1KdyrZhtwhEr22nzsww3vZh7v/wr0WZwA6
3IQJXaDLSLuYjoTrMUT6EmPsLzScGUDIw7c/M9qTdFsPNeKRlY6ouhYe2GxLqw3S
WNaSq1UfZAqhqacF5L2SJmy21VTlsGkprQAmaABozZiLLiwg+DGV2nO12VkyQIyP
nq7qL23lkDXeg3RuUfOpLNzbd8NgBhO9xbChqnRJxbjJPVTR6xLY1vQLMiVodhz4
Yne7DbI3fTglVGih7vB7BVFZfXo4aTb4th/lPU7CVPt+xiR639VwpaSrF1tnsryO
I94M5kjC87wHsTNOv0MJ2kLai3ClKXrLl0/DkwYFOeKi8huoYFjd+f2ZgSaxRJNL
gXKnYKBPQY5pbzzPw1sqGOVdoe1+aAVB31yWtFZbIG4s07P7LxPDo2K6sr4m4ewW
nxnupQ6ggVndPeMqjC1g9lCoTt42I6YD7FRSLQ5ZEoUFWO071kOb72IxDssCI6Fa
m4mV7oQ7emXGrmuKNn9piQW0ZQEVUwvFoKUnGzRs6gAbngBe6sqIAeROwmiN6r9Y
qVg6SSw4FQjO4b8PEHpsQixQNnUWGeoIIruP52B1LJ12SB+Yruvy0tYYVXO4AxBo
grfnIoNjIDvBUQ3PO19zV9l0lrZHdRB2HOnrM3ZW9zXZGa6mDMeQJcL4OONQ7+Zt
P5pWDAvUG4jrOXakC4YOkU+gUxRJYSuedMZ+QZ6B36nGCPNsu+Z1M/p78wKWO26q
cD6NY9QZSOVSUPCAEAu6e1N9iDRrdd5k3Mtb6835DWKP9+yeWhgHHeEsdoCBdOt6
iYJKIfDu4NRkfAImyTT/FhJRMQR4wmtcBxww5Pdg0HHPX3u/kF/LfSgLe14Wd4GO
7qgJ6RmfRdnkdpTKhIt9aAho02XKWKhb7d+mgXTeezym5mwu8IZp4BDhH6ncQ9pk
Y+hWQ+aXqz7oKoRAhJCoWa9Yig9KmO3K8ERpBBHgpb6cfn4LyC5nV4zk5Hs/WZPl
o335uHz7nFI5gBKIE3FNjgBIllxq0VZg9DxAt8RcebTFDhpsicI1E3gXysuIIOU6
/3tpKGGq/GDITO7sbhgGjcaIeaPJnBd4ZgeciAcOPM8OmVB20+sTwvYDodaEPV8a
SD0pBZmRMJ8jsdj4dW+WgabTZGL8AOSmdZuIB/6Peqf5nonJXuno7pruw3tjvI11
ZCDaQNTdDjtlAms3TMT9sJ0Y3jVp+5f0adMXQ3Z6k3BO1Mtzj+UuVQR9Iu9TgR14
UEzqQDYcIsfjzXcH6rbc+7uCiBG8u96ewC/UahQ8O8YTAIYSzFxjkGtwsdkjduut
2PBYL9a+Y456FioOccBOXGCMJuuWmsGQH4bz6cfgSB/hc1ZILojnm7o1NJftVt4c
ahdTDrBXTZmkdZZ0iPUcnfCZ6oRJZq9hYlT8YLRIvcjr5gALD2UC7Gr/ILgA999s
SH2RpVZDny7RRMJTyOKH0g2jI3nip4vHdsawjK8yKTz7+PXSUJ5EN0aJli/azzQY
04bb4rh11zHyeuHC5EzhhoKYGcbzRKfPeqV7vQdgLLzVCDV3cuAxM4d15peaIxnh
z9sTYqiLw0i+S40iw7o3Qd6+wV3P3eF9/dm6G7BzTPrCvlN8sqsCu5Pml/voSnob
F5x41GkTnJzW1eRMhwquU9ZzDNc2oru4f1GpSsbQu/7vPCD+MoECHLKVkDLeLLFk
TLXmMs24eMERa9k9w1oxFTXb+T4d5ovpce4gXGiSM+dK035/gr01LZ4cFKuWzZiI
Q13U4kD1hNqOtCxpPR47MFjlSnqOHk1cgBz7AVEdq/2uKb53UrMLHst7TfB0Usi6
xw7RCJvBqi0brf+KnCxuB66K5KmJJQAA5lpa+dgqb3P3cXud9h1oayhGaX6K9TL5
JjKt1KZ4sM/Qz8d/5x9NbNDOk1aF7oZ/wJeiv1oy562kWGNM+IOaxYvry64joM3N
bSZ5vEernzScY21CoW2sSFCyj8E5+LY1MU4BEZS3Y/8M4hIkksFd/gSh+752mPdn
tuVSWQ77hP+umLmOe88gilZDkMzDQzWklmaMpJ6Rmlmy5RSnLVLVUdgF5qzGVdRq
WiNlAafdrAiWZKA2dFKClK/675Szzz3KgXxjuMMaCMclBUg9/iAFH4JqWBjb0fDR
2kTKQDu/864OuqIPr898cHUD3J7lboWzfRbHJUa3hz2lylFw3hUJmh+H6Tda1Xtn
WwK6YjJKAMYLjfsnF5Fmnlh4w39P8pHIfvRAa9Q30IOqyT8/GWBXQNoZC+3wE7a4
UeOZpuUosdIvMTMt+VzGmbNl+1t1vTKXQIinH+c9Ny7aldJZ+Q6SjeRJ/e4yVx3D
DPRIMFfWiQ+LoSYfBIXhuVQGSbWYpmj/nqN3Nabp2HNVxh3c4mLsq2hWq3zkoF03
x07xuJi+TWZpuOk2wwgrfjTyXgzXJkAoXyvbcZHy562WRIl1tBif2Yf5CLln0A0M
v4ERe3ONhInqx154brL6UcrWfUnnUH2P8Jmyvp+DqG0c8hSLskmWKbtLxoAenw4y
XoeLyqvEX7+o6NAej+SxNKoi5x9g4WcbU4rjm7IJMg8OTSAAsjv5vS23V1nZmkR3
hlSX2H5Abuixa8RWM+nVNywPmQ/scjq7j8vtMYPvA3KGBEKYBHqKgVqnJb3o7VqM
W2KpJhGRtagkjrvbxtEurHkN9Zg01IDg9ZoBXx85S2FWcjBC2S3JJ3fSAjlF8AjW
X2FfJRiO3IePoSh07TNI/wcAtsQ8SjF/4bSgaXapcpgpC7vOrNx1ensbF7Ugs1Ea
ChrB3owyw+J+bLjFf/bmyvnzhURu+FX7q5WCeXmdydDxrjm3WO8NL9c25Fvb4riq
7pMZW03dNrpVBtzdDxLpXYzBQ4h3qS9JekKLle0CLJ/cjJPtI39Z48RkPFgJQuIa
69AFQQ3yeAiJqX1Gt94x/8YRYmWz5S+7JUxFGohzq6GeFIvhNoQewyw7wI7glacj
q3zeQYIqm37DVykq0xbfjZYwYDI5ofUclwH1Q+XWrB8jetBlDMUY4Hufu47xD6fe
I1D0B4ZDtR5bJWdE3mMCefhGR5wEDjb0DVex588KpYxbuELb2rvmO5ZE2a488y/F
+zLbWdkSy5Rw+4WKYY4Soq5uqnISFmIfEDQxU2ChCbKhgC3CWJkxueotj0XUSWw5
jDUaUL9yrGAjYPX2k45vaYwc9lH5pztnTEe0RLL7Z7mQ8+zRnLZ9m9dQeaFFT7e1
Tr6INNDaUWpLxMz0sfenFbYb9UWBmkdleinmMoJJI1ITl/n2VA0GrzsdLIEBq9TZ
pl7fMhZUNw1vNOGDOWQqaKJjOI3qOrjtM3Ix/+zYRSExbTfXeRIWKM3S/Mtkxm1j
yoS7bFaM99xo8kOlyT5AeAXjNk5KKzrSa0r0jKSoxn248VrlwR+k+z2FOjgoWv4X
D/ysoqx5NqXXUh35uh/43dGoooFB+5UFz+SX2mzPU4Nf2XW6ar2PiS6kk/ZLjjkw
NdFJKHmNwabYQ+vo3SISRRXHe2IsRMF9vJ5dVgJS8Zm/hkN6TPQnyiAOPiRLQH+H
O83Hp/o5Cs1B/wGkfG7RqpRuNwz+i5hgLFH4FaA3faQvsjhjUU4g5OeGlTMRxtHM
Pd/fY5rccvsu2aLGU6VtlA81G/Q1upjgOhhMtHNSguFuG9sMooj8QDSYDoJlUyTl
zTe/r1X2U57ma75HAsGpSfO54nG99y8bpyI+ahGUbdYIonDEWld5QhoGde1j7agr
ChrauGz8cyEoMb8zbce9T8f/Of4mZ+dHorAwTsB1tgsavztrL84JlNnUvvbxJswo
wTq3B5uWAot2iQV7eTM6tO3MdVietvFu42VahhRBNA5VwFqu+QetrOOYER9+V7Ed
dq6mnReLmbJ385E4WXYONUwM1VAK3YyHCyS6G9bx4DMe9JIkUaAUz7KCw26+z3qz
e6Lnlt34ZzPpSMS2HAzQ3nQetnM4a5wMKFj9qzRxHa70aPV5XjAI/NBjTMxgy39g
B3oFnn519z2O65J/ws3Vg/PFDbB1iusio/0h9FcmCWVVLQTqSTFwE2QPH4S9fpLc
/XvaHeFDwLmRt5RqKW5Xf1Gbb0y53TsqqHhSKcyFTDM6jNNHHu4MQg3DsCtA2cBm
3FPgQWbPV2y38g4dW0zas8udyIaCPBRXxrgTC0LWG5slcE9Ksw9u/cWZNBfMFR3g
I7Fv6csO37TKmXwYn7irlPaDauwpEbNNewSEc9TiQt331tFcvKGWw7NQDNc1NLF/
198+DFdDzrlkg/LfT+LLJEfc5Z7Uq7HQEp4b7z4XYSQpV1DEh3NYcGPGaFf3wJe6
+dWUuo43XO7j2iwsOESZld2FHaTdcLu29VOd2Oa1b8PWtFV5tpO8pmbG4/y2uwIs
TR2bXKKwtCNSvOr5jmypW+k9JvfoOZng0Dg3lKOEe/B+EpqiuRFEFOTVy4rgHK18
lo0bu3YItE3coBxWMxe7pnEgiexleo1PtUc68oSRvEdoCwV9x7up9Oi04ousjG4S
nIaCPmISbCVCOzMd+Yi9nHOEE40AtRgkJf6WB61PU36ifFEJtvtjlbh6yVLnbkbD
pmstMP1g7NQVbo5Agu1VDFg3wmnOJfxqGkCD5/gkOPXmSWuJqhYiSWil68KYmQtB
KWX9T4e5tsmox8/Drohmnzr2/9O305Fm29YzggSDuYXVBusBt748MCdE5c12+HWp
Answ4BaJ+43Sn/jZHHstfQ1u8tr/M+R//qwoN8JJ8eYZ7jqben2VPeUbE1EczvFb
msJpsEmOoh4fKvjbvbY9ZjYWJ/huFvAGVAUrFhsq3fLtupC9C95NJPaXET9bdU27
DDyNXmRikjmP/9xgon21usDNyXTNRxdfqcw0Ct9LOT3uuJOYWiv+bfN0pykYKVAA
Tz1q9dAVywh53EvsfDe/uD7XTBxcXbSLHDoMRAjRnVPFnbLNvKwegcrVeVUkWIN7
hLwdLUA2DoiIIUFtgKmG7s8V99rOXj2jXYCqCbJcvl50yoXckuzYFwP9MZcETzXI
eDi+m36gM7kRQUv07mPaoUrXmgI5b9CRTmrYFkMbEzUIMuYIokLHpLGiIcigvxJn
1WgPtuQ5/rxTj+iYFt1LW8eqnXH8omDEnNAJ0pXarZ5Zb1RX/FTzX+fh5P+P3cl6
UNOAw7VlQR/GzBdL71SozyhOxMm4+jEcL7EEtLytHXP5XNvzGU2BJljdU6gW2reN
yyDEjX/XMrK+KhBBzGFHOM5FY0o1z9Sx1kQbKrKH8xSwOh1XktA5F6QTaoL3bEZL
3ADpKbsTYehDWDWd1jbAqvQiXulXNE83UUXt2p/Y36a+REO1QpycLCLxAwya8g2v
AL3OdXz2bEKNwEvQushpYqgs+MMsczmc/jn+SzKSArX7sEB3za8WFSBIk/s5zc5Z
VnUY9K02qGw0tDzkxpE1evqVOkAMw1eM2eAajnqR2SuhNwu0PD96H2278zoV2m45
PfXz0uTRd6sAqBUBMxMJU934UfI6Ges1fbDW50PtZOEKP+Ki5Qt+edrbq3M4mQtu
3GGGwMM6ZZO5astAT0jgqHGEx9cI2y55ap5fn/RGcPCtl/6OofEClr68NHJL5+Hx
BGNur1MyVGdSrcYFgJHR0TqUjYp/xsNWjMpQwefdTGbVhsQjIlFkRW/y7eRjSyqH
N/qyfkXjfWe/69NKCjICr1VP1Tj5ZyIPHacXb8BPzfEc+wXfVtWW8yQ7IgoBnwzU
C3/GaY8iQ1G7LIehjsFMTyDfr0N6eHng9v0WPbZXsnFJSbm0R0Tye1+Kg5gPckmU
imPsDBs58Ynm8+v+F/tBFq0K4XFJXzaB2SlR4OfjXSJlw8WZbJRl19Pt2/GLRMrI
K/Ej1WGZVLLO/xDJuilCxjlOHWg+s9WHbQ2ZsSVXk39k+ZMLa9Z/NNGUioCWQ53V
wql/sIssUqkuSJowdKevZeSh6r4EnBjhZPYGt7sVji0AyS/XKNyEcFt6Mj2bK7nR
D1swQkOc5WSHHvoJiOSvZTrMt1QT6dlBzbuTmBJjuQKy0QK2GXowh6RhzozjhCQ6
k5K+dIt3H+nGARIW2ZHGP1ax+E1o/59IK0138gUZRTwu1uj0dzHL45dcH/WaQPnq
+A6Qi0qj/xUbxOaib18ff8RC4Zv4W9YyJ9QxbAN7mFlfcKX+qjmc8IkXv93ILVkH
Wqdye597VHOF3v2WdwhRkkJpI01OkWioX3r/j5d2xSvvJiE/0WAHx3iNKV7gBMuw
BHHUUNCdkUYDLjg43N0nEcal1P+tGkOzLpY5ZBeCsCiaD+aRx9TzIY3ilTyJBZHw
iMDaTrEaCh5WHbvoRbDSChN6oyM4wB3jCgLP5N6ZheOnIU8BhL74sRgSnTYbsrBs
tc8llpESjADnNinQm0112BzaNS3daxZHj8cfh2p947JB/4XJ+Inm6Us9BZ3GxRna
z03eR0DM7r43LPzcZKmD/s1YBJtujCR94Nsv7MhkIfSje/9KWdwOWN5GezGqXHYk
rij/rBiy6fPeDVNXFwNLjfYpRU99gn+JZID2gIgnku+PMMW2cg/dMNpg51pWVgTE
ka2NUgQaS0r/XIHF7gzt2coEbyuNdL7DBjyRFpiM3ULe3hrL7A5SyEoz159WRISd
uy3jT8zADldVjXsPt0n5RLGkrwECmER1c4WsvbIXYxrgNvTRoPJGlYo9g3jHr/cE
6yCjpoIQUse2X9EdselAtKuQd2MqqGFj7ZhwvTXkcLUjKqfpn5Mz5Y9aPggjmAwz
FaQKKpuyylHf0sZZSFXTmdYLwpC7n4RsgVMkN6Ur8hW2ozUWgxezKW9ufuZMb9oc
WmbepfBTEHOUUlJjVr9KayUBvGr9+owWVQyuH8jB0A/AMQnVqayTjtnKrETS9KU+
UAL19osxib/SdN8SWmps1JnxQERg3gnPVah0FVePD4aBjsxNeaynnTSqQ6B930T9
j+rZWge1QT3h0T8lBYiNxxKi8+mKCJQZsRZKEthEb7xU118sTijl4NSoEpGxumf0
hrddzl3GcPAcrQxzVaSZbC/9HL47kVOwGBdknHDlxuUvRz8XZYTGqcjjviIyXi4Y
pGYveeYMig44eE9mCX+GEZQtxhBSTr3JOC9R0ptQMJ6roXCT3k4Sbe1OQZoil41v
ykh8NEBsFD9VJRADjCQ9jdTOBoK4KCfR1qwyYAPjktJWYPgDExmI7SiKyoA/gyQe
u1SN/OnhCF0a54tRwe83HQkARbqFLEbz0enTOmIoGshIpYqLzcRAChUsoxjH2KMg
D5ZoRiHx70rmfpiIAyVJ6wv8j5zFYUJIEBDhJ2jflGsX0Frf3JPBH8GKTck+dxsv
GnZaLx5NewOi9yondLh8dS5sH6OxQSTc+T7Ie0txDoo9UKb5OGwVKVjAFLIc2gBi
ibR0f4r+ZqNBE+SgG8SXVDsz5tmUsFtrnao/OLLQ4EBW+QSkwE789JcFZ1PxlJEw
3V7nBWo8UNlIK8KOTsAHHqofYa2dL+WRwzZTgWA03OWXYmOI80KT3Xhus7bKzdZ8
c8CAggt4DVXTxYbk6pFzFRtSGxNKpIveA489eCozzE6fF39HZrzLZO4i6t62WRYX
9LLr1DdQm8m+EydtR0rDVMK6yRCGReOZfDmpukAFIJxTXhv9rHjoBmoJ2iVYj5Om
7LTc+cgkOjb6OPiwaFI2PxYAVqpJHM9ZRYogAD6vF204WWyn9PcW+ZnVrp5t5bSf
kVsAC133CF91NN+dXsx/+VNJz7sdt3br6rkDL6RHUSvuGcASH9bbUVy7U7ydOOnD
fgq0uac6hLXyheG4Zqp7L1tTF1S5c/NSk0NPnmyidn83sFtueNGnQ+658UXo/jE7
BStTlvckbk9q6pO3JKODO8EokT2x8qCt8gcKVTAV9MUVRCecoQwrMEY2xim2FHkl
2t6WDRmmSTAE+BU5kCtEvIBCsi4Ai7zTXBi/23Bk7B0IXRBseLKlWXI4/mgq1fKS
aRJv7zqjg0P0Mzj+QH46kxq8xHlIgd2eo2M91oPcGcQUWIohITVD4yw2FUzn2D4T
LU/jy6Viyb3+HFEaYBC9vjgbhdpoVw1nTUevZqO+IoDoLX1RRf+wMvAyMzWxss8Y
hOWDQvA9zprmCptOcT22xFYoZjIDPRZ5eQUmni7506pt2oV13grqNhsvfwvVpfrX
zU2CJ8I8QNOTXdB98S01wVTX38Gr9QWjxW9GiUQz7wSbhaAdaCp1b/2L0TFDv/Q7
reUId/TfH9lxOfmyMS9zJnGYI0N0D3dKzJLhv9pQ2DE8CDYkxPKcWM5k21/4GJRA
Z1rhbdT0h7Dp66JbTqxnLIfsM3xPVZFxoWvddJEvpc1xa0QJ/69w/Bbowif6Ny3z
kqYb0phk2vczFM3DFhGkN5HFOesYjtV3qgeFmyxLDodUG06KkTCaB/GmshFzJiFx
Xa+nghgftmkf8lzu3kTgioW3umD9cH4ifcWUGzN3yLLrgofiBfG5bwYhrn6wkqEb
Y4ZYNDtaMx/XAgv/6v9qKRGKA5vVTgPdoqVzsq9wYCfHGIhJ4pUUiIqi/5hTVpxp
nK/Acnhg2nwY/AbLYXLlwnEgThJHhPrm0VRYV5uXrwdYCE396hWEsHBftIuFkCa7
gHO117WUPprOifqtXigwsesdCmZDWnF8eCtpPqaNbnRjMXtpAJUa+ifAwB7mrvMH
YZ/uFjWgaWGcn6c7UZrP8/l52O/RxA1uzXB5vClvnd2XIWA25kZoBSHZrlIvFcSr
DaNo+jCF1g4v2oO85Nyp5y/kmNTJELnAn5euQOWwdZ0glt0D6rnBej7+btebRQz0
hnRSC7N3Cd5JAYqf1yoIcxyTAJ3hQvL+wdBejiRLJfdJmN/txkaPFAidbxthoJTs
I/hpoRxrcHOLRiFn5tdmPrsgpUStuj5JGCv/40o0se+CfFvZZn7Eh5sx7J8U5vxG
kpkksjVA+pK//1wXgHrOWw2L5vt1jYNsj1FS92bxX4jqFr9/RnT6yZ4aNh6ntKwV
fjMR1NqsZpoG2DG0zIw41sG+BJR6kSBeMJN+Jutoo4IzOQcwgu4AHUGtP94TLZkf
KGA/lWpwUKqFUmeyYVe1ylzYZBMDPrxeX3mJP9EBaTNwlQaTxWAvrDxDmZYMPSUR
ZanRLBqI4FVYhu4oaBDyRKyx9WqvIn6wI/uALiiML7Zp+EKmuoWXMFFseck/aPEk
PW45wqNREBl5AbPkLN4MumZ344Hafdcv7DyKvtzHoxKya6yL4WRlc3s+7TT0Qpsc
jm+SW+2R3I/i64CqCGtJqkjk7RMhPQCQgezz5nD8JSdz2/g8HzYZThpLkc2okJ4A
xS/ntRiC33FIo+LgGlGJxbHSA2D5LmWXX33oGovDmHdriZxl/Fvdq8Al7YYPKcdz
Dr6eDAKXYcxFlynpRNB8AZflVAW+wILvZ6cap2/Ey2+t7wkNlg32B/LSXwfkIqU3
gOyVGKx0n3xaab5I0cmWcrJQpB8nKE2mAsHyHHK2fGnx3DopeA2pK3RTvCdt8h9V
M+ZFeL2TlPJ2Jdn6XY2RCs60GaeS++vmIXHhtlylx/uPxgXakwxCIwNVVKDzIuo7
xLuP6wWyePHLx+M2+qiIoPG/Z4BeN73MWKCuS3vQC5yb3JpExsP7CtagfBpPdEEp
XuGDTNIFH5Me3icDJRCm80foLvKIxdmz0c4IDAW0TIbpOWi0BIDVS9UtalPAPQZp
OgWTuLEKTSvS7knctMqwK1PXsBSyK99gCC1kj1Vsh67A/IygSaSEHs4O0eRfv1ft
QAs3+3bi8EYglITJr3rHSrM91smr7hggw5ATbZhXRTo/XJmwRPxcwf/oK1JNwV5T
SwcRL+KrLNmmGsUPNbwk8/x1V0d/ZL815Zd7+9s1K6UIcozJslC+pUuavh/cGmT7
rGj7o7HYds5ICegQKS1b1wQp4F9QX4mOxKxpxGWJ/cxVcrXbkju+nu4t3fDqHrXy
wK7Dupfwn9j23vJChmk7g7kvsOxKj7+uBhnf+lcR0HNjNwwPKk0KE6i7JA23i4/V
yO+eHkyzqyVhYw3txgQrtpmfdas33sq7sL6rx8WivSm31TUfQ3cGuF742K4TtKv5
8FpCn6QeVDqxGwl7/FXJNmkbV6lCPJWCfmjeFp2O/b/OcXef0JNyCtoTHDkFJpw+
Up8r3u2+TmOZf2modHtXyJOSGzhI95ACl2LW3WFyfcIn6pGXffpqD5g3cH0vQ3Xe
4XcQbbuVMtheVl5ZFKeFNjcgK9LI55mlQJIKcWXVQBvyLPE+CcXkS1RBsXlA+7/Q
SlPUX2wlCtwD84zbDMu2v5RglZYXjy7G8ldukAv7QMA3vuVgDaTj9rX+osRsVsGL
a+AJpwW5JT76Xvq59eseUYufab8Uhx0OwtBpkqP6hWv9otz/FZEvJKihCDuLAcKx
w/mtFbWbKkpoheX6d9lcU500DninXtCO9uB9tnFvaflLIqxU4o1THySumLPKi1ni
943ZScxnKECxGAgH9PAzATZG6B4GtayW5GSvbDeZ/c/jpyA3iAlsObBjIkR3piLZ
L4HdQtB9tdub5bwrJMgHcABKDxZNExuHrDvnU6XoPAoQ4Ziox9uL6vuQxXPamQZF
SEgngBjZU+tX/3CfPicV7gTx/tHLd9A0+7JwPQTjU/y6Zvt+3EL9X7rhFBhujOcD
V+b4tpBMP4ZPR8ue//ULVF6ea7jzvq3oP3Km3ZiMk+ZgkenhuXmp9Y+2l39bAW8r
gu6Vgwfvzu7xzVPdZtqgeEPM8eugYGotD97L/A3zhGdX47Ldg61Iqx7icfxCtY9J
UNlzT+MyxJhrDs4OrkRVe5Zkv4JwEYF5TEZIVP7QSq1bao2ChjT4WyNU63d4Dep2
pCGak1nu0KHKfBHl6s3D70cN18ApIrTncf/HBcc3EAalwkq7N8czVSqlDi9jGTFb
3rd5jpJSKmZRhDG8j0ZCbzd+9ga/sEGJK3cJSO04JpVeBTyx1NnSR3fX/G/ZN7uL
XFqGjatsnO3M7sR5SL8jU/I2xemH+l1Dio9AN4AZnTV8AwaKqZr5LJsqRNdt9crP
SZohtVGIHzJsplD2fTxC3JL+b0iIDNNeztMCmJtK8uOp1+8PwX29J/X8AxN6QtKQ
pc5nSUy4m/sJxygbQJnlT4NYX7r/4GKVyj76bJDoa0/oSPP0CsAL240Mdc/ZhKA4
LxPvVeKIa89kjyak2gmuqBRQxNUBD1OxpxaG8NZksNyOM+mSQ704vxvOsIyBvQX1
yJm0ocDo2j7MnWUVQI2uhTwGlwTrgE6EaLId1qLAQXHWReNuoW4My+jHQ3Vr9B2l
Tox4ckLnaOz31/YCafkquE6ITs7VyCtU6usnHMi8bgTQzqGtgUlOHq8gZlcFGr4b
YenBn+8dtE2sj2SJgEn5bnVs9MuswX6XtmJ6FcAa6+NC/bWlwcPt2y0N6fpdKjRL
/9ljGiEVNSFhGBKCWVPK+WaXzRUtUVkL4HmbOKCOa0YpPxyDWeVeoMeVCYFUDODi
waUjyyuWP83+TTGt6hprigiPAxbIy8l8echxHwYMtfNKAS8F6euUjh1WRZIohs94
//GpHVQjoWAZsqIaHVT37m6D5lpU0ZzMVGTNY4m+QYbEDiN81MjBzfXkD1+H+aJ9
CbVrKJY9Z6HMBsWzuqA5AwjFmIScnLJsP9ljnO9u7QIoH2/SR5VME7mkFAG0MZYN
1mItEf7CFOadZmOd0Tr2hed4/2muysHWfq7qeHXPydQmmFe3Lvqkt+ZkwUvm9GSq
EfXF+g3Lw7v/Q6SD9Aix8GzXACGSXFusU11KnjdAITcOLnuUU7aqzCAqpMPzkghk
+/EW36qUgUH4wBbkG9dF/Q7SyjcDroGB4yHLiFyrnPQIB24CXAJjOf0dhGJcEh0B
2/axL07inyIuyVFmiOiM13lbRCYNh8LFfYmRwYWv3Jly9AZVtFDE/wfxSg5qBSwL
mOTkoy26r09nfNIIU6KlwX1zXJTurwPeV7vHGZJ1t6D2mnBXafVRjN8zg8EnB01L
1JQX5tAwMEOdMUIwV1mtHKUQr6MLnqMDK/lGkwsmBvdWwOHwaLuHSK8oOdEEac2E
HWwGZClLjApRNSfaamiB9yKc9pmqwVh1WTqS/ep5Yl/j5aDVRVCOuyVM2KpREDpA
mYJWE/raodfkzbBvqZLG2cZow13rHin/Ep2d1dcSJmBobTWmzLyxTWKGoVxjxqyb
jfUZv7VbXR3+uEopCD1A1GdOHDIM2007ycKAXNErJ81wT63o/RivhGLjlSwo8yv5
UnQBRHxfcR8rVeVkS+bAJOY3k5P7u3k35dwBLaRUfBWI8p1xrGl2ZoEGE8G0f3+a
2lzy1XL2piMMqYIn71azR2XpjyiQiK3Q8xmdsZ4rKIQ6do7nTO3ZpO3WORDZd0uu
f7jJrhyH3p1lyX0d1KSIlsimNBm5WCegyWWPJdwT4y3KFh4d0uiE/Uy4zhc7YlVE
xaSUpKR+VSj39n4xfDdhxFo1tWAGYaWm3xEF2aw+Z77+7oxVw28UgTseHQSZZlti
NJdr8g88ctt+hJsAB/hWlOxpwKHlAP/l420Ifi/5yi3icoXlY+fbCAo+1vfmsXqQ
oU3dxlQF34WaczGircjfedfeYCP8gLIuV3k+FB8W19Z49WwYR1rBBekod0IaXqm1
zMCnMx8MUVPnVASjSOOiZqk5uNp2PH0AxbyXIvv4nEb9rxtkd2kaZ8jRY97f72kl
drVQqLrWkhf0Wv17ij99LR+y+dz/ZjSBII9Evo8pj8FHizq5CrRfzOP3g5upnJqb
kt7txUroDGfpKObcHkRpFjRQBWrxQFi5Rce0om+Uocq1oG+zrrXcQmGjmmbcZHdx
nNGR7JdVm3wVLqCvMhcyu1tMGjQY4l14cbu86yrBFtEggd2HiXoZufrCMAc0N+fh
ry4cP1+sFDbGVpZ4wCR7MXvTjCqpQvo3WkEIgruaMtdIWzES3kZNk1bB0eQPt35y
wxWAFYsi6SlkyHPY86vnMJWGq2VNu3loddk7ebxVua6cGdOKdOQBzcaUT8nS2tVS
YgByh32YEMBdBs5ggqetxk9H1BYDe3VZgqjwwvepuD7h4hfiHF+bjrhbnHI496CU
B+vuBWo9Phu68IzhJgrppuc3yNlOY5o6NMrVOyAdwB1/pPqVPiRFBbATMUtpeToh
Kg7PMTUp5Qpl46jtpS4aHTZhBdGE9ZodsFnGZfSOGp7Kk3fAWtD2F9MO8SDbV3tu
4RmQ7JPNGbsninOway18fGhVgYqxiMOnOCnt7/QT4ykJQu+8ycCIrrVMIRFDyo6T
elLPgxbT16XYPIvKA5XITPcbYURiqQZIvDAW3qtqC1O/7EsLnke1fWOIaaT+xFYJ
BNMq/aIW6TzJZqvLDTVV0IgxjRr8F26VWMCH0wUDFl6kTaMiGYoS4g0KavR1wmX8
4ND8Q34txFdsQISGU44gEPWKUuBIbBB4Y1Ordct2n1Rlt5SbzQQp/zg8LI9VH/+V
MSq2SpezWxYrK6hAA/Ctu1P0+HjLyhpYO+sE26ztlQqNJ132Sl6hHkUwmUWlZpCI
fA5BdJmYEKbTSLaUv+wYz13gFr+bAVJi9Bcifyg0HzetQhijPurb1G1/lQEbcS/D
RCbVhknwHFS4LnNW9CQ08U1ow5DP+qvNCSUjQOjLLGQyNCGgNeBoz+mm0fbj4+hY
H5VnCONQPxmkbHc6at3KOXqU+6q40BrtQWMjv3Ax3FFrWQUtI1LlQHVZa5sABG9m
bRDi22O99TlnusGb9Vb5HwxXJOCgQ6EINeH+UJPGoRfsEV+4nCSq3wEfCqVa5VQ0
tQOyTdgpFEJv1SJd71ppQIt7+hS33MPMyytC26k7xy9RwfFHuU84ujKLVf8B9Mbg
9UEzLZ/wcHkXAISxD0uLbUfJniz1P2IE1sqVrk+q5DiilARIIJ57DSeq5y3j2W5u
qXjGLUab717Ty9kBM5LljpgdVkYTumtGluPfINUGuAXq/xzdkl9nJu04VMJRUPqH
Mi9JOx71qwTXQudP+433nF9TGeCPVLWrLvRMSu0va+UD8FTTmanxcFNgPObJ/X9j
0s2bVP0euZNOdDany22EZs2P3jys/syVmO8Tk+GtMYeF59CA6ko9L100vh5mtKRA
uOw/36o627V9eN92z5JfZyPFdvI+qmNUNxFJOy0e3ErkM2lul2DknfgovdpSmX+D
MBiQSu3i4iPi/rr5RdHc9gHsY7djiixNx54uVD0WIaINhBI4UlUUa6V2Tkn/2K+O
uHpRgneSLi/gO3KrWKHqQ6m8slnbvXr5HfOjoNGLUjmfx5IR+OA5FSZkPHUxRug4
EUXuKiNPA32V1KIArg6eM2qqClnFdv4yrm3vLEA73jlPoBK2gF24I2fHd5jdgqak
EfmV0RzI2XmxCVfEwGjwh39wspMj8zvwoupE7eWYLbnbDRqNr1LjSM2FuTWziIFQ
o6kPRol17WVqLeCfPwrZMVQfijw4RileWCtzuMwdIeAOaBi7aQT8QNsI3hdqqneh
1BTdGqPNvkf9+l4O9g6H/Zx1z8Qjx2zEcB+TLeF+1rDCcdh2J9RXyatzzrWZpL/a
MK4cK5cCsyrw5CU8R4Nu5AueLVNEYnsoBY1lGOqFnVs8ALIELPXQRJhGDMHPshGp
19ve1CdBDkCTGwNp9zbuWJjARJAjzCNGxezKWRaneGAjZVsRN8y+AhC++H/on7L4
t8uVZN8AcW9jfdmHqUyREFZTACNXDyXaIa1w6Oc3rcej2zi3MdmVNMZscECO7hNu
SMdGrDtX+JQYzow/+7iG8WfBnd8qOmnNbjU42OW6T39ZdpJ6PKLSumWDbi0bsAJA
ud+FF94IlModsmneM+I69Xj/1CQDY5rDZL802mIuE4XqKYvPcIe9rF7f2h6IJPn6
3vkknJtfZ2GyxzT7mK5WvK5se1j9irkIxSHxD234NaU/++HH+/YI5mXtGk6U84o5
gnxz2KMLCIUQfQPIi2xpyfzBRmy0nbpE+/XZxgo6ju6MNClMvlYe3gtJU0mPBNsn
CgGK7Tk2cxL+LmvflNdWOeY0Hxzes+slnYqljbQAwT26m/OIIwO70q5ZwOngvj1W
0/2yzjuFrt2bLh8b3+rjyWpoqjNvt9rN427jOwTBPW6iDNppHfMAkrXFidZdUhvz
cE9OykZ4M49veqDlVuvGuUvqeYIL058/j5FMtFcIatNwWC2KJAWwiN+qDhDLkrly
Dz1fKJ5DUGvvSqhfYobgHeB+oUgK8G/C6AvHNVWksWb2a7BEsoqyCjSwL/nkQMZZ
RcGRJA2caYF6GQOpbFIghoZhn8Rpa2lFsDu8As/cloyH7cZbHj7762tYL9oFbG7U
K+3OmfRObI6/HBDcux9UyQUQ6LzeXERzG1yPF9993rcHrMtWaNa5nfGdu4d4jxPg
EQ1adZMiCmPg7cMQzPyq4ZX9tYHj2pWP5BG7VvWdLPvOZQ2Uims21+xylglY/T/e
X3NfIapsZHLFKlgWdiX+YAlEW6YDoIz39/+ogygYWK04Iyb7lpYM1sfMUuaDyc9Z
YZtFT+JS/No/1hpefujowLtvp53/1wq8MdaHhykkdo/Z4mvisOuxNx/43+DxdNpx
5A1G3YID39KKfEnvpHL5GPJyHBTEWisfr3qM4LOG29kzjBL6MLq8dznRPXjSQzK0
vEBQmn2/rGwJyEUemiCMFhdY9GHPU36FhktTH4Nab75HG8I0mbmdeUl7Cg4kk49l
VSK3LUz8cO8Mxchl4Gbkcw5j9LA8NDKVMuIXgbGrvTydCZyouFilYzWnXAZCX5Zo
0HkyzxiNWHp1x6raWe3WtzjKJqybxQ4kwG8fTAxD0PqJ/Y9LGndihiKXPVrD+GPp
UFCB6XQiGuZj67rKSZluQHL3WUFdconPYchlum6Vxyca/tL1lHeHHTjDAeVlCEr5
bXl8umDdiSCLXDAZL3eycge7e/plusBSyiuC8tcyK3wD8hYvrEXF3fQrrvaVkK3U
fDVTejXipjWynYzmXzmMyzvBK5aezZhPyS6/be4bsUC3AK4Lua6YzRrKnSO22u22
cIKmGnU5WdveeE55sx3tts2XgPixLWMBkJFVYAoTKZplYerqtC1fyTYbt7wPq6Z2
RRiDuLUI0qR/X+8/EYV0CqHbL1KlrTLwuXgOVw55KGuCnyk3xSEcCioJX81+rIZp
HRc7pZy8/5Ny7mSL4cS3uKS2lUvB0/+wl1GwFMWyLUcn/GEMhPd6Ti0yz+y3N9qy
JXzBbe0lVlHnqAYFw6u4sHnc8ei9ErMW445riT+7fpzxF6hkuRI6aG0xhiDJgbAm
fhghd/X7Nac4vzMoNTgn4hr1FwSkNYlSQhVRrOMZAZxwuRCgdxZW4bdyfJ4q53jA
JhDnwwsjk3Kn9jfSNE4RqT++aH2/Nu53iKeHYhBl97eAKxtj7Yxd7o6GMiZbQV8P
VBxpaDiXNXo6N1SPY9ubVWM0KFOH5mRiPJFUy2Pb4iSdRY1FTpXmqhDSowGwK9fp
GMTcHY9WbVDGeY2ryf2v5tiUUDlr9dP0S1alLlvKHcCABgSsJ/6KvkRIMld3Hyjl
l9gTJbPsUSm2G8zVUFCihDgrwgCgv4exmcKxBDSwVZlpJNMCtkxAEZHMj8aRhKyA
QLlU1wHYp3LCcrcawv83xJ20V6REO6H0kRq94bH+2PBGP5Ic4nbBfmtK3pexp6pD
IiNFXtHEqLo1Wk28W6COo6zneXMZlAlNKTfMNY6yURVvxoc7DoF7RUIx5RVjAU3Y
94SDOPpTdzfs7adRMH8abh8WJWQnKYfcwrA/SeTHQrD+5hS+q7L9L3kW/J+BNZy3
7BUYPT4DNjMTZL3VoQnuWng/UDWbVWkxSuvFUrVWdh2voe0w7s4lcgPbsixbk7QB
OSFqBhkzxv/ryQ9dgCGrXgoeEM1SR4e/IXDZFDUdhidd6WHjZZkJ9sM+4yvRHRKY
+7bdJ1jjtR2XrcXYL4Cb121sIClIS/6VdwONJ3zSc+NqZw7BkmutQmUJ7OmRklBM
kh8Ld+a31dHvjJcG64dh7ki4I43i/m2/NzHb2mcsCKx3naimeQgHY8PqP8vYpmNe
Cehx2jbbxHXl8LKApcHB5INbcoz/uuvtgMHabPQXc+mmt8RWkb1klhAEtfmnAmkD
s3TGTEMmXoqBA0oz5thikd1N174grfHFCWBvS3l77tWgdtfD0EnsZVrAQlcdiPLa
2PtuKS6h5sGiimF2wO13nLgUxD9MzqWAJTjcKnjpTip9XJ/czihO/a0sRV7FBMcP
yEfRC5RHPfsIu6+360RrOaCV1Ls+RV7+jakPCOP1ufzZOyR5FJW7zGdLNBQR11XN
2S6bM/UiUm5XqQGzVfrCOoYAWMeY8idW2C3mf+uFC/6PxTj5jm6BGu671wun3GVc
ea9cYB21UOMLWZ4tmwETY/9TiKgWKOl5uSAggVGfV8wXObh1JzWntTmAZ6maMJUv
HKgbOUoXhvA43EbUjAD7qq73PLRW16h9NPowV7vBDxiJopUqQhQf4c6zuEPC5zaG
/eB16WWtcR8n0bNjejMbXhgYDd3h2PvRR4fc2vQY+i/sNsZRHZVdON7cOSmJldRQ
t8CwjgnOtR6BsI+8uTXZEk6hK8A9WvLkQCSBmU0p4Rblqm/EBSq8KhaCRLMUeRcW
+r/aIyzZ0zGZzCJvDoirX1WB5P4SrqeMNQXqgI6Gp6GYRo4T3UAu9cCGD9Jl9Z8D
Oifw3WOi2XutxeH9PqA33NU8J091t87ILdMn1DKZlQ22hCgTtvFaGjWqx1vpKe7f
bv4nWWUpuQjKg1XhpvYv0ZenBUuTuxeBM4je1nbgP6ib7n/8bc0AjPGdeC77cZE0
f3peEEmD30tqsUs/jyvIQ/JE34v2c70Z9f1wlG+/J+A0aA/kvhmoF3Wlsx6V+bXh
lM4Dib+tOOXcnTnZc0jGEXMrv0iMtFxBEdirS6sy7Kv1XrTDBZ7GzNTyxcVtnP7U
eJYpeOm6mw5LRNfbzyYMxAw+e/ZA7bsqgtPsE/X5tdc+Yk+drTuKPSRP7CR1Q9aH
Y7ddGunjR6qKAU02qvne5D2Cx+/Lpm8ZGZFZ4xCK7yV5wgZnE21DoGgA498V29wm
EeGKSiCTsz35Rz5etmkQKRciP35Lmpt+3H49NmABqyshkIyy3wmQuFoUBR32pOdX
1mavVu0tODZxiaTfpDerC/SjBjyoDisvX7+9t6yWXVQ5zsb2G43inIMWJn4cAJRU
bXz0hyH9XmqGJdqcYjzbHJ1oN2l8aNNHAFyllKZKb/oa5XwV6U2lK2dT97iCHFwT
n4lTOvx44a8iIa3MlO6r21f8kTUsonK1x1IJwsnn3vRfIcdGN7xSygm7owtO3+w6
of+N1Dmb5Ehoc7qHKKN0whtfkfzSXYn6r3wEWAmv95FW76JKt/C4y1Jno9kNpnSk
itLVBYabtOM8yL5SEG7TEEz7S8v/ghWbTxfQn+Av3kZ41dlelHW6176dNrlQCYq2
DRSx6akdhMLWW0lT6iXHMdmHDpMMAN35TnzU4/Cuq3ihqAPo1qS08TbIFeFSZ4Sl
wCwdM7B+Rn+nXgiR46k167t1bVlqUjMqmQY7a4aNfyS76EpLrMjFQZRpV5BBhETC
1Lzz4T+VzS5OVr8bJB83VNgCLCeMHgPzWk98Gk5TGi5LIfFK2uyxQB6p2bExmdHS
+OABkmUede8bxUrIL84JJH3KYyH/ApsykvecW78BIevhkgmdY8ofN59hgGsm623S
rATv3sju6u6HL4oluRBVEwCimUprdO4WvKlFw/1MPmoCl97QLIWHog36VxeSGDO+
YBBBxWJEOID6SECJ0RTxAaWRVOsmlpODpLMrTwJHmNbC4fShyY94GL12WdowYrnZ
m1HKekfjSAPtrz0whbImycxIgEfvt2K1HXqqqvDQQ/Q8fyFXFnlIMWToN3UgiZUo
p7gUjBxfkosaNenlZM4qYwHotonC1Kn/jT8Go1usf8syCbkwS9eHrsy67UqHiT2C
l8cswvWfKTdiYyorebj3tIPGxJkmTj1wgR0KTOCN6V02ZbnRXXH2l8353U6nqqWq
yAiq1wbmbvcB4fVxuwW4zuAtvlRjlyV3EOwkxlw2YMhwH++qhL62Pgdsy4hv98f2
iw07tS4qtdy6ueZdKVfwwO53ZdKwQHhKiiGLxfloHj3XGDtPUrtUOkwymrjIwjli
khNXEbYktXafy0PnMLs+nrU3T+wqAFlQLZlXv9P7bf1BAZrzshaakoFTtC7PQrZv
QOxuYaeBo7RSkdCLVJzknV0yargJW18R6Kle5yfdtDknub1xuKdeV8z8oxURxWyg
HcnBwQoexyweYL94PxMUjcIb40kS5roJj/H9lyD9FJkH5fFWHd2q6k3UyDt8TrW3
pNxuj1pmJ0+f7Y0Mh+M73pFQL5YEeu1OJZsoj+giIq0PGR6Ar+t1f3Z2k7e70LlS
yScyIWFBlre6hG0VSI8U9L3/P+9eZeqeuzsR6yxShyxGbnhBYbR48Vz/dSw4cpIN
9M0Fx1Y2HItMkJKmBHP6nm93g41FcSl9gbadleXm4S25AmXkulriudj68mRlKyZm
U5sAA2Wdz2+gu163qTi/4e0yz0H9I8oOXRzKtm1G7zgNOEg2k1bgRbiRyx7YaYfi
428M1/656M09hINHJ0IJ709c8BL8wH047c5/pupKgjS/Y/RAs9ePmsLtEabZZBz5
7vSDk4CBA3Utfkhe9kcB55Cqm8VzQ6634dNXmfvzLYnA4DylHvgdJ9nUCU9Y06+P
BBdLEe5I3RXo+GPa3SIkHmJypLspwVDITqaeOAp1XWdUx87vJsjEpy4zzBmROp/G
PAMvs5JKLk5qS/ogy6vOaCzeQD63G9Pc++1aI3GUePAPRFiELeWrAFFMERh4DrG9
0v6O/9tNWXPnsXWl1a0y9S1JNxDabQ/LwTorsL9kC/2Bb3WXT1YF0mo0JdBFxWWr
328scLXgQs8EIYeqygpkSwHcs8Sl1ikd0Ge9y4XsuKb/NChu8auInMLbVkFSRqcO
zmWCisE082vfCGYam64mFiF9eldvvKbEmElfV+mGvDvUyvVhimDxJOAZn6jXDIVs
vMLsprI6RK/3ponBag+Kz/hjGvozjfNS2+OEzDdJagYVnxBB9cDlG0+bOJ59mch6
7PC96KW0GHp+JoUA906HAsSbEJ+O/9MHm3+q82dUf1Crw6iqLanwQZ08PTny3nxp
PykTiuzgy7R7FcLEjLOQNvE2uDCIjoKcFzSOGEQclkbHJAKEBUzA85kZDi3E6ybL
qIHoamxo79nL3NFZzJgidqi5TmI4dJt3pctjNg2Swh7D8vcSj7x19CdEhKIvi92E
ilS5BPpsc+k1rBhnXRhTZdKjffSf8V6SOGS+RW8hfpM+rxOQ//KRlHCeT9xrfLwf
RwmsrccjwNRzY7ebOsuN/dzpXFgCMh0fBs+kBgI2xHke3ONBdxjBtozKPerl2/LC
Ro8keczA2BOCgGKSKNisP5cbRaS8ZOWs6CsmNBycjVMtyRWkmTXAoi1oTgqGj7X9
gTNPc1VcnmH7xSKGaqXc9tzKVq3IXe9m7y5urCVIRgM/zOYxTrNxlLFAWEjmwjIZ
GS/f80oDBERG0Qn+oha/takzaHF/rlWoX/fRBcX72+cWsTiGBCkxjRgCrWojZr4M
VeKDO0+z00BYWytKx+1WrKw8HMyVE+a+uRnyk+0WBb+Q/Ga8l2JhAbGQgAaeu2xb
S9jFrAs+xa/s0FohFk9XTpAl2RhoNT91ifsT5/GZqjtYCjCLhIb9PaR9ptNMPrgc
MQmVxfncfF037T86OyXtIoFtPxQgq5z7uo0aKC3ZItb1iH++Nf9nhzdy9eE2MCWt
RkC4ORyDg9Ry8Yz9nLablMu710bkpja9Kf8DmKqw/5/vr5hP7GJ+CJnVc2cCF03i
cAvscn3EMqa2Xo+WjJfCdWAuVgvqdEAIF8rigNqT/TVTlN3cj9kVRbg1Bnv5G0SH
ccQXQ0DyMbeA2SRCx6bS9GCzO6IEhxAOqJndVYWUenYILGiTF9+hRfga3cBR4Xr6
q7/ctIrRxE7B5cGp1xF1COocf/cIJwAu0hNFKuCWaKvkFe1OjAlrnnN0QvLbPs90
3Q0jZHvlhv++dL2Va3Oirh+xuYfuWvM/bn5ECe6t0VFKXrN8GnhDON4JIVRmAABC
6PSbXNhPJSYuRnGFJsYyvh3f+TPbMPXMvnfBzSBIUaVWLDZB8Xv48NDzgad4kxQf
0YGVBLL0L12kBH+ezt15LtUaG2mOID0BKy+o+AfPVz+hUf/7KJAJqfxCBOYDfcHI
aTsKbQBytJ4DHTfJ784+BEd7zhoBtXI8uu5VziqM+ArAaXWqrNv2Z0o49LkGxY8E
MNmGWBaoUajVJ4wqmaLvMaqfLjzSMxAzEK4iFAHqThn42IfhRhMDDUzs2nHLZx8t
O056SYCw9ABSP7W4cixj322T556rz1tRAC3CjkOQNZTPRvP08Em/XP7c5JDIwhLK
3HOcqHA/I+nd8Gm5YNVRYRWm5CQZRtknV6Ytg0I7HrgO373ifZ3x0nhaYfewK53Z
tRRpRVSb/kS/aU0yOQ3p4j2sbSgtOYsG+4KewDk5FG+99BJY2OfC5SVUXMFrSzLq
2IlHyuFi+O4zNbD+YhuT+2Zu7OqhMqhB2qsoAwwr/oUl4OYeMVefsE6sJatU2BU4
w2O9h7MB8fqO8ewsYOq0Bv9OkUyDE8NfQ8V9oARGCX17Fg+Ov/xig25/LKFo/cv7
ClhmVf0WBj786wMRycH/N95fD9vQHbQq7sUimN98Se38CK9+mI9fp8FVrs1zUxB8
4KXRJCLTaXwKpI8s4S6nfvsBJ3Wey7qYpYV8YaCXQ8Dt4rEDfSOtp7mATOfj6B42
ODmCQY2BjZsRfukfJuaIlwP2ur0WFrwdIP6hfvcnOqY2B0t0pWt6flArMbX74jX3
q6EENO2MOeNPDnbLp8nXozFuhl6dXZfW79l/7z+MDdeCEyLGpWqD+oi1QIjwbqv+
5Fy2uKY75wq7JTvC91E9Fuh1m1V33f9jTK5JSHAVxbVqP8NfcfZErc7LJLRvwvaf
PFwFG2zP1lLGPbNtcDwf1WhvuFVcna+gWf20X9t0DEgkl1Bi4o0IOCWjFMqhF+ED
pvXmCQSidAvOmp0RsYpOBowU++L4V9D/gAIMMG7yKrk5K9cNvPgUweUHl670JHWY
9/3SuLMuP8y7HQjCaw8ATqOV6c8DrUYH3cX4G8aWHsuANqylAKBLOQ+TKdyieu9u
vdVqnZtAnsBq5Mybv2IDCMcjGnD+6Q3GJrJPdrVuIijwZLM+oR6VPx8DnDmhWXcB
dAXmy3cQwklBIx8Hudt+oK8/OYzcDmgYjSMBKLEvJggBVOkKuf5vwb5k9d4LdHKf
WwuihQ3sN/n3hOAE0X6/9VKNZ/3cPQcByLoYr75hoT/5MJSig0MsxpRKPJ0iqatI
uiR9ZpS+9uKopNGeOdOaSQPZruWtFxn76P2RtiTEH7xN3/7FO56i0gSDV7VuW3M4
Frjvl5XijRWnbsklnFlRNhj/+G09yL1XcFAJmU1m64c6GH/0zT582nOPunxpC8bw
CDREFXL/qdBn3cc1H7PBxDovcbo3kqlcqGiff4q5ScX8g/JkwzwHlGau7/CXTvDO
2tuX5/vPO+iZ4ELvE/SsOZ6il0hxkCfHYaieVMTjyu7/uJ3JX08Jze7ZyL0ZFI1W
JJlkm3uHllYCUZ8PR6CVVO9+tbGis1JTj7R0bUu1iKi5utQS8dnEa29qLa4AUaG5
iJka7MzNB9SBF1YGpr3D0HeWRAfGXwQrSo46WqRhawLsLmEs32+nfXCOdLQASvsP
YbdkNOngqjILkHQQuq3xqu64vRyEdR8/GaGsu5VI6jLT4pte9RSNnczKu+a486IM
bJPgFmRuEn7+goG4CNw7yoLVSHPWznAp0llXNdjoYAyKc54BaqmuItms5ZGrnQF7
O7mDjZTAB9g1pjagX+8EvKJAmEbNqzgxrzeYTJ3SAUOGdbyV295Tb9FSglJJBTzr
zVA6eoE4/GQQUtSRr1vXGc0+NjhOsOVNi51yoqR9OQlyoslTWZxqxmr7raA/u4Cj
v0CGzCGAfZZHZnu8BTpWfN08oT/FX5w/KI0p/hziGHs5Fv9gcqYk+a/cKydpLD8O
hmoqOpmpAFb5C+hVKK6HhjjMzcPZRU6D9Ciy1Nkl51q/RWb0XqZQOhcOjWgkdh3v
RCX1qa17JziYJEWz4IfOlv+PwqyGRds6AtuSXkzFPI8OJF/qHHSyj0FSm0OC/104
cj2jn6XA7ciB1xQFn9YjNRqkW1xOOay/wpZ0WE7Xxhpd0Qhau0a+HBcXG7YOSckp
hwNegCudGxr9aTdpincM1O5sJZ0h33FkQdwY6I/AGoKsx1n2HRaUbLbi0ps29t6W
3rQ0wwRgZyDjk/bZ1QLElJSBiPOOkaJtW0S6beenYosL+ZHUFLpnjhqu0H/de+I+
wnjzhk7o/tjNgRaWi/NMA0IboT4TI2k/4VuLrRyJsddklHGnUX6O0LKXrxAu62/s
79H7u54cuLMFTQsDTX9RU3RUJg1ZHcNxiW8u4nh3nZ4SyaGRNowkdL7r64ob0wiT
QcHT3ys5//8h8wsZrOinKKCgg0im7UQAIJdMTM3NiqoQizKPtZbWmUhmU55i4TMk
c4CHcAVYVg3cYvv5/7OJObAzKchXSpuPHrfUk9oeOi+TNrPWgeiXi875Jf3uSqay
n17L54OhQowdWMXbqoCOLw1V/al5oz2800KrAF5y2Ya8fD4FoXKHHr6SDeKAT6tF
3J0nlcA3tuFdKGKzwHpeKwewYXRuV1mAO2Vh0BxjZsK4IXeWyVKQpiRPZRyDBp/2
Gft8OsdYGgGEi3w/t7YPBJsCoKxdu52vuJNqRY0U4UBBFSiBiLN+XdYTdZ3znj4d
pzctH3+1r8UNfGPvMovZFFkxARRe8tZtIBI3z0akcks3UmA4mBuTPDcW3QjI+e7A
IAnXGB/GpZCPbUy551881eVwuekdBqkMKKbKjA+LnQGA0XLKz1ZYEcQUwE2tDvCV
8OKa15AG4eOH+kxvLiFhs0cqNJzb1zykIV6KoWRAmDW71GYcyTkO/8nj6PA1dkru
8Z4hl9UMj8oBFUC0CYiDVghBP6AYxZhRGABlmAR3J8iG6OvL3S7R+RLyoAKuOyZd
Xr14bEnAjIKOEghddNVSFkH0dttuYMczI06FmktWDXHcQS/alRLca0nFzzY91OKC
N/n47CHaVXi4yiBPnHHWspUYUht75W7NnaNxhoOM8rCu5/AqaNXykr5J5H+HHvcP
8dAEwl97W2mHZ2jXd0czT4RWxPCNXlXKnh+oIaZbJJAddAJZ40Sximj3wtZ7GUCQ
twiq9iYkJT+qkvZ0z2tLWXukzduYFGA+eS2Wyf1CMpCsFDHqW1FDS/7EAXI/t97v
61y35VYImiFsY5OJtR79Db6kgZgJoZ3NoDCJZXho1mta84O+3iqQyWb0Gy1raoEd
iONxRP8VHa2paZrrpHzPr/Qrrrr1QS1KQZJkje0bl7NS7JH0+8Nr1XjO5N6PBUH1
u0I5wxlhPQ0N9MLImPYBr5SoHXIUP/kVxcfB4UFLzif57yhAcpZuGVK98BE+39qT
apX83p5DRTomubtZCVmioz4FxOAXNIYeRMewC6MGsFwnFc34LqoC5qKeiGFrQQXA
qw2Kd906hagZiRiudhgbgDden9xt9mBNYp2NN7AJ0NaAyMr1olP8YyZEjzsWgeAP
hBSOgp9wDhCT1Bqgo5KzHpg4dvGJ0wDgd5dGJt9eo1w2aOxO/muMXcMfz3Vvrg+o
QFXkqvMhCYkyYe5EZcwc5R1ohTxjhGKXLI8+6SJuOajeCwXoJxFjPw7JGjN1R9JK
b7fgjXwrcIpHEgr7/T2qjhykwb/RQKak0vd56xHCpZ4rESR5X1p82ESHBOYw+t0y
vOtiGABi1TJBZFwvHXtChwK8z6TcbVGaZu+blKhUHfOrnF1mp8m3L5mC/mWHgv2d
gIwRABv7m7UZW1EsrwIWpdCYEx175fX37bLg495n6vw2uInhx0KH/S8AsR6UJbzg
Ktg+BHN4TZUKSH08M84J0jd4EgBwnxIHwWz2PJB36GvGSPDymRNYw2ohogqxiZRH
ot47OMLWem7GQLDqwWHmpRfoGcR8xDPsTii/Hliein4T9H73AziSket304LQNpGy
UEYMESLf+WRu7JsTYyFQDs2lPe1KvLK3dqnTMF8zwQwBA3u0CNM5l+RicD9mIvJC
+ljg2QDPAizN4uamWUmufbAq0ptM22ZWuL8zQc3lmTcoCSo+YcLrLacQbW0iZbmv
UvdUI6wi2xBr+G1YbRRIxKNjg5UfQkzM1DwT4Hh5apxic6zNR16pUotpNKpwumWi
iHuj1LJXp7MERUimO3X6cyETlPXUFDGdfyAEiigIFpfKFRvW84FEH7w4ou3F9Y1p
0c6EA7BTc+HIRotWbAI3V5gUJmKMDSYgJaYo3j7vvpwABlu6mZrwLim3tBDLl723
1amFiCOrcjPs6aw/jPoY/Xpm8dndRjXH+w+ZiVJjAXRw4XbXJT4lL4uxGODXb/0S
KF50arfvEuBsyTZN30MLAekLLtMSFWdU0dzZx8ULuao1lNX5EV4hOz8gKXrvKUWh
DfdsPSAv9vSUGGtVODI62G9E/LHQMXxxRcH8ejW8uVrJEVwJXi8zN6RFzMWOAmyW
o5AsTaKyERTHsfncs/AQzLLF09ahy5kQK8bmlLw37uRq3MzViKKMoqnF/dmJ5y/t
rpzPBw7A1LhQEmClPqTzWOHNupvyYMbTVnDZMbnQT8i+pWbj5b90XEqJ336O1EVa
mnz8S6ELzF0+vlX0Q1P/DZciZKJLBAzZQEk01k1DeW3ympV4nsRPRwk+9F95NtTQ
v4tvcGVC3dfj9CdN13+GhaXvnpWJcM42NMHbdoRrsQGGElNKfer4tf+ScaMSeGSE
FfLib6r7MRSCve0MH/5n14xNMOMJCEpL947KH5R9kwTureQoZfz6xvqIcgVLwGdX
FI7ox3nhi1XAGSrsE768GaBsdoMTPhIoWXCvuXFrLjrYUSR8A8cf2AwnKXfQsCqk
Zi/Tf59b/w89ZAS96m2FwA0RypxMNXh4goMtgvqGqWCMr2buIp03kCPQBXvyTa2P
WpP1GubUY9/RsnV6B50y35mrF4UCPzdcUjk4i1qooYj7kHGIkgoB4bm6CgIme4qf
/rtviIREaFeI5Uv/uQuB3+fv2+nSzCI8H/PRE0U/RuH3GycglApA10Vlp69XW0YD
2ETEH1qzT2IFlv66lv/GXrE5/q1VDTxX4XCbIn+Fxz6FxIEg+jAlDo30QeArfVX5
8SsGr0S9QHAWlLDHaXSvRhOztzTmaZRrBmY1KL7+QsdgyHo/mggxsLG2q7w8ezub
HEKAAd16xcbSEJQHdcfIGt0CVm3nXUAcV4I2ZXVHrCj6Fc+NPd1pfcBNlCqewPwR
of8niRGxFqqIWH5onCeNYS8lVVgDrpiS0dLKGRnbbdt363md07T6gxRuvXyQZbeL
jHLKhp6KcAejqeszJY/g9pPlmlgCTFbTv25TMZV1B+V23AF4sJAIJQbGq6PE8R2o
X27YW8qjOo8vshHcLlmQDgYjiyrvFqH3l/pl35uxzGOJMBDBK1y9dIlPtKzZo6E6
7ZI65glrKMw8EwIMm7fHESslS5CdnAHA5JjWiHOPd5kXDmNCBxAKmCgZswp+601G
1N6es5/Aj2NBwaPIMS1eB7lNFpWHNX5sflI9VOBtMxV6qwc+t2xxwuxE2AhfW3n5
IU1luoWRetSapxfX94AhgITRaa5TzIspwajRBL5wPONBb5GpYFHHQ2Gy3bZAQb6D
0dxjBA4cxgoZtp4nXlGf/SSGEJp9XShhN5uAUS8yjn+qzJCA5u/XSNsK/2tiaIgG
GC27mvDoUuMgkRqTYwkJ1tiYHOHRNVxJYbNroJEb+s/PxItxWL5OwUYsc7RbN4oI
Z4Dc54IVFAEls6J3BG1XM77lkdqvMQLrMAURDvTZOB4FVMV6IsdsTfUOx5CWUQAu
0GgxPKSLof575G+lFw93jtRUWJ91TnKOtoLYedCuvGTxfjsKiXuVk2Jt1LZbCWTK
hqUYMdCHXfVKOmqyllPpcOQY3cWYYmF8iqfgoCppgofSJvbuBBMynrpIbii+Ztmo
FayTgWMZg/EuOwQPs3hSIAKtcZ4OzzncVREJgedeyMJmN3C2Teb72HS9pa43UAcD
9WMj2esTQ7cPaHf6pQocw4tS6Dr94y26uBo66lgXhRWAuC+qko1RHiiTtxdS8vaH
Db2U32MA85eP4WfC78rOufmarZuKoNC4OXKKCh9SHvr1GIbCgWAp14jJfooFg6CC
TxlSndbxnGIEzOoBlkqWxXy+EUQQyFom/9Cy7Opi3kSAvU88o+tRJdCpqoyCK7YQ
b4xh8k4s/k/IbViWopVgmExAN179z64maRFL40RUCi2BvYeSkixyBL0rA55wRTvh
hivAt3ZhegQksZPcQBDkRGpjolS/Gw23sozvY+9PWD/1K4Myw8xamjqVOu9DKm2W
4PNTwU2VC1sFes3Jb+44qJW5H5YQchJ2TDJsvHGMg8X/EOvkJ1v6E0AGf1eE7cN2
goRVQj84nT+bSz7nHLjMeQvxskjVDo+b5n9TSnplu1Vq1jZFYOWn+d5dU6qgS6rs
g6OoEoG4qOL55pm8Ygon8bPoN2DEI8E6RdN5c3qt3tx+vXRRMQHF0cmFds+PoEsP
RNKcT+jbuWjUnUMteoATQmnjMGzyPFmvcpXDK2ml3hGEFLhtb9FV0iZtzCog5Vme
XWvY2BK6jYR+fKvs65ubeN0/N/7dQkhS1fwkUUdgVscxvHMRbQqwKYUnMeT3Dk78
LVd9LHaisPuh3qbRG6PDDUJzl+p1fM68HueiK8RNPhgjmMYhlyzl8KUR3DLu51Ra
NcEgZe/rFpRVevBGBlKBruq3tiQ1lOIKoJjb2k4BkIRU2KHKgv4fhvaKLdc9PbVE
AATl3kJELnRUHO50282OEd0PMmW079KQISljbzh4x5we0q4NFtn4nIOSBeyuvKYX
rHDIjFXnSq94JDag17Qi0ltuesxb8xh0vnAfREfIQUYyq2IC7FYkbldgx/oDjN+a
f0yfKJ+0BW/wWracfekeGH7KlG39AZpyXy9p1bIHeZqUvHhR3gO3diT8Dx2W6Alv
6XCPhplf+Wrtis21MsL8Sttu42TJV+erqwyTmzJkvavpS53DherFuAgQYU3W7pbY
7nvYLUpXJh+dD69/hoMEx/HCgWzPA1N3QawOb4mc225+mQ3k8F+Pbq4hqSCQ0hWJ
NjfyhyT/aF7CZ7ZaTi1D2tDrFvUm0RZZOQwrvk5RqW7KpJ+Ww0IM5Joz2iAxMpTD
4YEmrhHRLRKUmSSZUuZuec7521uEOYQhwfLDrWmFcPvJP6GZxJuth0cCeQh02zR3
vhY/7vuhyOwJoP9VQt+PlJ+be/d64INRw0oZ6liWyyjwsFeEsmgkVTA0n7TU0Egt
L8Y3uNDwJ6ogZz+oy60lWyyvyD3NeTEiVw6Yp7eQqunQB+23fivFNpWQoQeSOrQw
Ib0DPvrl+cfdHjQoioPta4YMW6wfWQSPKsK53AAR7SVZyrWIUnU86t4I58vLWjcY
Ng6UzowZIH4exvK2rDpMuSKJ3bPcn7YDx8FrLAur5Xrme1mUZIxAE8f3vmrEFQvp
+GvPTp+NYszMOHcVW1+YnIkYWD5e4+elOeYhRlHDVNAa4pjHasL+TP6bTxCVFQhF
ekWgo7eiX50CJK08NOObFs7rlQfUYab4HUYnm+guDp0ohHZFY+Cqdf9YHP9sByWd
MI5ARFECijM2op+xCI9hXlvTj9t8ihKaIdhTc0tWsqwINIPzQGmJBLYs/bjicNED
wZxaSwE0pOYycLbgoSnkhRiTlsqtEKo9kE7s/RoZY2tZ6rXuMpy0IMHYY2lyFZx4
/PLbcrGWU4+3Mw+ZEe8YmG/sTGv/nHHVsgPQ3NpssPLdYthcPGTOlV+eAh2g/xkW
jA5KpGTGjWjZ4TUtFaO6g1ETYWBaBuLGVSDKBSsVy08426NzfAf9lpVhQKyzomYY
6jwj2fYAldSfGVrPIG6Vd2uziCV3oXX4/5BLrjTEP+X+Z3a37uoU/6Ft/a6p68kg
i+6wUUklLKVt3tun3QhQXKK+CyI+H0GYkjkjehmC1vw4iSqlkPtcmRPM/+aHZET5
ltoySgKSqvVIfSNErQwQ5oU7GOKpNCsgtyWG1u8Ok828qFCRixURX+wvuCtOEp33
FJNuWUe2+nTGeANzdwg1KPCrGpPMNEzG+j6l0s6iP6iHfP9+vuKk2wf9PErwb3PV
e0wcx03nn8YtrsyFpK8T5SHLkT74x+keK11rjcSWsJySzWuGghniZsD13B5RoSeU
c2cMfr623YR+0YdHQuyqvw2iiRI8M5SjOPCOc3gwqZ4QOoDN4pio6c3jbGkTX+gF
ba41grZUEG8pLpkmDhOCCHovmh4rORfnfNHFgA/ygFeilOcbe/gbrTwBaQdWtM1B
d+3haBLCord8TpvC0NnSRQtBtLpgJueYOm4DWxlrZNQ9YDF1abbaGaEB/K9XZnXl
Zi7ow1bq4aSGAwZn6CqR3dWYE8BGHuH1Ij/8fXtAWBmHVzjsx6m6MEQX95S61hrx
+idTnocE5UMO8VSb4Kpd4FddT/t/5HpetojOs8hz1gx7EFgrgyL2xQNqsMQRLXh7
iyD8pCVEeX9Q3gnTyANyFZI5JiVn2ptdKiAEqJ6NPOT/frqutUGfYg/6FXqL44Pb
3wauJ1cNH9TDkKTzY6G3tzkGhncmqu586Fa1qJltirhIIpiL7O9U19fOX/SLJSlV
q8Ram9F44jGiVFVtc0xGA6J/+s2+UQOQtvxI1WKa/5lIMS9mHIlEc5DZmd+KEhR6
W88ZHbTtRTEKCGMHXIhxz0dhKdc1Z0KV33vuUQ5m8JYcSSQ3U2fSe/A9IBfWSenz
zsIC50bW/4u0RxPsjwwfVArLWpeEBoPPsCgKg/Ka0Rk5HeBwchuVE9iZ8if8Rppw
90E9/yXj3fy/hVGaMOK62P7dw9JvTZVobey8JWNXjFxCJ5aP4lQOHfZ1MI2T+AYy
/w+BNBFX2msa0HjBUqarbDVmsoGOKuABiAswKV3NTT6aPWQW91zWK46aXT4/V0sP
2aNBuPQUmDSE9fPbJAkjRAAgwbyymG3TElM9wKjAQ8AQHkkcN2j0+zyQyxGlfEMD
IT4CuIOXX02I5ZmptqiTIrk4lGouVJLq8oSoa7lx74q9zGlvvEastP5nOLNb7gz/
jhG12dGssZIjMuC3MxPCzm8gk6ikhYejasPBPvMvD2YS+cZXuXHyWYeNAjmuRBVW
oyYIXIVnyQtKn3ufvHror/4/IKFHJaYdE2BokrhoH93Kf2gNwT2M+blYFdnNyOra
DxetE1af6JaSx2L21eKOolEqab56JVisgzpp4Wgigtd7fOCkN1cN1t8ifOmlUog7
K8vrahKQHKMdyZwcCOdCLDb/yt4BrTPKp+wJm0fkKjPJLwpPfK8RmNqjwsC9Ln+7
jh/aLJyN+/dp/9zxQcnnQI7oPVKtPVOlzIXyDCA0oZYD5F7OpJW6dkKP2b4jvIUS
h66Oi35pfiWTuR/3/PQLRbLN4wQPavMF7w/hcrKn/8CitI4vUgjgYW/3kRlRXvzE
mbp/lO3kIslvz8QCPCed0MSqjKuGFIQnokbRZrFebWIOuk+gh4LDJW3X6c3oERG5
oyo6BYTy1feWFQS5vcvjY6TTcrpMEeTdAuAtrqj9uUvu89laikpQb4BoTBp6KHpK
fhwyhaooLU48Bfw1jFesuI78ObNnrMRpjRzZLDNe6gdik03lYgHJ/BBksaWumim4
Z0hy9EoIGe1GR8g35ywwtGrJgOYdem7o85LcxanASjjAkqSD41QK+TNQeY9KZKRK
TFA9x6K4wUY4EslE9RUcZG5l+bJPWySvxutdmwEERO74Jd94VbJ+5Sni+R231IO+
6L9eWDma8I2W/lUwV4PUJB6TCw7FHQQ+QsYVmY4Y+TNlM6Lk2QHjcDsb05ZNqRM2
rffTGQAmcfnx6HUHmUTfheloTQ9Nm+UyKAtvljn4e6XUJDuPaTtaZaB4Ntsn7Cwb
xaM7mTg3HqzZUB/EjQybqYh4VyGM6lVYl8vq/MQEmyZOWkfAqmNAwniZEZccbLpy
NJJMPyifeD7fa8sTB8b0A5lqH0j/dS29adf+OAh7l7z21PNfodpnrA32UsOdw6H/
9RDbtHlT5t/2pUfgEBHAxBfXn1yzYB1frZ1e6Fv5HbAJiqtup02fqA/V/azjVqfW
OaWnt/40oFS86l35oJCtTgPE9eccak8Lv/ZLBU0YodeP+ypBMmQIFLk92AeNI/3d
AJjmtJ/6Ly4cnEWLyuwZon4aVG0GyHLXNhkbkHohXEFvcNbTJOBxQaAmp3ncINf8
+Bf3hcdQiL8D9Xm0FzXkTmXU/h6n+UNIfUtbUPdttqw34k/G7a8UfV/PxvF6zOvW
nalGA5suOCoUsGDFG8LVQbb39sYdJ9K6JTDDlBwX72UwTahYunBM7fBo2D12KoxM
RN+drodc2UqfjQI4rU7L8447Q0C+lHPqES8tY+7tdoVbGNho16ldoiX8EFJMEJyc
aFj0Wv8neQs8QLQ6xdq1oV9YmpqtcnFXuzi9fX/wobVOuAbsK+jIYUUB3hFUxHLI
HEGOyqNoeDOAHhRuujb3tN3mU7YK1ZTq8BKxuIe+JWcJfbSlzb53xRlnnbOA1cbZ
JZCyqdYx7JlyCG9Xd21fGTh4jeZakPMEmd2ZVa+OZFApHhyy25B91s/qP/tEnI/k
m4K052Q7XvUw6OkFRpJEheC1olmjFS2ai7PA+zt2d+XcypzB7Ln7gU0RuyVclALA
hXgA2E2W+QGNWhefbBfR7BPtKZQvfwTP1kG8JVL03L/UAM++Hf2IYu9j0bkh3PO4
7s9PbhHLWRo7ngc6znu95C7uC6VCvxIYiFIXc59PpCZMwee7i1vWAiZtSNP2DYon
94fdBOtt3Ha2+LauXwxJMJ+HnDuWs+AM6oGKNsT7AW0LmkNZ6pDrNB0JVuFK7D98
iUgXwcqnYwsZFspIjbIjMGXs0Y3RQ2EQwFupo8QtfutFVUgf5J4xfyqTFjJdyxLw
A/sdQGOQPnR5cCK/Jb5ESYY5vX8nbd81QYgk/LmKrmcREFnR3ISRFMUVWwktFVYp
VvheCyXiRegU2cYLXjiPaaqFVR72PGoI5lqRWw8sbXPNKjGrvaOwC5TIXrz1fCix
G8g4BokUmP9rydhM96rbZboS9iiouO8Vgx+IPVjYFIPH9tlsA92Zz8xytoPI6HxX
GPsxFA3c+7HBA7Ni4MzOUB1p57VmlgRLzt2NyAnktWRaugrNX9cT8w30e4iXc9l7
H24FB3h2w40obMMxktexViM1qCyaa2XDJgQ6NkxBR8g0snTVuQwv/em7/82xjD1Q
VQq/PiEB2MZFTBDWGYcQ37m7AxOvMtplo4oBH0psv3PscfEQDpS6tzijMFvXAHFk
4Tco1yyRQ/P7aou0Wnk2kO2HcM+lBi0XKB8+lFPYFivJQ+Hkba/aRCkynfSwzflA
1krkzljtsu9MIPVTl/g2F5V7b3FQzvHI7ijYodcrhgF7eKm0O3wmM4bXDyhUjR8J
mdamDkVJn74axGC9/DYniRCZOpm0Fbm0vuwLjsALkj2PoTI3DVDdySMqMUjGDMht
YqI07vSWjwdBgPq897idmx6W2wpjZpOqlzBq1Bj5QH0KzojAWt45m6W5bZEi+qFQ
3EuKukeMNDB6tM47Zi9m1BMxJkG5d9YKC2rLiKlSGQWNWK9/QvuDN0DgXTEraTpl
Lx94byHlgik5xgQ12INkDImviddM7lkUSRlROSPRAVD9z3ZioanvL4W2la22CEL1
AKjxMRkMkS7p9sswYUaPkTqkFOsbr1csO5rPOQSeBH8PVmTGheF85WR0k2GGWzd6
9Lwnd50XqJEmtKzuECaRJAmwmBwfWskkIkB7Gnc+gPgY5OIF4qBok99GFbKIaBxu
vrtnyjqiESna6+yJHYEhDnb63C1LZyZPeb58mR8eHPIMY5VfwgxhVGsZq3ne+5ql
qE6LKyttx8vavRWYyIzmTbcNwzN1O/A8oNlLx4mebvgU55HhAiA3Ar8lRrqRZq2y
GNnDVfKg7kVK8/fgapt5xN2SR/spOD9Mue8D77SxxOYnTvVdRzk8ItRJ6UQyvxfi
v/4RDTKB2Y7VzrWHFhz/aC6SQyUJATUa5m6NzD38j24vUcSQ5G2uLoveXaABrRY1
Xb6hrBF8jbbDI2+909CG7RGWq4ncqlsQgrGVyd/4m1Xn4SAWd0U/Q/av2g94ZWVy
2+bu4rCgCBZV6538FXjv2qfvXjnBAaT+P3Qn4Niy/UyvXZj4sYnU5FVKNeJLR6BP
C+wLtNUKGMewJNmMExI1MOjuaX3SqWtq3f3zmj+t36LeZTphzZScKFwKa/tKDLPP
G4UznzkLwt29//KiyK6eB2GMovIdx6By9hWGB7uw0RraMvXve22dNkiVtObiX1Jf
/XwYNcGxLQXLiMAmxoVuybvy6IYLPp31VQ6QPuxBNvrfoQQN+/3+mtQ6rNDgqrbu
zZJwlHH0Mp43Aoi3oB5MF7JutQece2DdOndsonsmimjTPLerRQQyTSCHhzi/lL5R
daqr0nO2wG4rR6edsAV9K5fGiu/rTpVsIJGGZlw0TChMIboqtPFwYR8v2Nj6vnoM
sLsSlkN18Yn164kfXNK9Io1avjQf3DyeQ7jAXr76IvbyktqbU0LH/wyeXLxWBgFv
qj66ZGsMMY9H6EeHcQf93uAiGCcaminpPOOf1sHn32Ir/DJIVGmYH78+k7HWHhgf
RjCd6UuyLHNLW0VQ76N0rURvSRYQIA+Hdt1Ts+r+jLDUH79kCixDPpjb7AGeDDvZ
LlkN62hQQGO9EEx4kOl9taiav1ZRFunNuOPxaPvebXNHPwVemwFodhKmpI9pvvSk
AL5VAK3eLPgN0F4YGZlWKZxQeGjTByoIT+hlzj3DzUpNwFTjSids7d92b0rCoyPi
gf+PLjH4QKofnsVC+nCoe35bWhT/823KzH1zSQ8IcEaUmFzE+KBcf0nkheI/Ms7v
+sjGyx74qB24wSmLM+4LK45aEnce57WsSc021GWCfkSfXv5ZxFRGDttK3lq2pXjV
e5NEONLk2rYN/l5KpLV6k4gZBvNDXrhBITyN0hrZDRQjDmCcmqXta4vvEz3Ps2VE
r/IZGySUW/UZY5dz9VBiqE39NRsjWF5x9AoI2zGyzJVoysGFCYysP5+EHGC6Ovlz
WSkoF1yQlsqpgAgIfLLoIGZvABVCEva4jw6CChgc9HDyVQS9VotgePM92A3oksnL
Fg49OoonIyj46ji1wuXirgOdgWqT65AfGDVY6UZmIxfosw7TfrlrzbI8XttXZeW0
4ZdcQGSeyr9VqVNuNw7YYl0vOzoOtep17psZdEbwxMqBkCQ2WYIxw5RhfqCfwugq
Yz/qsL8+fS1GQV7v3FNuofAqdU97hzkH7TstwT8Vs4Gbl73j7R6jy6NxZSxbMTlD
X25KK/OrMH5w4BSm05x8g6qKtxWkETQZwOWiDkE94jF4Vhtu6CRmAj4VEAAXFip7
lLHmu5bYhOR8ZtCHB7gDetr0EvuoKJ3y38IP9YQmmH4zY0G+m6GTNOFEfPk43zMX
6rCSbiw2b3FPcAiYLJec1hxtNzHs+7WLbZGPobIE6AJ47Vi6yF3yAiYusBLXXE5l
yhtOSQZrAMlrnPBIC5XG4vVaxvD+WRyKRNLhq6Bt47RiF4zHr8makDuz/VsqG6wO
OK+44ddBdlZyflnLo/QUZ+CdYi5YRU3syvV5meabxfHROfJ1oqaNNGAJSQHg6BQk
BxCVH30KnmUh0pFW1FyN9grGF547xatzPk+sp7sSvOcRJW6JE+SRLeKlVB6OcRMF
oIgXkZjPDNHZXVq0UDSaq2le5A/3iv4nx+nnCilDYmyek0GY/u5I0eq0+2r8qf6Y
rNkDfHSJX5lenL+bGzVbwLRA8DISClyRAeR8DO+WakEvA5uG8PIS1USq2nM9DrdI
0o0nQ6m6H0w3YkGYSTw9AAzpR987diE5/vYJwqVMhsm/tHc6gL31UCya+mQpm3rH
fQ1D8KYQh8Vf3Lb4qhTEYgvgfyjAzH9bZ0jdidAM4g5CWLwhI7v0lPK7fazi156j
rgpJyVzFT+PQbG9vyQKnzrfxekuCDWNXEzqlj1jsfViyxa1XoBqkff6+HVdAIKZD
UXbVK8/Bqg5FFIJUfBTqgtPg47aGEJlwX2PYreFFl57Uw9O24PzvgRqhl7XIhJN0
wr7CcyDYurWyXe9d1NmWGkFRn7UChox1wRob9GrQEVK7XQxVG7qJL+T+Lx1xC9zW
bRkvApRmz0As7+cO8BybCYfX2pkqfqFQa/4LDr+RcBDW6cxWILFxQYoS9pWpo6SU
Jh0ntnf8IqRFw0+4w8kl/knN7vDXRKL7OEyveEp6SmCxolA45l1jilobEGINjkk1
2XKeHHCHVO331+0mlDHE6tNjD/Yt6tdWM3jGP12yZTfAwvebbSVBXTVMLB06FrRH
L82QF3Gv798W3MNRFJL+0a2V24mFFM7FgOf2SSo24GCH3UJDQCa802MLlV3V4oOJ
lB3YfPcUq0rMKAHvJMsVU38YCxyi7wIBqhesbE377QfWfWBfHn+71OP+tM+LKnDx
qYeTo7QkDorb4MdyhimLlTJ71Diagra1iOpRdS20B92Qthx8fiWn02xUXmziD4sa
crMBtJT9Hx6+Rz60OfKpSNy2NwrHg56oUnOtn3XjWo9UWV2JE6IGZDiU737aUGNr
YKnXMtyy54fZG4ACbUiR/fx+ZjN1UdPxCN3xRXH2xFpY8MfiyMif+lf0VIv5m6cQ
qdy6L/GwF9gGlLvFg4PhC0z3oMCprZOpLdiZyjPBchZmw7fNz/t3YgQBTbFm7o0o
hZEQLympcd5vS2vz4wD7B1hj8DxnOIa0v6ZNb7VCVaXxVSHyj1AE4l1VsDmIWcrJ
wRaI9XZjN+Lb3593qPAEL1yFHpBMtoSMEEsZQzI4AjlhIvSfPCYoJl8Qqxp2kt+5
ULhleleIhEwoCwNl1/ryIozcwWU02CAQHSQmiylp/MJxMCAI30pt+hnhYiBUWKpj
9p9ZoL0xdffLdtdPsSZOiD1sx6P/Yf0W+VhRK5X8/YC6m3JgMcf/aI0N4qtPNrNH
YWnaUxlIjCcpB12fNh9RucFtFSXtshe/DEwZZW0s6S5fOdqIB2BZUeVXHSRVaTbp
GXVuVx84dCMafMT8DWlbhMwl45r0A6hzSeId/8JiHYejLhX6NMNq3/gsK6GWSJO9
YKU34+O3EOBN9qqe9PJE88+xFlQq9+S9bDk1h1FAjArUg9bjbdu1TrUU51rClfVM
oA9jp9l+tCVq3wenuylmrQ/MMnTDTFfOaz/s+cvOryspio/qzk+z55qUTFlmQKDU
ZXD+aV+fC6gIoooYHESk8q05DZJjlj1J7nRWcIYkSCuTOCfn7c7bFXUyyF9fgt4p
qGAOC4WGTdb4lUzWbZc+V8vVhgmfJGJR9sYAPlcdXi78usPZSXsxJ2TQDFnmRKUR
Ub/8msCFDpGBh0lxtPC4/XclSTzNDKQqcPOq9tNjk7i5K1tWIraiCfZOMwDdtkqR
wl49GpHEZkjbGAod6uxVnP5hGGmwDWJXx8wY4s4vW7AFpIEP9LSCvk1DX9XC5pBF
fxckLxHVrsszadOEnusFJiLpPkCnURshZQiT38OjpbLELTbS7jbQheGYfzATWMt3
lNrKiVUEDXXowvUdqCQL38HheG3gijBfndib3QedZ6UmE5hsQ9vLGLdZL6mYvJlB
lSyheMUN3GB1hdhDEyicoo6QRtyUpUqateCU2OLMYjhWH3IiQIg92KYjmlupoxQs
lLDfEivi/m2uktrb10AFLmZtYeMg3TU71kXkvjFgmtze0v+xAHzj4iUx/hbWFZkN
mIRiBZqu0Ap8Nv0QegnoTJ0c42hSyTVeg3aColOWruzqGEu6Rv+a8fYm38aZzyvb
a3UIomW7G2NZSnbGCRwpWr8qMk6+Y4jb8OFI1sbvdfZkBXjupH5wluU3Hqs7CUtm
wsUamK/oejr76AAzOz7Q+nwCJwVerawv/uqpWfb8RiZH8JqH18xIaKQar4/JbDD/
13QnE4e8y+aqGUFg4YQk6fC2bKrRorosJEwSfsGmcvptW6Ytq5hTob2WElE08m5i
/uyvqJZu9AyAb5MtNA6m8cCB3h3sA+xieCsl7Clk+iQlltMZziiTGI6ER6viNWfa
FcXycMct7HtcIrWPOVNEAXX0XZujk53DuGMttIHLC/5nvjt4xH1undbv6efCM739
BBfRncI/FGSu8brqJ7USqMeCGqiapcCG/n4rSGb70Gp4VOm+zJ/iZOdLHP/ZX8+c
HfDCy3oCAE97MG5G7OIu5UanJ1bjfUeG8WcSnYvvAdtAjatpCbmf78u4FQYYeinR
A2yo37g9esWhJKrzXM88T5ql1fhmXXTyw3ZfG8LzH2ffX/E3il0xEySmdoHpzNCd
sq13Ev8X2ourbhhl+85ryV47GFwPvwcefuHbbwz8hKvAKBojce/Pf9v41Ixu/xeT
kXJWY0+c74dHJHbATeTFKVDwCnFBO7SJFCKcSh3xI8J3T9+8I9s360pz+kTAQqwC
aCtKrInKMCOwEo9+xjFZTFXfwzx/TgHpv1+N4XMIudxrCShTqvKGOSzMGG39R2Hp
wkw0ZsoOucDYoW7oN/JzPRAcqUt98yJopKsIYvd2ANXdP++/eDHwXCLZ9+di4aHL
d7NpYOzqgLqwLjPz407fxrUIouPcJ7X5t74gg43z1bcgVBs6GU8cO14LRxaMdod9
NYUznDgax1j0VQiog9F9iU4oh7RJNjN8XTVrCcEw2+1NlmcnUlGO7axz63goMXLG
nCxTohq/zb2Mw8XheWJ5RKaC0Y8xz0hNsj+tlw3A7F5xQ5dbc18UXTnGb6uoXlMW
scg+Mky1DcVh//63nZYYXHjOi6g4lAulYY77apNzluWSV9wWhp9HD6zUIn5/1Vwf
7YjOE4Jm2qBVzGdHJrCGcNoJPJ/vR3dIKeKGk5qBHkGGw1UEkuPyWGN/VP7jDHCi
bV1p3n4jAmDJemcS6YDQzKrI54RznuiNmY2H49vC5OJU3Ra9ZwKfQ0mfTiGqd65H
9mONlmhNEVlMfhmf5FYWUfCXMY4U9tbQdMvDhETGRc1JJphhMNhwPc76ylFjzR/L
DVD9f42jeq3WbNs++BkbPNoR2wmr50g0nRr1twuSyL+bteOBD6rIpCnWWWDCPkUW
dKdDiy9SlrNBtsY2SiY50OjfTcRWnXX1Upi2SlBW1gaOw9AfLlWlX6vCKQsUFnxA
v5KvhPr2bEYBa/OXFZ7yCQRaABI8NuZJ3lTC/buzUgBn36egZBqq72WmnO9N9w7s
QQkCfs0Zfnu3ysYqAGYcCW5LmSBhui7I+cxJuA1igwHmzw7CLo/6jdgctKB2YwS8
gm6bAhYKziqfp3Di0KHZfIMnIeHx1m3nhv4k1I0jgZ7lpiLusr9fF5EC7At96Pdp
D1GkuA0B7km7u/PGtx44xYTEcfXwFI+SP2aXhdVJahtbJh7RHT+gmM5+D6LydGB2
0hAmKgyI34EVBr+yhSyye7Scdvfw4byuKQVqlgFHgE1+3mrTE+RHHCaY9cEzaPlM
EobrOo762bgW0pBNy/qZhnD/IdEio0Bu5IyVy3f1DduCgW122SJS3Pm5lzPfV3fX
s0ss9rfRMEwtzhw8CApD6clBej5m6EZRVfUkMXAl65HvzHx8U8ZKw6xkwyE3yzBb
GSJVOnYa9g7lb/dENHi/fk5xYzhf9oGOOoz5MZnRiDFYj6C9gZX+ikX0ZzX/REPz
oqfct+Bv1AkCi6wv8ppsM66lY/HMJL2dhYbJbgDaB4Rfi2/RC6YvtxTMPLMgcTic
kVVlHibbvs6Ml99qipG+1iVvIp44yUXQDqiRhJGsulXSHxQVs5YLUi/usMH8IlTh
KdhPCFf4XWF4XcJOKqf+Nz1sB1wGCDfZcPLywMEtzM7IJUX8YcG2X/PWN2K6Ef7a
bIPsHSyPgxollVMRseeRy/0qDb+dcaXak43z9nxU2vrnJvSnk7uJCZvAAsHfCNCr
aHetM0x+GTUIhbmgT430WiPwcLkcO8DKyChWCeYAc0OUGXp+mUQKvTgsulTbj9X/
9DALZrnr6Twn92V3dWT59upORRrveom9aEHuNo7Tq8pnZGthWcwDHCzq+peLHVCa
a85RTdsN0utS/Lh+CUOi8GGLzsafSwvNBA+geYoWeNrQ4j73tTHiZTvKcjOX+vJ1
OZO8bEMkr5RaVzeTFuHTi0jLku4sZLXF8uoXn7Q/zh3ZDEOfQXC//jlpVPC/Ejb1
eM7GOW2xCP/b9cRGRYjAAPyYJy6r42NhUuVOf/LGa8NjlD4/avTMpxoauzVSZjfT
rS2YOBgoBg+EYs7u56HzZEx/hvqmySDvf8j0iHBBliQNfHHElhV+E7Xkic9BDbzE
hKKgA/8XySiLnmOOCuh8bMXQTDdfRZ9GE/7V23N6ixsn2GTz+NzigjnT3L04Dx3o
pBiqMQ++isHgpw53/7gnDLuyZn4CkPJSd+3iouTgegoQS9IoF1fTp0kE9RPAWzYs
yRVKr8joDzcV9GZqB6g7pKXjWqtblHS+V+JetQ+L3TG89urgJLnZqPhbxunyNZBw
nRaKdkE1yQExZp0niEQ8+cgNT1XXRAO0I1PbwZNf8L5b6E+GNNEfxD6BzvXKQCXE
AbPbKfMdp7SueOwQ1xMEvaJuVrxmYH2dz72ITmqAzTRvr2bPKtcPBQQR3GUgVBIq
dEiP6t348WFk9khMxoqgrDRSoX9zYldaycC4YIQQZRDZ/xAqjjS9qQa+EBm7qoz6
WDGfkaIt1Dv0wl4vcITAIhjNj3nSBnl+ml/jZHmqlchDTJpVR4YpcfvzDCqJt6GS
s+KEaWs+kDWUQFIrSaSWPNdFvez0+w+nx8md9giKavQsJy5zxpQ10/I2huitKPZ2
YVMdGtvtIii6ByJxQ1qzf8OBbMm8NcpqbJAXoP7UA3EIiOwaHqWtJEs0fxKpDXSJ
qOsr2PTTJ6vgg44ZgTh8ubvQcnddGZSV/7h4npCQqs2SpmvWtx0f5W+AlZuaNRWr
Jq8Lts17s7bk+XUMOs6dTgpsmiqo+WZYLLWEtgfOEfr8JYRpDnPmHfseinw4jL1W
2UK4gY7CM1GBlq0WpHBq/J8xlGGvtuBB/mf9c9ryyH58t1QCYcGeW8h8vHwtH41j
CKhmyfPPByONMeaksfHvFLEMwwJ2glzKf37ue+YDW5Rsa9K+cXzKE7WF5JLgW09W
AIbJnXyzLQ5yeVZaYrnLhthKN07Wl4jDoIb8LpqoV78Mj1dgIYdJFcezw6NFLW0N
GlHyHuLw+v1Xp5dp6xpfz11IuXmjl5P7kzZIvr0TthCx3kXK0vzv4cOm0xnOxkDH
xSn+b41pBjwvakJf5y7/N3Chd6pSgLWRNkzfCEoAXw2GaMPMTdjvpApNLEi3eNrG
mgNcKPw5QaEoHFypoNdnlhqzuQAfQ6NxdMsuVXP88kQcNWtEnmuum3/DHDcFSHBE
AysG3CLZaaIovS80M6rxxlXOAdKdnbZAvxmxfCWHLXn8FklnqlgZelptlBpMt2sT
a6XIIsreOE8mwvThXrdXMlY7qOviGpq9YeLxtYQljdwVr++b3o/jIKEPUQDySyk5
eT95mP2MzLnWAJVD7aRVWLGcQX1XLMH9cLUMJn9bAxR7VUUnBGbJ+JCQfgr288cS
2u8X89zl8oyEJ6eS3iqSgU/MZW4YgXBQsFaRqskCPwskyOat3YwPZ8J9zjz09bZo
WZlbszogT7Sfz1TMyd857VUyqQs2lx4zipYegxVWlNqXYKtGO1IolrXvfxon1mI5
NNaWdFFkTGU98Xvy0wOGhLKgz3oPxaB0m6hCoN14AR/8OpT+Ccl2o2/p+j+pNIsF
Z0+3vUkGX4YBa9xOHRaffNnzzwIC8ZzhfbTZdOQ6TbMZA6aAHVV3Uqv7fisu34Qk
/YldxTCFKADGEWJt65IqytX3afjMs+gWhtYDT8p1mVtnaROXithQYuZXoNx4VMiV
h7vFOgLKVVUaw+CCVDd/HHtQnsGrqWDUW/cs86SHNBP2JO86svl6zXQERrvSD03t
2J56+TWisLEkgGFyeaikvp3+hhAqDlk3yRqHiCnTXgj7w6epr4uQSlD79/os6ZpG
MQ8/22UKMf15TOeeojTBHsBJ8fpiEGY0jt1rc9NwusV4y9GWSoeeyYwhNNAf52u2
1J2TCDOHvCCWH9zT1Ezm/6lt2AmwverjS4RVOs2T0AykVOR/rql70+KyFfEiictE
RwlFw2f1XhDXzMPJ9xVm3fk02YEt5zzTvNOvnDPYUceuR0U1HccuO9NOSSIOygye
hmxe5soJL2RCc+x0VnTQ5mi/BshedycVmjy00XTOtGQgtWchYeVa+pKBzbrnBQtP
P3RVe6ot9cZa1dYfzUdDD6lN9ojsN61/8sNDPrPiaW3LPhP1bivGX9V6qCrGQhYS
PRk43M1mUO/hHxMXiLVYMFNHGjBP/Cou/9Y5QHOHoGYNJl+FPFPCz9VxXebpbtDJ
9BLBS+JRpxZLc1dbf6glV1Gk0v0KRGPVpYY/IL8WQgwybYVYsrx8We8pi5BJ54fD
rfofhNPyaW6q2xiXZ7Q1wh9fLcM0rklPvmw6roYXZAhvAdfG9d5qtq8iY/zwNKrL
px4nZXJ9HUlV/JLfBG5qnqi620uhPPZvDvhlSDHoDZPZ8Usc9KQ2h2pdTh5fAQzw
Eaij2Va7hZVoBWMYdfgUNp9J7KJ+wxbFgO6gnTHOTiSV7QT7dkwbp5Y2mcEZjXnb
ZNiyQpvddNkjzIuPQ28Go7vlnO9SEo2827Dit+onTof9ay5paVAUPBxloUd6S17r
vCmZrCwTD+vPiJoyKPref+ZAAmTbOsBIobdynk6vFCF2uE0C8XzS2qdl3ZCPVPti
c/NJfg2cAkJXRLhtXfe7/mi9A/C40M+uqgd1fUaE9U8AjPcCndyyQQW5g7jPpWPZ
nr6ZyWEH1gcCc1wUBpGZW4w/jHYMS2nyX5Ow6QAxpNe+BlWbVq+fw1l3/DasPI3Y
hFACfR2Nh5PTUdi8jfP5LRfW8Kdfle5GxuHCpGGSeO15sODsmXgHsA8C6K6TZ2FI
e1d/pTiHBPxafIzQOJSAEfqr7zYBNEzjiFwKtOwD+TJ/WfeTbF/c70GDCpHsS7z9
5P342yPRulCzxLLK/teVVEU1eJ5ps61zQFFFYAKToeFsQU3yxGESDMba0PavajWc
LBwgLazDdNyxBTxm1tGLWFJPmkaWfWgE5dAzga7/bRZ0rOzjrwlqfEiOs1fnjk8Q
LCD/8QTdOx7+f+/D0ykOqlXzLEYtGbE8vZFrnoFyuTYtee4aF/0TozI/AkSQWkVI
NMaUFk6HlJTqus6w0Z1qJcETPvSAXYacSVEwBbHDA2QQYRZe0azJxXstdQ3Buz7N
L38/PhhSP8JMSahLBj91fz/k4ZKGW0ylt5WTdtZ+WayZAeS2L/m0odWmZbKbDTKC
Z8CMxvFV5v0ZiQ/mqiNMYMRkeT9QzoYe4xJhw9gwiA3nrWRVway7tm6xdwaHJCNe
N/OkdXT1qMJo+m6RoZuWAepaQ8Mab5UzKxELatATDofzRXa3HylYYvn7HQCzxItQ
dUmer0zsC9bOSEOYcAT8slVVxKcxFoH9KQmmz7JfhNiy42jqEOakrC8UtmWGBLc4
3jqLLSGDNANKOjfhbuZ2l0LztzVd3oRW6Rpqxi4Hd2aQoPuj1q52b/27RAtLln6P
YNFV25L0e0x7FiETnsVXmD+ZlH+iQ730qvuIHWEaRxvAl2yoYtS/QoZ5WbHxTGjU
2QGtUR+/wx6U6O5J6Bpj6Hbc4xLRzrt+GLuqdrc7VinOh5TDN0ppXrRXjg7uxrwj
3j72KeYYroSMUqaGpWRqeIsOEY/yPBbrxdiS0Y2heLoq36DSykhdQheFsIEPQMHy
mV+/SlRNgAfGudyg3gTYkm4EXdPrl03hIVBDenWlLiw8QKgqkNNhLdM7+f0p8Bw8
+kN5O+D3uN6nnM2Se2gWIq3CMmmQlvIJJFTcFk3HSUBtRC6b1wr5mGQwGymw/Ahk
hhvvulDslh/ZB5yQwbrUVc/XyBvDsh8+lnezVQJJ8CvfqooLsZls+Hs8yRdUEOCH
VZwFY9Lj4IBXpTFmu4Ie18MyB+t8G2ibFVjLHCN4SOIUMSZE0jO+zZ8S9MWkRVyC
KTBnT9nBGUI1FBza3X7KLaLaU+vMiL6xLK00q8+lFIK5QLNzfYzopO+JvrErHQDP
ouTrsqd3p5vJx92oz4dsdPFunv8pPzvNUjwPcXKPOzRU3LOUNGnK6iuQgu4PQkBV
YpW7aBsduwK6lFHCDmuXZfQ6OIilnySYvqH4I442mWP8+7vJjCjK/MgKEkocjx7i
ZrQqu8WTkuhOKcdgm5E/Di8m3kRYDC9hJEd9RudQl+LH6I48+5I76dJpFScb2kLr
5gSDEDR+gD9Fx61DNXyjPRq3OIhdwPfu+GlaV0qQHVFXC2GHkympELYFNfNqWk1/
aGu8YXW5M2Rd6TNLuuUaAhY9jnvdYzuwQ9c7BvJb83YyEs+u8muxnBzdGGiSKr5O
/LdBkafVOb1Bu/hTeyTzz+VTARu6kGpycGGxNXyXgrPW9jF+8n9R3GfLmeDg7L4B
sLm7S8W9pBBQXvFe4JGYJUkIcmEmguWnjiOerto3mZgknIrmnufdgLw1HNLGO/CB
GCsGaBlvF0aXV1+IVcZXhKaHPQTVdpwhBWTKA/LWw5LFFNRPGT+M1tiyfhXvfUII
TBEL1aj8YrfxQioa5B98hmGHaBh2wlT+osBPX4lhZ02Kh1N0dX7Y5pq1M+Zm2NGl
JuBf7fJ4MQShPAiA8KX9Q6nalL3LWqgn0z9Fisatdf7v40IMOBCs1yiFI+JfnNmy
1CIzWC6mSpfxhtS5AmSajTXUojisMabs+LQWexUmkjeCqvehclqag8fLJioGEOrq
j/2UDRuOoFoBoMBSSIbQM/7Zk96UDLDd/wXHGzE85tw3cAHMBVDXFXQRg4zFUWxc
SxfDjaBPtFiMv3lc5bN5XJjm8HdhHP5Jp8a8iAOqT2qL3iIOP04LLewb239ZjME4
ZwJAZvZhBObZXwy3zEFase6GUf/fsEvgw12zuF4o6sFRqeep/Zxt9Hy9UCq9l6EJ
/Ccvz6oUBl6UvLTJAsK1ismNvPww6NV9ZYkHAQrsDIHzt2urkNqNgyy4cRHXv4S8
Q+8BM7fEzNwmWRwC7Qg79hvijGdrAeyha+X6szMqjJJTeoZ9Hcz8lLGcO33zal4+
3Htlhc2QJg8U6fAEWjw/tl5hXg0S48sm3x5UuW3/0U6kkSBdbTVEvY46N2juP0nR
uYWvPpWDma76E+n1Z0MYRyCgPe9BcejdnuES2w36GVxoOHeVoY5mAAFIwHfLOghr
3kUmiiiXZJF+aCf+sQpqA3MqEs2aINBjNjvauqmj7YoKrmcbOCLPBi2CRoudiEku
NQMxDbLSriYd5/LrL4dZ5akephpRQ2gSQ6cPZoYHRAyTaTxKuf+An0FSo7YlytyE
BYwin5fK+hmAIXHlRXyEgzZx2zOxptDi6rY5sKF83OLckrJ30a0xj9L3cGZgu6hY
2NMVKh78yhiqtyht8z6rtDlFrJRG7mzVxDTcExQKYPTM1hK+KJ6kS3w6XNT0fSfK
btkhU8Llq2mKXAFHURw9qakMuH7MqAt63vRTn0Oc14i/1EHYbEUEHZP4LB5rJWIB
XwYiZ6DLVvVxsShdcH0wZeIh/3XaBStLK7Jlzq2CATO9iGkVCjt/FLIQ8wr54JXB
dEYxcmAGODgLTZAJrIVPz3yv97F4xUwjub67jfTJhSXVEQkq4X20v6fDO8Upuyar
POx9ds/u6wQL3IvF/dA236vxIKnyxfHwbBjcmkit9aTS2x69pABFusGHH2y1D8WL
c+3iWqXOitlQreewTPriPmjN/zI08rJmN4pTDXFZTRLiZ0urEwez1bl8Y19jDwfi
3hntPRmH20VmwvqwKEJqyUEHeVigNUPFauIZF0HfgcbjLRII5ZJrFsmt9194giDu
yn4pNPKZ2ybT5nvX5MpV43gjff6cyL14qD0XKe+eEaM7bY+6jEb7Hw1q6qkVoKJi
U5KvNY1Kl4GO67Ic0ttBWkfYh+TsXwNh4O2Vxwt0MtSDq4qAl8riBSj2RmgPjdRF
4MEIcdASaugRdQcfRXoQuCV3pWlvbwcmwSosOVn8vVgaOLMSaprAB2rtWT8qz0Zm
GnZ+5H3sewcXmUnojdIDxIKbesFPthvOmxX5+dfiZTKtZki4v1637GP9E4Tl/bcE
1H1zyV7DWSmpANPGI/yGkVGiLmhm/T1cA7VTzU/hPQ09oGYLBb4ku3fb+o8i2QpA
CtoeOiIenAIo47NTRQ/EfP0/JljwOgEm3mp83E5Rz1G0/bOluwTEA1tV8xKiTw1P
Wa4V2/xkcbk0YYVOC1YvXOIxIU96fxe9qk43IvFUWiXvvWbu11PuMbW3hl+pAxbq
bWpJ45SqriJCOarNbGazXGGwcWQncdwHqGCpbwRk9vIr0PDaVnVTsSi7TbXe5jxH
tUuWt8RA4qGe/hKHBdz1ceGnx6vbB37QcA550DS5BG/ejOLfJVQg3+k7HkzzmnDK
+v/+fJefGbJN0QLJFqDhvg6yKHJdSNvahqKQXXTvXTo2xyCmuxMhT8125FkiMLR8
lOS6K7dGWo89AqPUij78nItNK0JdNewhH2NfTEDaMMq7gojNg/oG7xCHO44vcQ80
+Xe+Ua+6D3GtsQP1xAcw1BNslNmCJICkrD2Al510U9y/djogy64du3G7llRjaiKL
dr8vg5H+tU/11xu+xkYG6kVKQYHiLL/PeKDLKqaSvKt8B7tIYXMOL8I+8ylntXbn
N1f5n3LcYkKLDpMSOzIkTeJetCIdKXg1IJEQ9j/JkmkEG+VceHf/+v9USemW5Iwq
5a07eOL9hUgnzJVtOINxyHmUVgEeuGvmzz7wCEvylBxBq+L1zPg7zluRESsET0Ni
udEEUeH/bohrEsjd1L7X/bbXoJbNa/pS+LY8+X5KyLk0LDld2t38XeTz2Aw7X4GK
dLa3v2mfiotiHhDjZtYlUutkDdos0LQLx0Hos5Mh+yotgfGCsRB46Qwp61zJSNr+
mejcU2ig0XovzVz145OnTRdG5A6/WiR5VgpY+skDtkw/vfA+ddQbKT2atMmi2uDw
LWwf4tJJQreYQoimpVe9BLigsmJOWhzaciVLTNI7FSgEufwADXIaUIEd/DTOim8i
HZQGYF3Ia2oaU5GGGsHXKM1QVMMNs/ogma76L/bNTVGPuHnRHeO8ONYhOZmNcaAE
Cr8lm51iFgCdDPhP36mHiB24ED6t8SfNlS7OhNeHEYRudfwFZstkfT7vefZTHgkJ
o0vItJ5qLdfvZRebz+CcCl++zjQrjmtcexSm5lZhxy9vVKIpSEf0xWPXWLt4foYR
2mgMS4S5LgT/newBe6JJyp7FNKOrHT0FjEHfWgMLQgUO1l3/d3Bjuwzyw203zYPu
MzW3RWYu4oQtprrKbfkJehKLA4JJ+ZmD05QoQbSX/sxuNaepV3/9Bk/c28DO9fHa
/UiklMdHrpFuZoqoxppBJNhNakLVUDVb03Lgr+eAExyDNNQYF9AMVRcuTQugShmW
FLxCXTVf31HPxQEw4JAKBsSK2S4zAu/2BQYSbcMSP+b5c7mQcd7Nbf/lEwr6qa6k
YxcLxWfzoA0A/abVjR/fYdyZvg7laYTj1jZXv7+Aw71VFF4cdfnLfr4JLOfqJlif
V9fvZwn30anju2TTAzlmmCkUNvkDmed1VuCD0jQxNyL0dz6/QJ6dz/tjbMeHTcpC
P76sShzhStDKd0rm9VomtBenNcBp2a+6NHNaZ9XIDeujLUDIgeNSaRPye12DqZKG
i7H1G9eVWr3lpnoXd8iE0pVyIRBKinOy0dNo8QUfWHT6KpydQRvehXB7471El1FS
eMPJoNJPrTOwgskvF1ylldwYGiEtpQCaiSlxaSNLYNuVTzAG99K5bBtSyVaH9Rn3
XHS/nepsSo4CB9kKJi+l1cz4bKivdZcNxwheKF3MuZXxWJhAorcvyGdGJscjLgmr
j4l0yIZLe7YqMLU07A9Nt6OgKr+l/UO4UxcpNQqSdBLWvbEiRUZ0rTu8Q98N3ki8
CMIhNxpgGTSHFuANoSmjWkD9kSwNHloxcHj+MgK9933IJp7PtFcoqGPla5zCmGRH
uR9dMQzqOBEn/yS8AP6hWvBb2UahqFLmwK1RkETkhZdV1gOEo9Ak0JXC8Ax9y1rY
NgcJ42qyz3+GsKuLmb1esEh0RE3CPkSc4gosMTPXzKmDV1cPtsWChb8Ibh/S06t5
81lTuY8r8Zh1JsyLhFuknhq1IEu2I11OWpYhJgXGlbyHcuS0DE7QfdWRbu3xUd/b
H1UeRtOmNK7+x2+EO3MIXEEZVe/sTMl0Rrx1VBefP65/ZDb9cXrnM1LC2adK8wK3
IBM6DoeUXKTcErvGeVE77IAzBYlWvGNZSMgb7V4MNVh849b3qatH9UOXvopjiebA
tFQI4owdWoY6cWetfV3DLquUKWZNB9VqTn5Wl5nozi12KGMvLgMtLou9vldruhsr
4lQzSVbE73HRoGdgCVM6EtJAlHzTp3S6BkNNdrn7MfsdW6vwwFLUeeNJnyPtVtCx
YPgMsEkRJOUdbBVSpkiNW0n80a7hOrRBnypUvJ/SZw7L8nUa2ZzZgVxthGFecngs
ddDf3h1c7/Vk1e+sikuDCEWubipLePSgu1wEap3UVWaS4uvP+D5xNCpMLWfjPGF8
cnMNqaXNzWusze1IRTPuUrMcW7MMFvV8gABmypgcPQ7/n++dpQDYOTslsmdgvkdr
Zv75Og/SRP5ItRXlSQPX5TLeXM4Ue7vxwwsDSfPQdOfMfRg4PtxSv9+V9ZKxuC1K
qRaaRgIZOas1cstyTc2UKub7GlhihoA8200rEL5Liu6z3Q+bW0AbfJVXcTuqXUSN
0E+ZegWQkzoVhcc1eaLocRPschFhFFI9bTE11T/DlSFW+hZwu1pyC4vD1xF3sBF5
mTmoQhe3le3QiwlJQsWkMprU9lkC3FhODKUwLARX+qYzB2XgsUxbiE5U1OUrJBUg
3ispMWzYA3ontXLfUyUib1VQsXQed2MaDKIRdcpI8CybG1wNMGSY7pGA6+KP6k+Y
gAjz3b2IyJkYwLKC/qPed8oaDBYhvS25tMYWj0j7LRva+FZLpRDBeWKzYIvkNPnY
VQZFL4VSXqVKBssNgCCrcO9I7RFW87XAJeSbqYUX/LqepeUs+oAJmz5he8Us1SjY
kIDbVcYQ5Thx/PaohbeR7yxmfQ1mWzOAB4tbjTb9zu2Q/SUJAekVdLcxi5npQDxF
WYArRSVAPEYv9XKC65qeIyl9rkWTNP4V/Uv2M6WF45ZdkKmoh5JK1q3LIjBoNy3f
6FHYfEcxkFVe3Ec7g+plDOU8Tcgqh5BakQrJleor7t5F5MtDwrR2aM/Wz10z32h3
/Ci7KJ+qekn0Y/ZtcPMRIgNbKmlPeapUdlUC10aKHWLHRQaCqlqP4Mm0+c8Sm8YE
JJNaQDXDgoGgAJuF3yYr7CjOkWOHB+Cyl6AorV5bdFP8In/042R0Jsj0GwWe5rxy
Gb32N+VIMKr4cUE31xHfOftkUYtlX4BR4t0GX39eTff7DEHZrECSlYhjPYVdDAmQ
bIVBF/XaYYzHexkttU/nhrGDSjztgLN17MzQ3SanW9jtT6WET0tvRtaW8k1VNih/
OzbjWBqNXsmSlp+cIjyxfU500c0rdnZlaJyrtCyeVRPmMKzKCy8s+USgbcNFL0JE
qtHGRhgU32tTdIrCjn+PgJy0qHGMxu/OHyLBs+dB+iupQK2T7pLbjGRfR+DUptFf
A4SfG74LZ7TyvZNbD7VFY2ReXd034vobns/C5DKU8xpLq4UucFoGmNTkomEiQBf5
WRqMY9xHGQYzXV9Q/Aww1EJWMVAX6Q1ukoSyiBsyscGhyLtC1v61seYN+c+3pd4M
n/EZmEbbC6Fna08K6gulriS77RLfcxyS8w6OOYlRnXXwxlz2+ngh2Z9UZ/lKvAoR
jut48xFAHXE1NUtw6ziATp1vgHPqrHvmPo+KxUXykAqIth6Vb2ezDbYaq2/vlIVd
IF5efw7bDgBYGbz5CvMcPYiGF2fOBnCdK2Z9A8cmi5ilPdfjVRHyz9Iszleb0X2A
1pxtg5BfDfjHgndTME7Jb1gseFIhbzPZNE07i5277pSUMy6Y5m94iJ49oQX8KEzv
fXTu6FpRMfuZnmU9Nsyi+afuE5rWAGrKeqGRh3bPiIROsLjWltLOv/2AgUpKLtTU
mF/vrZtNPrAK6oxmcsgU5CVSDKHqkLUrUxxtfHKaq3X9EAcVPveEfI5pMT1sKKpW
Lt5mNT+rxdf7Ls8QoG/9PJ3vyuBQNUPhxAdNuLt6VoTq/TwCnnfVZP7DARu1zwfh
eDX34FnrAAoRgs/Gklt+IbUfpvZDHsFoTCrT2/QH4RfD4K55hU0vTqHZ18OIbLyw
DDykQJKBKGICXdHn1hajVgU+zfl4CIq5XOR/b/GpyxHEwu2fUJt+ukCEzSghbt2o
Y5k+NkeY393GHT5zINFgPHiJOSdupLV0tpi/hCLtNcJMcDIHbSZ7UJXfnnwWMJod
ndH5+IDtZP0B2OKJ7fWjflRnwdQF8yZ1/FhLNoyOdvpjHtEfBycx7OCZ6nO6DZBm
aPc8Oh2VpeO5oFW3l57/mNj4i8sy+gqetandRVH2cjVgdr0/NftXOEFoHHi2mq9m
+rjgVAeht91EEKtnuUxvlhgdLZ5h9K8cgluKFlgE7ZX+KUg+sAWv9scnZwCjl5kV
OTfDtikHD+siWKhlORjUZ829429aa7ZgWPY03cDVcz8rNzuctVG72yq0SKUA4RmA
m764mhwnbeNSUxscwN666aZ+avBQsPsw7mUTHND8iXqlqzIJ8rWpSUsRW19k1A0r
OmjNDn+NPm2Uc3sDc/Bw9dN8Y3XfkZfGNdwX+PndBBbXipMlyVTUebiL7pqG4OfS
dfXtn03bPF0XZ7EDvpGMJEr5Nu5GdgCm5jmPR8rAghsPfzF+q/3IMt/+UzbKcva9
VyL6WfB+AhjuUoHOUgiXuoqniBM8q2bC6/xIAHCKELI2XCAQAiIK3eOMC3c29qDS
C0Be7uLhK2uOyiNKNZOoJu5C7jVtA2AwhMX0VP9t/MV1pMPeF3Z12H73Z+/ZUXNb
LGeWVcKtiJwooRcJonHozR6/w90oIZjwAL/8XeLnk7EyYZyROsaktNPKB0QRJodV
aUDvhtMVrVNO+SV/oMPahTgDgMTb1hlxZUzZ4KPA8xMj6wIwW631ywqFn1be1xir
pV5yRAP5UEzQpaQS09GEGMTIRagB/SJmwbYHggvzOhdo7oA4v2J4Wdy2IQc7z3Nz
VuyIdykDAwwNOD/HpC50WlwpWdLyzB3S1PYGm4u15lhG8zp1R+5INfPxlE24WlEY
qWwbT2ZcZATdta23mXfnCMrGBoa8r0Z5BI3s8FpR6xBrmpY7lwBhGWv2anS3DNW7
/igxnhy+xYauftIsi9UwYnFPAv6urJM5esZREsAL3KvRk98bDW9oS5GhYUqQWs+e
aUlF7s66dApjMBux6jt1zBmCBp1mNoiVo9DN/ensTbcLB5oceJAmEsyUD4lr3BlC
8bnDBPqZQbleWckd4HK+TWkK9aGZdIO6YZyuRhyK4D+3CesmFgIhrQRVGv+uLAQE
fmIukhGK/T66357CfYEeODT/6GfUuwB9XfqAYCr0fcGovLOzUciN/dEK0/Y9/tIc
brAr4PPLoJb0S8VP6jbOnIRXjGj/yh5MBk7eAZBMf0gblMMusDXf03xbdotv9FI1
Le/DveNKFpzSedERxesEo3XxenoCqECC5qbSvKVS6mlhGfJDx6Gcj3ToEQZgs4XF
w55cywnUjliVWcfCt2NsqAuHAa+sjq+iaGSSSbaYcmAy0RjW13O6sgBpjHfjHO0S
iAqo7zqS8/YX+kI/jNykEphomP6AKQsRZsLbDfEd7yBMqF3XwohzYQ7cjoRjrsel
t8wV70ql4LXoDpzW3rSZSNx11lRbXOalPT9CZWDC8nOltqdbZJV0z9KzsAXO76eZ
DojWuzg76Wl294OxVOTQ31gQEuXvHHBmIr4GsOg+p4WIbOJDn3Ir84TbPTK1578H
Vk+O6oyeRjRRw1AkYoTQ21FVG6ocYVTv8SZvwY3y5a1tTDehWJpa5FIv8P/UIlS2
AWL+kvEcB35VU8ggksyVrvwnCnL0L8IkLUJnPQAbIcXXbl9yU3ZblFIszcKWhPup
pHA3K2G6OtuwAYTj3sbYIEItU1tuMcHXQ5TPT61Rrdy3qpx500urEu1ttPeaeGDL
TLn++vBKkq//lM5wlgtWTJWdYHUiLTPc8S5KEXbpAlxIJxNtEDfDJ42KJxVwA0Ma
O9j5mPy/rM3dUAq15DZVbM0i634H2lg2AMeScqKnfcYXlMKOaSxPwFwbq1D8SrE2
v/+HGRftubdjDm3LCHS1d7O4+XoEx75Khjl+nNiOG5BeikdPSGR9TheLKrRkVI3i
hAvH0++J2CaHVVPz+NK7zjGuF7YXEAnS/Tod3KecYxwXDOyr/5pg2DdqPXIaEyWo
mQVHpkVJ9Rs2nKVt8zJ7A0UqIaQOfN5sUXEr4SdvFrzrWEHqU5RrFI/8aJ06aagM
XDpx9yeV4Nseo69P3svPwFQyg0Xj8w0SRZIgzcCl3lPqWSqtMRpBGMmLJa02nAtV
WqJErB9thfxnxYvSmBwHU8ggHzxhOTGGyqpa8tgWnNIekDeRYXWGPgwNZiyMFZpi
eXW1V3R/HJg9YNZDE/abkWWrJO6nrwvOyj5Oo980B54Ztu+M+Bp2To3qjaPR/nu8
Jfkuy8iN+qtD1SVF1j3Cq0zs6KiaIDO9xhXnhDHqf2CjF62SDmTxktTtt0RGqcxf
pcDi8L4cejRdMbG/6sYZLbwZutpnm1QSiRl/GdAX5H8xklmquHTPXXBHaMPgZVIk
hHB2q/7pPiS3uOuv2tXoPur9dWufyCTuhGq19WajjW3PfS7D6Ki5UstL9h7MCZ04
960+1RQ7S6UJGSlVWv7KOFyT+pPlSPINMs4EQ9vRd/Ju7RFqYkNcUilmU74AqrEi
eJUIo6FrJtP0oSV/nnw+hPavM5o1lLwBApnipAUW0RwQxzVXgmxO/gS4ocHP+0aJ
xqyrd/tCP9ZXwo/46+pqLp1Tclyld0Tt8nav+6VLY6XmlyPjhnwffXC6htWT7nPP
GbQY230wJPr/iCDt4g9VF5BuSKHT+Nk6VpD9y9yy57Wwsk5ttOf/11v5ZmrG5D4w
hZ0Ixm1rQ3gjpupC+IaFlH9EGFpfitIPQbYjfIj3v2eZAzxS111KYR+mHQLgYlME
GIVrZrUrBjLuEOs4xybHjHXd7C5GhGrS9EBDdCtVpCmKthwnsQX8lWlTPW0xNdxT
0Qi53HSqfSGSV4v/3jBbqS94IUEgHh4ejM1rud8nyxPhBaS+0gQYLmTjDLCeDIMc
+AFxOuI8UbqE9Odth4mWsF2rJXiErvXTWk1+RsPXz7IRDWR3yfkrHoBeu9bA0xmd
XJHdK1MZL7i3FxA86OpwFEkixpwH4k1jVCmvh31aEQrGLpiupwehD4ofejkqksa5
mSRB81LxLwtpe/rGo3D15wDMsaQYD1CdRcgvEGz7TgGs+T9bBroM9h580h7Z+5ES
HP+S4LM2U3HPLtL3/3thDPJV2UB0bVVcVm1XgM1H6EDJA8lVNDwrFE0GAkBfRlRg
lY4LrvuCnvDN06lhRQhj3mDcRKx82SpWrcU07nn3pEdghnrJkSMK+im2KEHH91eW
3iK5JaTSWrzwn/O/j3KUludhXXjcSn6Z0MH7ea/TJCp0zySCs7UBpz9qxlBlRpGY
j0ef8i74NhdcyUQ7mnImog2xzjEzgaryQ9GAQC3kSiCLQmdErEuWOBWTsHs89cZ6
VgMdN3mKYABIz36Yv/5lZ8xYyCsA4W95PMAkTs4aFpvEuRy5Umpl518FVem1O3OE
et8OzFjXi1Tdj2J4YRHlyRHQ1BSRNhZG682rWAG1Zod20LS6+Z+lzmA9K8l+bJd9
uH9eg7A8namf8zqyV1heVcDJZJO6g0X3nfyRD+Rf1eedrDrUEFToPiusWvxuxI8O
DzDi5xKduW7KP+9/yXBz68sjeiIJgHt3uL+fxphZyUmnBrukMeeF3hrFzZg/PJPM
qFhZ5fK0iuYIG39gl4GEg0wZNK49L9SQYUE0QY5VHolsFy+RShpqaExpLqsNCm8C
i7Pk1FXZ3J2jfSsY417DHEacBzno4M8fTgHKQeejN/sLcRvUrSmKU4baITzz3s5L
3TrPbvN+1l4xAzR5SQs5vgfF39D37/BTzvBdwZVH06qEq/gzlpaydthooh7BMdZq
ifr+35Pl8Dtqzfo1kvy5Kjl+bugwzCqeMqQ7m+2rumV6lbukwbdODjmkB5ob2asI
WUyF3KWUBqPpjGp3jn3jsRfPlFcyCepL/7ouO3npH15OzY/cGUwZSa/rZn3m80/i
xVA6wF2gMevtJ4cBENeRaOodDPvr8id1Nytgoc2/4R1KKGy4Up8bo51hzz0HEcLz
SRiPZzrzxjV67iaaADp5ecCO3kdCnNPO2IRQZuhh/hLxNjqo3Z87kZPTRjwKqws/
rQ3rVLL4jcMW/OZV6/dPc1cX7DgTw75Ctlkaa7gaTlD2Tg9AtqeJWduIdTRnBjlz
kdo8X+bgtZkQU4Po2s7MVz2/lT6hTuGwNG2BG1yKPQ5TLl/sbVsH3XPBWlCThY/y
Mi1qvBqULlTUTUKbVbHKUA6YPqdxXl/fuiOcJeagkfi7of1KpYG9jmeGmZ1DHn2o
YIr+8bJhhvncfHURT+6dHcA+Xlqj7KaS+fKrAh9Q2ApIakymT9q2OhQt0QHIwHrh
1sGSpfjMOs/T+9POYgKYb24ZAD9RHhN9jx8vEM3mgt5qaKPq+E6icS60hEQMltZK
b4cNCPab9sKbiyg61wBXn0zLXQOiT+MGeEwRenXuEIWgNWQt8Xtqnd74oL9ajs/J
AdTbe6Ves2EqbkmKJTfuicV+SGKpaGAx/q5FU/6xOefNVCFxxjjA9oFa/I6A3ryV
o30jOYob4H5mRfgX7XoRQjTn0S0nDTNgK8YT2S8Vz1XL5noyl1ZYPLia/19ek+Kf
6OCx2s8mJEHqvLAO2jjifbr4syjSCJP56Y87NnL6fCqyAVRL7drnayGenkOSlUi8
2JzoYQKq2bHrZpZbRmZ4zsEtP0o7mVSODLthFQ+ORJ6mMQBz+0loki64oTLD9E3V
QmtGQojmQ3pbTMeXYntdoFIjvqpDdhS0lqzfK1xyfdVE2xSz5/lori6ROR4RM+vo
WrB+JeUQ+fBj8qZ/7cvfGpLExYrSCWQQy5T8rL33W93Z1qXMi0C55jE3T3ypFQu6
SjaGgzFevEdSE/Q/tzmaLWRINhpePcLq/qV8GmQ1kxqqAL0GPS86uP7RUArUZ2+X
dZCMHP5iBC2pZoNJIhRNCk7LwuO9WJC14JmtMrFXwSP1T+cq6J2kbWB/4lUgVlTQ
inEv+6ViOVFWM6qNtOhKVWLG291SGjhIBAwI9O3p9neTgvxOiXSIAPvif1YmRocm
H0Zy4z4f4BXCWyxU+ec/znOyrcZcWO5EigTSAKPON2pCIB6qmAuBBcvK+yo/XDT4
ceQAymoMmVvwYh+hduN308/ZMvTYVrvkwi8LATxqg/d69/8ErzjvaqX3bWcjuzWQ
Bl1JE4vKukQl+EySApVDowHLoAK/q7FG6E9YiF2TFYa24L205/hPYmLRXq5nvvWc
81cjAFeaS3Mt3Q6JZoCGNXjICMNxSRUy8ejQvQ7mmc3psMzuJK7U0mrlT17LGCjR
/aAivYJOXoom2XzWl7NMubVwR4xflbEGMJJU0tbCNF71MM1ltQiY/Tymx1s+d/cB
0YpYVtulnT5QJNg4ScpzaBPOvDbVhn4YUZDpwFkrBakMhn9RpSJVzd32SkTETZsT
SWj64SgnVcVganCr4AAFtuqoUT2kfSnmUcDUpx55uOvmrC1IiQYxOiZtJG36ov7H
IlZbPqxRYqHQvdCithBBIJD/GzkYMxITVaEBtV4FTum3CysAoPqMzHFluTStjkBP
uoLxoJDyuv2fbZep0iafaQ07B+KFmKUazA+t4EgaAt716pVjHFFkbWHguqkzxDtJ
BwySooixdqoxqAstvX+j4mjkrwm5fbmfUVNNymD09j8KbxUs7PU98ApJmOQnlAUU
qoBBh/kaG6BGIIWDkd8S1mK9cyatQI7RAirzeBO3Kf2IC0Q0+xMQ+Nk7lZ3yI1T5
wZBAP4K5ecU390tNn0UI4hXQ1LpUDmMqs90UdBmn0UbfHnU8WOUPm6LX96FRUifi
hsOzGneQU8yOcU48jFVhpZGHcPanH/hKDZTumnuVcFNUfsvppafZhxAvvtprrgZh
op0GhvP8s9/YeNDhllE680nlr1sQQ6PF4Zu2iz2BZf8ucfne3MyOzHwlxLoj7raZ
jYHgPZFdR4Pn6xKSZaYQIoS1qxm7oRcDN5uqAZBvA61kISKiYsQkolhUxg1PYc7F
rw+Sp/yVdsbRKve7x/xShucF7pXv3PZiukmqFHf78aFdfG+hBrLMT1bZkcXRuul1
2EweUmu87IGrlaq5LIp3MRc5AxSGz8pqz/JJuB7R+tV/iyTS01uW9nrO0+NShwdu
kQZyAd9RoAoIHDbCNXEc5UV7Wv9kHbh1kv6gBflvUk/7Wla7PY5S3xDDxsoXISLm
sh3xZ0mzadXe41zudZ7wjlOiy3pln6XfCPZzAJZaWX8kejt+eGEUcIUwuCLigIsZ
z3HCjNLyDfrMahKUFCBPtPiFILcYm4T8dcTh174tUyvXjqOPEfDLeySl/jmB6Dhu
mSWojRQAS9TM9yVitHXKvElaclSOFvxSVXa2vfFmz89XwPz6WmDw45P+6rdaN9Ua
4yylzwkTZAIbCUktalZo51kxfutftlzSmnWszh34k5bHeJOPMawVsA7YCZDnfuJb
192CzOAndhbEdquyu8LDB+jZzYrKUMCF1pnttgo6z4jluA/UfAuaZVXuz7fWuEgX
j3YmpdYS7Ft8QTKDUouHASaXU8oXY22Dqe0IcXxdoBKhf8A1yacjjUdDKBnfyK51
Yb7Q7sruEYayoEviYWQ9gDuiItyUyYG+d4P0PAiK0MEbWNx87sTP9YYP6RY3Wesf
So9reLALogcn+KQnhSS3YiWywvM9xfx3ObBsKCelX7q4L+mKCta12bYo2RQid651
osbqQCSVP64LBM8doCYlhLiNwQqpCoZ4o0EDNFVSfbd1pMFSgdYogSwhBet7aJ8F
Jz7pnHUd+C1iz+UJXVvEH4Vk9gC2MPtRCSIJ2zdJDVnUfiR8I6NCk1REeRTZrCsf
90vfDFPEfU2it8NLKgcHq0FhV/1AFZPPsNkIE8gu9+vjzFU9Mj/NJicFGg215USw
ncJBKkJq+IXDaCcZhKWUOCFwcyqfTdXzdWn6372GTDIFLz+CG4qW9FXfWmKO+GF6
E9MbzlJ4nBMCzxeYfSAXZ2ki851iO2OXEbbVjdhkT3xGKD2LX41HMdkvg4JEnxk7
szxT4YAyuoFhzoRUq1R1R0jZGHw4dzNjLDRIvwTTG0X2z/HWmFC/DYfov97xAOtf
CvM5XajfeS1xIUV17k34FLqmeeZnKnj9j4/Z0iWGBdgqp5oncmefAXJLc8u/h7S3
IgOi9QnITk1LA1lg7XA51Lv1Y46XvdotmjlZMziOQ1e4shPyDvBYP2NUlSAIXrMY
pIVqmysJrW+QllQrqs9wTEQz6uxs8hQIgnFCGyKENZE8SioszZe0i5o/d66mWqG+
KLGYhNnQhQP1Tdm3r847VBC6Fe3AgQW+Hj1wPL3tUPUAZXz0bTNZ7MYQynWDKHoz
xo95N/9KCs+ae5c9jr0m9yN6I/jhlRg8mkB0BzqOHr7gbyjVV3ly8tyTD+equYvn
u30iyEJI6alEa57KLPgzj9rilSQjR2d9UIsYcVeNNVKDL5jo603M0hxsDM+k9zXj
FlY4oWyA8Jg2GZGRczBOts1cADBI2qwu2GjzfMozzHn7IrYLRlmDcPt50rKc/lAr
2PW3G5sMzgk4jzcdBy9HWaqkc6m6X2jp9pUXhBaFtglvK+p8iwkmFq96kESx4MaN
crhww5fWR4cxfcGD+ZCE+pkXIm6gS6mya97ImB6G2JYGV2URbM3tit5YQKG/j88e
m5S3wb/Wa6e4PYK0KKfpP7+WwNWFFmY1CDXpFpKtTDp++118fQ+4cs5cYSEKryBi
CYZhGOQRyrLg/K+PPpnBxFZmstiQRfcU+MQ2aSc98h8sHUKRSSeDn7Sb2BD369Lf
hs2S49fIpJtPb2TR/3VvdrBclEijzmtAWPl5udFKPyW1qVFjPqVe/FBegHM0F2aQ
+5e48vU6EFqNYqNDItlSavrxSyLxmpGxWh/0lKcwKCLJgc5OOHDEBZsTwnblV6lh
fBFWeT3SskPYUrnByl9IbfScNlm/bbeTJjbwt6lmxXdhiCJo6uS0ek4BPgWx2Zvd
O10//ISPRkYukOCx1Gy9ZZrK7XbRlqnpN1q3ErRvELTOxyX6PFEN3NlRJBx2m49E
VJutTWHNtZ9SOmWlc1lj/LAyzNnqbQR5U3/qyKD5FspOTp/UwPnACKJTSuGs1I+r
9X4ozrgkMPcwNeskubNTjw3lNVRX2M6EDwPOoed+MAtvAwigCLK+E46YUwMNe6Lb
9kT6xsW3efHNceCVMhn6F4tfAazkljVZdsgF9pSC9KyH9iSDb96qQv2FIIkqi/zT
i49z1CJTu/6vurC11KSBGMWiiZRkvr6fngRFZZiwkHgFzf0HLYRTjFXjPbo+nVq2
BQ1SLg+rxWLZ5uP81fgZPfFk1s5HrwQEy/3K/WkCoZlMfIN6kZ+bbibBePkbxStH
ifPyew/oHcWeJ9R4id2yd+pK7mv9yi4EeFgpYEn5mChGLclvZ8nuO45xpDuL+fo6
WPvifJ9a8v/kDrFwwiCw1ePqBOfYjlAbeE5OZMUTvmjK9yy3W9ULd/V6w08ip/PV
u+gbd6825ztRhN2Uo0L2BeKHKln1UFeCysXT3ovgwzBrdsOwoijqtXkflgp8reFH
yAdCapGC9xqHF/umJA/Jf35GABJi+hP/7Q6Pb9USF1grY/f3kyTZGIA6PVdMMZUq
376WSgwLcUH77MKMQUEvgrL0QFtM69EqmjSiX8DJr4uQ7pIvWbgeIax4CH44Ektu
WBh7p7/k1FKsQq1oo73RAFpidId8FZ/fWPKCWcg70IPNlXjW8frw5oL5SpjMlAUo
SMBPY/l/K5N7knh9j5vztNIfJ8IMVUszVBPLMtpmpbFFQQ432MQ3ScteXqcf4uYC
oU18YfBIzuXPAe9GdmXa2VTx7GerA/bT2RXZnE327kpXBk5HgWU0aaPITyrz2J3i
vlTzSIj9t6mjbcK2C04IoVxi0DZUB3Ls8hamgjRDTO1y9FdNtWiqqZd7DlXEWjTv
tgWPCGiKS1nWDa+6EnsMXA3yJZEw2BirIHUw3rLInoNb/lIbfOcPpHH8czYBKw33
eZT653gRbasfbeLjmbV5ziujueqnPsZJ+VkVTWkGG15nmTzTBtaaycAA/LgDHc6t
jlbN3K8AyizA24vq3qW/2WLGNI76QFzz5Hzdr8oId9PrD+sqzamR94E8G4jQuIMv
O81qQligor1a3kH6vhAG+T9+ROskHFwT2iTIRZO5xOA7SYJRAK+8eLKdIC+Ctzz0
bECD9NYK4MSt8mnISOoDNiQU+wu2IK4M45ruAbFpUmDFjvUqQXbas0xBmn4Z6M9v
H9/HquCD6g6j0tDfi6iie7eNVGLG/e4T7i82wxNnJO8eOTxE6XYfZvnNNfUvDjFG
A1NxrkBI7H9UAFgHCqYR8J3SIxqc3/Cc7XrdWKof0o2erXDm/qYtZKubK1AgiATo
+oK7o4UdQB+gNPNBkUZBX9TXqGM5baoGwRI5ymu6EQy7LkgrfLE4yKyWZR4bIlt5
Pk3fzHtk38JxCCw9/bVwjqptChnhdr1pHSYoiJ/czXtvEjX2BAULBdTk1YP9C+Kp
kULo8c3eVsH2tZUhM9sdj6RQ9z7TllQFF1oqXVou6XXVfOzfCw1+mzRVSx2AwjiP
R2RDQAykx/ZrreH8d1twDdWrDLc7WqFTBgpn2CVC/+VxF1K5gZTT6nv9zXaK38LM
NfWfkMHbFMU29eDNu2B8Uc6gY3MXIG5Y0OdQMgRwxUcqWmk7CpvEsarihIcu/lPw
puOdJ5ZvzR3MRoFc7QBRQSjePxeJHft3Yy7OhPfMn3ZaMUZwJSF4SGIMy3Qw/GSK
gKh2jbnoXGrdqB2zXAK6OSVIOlQo7Tkj8oOwbe5hDYm2hSnRwmAoZADjGFhh1R0i
h/wwIbVYbNUwrfQ7lex8GBzflOB1361YJcdX0z7BAkVAwt6eyN9tyAMYo2gGh4um
9MNWkat+y8anpgqf5o3VoTxDGeeH7gsqe+JpPKSlb7gThBJKwTeLMFyzOzecNejY
WHt6hLof31iuZB7cU7VMfj3DrYnBWsJ/DqzsJVG9hVCI+LQQU4CZ3/LJb/kRJihM
nRKnscCti8QHbRxY6dXo+KSI6vBqKe6W1q/t5CT6Z/dXtb51tkzV10NlZCzk1evo
yyt82iYVR1LV4E35846cF8DW3GVP2ksNb/PX62DwmHQLgBfR9ucNppnqq/m7IaX4
waY2TsvMKSEgOrr6AVznxzrCZtUQ9a+yil3NyHoF6Ah64wJ7tHbLUIKz4RxlSeO8
zLuJR+V1H3nIy3QV1lpfTA8I05f37SnUf9ZFlhOklHb0mveRvsQqmDtFBtRcg2jk
CP0hqLA4CNzgueUE9VvQwdLfjY/b9DULs08EbExemtKL+4je2MjDytlIXg0q3yuW
uBFe3XwqznMfts87V1rpPt5/YMzxpg1gBIYBXqrHX/O1iQyO8UkV6lW3iWoOOicK
0ORJeIodxymFdvCZ5Q+4Ll7a3ovSFXdEsEPdfemoepVl96WSfKbjgCWCXeiNz+hl
lJoJxkNLiZ+ch9cEk9o0BJnFyq9TrAIfnyC5WIxX3ZEqFbENMJmA7FkgobTXbmv/
8fwlMqPwbthXjeCQxoAzPqx5ZIBoazrPymvCI2HH74PAPdrP97KzFxmTjLf7TKEX
qvMQq/jxtSVdy2j1SQBCQeBe1o4z0pBihk/Nm5er7LcYfEBU1C17iMBOONtbJl5r
p+1CcdFVVW3BZChXnLTqQvl6fth+GM794dMWiZotmnUWGPQblcIJgnVnZxsH5yny
/d6WG2CJw/qJvqR2q/+l9jknbEUrDob8jlHtjxbsQ4Dg0zSbaz+TUT4hmAd+vmYj
K+k3CbqAHJVoDJYnpRQ5mPRpAuHN7YuUedn9OKlke5a8IAtLT/pEDJ07BphNJj/Y
9iyb30l1L9AtcVi++sst3VDrcBL4gXa1LGejCYFK8CyFEDmw7VjZUbZm9Xo1GbFS
ddeoEFUWHIpJGUgoqMifixpGYA9jguqrj5/3AS9BPjobuEH0m/uoOMdncUN9G4Iu
96AOMFcm5T87oMazcZEXZpNigqMT/U2cJLU7J6YVUyjUApNQxkEaOt+pvdU6FvjR
heCOjPzwHA+zNjY1jXg0w8Fxq9CHIsj1/rR2ZpghDNPCjbIBny1OGt4XQwH6PbTG
oxD3Fh/No4VoajHRd8Ullnj7SYs3KI4w0SSaU5gjhsIDRqBQbKg1F58if5lr1Orb
Udp2nSdf2OJgYv7fCt3Dzzv90SJrTXjdoS8EAf+my8jV0rOCMZ/EqrIj/IjQnmsl
3M1vp02GZcgkJiMgx81vHCdAMaQ1R0x5c2H6sCIL3diias19w/D71iiIS0dOY65K
hnqJ4rz2C5jKLOt9deXa/MheSOwxoZpeOJUfB8goAkPl9EHN8vlrs7nM4CUw4zcj
MwPARQOB5pkxwaz2So0rGUlRhKFVHdFisk53BcbDS/I50hHCezMtnsTqNNYGVo65
wX/jyVqYerTuMoQS/0AzM8kNUP48WSqsAiw3k1cqXgu2IJsOlPqnIZz68gH+zqPX
RIOVpZ8tQTmZqTfl6J9un/sWwSAKpULaOkCanhCXTXi9SWVTrMH/VSqgzr1pz3+1
rlwDDq/258rAiiG/hOrO4JEWPoAb7WQgGMMxCFXaG1PuuXUXF+853YaFV1GGY0K/
xlfuIgm6HRhaS2u5uT8bCIfGZ4Qvryfpa4LXaJFaWMzKq+HFq9r0bn0cNmRv2CEf
1WGF7DDZpT1pSnchxEQ+0tjZsQWMP3H36DyvguL/0U93pEoJihhQJIHLfLgxJQw2
+FM1KYNEjbptQ1hOBktddzib3O3KL+urpY2UB0CYiWCbKr8BcO8n9aDviGLy4tm7
bxecqBcfajJVprgV0seKZdBXR3vVxcRy/0xGede6/pyvxGCJXQwSBlyP3EtIGdC/
IyIFrXixfDOr4A5HoS2XpszseHG5l0VuRuKj6cvl+dUG1XwICuc8lEi60Fkgs7u9
Cc7lgBzX1+CJ+RXPXbJCGdlrqfFBm42NxbiRlTtJ3ICBQgifDmmGOftDaKjhAdwQ
Bu7CN9sVNdbCK1ma78ONsackYzQCwYw702inuM9q+28tDyednLjT0YbizUXW5Xo8
4X5hMJMK+RuEJN+gzwdu1HgOApmGp2/rWPMc5mbcqPy8Xct8KJlrK2sATJKsgZT4
2w/0UmwF4zFEkKHWD6yV0KJmrlDhUrpn8fu5ydqWVYredBRjVjO9ugWxrJKB9lqH
5C4DneMWRn0Pc9hlh2/aKobHeXJIwVRpytp9Qdnht+mbl3tDxO4LTEX4qvMsD2Jf
m6rEtRRsbKFgHV8knVnRXW8SYO5z3hoVMAATM3pX5cF3H2gMj1HbJaukVvqUBC+r
Xl6z09NbpjCDK+tZxCUuomhYlGHi0PBkBYAo0eAWhNM8uB6icBEsh3RtvQWPK81D
+8JlO47rYq2i6KPKBpxspqeJK86BvX1isAhHY3h1yzb66fbmFa7dIBjDIYYoWQDV
LWc94O3JDjDxXEt6m/rFdDp5Mnp0l8bCv+fBymArr5irukTqB7FUyQtnUvhtUc5s
uV4yj2J3YtjIQVRlYe2bMd+Vblk+8kF5KTdcQSTvCcdEoo5AxK7P3u2/W/Nnb0gK
Q/UHktLkTAG/4AMqx0cQSl9EnuW4XnTtNi2iggBlXLSg35TaIr1BW6vVz3ovbuVJ
OGIx4VHExOQ/iSog4G//o++xpksn3hRdPjufx1xqxqxLbdzNvgXsm+6DOC2m2T24
nwMXOMuQwbdB3QGmOI717yyGh12V7nhk5Ie/V3FkGX0+Vbv5s7dEEXmJ5CeGu4/t
SfCdGzWO6Cxvl7bjB/QUo9vK+dkqyMv3buRNO5m03IYH5X40lAIxpoDLFfkbIhgO
alHI+FaqnX0Ts8UKk12wDoPP6ihcHDhALnYyAiKIJdBb3eOPFNKTOHi/Wj/m/RBi
PLgymlbrGSpnlghXOy2gjN+nDHSYr74Smpiqu83SRpeGdo5Gq9VGKQtzYdMeAXVB
YiKYy/snBHhOb6z9JyZaeSqlF58USbNF0AX/RqRij+paT6qD2uXC14fN2DJUzXE8
uPgUhEOJ2EgKUCy+qWOwZASLxfrZjJMD7sUs3iQXaD/VXfLfyKxvx96aokOg+Nhw
xRLcl49fnh9Xj7bBluY3lz3tP3AyKlpWvn7F3JHtUMLbzRQOwTcbJJeJ4hO4opqZ
ktML+Mihz7/pX8omAS83V1RZiIi6RVXLZqL9Muuhz+i7BX/xLaG3ldqTPbI3Cnko
DirMxe4Qsd78j6AAtUC+ZAU8k9htUdoPq9UvNT307+ekK9p/f0ArzoUVaqpnkpf2
jviM57ZVVvSRMsX2PuzAO5W1AwEpC9LH7bomXEkaWFja+laTOMT59b/JWGivz8nf
rkUu9SMwm9aM2Oy47dwx0MAprkeRRyJDdEXcEy4DSCrSLPxdxDJdqHXxBNlYCSzA
esxvBlFTF+GHSSWJte19Koy48M8bOiDXzwj8HfGOhnae3dN6U6JZZ+OhtSsMu1HM
q0oyvmeIQeZ/b9wqE134PHvMp3jzmFlY30eJKy5haON+cD4vJf86F/qlGiQKS2hy
QRGjgAw95YiYXEsZtrQoKuuKdN4o/beYAhxu3YXKB6Sip2vwwgBH7pEUI83Fkmb6
00sqmDN2/NYufa0+J6+PRn9N7asxJa3C1M+acpOdIfHrSwFSjV6GBJX0YqBIHVfh
4X21dIYOu4nE4z1A7VT6MVx1dKVIEHHsfuFHT0AemXzU1F6VtB9bpjaOj8apO+K/
KC46rOWM0EKcZxm1PdR9BADNk4fHlGEhm7GJrh/1y7oy7tjXhlnPN544G3mFplOv
6Yp3//PG/pJgPriZt2cawn1o0TAaWP0B1a5htYgNLBrDuuHLZd1NVvyfW16Wig4r
KIUNlATUUXi9CC0EZqBUaqGMGIn5c9ibMkV8LqoddT9xyLmzEHxN2Q1m5+LqaUJP
hk/RVWpMuTCqSEc0m6zipurgzHSymZ4X32FIfLBk+FNJZSkDmbUXFIF6LguCpf+E
UohJqx4tkER7kZ3Ae5MB4dLYQEbQfI/2Tf5mbjO8zLfxmJ9rymD/8Rz9j2O/Y5Cg
h7Q16vTVKgyDBp5bJSHtycd0jynP42WoEIkn5kp+G4bEU6/kR3FG3dTcJzqTSKC7
XRv+A2rtSB3ePVX3soR2hP6q6HYIEVcb7tY+vUdUhZcsFpG6Hb9blQ06l/BqMz0p
Fo4qWJCMqkHFGGn5fCs4J8qY66dA+8Zo/0qTsrjk64gvOWfms2sdIl5RxRdgBjWs
0JrGpTCkvw+QJZDwGpoHS6+R02pYUNIVZjckCXUZaSMFuEmJfKgksa9trYS93het
v/9aaQLsyLK3znbPiqqiG8Ddn03C/+ukchG67RnDy6jtp+8iIqpFeHuxiaAXYy9z
MT1dHrkwwQlICjuGVqb9vWjbNcQAY+K201EUupPV+TyMRlSl1iO7U2oO2AEDj/ax
b3TafMvuCvWH2HHke15wAPsHM/qThzo6zoN0dIPd3qT7BZW1NJe6vHwiw0fjaZgu
fS6OqnnUBpWwFpmedZ5WD07ZmFvTINVmGdwP+wkpnCkissb50yCFHXF3oQ9csvU7
De29HUCGe60ZPpjaSfCsKsCZonEQG9u4uL6yWcG/ixMK/IGA1BU0mkGp87seAX3H
O4oKHv1XPsrz/ElEcg2lEIr3OF1thLL5xn09p/CgKqb3h+E07kR2DmrHBBltkCca
7OQa+hpFrYdpPGbKmYSfoOgIGDXiYqI+0R0aOtALR8Tszjhg4kUMRbc9LaBBOEB+
Ae4d8191Mn4DCCxrRG+8YG6KGT4jwZsK5GjqxCue0n6V0KmIEzTUEBRjWwEBHHVq
IpzvEiFSPrbjXC+daLysDerFxLAy2CjWYYwyexPUr3nw+5Yy1HSz3Wf7kqSb6oze
E4Ll3En7aTXG6G+/eEkYFgeWnFKXnhTu2qdHIwGIEEF2U316zmMURIDEbkdenXCB
0eqkodLfJk4cYnQMZQPlfaQi/uFuZwSDdVYIMId9SsTkHuBV+edJ22e8EKyKSXS9
8gZ/raot7zR+DJtf8TibrfiX3Qq48NAFA9Xsh7o+imJ+SXyhvi9fpUZUP+VgPUca
FdlIM+TOvM4mlvCtfeGSu+BYVjYpuM0uvvowukRMEGGe3U8qnm4sNpFC9+2fR8Wj
nkO6nCBvY2vcrQ7ggqchBuGgShoH/QqLWUzMCWzVfRebAUVgv6hEReJcZqaeIfVu
RBkeuEu6mR1lXOKh3hy1KN++ig8RAzv4LDOZdQ907g6q8X/GTekV5xFHA3ccUAKU
f/f3/9mVkKs1hNWCuiN+U3XNy/KwvGaDjZYAHxlojNiFJyAsHWVEwT1OuBw6PVd1
mLyrLs/Z0JPyZduSa8Fd9zBwVsWqd3EtlHHblFDXWV62aTTbuf/Pitlo494evEWa
/Wlsr6ceoy59e+Y27NW3u3lsptWG+Ub8LL1cKlDNNbiMQ09NG8VCUKaapM0rJZjc
xb0p6+onxDU1JnJvaxoqNCgUMVj2ur4jG7SaQWNYf9d327xFQ9hcpLabIGdVZ8Eu
+xBQZgcVuIbUQOcznTS/mfACZBU4YlzUX1yufe0wg68cuWH+vLNHS4Ss4DYOmIHz
Aq6b83PKkdv//lbYWxPh5lXK54Mv0UVnb2k+mMRyASZQngL5GAYveDVWTwTTHwrY
Z7yG0xvX4yFyTLkwqynfCqRFp6NsfDtENdjkrlIhNDQ6257ZIhoU7iyyyvk9or3X
TAqwKClb4+6tv0qZSt1YUX84iptBk4yvDyQIJkaZlQKFStdTlk3iOsnnisQdc260
SwZNG9PNL67He7nBzW6M0oTU/E9IhVthGIqjSxRFDyqWe9vZliDWWt327AYhzjOd
OpjPmULHFaPzATLPxjOjcW+2OyitXs4jeEuhKkHpAQsn4JiK7/CZPwV/zeWEYcDe
X/bX4fXXqwbJ1r1rid2fnmsORgtfONVEmRgBHIDxWxu6HvSNwdBUjl7Q7bJnzfOd
t+JTCYbLinDSoJSNI9k9NDzxCSm+GxbxEP+F+asWLn7Qt2ZFGb7XHDwJ0etpMTO/
AEqoDr8yfPe9Go+Y4X/9D6HATVEhkYZ1gDY30AtVt/a38AZqOpXWqIcXOQnCHd1r
zKrrxquOnxlYMd5jPI5a3fTvGqmpZf09sVRjEK8+QPr05upD95OEcq8+zr7uwjTg
vYuFTBGdHwmhPEd8lbLFJH1jM6Pt9F/fOzU0gJyu0Qi8pzA4yvALsiGlhxYfoGjw
ih1oDVGjpAV2FGxqzuEdjsZcXtGcPPM5d87PN8qsDVr23oI4GuXUFJJMwoz1OkO1
xxvNrLAGBH3vsCKSqbjUvX1ZWIZGG9RR6c/fRQ2SNAfODDBv2Y5p9YkxWHzd4xOd
Eav//ZkfKDaG1OB924jEbpmWKJ6Cum2kyvgeFQqjRvHlsQxtfsUji1dExvJFHoKg
Pzvr3upWvpGWf2oDq3afnLlzhH0AI5FBcWxbD7DmTGsrZ+SPqdJ5dBQt5QmhnYI5
6nrRjKm456kHIjxgj6E7v6JLScrOysJJscBAPdb8VuocawjhcCz/n50Sl/MycSLd
naMqhckXcgmgJ3QFEe7flayfFV/Ky2DEvp90r5Ay9+E9Dp8KW4jv/NVX2h08v1hY
+jS/lc1L5iFXGmmmxbrrsL72slXGr2oXetxqx2n2ACQaOzNF1O+7ZuNWu6Z0Pnxi
Y2p/oAuei+RDm0RcMxIxuvhc2qSi1bAQs/l7Ugesf01qd3zlRqTlJhTkyapvaAeq
zN7sNxuSEmdWml7VT0c4myXzdWNU/wfTz/m6y0c+rELLhCHdiAdcnY/vgIToPoaz
9VOAKXylY5vH80lgZs5by9mgiZ+Rg/hgyph6tCbCHU3IHUyPAysqYoThUyV/C91X
KoyzYcxe6dM8gLKWw/GQju6QHQG3SJ1gUOcbO/UCD3j/oblNJKapKYcaPF/u2egi
BvcAnbGY9UkWifTUfzve+s18779eZHf/+2uBKIsQFleuiynlAkXPfSiw3/YcZ1Qo
Ox78UOxEAuunLunRoYpwYbl9MenGm8VcDvZyuwtOyHeVw9b9rCN67ktuutneLG5I
feL5aOIrSgFwKyOZos0fMioUvVdrFH96norqr0SjutqoYA3WEwaJ6OyFTZV3YTDi
w0ydkzDp5Q1TBmRKSGnNdjCegP8VemSc3W9afquXyVKJ4joVSMdAP/LPRCLHgLm/
+FURW9b/N4EWVpB3+7GsklfdBnNzRfuo2Y1bZUHwFqiq/RNZJ+KAsDNewe/dzbaV
lGTwiwUXJ6pZujwQHM9gKcL4o6uCt1Oyhe09UflBTBco6ZiL02KyljvcyV0pebCd
BLqWJQ46OSbs1eSITiUm7dYQowa7/vFXUnIRLP4tIy8i53YRC30Ffea+9M7KbxPN
BCBDlObSGxBUdQxpLQoS2+wu59VoAGWPMe3rhocnj4hHm/f2J+ev77auYtETCVys
W4OIFdjTcgQLZqFdV6xLj2yseptVBsH89cqQKPyVfp1ziMDvyaxn+ZnSIpkTfvXM
47jINmg97dSmOboq+pDIbZYGjMC0yxCX1N0/JeIMZtq5lBngORDrqVCkwnaxzHbx
nv0rdCtVmJub/aaR+WvNJpxxRWQXDqYxC+7EugOSWt/ufeAbOtMkvCfUVgXmhnqp
vEeyKWqp4S+aw3e2qBKFAMOe5aTFDpu6WbYGPWNLEp5PEqfTc3vvYAvR7NtvhvSv
UXwAPgpg4QZrAsTO5Hglu/mCiuhO+pgnFoP34OHxYoEbGVEqSVCQLeqB4tH5tdeL
z52S4gQ9uFzCE/0ILSXqHfXZ0nrZgzEZi6zxYY1pU/bSFMrGLCT3u5nVdlMGzzqC
h3W40y6IxIJ6tFTUqd3sPsJhE7JAoH4nn3RoH2fcWbdqY89HpjaD7eg7E5mpAWNu
zGz3prND7YpAeu71IQndtEHNosOlN3690663NlX0HZq3D7BfT41/TI9SoENarcSx
JYWULEeW2B6ODqucI5gCc4PbDv5VH9ZY5naYOt4645Mth4K62ukp371ijep+y/lp
NxGB2EaQ6kiVnb+u/y/TLBEJfdwbFRPDw0+ilC2IJkbADDB2sGKdHrW3+P8JZe0Q
xi6llA1MMNbPWzKX+zkJ8W/azEdSaHLq90itEFiLvfJMq3lHyrqr7fz2ii8SUVtH
6CZ5CnKvmSrwr6xc/FrRqcYB3PJBzCAzTqpf7KFsXgLmnplHDqR/Zd/8EyXq1uFX
LdaZqHqnmjRW6UE1NstipcE/eXyq05+EvU8/JjkRsaAEBMoSCnm0z7zALQyggzWk
e70MfZtF6pp42U7IY92TJ/PV/uo5poQ6+4b5rG2lrzrMRcRTr7FIKcg2fGh4KrFF
MkGjCCuPyHldBgpJkvzw+BaIYrR349pn0zjCZ/HPDo9NuWpMzZMgm1RlYV1PyGu/
RVqwahtH39yWTJXlcsnj8KR3XkfBAzOQTG/j4kT+/h5XTbuNZTXdJg+Zuc9JRGrS
fvl0TmoEm2Cuj5WjEqR+aVTv4ezM2H9SuamxrR4XkpVThk2goGlqyj6de6QH80Xa
UYHyNA9RW04qVak72jf5DyXlq+IoZEDsVd+CdFzQQdvQ94W4zWFFYMVtmKCo4WAb
sCcLGy9vKL/qkHtmN4jJtcQuQYbxXGDgiiG3T8tirSkn1qrzsEsnFZr008/GuX/1
iCfgHwEVz6twoV2DGcNS3DjeW9gWT/SfoaCKE1DaAeg6ypK2RPhirSzbgM8dKiQQ
NVnWa3BGdcuKGh8GuRd8CaWXyv/9wrY9MqYePJh247wV5+mrn6iubcW+7MPFVmLu
97cnaFbwFNs8/2xZLmhY+kgMtHRZ9gOp5bEL3B8p1Z0id9xgmoOwc3vnRk5G7cpn
CJbKvvnORw/1iWxQ+MfAe+T3w5OefrsiY8Gqb61tOtDUPfB7OIfRz7oTNHXndmZ1
tUqplp49CU4E8W+7+nsDoMHeJyYjHw2vL/3gmv1HfnPuksH53P1InhFlopQ4QYL2
mFuULm9qRXSBOCoG6ptgTTqVsppBOfK0pu9gvEwCnlLrYzkbwi6SB6lZ/oHkGIXy
JPiQROhZ7/M8K3KTK2p7LOhchpnWt2ewP9f/hp5uH8qoNhl5COtlTJDv67I3RW6L
fLg8UaYdVghKLvoG6Bk9LrgB6NFc1Gn1n6vT7E66fC9haXIVdJu8hOco2uBNiSTy
OdeJeHFpp6OZVBDHaQoGjMTy7yfdUrl/RxXBVsMPOQT+/dCcZPS8njxYlRXpgqOU
I85PzqdfO9NTP1y8TAvc4I6beOKJ9Li+ZbhPFDzoLpA6iJeLR29RuCCZpecLyZbB
C0JyEnx8Jwda0Ddgx3INo4Iv4pAemncqpBGumCw0yInXlHWmqr7LKD5sraL4s513
J1XAFkYWcZjbPPuTDYxmgzESIaa7qrMrhddq7o4ojDKqmJlyKhLj6a4W6pOysElb
f1RRpVkr9lXgBZfQ+Rvu6P/CSMymtTsYPo/OloKBJTy8IIp+x73BuLeoDVztUA7m
UOmigxYskGJhyPJyUiOWaTCRV0A93angLwiTWAFCRq575izvloyhdszZ5PTBF2MI
AbiTwUUnQVouy8mr6BT+Pk4Bvbo2YRvk8bHieJJVnP7kmDkcmNDUESzmAN5SHRc9
RtyyWCooWu8jqA8epHVQSSzRmlltOOsz7FBuIjpn+NBCC/NxL5koSAlP6JUeuVsA
I4exTlJfaWnZ8/AY6LM6xt8wfRLwFpr/2MWOJJM6YNe6zjhNWV8/wOTr3LvshSmT
IrITuLZH6yEgSwx97815mrgh4aknjbrAAXGwunIOKfnz+EbQSFUhuy2/0YldYG1m
aZn3Xhmic2damcW7DVf3uizaGLV5y78s1Fb4UtLwlKXZ1B0hYoWAccNsYNR+OyKd
+sZ3YmbEii4a3SVdGhXatC+OIbvXuI0Yrao9F15XV85BSBvMVQkMYqY1/nZRE27D
mfnbeedjrJIN3Nj1P6bq0sisIdcD/8fJ40qBM+RXqQde8u6KuSfG29cqrBrfSbb5
SJZcBdSqM7hy2k29ZBzGmiE/ZRV2A1d866EqgvjKpsLAwBugsawY21J0w8lwIPqJ
n8xuLTXOAgs6DXK+z8r6FxzvKvXkillgQg2cKTku6j2EDnIlSI7RwkuvNLxOyM5j
C7CCrZ62DiExDxKuQq+VTkwZK+A38ON8lPmqC6QfZXbKlluysUBSgi8uBoWN27Ni
GkxQLKyaUjy73+W4AbFTJKrcQaQPv1Tic4R8OmzSn+JFrW+snmOQ0etdQMub85JR
BkgmFJxCUtN4KQSNht/plaJ2ejmODP8tG4XCmvtbzNCcQuQdtM9+HoYcnxy1Zfvm
ILpOjcSsiEVSwDHIeIu+IjLqFnYCqzuRwMD4f63sXfHve+u5W0yCSCCfdd/Ugw0u
KkN4LKTFx1P7EoYP2/SG6t3NjJl/2rUHFcX0dcVEGnV9W4ac8hgy7nFVNL2EMCsf
07YtQLbeXNKb0d3AVwx1E19I5iSilGsAVKrYQv7cp2PutAnR/MnWWyYVowMea29X
5wpZw4ZWdyd15/Ny03rCGLURu4bnowYTFjmel4XBI1r5jub54c6Mcc5NeUI7T7wg
NcsSjS3IaQwRGqEJNrUpMRL+cXrm+u9kQLk9TkJC68JRRbtCnPQeqiIbNoSk415T
pB62rxz0GjCvZrwxjsrN+jlVw3g0FL0T5AiA14+jN/oqszsCAjZDa1egEjHCNNuK
FPXsVJJGdQfZuXDkiULLKlqg3efJjS3sDN12gfROGhH/IxtbA33JvF0hcnq12/Rj
T9MMTX1Rr0iJbzrk+gCMsHaQmGfFtMTnqzD3FwZXB2I2Wo0XNdI3FOaK0BA/skdG
BCeC+QtZjUxlQuFaHr52As8OZlMmYfm9F4xo8pNR6MaGR2lslI+DGV71CEWCX+qg
CFM57zQ48SZRlX+RkAtINm5pZa36h0puN1sDL99ZC6eyabAZW4gJRafDqnmLC8QI
FCYwvVuC7vK81JP8oyfavCdq3fGSGQwEWAQdQUno9d4bhqGebXp4cI9+u/bglKIB
t9hE5RJW2bzgMwroQ2N0Bq4pfxOW+YGLwxnco8W/7aQM2Fd9lHhXT9iI2grX8jty
llNYYL3IdoVQjNsq7DM92szFuYgLZyoI/D1A36+A6dX+/rO+J+TROWJ5sTrVYXmQ
kcJAXJEfIkQUn/+KUU9NcL3T+/gAPjzIQIU16P+TUhOtpkjMuACBTwio248zCeV3
Iyb9WaLs8A4LNec8omeIHTSSdaocKLKJBcmJ9butLFIjf1iPpM7b9z0QGV6w3niU
94ZX8HF4u1OyCPYM49U2vxYXL0JaEGDR9IbhWXrfuwE+E7Mn4P9unX07GJ4ZVVKo
LFahRIs1QbG7HdrvfEj8ZW0II8R8WChkZBFZ1Bpg1Oa7Xx/T5tftjTMkjIgmaEpb
hd3ewBpoUbU9VZwfWUd06J/dmZsZiQ+aVtBdCSclKwoDfnNoQiYLwzkSnm9PdfVC
Qcmqed7AaZaz+i00C99fvjSstPrkaDlHjzAOAq6awxz5sxLJllcvex9wvTGmITRs
GtEXJgDmQxIvd5U9Q+E2nOmmEBI/tAeahGtGcnTmJuO3Zs1SnGD0963L/EuMzp1K
b9Q/t7hoBsQgN9T32xsJgCYRGgyCbJcpUdJOEwJULNBM8WZ1yvUhVsYE8smFqZ7k
spgt7H/VoCJ/JR1ww+rQRsfYVaq4g4wXDNdNiGNAdamIuCL/PsS5BfnPPS5nMuru
7+H3hB+oaEB73Hl/XJ7PcWLKv43ocKMoGNoHiqVlhdTVI/bySdeTDB0jlkIbZAT8
PSJ6KWBih8pY02PltcnNSQBu2RZptaBIN//oyvvzuz43nU3M/S6302pcyfH+nh+T
w5PzFq0VqvjPvSs39waoE75amNbIHUHV7qQP9uDWalUEcNvgpIb2Mur0Oynxh4Gz
0CP8hRPUJtk36Vp5ZLLd0VRtu0hDqfJmBumtJdUjJ62ddcq/NjsYrGVouImdYR02
YpUsxG32vCIlvaie6YdvTPQBexT9RmQfn1ZzkdNAIqzCahosdlLxFZPL1tNTAFfb
v4FxwSWpfQl6lRYIJLKrIF9eCmeiuGZh1IClMIHX/qECIGpuEth1uMupBlM+iAgP
te5VJ/jF8I8qUfakFNamNyOCoMwgt1pjq+J6ERPH0q1ZITTUQUOgk5zQgLa6ttfN
2Fn96+WhiJu18bSlzDlTd+Tur3koTi3WBz2PcZkgb/VMzwQdT/j8TPO89unZG89F
UwHQtCBPtqAikF9Z/1IyadjEZb04hdFMN8njXNW1XS8vqgQcX2YUfDG6Ng6mPHE/
5Vgd7fVn+0E76bdwwbGve0XWlOto5BA8+6UxHPlagOYRq/eRGRggKMbZO/gFYlju
jyVfS0oTpe1dwLerTSQEEwd0SRQ1Yt07xUiCl4hi858P+K8nqlnQj23Ti8UaJsE0
aJsy6II3x8LWsn34DJhc4JogvZVxY/q24n5KBPrV/UaQ4M1YZIRS/xojoJmcBl6C
meu6wawQSGS3+V1JqVYUwIrs4fSY5kOT1VT9bR93OfXmpTqnWoUBUbzQ0lfrpf5t
zFyCpL68XN3jeM0ZWJBQ9NOc+rbxZAw46OsJ5Qfc/4/H344gLvZqLjygzKAJeD0G
vLaXFdThKT7EoVhTl9J9cmP7vif9bnvwL49b1Eq3wRyOflX21RyvmMF8+e2Ifcsd
FPiWkKzIBa6TeZPqvg1MUiA7UvdjKCDqh2TnPFXcw5OrTbTyFxqknGIN3aO/6yQ1
s+DHNH/I0JaoKsPF04ngk0YQm+GQ6RE4+QrYoHllo6rXMjye6VcYR0GABTiX+lEP
yuEZ9Cc137+r826W2EhtZ/APiGNOghviTpSgMRo81anrUqGD539Ts9poFFN6k/+l
zYcutk+eJ/eqZ0j3QD6Mf50w1zmLxzKkleu3Q4E8Ku4ZMvmUszf7XPPdUSc9x78A
Y3/8B5Dcf2Qi33oX1OqQ6TkcFi4Ih3Bef6DhMn49799Cv/3miTP7S52K7QRE7ZZi
M21djWgDqNs0pxXhxXzAKUjjU/xZ4CYkeKNBEtUNVHUxkc43regAxycZT3H9VnIP
/iEAs32m9ZI5eoS1pTKrbpiiI81ZGOcvv5yB5UqNkeXZA1DBniGA25UfRyu1twyS
dkQ25UlqepMEIkbWlSG3bQVZBaH2au+r9l2KMDy4YsrWmxy19MwswVLMQMA9rkeT
85jVqAVaTe+7exthhgky0ikWRUz69SLsUPihjbWPbcE5Pi3diX4RWQOojq/CuifM
rRKQ3KVd0A5tdH4Ka0sD97w0oRCNBThCy5lZqrHdOwGTtQec0yhgr32poQu25cin
r6fe5lZmcSlPsuRCzmWhpROoyTx8WYaholOgnZK3G3pjMkuXTsS1WYJDw+1fiPXl
3dy5kp9nIA+/94Msyx2uT3kMIZzs5CLWiI8FWmsn6UK+g7n4qcHL6M7BW4yEtcM1
HzlIMwdwtrbl4wwNxtdny61jTmR0NUpazbRjHZOsE1vH2lvsPUAOQVygEsl3JX30
Q4ib2QaW0oamd6g8MlvnlYBYYptX6yatJYg3LrqzVYqiXYcI5GBr7kU4JZAaJ+lC
X/MM/Dw2RDz37GYsi0dn9xGhRZjxwN/vgX8WMSNg/inczg4Oip+YslQTSAkY/46S
wyevUDUZuViCiETxkZL6rlinfTLcYyCOsbuhI8oN5yH29Ah0nxSxPnHHIcLqCJFk
vxKnxKgZrjpYiNVUurZx4eW7/ImP7NbvvGcUZWlmTugruoh+e6N+upcHQ5Szyfjb
UuF8Acxo4YPNf9CJt/GlUFT79sLjPFV/K1/unTBAH2+yst1HPHzZ6eTbq6rBQX/1
wJeqrzvDVZctXmqcnMuYqKyfrNXs4cRaRrDl+9S2JP5S2uigidk8tGJM1yzCZVll
TIBxXbgD/zHOmspS02NSZRGGij43I9nADyOS0DpXrNWmhnJUvISIxLWWaZLSdX1s
f/ME6tbBEXqXwgfIEBVTy/whnpNYLMmHBz9GVClP4DY2wqx5BWbK6UBG9P2EgSmm
fvmXD56vOK4l9I/Ez+g1cqN7ju8fgsMsRUcH3TWwH/VZvE1AYdd64Qxq/0sJ1hH9
fIfCgzyDt7MRhh4Xoh8ny+dopJaIxVafRY4IdrL5kDr5daFDhjgBy8MH7Utb8QHO
LMgMhY6gf1TcUt5NeGxThzPTViS95koTwiL1IhtY8TRMq8m2iUtEeFYj5EPvlqMR
FTi0dL6le7OKfy5AVHQhzU0o4keaQ+46hA5NUlgQqyS5RULShKZ0cSRq9AAnaX4h
EYMr1lzxo13wTSSxHQevCqsnH+KESCozN+aPlEJ9OBbS0wnFYVjnbCsC9+Co2t2U
cDKwmnOK+ZQlSq34zV/dWhXo+FkQXT5T1McTZ8jB6Qhpx5OTf8ucwNadEQd4jdO7
VQDEvSsjP9oBgJDAHQ/3V9D5jEu0c/DpAqIBSZGsWFGAf+WkSLx8zurV/aNu4ZP8
e+Tlwk9Y8S09P/T7kE91OKHA1KW+ATB+ZyiAY49KiIp97s6DYZ1juZ0CT4A1DClx
BaE2mNcZvOwMqihjrQSOUkiEWvyBzqHk7IC9RrRb/WFmOOc08ucwd+tNQH6dfC8+
ShIf/WEB3TfjA0eR8nC1IL9SLXce0ffsXAwB2f/hgKNTVG3FgJFUX7lGBEr0dQfp
CZcWu3RajqoILO1E3znhuNKivBKzrlOifnE3hhbqXKmzTHiU7KiBEnd3pueGE3fu
HNPFyagsKL39NmBhsaVh7yRjib37uuNXVxpCxM1CziIObfjGV0xNUnBRZ/hy4iQF
357dTvVNVmEpURfMqaNuXvTRKJDR9luqG1Wm3UQjoJUGzZ6zbXtT0aRWf0cfsgPh
6yroPcKxSd8em1dBSYYI/00lN1XkHjbafhRzaw2PDiELteUxqXK9Z6TXkfU9yBKn
BY9gTXoOk9tXSYsGz2GXKovAnl3VJM5IfyI2cTnTQap3iCPBaDPNO3Kze/B2OFA5
genijAYgKHiUDhmvHgvn8LIZ5ZkyYK8JW2lmi52tO7CiPXptNIdu9h0qRBV6qyd4
lRj/0e4M3qh5xAERWH/FdlEUUqXfxxA3T0dCRqJACNbuo3ORTeUcmKa0a1SabtXp
wtvVrVf/vfOXRwMEc3XCX8JQc6s+apuJ2pS+Jw7RZXHbJ1/C6nUPI8OT1Vkxg7zd
OjpRqy83hh9Myaram8+Sou/AYIKVgV3AzOEAO2Dmx9BgAj2h/loO+P2mGZA83JrH
jJ2d3OCZ3roXrAwwAhkFfxCXrdckc7XvoQptFG7FHtKF5nIlqdXWZF1HgAvMt+li
K8YLRKK0jIiwKLH1xJAIcEnAhyGz40Jn48b+KmZQb3of8ChA8lsrSKMwGXwcOa0/
SdZZqVQbwowvutXNjHAZWQu66JvY9jTOMe25pwwN2f5Y0dQLu5/dI5v+Iyn1ECz8
gQfS2TMRtyerrv+UGUbs+Oq0S0XHy8JspKL7I5AemK0vMBHb0g7Vs4unQkIDWCqb
HspNcDZraHNUxIQV3x8lzA3XOQYSbRrPMVBNk3JU4m1as+4TRugWGhs1u5DvV9ga
OhOUi4CnAgxRUMV539T7AYx4QovO6UDXt0771RpJFiRIYxyE80EDdasEz1nF9mmi
hNS0sXM0hEBzmHsPDG+XD1MOsmiP0Bx7FEor3hAXWNVkACI8wQobpyuw+IJdVdvA
GdHVXIN9wXu82LmzvQ72904xaGKPb/YChHORQdeep1lb9oEpia6RZ13vsmryLo4p
XY3MPMSXou8jPmULO7VCncocRypoky/ol+LiLYJgl1bBipuqDzAX2mcTN1Mp4kjZ
KvGfDQj0uqOjwpF0DDAkDrCbJHy+eQxbuMQtizo7kWPW4riUXkGIGjpZkIFvcKfX
nltlRuoPnui7HpUIaG5nJQSUL1NTKKlO8g1u8ry9PzJeHdLJVz0MEItKyMJEpUcw
LMCTZ4klbY4LIa/9t+PxoCr+nSkw5DOK5j9QeHCIH9sL6zwSegrytk986om70666
zi8SQ8j2K0mqd7Mofc0Dj4tyMVrqb3c6VFNk1aFMx/ydauuZRjE9JdhQM3Kq33el
+jL7shatYOUPl3Gm/53Y4Gyc6ArNYkloXaQrNOVopAkFCGK+3IAmPTCsLvRDwV3f
K4SWt2zgQp/Wbhawqkr6/fqW4KUSmenItV6TCzu35C1bsQ7bJQMZfvnx9GQ8osQl
R4sHFUEbyvTwUR997E2EMHe2rs/GUpiGWZ7RQe+oNz5yzsRa2JeJCbB82kECOunZ
Nfx+6LUYQHj6OIes6vVtd8tNeHRFK9IBA4O9OL42osK7IZkGoGGZNiP3kqcvpsnK
lQLJpQIYf3jqtLQQR2EvlyoDUKK1jJYE3p7WryVK2ttx3yFHOp9bzNgz8VUEzg9S
jM0dEhPrynEeDW7SgBPgtwae5TcSG+39Z8aP0cqpxkPuBnTE6V8yf/6d6Frv529Q
4SfVmHg0jaQGhupCSB6jNhgJqJ8R6XO6IAeskA5/0V6vbz5a2vJVCV1oDOsU3gP5
wIMtbGb4RiLkch0ZiEhzthQFwBRtSUH5+FGbIoxtouBMZorX5zTz08xVrP0tGzPD
ELVVqIKlT5mszi0ck63Aj3EpChHla373Advv7pNU0WQ59Irg6Ip6+LHmPFLiwUvS
Ig0HpUAf4Fsb7tql/ew665dESPms9GJ5tN5YhlFxQ51OMpobzkkyTI+pifQtDUiV
ZGtf3geRXmxfjlpinI0NeLeT16Y/p5lATGMJkhb2SXo4vT2TVFz+Upl6kaN4K0Jz
FPpWHwJH86+MbDVCDvko6/X/08wK3aB4X/ELy2VAPSxp3D/u+gqSZXaJtSOaE+oW
pJrKTXuvkBXxoXX34X3o1b96z37LW3uPEKs8LvAuUyJk0aE43tCrSZRkhtJz7CbN
Obk/bxHdd+acMPHFczMfWEq6a8rzl+rKx7zxc8QKLPl7t2Un5gWYO2hExGlEDI1D
VI/L9Tt3ZveeDleXdw2c61qhizbILmGdY/2AHHNc2BvGKMLEX2bz7mnK8vRBBn9w
45fw6KbQaykXocCfFCsu7VQHEQ8d62TIwCjjM899U4seVKromLf/Y8XNHotq9HUy
ojDTu6lDcDQKKo7r0Qu9ktiaujoof0spsdV+23w8CQK8MvL2OuwF9APTmbBhahEd
QlTcd+CAObTvrfGGTqPbPJkMB0rjsA5ls2WiWjbNKZguAD+E+hquCjWjRmLpQuHc
Ea1wDousq6+4XElTpH5Vx5+yivBVB3xFlRnU/u/Vw9Wf4bIaOmnk+LR/kr6SuYRJ
VN8Mq4px5z+m2HxE7roP7syXMfr2UTXeq9wJPQgZH2r1ZWTPVx2h8ZKuiUYqncHr
IRV3VpZfgCWhdkadbYqIptdL62B8nKGcrX+tVZ/KQpW5hmgYq31P2+JP58AOa+dU
Uc5Ruj1ljDiA9C0tSaofM5nudoOrt94s5SLILTJch4zsjhgLtrBPbu0ofLcIpYso
629Uybt2y1iDju9p5AnnCF9TOedTi1YO5DoEEPrpE+EvCPZ7+WekUXAUvPgTvbh9
H99dZ9d4WBWmUYUyTIk+plEQTCYxQQNdGPH3RoK/J18YHZsohXBuFqpEEH58u0oP
/6CKIkBMHmesrWj6l6RXSCMOoo0OJWEsqNdWLewZICxMkMQ6374HP4JGc4AOEh9S
WXtpe2XVBrsblM2OX0gGV7cPnL/cZNUBAQeGizEbAulLx4vZnXH6i2WDo1B2vW5I
o9sln/SfcG10OWgy+E6/6OB3D6KNQZo4A2vvH/KFsgzwX3/Vli+lX9RcHoEtkek0
oD3zP740pqmtzNgsghMNyYNHzxAafdDhB3oNW4CHgHHx6XG7s6XLIm0RZynqzcHT
Bc7GJDdYEsQOsm/mPOguGx//QUxgjmB/KzOa9NZjH6kra9S/6tyP81Ryy3OX6tU6
HsvNZc/EIMvXgLfthCB7iuNtcRuHWqK7DssRDa7shTDeeD4gx7fDuWe14CmJpeyz
rRmT26kohkn0gSPo1/cntpListfBMN/B1EjJ4uIFsEt5qCAOKu1mklOE9shhKTuh
v5eMTsGR/Ag6YDL2qIrW5iiRKvA7ob7yaCUa9E51tFvpySDqdknVXLTFJSM+zgB/
QnteNbp1mYgWXJJExOWUQ2P+IUmTGZ7/p5gInV6I2KBVdh7CiNhYntP9napvbn32
GXCue5QtstnrQ+xD2TbMC1nypQISJbRTaAzeITOlM1PGVa1aQooCfCDX2Xp7Vnfb
seNVT1qrMUDclPrOJSa1BBfcNkWX5wa8dQpH/7o1yFrTvVzLVdbBJgHd+qCoRqv3
vGUyUBqXWoVjVXb/2XJCbDh3zeL3OONZLHjYJLxXF3UwH+ZiGolX8497I+PIu2oZ
N820xS7Qti80Y9GWpCMFHCRaG9XjkaVwwTSHLcCuPxZuAPFseWvW0dzXq1ooyc2i
D3K2pSFxqf1gYs5jun4+YUMd4e9AwX4yWuBYJiaYOa+m3ENNDYURj3GhAUsthn+p
DGo4/lJKujOfQ+o3e4oQWh0g4Bz7HoYcG2uxNhtUCj+sgaoWwGDfX8REFRYVTvag
PJOJPehRg43cGusFZyYGbJtBHIuFsN1RkxMIOQDTmUWrnyEmcFkt+mAc8GkLbGe9
YVhForN+0VvNArFzALaj143CIeAmEt6/1XAows96+J0KlZQ5DY70CvJF9vez7/E1
ZsbKXC3DgmVr7nUNNfgXLxRxMifxMVN+FSKGzN/AJVQjrIKYqSs1gtASBr9IruEh
4iVTbdND2gl4acwE6B9e1RNWOLzbxc5+3toz4psG5du1NwrHRBiZssjpoaat3Mvc
0/ACXyMD1nrZENkg1G7f7AdrNrAZKStxEhJuAyXOjh0l7BNYQozuwmcq15NdVATv
xjSBuhq/rDt4ON2GyEzkle3mgPLVs5Ovfm3tqVFThMrHYLnJffCoSOeteQM5bI+o
pqGX//Ytz64YZXoMPwmP2+cgeZK8p/NIAT2/vcddy2n4cGLIaVzv3UP1AEO86PS7
0dT6vdTngPZ/kkgkwNIDcstXLrdyrJ+3Zqj+NxVWyHrVb2fuk0HUzC1Xwnrf6EfH
5/WKtjjgTN9jlrUfVPU7aAcM2piG4fXYnVayc/Pta5vMRBRAd8JB4OH2BSaplWjg
odUvfxd1SoEdceC8fFc9Owy24vHBKgMpD7HVkXRVmettechaT21CSAJz0+3E+1L1
q/Wm76Mffz/buEdWyPIRcmXQ+3waCkUpn/MmW0o4pXpj9vr1YskXxtdkIbGJODwS
sPhgd7Ds7/+Z4SD+VC5kGoDQPMNBMknptpyv9k4eAs45KYlywjdcJRJaKjXLGMSd
mSj4Dee68WlvweOA4JYS0vlcvFBYJHKPEwMkCAFyUp1VDi7B22a8fiEwe2cJj8lt
85H8kmR0pZovAgcm2EF8rtonQneDadsMOs2FWRMVJsYRExw6DfAz7wPy6c4kCh8F
M0KXf2MLxEkUaQz3t2D80BO3g6Tqv8vwH3TNHMrRAc+5qRnIuKL+LGKPtRKHs7UR
PArFhcNbRE1s/8MeMSxzjnnlERM+w5/n9ZBckYKtf/rA/iLKruJLGE/qodVzSqcs
eSxLKBbmarTGjrFORYHSN0yD4a7DFz0S7Vj+6RulteIUPhE1UtoB7qNxZdiR0Yij
tWgAFLcfEQf07GtB2N+40NCWSEYPYtXiUOUL+XIN5wyb5NVu7Se3pIg+pUk74Ajn
saiW0zS9IMEcOSAVrNJ2URfwwb+SgifiVtgr5w7/3pJ6JuKmACSBFIRY+STGB96v
EkvWL1Ikwu4RRsixf62lK0dHYJbe2jtBb3of6LPYaAreaius7Zu33pu5WsL1mEi+
ZCE7fBTomSA/FJKOnD4cMr5JeaI6bBBf21wCpkfCj7zQOEEeiJ7gne0QmZwb/F9k
7Cj84UEMvmh2p/I3D0hfgqEcoQjjrNOSI9EAE6T6r7A4HwiLPvbMHO3YnRlmecto
U4rLZEAQcyTtT726Cy0/p6eJNkxS4qWef11ugHxQgrF0d5RfrjwMR6az5goNGDad
csYXeRfCU+e83UL21Z0BHcofeTTynHTj+GyR3zk5Fi9jXIN5mrpQyLm3JhKa1sxH
IR7g6WBBDrCGtMhGaDSujuG2NBfvxzVmKh5Be1JUqT2GHADzBYNtpZUt0oYe6Iv7
9OT1IgioQu59VFBe2LF79b9XF6khzSvcdACRmq5a6PtOpRZ9ITKL63+cd3mNGkk2
WZ+r5RY69rCEIssUyoSIkOWHjAiTubnXJe1QrSj54O7zB/eTvCZPXgJeoMa3FYka
Q/hRxDAIEYPlS4XePQZxPI5lEvVJ6wVrMyDGxieuOEHgKDshC+9K2dAfgXO9F89h
Wee5h1ZLSrETo9hesQYsjaykRVYuX0UsRScJidb5+aRvdrazuDx41gB6TTVFZF6R
VPCTulow1BRK3ZpkS37BBXdZqdZlnGX7Xx2hzg/L+I7tN1G+Kzq24ReDclIHWOX1
BNYs8CjDztQg/CMF34ieIaXM7UVtEbtKItG+A387wNTC6TulDVRPoMoeoQy3InLG
SpZ4YNzlRPUNCQZawciIylvt+x6eY1j1Dk+PR/0O8a6/ynhtFknPP80Izrt8i0BO
/2XnlIXVYSFUSwTVovOA+VxRMbt4GGLJ9lOcbufryXzsElG0kGWRpIoDhNi3+YS6
A2wGM3MPYnc12wl7VvxV33rwapK023da11VqaqjO3x4ZYaXRfFcaFoA/MTYEQuAJ
jk7vLLlDWQW7zGz9YBsvbULoHpFaX02mrLKXJ0SsnGN7a3cufhlE/CyXCB6MN4Jt
Jy0cDV93EQfslVe+VY2TXfwkGRFDCsV5LibjMljmeDrNP4Thm5SMUIqP0JP7P3c8
Pcn+btyAe5QZhHeuWBFCiSP3zJnpEoz3kRnA/GM4Vzv/a+mfwka75AXcKV/fwgg2
q7WE5fkLFNlVZo/oqEBY9g/ruDhQDwkOwmZHj+QVGJkqu9crARyNb33coF8a4E7w
p2ThLGEOw40NOXaheCsSfUJCURQNKA6hY2uo9G5q56SsIHchGWOVjrfgUU3a3Htr
y8W+oKDKkpN0YCle9DhCc1UougEG0mJl3MUEyea4c+cKeSnQr4Uc1OXPArYeTv5D
gOJj2DPIHQ5IaP+wpuwYD050YYEnSgEIJyL3KzLUAtwOkOjTLgBbsFTDcqLt8Cp5
fvS6Qdau7SseAvKph67iSUPEXTYssQgHaFkak2B2/nYrkdv9IVv92qClBmq+MZxB
yzg0wyLNNurDuIjq6EVwIs0AEh/QS3alK2dcnw3YWSZ95ZuVTfVAsIVqDzVjdSPh
oLcemFXWwFxMtrXs1ngtuPjx4QURGVdT/BiaE7xY2je6yTiRrG1+VbIQGPZ5vWv0
3NNsQZcIw1XRljmZ0I4cGID0ulefg6qiWjvpqF9Ta7t9G4ZyS/GIJowboh3XnKgO
KcBW+2SqNxnP4diIUZ5sPn2QImmSq5rw9H73KGrLMXQFNwLAsEvd4Fa3TNqkZ9XX
7SpRQjyZD5YrR1xkDyz/VCHKL3ZAqeveLGMu6A/4RjuVc3UyFFv/dXGPLluKATls
Ij1yjv7DWV4zIOxX6eJf2QKuR+d4A8IihONPELVEUOKuQCFu+5na6FHh0sZtBHh8
p1bzI2bN59as9M58lXmrrV3O2LmHTP8At3v+Qypk6tbILYRjfB/4GDtB78+LiY66
5JCH1m3tP7CDm+AIQ4mPVDKpNjJmJCQE9W3sfIybGe54rE3fYy+9zKSe5Avww7kq
0zL51+y+6pAh7hfflyiSE4OJGWmiiwzJI/nEaVv/1G4X1pPR8mnFE82ziM22+5EB
jmTWlZK0OFDEba+v3/dJIIO6tj5kQBynzfcVpbtSuDX2LGbZLdA5WDr196WnGlpa
96Y6/+hXC+BrLizjTIDVBJtBXRxvQ3JJHnmRjbWpL6atgfKIRzIWgofZbuyaTozC
S33q0vm6FWvdvYFuxkj9A9GWXP2RzjWWmyLsFg9ELcz5/HLfDuLs33u4HM2KLFlw
H4JGYdHxyVRCT4g+9v2gkekasxQHEPSDQXb56s7ltUAnjmuw1P4v6IMECqxh7zhM
tIPveyPPg4YGv9Ww7jY8TG4J9wRI/ISMTZOxvKjXqg8FuLyfsWcq5RWESIDh7pRG
sLGPieEdt1oJ1bvOmRxoP9liLlX65NBMDdf9XyWFMCj2x0gt+6Psxv8J8CIM+A6Q
sWPlLOiZgpcfSDmrldDgZr3JOKCMSmWAIY7CatR9thJch2LQ48syltWy3WQErFPV
HVqFwJKs5v+XBYRNcNpZh/lEjPO3yp/v8YJJIIGoaIr0aAOX3iNKoWTFbeSbeb2p
mxp445FmIjqSNtd25/2kHbU/vgM56eUpyPw857XcoRg5xcfDExmJHjJ0dgsJQ//G
wllAuxgPUusMd5LypxpW5wiETqMcrH7WYRxk2aMaO+2f9JpovSNHpm2FjmeNhyMz
hHRPazDyJhd5LQEOo/3hntMapC7NOaqGpahmHpAngACpH4cWnUIIgOEqZXIZfb0e
SDBXlBarNrke8B0RIqnM47FWXKwkIh1bmYAo/ljtVeFTxTkliRH1hoBkz5RPU1Tp
zE9Q4MCFDFHEK5rLKF+Idk7Ftrb22CjXHpKQkvjt0S0vyxscaB9cjpxQqhZ65cXt
e+qXi9dBd0rOd7UZlg5tjwCkgVq1y/9NNajcpVcVCUczoi+FOJpCFJ0BB8XWTz7s
PpFTXvqN0Aha+3BB+Z31woEgZ1jUo2ktK9vsgJ4q0n4U3ZSsKHVBFjGsIWRlN8Ip
1u/YuL6+CVAWKakW2Lsuwj6kfLoqnZpPMoaWy44bMXrI6sma5ub+Lz1KDGLHsjd3
VuSSt+LxA+N7QQ06eOh7VLc5gD8K7JwmThscsznXQvuwKT3iMQUemVs4NouZZcT3
3RiilP8lZORFQW9sqFUcbedI8N9dU3nOJSpB8pY9mNYXnMiujZQyN2NxfhouHiUg
7CFS1B3UW5VB0fdeVK51Mttzs3MDWpWklRjn6o+ZP+Whv+P0TtOoT78yept+5QfG
DrQ1hiF1ig/il7Ydzk6nt5bdULiLL5FhOiYmQF/TmyMIFpljKdg/vhrgK34FpyoM
j+VETOHYvCFhD/F69Srq22I0aXK/9ZJUcEEUyE4TIfEJOzz1abI4IgCaYySlnt1B
K9Taoe4XOVvCyfKhARf+YrLb7hZEylOVCCKIPaiAbFdq0CYe5dzc4u62TCS4Xmad
mRjop9+XC9M8Q0D0hvPQfrh7xxl5vws9m8jhP5VPftxrNahmeM0mgiaB0Cru7o+j
3BhD6te5basR+Tz4QiIknnmy+MHUdoP3KR78zPFTdOV3Khy1/Yeom18mLVvKml4d
PUQxIfAf+6FRkHSr0F+5kghwQDZlIC7y+Ch2/o2R/79KJEyur4mEMs1fZzeM7UIN
4TjKwSE2TMRCw06FjLuVU5VS/SV+gQb5f7nb2wH6FZ6NIBLSP4rlgQKjhH3M5kqC
dCQYyheFcbU/4f2CAU0qD0C0jS0moFdyDFrY5k76k/gxKuSG+7Jx0jpMr5QTxQvO
DCqN2ocUFOhAt3pqeA2P4ULC4DVJeu+uOqDx5cXO9jzSUF190nrE+QGBXcubpCLp
05asJbCnAhjUaYf6ReDRl970Vjua3WkaKWQfvh3vGZA1qznC14CiIemZiSsZLvwZ
7D9vtfBmzcDkdSXUtzHEqzYfZvWhNwRLocLUdKJvufjXHU7wscR3gqpjWDFjPB/n
LzDBv57csd+c+B888Vxzsa9ajdzjaJ5FVI0HwCReCVpJAm6yF84HgXIw+x2Nt2wM
F7RcNtjQKhUGROK40shH33hGi2RLS8xvqJG7nnLQZFZDlLTZvLfssEnGiLLBsrrn
itS/0wyzd+UV819v0RQylmgR9Av1yA7Hc5l7HFLhRqSyWtl9x0e5wFzfeOY5rDup
txYvzGQWh4H7Wp2zyjSuXxBDL0gVZWWrArmD38xIifCf7Klcz2xWDNvepp0GhpLa
sm4k9kub9gyybJwLkeFvoI4Fmg1W3zWWYtgSsrW902iEhOStjPreYqFnXIEi0Rey
4xQWVUW6w0D0N7NKJI1syRTOqEJIIQJxbhqkT8e24XaosQBiovDM3KtRAdG4FwRw
DKQL+zpH9Rq2ah2XpXNmgYq6Z8N9haPrNbWNTwpE0RUqWpM6S7I7JhB/xXPDhHm5
JnKXfMpQtwHiMiI+lUm7Xs19hqQfVP77cecxUSyhMx4YiSsmsAPLehapE1JW/Ctu
DNi1m6MMZNGMojkgB0b3yFYaJhq441RDG1qEUv9jB090xvwJ2NQdS0ll/4AA0DJo
pD2Dkw7IPskBPv/RBTH7ZNBrjody193/pUXJJreG2DqeYlFVUVXeIRPReO2o5GXD
r79Z5++e7cHCUnavqLlwaBFDYflITq04czf4mO1+MSX0dTVcAAB9xtULrE6z01vR
zFvB47K22XnDuYaV0x4dvOnu8SmUJpsywEagfYjmezxa7onn5ylZy+zRNswliQ1h
v2blL8g4e5YFrEbsmxYG4USBAf7p76LrBNn3tInJ7BzEAdwF/Sds9iVn6FhtkjJs
LCqgYTe+EYItXwlp/3PVvA9hQVAVgG/77chzQ3rnj5Ab2bfhyvmqicaCOqb2FDKx
xAFVLV/yZbUVWg0C/rtvj3VsW8yiprzVVCM3bFEFXXx7HrcSEX3fqCARFHr0tpQ6
6/TpMr98wcpOlMJNO4Yg3v0ZlhiXR3DMzS7jMRmd+5zTEPCf3QRiua9DN4eGRY11
HMclC5EiPmr+BAQCy9x4xD31hjnPRVdslc73Tzm4MmB97CUOrAjA4WyW6pwyH6g9
rqvBcQbsWueeuaU9PJSmAlMzhoqmld3s+LEnLQFuMBacM5g7zXThTgtHriKFTZdL
4MRdjeM7yUqaidGMpDbb1H6GhMQxUGjYeI/hso93RzoLjp3YU62amGhnPLB2h6Fm
RX4FL3VTxgfgy29XttC6wdaAUioThF2B1PNh9jtDSTMAk/epTWU7ZiVdAFIztQdF
XKAai6/DatFV964CKWwGZsNUxDSBpgGokcTCYokPjkqlyp1eGqtO/D1K9mqhyaVD
wj/oU8q8Mx7xnADTrWQt73rabF2GYvSww2NVChIghlSaNm22m9pRyXPrJpT31Q9B
m3DERCHohPtEbBkuIlBM9xGwpZKzn3nPQ6wvBoOcWQKDJfwub4sebLTBBhPqiDob
+ktEWoVEqyf8UyL1Y3OrFlPByU2qmqNputMsZThCWxKBaIs+1ESkmuZYN/cXWklh
TD41Ttke6aaOalfXMBCWkLgvHRqOLwpVchxGpifyt/5bcqinyNeR7VkxKt9Y2exA
XCJo0Uki3izds4Qgi/c5CnQhxtbiNegrtJIERu1YfM4wynW3yVQOx3nSMEg9L/E0
PufzilaxCxjqPvucP7FuFWEnzAYX8rlTWweo0xkS9gDIl+BFb/rdEETR9h+bPALj
32pwmfGlTjDsUgbx0+ZSkgxEzpwxKGBZvOicagxaK4wEX7XaH3j61ospjd+QWndX
x95YX6SYq2KrVwiyjloimLPW9sCGSLRNcpSHT4W6QDpUpcgqI4iyT2jXc00tINpQ
K3KTrM7kb38t2IWtMi5jvJ3ebSfmeKuDU+/rd/YHbsm2BafmJUMs4h4xzWtbgNGH
0l+OBlw5+i0XLIj1pm3BRC9JgJBf8MG/y8A5TkugREMQhJzpw96+K1yuCCFMOWFr
5utBQ0rc0RUX94Csbk1dw5URYC1Z1vSwxGiqpdhfICOvoZRNLcRvV8P/8lc90d54
fYQZRj4xUmY0SCgjGu2j8V6WLUwHrtJpJoLh2mXIfEFNtSoLfLdgoPVP5VYTUd/H
4sHa/4L5VO0VbKHizh9lKBLgruKRL9UbHSUqJstoXc5FcYDRF2vJKigJFmDH8NGi
IB0qR/9FeWJdSxDjTI76CDU0c7KZ9+bkgi/ldg7fW+Ij5R08TRYilXja3Jymqi3o
5BC6GG3d9kyZFrhkRKf1DGO6NL0Tt55fqAr6+mS+RzyfWuw90BRHCvnvVus6IvW2
MLXNfJpnKn43Dp60v44nsl5a8tLljDXW4gibDIffW2lI3Z8rfe27fbCzJXAevo1f
6qeQQ6fWWhjeX63DICqXIhO9OWqRMLH8Kvz3mLl1Xke46k1M+fzdLycmePnTyM2f
Bl0kc1Rqq0pm0AS3xej9uWGBtXC8RPtDm0tyNXzKSC+VJ1TMsCgWkCh8qOvzsBpi
722iHAhR6l753kVI/yMkjnXxnSgvSYrGH7ddpfxal2C+x6Vw4kdfcWByBPS3bQPw
rMiPPD9TQtNWh/OkC7fhB7Xzvo8EtddzqoH/cotEq1sCVngUwGWbDhJrs8yq0wPG
9r+sQT9tArYTSG4vjH+hw6zlcAGiuWB34CL8BG1+4SjNK0yzXMtOgTpZQk3Pq6r0
4Y2DRRCMlisCreLPxWmDrdeeRc5k7vF1SMLUoO425sRxkCnKfQqyDNPbZ0YClns5
zUTakCQCSRZsjKhS8U4knd8XtP4GHD5Ac4auwbg1LoFQD8M/jxsU8JpAMg2+vBMC
Y/ZAbfHvrWPIqP598aRJwpsFoLq2wRzzFrYdko3s0BTHzC8nc923YHm/MlTjsgzs
z94EP5/IMZDQNCx2CUbTFw1qtfK/l3oqSIIYEhb9+CQJyAUsUfWnJ1IC+ICzqGCA
JD3Tt36Jiu3FguY4yj4iJSdowjPqbXx0h/cKHZnvVsj4rr91O359+L0+EAIQhyTV
OJOd03T5DvUM8U4I0u6HS/DUvQ+AEKDTuJxW9en4DRjlNavugzUyNUjJBpwSTyTm
XQkmPvK8VHcQmPmSwM9NhIEQyuzNZthxKj6XbvDXSWdhRgYHtKEoN0iCcSn8XZZa
AmWEdi9k19WYo/ziQjUj1wmQzgCiYU6J70eBQRf0qzcjSlp3MdD4kJaIi7J7gIkJ
I4XNZonsNsT+65ldeQXZVKcPqHN1be6a07opgGskXymKhge2/AuNif0Z+I72tecw
Kby/m8j+CbsgPnE69cfn8BbNoQB2uYISYGa4FyTsO6zA+2ast9fo0Z1f0tV+uVa3
GFWbiUBoUpekn5kQUfX1OQGlgZUmWp+PNt4nbRlRdL7XtuYrtsKMRtUL6vWNiyJj
mVsGOLc6ApWE6aCoYs88pm2bobpzfKs0iLB3+iVFnMyOiK/Lcgg/wKwDHf6hsCsU
s8ePU0pJ6he9HqX2xXyemZvNJJeHwhwOae77ymdHZHHeoqG19WjVLJmliyfo/aO/
8DfkX+L0Ic3AWr+JzoQY8f8X4yl/fhHuWB8eGriHrDc/IPVGF1f0W/SlVqRS/88R
Zxr/sMN2bSsL/rgUG9bLg1mVR9pQPoiAtBN/O9kWGQsFPBKqhbAM8EDhYM6nF698
PszPNa3anLYaPR+BRCjiELU7DMhbIm9F9fJPGAWu2yVsw5ppoNO/KNg6aErGQOKO
nnbJeHmgZWdEEraFD2n4DHT+AJflJvetM0lavGQh+kufwXvLDXxtrJI4AmNkCijj
hZoRFAlsYJLL6ufZ8FEboJblEX3ohAhoFNjZRX6qTPPcd3OD1E660SbdwfR0n2C6
Xa5ZfJFC/z0yrgZTgyVoFYLuaU1jhkJNdAfvlx+qbWP7UoWZdcVkG2KwQrTzJ5yR
LRR57uHI1XUQiHSpQ33ueCZuVmYqUa7xupUeLk1jvCZt0Dbjr5tmJJXTmA5exuWs
wh8DdyVrMJ0qKxPEeujlmFb7XKqzPwURUL1fJtlCG8CEzA7/9Q8nfWeAFI4o5alz
lmLvpd2cJauA3be0dAbkp0V2nBcXY5wH3ccPuGkMqyhlADvfGAtWhakeCBVSqcee
0kAC8Fgh4rYbkPCDsiu0ybszLN63Rcv3krhB262VVTria0p8ubt/JNjS6bVLK6W0
POYYy62XmIqoiybPNTxOXlme4swEgIrKCDW06AdMZs7U0eMWYt/tYOtfwd7Uhf2T
A68rtcasJvEfL0KkHIaV0kBdq/84Oqd4kkkFWoTX+hDe9UbXgClLMt3kbxOzdJiQ
3aQSAFqtpzudbQfwMMZlU8W3oQvehYwYuqgtxS4ZDyrSgJpjsarBAQWqCLEudIYd
P080cAaeLvEkU73k9LOauCCT+1PgqJYbZsK3xXOZ2siQq08KVdELHuIVwhDaF28o
r83fHIRPpofjbbZ87JQMDsDUhBRfSGLuHUid0JOXL86Ptvam2MeQrUpoxokmEimP
Pfm/5rtBNIMwFnZUF/ch5HEvbJZeFs204WGfSh4Qap+ypBqvtZjf1w48b5oJovWL
naEvLXK4l5jv6VzoUQR8iPtQsfJpUGr5+R3BgYGWsY2jU91sUKucW2WQOCOMkK4A
mmGcqMHUkkD1O6eu15d/XG7jqu5tge2QoAlLgZR6kq9mywSeHHC8M/d4LRuvRGEh
FAz71Mj+vmvRKMK73oyuTtjOkvEEChq5Knx/icW/I9+6/jcJq4SCVHNmlFLNk1qW
vb55QUGajuiA7R3WJaA9Bx0Ad7UOLXgl34NDxzDN59mJ4OUo5ybRMWoJ2WQk1hv4
3+MT2ktceWxdENHuYOYXqk7hJtwBoNEuyGqUPVuEQMv9Z9V3rHN/jI3raMiDNF5w
ihmNN6QRIhydu7FOY/XgtqFJvq2ftwA5te+nTcBpBvWXgMl6NP4Ec1VIVwo007sq
UljfOIaq5jV3jY8nnFnK7dvVbLrtDIqzNDGJXMbInitsm26TY5WGhK5pSguyqsOL
fX9D3d6fM9rcYo3ON+qMdUVX/eIp1dQoaYuap2edhTfKkFzOlYr5YBYCOzROc6Mo
hJCgBCN09n+bytc2BxoFcv3G4OdbR35ZfJudszd5/ltcsHHCmI/swnRJmfr2nZCE
EemoVnPuntqS4fUm+YQa9WcvoySU9+EUdf6jU2Dqa6iyPJPtwVkK1xg3pyx9D05S
pFOtDA05vgloASpJ9EpfVWw0ORly9utyuqDZfy5T5wJ9LjEpUIV9tbURZABdVMTt
ApmTGiRQBRsLyA3H1anYBiOYgOv/mWH1uU2N0Q6rCBET4j1G6pe6WYk5hWY2Y9iV
fvbapbOihyNKifjX0uNDG89N/InMKKTyTEOuX48z7H7Xs0CMJj1zypnQ0LzrMJqj
wz4PY/2A6dV0Kb7oj24po3S93Yywu/4hIzawri4pwAt/G9aXltxEMqDIWuFX+dZD
xHRZkwg6SObdRcG4zDasr3dsdLmzSP23g5yIhb0ecNa/XAobhvObUaj6ORO4dmIS
pjmSYa5KlvqAaW7iZaW8dGO1gX9SaWbElx6XlFwwuNQ2BaafhJqnAd1eiUy8om0U
mL1v34A0ySX0RvUbNoG149N4R9J1hZRHX8dkxzbrmwS3oA0XrXfOV9SHbJ29E6am
p/bwXHtddDE8ptAf4ve2/BgQKalmogX9yNbiIjHXEfuQNZ9/ztsoISmC3FYn9Vq0
CPfvyYwPaYqm8RXcIbYc95iOS+THrGhO+X3KjaYjK/NPPrji9j0IMyYCZt3q7F0G
QD6mCaEY0aW9OKPLj5ppX4/cnujxWwlsYgpXKJ+W0p66fbDWtzj7KwTSIfm10uN3
t47zTocrswBHvLrJkUIypHoZOo2+qXNY+QP1ShDpJ5EvFLLheXvQpl6cLBU0S9me
Ps1eVlAyNqtDaUI5PQjjGCAJwfrc3DrsHfw432pCm/2bL+kdMRxQKLeapP6zrq59
rVGzkAn7ojGE75bIMl/sIpbPqxdPO0BiEfRdZ9m4HMy8wg5r0TAGYOLErYhrLyPR
SO5I5/DJP7w04Gvj+pYD/Pft09YTBMG1W+id9nybgFC9vLxIKQjsfAEGyCTS+WJm
/4XRTnutc9cu91EpBlIcl3pCKXsP6wD2uJiTndOIXk12dgN/DQDk334wmcNg5E72
VCTqqJ3vjsqjxck3vi4pN1r2rKz3s7ioDWmFjjvRabbd6VhZmj3nTTXkmkNGue7O
kiZjG8pYGHS040kbrxFYLQE7cD6yn6CekvHuRznKq3ZeyzRIIrLJVxNW9X2LP8L+
NqOph1gS6BqW+bHj3Zv04i4q/Nc+5u+wkXbi4kk9en+e5V4yYhNqEPhxPTisU7kI
pl+yoOKgkELgFW7hVaHqXTwPF0B8PnarwUrZaU9ZYlayrUTxcpoSwLSBV1kBvWyY
VdAJwA3QmPA7rxCEfUZXaVMxSQgWTcpmw71z7Wg82koZlrAXfTE0YKx52Us5qdUj
H91mWKR0JwH2c0NUd4HEy3PLsIxz1ne/zKBbKbE6LpZdI9yZb49mmExcNbOi2KzG
1rKHwh3QKstvG9xl/Hpk7WbMgg2g3qa69BEVXcIN+rAqsQ0xvvo5ZpMJgu64DRXJ
EB+IUdVaV0xVhgjddIJfZMrbblAjf89HeBkGtTMKyUNnyxJueN6YjNc604WoijkO
3Pg6Tn05iDrrUzCR9GhBmqsTqrBT1JfJUt5FzdIRNjwMsJdNN6gQv8rChzlXsTEF
/1rqaCy/n/qYMKqadYJ31xjMyVcVDS+Y55uZ9ITqbkzm9V0016wd4DPtKOt/cCPC
12IYbLbWhkp3WK1L2ypKZ5vLTJdqinWV6NmK+9QeY2lIzYAEQgkgT98V0PHN9kAi
ObL8F3KSPeBKZbKFCtrsctJkmIPUBHAR/2VvCCcbJ0+u5zN55xH/lDvvZxssvNSt
cAPHwl5/2UpUTeHdnLtB+ns74BtJ4zXCir3i9qGKTxKCA/PTgN/Ux54Rk4mnVAzX
YjbKedQQZt+GZhZ7Dn1aMMG6t/mPwi6GtaEl2Ri+DV31zhbo1rxT5qESEJO7Rs2n
FYDJa5M3PjICwcQQ7cIo2bluB4yUhhk8HZSx3BObMKmNGynhIaAf/11Y5W7/It60
Zc6fv7pVyxE71Pp7jgTYBIQe5CrVTxywqB5Q4xqCFi6x93QWsNm6jqM+XNFY++oh
9XV2fSWWVFtmJYD4YIMkqG+SRBJQcC+J/1XIe69w6xifrXRIIDJpMi1Dh51Aewg2
7Avm0bYqm6Bv1iF7tW/+gtPOuGagDXHCvcwkZ5jLyL783+Uyb++EK8v2Wc18KsY4
bPHTpV2JFL8HwjzPst/+9vafv8fSfN8U8NW0ZS36o0yF1enxcMO9NnAdUCnSMCX/
bBVlGvdUdRf5/YCooQd57rUL5rKD1N3Ped/jPhjMlKS4BCIcLRPUJnz3wPXzv1ic
46014OOWcIZ8jZ8ljfsrXJu7oNIfC5l9oZ+BEYRciSO0KNY8I1bAi0q/WGLD/GA6
LXq7tabZdot3X3Tem2yY//WwVuCyB2slJ6RCl2y5SpIJB2+LXcQRrepNRF1zRf3g
SGvcZ9fV7FA4umun/PO3F2cfvPKy9AunHWLC5ustbejv8PZE/YxKUirlVJN+UOtL
tVJQVfL9JvVsIPJP5VKSDi8fvmcaildUHjBwN8VqbQpWkKKaivjGEiueF68xvhIs
ZvrOMFYR7lZ+qsyI1dn/Tiy/Df14fuLPpQLcoeDqoFznrdMQWGwvhpoJrlBc6XZ2
cfXdHmJdrZ5mGNgrNgTffVytOZ3HQtvMWLHX30AV9Ha7UTzm2J3Kkd9fA/MHg+PX
wk6BOx8b1m9KOWxwmiEsyYEW7AAYtQRpGEHEqHlyU0K4BZFaL+wbFI5qNDZlau8H
w0bJ4IZ6UlweFr0LgETwOQlOtzcSFlZlQP6fmmss75iAuht8jtUVKd0JEd3Mc9NB
l8PHgizBph7Ag1r6tJppk28VhizEyNNhHIFeBZ5DfCv9Tw79INBkDrIX+dFjkS9X
3BccLGmn6Yg++nCisesbx5zyU9O4Cyo1TuRlGo5I3qyg7SBA/QeCnMqCNXA6lLgp
DangxoUn9Z7EAldAfpeHW92vXuGPIXKy7O0plzFZMzhfPuBHWmHz3JOroN5OBwyh
lNuycYIrtEyPX7m6fifVYh5YNN+nSLU8eJjlbqC47JOlFaeJR4A4SEtLKeo350if
OaoqD7BQWE3T/o+rz/Fo5swkZMFMMOQ1zGdCWwYG9GWEQGCTndCJd1jAvHk1ABq5
3mYuZr8ShsKfs90dl5se4ktM5c2fIVHBW030Ei/njWLQLgtUhup6d82ksrQHP7tF
UXV3hlG9+A/qu71+2rjQO71eaKVOdOovrFrTf4Snjyjl3zfvyxuo6vJ+DCv26Wu2
dfTGrYAXgik4BaUDWKT1Q6AZAiiDAlKpd6CoTsEn6mOjPvHTcmOrMKxHg4mlUWAZ
cwpSKd8/fU/afLLNKF7RRsXmhsc+fvLkPQ/14TTSXbw0psOfU8XJb1uy7wzG27jt
ReDP1XGpCVBJHOHvvmXy16295BMoP1hR8g6z+3pK9w83txmlHOjBXQN/vtZqPqru
iNhEWZPvoLvwzl974juvHg7Pk3lgcAx0BTpVT8db70bhoOwh0I5tw8h/hV3KiahF
9Z4ZZY1gUwZGaWY9wsqkc1dmnakYQpdW/6maVMDG6ejyBEBB67/9jHIffgVNzCY6
Wr4NZZHe3Go6N8wwZjLy+yiMXX8783E2z6S6PcShB2gVJU5WBMB9z17Lqf5i4pCn
nkgKJxuQO38ZmtHgBLndh+FHkx1CDY51bmmPpyJzTREXT3M6Xj4SH+5FNcs34Nuh
0wIbsfgHtVgymD/Bss/FF9JNIU3DDHF+p/fY28nd4slljc2zffNOwQB0nEHq9nJL
TUGVqYrb8yLWpdZMoTEduy81TKZgUJp23D76oLaFKhugITb+R9YLK0qNB2NQPnqa
jn1jTg6UPB4fx8aSNRPrKe0CkLls1aHAyv3PKvarYEpOMg6Cy3ybohBj+OIQkQa8
+AlPnQo34R9ETL1MFekM15nXr9oMJt/EXtKsXpSspILavxweL/ZYXq0tGubsASY6
PUQNzeG/tOR6li/5G0gNJ6GpUBHdvGSKsxoiVf2LHFuStGzdsLzZw7bW+/mI33Bv
ZalLIgl39NL69ucgn9x70fQsWP+iviqxM7Ko/so+oMxfdkEDQutG4h+olID922H3
Tp+1ol/AOiliLYx/57XqYn7yITy/qka28t1zenhMuOCg2qfgcva1ofy6CAmlv9gq
hqNmfLB0qXaeatOy3k1B8Zrly/ybAcQiYN/0P+xPnMzN2zhDmK1aX16c3fi594Vb
m2P1c6uJPP0/3Gr6mfgxiz2hNh6XK2FWY4efeJq/O9NUHPXnbYqN+lQOF9tznp4H
TGLgGZONKSJKrjeK7+SZzFeg76RjT++JdO1OqmSML3aKrLPwWYmD03zmSR8g1ZqY
qg7AzwIDU/81mEJCDBUgp4AUeotONXycfLxHPwIdiIXTK4QwhlE+pxmZ2oNKRKZ2
/j2qj61xTG42V0tkwUnPTs9IuCltky9B0BrQ3+26ckwUXBBhQvIeUMIvanfvxS+Y
vB2veStaM1vC8tBqaoKQBybtawvPg+JEgXoNyD+UKOaxprjSR7aS4UMZdX5Spux1
W8njk75CPRrRxyt9XtD2mVH/T5AT/ttL5XnA6vpmpUzhWjZBgYvsC2aG3Edya0sM
56JJYdjmXK6ViHmMx+J3A7D1tr5zlUotE7YW+NbO6eTGesfaTivJbPHiXXecPOAY
/5y9YkVHyb0qY5uAzbftU9eNqlp7mq0hqKgnIwLtVxB3B9FGVOH6xEBEyBs0c+oO
9T/zU22U+qUVdQ5mNczl7PPegtSo4E1bwURuFPPpOP8jm1sOB5e54mM9HW5ukVSM
QGImz1pHjlnLOKmItST0M8/z/Frb0MYTbAfUb6eEIT3nXuXv7tRqWaSz9WizMm4d
CxBFFEpCSxDrczneJTODgxsHvURh3g7HqIVpB6c/SKdMHDFd1J5Efsj82aQSLE1v
sumvXrTjjS0q1ixcZOpwz0Kb0Lr0IWUPdWE3hN76+gvARlK8Mb0fYGwJ4uRtabSd
jcMDhxwXyj4oMJIg0VeG2s/pboCRsFZditTrULlGQiBEvHs+X9sKpsKA1AqGSXtr
4l4p1yP/qKx65In2Xc9LU2avU4C3elQKN7FkhH5zBa++SXPpnycwA5M8VJBIpdTS
zmvSAh+woPZ1JPgRCDRcgHYoXgSraRGOA3CTgNVJb0vR5FCyGkl8wevZlF27w1z8
HgzbGTrhovI+xhg1dCUQOesCtVhG9RUPXgvjXfU5FtVKFCmP37uKrSXSfEFJfGAG
K+zdwVd+xxnELuxJAsK2WMGD1fWlT+Xk7U1mI1mGz8zToHdpmBHoLJWYW5aZN1S5
xcOzi8RqJqg2KgTIQzttcSVws994IY31HgMkV64+jEb44vSpdnPqxQ1pf2Wba54e
nukMX5FSFnTTUYvMj5I5FVsQoamtdjzz3ZvY54DbesgiGtNLkHDC0burHjyRY3p4
BxuZ7CCrzCAVwhysp6WjjE1Li8gQZX47fh7wNEi63/CEivvYaHRXrRLj3GvAeIqh
hTyhwKLU3iLz7tuUevnW4bMQl8ZScSFUHeQjrI0Oeoa7M33JcRZF96nWgWfxMLtX
cZ9UGU47HXjeYtVU7L2ZY2ZCL3w4ccYkLCfTNRJkkVqusR3mVvltiSm9IP+8AHgK
IxH/meYaM8Pw63wa/IsTSFqhsevpFn51mehykfOxm7oQZhwjLWH2GfpUqqbQf5so
/5e5QU58ubJFQy7Yub0J7CFOmciFTeNF/kahJugb3SRf0kQjduYJ4sO1kpsao7pJ
2W0l28jOF3k0GrCNllWrRfax/PiwRq/VSieu6nnJMONtddfS05jMuumKM0fzyMOn
kxjhon8lX/LEz7KcfngK6wmEhys3pHBaqRwuq08LqpM5tNZvaXSqIzKuDOcNSOP3
lCYmRNJ0RNe4WrnRlGrrSPxeA37xbYuxqFLwNAeQ9BOq2Fpj1eegNkbbnfBfCv4x
o8qUSdmGmh4LnFWu9jwHcTGnAKUwpT2CTIx5E9SWrffm90qulcOai5VxhriTM49m
Nmftg/CSGbZtIWMKIxFNAf9EnVgyWtfpILcWFIBEnhOHfx+Pkjx+viWjsTjK+4gD
1mog7UaN3AovKYVTl78zoE+LARpsuweriQzupl5T64QeJuVy7fer6GnT7htXpv8v
AZlLLOu2hphl6OjpBf5pH40ZEfHrg5EaHUYHAtGhAXMjhA+Nwvt6LQSXEUiSG1QP
84MAkYAcZVygZMEJBusmsblQsmmyZE1mMljg3FjQucDUk/AyLNBty2fkdQMbjlg8
r8DUw84Ticx/VFEVkFMFxoz8o4yH/wbYtL+JX2veLM6LQSnnCtpxZWH1HFz2iMrw
RATBOrNkzarFKv0i1k1OPn3BRBwcttAuZS9u52W3foFt3z2/QqYd8TzQ1TIDfSjq
c3RPmJQQl7ELt6lRHMAig+6j017dNdUUP1Trof3M+o6+zVViip57bwJG9CFesw6Q
GUUxF1FrV3/H0jJSm4xxyszkcVdgYhTqFou+XAzi3vKzez/oQxBWeNxiAZsQ2X6s
JokNPeZhu1PK/x0HOWpHF2SlmRn4Xn3HCLmDQqbHz0vN2AqyGoKnCxEAlOr2eSc3
sCpJtk9J6ks6x5XHzBHqOqMVjZvw0UndHymAtah0coHsJvkpg4nmVWyY3eCN0bjY
OhPJTGORnWWHvn1pcXwIDkpOvgQy9sozOeQFnEdvF/Kfrjc94LBiyhlet2bNc9gY
xfcsw5z5UgHq9BLcN/mqj0bJxy7xQKY0t2VEIkWXmD3QTcnRZ9Pn3k4JXkj+5kmQ
iwdQBPovlyTCOzQV1vEviW6yOZYB1OGzUezUT902Bst/YcxOkV89tzHKC+Z5hDZG
Qb5xsyhzu0nbEUjHMQLC0C+uOcz126NJDSSr3qVo1P+aBHcLVuBH3sMN/VdK+/MN
49fmgEmBhEcQfFD+X15E3bpnILLs0qJE4Z98Y92cWhNbsDPt/cLjznQQiAWa65la
U3WK7bYF5U6HVft5z3Dzn2EgeGWsIQFXMJBs2AZrbd78dxcOGDwoZnxsGGtGAU5D
6J7maObFZWTLsOTjpSS0uEcaHdAUuUxu5HbVtOw6jdFhzt7mR7Dpn+p0gvkjLLl2
BBtTDKiVsvcaZ7Lf/ee3Zr4rTCJCpQiwTzvquQXzfVEkL3dsVOi6EKBwY94OHkWJ
sfLlKNcKVNvJvKneXA94NZY53covP4DwBnhD9chSuNTxfB5HcfeLhIexoCldrVs3
DCkRzERoookfrvuga+0bK+0SfCHl0YpJg/uWWmclvt24JqhOfy4ivZTHot5dQ7qY
UODhG7w+x/LwouFdzwodgoSatck6SAzZMX0vpbNdyGYHk/OAtvK646tCe6IbRKnU
YJBsU0vsHrnTilDes46wVLiVdLBQPE7r0MOhMFsuw+UYTv2Y3IUWXj4S2omOocDK
XpLSTsDfXmsS1R7zrpRoo5EqrHOUd7GdINvDD98BaHRp2PMhZhwoo8UTgSGDoiFb
A1ZXaTZI9GF3oLafZ+xkxqpiPV89uyXSrJGsSBVzgzF0nkBKqlvhG7xnffsoadcg
fufQkAb6EK/uOOmN9PyVuWMl8C36wpm2dtnL2E2WwTl+tT4SMQdJqNUNGRYQerQT
8gp9sNkrwOeVcZIz1QhIMPejMuJbhSCp3p7TQpIWcFns4DRdwR6nXTwpIpiqC5AL
vyKHxb5a3cHxbz9MSEVp9eSMkLsLGUWBNepRgdwJzuRt/Qe5v07p1x/1Cmz28pMz
1g//d3lK5Ll/WF36CLGXv3yORPwrrLceXxaxsSXHQcdYeZsYytTRYFiOJy1U9P5M
GRwl5FPZEe0hLxD5EMxhL+oYqPMPq7UfP/OsuxKXdPdm9O2L7EYexnzscGr/+iQs
tNdTJNZGE5O8y5I+/tue+rs0P6JqQiQDVYDkyFgSkZ5QTkIuxFuN7pc7K7lI7sYw
rguX6ifzOXAfg3S13HLWfF22i8XdDTxtqe82n9Vf67Nut3SP+V8a8fCF/i11vFNK
2irOEItIjsj8N8Z24K8C/R0fTAXERWMzLFqum034lVpAnoLCHlPh066AutPyu5Qo
xPZloH3i7cGgs81LJUdvv+ksB2bgMshbLb3gSL827QiZrMdYURvPU6sazoKmM6ok
pGADdIkxgeZPWC8JwX048T7sOEqOaqxQBZNqv3rGykGkYt4uNPdABrfheQPVn8jH
hLpITOZc9ccPucEWA8e2Dr0yiSo2fMyobCNltRv+EQFl6h6Scw+KAWdmMTaQ2Hbc
QOwhdftV8bQQ3pNYi83uFGZsWJDhA1RMIxwDNfmxBrFR/ZsmZc7L8tTEcUWUa23V
KKoIlHEpyZ4lDbVR9nu2kviOqwiP6vFJL4nzX3LuyeYkY9n2PakGiZoCdg8e2QIu
3bxYktn+TuJJDP231sqSNASgDOhdX3Z48TORXR0oakbHoCgI/wi/JPL+4RLTlyc6
uGOgRK9A8pp0qasvZ3XJfCXhgr1VekIaDW3hmDmFQg/aKZNiBKdT1oSvmPPvjBG4
Jwjr5++EkOsSk5ArghM7R5cb8KCyO+KHzCVgwLkP/GvikoRav2pVSORxiG/Vunc0
gLSkdm28q/XMkfYtJHPotR62r74vPis2Z0f0wkUyMGy2xVbR8bQJb59vYkIU0nD8
otMexoEgD8jlObd7s/hx3POUIlx/ZTxDVPObNl/DsJx3SVrh3Eygn+0eG5+zy+nD
4lSijxM2jt42pd/sFenXfe06yLEwhn3B0nSdp6yVhSc5lJhnuaKnmOsWkZQt7z6N
bzp5hmabxYdiulce8+0lWb6thoHNcq91WwTjilqB13fG5cKCrrbpPdwnPilOIcE+
QTUQE9iGp6G/MW8IuSz+RArY7tEgDveMZWkptb3IgBAriFJwTs0Yh6YCvCxDSMGd
SQNWREQSsF6oRzgPvNWE4Z3wulrv6BgEhZw8vyJOYkGdqUrMTR8s0017g2y92kfy
hK9fXgyp8pFMdot/ggeIN0bFukgmI5Qze8cw40ntXSKuFTQLpTc4oAsKgetjcVDn
nL96xP5Dely0dZ4LMpOsYTTTm+ZWgvHo9nhU9LraI9B1M29K1QH3IWndF0wygROB
GhtQxNLvQ8X6r8Cm3TTb7VOx8BbaaKKzSlKJHwirIjCU+4nX7OblGqqiRwKjxeWz
PdZcTxgkyDa2t54gQmmepyA4bDRgckNemaVt5fcwjZkdc0tkXHS2Q6spf975PgkB
JpZUo0lqaVG9PsAaTX6yoTzVAE5pfBv/gee8yWxPK59uIb3D+ZWu15xzofDhu3Q7
GIbTOth+XGTOY64IQfiY7cZrJQbS6zdcGyHxYE9t+jiRLxYLK76nN7wH+mfoinUv
BCU4eDSAgyMn2PIAYk2aWkzTqwmTG8pNGIp37IfAIGO48zD/cG+XDF5ZZHWS81GH
HLTsSigCCfiN9Rncd1vd0/5i4VyybyiJQlTTF1BvFSDoFWe4FoWJVuoVNv3EyDAD
SWF6Km7+9ExC0ft/HmYxHM2F0x3L2mqG/sjCl58fS9/fIuWKYDndZySDudAl99Ns
7aS+p0rkW2GmfYotCKrLI548o0asBlMJWScMqkqEjApsnwXZ845A3Sm9BAp15wrg
OmUZIuipa7Dkjqxj/OVkxQLrhkZs/jvQ9OE0ijIMSM3kNfTV8XfI2+Vtr9dcsKVB
TA0mNWLYioaHXaRsTZcMJ+1p2TKz5rL4RSKOdQ9sxHvY9bc9WXr/4Fk+d0WrscuB
PF+s1oFFyGnmhrIAOVhy5RLD9Ac4C93X18YI9XCOsD0Ko4v6hwpMefgvznExwn/O
s91Heipuu91pc6QhcoEDkQplo5HR3Y8wAnviiE2/+xS5LdsdlLmuXPqTtSVlnQ5l
oP09k9xbZc+bqSZmJYAfG2hp3g+2D/r+qftdhI45fTllSR68r1bSzZP+cPpbQVet
rJh8bEkhkrdlUYdQRF0v50HhmX1+iEQDh54BkgnCUfnYBwonu3Zz6U5yRHPEOV1m
9kNoZk7PhDIEe07ENr/FBOZKIgyvj90VS9jXx02OpMciw73QU2IXVN1RgfQfPrvL
YdJPA3fIJO8xZR8x86m5OSenSUSZZ+qM6bV3rFg4wrTna/ykaUvfn4cl01iZfnfF
SNQiT4fYv9sDrK/7MFeDGoymUG537GIjnSBh8aooGx/Hm78fUc+sh8JwfUZF80nF
fhynrNRiesBqiN3bmBF0w9tb/i7V4wOaZCwaVuEaJ0Pt3cRehjs2r4xRYe3NR96S
CILkfHXHY+I9fkK30Ov4Q1WwVW13nIjAzMlPbaaIGox4hz7YTWfDFJMhVM6eXqVy
SyyOMpGojUPK5PuRGz8O/w7XUovldZYCSaQ+D7QH94svaW/8K1qN8iatn3R4Qnfn
BgkccYff4VLQCHZByQ8tE1R3LwebMNg2MsJz7uVLgfPQ8nj79ZLcDwcSWtiZtzq7
eX1kf8rChB5BxgwCY4t4aQ+u8LMXueI47TJc3Pkb0HHjC/DpgA6BPDM8NF0ci9XI
bXlm1+lAQTtkyd5dOdD8IczxWO2MrFCkaMBNlky68IanrDi2J6Yq35zHDhM9Bx/H
iJJBZyDo1mocs6YHfJ6os8E8sCSK/FwpWyhL/ECVYj867t6KtD1gEtP+ElFDpb3U
2pmZHp1/2AIrw3ldquejjb9wTAM3USQzCdPmC/UBlj7253CpnZINjPp8Mrso3rTK
IOz6W00LSnF954lRUXREoB91NE6eJoNMv0zDmHwPZxmMFSKjqMllW1Xpn0B5Ijkz
o9p++CeZGGMWqOW5PDH4NljpeQlxx6P5phl0WqUV+yJZsWt+cwkXWjTN2ibGCRJX
IFCTytmnfPzCR3x9BL2rzhfQ12sXvLAig65hFAJgswpbFjiBlmN42NW9Hcsk2lxo
YL0QjsDiJ/8pyWwbqo2a9n8/tnEy71p8gCkO0+6sDFneJ1NcWzzzOkuecUJJF0Fd
7DNe3AGkUZ7ZK5pRZZruDlZfCR615ToolKba+uBwQec1BeVml/VxtaZ+uVAAl22/
oVK4Yxs+Rc3sVJyJDJvi/Kf4Lg+G3+X0IHVAA+6x6USuQq1JMFhQ+GbQxJfAQfxJ
Vio131X6y5gGKA0a3oEAt5Oz24gRUtaYsDB7TncZFC+O9FbY6aOF7ZqsfTdg6jaz
BLZXbNuETrKfNogrYa0DYa+JThz2bKLXVY13guCAUXQsTRIKFwtjS3G4bzWcNIt+
DzpR/P8MiU3rf6HVYVQW8syROTL2shNtR2UdmCPsDGhgkI7yy4mDqv/R+GP3s39b
8D0IyT1FjpX5fl66UDbol5wzo1oNEpd/CM16KJ6uda/W51X1qZircVyTFQh4ehCF
W57fPGFHxWc5adtgKGxTy1OIRkkBJ19G4H4qNvOC8XzFc5m4KKQGXPM+xSX6cANR
9MNdBWGevk1tXRPKo1skEqcYGl7Lfs1QxA/8fNXimErDWFAJI+RT6C6G7q3j+xY2
93l7/I1vx2gceEY5xJWoogLw/9zhnj0rnFfpbZ2oc26EcgurjKj4uPcrkteVgHun
GIrWUiT4EzauTsvwKCGOUYfEsQydfDQWsxGHfKssHoh5VoLSOfZCnoJknVzlJR6X
Xjmu+V2RgM7+vbRenOH2MFrLzsL2hEGkG+DcuEUu6Sy1RqftypF1coCrYJz1uPZm
Q3wC32yIOsrcE0qwexW2RPcV/LJCcvWznapifokkDYhU8uOZ0HQzLzYphDyhEX4A
fJ4BaZbON4mFF1bakZ5gAdc8BeVTYC8zOptuntqNdK7p/G5l6828g/JCLBsw7YBI
Ic1W9xqd/1mLTpzcN4Pk9YGGVvXlhZqhCAjRhXVPR0px8++N4ojgZN865yTkw7QZ
/LuuRpiSTBYsgPuw90uxji1wuwbWncUsg2cKQQqc841Oh9erpcuXv8CP3m1vk8r/
mZlxSx6RhAl0QwGAn5dp5BE7HzN/Tu2DTOyLv63R8y1JHIh9I4IGW0HbYqpTBvwF
QvLvMhJFxIJySg4/N3qhdcgOUt3rypeyKKYgVdX9wk06NBfgVtTq3bAjRJC8mh2c
CQVLFVit2tQMFG/ThrQEB/lPoEcaTbRp8+QTyOB6do2BeuleVtAfI+FYD6256l90
6UR/NmsPMBXQm1tR8jebHAlneeS57uU5+KgAxJ+0GEoZ1WMghwP6pdaVxfDiembF
GpXzn7QOe9u2r1aWojTmNUuKOFpVG/MoptpdWlp0dPLpc48GS5RJH2J1u9JFjQNM
/7w+RDxptVD9js6tdnVlNzZgTMeGoAcSvX8bEU7L4y5QaQVnHh5ErSFnEW8wM/+G
VHziVoDsXEgzGg9fOiuVLLjB71OGOaiAFuBAK5ZQ2316pHffAAWrmmpgt1/VDrYh
vGbRcqzGs79tkTnVsXKomgX9KnTJy7CtN3Ufv9F5ZRUcaqGqISzjOYVZc25yyHzo
rPWnaM8OkNiT3VPZEHGCi5Da60hBY6HXjLBU804fZmGbE3ls2JVFB3OeewnUzUi5
4eJsqbnvjNf0NQEe9C67H3bmvZyaxx9HtVfPxAIcThY/HXD7NOWiZE+O+6uV1iS+
gKzYskovfG1G9RsAI6bER5SF0RIksJvYsk+iqMZH3oBi1vR0TYeBPSQJ+Vr95rwv
RCAx/d1fiBXtRgZsopf3mdLCrTllohuML/Bbs+OMivpr2OegkU1WqYBybES354E7
2HAkRidxUwxIuDTUoDEug06lOdkl03RcY5VXDcbT6hFFi+Yx5b3XWyCDEHz+1KBD
rpY4Z/qnjHA8Uxrwtxwu0u1z2cdNgGrmZAHTY6Okye4z76NYyqhP2LlpuYZp5ybT
g9ubEkSUpS2r712CGPPF45ngffP9kGsN8RkK1AGfn/vVcCHh7tRwMgjHaMmwhvJy
h2twKRqqqnGAWKIwTtRpQLdUwUQGXV39KK1xFmINHbcXEbYloUg6zY0dq67nxbRA
Zvyg66ZH24bFUcVxaCglDfYKrFtTo07LLmxEJ5swKCJOrUrgQQ+EYcVBjlF7OWDp
quXfd1O2dGazjEgBW1fXn0pS26hWV3/L9eaLEYMgjC3Xs1XE2zntIo4A0CJjrmqB
qQzL+RhOZZqjhP4bvoOPPnmP1CQ0t2dognG6VmtxU9LMVczo3lFWmhDJCFzCfmuZ
DsAC7iAMXa+nDImGMCP9joYWBVo5B+N8TWrvZsOUoRhLrtDCeYeZDCbpRENKe3qF
Q/RLcWZ9t19wvuAL9MHaNYAOSDVbz/6j8JYvhPLafZPA8UjDdtHIJblt2Ej6grl4
7aTqe5GRM85k59yUIb6AvGD7eM8ueFWs/eVwUdcxgm8DGXx3Op1jiPOmQOBf9x1H
Y0Irl9/30NoMRHcHU/i30g3KAHmCt3he64ArmkOhGX2ahJRmFGYWuxfRV/POok35
CmXZJMpAN6ntIAjAMjGRiuMJhiJ1xPg3dnpw/w3RNxshbfpRMdiginKno2rUWrlg
e96P5Wxy/FlHk0SZnlnZ6KTf80Ky0xU6soOk/eFIlsr6dCatYKegMD5khHWlsz1/
hSKRg/sGsmzeajbQx6JkQuRIS7lrrMy4NQfH43RXC9HDl7qtwxHcEIx57aRmDMFD
KmDAv4N4Y+wReAZ6JRZf5vam7jQxxK5UpTSP7awAfgzPXzpAQOp3N6kWdJ+7qgjM
U9Vdv7kFFndSk/NW8hdenwMFFeiXzVqwNa2sex6hJ2yvTjPMtZqyCG3+Q1gPm3A5
r9BVx9h3xO0lsplnmAa7I5k0z/0+8aIJBsFo8CJy5RMY+N3p2/dxHeaTHdxTcsa+
ypqEtMp0DUzC6KhG3ivlbkx04Ymvq7BL67KMrHo2tzGMm7rVfE5BzXohM+2hBj0R
2vmaU+YOsM9KVWs+jbg0EhxMYsiBaiNMIs7iburt2diNYPFBX9PnkPutjNnXu/4V
1TGgw9PipuAQoqID3Zl9QjiS9iopmDkvmFjNAlkcpOdQ8YWT24QDBd5su3nSdqg5
uJ8wkfSv2Vfswd0GzPppB9p+iXVtGJH68iDG41yLGF3Dvexs2QmspNFHBpKfTgki
ZfI0o0c3BvLIzff/QP5yi46WiZyOQQQOnE/+c8ll4bv7/exp/ecylES9am4hsKxl
e72ACytzn5jfVOw8Ob1xKU0Ip0fKYtKJTsim9dVIvOpIAgQmW7nimFO9g5doy8hc
Vi+sWVSpLxRbNasfqpAC3mMk6fPj6/C1OsBjQi6z+BLo1oPtaDRLF6gEU0AIORFj
5u2KAr1btc06XfOOQNg6lrePAueWy8LcCEGbZ7VJjiR1XWKbf86A6D9UaUcARSmV
xq07GTFL4P+hqidCAQbZZJ05Wt74RYvi73wdsiCrdwdI+VwQz9RHKKVMOInzr9Vs
Zinr8YP6mZlN1gOdKeEXRnY3neTopYzSHM2kubcx1UV8s2qCbAFiOzKRVJrrW017
bBq/GBlHFpu7OKoY4P87sDPPHW9SIhb8w+prB+txn6V5yLKTqYlWKHheK7ed6f4w
zL5NsK/1Y85VB5muAXCCwfccG+UnbHnu/rBN+WCgsbvIKjic+jKf3KyMYDgq5qk3
WMGMpSaYyYy62PuwDPDCrrE4ghvxHm27GzZQflmDSj4/Vbz6+PIVKbMcx6erP9OL
082qmuDsC5aa5M9+nVptZEd3WRgn8hu2gfUdllMnfpw2jRNBzwZ5yLewmF2nT1hX
AH6ZByi2I0W3ktr28Oi2VfJGe5r/2KJK7JdhjGrL7K+2l4jBaf9S6/edhL77Oute
l4zidIzcgQgtJnI0spZPRKHIoFktGKkPcquibR8lT3sZLRhknojyXb8BdCDcLdV/
w3w8mPcnP3l15Ao7Om8nP0RpBZCt1cPcYW0L0iHG+PvR/7UNwDkuyA/N34svFrm+
9zIuPXhxwgMJ0SosOHqXdFbTQspOvmO4ByzdU/3Hcw8XMpn3qfuVqKO8k4fqfc8N
HKe7basCH/ke8rwI1xMfBqCqpaQJ5jarQxxXUuQxYQNCav1UF3txu1QiT8yRLTe+
OF1M+05b7fWM1H0mNQXFh4gIFcAjV1pFHW1WMYrj7k1dnAItydrqa7xPC6mceGSZ
0kPC8Vm4wv45LWx/ImhalldmP6sUvazxPz18eNUC2IuBVC8wvw8YnKAUHHh648EL
tkhGxi0iU9R4wUNetJdcf+jAPgEKyC4/fnr6dWDRARfza7NHCBpNEjKwL1h5b52n
qRZBKoN7fR+LaO/2TQ0sBbi4hWK9aIYgYVKBsicSqGZ/6Q7IfZM2uTKjcyaQTHae
6QHDr3TY3wQQOt8QPRPjPFeD3AssEUP0yFlnozd7XDEYRYTJPEMqKM4/4zjsBIjw
5EFHwZxWBlGadj6Z3KdskQhSFHbN7yYgr0wBeGLuYIX4o9j+iiySnCn1UxL/d4n9
SiRo18NMH/3glITyI6W6jYiMTd3x7gGzmeHh7+r3iLbAf58IAe7iHxLxxpM4eynL
W161Ff7rHQ2kXe1AyFWldUMWjXoU1oKLPwV8WEERuv8sDh25YBclQhZ+Dr+t3JTG
vurWNb5j2EiQYzr0d3BW4KW9T2o6pABBqQL4UZHEIQGyTYdWPRi+LrMzLR9ZDLcz
zeAmrOvqytYpgkDhHDr1yvgleLRaZdSynZcL+/9Qleh1Mu9IeXvt088e5VC3xMbP
jF9uo/HXEXbzrbur8NK3lfJ1s044p7AuxPcTd0f5jR+OyaDKAzsZNw/Rc9MqLoUE
7TxNFgyoUOzZoXvHNJD9XJ6XtHnDBWLjeLieQWUm2oz/QLW6GnB6pm6/fIqwc4QE
Gwq7VRI/Q0llk+vDy/pp4u+eRrHJGrh1xY3ki7flhMsO4Da65IrOlRKXQf/s2Ao8
isBwTLYlEnmaZdfOvHY+hydU4qYFpbX3CuxQDyerFQr0mqZMVqM9MMIscxTXBwqu
vOlIAcAPzeoahTgf9G3P7mmAEab+G5TsSL0UU6kroKBMkylUKyRLPTSkZ0vt0UUJ
XhRyDy++6dEhvyN1O+zEeWUtMaRrquLh0rWDrCgLZ7r/5tDZiCEIqguGhPOoICWJ
0W1WaDWJ45AcfD6kOYjElklOjgeh4cm4nwPxfZgVo55BxXN+xc3i+J94y/wAuU86
7MIbJfk+jNdJkC+UQNUEr7LTCVq9UWFNw+nC+4nFE/IiNcmEdMrE+O+EYSTdUFE/
d59kJpBY8hBlvOwG4y6RJ3zX53dGp5iDTX/8XGsrh2LlHjzdfVr0pHYvVwiwILHs
/TNXZp4Fm4vBILukeb1vwc0Zr9mDACzGoXRBtLFsrmBDuKRhYiRtFXFXqzwAGpA+
sVsI9ByQmSE/edJmNPboePg0yWY80+gB1Es4xbRvnOxAck+z4xkhNLeFDr8Km5VN
AmRC2Pk6jfSyJSrdImms3SdoxXrsK97MUpj3GzybJpiOW4csx/BDiPE8zKo9IHfL
6fBFsuK9KZRkPGzR7EhIoQlGLqfz0B3PXw2ZMspSopETrt3IL+zE7n2FApfH3prY
wHhMoZw5m8/u1VGZUJGv9ONOVbunTJOZ5GpqzzW3BGPfWrlDVwhXFz6DldB4Mx+q
m6rO7eeivMaZgrSv+z3Q8nyBXo/a4hwIvLgtAeQQucqh9wUIP9lik56G9DhKO05U
WkXzg8lSnVMIQ/A1k1gxdM9+jJudfjRgRUeMA9ak8gW/hpdzl0ekttnda2Ck8bOm
5Er/yQDocECgFKLZ6RMZ4NrH/lRjFP+zpnpjmkPsIzvq0xNA28kAScZwECUOAB33
5IPoeTk1TNTmFDf+LVOELnwfv4M9vyXox/RHeB6dp5UA4xe3g3ayMcyHL/cEOPw7
wGoKGlMm2jIykewfOolHXp8xUFDYyS05oZYUGPJBRzJSoEf67GLV1BaFdlxQHL8v
MYBGdsHGwN/X975VkEEqtqhU4qvJBuUznd6O12Ru/WfTfUODWzLCcrOhd/DGRo/3
7/4aGPTv4J1qZbZbOyqSXMj8W0sduD+ksrnwwngfu6dlNmSljcidstbuIX0mAV0H
Do/mKe/Hk/ulbbSr+wB9qYar7Y89uji+osor7mK4Pe8N4awfPS5/cbH4Tx1Ehnd+
JBMa/TwEv3TFSbdqufpkx/ppgqO6nSbZQfvKZFw+hicbF+migidmNp5xYX8J8WXX
hG0p0ciqHE+VgV+WEUc5ObQ9piICYfkMHZDcgVi9KfumXRcmnNygMHLaB/Z0WcAe
nq4QCj6lgPIdEUJcq+nsSMwpXNl9lVWHGakleBUyRIFAEggDSKylCFvDRRC5mifc
MxI4rjfRjmyyCERUP2iP5KmcOBkVIHTIVJr+mzjdYUj8VwW0P+9ZUnp4ZcSSz7av
iZN3sif2bEwjZFL7ZLBwuqNnIOrRLDqphzEutTKXClvcFFtErL9nfnBFRnRrud6L
/t9eojxf9uKl5cq0giNQucsHmCwRbw1lLo6yuZcN5ucNZbec9aPpIF5aR22OJFA4
JxgvucK2VdLSJU3u6jrSjROJr1UdwwuAUNxOOeJBXpWg5Ahyes+UsvgnEcoODpBl
ZuJv1HKBIcL4Q+SgheaQXZ74DJqR3rCPGLkWApvv3SEXuX0w3aN+U7IZqgpvXtuC
LSpnB8TTSZI83IQ1+Vvcj9AykU7rW1fmZau87E6MISCsNx8dZiJk1E71n5rz6pXa
IkBuHboNuXVnE/759y0LglSfbiqgr1ZxoIw1ms3GrcV6G0F85wUObi1sNJLa7c0v
bpba7GHA4u5Jvf46BCM8amI/dSclTq1oGILxdcTfeXSsE+4GE0of97TtiYN7A/gC
+RfjpurLH8meX9/kwItFWp0aZ5PWfeWgUq1qXUJ1rYShu0qMaTFAXFm/OoAptHgn
G78S8tjqBeSb1FgBogZqOzwtD/v/jcKN0F/605h2wIMN1QMK+eO+BcpNBL6yGcwb
f6L/6Y3SIoE9Gwf9ualmGExvcEwdsrk3zTPiImdy77q6jLpRzywUywiGyC7R6w6Q
pnYNYxDpxeRuUXIABiQfE8+FaoR+8i6g86BdgNo7CzxvVedo12iHaemWpkrSDNB/
19DNkj7X1Iw54pM1syywS5vjgo+UZGeJxw50y/WvCaFjWiZY7+XOKsHTjwRCRdF9
qg12TYxaGfNhg1cXPEuxedxk5EqbF3ZYYS5ZQPpVjvte6dZPHaUQqn5A5ETcLjvA
bOaV/hUnF4S3PwIibap2sl0ZYwQ06pfPn469PSvO+ERhqsysiGhuZLksU2fLwGpM
TGYBDUcL6mDH0vhTn/lV7jhT+ryRii3NG2163j4+w0tQU/IUpMtQGLQqTnq6PDTC
Ixl7V/xEG10s+9DYo+CcN1Cpme+w4GP6HMtSOtK+wgBLKdFup8ZuIC5Q1CUx5A8j
SqEEu9mdF/IpzxbRx+GvXQYJ3oWKvPXKKvIWfAGiU2kYZ529J3cXLru0Myuwo6yj
tOc0L1dhrgQCtlPnru/am+pcXzYZizAWJi0sUeW7FilCnK9OC1429xioAat3Vv5f
UKrJDx6Sy4ZmHpIn+5W9t2dOAt3ipFnpB/gcO310Sb+1aFLB1dwebAyQuzkA+xRI
w6mkDTOFN4JpN/wbXy8f5HUGj151JqhBxm91t+8F27Flpb1HZvKDK5HLG88Wya/W
Me7fyRq9kn3UuYuOO5c0w7DJ2C95Rp95I9h4c2p25/8vNsh3ff36aYpTeAL2fKdg
TvmtxKeZ+3nQNR+okYZ9QCPMLrk0r044BK19uycb4usL2b3OZt0l6PRDTcpiUM3k
sE788nWlvECrEnUtaivHupw879NWv+eeDFtdOTX2IE6kfsH8fhrbaLD5dF45928c
FunDqy5thiXldbZqAg3z6uADS6ONrxrmbL7ab54ourWvRMFeg0yRGcqQZZJSkLaO
Wt8UzwO8zTDeVuSBfmrzQNJba04aZikC0HtsnXxEDJXL7HYdp5W3qIbWBb/pC5ig
wFK0oHMTge+NADWyUA/SKmtbHDUdJP40nBYQzu0JmEZV9OliSVNBMfbKpIbYXC0x
uix9HeWuTZbcfKj66fR+opHmcXJxGZFRUQPqwTmmZeCqCxUKP3K26daTsWTCLbLY
63ytGFgo7PhkiHDEIRR6OUgOnCSiG4vfQdO3hmeYdNFvUXWIO1A0hR30Y6i1sZrA
9UuhFn8swdHqPhAlvIp6dv+1KtiDoOUUKO7sJ2HcQp+ZeD77ZCttWN2yFi0ULrKy
Tlb/+I/oXrnAO3NlJPOfkvX+cLZi3JLOrGkjb2mKhrZsIW7LdGsriuYB1PQmTdQj
EF0VBNrzqINcS9R1rgqaoFdVVxL474pXFhe23lXSznwwhU5a9Df9VLkwgRrAGikL
rMnC102a4VN5ygy9BzgikgduZiuRYKSriUbc1eL1zcbQi3IIzdmOwk9hLoi+N3hc
WmQtjB0E4iyYdRqytqaqL0tgoo1EloMVBW1GfGCGIqWkH+dzGDz13zvmrGRODU/C
Fw2ikRRBgb+T9B8hbV/GA6QNAOANiWbkfB7+sJU3K79tqGB2ZZemphAnjFjRRuZi
0PvxEDIzSJTPEmKnGG0wDxfTWrcx3IpicUttegOQpSNpOvJ/YeDLfkQBC4sBr5aK
iVpB7r21Uff0WugU2+MF+6yfMn2n1zT/2ohmeQ0B+QfpJ2D2t/lt8NMXniDppRZx
xRJTg4CNDxSqXvXf8LHDt5Z5AYZ9PynVcPgyXRZ3dlM4wDffORqGjBzQ/LkiNzz7
HrHniqZPqW4cMrwhAy76EJchWoalRK7B76QMkjj4G/8KrunhjY0hu6mLhIyup29W
XxfOR38cOE5yP6ik38GioXcb6g9B3bZ0kGYCHb6XnCKdDwt+MGMIoaMwbmtvseTV
wVP4TzvzN3q/nHWMyGU4t8e4oP/cygB0yRuG2NzxcKMyOeZVbCkDK90/SROxZZZ0
O2/MikhS3etw1+Txf6srYt4yy/gtgCsQnKBl9NpusTIK8KrzFQQMsNeotSaP02kE
nqNkqdEBDawYvcZLZRjI4hUqlnD48euRTz9IQGd5xCVROa4m1BHUO2JZmaRyhO1e
Ho+YofIjE/o8wcF01Onzrbpe7CBvmtGJrQbaQ172jbec/CvZ8NUqwWK3tQlKtMbr
hIVxO09q8TzKc5lPi4CT7Y7iIFZIm4uAPlNeHZzroHirnoW6FDvchXz+RpT/gVrd
ywaF0lDQgySVcXMuz22FpYgqMkYuQYfUwOLECwDqgZoL00xi8d7Qk9RWIY0D/kF8
zCMxPFxOQZrVo/FCVrHex4ZMydoN4qy+X/0gcgoovdkKoVpu1civyMALhuB2KFR4
3JY8Sks7lPoVsf9mIIoiy5FkWJ0Jnta9RYazXN2+n4fArgI5LrRpFq+K0D4pKEGT
Y+E+JfatVcSNcjUnZtnHNcDcybQQlkzafpBDBNeCh61xo8ILvy7cLiXoeSm6uj16
mavHWIIF9FSpna9SvZBh/mmMzluD9SgbgEXm/nDBNZFTvwn94u1+7SZC8b4aG/kY
wBw1FnKOeLHuWPZ8vPLbLqFMTAymtqygVo+bUjdVRtmm/3ATtWFUOsZBTFrFcE6J
05K7JBQpsespkeWNgk+SKZ+GkuydQEaznz73kpWimFvExlJcLvoqocmN1exr4o5F
je2raPwAi8i9CB4EmyaWe/wDQ8JQJRV0HnlpKBiE+MpceKYNvdY3LlDFXc6ffL7n
tWqOMAxbSsOc481aJSVzX6hliI5d7yME0xJmQ7yIpx0pe++ZmSn3EIYP+3iLnQwt
nidp+Qn9BPQt3pb9UNOxpF7EenDVJFMOm2fCejcE2gDejvZ3Ec6gUPQeNQeeC8aE
jdKV2o+lHbmADfnUIBJ/kZBCW6diY9lnOdIZchThlZW1qK9i9gTJNqt8a45Ys1Ug
IuZaWGvZGbp3q0G4w26L9buSIZLEHKcqtNV+F1QmHJND/sSxt2NfY05kZU/evnQ2
sx2VoSEpAEKeU7wrL4hdpjHOuFEmWy80jSQMuZoejFg6y4db/Cu9vWYZnOoNLlho
gXlNit+P+y7fb0VXtV6lYngLGuhvdvYrk6e9/lyK3qJaPv6Lk2xj6mHseprN+OlL
pKqnKG+RdK1UHIVwXAMXASOjM3f1rUpA0VYMOsaMNscH8NvRi17gw76WITbaTrKP
AWNE4rihFjJ5u1y4JCFOD1UfWlFCr7rBLquvpC2zlfnbKF1ZPlnUQ310EPQ8obNG
W7ZDM0Ze8REW4F9SduN4NGnasLkVPBzHtfcv1CueBFDoQQ4naCRhVHe1y7yDBKxc
0RovFr2CGdxtcutofoU+Zmd8FUlF1L0o44LYfQ8W5M0uSN4AkGXc1dkEIICcSz2j
l91e9oIrIpwplWoOQKCjfsQfthaj8sA1L/BYjMI2GBY46bvt/JBJLfTMPRzJ9R3h
i2fXWt4xibgdTQ6upHm1RBzi07Fa4l1uHz2NHsQbmOVC6j9FkAAFKjgCmI2oqp7U
37/CEqMx96LJz/sOUojZQGU3XwZHCgkKXo2BBnAw7KZFG9xcqSEzCA75+9e1KlWW
6JB8vpwXUmztZsXTiaO13XrwRWQNBQOnr4feLVUHMibc/miZ74puEfc9WUOB7nDs
Mmr6YX3rB7xDzzSJKC07Iq29tQsKGOEHzNFeh7o+I8BSXE+1XIan5CYiYrcwMLwr
zhERwive6FIebZClXL+AU7nDjX0gr3vPWLj/cE2UFy2pNZCgs49hNttj4MAvFQTB
uX22wb1NyGj+SS9LJ+kDGkEw2xEhBUv4mncgvmLxFGFpEY2x3+D3XqWocenOOeAu
4UTO+VRl+Ij7D7S1ajaUwVJT1HhVbFecWc94Aeh5Qutjwxrzn+usyuLkIAtjUcaQ
VHQnaWp8SIU6tEuK6hwiQIEoEI1kIKgotg0YYRlVedFgLHHq5axmR0VJ0+HGGUB2
MWnlrwwCV2PYM3D/sxYIGtok5C4ecpNF3V7WbYYRGkaXaqRgnm7lrASoRNHc3ghN
3GZiaelGAJOUiOARDasnCEJREWb6HL4u8kgAKkJ8t8yWSo5cErFTf4T7k6BL3yNU
Q7cQvaKYFQsdS46J/WeZCEGGK4zHuuQnwpatxRcauiMoaplzIJSJ5fP1t72NkbQ6
qSsr4+gV88T0FVJqF59Mr0yDjjylKg4z1LKqabz7jzTe7+7p+voKQLD5NSn9qS+Y
FQsEQHWlhnlATUExVbOTRuLZi0c4pKv0QkeHqLSVmGoDXz8oggpth9VrGa3Cyovd
/AvMkyL63xW/5u48+4xdQ2seTV42YRMWXapEVQUmvc6MQH32Os0RjM5vkhnFlw5G
PcjGDA4a9TChf9VqM6lv5kOFh7WgAK6wz4nMtv09WNzhIZK57libsfncpKuhSilX
LBwGiKMA0UdishdKL840gW/+MhiFADB2v1Db64d1cz/yfKOlUHHDk6qaO+ZmNGrV
rfzcv7Jv3FlpluavrtV4MjjQtBfLD42azY1ijtclVQbFphvXyvXJ7WLbiZAtG8wQ
85JLdXsDMhoSDxUHGG1WN3IYI2JStf7O/fqDtkFTRd0n33kxK9SPf/k+xHika55o
cCPcuveqnFdiIXD1OelVp369M6byfV0sz0ZQn1Ptj8NZahG5v98lQYMeY/F1LtM5
X3tBwTVRHgySgnc/13I2nxkN2zzKL+KYU053X2fl7KykXE7sOIuAtHOMqtPWnCZ3
V5DphdcKgJjBKuECqXoEX2e9iVG1Hdmavm0C4iFa/QOIMW5ecNq6+q6sFIqxvGuX
iEt8hc/0Mx/tP31SlS3tbYqqNqUrUZc7iKKzAOK/0yNJsxZE9qc22vyn15x3rCbK
Z2lFQk1fsaLmmttm2eAuAccXxgyOj4Tw42zUEMO3SpEbQAgKz5bV1MjRNCyvyt9h
SttQmfkwmV3urfKmpq5Qk4OwrWcK49+dJuAIL5XoDseeLCUJOkwlkIQW1y5q8kfz
8Qh/ykfFuCXWqbzC9LwhOaZin5+6swkUslap7wTExiOjk6S4WUfcpaK23njEm0W5
G+1LWj13GbYTRcVUP/zfoF1DLOgm3H8ITZU2BWlgFFrfYa80kMakgnKd1M6EAlsS
+29j00qsI2JVXjkbFJmWsaAxJOHpYhskz9bhN690fhs/oNWS2I6h6n8eGTMCjpd4
nTuSDyvFaws49dQZz0fyCerEgtIzoacC3z7jJFwMhFBuXn8qTvzdAQ+yeJ3zP/2N
jjfhJiZZbBXSxOeAE3PZlWAjsWGfZzmXSk5BDjYYFss9OBD6drjqErTZWbO0aCi5
Jz9sZGODU/8Mog6Fylw2AF+3H0mcl08mW6XF3VoAtPBFItUQWG0xgspslcRjN60P
LsyS4ceAS8ypyK55OUL2Krj7kRyf7sHVNCaZ6ggEWKTcYzHlbngU+OVrSfspFPpN
D2vzjA1Z/df353X62RSWLwP73lPCIQ1BY0+UcM7uXkX4tWG2IJtMDsidSJcLztOf
27XSMx8kUWNTHjH9dC4kwf3lRvYF6tjZ2MqzFUpbvSrqJgJ4ScQkiQKzACpE+s6E
v5Qdv5+5eSIsWQMHXPNaJ1iEsu6PXUMSLonDedgoNdMsDymRw9k27hoQnblvTNce
3f4xY/JGlnZxMRoDuRtTKPaezmcLY37V+HY357ZBds+4NeHFikcw+P4oqoRUUB8d
Wd8WzBk4UUHq/agpmzS7AuN6UI4JfHXv5Q4feE8OjVWytjsekkekR+3II7IFeFbq
476tHAHTjbhhpNd+uJoF92zssD1c4r7wh84fuKzagh2m7Lk657SJDaZ/pJOY8Iqh
/ibD6dfOyklwd5ds9W8eVkFcZVFznWVSYlsgsjc8+E2nYKCq1c/wlJMxsnceSEEe
2dqxHr3t/jSkkETYnS4DULvSraJWBjxOnAsnKHS7/p5W8bM46YZ7l+UIRYuFS14o
Xbx90g10aqwRGZ3sxnrv6FFuHWqZi1nmbXSBvkDOwAO1vuEUwxwjpZfwzs7RFoDZ
sdXf+znPPPZT6kXP6b5gkCUYClxbCA7soi3muTsJWujU21/rzRJiW50SXv8M0uPu
F9Li8d3gaJWKp0psZGL+ASDargWoQTo1IFCxGmTwPI7aRiUw2GVO5fP5LeH/GSaC
wuZ6bNWXI3ib3nlJpys9BScw2yPhMgC1MpVSijGXsgHSlI57+2z8958FtMTsNCEC
o6wo7yJWHHf1uHgM1pHxcgGYRnvv71pPTEFiny7P3qkB38RdtSRzMqLosgM42Mmc
sDOUETtOFggDzBofrT13TVRHdkmMDN9t2yBWn0OiF8oEmPxmNICT/yh/JwoTVThN
e4KnpMym/YHOZMF8imlpvpi5c4dGfCpIkuWA4i3e84a5r5yq04vLA5vNcboTxvyp
3Wy9j+zOAS22RFYvTIbdj5tmPOkJZO/A3Hr7i41ejWBXEY/otEXdfBg1q19l7m8f
IBXJMi4SuJdds9AQnAr+aTFkfcGIQfZCyCDXvx/2s6qf7quGhc97jaeSkTaqCREU
qrf4RYderUl5agh5HW1isxPgV1xAhhFFr4t6x4pTqZRdItoyhd6qDo46hh7peesH
Yz8O3tBLL5ClvpBWpYNzV+qwigGOzuaxxDDtK02qcNO3GySOG/WpayOyvba8/k0B
ZyfkDWGAjyS9inNV3g6DfU22RGWIgEN/X4KH34W2kxG3jzomd45vTJZsOYbKpLDA
5R/sjIgNYCviunX5G45/SWAdInhdvBewWMZN8Jlz2NiLjcZmut6ykyGZZlQQsUmn
bDI5I7dVWkOMpRj84HPWi4LeSsBayqg/tOuBNWa97di1jWU5RLTBkoN9aHQrM8tl
uci/S41G7zcEw9+yO83jTQjGizG7h40bb+WwpBjnIGWK59R2Ee57B96gIbWS90W0
dMBpzgW9yGdMmgon4kbwc0W2xoa+ClTLXoN5ACNsB/Tpx09hkRib2smQD+yjxwBS
NH+rWg6q9+NZK0xYo9/m4ZFkbsaTnsiBLyTjuphDq9lPOrdUXu3cUkbns6YmjkAL
X4/xREAaapOSk9MrUjc+M5jjv+eJIDTkRDwg04lLK4a2a3hAWKmZJZxMq1Nj3SSG
dHWnkRtZc9qpLG1vQ8g1xr602i4TBYeFDqhyX0kSNgObuBPOb3/eduBUmtQsuJpr
G2uCqmpMPTmEduE4RuZY6uy2J8yFeneHtPG9jL3+v2XDSPWfdSkwLCyC5vdZeLFE
C7YOkNakZ+ZlDWqUEcoTv3FD8EYzrPLOgIWT7QhYKehbR3i7RgJhlnLGteSJMG5B
W4p7EsHqGfh6JmoNd99gNQpsfyL1vxRi2qxEeuyAbAwAJ27ZE1CJ+3jjpOYc26nk
oZ7PVprucpgS4xF//hsD75GIYN9o6IG5WJtsVnn2uVIz2FEmdVlGtRSzgMOhf98K
IQ0LXDUx9YNtjTrx/agVMSkuv1y8hzkaZvLOS5tLdNraSVcRsG+9YHTZI//U3FKg
1Nkgda6pVO+7Yw9IHtvBkKelTs1/UbvgZWkO4qdPAJzQdJjjjCEhOo0wqhi3dSsb
dYw5mcICJFBxmOFAedKKhB1YYDpBho5hhrtdxTJDgo1DwhMiy8yPa6eqpncCJDZQ
6zXZtfjlQrJDxSASut0epu4tN/wn2/Zc07i2aD3DOgDsbOe0XVPFYJhpFHAn7+9G
Plo+Kv0985/86Z0qlyfXfFS0xHAMIOzAbhxdhhE4G3p8DuuFE4FhKEHpii3jhD67
DJFm9ZLv81wOrib/ocZO6Lq1REya73y71iSsC/zbC5VX9E0Pv9eYOXaACxP7wefF
MwXahXWG9yvLYibwR5swBV2w81k0yY/l+IwZvxusqeHbXuviai1GuwYE1yQALWpl
ksGTBUNQ/UocZGW1127+dZaSLFSj+i4l0wCReJc4kGMix7Nnqr7m4LhbZIswvL7k
9WVpWNApDcMXNi24nGgpeK8wJIYjWRRmcAmY/Aka19+X8xkYGeiWmmUi6l7cb+bH
i5y+I16/L0nooXQ88TKXaYxXcNRQV1ntKLQjmYfjlBWq9BnQrqN4J+safDVtD99a
pW0N96fhXs4WwR1nVHFSTAiUwH37L1QnkhlB9evW2A1DHnjddCLh3MT9YYa7WvDq
EYE3t0dt539FxBXbV7sKwBmgkIzHv2kxL7VzTlkGwOx0qGj78DYxPQnN/+Tp6C3x
Bpn1hApGpsqT8ffcOnCgh/FORx1N3J7LLd7HaWEhowtXa4Mwd465AUIS4PU68m5x
Ghbz6t2FVeKe8lDSKGhT+aYjB8h/4rHnzG9D4UF6HuEv4mOGFIwLoYg1r+vHOlZn
lUnBq2TFDL/4ZVoUBNiVfmktJI/YjpCVSJlxxbTupk0wiFA1qUIzTJVTQnJYQKbO
zG44hsDv2rnrALYy9BFVvW3wrSCFGDkJTt+nFod6vKxyVFRPtBtMgW2MgTTQd+oX
DLqkV9ZVwyyBtOb0bdixARe1ud3GeLJEjCAvL2pRgAxfHeJMVQrX2VKJeitpu0hd
O1sGEFBJK0srsj4db2xrfmStA+6+CLeFaTobwh1zPq8LSAnmEkAA5oOWUb1DciRf
m6UV9CElqrPtmY3u1Pxl4WNOkANTJ46MamYjl6JuY7AZfTisaDgjYY5sZBiArfgA
pU98Kug8zyw4taFHmqj7qbPJbAnGVPikWsVDG5uK2WqTfn7xzL0B+mpg+F6Vq05E
16Gojmpxv7woQob9+cc9IK8J2KXm+pNBvKBGYL9Gm5oU7caViQWtHQsmbVcqmwgM
5fgDZjyo3AujmPzxDqYKHxXqNXXb0xLM7RBxEIX5WXbHZWeTWN4F1q0W3TVzitER
owIxqYkUdBa37U6tynHwNPaJJWiu6j5ntwdF1tY/XWFrws1WeWDdVqwwWiftqMMU
JtWhi8wS/SXVqQmHQH8Z1vKtoXL/ALedtOBBhBHgk1L5BMJuFq1Ml7EWZEHJJrKy
7YYx9ZvisIZBKcTARCQp9rzXXaHhACkS8nkH4h59Oyih+fpSIStJhUQ0cfZn79CZ
Qz1cJEsdwc+ES5vro6eytykQwVjU1+9qmaZsmbmJjl/MatOdGa9u7K0t7Cvz7VaJ
yv+uFhl4NH+KxL6uY4+acxuKTDsSJk4jrUWtRau6Zw+zPb8Fd9+2gEgalPc9VRoH
C9HDceN8ZwdLog2KgQ7OGWPD6sWcPbDOS/1pelRsbFVL7dTWoVMlrbpdB0qntBJU
W5Akqd+kURzKI3p+7l+7dOpk5RoYpbEJ7tKiZtiav3tetomgMfQzgyeE8Ia47a0N
8xeWLw/hwnMfkTmsBenT+/vS4+6ZIJuVy+HcADlFhGFXB9PYvad+dMlZk1QRXs0o
CeH85tucbrU2uryKoLNa57koP8+y7Y9PDMauFh5t0whi2Lexogef263d6zdwvIO6
gdxovyI33rwM/6ms1ugudchqi7dvJ8zuMR/zRCUCpPhb4+DRZBlWNK7gKcPMcls7
hw8aMPhKe86f/Qoic9+mOp32tOIbp0TID9JNXNYEEMaAB5HXrKp3NkQsavgRYA0N
TzUOpDFbntfUt/+Xv4eC9Rc4X6ADZuQzYQb/6ZCYJRpww24YWe8kdlDByaG49xxP
QWPnWIBKaWqrN+1ZEAM3u6lwm7Romh5gg6AHefGVFSODnArfC+3d5FpZ+lzVMywI
NMLkR53FCeOK60P/jxWWs/z/ER22oJ6z68y6KQvAyWQ+eVBr5CEjD+yQ24VaNQRv
LNL+Gktsgg18m3rfwe3rCqy4TFQmJLjXMrbMFMzU5iu/BB5CsMSxE4RqdtaafILd
4x/SlQygUMiy9qiLz+E3hb2UPQNH64LGxXafjagBKPdOhEx4RTrhIn3DVoM3F9Ow
GOvPnR8lgDVoiz8okxtROlSGfrMegRZ9B39YbGD45B//emyqX+jt9FxrjvdM9sXJ
q1W8pRLAM2MvAn4jQZ8bXs+MQfphYdpIytMQqM1Q7/YP9mPDOAfzg/8Fj0rbnoBD
c4LWtHeSWc4emI4l8pN4zH6WFY534Z5D7bgyBAlHmPKx3gBUCvT8H263QyoBA0Qc
At7pHEEyDpO8KG/OFamR691pGIaWhyzEyiyfTjSK/X0G9FY0d66t9/yJWF4r6JN9
cU/hd2Kui9VV5X/jSI1TzodqB1HPMiBFjpX4LAH80rdeZep9Uk+0QclbpjLYnU9w
74O5a43sRxG5mmj5EDAglQqsi1d9TlH1zqTLhYkw9qpxt04KyjCDrrqweTHaBiRY
d5I9mmA7wNHhaScNMNAXaDeLo4Mn5JETQ51dCp2H/Xz0/4L3icbsP8x1IxlEFUVh
lFSud/pvaC7XIs4HC1LMrCx6O2R4sWNzaE9JyLWdrvMOZPpXscafSmEHHQ02VxWH
/SRJg5UfcR+4d4cswbYEabomaZjyCsMfB4yklWWX0rYBaVhVjUYoCLrR7WV4MJ/O
6gGtfH8wid2aEZWGXSCylJIn/6OL98/ZVcx9PZkqNXoSpUbNxPJHLTqYDliKO5/w
oAyUAl3ax+7VRIUMXrmwffqfbot0SKHe8XDRdrbcc6tDT5R6wE5HwlJhrKX0gPBt
JE4oHytDV596coLHp8ji/PuyBw7v1fEGy6txqJSP0FaNaiUHSxrTDWZj0UVQqlke
XogOcAheBSYdvrr99pqgYY8juzo2crKUvS/rTPGhiB+LUubOQloDO9BAC9aVOimb
iDyX5aj5tInxrwoZIbKI/YCLldkcfMFf4ha1po0WpEJRZh3nD8zRLDKR4oFFFFlR
YLrCX0ou1cAa3htGTJtsAwpmOfzwiJ8O6Ocy1f32XcsjWrNSB9gSko+cwx92U6Nh
dTjGu5EjRUR76+fr+nOWWtOn9/7mczPaZe2P/G3D7jfegd0jhwPghGyBeO0IoUpo
JaiunhxavGqSyRmRuEm0hM9we86oxd9BBXSykD+/GvM6kY8oftyOCaIVfy9rPEWp
PACTh8Xdqk4DymhzWT5GbvfBP/0EQJPLJnC4BWSTa2lFu9I3b2z7Wr8uqzPTZ8N/
hb510wreq/kaQyhUPlrF/vyK7uXtbSy+KAfI3omyg1r1DEZUvIUerb9rhA1iRxLk
Azpe9YF1fHDQrx/OIltUe13wTq/icJR+0bB+wQtn5wbr2Q+564STLtlTlC0vLDzi
37ldmY9iczr3ubAMl73eznkMoFCr2yuQJSt7WYgPQfwLAe35G6Y+5oiZvB/L8pu0
zEk3oQ2uCn4qD6imyRF+3W1LmslcCjBcTdU18eqlYuuN0DGYwBXH0lsDm+okJwu+
L9JuFDP04Ph/qZ9SJ+lJm+baz0E9d97KwyFIJ7qcbOeuBD90PsOeczSOpIJ0ybGZ
kyRX7dYYquqfdFWmEHvGethvQW8YRie4QkeqlpM4SmjegE13IhpKJLoqQbxQgjv5
R9TKQmMcQeryfCpfaQQjyosXmqGzS3xtKpZi2mZ6u4E/O56Nmugxs9Ak6sofCkju
U0rAwx1mLKN+sRtGAIfqzLMtZfI4GAKauL//AsvrWoCbjO7iC/z0ZmNln5bYYAJr
IRTuHwuXOH+/oFyfQAW88ke9nXhU5mwjJAGqdYPjZnUdLaVKve8LHuUq37wMqoV+
i6sxwHsJztT3rRHmMxhvlouUFxIhvc6CeuVn9AMn5HJ3iK/Ng5srlK+5iwAdtxvK
d6NytIuUhmBgxZDSgpaQIw18HLgG+ssZm/yT/WThMlKq18TEQbFKYLIBJbI6srxk
niXIZ0j4/Y7WP705fhJa2zTz+6DDwAPd/fzgEhmgqxQ9Njcbxt63sU/gBawCLb2/
c1wfb3c5gFdgahOvjnEtq5gW9KzEMAHKlZWgPDTjJqdkD55Bp9U8JGZuQPaDnqqM
TIBRmnMhmIcZgbNbXfprh5Jt9q3TxS/BysbIDPFx3/rq7VhDVvSgT2G/b999DZHR
MMOis1h3gQHg5S1mLuMP0DORi7C+AmalwJbLyXwJ92EsCHGSPmsahgf9QpcXUDe5
VARiFrO1ukZkmX0UMNMDQA+j7q3rW7OBXkNVD0hxDMsfQNdCNO0GR37NWzqFYKCe
YRR7oqWFow/dlC0ayYb2/ZIa2ZhdqjbMWgj1C16NsmIrplv3KFjV2H/juKxVPV8X
zWGGuoU8t9z2zGi7vq7Xam75mltYVzpXEI9zZbc9urrYjWl7B4su+YXsTtIyYQCi
/tHS84h/OOF8qseOP0gQkQuHgA7WHwzViy4qOi5bZQVeHPd9H6ueya72two4lzKr
FDlJCoMP1sgjMh4Xfx7uFrbkZbKxG89OonF8XOO9xOBwCyVhpjph9RM3doQBOF9H
pIiFN6xI9vutfYMW+xayEgexJCYVzOum0TcR5vckjsaoLhTA5lL6u7DLzhrnlSnb
NSF7vn1QDuZtfxOOg0hd63k+QTIYQ+2FlcamT0uZQS69jMWTjQ/gHoaftTFYIqjI
Oh3JDERNS5umZyvTOXF116eQVJicCcJt09hzLNGX1Fy7tBZRaMEG8akOYHChv1UC
wtkkM5u5I8w+DhTERM6pEVdcsuIIKjj6FJkhgISjmWsYoWdL5dgmw6uG42KPpLks
SOKk5oYeUkSXpU//Y4lCz9dg1/NeEKSTJfkDgdbe1WGLdcb7uBUDRo0KBa5a1tNM
/Uf+OwxPBKLfHE1OW9t7ikGjBsk2c8SKeBkmPNaD0d/Go1nwHBjmnQq8ssWyrc3x
wTwrITiXlNFuXZPvhpmTUjllwUwWlYPyT6K8sBF/dW0n9moUqyrR8EP6llo51qIH
eyu5abFRAa2U5i2RhNsR3zTtghzrWpf5l+zAN15B+cGOhZ+/PlgHxAtBQPP4KqrZ
HXHiP3ZWR1FtOc+ndxlzvLJCRUU0hZFlvFRrTp29KywSktG87bDncct86OMpl6Nh
F0eUlMxE4nS99A3OMO5I0Tsl0IkeXtIhIb1x6a5o1hUA4EYpCcX1gNQb1kBFWcox
Io/IRWTqSeliJTueQM2HInSFqWTBlORhiuyOSeIe15opoRIuQP5RhPbCO31ygstR
+wcPgRCQgtfp2rCykdSsE+q52Ca3og0zHPGz4Mn0QWFeySo/FYeYadYwY5IHR+q+
a6M22XXYD0Rrn77oB5mi3uBACqQcAm+O+OYDTThkGQfE+9+9KPWFwnGMPAxSPBE8
q3ZXeSz2zzoSxxU/G7c5DX5IowDjXB3Ja3Z3kB0w8QjK/9TQxayLf5zmTCoXXl8J
A5EsJXLNkAW7MmqmM8AlyyUuuGHbhPFV9NcP3pnadVpqqzP+1AMVfRg2WXln6r5i
m7xunGeHOTVqq0cQU4eyAKnNICDlcnMB+CBwa0mk0qiunu5jiLquy3bMtHidQf3V
jpE7Vzj1sgbeyWBNcWnkGD56C46N3c+eXgNLkRE9ieJsZMqm+oPOK875NXc+6lfq
SERUlJKxQ8PaocV1tuySEg0H4dnm04sxyMM5fdoE7UtAwDPAjHfBfXyNEhGa9og7
JNOUFllNE8SYD3PllSNhSBA74KsXW6ajg1ALe9lk32WgCZlRxl1sQxVX08ttQ8l+
liwKWSQM+jX8PeS7lVtb+IZuo9CDPbbSsWROaElQs1AKOt/K506Y096rFRmZkr3S
p8yVVggm1vPwo0ZQzK4uZqYAtTD5ChmTN8frMr5iCBUh2oj7FCZDaQ88bpd1iK03
ZuM8ZbTgh6lymayrOVbJiKgL5rddzaFM4RuyJ/N0nbUhjsFREZefexyR6IZ4A73F
04VBUg0jJJNxHheKhFA7Ej5e8tuZQyRe3RQctbZoU9myYd1/T0eZ0E5UcMxKtdoe
TZ851D//KT+G3LkFMQXsm/mQYVmqbm5F8Lb6Lq/OjiEXvBzammZJrf5KSW0k4Uaq
ihiOhE3917+d7w0NsqLDfN2kqyDpbq/868B5G+kyTBEyciEw2YWro2MdtTGxbwHS
/HHVIe+x69u2NkFvYb8ydrjKKsjNU0PHGvQaat2xr13w6QoLKwkxGpHnORC1HKSr
FNyFBab4NWQCIjmKz0mT8Y00Mke0/dtPjNkLLE5yvTSXI9NdQZgSBLeQf/+IcImC
J+OYC0RsgQ+PxuoGWQVZhrRkGvWAhD1zct4W5HC7/r4cLHFDNXHcqc/Pt3UALW5Z
UGXbLg9ZPWH37DObJO5qI7ZMB61uICxPMjUfL9ChUd/00dB+To6HEOkWvuVwkobn
6+vZP4nOBpdgnUXK/2/Y2KacmSrRjlaA0Ukr0M4web8r2kL+QsucPI4VbcoAfqZF
AM8aVKTfABdh8DmSdP9+zPHcYJaqzWO9YoRndBE7i3rNwCV8UHUDhNEe+B5fbIHr
JJWTRVmd9JlmNaNFShoJ927XmYRSHW1ooiExMaioQ/7gvKL2KaJBEwx/WTxbvfYb
UrSHmy3B7y+jgpvrvLRFYP4th7gKSg5xqnQrJTuKJ4kdHbr17HJjLyE/8tRSCyhY
3aZRq2FE8w9uYDoV1Y8hH4GXG1FHdaPd9T5aAMyqyyoipIl39pmVmE4uoeKHNEmX
X5U+/EfdiGCeJ9TOixDw7sYiC8Yj8oyPQ32ThuXULSq/6TuZFP/bVtlbr0crZh9V
bRZ5v4yLBSXLuzAIdvc7kStCtHGEhZ/bdcqC/6BoEdOGyQb19DLCPVqUElpSbZ6Y
3af2Ybrw36D+bvLnFJaHgEQqeeKbKvYNe6jMv2zQANAfMNAbQZv/SrUGpPi8Ldvu
aO+7T9JjPZgNXGezuM4pkH8JoD38HDellIq0lLdeNhCMwoP7viPrSdXjU2QRFIlV
YakUz3hZ1392UZbisSMwrUpuGDD3kJ1o9qfB+Yuxq3zqmKyP1Vj2RQ1GRwSGe78Y
YNc7DqJAml1TZSWalOtDLK8XWeYj8m1mUJ8P5yeS+jYeuVg7H6Cocy8oQpf0e1no
u+SNjnVrnBeQvbnBpP6LJLLs3RhkNOGVJ67vU3W3jJvC+sBRUI2l8S1zNAmx5gW2
0WX+Y2Ki2b3lj2ZhD1OWqPwBCWt7cG3LRgzlLXetNhXqbsxSksp3bBhEnzD35PdX
44DttlBPF+Pm0rhFfG3d6nhDg5wXKyCB6C9UZuoSzt+VCvo9ps/Yt2Fnz53xeh03
/ew1W3Gox0xSPU5xNhOT7Z/d46NxP5ecnz+fjIqbor4Yq38DAGOo/y9FqhN12wrD
epNRhLgDXNLINvaP6mejOu5DQ86dX6nG1sWEu2UQgmSvMxkOfMEI6f8GoJ4MsENt
5E23msQcTXykLiuY05oxtVn0F2TSqWcWbPAv3U6v1U8AVNGuS2SEW3ObdhbjgvCU
2qJiStN/z0kJG0+41qloNWUrVWcUb9rOpdlFVAltR1/0TCRADt3Z2oVyFhW/8GoB
k5/2tW03/4OtUCZB9ZBhaLVtEJXInr6+p8HcmdFJKID+s1l9OWzARsqF7yo5IHvt
yvwU7YpBT9cDwX1xOvVBq6gFP6kCoRdhXgPCXs4NSa4NleMHsHYtpk+1mHMzg3AC
G+yQPhqYG7S3ODDdhsOm1TxjsCkdCnDmKiG7UZCDcCZnbPmXFbEEZmXe66xSWVnj
MAqmMRoNW3ukqLKPItwg6gDjMrCok7ss9lbQbQnuweUU0kyOrib0tAikiSCv7FXD
z8u4QQ9E+S23XWZY4WOWuzru1VM/hqvR2wPoQbTciuFj3r3UtvGQmVPd9dHxj9pB
OjfSvpXWxrhHcPClDyfmsHzPgYeqZnd0jRtStixdV6ksXNeET54xExIm6zC2kWAl
QTJ2/X//q++1OxJHDW0m4bEt+eGGBEpBWyGGqiE5oeaznHT6uc1Ml8QEB0wCNnvL
2osMXWAd91sK4yYQgftW3xHsU14wiQQA4fnRhdUrF+GMiY1mPMnqR5CRcFRoVLjW
aDG1M38pw1dcWDhEKi9xycE0aHOqoM3xLZ16ZXAIZC9KLMZS0ePf18nI9+Hygw46
XEoc/WQKcDRwdMwPF6WSMX92YTjExf+AQgdNnwgtCjWPV5nmkTR8UwcGxMQ3kfvr
sRe+Lvc2H7m04s8riEqwXF6Gv5yjuz/ZEJ+TnwDzC2LBWtSGEVD152TBW7cinbI4
xTeVTUs4t/gRGjd0Fxv3v60E0U3Tvt7H7sI/CCknXw/vSNODpxBp+Y9dcO2yR2SA
Z9wyXs7EmXbIiWXEdfsQ2+/SbwQPmKiaXJrjCrPjshd1nFkitQC+Nqa4Si9rsgI6
CkP/jWjWH6FYq1AwR5qPRk5iVsoBCEIJEMSvLgskOWXxLsT2ZOombm+uneyi4oxF
6LwooNlrVx9k9+YR/veSOduBKYQUhvzGSIqel5qRyOA2cFH9W3u74VivdIMo79s3
nRWqcHywrKWG2AiWvxyOpIC0eRegprGkpXibP3w6VxIS7SybNzFOuc3hTZvX+7HL
JU/ykoMBdHAhwFKg7PMPUiTPtoq81JhndmD70WARaf/dFl+4e6rvIxL+NsbmykNO
iZVKuM21tp7izDAkWzxoK39dqCVqviEbf1fIbaCgM0oxkuTrmvo/yEN7Q0e7FUDQ
+Zant8/AHGmbCgHaHkJpCabqepQ3/zzlnOzhCFqxH+qt6vGJqIkU8nELdfOEfB+z
+qvVSOaHQVPisf+S96BXIFgJnGAkLIiRKWRtVenXranvGoFFKQTx3AaTnL/nzMX9
0zaK2UxCKGqyhD41rt3uXFkx5Z1XyN08lo1VyUt79l8YogoDv7w8WwW1K89m84jE
AJn2aqQxOndACCDdyO0brqKW/8jbO39idgZxoe2xORrt9vKubyZkVpbQbqwByO3E
gfaWYV/iTd+cH3NmaUS6Ij8Lh/OpoxwtznatSy679Uc7JpkhgtyCUqDGG9dav7cb
VX7H4PKeJNc3lKnHF0L5VID/zFmtd0O5SjNQXh7xZ3CVqp7ImF5tToYRxncmGcvr
D8PemUUPnsYLt3EIWKgbV8siQiL3faVpxNkwfiuwNi3Uzsg0NZoUAn102czZZtHW
tNa91JDvfhN8sLhjQBRrpyjQNvtBS5gs/oqERw4tQq336Shbl+yD4MT3OuKjL+K3
A2iatSfhQlmkuseaOozkz9dlOo4SDam3JerZYUi7lRm6dyZMoCRTix2+EQhLgpnX
Ss25xGgxt6tGCmhaKf1GMB81T36/KUaYhhnmTO4rqUneoWU+BxdP1T2+HxTLcUi/
wFJ5wGBEBajF9kWTMyAm5VPuIoGxEVQk1HbqIYuTP38k0O3dtnTOM6GC0gPOjLFh
E/oJgyIHfkGc1d8H6MMCAapjc+wwTZj0+Jr1LzcA399YIhzwTjyzU7mKt8SSNMOq
l3xIp4Idf6MvZno6KM9u/paWdhApb/5tX0YJmO46vPCXhbnX/jCp3RdQEZKF8Qud
YWJvPk6GBX5Rhh4o9RFJ1XrkVr9vBgagwumMt75+/jWY1La8HPvToBeEgNLzkJBN
n1nES65kbI5fmvqyDkuCdzv+eUk5eqAyY6q3cMXnQBmu7pXHyFKrLcDLGS7EMZGR
ZwGlzEH3U1D64rIzH2gA+poJWgSr/TnNN9ePrLbiZNZwO17wAIlwVrW2L1kRiizA
fxTTkCrwSKHWbULk0THaUNA+9WMDq9cQk1RK/gm4i40iN3ECrLdOg+qMdoi6Hjdd
o2vV8orhPBuV37k1qSPJhQa6kgxOhcDjmDdRkmLkT0xqCjR0IqMZO1dw+xr22ZDp
ynQ2twR1Lote/1YSGhxNYc/lClHzhYlCDJu2Txp/ld3g54T/pbRASXAKrSfeCwsH
qjZ4g2adaS5OnmN/J9KA6EgiaNUIBfGMEJOzDnlzu+lCHSXYzEJJ9yTEWREGLdvO
avvqmCjFvuqJ3E3lQumVMxgIvEUXi5Uo81ZdK/AEPAWC7WWo6/h2KgeO2i75uaxQ
xXcabgmlbPA7NMGPMwgqwjSlZcHtX9NCBNiE3v+LmfwiLAmfnRUm4qW2JpBD0p2e
SxC4/ti5kwEzt8z2y1rC7aymiD241V3XtgMlyWHJVTcqEZqHAv1IdO0ypalZmbkX
gfGnOuhlUzEA2gbcuR6lKmpU/AahiLkXRcaGKMVXZw6YTImodVDvCaJ6+6OdO28B
nizfwvLCG3bWS+YBqLyHW5C6vBLviaZeUNqpcqjnBqt6OxJQ9yLts7/LAWAvUGIU
VxLKPUgMq+WB4g3/LXyDhY+P1CYT9WpHelOqSnZupW3jO/wokXLn0/hCzNMQyVm7
UzT429lApx1VjJtZ6WqxcSrrK75wrmBQbiCMMl2W6vhQyPAlRWUpvtvyjmG35cfN
06ebXpdUO5QBoc8dqN9FJ/e6TrYjvcMVsSsgvPHJYfjb2wbjlqgEFTmqx/A8gFZk
/ukpDuPEh6KAOv98i44w0AeWNfQ8V9r2TmAwzLdlFx7Mq9/BSxowxzRWxiAcPmI3
fTjXiYc0YZIGmRf9twsV3UUbZN/VQ+SnoNVaRPc34PYdHKsxlTTuxAfMgzdAcODK
4ST1Hw+/q8Zi1nkplmmUuBCP2F3uqkcQVpRebIcEmqhPmZmyRid+Z1M4N+Z1ltwY
e8a3AbY1mhsyVDi8bQ0BWtcbUXKO1AkplcmgLyT6xJssfCaxKIuTG2dNKm2L4TDN
l5UHW+vqIlr475tfFtTkYsnn7Qa1uJmV6i8AnzEKG5NCKb/D/t4JnUCQCHVsJJPP
8bYvinBqfjjethwQYcldHzLEpPWpPev1yF3bJSNk3hfT+Dwcn9JAqzbQdfw3egpr
5T8Vw61PJud2dau7lrj5RBZKTTyMR+qK3fEe5D3XadlEcyrAYpbJ0N3BBXwsxF4l
hXC1sSlWGrtrnc79AagtkdM2yBaHEusCc7ks5qwjVyzIrHvxw94EbrWDc1vDa9Z9
9+2wgzVpkybGK2LP1eI60VTtyufoP/G8k6kvIUOZrVWkCyZ8P/DvPkuX2V7W/nzn
3wx0cF50Qg8wB9gLq6xf0LKhWJyd7Rq0NuiiVpFEePKenYD3VOXvbYIg87N7vgQP
Ah7VqQeDeyVuVZ+RQDYxvYHPKXqYSAS4z89Tyjvx1ZToqKxzCyl0U+/qf9+NcgYk
LBiTnczWxguWrcAJ1BpPUl3DKth96iS7rpalKylhaoMsU/f0TiJN24LYuK+k4GQ8
HLalZ3gTPxCD1hniSvPWz6J5L+pPPtljf0S+ZCc49nVe/Y8wMUrfOQtB+tMmJp9W
ebAfN0EM3e8akJsxwwpPeXauEIGH56shBbwmJbTSOJ/by1CpWoBxmzsQJhPpnfoJ
0gTHMrMcAOWrZtzxpOBiMFlrDQTyS0Ak0pQqZaE8KszHzZX4wDCHVcEUIXHVwPb0
LFLMJqow7yzz01CCoBu3pdVguhXEqHdbonC/iISPWZYOSWLYKHlRvUWEjVVKMHoP
MGsShzff2+VWJ12UqQlsp64vKMbTawicwsovBKlVWaWe7LsFPxqz2avMWXc8QMtz
t36Z67QACAJr+907Z3XA7sMDEQna7j7+xkJBp9YDcOvbuvbQOPrDdncBrA0nogmE
wr5x+mSkod/JwBCeoW2L66XIiJEpf0UKgIaYIhuzMQFo7nT6Rylv0o+N+UNc+fvi
vY78K1MzTB7pgqC5YpZA7b+r0SkQ9xVgtOqZAJAjLIn0K7fadgLNAjWD08JXvHvM
BSkaFHMQjbfGVborNJTP2hNQU0UtZ9V7AeYmPcJtONAGdWG2teeYqGQoKpxj+/SG
pKpZvZb4ZKnZm3dbF7vMBKN+siY1HneAMnKAOXCOrs+JCm5KF+jDSH15pIU954he
9sOZJlE8QYzlv1ImRk82p8lpL2zDwmupjbQvPd51WuMX3TZZw6k9NKt4991xzRCY
kVeIX1DnnYIaepfjhYhcm8AjyD/cpH4fgIVsutjAlZJ58GSCRS70BzEAmoTBJcJ/
hurjWS49tw+nBqM+Y2VT4+5yr0oyOC9ZZHNc7as5bGRgt0n9xf1o4AjntnmEqTW8
otLaTFE+AfLVIxSYfA5/MCbNXp6bkJfBR+jQW/p3vlx0a05VgKfndOckbF1oIfiE
DjuxtWGtA64fIJCYeGsuxSVzkLVw+1n6NOVKalrRPCU17M8wWG3I2qI/pA8vWRBU
k9/W4F9WX3wCpTWI4jy1ME9vhfxjUgs6MYqbZnbjS2/eZvi4s1T//IqnY7Zqdynp
m9uC0CXn5rinwVk1+y8ZTbN7vMJrrWP6wGJzL7hR6Gukmt6E9Uxid5cBrR1X38CI
pXWqTNpdd2G59hfRyPm3/vmRdHTxH1Q6jZV4zzSy9fuJlL0Izvl0ShGjfUc4g+cF
1FMB/7YawV7bqQje0fqcjkvXMtzEIoEwx//cvr6syPfa1cqyq6QBOvNyj5zwB0ay
o5sRWOf+vVX+McIaZmGMrG4PrwbV9f92IN0TEgxOfBopR6x+tZzMMW60wphrC5hw
80Y5Yy2SyjdZETHn63Ka+ez4JocruXzmRDoFajUXJBWcqNzLzN2InP/m1SKyRasx
EFMlmRez8t9YYkYq4Tn/Tp9oHkhXKC4k5M3kvcFdNhuwlkwmD+l/Rulvm8u+CMke
f95b5YCS7XK6bianvtSZ6pshEAWYprdvwfd5zxAe5xhQJ+2i+/CGEtm0aEb+wfWX
At+qYbfrKLP4QO7Hln1lvU4dz+MJLeCyYobh2tPa4kf3ABIpQUbKOCaq11FhANJo
KLAbNzxdRNXDropOfUfJoGyD3GbBJYODZKE4nH/qjgDvZZvPGkozO5JYAlERiV34
7HotJwyhMP3DLGsjBXjnwuemkf2DYYUwbwi0usR6hUijIoJ1OMxoGknkpUM8BEGf
uR2XC9pUskZklJ464EbkQcA7lykbiUrz//zNan1o5oAfrBbBRM9YpVSKrEpBfBQv
Vq4cBQeaj9SZcKf4/xesox9cnlS0VIzaIE7NuYV/HV5J1NeyuZpsoejQ+HX/Ka3r
wgNnRH6OLAFVidmdsjCDwDoL35069QxfYaM3n3e/sC6KuEEs0AlIw1cuAAcndFCG
ThTaq/xIfjpWaNFTRDiRP+hCMrXZrv17EjAMwRpBuRHnNJg8nMOcKQJRtwGfCaTL
DDBQrnAgDxi+Pdwc81HqHq1Ij7fWRGX8HCv/n2JBchWPc8KPRPeXuZ9Udvd1jfQC
TxTQXeemqMbyOwsfMYMlK5Z0Yim+zDLvow9zNqh0a68ARjDkxgQxiUyA1q0w4GRj
IJ9WdX4HOgzXzCBUObBi4AeM2uibJ17s71vMcZPkPitrSvPhlUS4w7qtce789bCB
udoJt4KUpG/9qjH5qe4OA7f29fxAWWcuZ30g0bEYiCCG+qzuuNd8RfYocB8MdQIX
XfEElrpH4nrhtHefeHjbiRX6/vqgmHSCaRkaPoIztwFdNVSUSgN6Io9koAoxS3Rx
Psf7JyryUafDGZ4wv5LQVx55+ReTOZxgmHBH2tjLJewxpZUkInvVC4PmWvpNT5s6
FrwgirCbK0bi9ReZLThUDYSdQOSw2b6wVYHq7IYigUJwqWDcFvO3UIgGbOqUSqEO
EC0Y0cY0bcuo4TnTIFOEYc8QGgXtubef94G+9BOMStkMJzbWsDCvoOsddpXEXWSd
Go+KckS4OoYTS/2Xt+QaD0+gOubFnl+oQLZNaciNlUNEHb4r+YnEaWya1a1NU4zN
PbXTlR2acmrxz8mrBmcVC79pTLZQ8eVs9rSlGNTncoHhexMHL5kKpUb6fEya2MvA
013icBZvSGrqhR1fstRmiuE5lmMeNWG0Pz9ljgUl4eCA2ezlsI4Hoy4qwbgOZY1r
yh68LT77+k65B+GUBL5qLofAhm7cr4ME6B2QyBTdCjpzmrDDh0dxjy5xvDtzaBn7
Hx7sfIkOSgO2qDm14ZdmJi5B0Y1G5G3dLsCq64w18s1Pcx5Zk734Ilq/bLxkuT0A
qElMLPnMI1OpxY6IE+gHp8jsU6mWW/f2sQjvtAJTtJ3uhU3oGVLCrXXJ49aeqSCk
I2N60PIu4/W8PXG4lpeQfgW7x9i8SJ3WL5DbKOvIPDRSaojojcJc2xMOzWG4ZZ7S
r3eno1OH8hV/p8ZMLCGx40Ij7hHmTwdlcWcLIDbj0MuO9wosmtpRLO9Ba/Tf338f
LNrIkVCrg1rKMSig41oyji6DZmxTbzggKHuK7NwCMk1L1perJbf1s6fn0rV+LHLT
E42m//I0bUkCsye+1RrtKpWY293L+ZMekP2hQSpbv8qHZqjo1pgGYl6p1bG2EIej
Qgph02OKQ7iLIfkJOEDxwajhofmRiH/if6WYum2/yx+wRD7RF8wrdCO924/Furdv
HMUKt+D9GFOAYQa60RaTCvtMjQnFObyZ8cO8Ir0lul57bD7ZxD1Biij3vzaVz56a
sX6zOrVXTU/Vr24qhcMKaFxB4D3i7RbYliUPheA/b2JCRZvrf4mbI6+1WNEl0P3V
rNfuI7ZvlrqdLMu36gNv1Br+lYNGb3UD8RNQMv7NqXEGxJMbBzfoKPirV1JC5e1b
xcdw9QRMXMt8hgEMNMnKxf3MC8hPSseQQ+j9C2VSIs3iCFdzXf8BeztlERnQXSUa
6ETTlvyPePcU19zPTvph3//3Th9mPcd8kQ0lOQz/+JA2xh0zJO9YtxNK+V7UZqgs
zUv2CGoWEjpoUsDZBVzTSusbipnLoJQ9k1snnkgOFjbQoO9RDA18yaQKPh45TneC
9IxyhvmyFJUkaCgyJMorcLsLqcKV/DHVYwbJwxqqK8gKPuN42QlyzFK4tyvawHEo
Got/BZ/RHFCmcAwWer/UYCOfA7gtmZjV61YB5+pmwH1faqw5Qkk0TZJ7GRZ2Yed3
W85PqY5BJauAXqVuNIELuiScrPTUtq5ryA396szCcRHrIHt8SKv1rBwFtu7hAn8t
SjERDgtZPDm5Fi8jUQ5QClL5znoXiU9tjijeLQrJZ0P0fBtTeFGwV0r9U3XULAT4
52BdW51OK5sDANUp7UqPNh69KvHLo987yWTc/wWmFBgaDF0aRO4nfJ7oetdnPUCc
RaabEOdcpXLdCADYVYP2MiQ06XTSULa+tc6/Abd3RPCI8y9yjznMv+x8Vf9RRLLC
ao6xvvK9KGrYy7Woonq2SgZ19WjCeXihCGiNdPP8XYu6h82cSZ6CpxmyzZAyjfUO
egYYXIDcGfXrk6f4ik4aUWc+GPTSVvk0pgOXVgbYJ/l7UjQi03T0k8EZKxhk7bdk
Hv32SDxenfwkQJUW1Bf4T08T4f5Tbb+wE8PF2BmXDFAI2Ld+YXL/A7m3FX1WVc4Q
gSDZLooCrCzyP/ZQCYfBb7yd5fnwSRbgWDXv3RcUMf2b2Ty/MxVx/YxsQnzxeASs
mlTnPqQ/GX+wU2hnMNByRxeUVwnCrllTllFzrkCXaEnNXTQi5+QpHpK2wG89lTtf
fRjBnSQFWV/R3KuW4nJawOMaztMiBminjB26dYVuwWataokRpcM5zyGBn5Ms95xP
Gq3w92xrS6weGR7AF7qKcDJFMKPo/o/XClDGlDzlkClcvemWtYOXIs8MTeOdgnOL
+BF7AXkezEZ17QTU9cVjAFmRuYwLFyNGUjUkIrcmKa0GwWE0SyJKvE8jHKcjDoy/
J/OFevKUkYoAkO+0H4RJUcQVEyaKzUzAfJp1cXDNel797ACsE8GYCnEFTOk8vEH2
RV3yU9d3t1AKy3hJMpJCvM6CdX9MROvAlN/Ihl3MVn+wpDRk9VU+5ArhxYFHieKn
Qlo/m0tLr1BNYMtnCBMMMkXyxeSsv6nf8R/xSdFwDEMk3kZIEVFLc+OXzIxc9jCE
kJZuNMqO3kWeCmlY2wlN1157ZWw1vTBh+w8S842QEZwn4ntQyQMeGq9dvbgnu4vE
0zlDjVz14nssqPDZrn/Okpt9U0euD0ir0bqy39f4Qt3ggptgnIN/ms2rP7P5TEZC
0zlOHQIPGqROZBZ1DH6k3aydVEe0NIYTCQYMMnohoNFSZcWHvHdwu9u3Om061Wyi
zCHcAVhsPMw13QUnAyOUhjSu9JDqyiLVkwIvN4Gx/PVYKZsnRJkgS8LIU6m0ylZB
vj6NCBQfRbO2rvD7ZcHYZIWm/ig+kmvYQjY/S5ZxEN5Sxfd96x4UrIdu0h8X74qE
s/L5r7CFLD109lI3bMVLxy94ig2iXQF5dzLDCTS+mQ1qTBSKgmAGtQLLiVHvGqIc
ySOslRHMWoxT67RCzq5h6zbU6yEZbEBvA/uB/NkhVcF+Xc0mGLDHu66TplxzgczB
6hzY2gvcPzJt4Cvq9D6BhjDsB0BZn1Od8t7DgiAPKmoFtSIeWVv4Pt9AS1+sOUQy
30NRyNbHPowyNHERbzOoT5lFrzdDQJ63mZD3e0swrudC6PsyyCap6yr43L0fTi/f
iDFdneCOPzNhO712TiTEhaDu0PEU0x72n7b4fS9hsf2XUyDgI2CxeFtY2lLJ3d5R
0pk55mObgbnKuysEmaPsltXL1P8Sb3bgZDl8H+VQenXz2QJfkQhmSbdM6r2FDVuw
pQnSaqBe/VxWXsuld6NmsmVuVI1s+AUTjObiiMK/5KhIv5+cnWjGBPYPK3Y2QNFo
NL3OAsNFwCZMAKudcOgN2L58rElwG0j5ARm2TG+16uSNklY6QdCp4HiEPexdyiYk
PZm2zEG37LlJFf9WlzmLrOEzquxsGPF5RS2s5SVR2y7Euh9DUnSn/SwDb0OmYycz
mRINDZaoCnGE1l1Bd5U1EzwZx+AMbo+M5lhBfFVtDSmx13vcJvgY/SvtLNcHeMh9
zrJA1haieYnAQ3fCPbGm3R90sfbdqXvtU3ko6eDtopdFT74NECEMr80xrNxz42HA
QDRYtjg86qvzWUMHqiTGX5iWw8yxIhjrHzOKgsXHbQyjUphnc8KI0An2uQ+82ATo
NsWbpFe1NAumPSAHX6mPK4rsAwulmKlDhz/LshUoURWlNyviSEiHqRTOHlIVnyuS
J+ZHp9DBpnNPFTRxujxAsJY+CwrK1owoRsk0eUAc13ya18kLIDa2qBvD7zvsqJjj
w4PonfeUVd65jZ5GK/QHRROd/mbOM7zmG1OVTit++gtZ6koaJ/kYHvAFrn+OCz3h
4GVf8ZfY/HG6/HFGe5rqvarKZXDRdnxR8I3c/XH+NfHoh3B2LpDjIJ1mq7uH+DVu
HFhwqOTG9JpXumm/igedB2QHoKkF9cZO9HC/oe/QNB12NI5PFIvHtJMpY5l/XRT1
wkONHRbEGbWPqycfsthJ9R8V1y4TV4Yc3uGNKA8512EeYT4svNiKha+B8mKBTcBn
UGbYTu/0zeeaqvG5ayxWY+00X5Ku7Ar7h17C92zRAaEa+K18GO6AWwx+zrec7F4v
nKYdEm6+wMIGs3GyBwFfFwmjbLczDJZS02OP/DDXZB3S96JbPSGzWkIp/6/crpMH
crvn0prIorNOLDv94jVDcJQoNAed1aORF+oB8we7EAmylKYh2SOaSFPLYzRRw2On
BLdOZO559zoama3nCxKVv1Z8i5iiX1GLBK2k+bfqQFYVzk2NGHMyBFyyKjkQxC0D
ecn2Qd0otMqIkj3mKvjQ+m2E/C6FANOeHI+XbyJEPJD1MQ2vjxxsd3RRCDdvg/zp
tl2g0DeUej+S553Kk1LU8/au1uXPEemXFp3z1lWcEwcUjXA+k9qDtEiSkwDjbUXI
vZCuYRC0I4uEE8KE3crI29M3Bq6CNdC2jOpycw4wYQxtkApojhTEvlVoX4cBkwfX
RzUjNKSouiVWaaSIcZ31/RjaJpnHdm4bO/TcYn3apoxm5B+RpaGHEnrRD0Q6CDfD
G1+vB1bTrcxUBkOo3Gzz44+Am/gVDIJhNZRAU6kLpEKfwJRTKbNLYj+selSTclqy
WLGnPddT4j1qhws2zyQms17YnS6haCp32SaxmDsEumdonRsLQinNMHdZCG3myxe4
J3R+UzcEC0laAzmY/Y4KyCKp3hNvttS8pces3BSpN+gLHyneQtP3zBzsEiTgB3++
VtWpexTAkkvSuFYhXQ6ZkhAGU6UNctzZQ/uxbnrDTSPqjkFIq5FLsb4USCE7KVPi
QYLs7VwvIpE389XTXcGyQqxtyLAtYLGe5Pl94lnmO3HMzytN7i3N5Y6CO4JdMoFj
EHpi9eOoK+NWE9laEdFvsKN5fZVWJDqZxzQLN6CfgIpL7bzK4csTyBmorY5HuXMU
ae6AYCrC3MkLbRBbC0VHSqA7cGyhBPzUfL03yKobOL5/YYbQ3sbTStSnZx5x0Dkc
ZwDDm1HB+oSJNJfcUt2BH0R38gQdqhW5A/3QV//wuy7vgZhaIHkDKlpLX8K4wHMs
Ig6MUy3RVefDf9L7IfZtBHU9XoaPQmiw7pnwqIw+Sl4znX5R3Vdl6ftwlj1/2qCw
qMxoHxCY3Hcr2suBvfG68LlDsstlOWfUrgt7oONkOPIVLcGZdV1m+ZxqgnEQLX40
bYM5pxzs54P1C5C2BTtYofkSUgH/CpnrHFGBKIDlXMdNQUGy4srp85NdTXS/8lGx
+lCFMpLq5E1xSdW8gG+sQtZZzhorVL1xNbmY6vP32oC5X/Wv6cUNokouz9/MLCU0
MSGXTRkmntzTdms0gEdXUQlD4HRlIkw3+80FqfL+cQvlvF8NBN7mvoUSAz+eCP3x
swgs5kEhnHB8X0qAlvwPnvTSVQZMKqbokAM8FFv1trR974dHJ5H0n8GrLR2pmhU/
7VqJqQLzhizHqMznBSqdfp0ohPYvUtFRdHoB6K14ceWxZ140uV2xfJVchw+fnT2B
bKtgm/S1JlYmIR6ZJfw0ikBFXTP2gHFN6mM7cDmTZOReS9wLr11ofcPgb+9vC3dG
kf65CTqTvElczZ4FXUdNoRAKpOqN95hy7xPr6l8qT2ZpHvz+jKbXwTKrAoZfGGNm
isvTN+3iMj/xB+M5M6wW10J0lXskyBxoEWWd4og23KhU3az7EKclkD4V20tHNAiB
Z9YAedoxwJ5OSErVKuNPg8Ae57Kgu01yrN/Xjl8FHE2z2xhPLZkjDmvW3gFIpeaW
HcJrlWetRcNo1hcMuki7LPro6pjRQp3pSrKLm3WF8tpFLBTcrlpfBv7dPdHFvYAd
Lp2EWRdZQ6pijr/gi9iJhdPHHdu6iFeNJR+U5M0f+5HJCLSAzUpp3ahHVZRAawI7
JMv70TPTqWvinTOJESFt8j3wxwM5ut8VfAz/8h2Ox/uHnkqWNNsm4zbU+rnDbPFH
S3eKaD6lW0YCQAaSi1Bz8Fy6V+a7Se63Q/wDrFTkZjDzccX0816wbae40J2TD7+S
AXpsiR8SxjlPFV8H0gVgRr0QI4psBgOQ3dh9DoRFkWvQ2G1CzvI1UqlojUOfSN8K
PMI6bA5/JqKrsNcY+Ot35n46Hv2u4MNZURnc6NyphtGrf2wrC3WV7MwxXtUxp+fp
EpevGFlH5AvopZ4V5A791ctcTSa0XH80BUSOHPL2EOO7eykL8iDLM6pQT2nQGjo9
Nvuq6y39RRBk5FWuFifesslkRJrftbbfhmDUy3havc9mGQFvewdrM7ZCP3gGdR2A
J3HxMyAGLfdR0naD1GPjiiJgGi/gUabKU3pRwFZo9awbQRQE8Yse3T19qnm3poDz
yrqaK62B49Le+HQKb/k+Bq5/eoCj+7pSDB5GAdiWW1tLbfNFYmcvGFMnsC8XtdTN
M7dATpQ+SdoCfqwPQo/Y9yf29G8oPC+LUBzKnag3DN92i1ox7Kq24XeSp/gjVQk4
NP2upii1o5zz0bCo969RgCEbZDH8tZ+zajEELTIHQYWM3T2Cb4g6r34Cs3sTMr4D
swDiWZxII3ZLBiHetBzuYFRDsqafFNNdLT2Yu2q/TqzAGd5zGR0+5lu1swwRAw2m
00dBRYJ7KJCpkTh+pAZknNLrCidpMCI1LOpy09GSDW5G1XDSp0CXdW67yL5bZkNa
rMjkUb3r1YWnMi4I22CUqW2Sh+r1A8D8XFQl6pEW02oRnOMt1AuU3NSz+iKKGgf8
XswpPWXf1JR1ruXgj0IQBuTEHOifrs4DgwzeNUWhovVvet/d6B6v4kzwFENrJ5xO
PafK8x4CWrdUq2vPwqoxsMAEyjON4tHF326qy1FbkOoISBgQw0CaXGVUcjgktzYn
k/V70ZrJwSBQWO7BfoIJ9G9kDsjxWOnnYgunHANkEWG1QiI0bU2EvkuUtP0i3Gt5
SuF7fS25lXC5NdsVGIhYAd+idV57VucsJEngN2VCKUQM6lj41yAQp+KZWHdNuNLG
rJDQO8ul+U/fVxDYLuRObGI7DsWVa2+nI6KDt3ZsGyMnqL0TQJQMeXXi5IjhVtnT
7xbzRfGCZBotDZxijlYcqCxSv++0M+JExUW0mIEPVePCBK3BLxEj9EnaCLJS/ELm
FVYnVGNkNqPGlTciUVYA4/2Hpifc4JQ6Xojmu+X3twLlQKYwBX4VA6ACgo/WGOra
5HaUoc0gjVQnyli97D999wG8x5ABirttcmVg6A1tPflLamFdtV9rcJsMo4jP981C
2FLyfRPi/+6F8DmNM8Vk0PbBIUuo47eMDQbAjq5Mx9b4hG8zuAdsVIDzVVzETbN+
+5uR+KFuH6CStOlV3MxVM/tgbJCJhA7CGAQfRjWujyOvFtYf/QTu2/hP2YDf2e7z
mZ08Wqznw3Y8C1tDth1NN3k4qP3GBjBqSyX/3LJbtdgmRf93Akp5mJ07pNdDqyni
E37Fy4vj2Lth6tkgY791oGpOSnEkqB5KhFoMC4RQZ+JbJzPYGypQvu6LS8H8mFQC
Zk6hzlwNr8CiNbZkeqXjz/daKotTsO9EjMWMuYV4H23yTvxG48yLGXfZ1WtGWrVK
1taLpgs+sxRvIqK+48qIlGRbZ+KcA3d5Ohoa61juqQNGsu7WEVk6ssr35zxy6IFx
MmnnjancbfJWCZMDZHqxJSFJJx4jwKp3kKoHrEt+BSWorenY50vGWSYqd0oVnt6x
azDzFknuAjGnvGP4y3B820Z3y/5NaR7JPSEsll7NuuOzNGROvrezf7gRrdXXSlhV
5NlTY7bU3Tzc88074W+DwKOIQxoy0dHBGyciqxwnza28gH+U0M/o5QJtTIWCT7TC
o7khfZcVip5tyPs4l9R91aUll0jWprWIqgxD+ztwVZaIikz2Jm6MUExhHlxD77Nz
HbQmM0wlnMJZ1NoVkT7Mr7DuxI6T662Pq3SDcetw9qIZdkuUaN32KneJHRJAdbms
2J9gOyVnez8nuEQFcDy+fIwb6O4kGXiUulvp3e/98rrcJe5DdlclzzUAqpxmBpl3
UJ4V+137VcWxFRGUMCR/W+prxZ566OyM83KPHnKLFZ1wkwe/3egMgbf+ZX0vWBwO
WLVlGB8oIgUMNrKOZsP40ucxluTqR4IKvfZ37DdackiHHjGdtngkDg1AgfVYWsdP
sNzv+yCVEg/w/zOE+G0i412klaauf6MrxBNmiiLxB3TDKwfMv9wNsPJZ+d9JcmGP
a8P2nah34OXWn7v8VPVe2IUL8K5imWk4Vlvn94o34VeZzbc308UWrz/A4grYjgdR
uEyVRNaOJDU9qWIH+pxA8cfknfrbSGKmDD9oCuyD64LKBACOUsUBddHgOseuxPo4
1VZ2WSOyNB+or/v9eX82zWrFLl+SfG4KgIDcOKAKrm73f/ZkU5P8Oa1yZWK1eaNM
OFhzyoBpA01uYd+NsUwpd6GsaUDGd59UjYN0yN32WAaT2ZQXXYe2LQo00/3WU+j4
5j5ZoGp4YDt3GO1GQXi9jqGnBYAQ+sObKv5nCL5ElxXA9n/U/6yZnL//W2LA4csb
nIrrdynKG3H80igFfO7UTD0Zq4uXCvzSwcMgkxEbcMlrTUqZkzRs1skrh8tY3Iyc
VRqgFhY4JY5NH52x5AhFpxji8l87SZyF36ek0JkxoJj971UCWxjKGxbrZ7VzB+8B
eMNbc2Ykrhcl8OV7OhbmxeCyXlUD2iTMk0nMKW5OZP2fl1WcuJPgzDJ05XXnzYhn
35TDt51idoJswkX7fYXN89t/4b19Bbfdaz6oWMEWkmokivpHAPjWr1OUc5UXmQGc
6PcKRFGOqj4XGEcElHyY8niM3kDUQziIhaa/LZ1aoKNfe6TuWRXdnZBoxJtJN6jk
wtLEeyRKOUzGR0GSRYlKCksh3Bmq4+w7KDCEzyyWxz+SLruIlQ9d5ONYwfK1pcKi
WpLj8ZaRqMsPEt1Qq7YzC/LuNRghV0Pc6nYuGt947kkOcGDLqMAS6tv06ft5bwqW
WIrrjVFBfliqzPPCMkw7X4JiWoyW8JQwllxUhm270bfpsjOHTJGJu80hSS/B8f4y
QFf7qx0lLxkhZxuC8MsG+G656AFEFaZp5zErfFy/d5NWL4j7ObjEar62l0HlIu+W
Zv0ASxiiLsLcPle9sKLs5OqD6cXs+OPgrbddrxgUhskXNIbvXzjs3qaYGeIvzfdh
EcMmAdGhFHEUkKGbyETHkdlBgEvLQVFyeRUtUwihkEbTuD+xCPkV6ezV5azxASrv
yXjqruXnq0HRXQ/rALqizjF+loZ4UUmkwhQCHDQKDZGtuuZazPEWNEGeO0uyHbzq
uJsQ4jS8QEsKfwQGwfvO9LCZURevyBm5de6WEXCcmL0T7cJsgv168lj6qQ+EOfsc
UdxyKKWY6jB3zCoDThfFUf4oO9UiWtJyDcBPritiLYnTUe8nruWkOFFn47TLlO3E
4hJl1PW6vZSkJKO3H/AIBqTbasz2AVqmdE7qra8dRzImmIHfvY0XHmJeP4e36FHT
6/uj1Xyp3D9eg8nb9ReBCykjxKJhbNzST1+ckc2cJFLWq0IV23YBh/ubC2A4Q13e
c5I1JvnX30iOB1mosRdyw+vZD3wtKkUrqAqq6Y6gsWjpSksZOycsCHApMV8kyGWb
8xqYu7HUEk0q+niaGxR/Kyno+ZjcCMcsiEl8g/uL0lREFHDsZ+EdjaNsAFYR09aS
jltshuPw5qOCB/KYGtKTCB5trjznVvJ+9QazPqdbmtqp8aZp8BngCdkhlfY9tskR
EdKdogGH/47JHh9c0UIUllxqt/gxfDL5Y4Q4YCdqH93RwQRFKYQImusHue9IJ0TE
OqZq9YhnB8IpkbYVMJjNapdZdC5tVhHeZ0RjmCUQZi72ksrTn9bakvfpqcQvPPYS
9DVmX8hVbbttR6pRent2VBnM3DJhFbePE/GFik5IqdKhsI8JzwRmWWHHjk6zsBl8
u4mLqXFWwuDHOUG88jm0MYKQd2+hgN8+tRTYqHqFbdhyKcqF71QodzXMpBEb8yed
PkwOtnuzAq5o2o7doL5nsMg8o9pVgJFbhd7PK7VAIzhWLDTvrgnNd/FLZV3kEL/J
Yd2L2MW7+mkafhONbjd5BJGkPZo71lredQmRGb8eJ4CgxkwEUkH1TyAuWv2vuENT
QmHqrYI9ZPomn2r/TME6PCxA1s7mmwDhcL9LsUxClJzJRV+T2Bgw/Ci05v9Cqej+
Nwxf/jUKyH4FB3/fTz10bc1CeIisuEfIDdwEFmsnoeceIODeYQtiy+uju8mLSFOy
wvyxZaCP7J0bfc+5ahNjJZJTkHs88YaMbyLj6gB0yiy6/rtacIb55bSvc3cSD+gX
jQFAvyYXCn2ECJufzWyuqeboxWwhn2cBoxC/vmE2q72/Wudoy81wcYdrRET+Ym7z
CIUOrcty+FYKUw75/geonvm3T9HkXphxZeh4RrV1n1MNjSqK17BVP0TLkPmhYkRd
Y9P8w1sarsOMZqTKDFi5N8T0VHiU9N17wr1GBwEpNUnZ8Vnhv3NI402MxsFm4m7U
iSbzGTZq7hOFNn8D8n/jltuIM9tmGlampBO/h9d9SeacuFen7eB8tdQ2rlSGXhQG
rE2V10xBh4QVUdwBBQFiy5SQ4twA3/KPGuw7Ytsfc6q1aktxz1EdrIgcArlFsp5P
jukx/mb6mQ4vIlr7lnoVcnZOrPSdKgBGE61ID/PWoxxJrZjRhxiaUnwF8i1H8XwB
BrbJQvR82ETXe8B59b41g8GMNuoToU8CPZ1GIVThqZ8IJaCcxG6Mh0u3FAF4iuPO
S4l45/gSMdt30qqDy0dnZU2AjSZPY1kWZ/1dIJV9obywY7lEaRhw4StLvzRdYZ/v
E13tsDBENxJQ8U9gBN/nPKAzXjBV60/St6DXoWZE/9ptQHZWtfHj/6sbXZOqSu6p
ik524EPbWnjyuRz22a1Enxo0J6eVUBuRPX3YMJITmF9oYz9BqKdYxv1dJrHOVwyY
Mx8PpVgHz2YC3c2v8AfPq+HDMTPikeslnae+21Hj1M6EymQnIAV8bTdteCe292M6
jxY3nu9AoGPeyVdpvKubF14bmiJfMMdTHJsN+BdjwkRaEf0VH3brEGb+zqpmpWqY
CV4AUw70I4MPAs4haVXWwSGONS5WB7iqvC597UhwWDwjSWl8BmDGekuDxBpwNczU
TCUZAdHzRkLZJm4ZKlCQIdCGX3LZa3qYYliiMLr/HM/qcG4QmtncrPmHciKm0A9z
L+5dy2uOtMgELGSB+v/uLLyhTvYm4lbmR4sUdD5kMO2KmSUlGGFjUQsRGIlXSeYA
PwCulXDoSeVupAKSDaL9Vu8Bx0XpA0tjCBMuOcMXplS8d4r9v84MugM7rp8yWbnO
uGYRz72nVOt68cauXDyGTnAnVmjyH074NwDQaKsiXbwcu0AkuoQJ1ncalRA6Eljr
T6lDGAoIzj79N3UfFoXqzqYCz/aqvTvcuMEgVG8AslAE3ePxg61CXFEmOvU8VLru
5Y/wBksj//1Q7+9ZqXWtygG84AcPCSEqtOH3ayIjTdGbtkFCokgKExYY2Y1OrS6I
Ae0oKqPbGzRiQ54gx2fSq/nI4m2eQyHIZZyYxHgWJUFO0Ln6ZGIabt9ef45UFuQQ
XKY0wTsb+Rjt/V8QDMS6C/l4uDavgJIPU3QQLd41hImYV2+9utswxYvQG4FdBxgG
iZ5YVKXjT+H4IBKTUEiYFftwWOpoPnTgjJBrFXYzeD4GZb1xyNmT+Q2Yg+tw6OS3
q3JTSMglVD7S6ZulUp0dVApOAl9vLwLDj3BoyUS4B7CjO/7PojeSxXB/6gzramkf
EezUipKJVec+TE/7fhq+7A==
`protect END_PROTECTED
