`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHzFWMI+vDV1r7dUky+TRyHk3aU60ps1mnPpK5ebciTU2EZhfTch87fmGYLrDf9L
0pZU7lQD2cZ2bFe9BPsPjXmtarxQGw58ZLpUMRj5pqcLBO+f6tdEw/hJ+gW3WNFu
HYb3oxEylpBb9ZaoFlZTyteGa9Bq+gX+bbxX1+a3GbigJa8KM1sOc/O7c6SSgjUm
t9NYJVAH9SZgCj4IYPwNJ+EJugZCeXUDMt3moM09L4IGefi0tTHmASTWZtDliNhK
m6QW2MLVAjD1H2VhAyo2PCk8fl/8lyrUp0J/r7Fwry3bOHTQ8UbbvU/mqU3KFVbq
cJeLaU+W0FVbJrhSdk4PB3dxhGNnD4pcqaZVCec1VLPEqok4JmFR+lnyWblqlB9q
sSSZbLuI3YGvra/jtbo+nLtnifmAaYJvbg21sDI8+CmLwtkGvSGl00TY1tHg97Nu
IaZLpd5YTWN/rQCgPb7g8a7T54nKLj4GCRdfSgz/cMdK7sQ+tVanbe5/m03fym4u
yi497XWnCNjFBfUaMFFWaNv8XqGYjezgTS0q7XO5YCYqI1IkHBh3FHkLLnNZKadq
CcFWcKak04zAEtxmUJZT6ZAcqOVh8wdz4/u/gL9FN7MK1PG6XeDldBOFz/lyTHih
AJHm5nXzJ3XkfJM2aNa+VyQBNsS+v4mN8vKpmqqYZoU4Uk7TaJqTXD+2Bz2kzRxf
nORchtbErM+xlPMDGuaBonYMLxPXvEdhWsSE/7CRPJorJeU/MSUxP5tVM0TmWUw5
mBqUVrGM7uBnTg3EPacyKSHrlpIBcnnRRQfejyF4HKwVCoaHnVbmgBNVxVjRujcL
GgDp7AXkkyrzdnGrMdx2DxEtfbIUsYe1JIg9yKlKv3pS6JBCEp7pOg9TmUgokhJY
7qSp4XEEa5LN+kt5BhuUz+Os3QLalQBAkz9krePFzTWTzAo84f+CobQOHn1xKg/q
nZnsk5I5ywQ3mDCSPjHe+zLpK3IjFNKILmIpoGb/AxoAtvywBoC+hjUXEDNv85rH
NHSECBciYnxBlEsvGl/L1XUht1IsvkEG5PlMNo4h4BRDlfF6CkhKp/j9pP/JnLDp
EtJB2P5qpasb4isT/PcbGysHX6yS0CDbAs5K4D/a2KjPr//al2lvnO/pK9/j9K3X
Og4ZE2mGb5mheGljStwqkciP2T6v7R0rm+xHN8eSjESh2WtWtsrYmSCeVgjUFMz7
QOFLH6Wuyd7dAgiCp9OFJa/op9jiLLnWtvNd7ykkcYt141NpzSSn3+yu6MeTEQOG
I4YH9/NdBj3Krqm8Uaxi1gMwbGFuvT5m6OkbjM2402z3zIkz+drALqw3MsovA62W
kuvUwMBWIijTxOw5O47z2G4y4VVoPn4GTspxzLuPzkOCXCerSG6e2IUGbt/B2O4K
RmW0PVkeIJcQgAzT7X9YU878TxgGpMM5aL/w4xi496RJqzYZN8/1Sy+SByT1ho0i
f96vs2/GQZzt7mSqz7xeKKip/UK7ed/CEoeIJpZPuWhZMzsaSN3C2gcNp3p6pyRo
OaXXfX2Z/ilVLydIjBv6xflyBrJp/s6Hwg8YVV9ARmuTVf3JcpISpIMMh2jdSMBm
3BgQjBhIc7a1dc656Q7VZxQs9QspVlpzKYNQrkW32SyrDwUqowu1Uh1obD5m9L9N
HofscfVneFBA9Mxc6aQFAoV/pXMTU6L662+/jSz6edVyZ3Nb77WwaZ2NzhF+8Wda
JKdgZqR98tg49XbCSM1l56NWcWi6T+9CAhbuIrEivOHkWYnlElcAI6Jjk+pdqypx
a66/KA4gKOadBqARzzqPE0zsGy1oj8AJVJbCmATEP/QVexL7IkB39wiizT3R27Dl
6442IiPUxhJNXJuc8OyyrbSymmElWvapZHEJiKMn7Dq4saxd5jaJWYukoB/+oGat
Orsui1Ku53y+Mf5F0+nYo9orrkWAA4R/MVH6njYgnLqCSuJMmH2303hd+Mvp5PtC
r3+zO/ugurf8xUtfVqCGAUOUKzTa27AdyeRlCwq/ZVqvH44sgVhklWZtjhp7WvvN
q7G1lHDEgt7z5elp85Mgq19W1jaepv8Q/FL5j8K/A0fuLU6QKvPjA37TdfcYeDG6
tFDwPhS7I9dTmWGh0wxj1pEm3548bvSltCLAoPTbM+KrNcSL953Manv/qTZSAm11
80FzG4Scag9NnFFEkE9yn/TSG7/UNotMJvVjy23JRENZcgEqPpmXNRorToXZlixo
5E2E/PSzMMW1OpSE44c+0HD4ZytZ67vTs6gzm4PNgnsZFtUlxRNi3KY9fzZtCIxH
dwm7a69bSfsXNePkzjBbXH9g4NNKn8ONReYBxsDvRHHlvp4Zef/M0e09u1x7osm2
AaUiDw6KzhJI42kAjdFPkUkQ/iVLdaY4z8GrDNWru2wAxtbNWQkYqpm6/KFBxU6A
NM4caVOYNa/iIVTlgFY7buH+vDqj0S/M8Npx2JF6CXOybXj2o9zcP1TNQ8LdOviJ
QVbzzSBhh4DUEQ4TI01JX0n5ZkLlstQVQ2/ujyFIret65cHyYEf3HmmCkF1TiY7n
FoFRAmr9tv4Qaf4z2bbKRRCLjLM1+Psj6N6yAqUecRkoXe8lJx/Jao3hcJ5KAlsq
Lf0IYTndI9Zds1nfOQQUWHL92rKvIASb5Eti2m1ffBkjwfWM5llYDl2j1I8QRTJ2
zzW5rV8WHJv/qs5w2OqphtnQ8AdYtk+ar2ULTO1uKcMC60+CQLpveK2LqXxXm+Cv
rRzhu8EVXzoE7bCy+nhLvRMrxofFIdliy5vllILiSUSBpJ+dJMGBGYOfO31jmBvA
toWwnRz/AnT44fVTj0O1V1lLovzKDk3v1pKZs/OYYx3qf3Mi/NiUHSXYOb+v82FI
IA/Bwo2HJ9KSCGb1bDVOT2xLworesSlIldbFLpV0gIvSMc1/QYX2gLZbqTB/KnN8
tAofRD4Cqj8kxdGKWvjQD7/8SFv4RMX8EU6mKdNRzOv3gI15DM3SUmrGVeMycZtv
zBdNKK3BtgnNWhjX6hkGXhVQ9m4t7NclPC9JUVYupBw=
`protect END_PROTECTED
