`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q54pH4AIO+Cy7uv5zRyj6t3mrFL//A0TaAszVum1VrNFkAJJKO8UgkfHRHFyI0ZA
2XBLcAbdyTbk/unFg7AQKKb4dlRb2iSdanp1+yHcTBc9KVmn/KjQtA0E8+tL84VV
qf1mBGolRIT24O9M6iafV24H9md+RMvs7g6P+tJeKDcWWF0+QtauB0I12JLDFbyx
uugULnroPxGJQiJODho9qwx3YhJpXc5+wT5liK48NEeo7/I2Vggrvi0pM2KQ4XUO
JoKEPiUOi8V6+P0ml0HXL1jGXvh0J+M+0KDko/17l81og6HpYvmqiRWXnJwofaSH
rlB5lA1pAofzuCkMICa4DHlCR576gCCvAftYW9ww+NItyM+Q122KoxgKOKvnE3CH
b3XW3Nblim3lMw/5/wga9BdIZNY3JDHJQg9xdEkPhqkeDND3wz5hnlgaAmhmG02/
KV5lbGp7OwpnQz7DVCKz44vCD1LPB4TsxSnfgl7LBzbfHcNj16bw5QNV1wI+oe9c
lYZnLEWQPQnZ/7/jQrGLtA==
`protect END_PROTECTED
