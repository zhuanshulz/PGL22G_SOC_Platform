`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oP9b/zF1XBnwmdz/b592kKdYEEIoKATa6293GmvPKzyFoONbdlvKQ/BAZN3Ob9up
Dx79STFf49aUlw35SmXF1Gb1qMu5aRiANAkl4d9vOtFg8KEnC8p3e3yrfMv6hYI9
6kqSgtRyJW+0n+hQgmpkauGafwPPo/EqgbRL39lnLiEwirpDBxgx7I6AkF22K6Ny
y9nBaO7xAGsoXFYkouufpvczNjAYyPanZTq2Dao4r054BD88FiEAp0V7ohU/8cv2
XMcAnbr5K6HUZl8EqAXH8v7w02yNpsbDUa3Jr6ZoSzibkuOB82kahsBkFOSK6vSA
5q9V5ZiG8HRb1/LNW1mcbMvRh92k5cXnmCKCKL3XpnzkUCtF1MfZAE2wEn5kZaML
TD2i0JT6CEAQkPyaCBxAC7rqqmsQ3ceW/pArgjeHPmdgwDvEEyVL+kVzajzBIOfG
fhfueeBYG5TN09VkPspN3fnGSab9lfCRvNxilTP4aIbEcj/FVJugqRRwKL02hDPw
dAK4rXzK19tz1DB7kqWD4JXK9oEuUOibW3lwO6HEmTKDSR5FDuIfLKBDYyM6udgj
sJjmfBTFVdKeXBriDTK0k9qWhncDTYTBI5002JBKlwEBfNQ9A7QohxaUXn1Up9Cw
lBk468GvAXkHWoGxZgiH2GfjvTJvHfm/17r1KqACCMxca7bdx36JpQBMITcjSVvR
3NSIVuaKp3dGSEZ5jzJB0nIrGtr/Gs27DQCKF1Ek9KUDqTjHv5BSUZfZ3UqQKCHW
nk13uksyTkgdA6+mR2Y/WlV1QUxmIIuYSdIfsM6tX5m3y84hhX6hnbOlUMcbUZYZ
/sh0/0D6vZqRlEra5n86jA==
`protect END_PROTECTED
