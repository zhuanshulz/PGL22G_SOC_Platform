`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DfNjULR/dqwNntbmdEwqMPLRPj4MyKZ5+JwJ+dOvrFA+xQQeFBQ5sRh63/w1aZZk
QMoxBm+aLWpDSAeMdbKgE2rnhZCNOelyWwskevEwvcSjkzPWEcM065hoHED3oN9e
FaewO+VhAt8sjyYPtx5STtTD2qbVHtctI+2iPVRaxPs3uU97EfFp7nS/A454hyjA
6TtAxPG7WvZaZFSLOy1pT1zF/fABPS/NAxbIo4W2dZuwaxhciH+cOMm6jP+rbLR9
hFp1CshAhHc0wZrG6/nnsgjKdW+fSocNBcrylXJ5VhQru2HkC8taYcAQPmN27bE4
WBSH8eS45203vxCERqWFRmUNEWaUh2l7T07uwh16Fy4xjudGZAjVynUm37LGHAWi
ryV13sGBP1+uk24pw+/vMz+MZWstJvPXxM0evBub8jmBAgv/7f2hrV03SyKkPLJy
AF+5+HuwRsCnODv5hiIE7fBzYWwZmnfDofyhQEYrHgycckyDufxI+RXXNBqaZnch
Hfnx1Wnz57zjFLhhoIc6b6ECvcch0XZqSJ4S76sS9KhzG3R4bSoq55JAmyni0to1
mfg3C9aXRzPTNzlF8NAcM6VkquKP6e9e3nJkvgq1ZaZPUsXLeoSS33a1vz5KLkU4
EIzm1IbWzs5tmDDbmxn55e0Ogf1v/8MfPQ9/2v78maaVW65tqEHwJKz2gS2Raqz3
VF3UWuFqzLHzVBCU6rNIVaK2a2j5cPBoLpIPhqvBMj7c7t0veved0o0dsNTP2smb
93XQ/V/hUby8HnFQT4JYZt7/5nN+u6T2UWDfdjBXXmQhvnsfda0zPDIpYPXg8IrL
iPFJgS5e5KAtaR+4usnsEVqKub3O2iPBDt43EULLrZl8Oo9bQuNHjFzDcMBGwFuN
DXPXUbleiCHFIXRDVumzIsKnbKu8OSyzEleWQ0g6/q7q/UiajynYGjk+waYn0a0Q
FCuhg97quUG7zjpguiQhmJ9Nn3F59oCPwJlVlz/UZ7ZOSZYn/FE2Q0nuOIIQb1El
0on8zeWxBG/eOz5ufuEwbekGdRcGsUTceKFpPJIChCaM6v0/nGTHsdD1MMIwE1Wa
m9+TqjuOdWQ983XwHjtakYjl2ZgwiIL3aGicSX3OhmtDRde5XmFIMn+YkrwumHqL
2uU2pBGpoRirT3T1iQbnZ6GayUOjRjYNSFwkznYTOlJSAWkDmInSVypZg8RI1opw
G7e4WW8P+B7j6wi9zSnCQPNcmPIKu46XGQt4gswpm18lGXOiSYkk+NLRMfs2LImk
VFTgGdgwsZpGAX0yKb1XYF6Dui1gyslIbB7L2SDxqIRyJ4ijAWGSEF8jXdwL3U30
8vsRLT08IaaVo5H29DKkOylqofgPltryx5PrTDSX80uO9RJBRzzLuLVI17QIimbC
1HcAG+B84Xpz0LXPOl/TRXwp4l2txjgt+qiyvYV5J2E3Nh8FXFGl5DhbsKDUm/Bv
IkZbYA3X0MlMndh5D+Do54WZZsTmI9wMX8njXcGLK0wRQAeLRRpjH1Kea314/frw
WUG/SMz+fKU5ZPU+bEKFUKhlJT0SEoyaWTid47n4XNZ7w/7CvghmK1/A7fxRQGNf
FOh1aJ60BAoWknhoY3+Wcrmq5GFNNRmnii0CeU8mqAzGa0tMQN6+ME+MZuyKdGA4
KYKwtnoJ08uZTHiXPOEV4Fih2pnTW4dn6vfmGDSSHNPifgg3UIxpgx8/x7mgZQOS
TkcfpYWSUQAV5Ib48ovc/4ZMrI/+0NJLZZ/9XtOwLfnlv7/FFN9tR1w1BUK1Yfkw
1Rozr3CISimkAqjhCR3Z3rATusy0cMTk/TEpyTGFk+siwQThoORwFbw7/CQ3NMyd
8mFmFWtTJa5bU511fNfbIfhAGBbMMkuEmxNWx+5KktQII3ixsC1sZZ5t1MY53nIk
qrLo0/WGS4jp4xGI/3P1NVafkGLnWmrArFMwwm7rGENsfpwi40HdxyMIZxX4KYWK
oPETazzYfeApkFwD9Q+yaGmrbeHXitC5IM7gkFt0m72vJS7SzbDwytsYBVRKLY3N
IPdnrSYZizYImnkMb9u4bYw8OfB1U1r+SYMjO/kaHIZl54pvTk9hBdnISUh8hoBr
LtB0ULYOuwRayx2KR4kz4l1lTukaUwqcVC+qwJzre/xu1BrQggrWgON+avsdwEKk
WlYzdq9kFXctx90e6OnABWNsrhaJHhZQeJPKO+ysodAo3GSXAhu18Qjq93sOnwvH
KvD4go8TsvFMuqeP7nZYEeJ6m9vBb3esbOy9H8BQCtjycD2TuepQD1CKXBF3kHau
+9JrJ/I5Y6mSrVb5RnjPex7CPk3Z9Si2SoocixIW7UTQiwtUbO6NjDzyr+w6GM87
cWecEkpzGqCGN9vowKRg3YEVdW3FgSHLX9JResxxVuEoyzBGYgXGGBwLx3XzEUYR
fa8PispRRirkGL3kUAR0lU/1r7aBgdiibRQlAVxEUXDR7fH0Qr7QviFcCd0zbOsZ
6piUsWXIRKTJsY8Tqx9BNVz4od0NwpLn2kzVcl3IpSekjPYhLd6gJ7BAuuafoyZf
21wisR7UU3ZkcnPyg+LuutmHVQvRgpJNrsTyMqDPmvdSMrEs3SJIuodyZ8/F1p4T
X5+SAI7GKk1tUSSWuZnJpKRpw1aBlUaxU+gkwfurunjq646N+lbkig3LgMlFw6ch
RPBvzVsw2zzheSH8YDeRERpheI+IlA8WZUV8o/8b3cY54HKcckSzvjjhIKOvjvnZ
VFYl7BU3t0NzZf+zF9lsieHCxphEirUkigJ3+tNU1gZrbGUq3JmgGN2NKGGBzOHl
5XtJqEn9+tWsYDgXTJxIyTn5xEPhOogt6Q0L2TsNT6SPPSbhDuHtd7FoQFf6JgG7
bQahqcHOpnl5Hh+iEEHFPV55UBlrwpqqxEYQcllgL7wPJW1YoeRApUvU6n+GMfdt
jPR7UNOT0LBkv5Ac++baU1XvdqzOJmXK9nQoZi2qMQuRwppsWAX86OM8vgwp4ZnM
xRmslSOdjypeVfCrnU90ztd6uKcVk+RGGbQYbg7UrmrxYfKOLxmTmlHyMpLzbBZT
vyi3jJ6eWMMQcMFKzyNKoxdKwlTvPwYJAkaVXIbxgUwQOcAqrVE1ZlN32BRgtSXM
/n5wizGgBPS4CO+RMAJVP9E4r5glfPVf19a9E61udD9eettlc9XmFhXpnFc9h11/
vj1EJhGP42/pv5m3XQxZ9Mq2vFofhNuvm8NY8Ix0luSBg6E1QlMjn9I+KtqQm328
fVLkF4pzcREfo0C3uz8kCt+19NgDT5CDR6LLAu0qRhM6Q+AGQkyLEnttQOUKJkJo
okXh5b7fDCJtUTovM8AmLw==
`protect END_PROTECTED
