`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qzewMuby+iOSUDZQ2HjUyLfM/iW34rwQGuXG6bxDSakntM4ZOy5tp42W+DEj69vL
cPD5NXWG3RNx7TDf10ytlULj/mJrk3OWnonmx+Z3wNGqOq+Rwax18tsbCHUJ25QB
ReUG8554rjYhZDZUg7Ubp2gwGYcP4tKbAD8feHWWIDWFuwgt1LsF6B3k3QgVY3VU
GLiw1rBuRzwBkJIwRO4gTs26AHteIITgE/Udp5NjP39qvwosZyLsfBGjOWTgvyfe
kadlYXegxh2RjW28fuH7kgGZhW5cy/3FK18mwHe79jLG+8uw9P/1gP0iN3jMH8Bs
2anfzLk64Z5t3XwD3OKQfrbl7ElDyYg67XK+7gkYbPyMk4zArunBC46mOmwRY3hA
F+tZwu7//VhjjFW9dCqkNMsFvFtr2RM0v2uzp857XSUQM2A5we/R/qMM2UWRBBgV
37sPDJ3CAZKLCV3geHY4Yc2nH6jXQeYzpoXWqS1HzC0i5z/OiFv/D0fMegi0coZk
/0JzV+lmfOgJPOZE61aun/cjWjBwMmJ60g3h/XDmt/RuuycZApObTnu2rmT0LS8n
s04+v+UBde7iXPP8rZ//92VOc6sWDw9bUQSeZZO0Y169SR4Y5WfWnYq+Oh5J+UQF
SayKcfdtc2f3zV28aqZL93wfF2hD2wBicn3f4g8Rsy5h1kldlES3ycHZKBdfddlz
zAqtG6/9XYTaxKmDlQVq9zkLSt+PsR3cYYoXlHnxR2cnQfmz3Ccx2wTwBqNJZNni
JliyrBlTpmSnj4xCPRTF4QUqb5fRb7kwBaZlqVAD2QrMgMKYr0cJq6DSKub+jxrp
qvC8Dh40NA0iV8bkE62POtVc725jp5tLN4dDDHAbCCJIdVbHheIr6bVju5RsO6m1
rVqL0tCO2SBwuYpdZZl94CDmNAgv4UXiqacvEwpXDJPxMxcYdp+8yBxf+A2zn7Xs
dQVUtrf76grTd3JBAL74CbmhFhNwH56wWTPeRJL8u5jwyDQzZBkZNJegZP/bVdiE
aQxvaX1kui9Ug16Dste5GjLWkOKutMccCUaxENL/NBXiYyMhmbhjNNbQ93ACZGkS
xs4AkGvztA6Keeo+WmFDzzPUK3D61DptSz/l8ZF1HWj1CIcTIxqMgNLndUbxnPFs
lEdb4znyrUCQDEu2KfXMMO8mSDbR8TuzEaj6U5uFXXJ8vQEW+/Z3L903sd2FN4iJ
n8RG0PMgmXpCq3wc3JNM4vW7gShbjXil2cGK1B1FqvLr71+3KGvGex4XP4VIEwKz
gvF0LjxKm2GnGFgVQCpvQXfTiE4hC8ApkdaF/jHhGC47/eJhhNU/s5mxfOmstR9x
OiGrn4lgx8G7wyEQu4ki5cGOzyPAObxxr41UaOeZruL2tXxiyrbEIkiWF3ZMpW7O
Gznri8e+10WMFAT1XrJMZLEPUW2QpyHEdszeUc5dCJiz32tO/tLCUmOsginAINWc
78njUraUmCzjCVdNZ2Q1iJD6pahUIiqz3tf+7FTBH/R6edOvwGHC/ndJUgYoDc5J
E9e0U5SPxFTNUAnR3OcwtrSt7IyxPZzFL88HHbY9HzX8cd/mEVu4oL4vCVBjlJQM
93sTJvLp3VvgJlqRc5a+hNP66K6AvR2KRGPJMj+U1Asa9+dJG2D/rvUFcNjaM/4/
DZAFCWOqL0tq+LrvekwacARju/z9d1ppD+oLBIjJGPZzNaHdAJYPTsQ2EaFIwizZ
UGP9eUFU4/FbQlGAbBuNERpoPh0ELFxZ4J0rZeUJvH0qyGyjCWzhjl0N3yaqu9Ug
1rxzHDEa9o95448wlNxu6JbQsRxSBxiZor0Oe/6UpLfFReM8itxOEG2UQYQJf30i
WKVl1o3TZCZrJwypPzo9RXSdOfnq3UWgRYxtfEWjstzg7RsrQL2/X6N4UoVKQh1z
OtRFQcoe7UUbn8H9mb6YxC6Wn+qtkgOkkXEfXFqLHNJCTckPeAw+KGAxF4MW/Sro
hMvGIa3XDR5hQ8PXE5vkVCCK5ciMMLR91Pm+4iAcFub+s5VXyIO1PZbZRADkksNJ
E8KCxzhdWJWhu2J+sMC748JeBudQur7qwMP6QeRu9lVVOk4Jq3zi96ojRyWaCYyQ
mxZ0ZQSmWTuetI2xKXpqTJxHObtou2xKeDkt6rVo+3hrXyvUyjibavlZIgTjpImo
fPH1cBPxboWp9LrxRXNfpJOFsRKAyLnY8Nlk3DglvSpRMMwQxL65nCkaZYDacEGL
eySwJ307a7+nkDgFLzplpy8kVlKeVDJ/ZX3EgtgKfotC0PwErPsBQIALxMUCTlLh
+x9yEOrxeh//F0gn3B21t8S+MF4QsjH3vN/ImmlyknJhV5d9MsoEItU+AOD4w+Yy
DJ3WWBBMQVmfo2RBeUHPD2I1cm1GzXOVd9ZfhhdTeutrc1k/BFQLocSl5k0/tubG
SEhUWysARu2Ad8g6JJuH0ZO2b1XPxiT3PJvW/7WcP/rKF2Ob54gIwFrPUqV0SX6R
008/y0LaySQ2BASWQzFbOGtLm5IhcFuNgQ4mcZnEUVa7fzhgqm/4QJ5ykoVBlylL
2wW+HpQSXFjPBYl0MVhpczgYZLSoDz3WX9GaYXoys46ZkKmfym/j9oq95CN4df3q
Ml6QjbCSUETU4+RcvrJz18BsxNkvHUdLRm5nBU02TDiMbCrIkr96pBCFV2/+pvv5
xscd3NOnY9SZSXhZS0RK9n2mDFhAL4bvEmtpM8FzlQq9cqA7RQexiGb+o+7SD/dG
q0TTMjxvzPCFDhrZlAyeeV+ogxF+vTkJ5h+krpvHtl7sJqDigun5nQuCrlImpYPf
/Gyj/BZ2bM0xXXbd28W6tb7x28D45XpMTMxBfcXf2pNFdnKvGbyyISoyAgC3/mXP
3Cn0MBNHUKeJ6moUIrD0LFH76dYcSEtkhJh+IYYXpPawTl2fHMS88Ugm/6bbKzXG
1FiFDHMQc4FEoLz+0HZYrkpXqLmULgB+qlhLzoE2NwtghD8/h6hCPF7oXlj/21KX
rbRYFFFUJQJKOyJg6zQLgLdr5W5ZIWbe9Blhm2JtZC7GrCr5aW+qnTitf6+oLN7b
jx7mci54mYTjxWgyopAjEl/J1Yacqdl+sm/Q+kFLvPjPLhhuTf0EcINHnajIk9XY
JYYBbzill6yCmX69Un1zNOrVQhTjuYS+ppgc8YwjS6imMf1ARCKXkUcOQugCqm+g
wEjq9BPjMHrhTealhsPFKKocT4BPn9jh/cb5rRT1PivPZl2XId1S2C7g+w7zAVHD
bn8lSTOVL4tUXU0jf2UWtpF7DDMMwb7wLe/Ntp2/BOYRzTP2yPGv/dGjl0fCsck6
UrraATwfEP3XPNlklaD+epeqYJbEu0/uR9LKxAVkLcLWqqwKaRCieqmpDkZ5HojW
vvC+UZIH3ED5TUuQo+BOouo1EC+6NMtKXQ2eTb9eieJvXutyaHhIopsSrBLaJYzo
0Y5BAXJmkkOkdXLeKTHSbk/QaowUitPSQ2UNrH/8QBvKacv4cdsKcQPqv9ofczK2
7wjJx4mPm4/4Xfm80S+hPaRZy5jI2qgp11VjIn1R3Vwpo9NK6Stv/LPQHkrmqoq/
xOp+Ky0JXAM/xf2F7e9IHyvEB6zcsBmvLeEAE6Wx2FFHQ+PUO8x9tzg4Eit5GTHT
4Iea31HyDCn4soyvPUx+Rcal5IUO6EYPyHg8eS0182L4cu6Dxm+ci8R5fVsln0Wo
DaUKS1wN+KLLaBxhihXjagPlE2IkI9YL7cqFarDDPbVREbY3qYDPdDAPGUnTCIJT
wVE9feRZjNttThHjmEQ39No/TU2cXiwI+fqDStf1bYam3BrazaQn8Ws1kNfyPqjk
/1VsimE/0Xt9JXv9KCSgtQeCjBotw+XNOIKeXkwhFg/eIOOasnAJcGtN2y6/5y0Y
2N3modoxOA28bUnZvF4wMFlk5cO0MfKNkO30DNB25oA=
`protect END_PROTECTED
