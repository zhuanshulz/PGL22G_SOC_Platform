`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QIOsl6UZ5MRXzoqii0xnyWIof6ZvZUuTZaCaqSYbxJUQI683M1btD7JMlbX4tRPT
vaR+qcx+nsgYviuHgUG54eHXoj2K41FiOC5JOaN0RAmPj5P9BmyxXk0krhwnOLPC
FqQYy1rFcWJNfx6ravO6mfVDrLfJbI+ZOWWl4s8q9QRvzDpBiGheDyAjGGE/f78G
9UQVDQoVEzG2wLM/wMZCBugguyXCIrAlYWnN3HOQUoK83KdOx42mpLUayQi/4u55
yxkGVY29TT5cmqCEebbmLcJyIDSU9mlDBcL80R9YR81sBAK6InZjUyRFbtOzWvxa
IP7sDdB75rUIBeEQ1fag3mWVPQN8odjXAjQfa/yyNJXtrHru5QC9vW862DIxqm5E
9ROSJU8wobgTTI9J9rRFyE7e0evaJkSN3IRwt0sUkco8hcc353V4pHkQBlztp1D+
iL378xlykGPdKJzJTxZFKIjh3JepRyLZqKosS78pS4GLYy9jTy25fBBfz4pZaYGC
BhmfwnvKtMQqOrjCw0wVT1dzbknbaKvIfs6krUUvT0v7/FCXStU3uu/1oVpV+GOn
7G53Lhj09YxJRovQow1VcG9abHLjqfB3HIaXy40QDLUiuoMTXO3FMHPvgAey3xkh
rwDIsFAEqGYTi7+UKGsU1GorCrpRuGImENUvTpopoI1i+LELN5G4HENesdSFxVbc
EDA5Q0puBG0/AIaswmG/qqFnxh+y6zekKRP3sA1YzKMg39Q7Pz2ZHeQanboQfvFN
SGSgfzDvMJoWLIHAXdTaqgU0dqPNGDwzRkRFGRB8Gk1sa9+quQ5NCOpnjKgT5HnK
1d9SDPrsksNS0/dZzdvCGjH+OPIlls+LBz7mXvtswMczbkBhFeRUKqrGciLn0Xse
EnbRttGN7cqLW+hgyDxuxDQZaL0uyukqfXyyiJSYjp6JXh9KJ+FnjuHuFNbLsXwb
mDceHxoaJs2VpgetqmshkcgSMds+sT9PB3YlgqYfwrOANlEHlaknO8kJA5O7UveU
OETmCh2tGWUM/fF5a6PhJ4NfQmO3JXUDr3zb/BSChab3kgmtFv6dRb4AzFquyVEk
idoVOD40YJUaKstjc7nJjqZAcTeakWaosUHdZYqxnSK8l8UBVrYIAmDAV0zstmlJ
rPJVBdafKeM8sA6bHne6EazPV1kxP795V+T4nOyEmG6lFuUlMMpAcIyb5jXpv4Zk
2jSx4zcvhz862b/dynJqzY3IArsge9RZJwR172US/B4RcthsX28zMFHgDDOgBL/2
1BYEzdTbv4QsLePbYP8yt2JCsbWSr4XG9ynTYZo3Pzxzk5sWUk3AL+2IUiPdPr0Y
YoyyRXt6hv0dmifnI7NF9waU7sq/ek6a8O70cnBuzVDTLnYNiHoLOnZiVJdBfAF+
PZMYdTLT2T7JAiHWkqblc/4F8c+OjJqvND3cjUr1Dnobl05LZUInjLyIBtXlqIAe
zJ+O8YJFrXpqwBr0QF5y8WhnSdhV+gl1+QwAVZkcmEehMgqVU6914w35e50EGFqH
USw+0Te//uqKdopxGQd4o593APpPJqJ3S9dB6EaOOf9S2D7GJVZQyqdzSxFUZAaO
5o2z6zhgCK2hF5IHLagQd6WWOPiI4I2EZzs2MCTUStWGI6AyyT7fQgiBwkXAuIz+
+VQzCGNGhf3r7DntIGRveQ==
`protect END_PROTECTED
