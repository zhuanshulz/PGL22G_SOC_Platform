`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahEF5sA5aoazXTtASpA3GwuBVcxw/GmDQWsdAYoWR7N0tCh6TqQNYiROXgqDzFLH
bsbXZdnLgWi2RIShbaXYnG1v4AWDBQIUnor49sypZ3iQOgaULvRdjgQG6h/3R0z0
RT2eWewsGlcO7s/7OTZvkrhNkMMJwtAygWCsjcK732TL5q2NlayMovCSYzyrvo1l
3adkxChnUM9GdVskYhl/TpmyUbCBzJXIXAaCl13g2YsWmnBVFWVBiL9BGNtZMFf3
QGnyPhDWOrXqTPokPQn0nEoxOiizwdkvBzdEHW+mA+kYh6TX7S5PZsQw8aPPthd2
p7Pgp2DCEAtgnTJipkcd/+X/Ab/QTJ3juqzTwezBI9fPTGEK/fEA4dVbPiG4r7dV
SeDpgJRevM8Tv7Mvbnk/tFY67x0xpILf5vxb2yqih/axzL+lrla5dI4gEMZNzkQ9
SmFSGpGk2GO9y9I+JUqeDEJByFvYVfN47vVAAUjHAfFYA5xokJTuQ9sWhEr1BKrz
XQqBwan1beSXJgKJdtkm38XCtrWPn1RMq/jd54i2Z7lNFWezKycJdWvt/56d8zOg
eqF/2/Y8rGHo70Tj33a1zOFZLt10HkIA0w5OjdG3nIPWfNEA622Iz8cQCD4/PHMh
C7zhXkYyFPa9Z+sPD7W3DkwbgrP7PfMFvkzvN7dD8W/yOTv1nLpj0kfN+fV7qVQU
GSBob6Qka4TPAzrCww5es5A+v25L9B9yeE4xkGw4gSFxHf+MHSuejoeDlR0VgE93
nFSnt9CRhea8kOYduyK2JwTMjmxOr4rzTtOJqcx3i2E+lf0F5oPQ1mE+zAv/WiXr
Ol9NzNAYSwWtteX8YrJUlLRP1vZZy5wRdgwZ3Emu67MPnnbdkMM4B9hvnUJNy33t
`protect END_PROTECTED
