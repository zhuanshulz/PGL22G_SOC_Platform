`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0PDWGRrm7CeDvv0fO0Io8VJ4teSsxUgxuE6ikM3hEiBcM4dzEylLPvPrgOU4NvD
Qw+eCMM16Gy8l5/b6fU/oH+59MnAD+WOF0oK11la/pI2eAGmXzFHcATQYzEymHR+
FUIlqwixg4AIPE0xkUd34lwCPDN1y7peVFPJcXGkdOZatWa7cGrAnBBv4iBccIfq
ymTowMzgrPufNQdVziLXG7dPwUlP1DibbV07wY3dZar5lw2oYm+5rfMil2qDqGyM
yG7CUv5xRcCw2Wfq110U+w9cDSMeNHYAYFoBeXXznxpVQ8nxYU1op+/vmIZVB0iC
+0iU3tDLec51sYWVVRFXSwn1NjnIy6zY/etTXiC8HJeQuPR6AcTYX9iG0N4/4Lwp
ybGajEdkCFXOPrQL841cvrVI88bwzd+vMB7neR2W+1fLP2avOVeNzxTT9wWAFJri
PrbyblqEoGTLD6Fjl88gTfrhEZkD9/jt9mYB7OJSPOPntDcNOstLJv6m/VRhu6Hr
fm36PpPYg1vc5UBooIJNnK5TUsXNRNHcfPPaHJYOk/Hw/ehRRVRPo9q2EEoiSDkA
ztGTFR5aBjNKnPFssPT/ZZLpSpRvvkPS8+qra7pKEpWSyB/2fBfmPH2MsMYm2H5q
dRTo7FLvGeYS8A6olE2l3BQtDhhKkyLyIQQZKZyDyNs/ubw8ec4nON1UhL3gClED
LBdD5dx3nfb/6Dvb4YeIZebV8Pq1vZtr1mifG2iR44OtO1qo5ev19XDT5VHaktw+
WPVzBorwPYktTx1YUQayAzCQFKod3K0583BmIugjGqxvd5//8VxThWmKNXJnJi/j
zClSWXxwcxKn8mE3q1mOrD5JJVOlhC2d+Lmn54xlPQ/+BkrW4XNck1pKX4VeR+9y
3BtLuczdPQ7lESrEC4v5aq8zwdZ5erng/P3evEUYzkbQpdAqrl6rGO1A3B2lQdJp
P2Abe20jocXrc2qB2YEv933lJLEMUBxAEK+sPeK3v70c9tDf53FJflfzleRYTH/2
V3OIK+gAjXKfB9N/l38x2CElQGSDYIp4nWDntVerg6nR+yPAUh5bSHStdZ9veCWK
4nzoN7RzItzpVE/Lie34D82pqScc283rSEUwtIEmC2rtvwMxPEka1FsfXjSws+Bu
6ucbTuzhcacF4dq2cWKaO3wNCbcZeoLRnrVA9PINu6UT2Che9StuRoY7ECMc1WT2
bio4m3w+djuJbnGy/f02kJFcpwAkxnYLwV8hCJ92bOjqXcsNu+74wIUM5yaLPXnr
kcJtblleiq3aC3aY1/bQwkKvxcpjNhvPa45wSxad21f+DT7nGTY5AhnBpd+coonq
aBTKvAzq83ntO/yWugeZow5N+EW6VgPB0FSIt63zxW6igE79MsWcsvI/PUVH8M4B
tBQZQRxc4uizRgZUZoXa/Z6Sp0+g6ZC6xGAZ6Q2SKIgqXnP1aG6BMznRMY3+yKfB
guQjwNt/22AdcnDR2An+DgMbdzSHZ2rg8dnoOsvlpYSg7gKNbVMgPJTD2krvxfoT
`protect END_PROTECTED
