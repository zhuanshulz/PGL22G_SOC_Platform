`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3l7uKhKljCguOjcJkGSNc/WMsTHeCv4qc86O11+/8KDX19zWCMJw/HEafDenS90f
RTy1dWsFIQDT5guIJaqFTsH6PJ/vDVvMDRbHfX5FwZlPUqBBIylkd79VtaHbmnD6
oJ3Uq5iZa2wkQKUI9jgwFSNsVFhAdgrT8yOrXc+wNjsnd7dY+p4QQ7TInKqSuGLS
Je1kcg5pxyWaXGL+tyudSgy4Z5QY9WYYefNQGTo2mwpQAgpn7moVgqtV0Jkot7Ca
LiEdTI4oVpElzNKeipQX8VWi3pDgn7MaHTnFEMl+rG9SMyt+caUXG5IuCFQmdJlx
+vw7FKenRlw6oLRgYVMvyzntmiuOCiQ64IKlrJUl5/ySFsIaEjK8OOsQWMoM4huw
ZgrxTM3HSEMV+TWVc3z5Fg7XCa6FvOHoNO15K8rZilY8Fg+guXKt43PI/8hZ7uYc
RsmAfViMhOGRwl0RNx/6qspHiVVddvFDQPZaciS4F364uFrFYH2Fl8kVzpPq36cv
xa3Dr/I+CSOMCK3TiICQh1ZKWUZthKbMlQ08uMSbA+3nuuDE3Xd2tdl74BqOEH83
Jz8aGo/2sCcu/wu65fwgurHvX2L7Kz3FLErm2NEPTEWbUhmtBL4sEYsQ6VFc38Zp
c0LmX/2P59xMfydHvOLXQs7/EQow7bqt5FXCsFHBlc+5/V1kuy7uzHSf7c7rORUJ
6NEyTB/UCgxbzhqMeX+biDNJR38JdBVsyvT7N6Tv59pfN1KEFl1WTm2P/BYUYAgg
h408SQYQ1+/m7aFF1b5HFIcD171Qc6/oy6p4HG+k3hLoGS/Mt/FoWAVMU+17CAYR
caw9Y5ovJgdW/srJCahz8a2a3Qc6sGwDA+6URD2Y6WvPlxcgCc4c6nMolZP0+vtg
6R/Z0sNgcIau8Xsd2g+410LzXlTz70Z7AY0XAhlq9ubahzLomISXl8u4xMyYET3L
H7lR32JxJ9leYn5mn1l8FaSIlo2kTxj7Bm15/XUukztKwotk6dUiOtjzig5yh2uk
ZEdQswJUVKSCdUo2/CSlAGgAhhl6hBRNbQ18CUuFU6nuGUTrbt7/87//4E9t8ikS
VU4vFPy9HYtsqvNJM3hwrPg36dN9Z2SqEJYPRhev8DX0ttmzt+VFy94q/0mYPpuJ
3vX6VcGJlD+mPDxO+fOd0nIB3sW7v6eKYyGPeYBfR5la2hdRiVE1D7DFrp87HBOC
G4rjfvjPs0KeqO4U4NBAeaJd76Q/RWaK/ehOsh4Lc9VQH017QR5/2oy6BUUIhB+9
/D9+wfdyUg/lzVuZTb5xJfqvUk8uQ8WKkOuH22AYJpYRVgiWhB3xYoLS+pWxQ2D4
Ix9sjGjbjWAKN2YV2oOPLQ1AqKUXmT1NCDXlA0TlEzCC7nysKCcIZZuo796BUsVY
NlMEvtWN/4qYq+UgPAMpOQKPU8x6ivLVbcJc/QFZERBkGgdz3gCams/bD9C/r7UD
Ahpn13M9uz6Ct6AndA/VZ5cWk5NArSMgjaeE5/vokVB4cF+hevuR9cskkVMX+9wc
p0SpwM50+ULiqnM0oRxS9GWSww58gXsjXZ+/jXPBuEDZfjPOKNaXGJG2m6A1bbhH
q42X6SKQ8A7yex0jXidJK0OrPmUua0F0xwpVnPNzoyI7XzHQB8Da8qQJT+Uo7paz
zvJoFaDO2fWs1E+PiC5uUG3TpOUIVMI6MuWZ9OX9HdKnW4hugFRWg27EHFS0jUZG
PNbWIc05IExGhOHykbWPtLjiutmTv0FVbURnbgX4b9D3+tpQjsSRgZn0UKiBTGjL
xhXZpmvv1OzNYhn6OuiruageSt70zBWEMxh8jDWkbbA18gqqZ4EPWDrBHxxwgXnI
U4unH0WGBH99O88F7wBg9pRKv3Nuy9Giy+Vxu3+g4p7YDUuc4b1PuuQnjKlsGEu/
BD0oeNVlU+Kir7KWcSS3rty7T3w1qGiGU7F9XX5e5ZAh+zky9NEGTN5I/XajeQ4Z
75WijznS5drbxf4eye+PEZ2iw3ZPxQSVi/HOMw2gfbvaQOtxHzWTiQksz4y0cs5Q
rkSTBrCKDeZ6zSftB3NI3OenFQvhoY3gWbnzfUMIdPEIrOjbHFx6B04W6blo19Sk
DV1wImtwhKf8nJaoXrKPXCi1KS3X5kvTAbNZTTxx0qcoArxO+KaMSldzkvAvsBdr
r8CSO61r/9TsNN4CNno4klRGikNNAaX5/5/x4yrajVo=
`protect END_PROTECTED
