`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/rFieNpu7GiHdr91XAZQLK98z9d+PdtfppVWg+jP5/lvA/WjG3azBbyA1K7zISni
oKWruFC7jAYIpVlN6BH9DNG//HB/1sUVGfOJO62KCEG98pKGVt+ZQ+MJiAkyDfPe
//3K20hk/kod8hkNDxk8utSOqBY/CzWUPM1YrF36r+VA+H/X7wK5uf/zl/oQWh2J
D4IM2PuRGdkNANzoUiqLP+Pd19AoHPX+EYSWb+ezOnq43M1zy8/rD20jx0GVVQUu
2KNPiBOOuDLgTUh0HR3v1UkiHR9AnUmn3cksevjRdjobwTHcQCtRbmRKYDkPFBwk
LXPz/9CB6/LiPf3Hr8PY0VKokGvp00NNqviaij1Hsu69bQHxsqw/xTre8M1HAnqo
SxynjiICFDX6IB++O5Tf6n/y8Oh7eOjWTG/d8Hm7ddA=
`protect END_PROTECTED
