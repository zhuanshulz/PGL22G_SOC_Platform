`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VxZMlga1cFT++xUKQNQY84KB4JqRsAHQCtnvvn8H5XJ4LoOPsyHwyEV6xblUoeu2
NzP90PPRD+AnbHLfQ+LpoVjMMBo29nox7Q5FIQ2XJ5EkaKPybQJeQVyPW3gnoeRZ
HZ708Xdj/48EpraTS1+9c65Aah1S62FUtU8bfP+rrXQtwL0ypewtEUgonDni1806
pVeu6FS2AarTZh1pwRKmJuGI56pqnzUidPkC4IqFyh37pAkWG7/SWgKhhFg/m3T9
r00lOW6FFHEjrtnjSz2xKhqZTUz7BgBcm1kLwcE5Ejmm2fmRSedAIz0H054GsgEj
2UUUmika/YyH/E+J7oknEc12gc2AKsiaCssuxrz18nxked/2Jy/dtjiWltUYgziX
98ViH+ZliwtsZtWb47dPstGhVSUDaFvpFMKrwDJXP+2pi/zsaRFOlZ0bcIBq4jxm
+B8azEVnpM4c5H0QT/jOk2q06p65Uj6/4B1u2dzxvSI=
`protect END_PROTECTED
