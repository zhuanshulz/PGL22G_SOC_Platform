`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zUPQQO45s05wmHer9mx4LZRzktt/RL7UKaF3wbXFZe7CZdmOt4Sh91zAg5WwZ+xI
lq0d1ZRaXwTXI6syxc32DyUIVH3LqhmT8HVB6gQptUFX1uLq4CMwdvzXxqSK3fjZ
XI0O8EHcrzsnklwwGZlmyYQ95CqfnLVFAsKGTvHlbGTfpyuMkufAe+YDC0OE/ox8
5GmoEXpBqNA3LyXe3BVe8he00rPevfG1YvyCJnI9r3ws3sow/Yuv8IFVnScXfvcZ
Qe183iEnje4425E16eVlIUXtFJikt+CX4ru+hRtZ03/AqJ/kBlp/iTPGwQIMLtvZ
CDf9F5DTconr/9oU+a0I2nRcBXnzct891RvsHKTE9lowNgCDMt/CqA1nF1Uht1la
LcpBTapPVzHLEYW6uXyamjy1v62z7nplCjw/V2Uov8HaaiW9ey7ppZ9D/XqSCoWA
yz23lOlCO9NRGk+hES8MuyjTQoZt9uS+MXC7PC5n+VDASoBHhCpnEUA6s7Lr28je
O7kwuErqFx0n3oaXN8S/rV86GKJPPI5++c3SnjnGdIg=
`protect END_PROTECTED
