`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+zzoZl/t2mcU78iEJCizKQeqptWFtjUrXQV1h5+MFgSTGKrdKc5Di12+sl4AUTfk
Y0qRv3QR+q6Jay3i77P/DQx8cyuw5qNEZ5HUjU52QynF3crWB/jcrU82I798+MdK
MZWd6SfiHnGdatCI1i+PrdvOC34u8LLgeGrEGcVn2Ytqmsy6lG1A+rNnoVQe+Wyp
88lDy+pwvuKonn0JheyN4m9Ou2uoScJkF/5oj3jOurBPERsLBxn0aHAMSM3qIrHj
6L1LO3wkvUg35hRNwXsmyUjwNnx5l25B8cphUh0DCy+h5Rp7tKeLhrfOxCpRTFW1
XUFbPZ84/Ebv4Wt7PgxSW0KXs3H3AdkZ8tzZ+ylqJq/Vxc2L95wGJ+x1lA9/Vc6a
/GBWp97DYNJfW/4qTwOm3qzW0Xbfy1WbroOGa/O1eSd3qYcKv+Mob360cOD0Bujh
ECu3hq80xetD9vo/VlYDWmAhH8ND5p0JSTfAR3r1e2i+/Eje2m4vP00oP7hazRnS
s2z2kEMH04WidOWp20Cy5bS/G83s5jZoNKpEFNF7vyglr9HeF43puPmL0CMNroKY
h5z/ycXeu6skYIYQLL9w1RtyFc26l80d3tgZfAs5yIjh7qzUQpARa9+10OHB2imf
UPtWadEs0t6yvLtTDqG5vMcHl1f9qvwKjEaYnjqN1OSHcE8rdMZaf/qHZLfnPoIs
hpupXD9Ag20G/10+sAnTgMIb3Dh6iisLYHjPiFIoLB3FsJL2SMn77VNUlStDuvQ/
Ydnnn8MIwnSY+g2nh7sJcjZIBBv2ItxQyZ4AAJP9Bc8R8qASU8y+5Yy+UQVB5rt4
V6I1Gik75HlykbvmWL8sqhZed6OpmLcI1IfPY2eMnh4Bq5vaujrqGPXKCy1Gy/Sm
qPOYy2CEkJiThgzoZQgILbS2grvsK5muS/D9Q1vuB3jFf7DxuxToQ391vZT6pz8m
YiyzeQRguvoi3BuCwGyDKJkvSBD0nmOXNDrgV6sKytdPKtyt3Pn5rxztno3Vuk7O
I94sskvK5oQmA/8lp61Arynx0DE4zgXPQ03MoalY0dE83KXoLSaDxiCJlMy4XhXO
wzeuOPhd/B5IkkMThsS+n/Ovra+S/WJKk3QO5CzaGPFhrFphK9UdmiHTUo4Y66yI
22WDl1kVdYhy518xxJWUQjK1KXLhLyWcpuWpzjtFQwbehuIRL5SznJcdiJoGg+5O
DywwvYt3HcwJDvw2ahnvUJs95XqkV83bWdTeR47IGaO7ZopLcsh/xippuvgeWLGe
81OPhp1c3yWPTSugOMH6XdIoRynIajX+Xfaik5p5T1DFDH9OvjgFlIy66piiOb80
qBKlyxng91d3TYmYnTBwi1gmRNBok52w6cVmwSu4wIVPSXBSU6InJEAHlGMrTgrl
TUOX7dndnOAvxZvocMD18eFXyYXlK6972Ewh/+yOygKprQLxQkT0amUfJ/8QjDyF
dBuZVI/nlnnkGDfVizggmtF0Q6wE13vQeTV/JoS23oJeUajkNLZ2LxgQZ3vllIyZ
pJHydx0b/44tSgPPpH07wtk4Uix2n0wNXGwzsVp3WbDtURpu+MFNb1oIxDpdFJlZ
WTedeTGv3PMtqwE+pVnbLIZs64GQCtlChGHEFE4PfQRFkkvT74pCTxAlnO8Ezbay
GrFWrWWUeOYUhhEE6Kntiy9RkZSc2ZsvpyClP8XibXrPSjY/YOlkefCgzWWJhslV
5XfIwR7457aq/N/Pl5FSPi8uTeZM6I9Z2WcMY3vzId0jPjkuo+GWU9NZOPplBdRs
WvkTAfumhGdHQMi64WhkvR5oiw8wiUzjNI9PJpmQH0cVFJZEzEOBeoAFg5bB3FZT
a20kC1b59BpGNslZdl3vZvMIqps+9R2irFG2E5jktYxyOA1KI4pBZjl2SLzJVTQ2
WA23KNqiXI++lauTzsIrGRMV74OEjRzGBRbKVBKnmDyGqQS60Vs/AXm2eJCsewgN
f1Tqlrmql2xNbHkP9ed7j6t9vvnu+uObKxJCw29p39Xft5FTcZbje47YCRg9dRKy
8TKDEJSeNWAI0mlhTcLJQJn3v23Z0X9Er/p+A8LRHYgSgdX0Xb9djq/5rNu0s/yi
1s1ZGFk+snCNamSJacgJASFl2W3GNOUrwNyGnCgoWAj1MuQZaElLijd2Yz3irSl4
r7X+ySxnhfmj+4BDw5shqNpK7TdLCp/mi+eMSdeDn9y70ljBFe+Y37TDvkgy6iNb
fcdscB17Dhk1qowtlBCzWZNB1oe0OmLCNmRh1W7ET368KTcE+4sQsrgj3UNi3QF7
NsGVUSf8DTAZkz/Q/lnd30T+b6r7FqaOH2t4KxsiQOisYz5upfLnBgNaufF5CBbi
1qpx73LLQOmMFAMARWwpGU5ZLzZB1Z88Z4shctCApmAO9RdwJxh3uRWpOeoWTezh
0K8bKv5xugEu0O/yDK3wsedB0+lI54QL9BuqItx+yyhQItrnMaU+qL5lxBEArZ+t
3ayJMvkpjXzHERsKkNOpHYKyCC1shZgmmGqsK+pOgI86+u1CUvoGqC9I8Je0iq3f
TtcpwmLB3460686/j6I/RiN2Ga5SQAfz7436mP4m612H6w4BCfvtEd+0O5oeuPHl
q0JTO1BL2osX7dd4c0LGWAJANgirDn9Ax/QFKLSB7jnvb/PkJd5QSmGGHWtUJoS5
pyYRItrDEaPubJKVZsg/Kp1bUYc1fOvHynCDJEkpFze5d3R7KcIWwL3prVzlU3jU
uVSqnQ33RXgZ8ecX1h4QVPUMu/sadU1mXosZKPnvbhlBm/j4sk8OitrRHDd9vbtD
OEONDeOxORwQ2JZysmsfJL2STUMSYKJvpqbsJiLtvwV1EBrpgsmPeiZUDfW7NVxw
IjZMyVejIB77qzr29Whbl+HZa8sbBLICHoVeqSQeCOk021BCLItAxyC4/fGVS6L9
C91r30iiKS9OgcB+AWDVUSTGdWDt8tVpNSH07ZgYPX3AX8qCE1LsrlPh5T5hGBA6
h3cIZCDvzlVkqH22wIeU7EbEfMX757yInMkyel9/sGi/0gSmhd80SIkM/2GAQBPz
9AhuolK208V6YcFS7qVVttYk/6iV9+bsxZ2XIy0Sc0OWI/lsXKgRM5JfeubH3bY4
zYlesVbqEKUkfR66JHeVy8+RINt2AJndaZzRRnox7VWtUJID5Lr4WZ2jm9EZl+jS
8cYFHlzRdo39xnIG8nUwUjRbuiayuemNWqEhAvutg90BGt2VQUKwBECRnURqK71v
oMsyaqur6XI1XXA+Rf9Bj4sSbo4VRGKS3R+vumyK5tHvccaPaw0oo16YTMMxr8qg
0d7BdmNn1pLOiiZKM3lYWTOszIyAgPflhiWLsOnMMTkarU1LrlAF8uZWkmn8pSta
74v+s6jcSKI1i0q9mdGl/CYXtXPlI5ysXpByBCpL+y0+EacbJMEIIH9COI5yjeJD
bRiGHM/XF5+WclN1CQxeDDEVDgld2Qe/xx0vo8VLFE9+MulNorTMvGesMM3JRZ3D
g6IIo29cmY+LBRG0jzCCsUBAHGZlStcw7cNKDjMxF+L2vCbvjl0odaXMQCCHupLN
SY1w/asOZW7MdYFtB+9mliNLwpepMO52wHx0XTU5h19ryZh/RdcKUDDpQG1bdGiy
ZEVC781oKO1APOsFflEbgbG8WMh0Po13J9joWfkLKdSSpgJ2AnU9redHwZL4zwNa
gj/ehj8EJpKZM6xL2GEr5mpzpAy7+wQDfcYtCf3a9J6d6/X5YlFGuiguZuF5pjBm
U1XQbYa6bwdYcWvDifnNm04CH4ubtPmiTmET3muWRZ1u9fXiBwZgK5ngcKPky5XO
Yd4xVGOPVrDVYZ0ri2DKPExli+FkkMOzIFhw6CUVi4pd2ZotOIB4y3ayRHNRk+kw
qsG2C5M8x0F38kMg3bjkTBJtomwFIXFu4Q65AWCwTHZjaalG25fJ2fwns1HntAaL
KaBeNd5qmIDgGQul/HKpKeUhbVDEOpDwwDGjJfs6YTMj6OCvQHbtRN/1+7CLqi98
W8p0EFl5QlLXW/1F2hgUx+W3POIC9OxTV7zlJl/iB+Er/ec+W6kx5Fl5wVUbb8Xy
/ON0QVVaRV6TQySEnklL7QJ9k3Enz7CWMVoZocTe4N4xX1Yu3tPEVo2MOCTLcW1T
OuuzP6w+pgJI/mUEA2/BL0LPr+4IbTV9+ce1GTa638qDtznSIX12dTh7XPz39jNx
eW2/sfGfMnDrYZfuvGnGnth3UupLAC+vl/SDKJzBST50w55ofhXC8Ye7ULLXNT11
XqrrBQ3fDrxhs819qz9XAzhypBmz19hsknewGDG/S9JDkBnWpw1n31oyKoaCDu3N
gH86iaLpHGd8Qta0koxNsWNzgx0AnBEyRlZpI4rR3KSz/rzMS6m0XixD/LgsccDh
qUazUtw2pF8m6fNPbxT7urbRPBLv3m6LgKkFagZUNRoNc6zVqdzO21YPpwNPIDpj
DGTtqzrFfnn0OtL3Y8jrV71LMtCVm1qGDytvJnv3BNwWtOgEGXh0rJc68ozOTLt/
mZ6ZqJ8I8RipPQidYOal/JupaDeufuotw6HfWkUlV+PhpaD5LPmCERQGAhMnXZV4
AeDn2StYN4dBn61BqSg03PMYdcyP9FFuBSCnJWzrmCrx4As3/sF6gOvJn5VE5UyS
qN1BTHUWGZ46BpgCxIvHJfTy9w4dpsfnQk1NM/jdqv/rCetm1wuwZ/prxpP+k+p/
ChSLmGGvl8kKgK5+whGs1PmVXqRUeYdFTbQvBPFv7ffU9YTtgAjuPQC8SKn+/UxI
pEWE0hfpd8pk2YnzxlsZUn78vizHxtngUd2zYx4bEaYBUwVpl7faes+P+Ie7pEph
CJHu5Ad6K8InrXwRrW/z4hZYq2KZjrraXrWgdcUQ1pq/WnrBQqEAlZVEgjmBSfXd
QBUwO+jH1X+xk4RzO32bSYViCtZ1vkJZDmqGfqP18+H8JqEym151N8/ArJEuZ3cv
9BdQ/OczTqhc8ehcH52mcnqCWEAZ4Lnfxq2vCkxct3i7W7mIqmKxE2KbBXCZYmSO
Y1AYSJ8TTyMAcX/bGLqhhad5Sgz8U7qLBfJcaoJtF7XKvsQ/gqCPyqmwGqb8NTw9
DVzpouNUnZmWu3NsU0gPNfPWe6V5CZcDwjsNr3jpyUhv+LQdHcO41gsBIc12Mu/c
I4vlvhyYaVXkPIpstm2I29rHio0ZCNr2C7gxj9STO422A1qMhZLfdi13Jn4pPDjB
ViURJZ528XNEEsCxDRCBZS4TD7cOi9bhNhmXYaMrHnhxjIHJzwSIuc4mQkS3iAAl
rqkCe7rbX1R6kYZnBvBTsPsuKMKVKFG6HlOkITX51JLPfvPjkp2sBByMK6gy1XYf
szN1YPGQuyjGrA0jC+sHd3S7VYK5JTpRYBSY08JbaoYZUVwkId2Jlz+Pg5oEFD5S
aBJhuSK0bV6jKUlfJTX42R+BwlEQVtzZsDIR6/A6/bpWfQcPumBVlhcXIqIx5tXp
E6SPpTUcGQPkSxajFLGgKz8x0bnLPzEl/N55IdohFUzXc8LeaRErz16U1NmbP0Qw
xxihX36I3n4l53xBb7cIGSuF3wM3K3Hm3O6hlSCD6SDXJUoOthtCs46a2jFn37re
SxkNgilinrAz/+mj/A9ANXNiJ8AxG/+0/TpcY2xfVM+XpzvOWUN8ja82P0Vy68ei
qv6NJjj31sMVVdmlIedxhEBkhqooaY3cmdA4uSjMCLDy2HtT9RKpbdFVStX0pn5S
XLV59X7r6qOerefWRBWqp62D+HUmloj9YYkOCCJDT0S/ZhUplMbic9fDHBgB3UYD
M+JiwFeCrxXCxNg8YhZp7Vc69e0RsR0VeeFwRDpjnXwej1+x8Km25lLc+T+BJJGb
Sse81TMEPrEDNFNvQm4ylrSm9GW1cH3muvDZmM6SiKZ8Na8EdlAuz4Vayt9W5nYe
088d4XKtK2qJOllolgrCYBkmqge+zOcnNghwBkIl542+spEsNeSL7dNIxj6NQjhO
k/D72JpbUFcrCRqGp54RA1xJcX9c7+v7wRJY+ENe8l3u43jqs5OXucug99Xhxsqa
oZFXBwPgsLQDTbfDPcH7uPmsKFrO4BAe6+YniFjY8uUMNrJebhJH6hr6fsEjVDsn
dWfD5N+LxNov1hWPN5zaLr527lg6magMHZCbSAzk1HJF/4VQfve2hZbU7fX6XrVA
qOl5hxC7GB82xCaGesj1FAPxWz+gXbgIQYAvczvgLVlj6gala3ZfefGyQWPu5fnO
YbVzxvjlFc4b2oN9lqkbOm1dimcBL9ZB6NFs39U4D8G5b1qq5nznewfMUPbS3znu
UtYN+5I5TJ1owCJF3NGBBkpWBycGd9GPjLb3ZcKRX2/fRzSJQjC0QB7OUAmga7tZ
Cwe0++45pQ/ePXf4kownftDMCzexGpB6Nt8IQYDIYMGbjuRuXT0Vu4V1SF3d6StU
1bGoE5dBOtPOoqsuKrwElNIczA4VavL1R3IEd2Hlua+KMUMlaCKN3aaff7/bCLT2
uSrsi9NHUo+HM+RvgANmOAfdKLVpxSv2xraH1By+/jNjPBA1kjNWH3yNpgKEy0tH
f+kKY2/yV6lunTy6JNA4UdCNDm4YL/x/JQ4qS1l79yJQ8Zi7vcNmWlv5ddt0/0zp
L7eh6ogXzpIc2cgC8fONWBNt33llkyWJHWsE1uEQKDqyN26t2XTLjT488lc427yp
2096Ot2DdiftLafQy23eEvU8qx+5QPAePb3AClZsWz9h1+jCpJ5rdn54Az3BQfo9
GINRToRdjOabXO4Puuce5pSW9ySmyT2AdHSdMtxOGboFa0S52RyFr/jNSA228OrO
BhQiPnsdRK5dNaXiddaFQGSallAZaoRi+o5ValRZIw/mxmh7Auy968VnwWW2hzIZ
3OOHy5yn0b/eXpDyJZLV/14OAEw/Di0PNLd1D+R16m55lzb5VElvCrMaDhBFM8wk
DdiZRlxwtZxJ0EfdQoQpMnURd/Mvpa0SiQrOhFq3UVdE9YywG955KPmMghtCbuWX
xiHtW1iVCF9uTCMaMvrXPOc5pFVGsXriC0znUqWwu16WzWi1MU6E6KOPPm1WIRCv
b4yTaDflvC9GNQ4q7UlhZMSaMbzns6JAU/6mrOTXXZHZk4UmnO0bI84AXlnv3Zh/
aFcA+T1v2cGX/OVTwWN3grzCb7qXKklcgnrtpleZ2D/urbOvfW0CyEtVE2tk709d
cVfb25Nm0wxhDCkEmBER3CTgsaJTYD3jImbstaSmOOhnY9ywfb6JYpKFLcZ+v4Ay
AUyN+tYePdYTM3v7mBuu07TcPTGutr/PaHkHFphSIdQwkDLLsJF4Qthx8LwT21H2
zxXrpxc6RD5vA28ednf0gnm5o1Gpyl3VQIwoX5qoW7iVEgYIAqwlr8g+AZ3QUKBh
bvO7R3JxIpt+27ToeiA2xUJCPdr8wzt83y/+Okj4VdLj+QCN1PHrADPwZ2fQTm3F
2lgWIMnypoql/760ZZiws2M4O5fjsouh8AQyjiGrNwLiIhGuyTmW2U0Mr5nyp/NE
qsdWg0nhx/pIBgDwat0TTEz1zXKytjwbRFk0p2EqLTkH0gqXua3NCmcfIYE+8TA0
4IuTi2Tiqm+q8EjtbQ+Xr0ogSAxPcqop3mZ6ulrpJ0x/HbD+/JJ1tFbFo9Vr4fa2
gkdq2kwtHVVs6bmxVsJhWS9qN5Hwt4Yp5jisct/nSxmlr0ZmPxTV2a9MC2ZFaN5I
GO0QuUT+6aRr2KlsY0l7L5Yw4rnNdjjaaJGbp+akOQ5nsJJ3voBkqrXlY8NKvSzS
5e+pfoIfvTAbEDdgnJbeD0hrRD0vlrz67mGjA075WkV0GQpU9QCcyfVuA29OFa4q
JfthXF/WFRq93ckiDvjwDSyYF83NAd22XJE7E8nJk9A=
`protect END_PROTECTED
