`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXV8ZufSLIQY0sJa2bOZ7DB3PcDq5Rgqahtgrdji9fuudNxyNKAQelVCsl2/Yd3Z
jn55LXAawsqJpdEDqetceSmBp87r5CK0MM4LDadGdHb5WE30o3ISXlK3SbJrj9cG
qfp3qYvYNMG7gkT8BuiQy+wrWP+cruqGeUPvoODsSVVg7oVF23h6JmxCjK71UGfG
lwQPIi7thcO+Hv+K1YtMrrTCYaBEaI6ASYdAQIkq51SwTb33vIetlsw8xmcY3xfz
b1bLg0YGZRf9+OMY+E77+UCRTD2I0quHvm8zcuLobKVE5aCDeDw0uvLiKF5xD5W2
kJ1QEPt6usBukAeHsVP3qV9uefl5VMO0OTyP3+SC3571OtmWz5E2RQmdyoDD45/O
sNx4Jw5xc2qTJXq5U8qw6Eb4ZI611n2EzYm1AHtVqO0oXSZmdt0bzeUy/oOLSIZM
Xv3eBxdmKmPC4PYOEhjxfuU1Ffq0w2nLkJJHAsI3DSlzvb+hQJfQUkjXSpyp4EEQ
L3EAC3nlOFqUplICUahzQZuX+Z1d7vVCbssqE7l1aToUew0qS1quvJG2LykueoZA
Qh8/zZOkCdmLHBNKoLjAPtHz8fkLSZ+qzvXMU9M+zOTPjGThq2BP68vMo2KgfJzS
98xpfzvIHkHAi3Vd94jPcMlSJKrYB2j+PP4as+/BK24gU/rhbnJOrXqNhP9vcBEy
6rduuJsO5KYr/0lixUmZMldX7sMieWPMiiFu/2Z/27B0y5VAvsdBD4tNBrITOEJu
wLHy2UpbPoPIzCAu/BiUszcmMB1ham2bl11vT2YQF77Q3/rP6jyady2aqiOWjBFe
RUkgdWxVGJEIh8Ja5duyg8IfKWPu1HcHmZvgmBpZKvrLUr57N+Aq1iBs9CwBYCQJ
xTotHWrIavQiu474IsZwosJeCgO3zs0uLQ3n+ByvAY/ko6tJ8v5VdDzRAg1mgj3u
gAIDKHanEWDnuL7OQeFxqMNF8uF9byRNvHb2jucbbjNiuCQX/jwUQvxl1uBjcTvP
wAcGIJI3cyfFMcic7PDFqNW10GbHu9iFoZQxOng7jtOVPOJYZ/IvXg+LMCH8qJo/
WpGmtYSkKP+8I5/6LAbvkM2aqs8uvsHvR/yn9QRUsG8BpeREvPkMutabw1ErNC8N
rmmeuYhqIwcAkMitFZsTW8zBgNKStY0HNsH0L6V58uo1DN9oi6XH2RistIE+qpia
hn54SDZEqfmaAqhcCZmtxtUacp0Yjv0k9SdvIIZoPs3SCPxcnY/eTBILUULMsCyA
K1L0NR/04KCrIJkDqA75hEFa96D/yhtqmN+PCrJMwR2jp6U+Gxj0JIiQlJNCSDAZ
aows4suFu7XVmor1RBJY3D6VXX9wB3E59zYzII71tNKAZIlM+Ft4rk+/dSZfhqsB
Ege3NffN/6hBLMXpmuLzOvTJuQVqjVGeRCm3PgydWgUFfVMp0ix6931J8z8+93Gh
WbX1C/1/ppkgDvQ8NyrcRuz3nWVoylgKR+nPi1XZtEY=
`protect END_PROTECTED
