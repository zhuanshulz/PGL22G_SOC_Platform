`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F/my/NhoGDaxi2UzhRaMWPf8UIk9g+DpbFL7uPHqEXVP2ngxkdt6Wzh+DXVrUrBo
yT1Ji+3L14nN1QWCcwcOh3iucDIqCS2aNiDnxiMg/6P9cKbb9F2OJMVt6pQDyU6+
GCOHNR9vuVWcWreD13dmavNNUuxcg/Yx34JzXSuC4URg5SJBvF076UNheDoKCUZB
U8VrLDTDBxe809fz8o+zgm7ejTbEt9L/ztRX6WG3OoQrY9+HrRIas9zUgYFhoW5Z
CRdvSXScHDLVsXhYxHTrB40wB/c5mjBbHRXFmKB2x23t8QULQbUqefgotPrIv4Ke
VxCtQ2f3wshlpYimLHGfP3FxE78fYL99tyc7XViFYucnm0OI5acx7v/cIKBylLp7
05euAr9hdd+4aq9IRjjfpTjNM0EhQxNLqXlYZ8+yxAi7znKusI3NvDdNlXY1Hc+x
dsOqOTsQrx6s7o7IuhhvDXXAE8mPgwjOyBD/6KvZ3da16yUwL8d59jRf1934CTTH
iogZRuO0Tc1CCCyyv5+TbI9dOwD3KbxpSdQDevMZIiMQx6Aax5XrRB4mv3YRTLCd
`protect END_PROTECTED
