`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nd9YTiy7JoPy702HQXhiHM3Bx7R2384/98nURIWFbdGC/VySu+n9TODBWO8XHtOT
Rucq/OwLqnVwNPy4/gSZzdrs9OD8uxGIc2UnHT6EEa/BIG90RmZvaRvAbXJG4X8S
V2pJ9+9g0u9EUdVbOeGs8ZpWfuie4CL1UxWkbbUffKRCmUr4OQxHFS9eD4AbhNHr
BXpSK5wUaEKzdx8gjHzyS+tpB9Nfd+Qjd6Oh/xC+VafVze3JOMqwSiGGsDcrsViZ
Dr9MwUZtsP4ddubpSlJ6eElQDPoSJ8/9wYKsBbelWeWEahXattwl0FsmRr3p+id6
ygShYlt6/o/8ibpdQalDMR759ujbPPD3gBrZq98oRZtTwIVLGWN9kAWrSaC8ZtOQ
r7F9RwvDrNzVyKfQ1NPCK77BNXYcavFLWOs3jeZVvbsri5NOD8Gl/TfohTGjCb3E
UB2EAb8WShG1JFUtgKkUfSk31W8mydz9M2VOWU8d7Lky0Mio1cF5mMtdp25SdE1l
hrVtumRmg/gGslBsFfiJ4OQ2bwzHp43rP6SAXNjus08B6Q1tvFfKH2FamIm6Nx28
IqYhPOLdTwIdoncOZnijhQ==
`protect END_PROTECTED
