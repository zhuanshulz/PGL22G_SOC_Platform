`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDe++K5aN3KIlaA8dHs8SXNPUzJjAgbIqdcS4krFK0EQ4g0QUHkmrdoeIuI7hFQe
yc1VL96Q5YsKMqbx/W6GpX2xRCzvxdLXvCHzudO+wjdRaHBMMfl0hJi81xdw9bdH
hscJ63vMpaeb9Rcxxy/gTrLAg8I2y6HJVfZCbSsIXvNXiT+u1Br+pmPnSmf2Od9+
NL9wWixJrOvEegbUObuFJma4m+XrdNHNOiJA6Vp9IHfSt/v/xUoiKxLiBtRGdLqm
L6UdDjx5/hrub50a9MrvGDZ2AHIeCAAvJI715Bjt5Qa7W2b+Z2+eCjcy+GyoRU1l
RIwfr+QoVsfGngMSoHAeIA+raxCzcaEHo1WWr8TSyTNyRwaB7gtB2JQMFBx4GCpu
vrTVc/PLb6noL/EfWNxChbMdlU4CJ97aw54LMJxEpa/StwRhFy+lPPsOYGcescfi
SvoSR2NTx0NEAeJC/5BVfU8DtRucg8Xpg14Hcdi3jTTiduB8W58xFnlxwA32r4i6
PZegM8WrwoBNEIsyr9gLIp8QtZXWNRvlmTeX//lRXPL9hZgL74zLLrDKQuCrlMBm
JKvLonUeqfAHpBP9gCOhlw==
`protect END_PROTECTED
