`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
va/uo8wvj5YcbW5uS9EYESCjrs+mhEIAcqSNkR6faW47Z5Q5LoS03jQoiujNtw90
EqjvFpH7GTxKFvEiKQiSiLTepGNudESAblMbA0nsv8wWFfRmE/TmB22kAid/T0Oh
gNR1NcaY7yDcVHG5gGg7xOeHb+BouOeLrV8JiJXGWFOtLBNkS0AaFaP74MDAbxQB
RVNpf8o0v5VGEO9n5+Mlx6k2/EFDmgCOW4/IShpjeFylvl3bl554UwDbsDxf4Nxc
iGzmQ9VLdWRnzr5mD39WYjzsOF7qvvfMzT06tfo2uaQw+QHat0CB/3j5kiei4we9
OeKus5Jovk/xwgC+2zffZwRi/GyfBC+efSsKHd8KDVmS6zkX9uLlDqv5EiJ7nrTE
v9kNgpzwrXH+SkHy/rbyK+tdK5BIepMaZH6oHLd3R/kxCwAz5ko1unPN6eegarmG
`protect END_PROTECTED
