`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DCUcI816Zh/RUIL1/+50Y+bnZOjdudxvmXX7BapHnVy1J5XKYBB+qlcSwlt7G7o
FyuJwBdFGbC4H0/wVH/wNKSFoh/8iZAf3YAMoX+ngVT5emCUqCUVV/vXnj8FMGMN
dWKrRqLsaOivGhJ6oO0b17n8uBgTiLfdHqBjZG2mL1JaMh8SsC7c8qy8k80jx51A
hySAorsKjI5p2UEzoYgaZmtWRpdkSbYrmfU7oYbcEZcbB8VfTP64LR0QvM+BFNj4
9IxE2/y3q7fjVgppJaObFysWT6MXFoBQ9hIS+37CYw6thNktJOEbjkk6AOQDqL27
LslInIdPqU+mAxlmbFEsB64MTBXv/1ZKu1LA0Pmv+xDnndZxqW0tKafWJ6yp6rAR
vLL5aISnn7Go5hR+o69G86PljXD+LVB79ge1bbASu2YVWnq5w7i8RqXHsJSX2Mya
wl+fGg/MqTodW7+/6klTAO09E5yHn2qViqpsx0GwRWc81+H2QJaTBfG4zqB4MVLS
b7cuRm2SBXf4npqYCVhHkCbMlGKxJIR/S4RH+rihN2s=
`protect END_PROTECTED
