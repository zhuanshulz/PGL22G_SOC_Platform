`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hm9SLPW7Kop8sbKthnNtxJGO5BQp0NyLTkpQ7yQg5Uz7jZcwPQt+V1B707mzdggO
T4yU/wEmX7ly4mT5ZGP7UpC6Onw3wL9gjE9H6x3x106hJvY6d5qx14fdW7bDNBWK
KdpijREHnredXyUvYNKITRs+OIhJJoCeS4FJv3RPlDbXIdHxokFa6kShRlQvzG5B
pvh7X7f3PAns2bRRRK6zFDMDFHNRwhy9CjKNOYQdtrDJYZzYcmKvKtWPkTT43AGn
OmYRq6SsQK3Skk3Gg2Ju40+deYgXr+GyPwErViO1lLf0b6lQV7Q2O1pyU8Juio8O
Dh7RJxSMPa4rMhR3UZQIVFTiquIpR1GcdRxpDfRklT4BbSZXJgmBIDu0viYZypVn
3VZsTqKD25cUmbZWVZASKMgdkfJ8wB3DJIXCDTvl65Mgb2YrnBihJW4XkdWFzpO9
nEPGHWhtFCwF60BGUiFTXi5oY/aqz0P8rTCLZyAsnjTrXCn8cD8demNyI3LxC7vd
a5/Sv+IxT5/s82qjcdu9Pb61s5r/+yJP77fw6yW2k2gLuYAtLf5ecfuMH9Ul99UN
oiCT1hLk1oZGhEiF2d236k9/v4wqaMA2eULJrAFwiiKu8IBosZfsiZ93szrJGQ9d
uiuHFrizSiIeKYtrlafMM6QrNG4VtV6sIxl67lgx9xfNOaH1mFHDgRQA+HNNIH2a
pi+U+n3Nl7X9GcqT0rYYdE4ZG+JyTwIs6E6ILNiLSEIw2RvOtI8eJtmQR0JfpN56
4+G6bS35ZGQzH3AsJlI4ESK7Xico7TTOiUP6tIJEBvi0XtisjlosLHMW98lRX2B1
6/IQmorikCjqeGJzDDQk5SYRjyuLeqagaf06Yzo9iMwkbuqS91ku+W5xBE+zEGDk
aTlJqiDxZWfWNrrCF3dY9R38GyKW0+ySqb6C2cKQnJX5YAr5nPYmFOW0rY8IjEnI
6MkwybXc21bVNqO3D8iHl8ADsPdTaugHzLBSQrEficv1ip30Jx9WX9/Dw2Ga62Jd
BGGW6H3KuNer+LPoApozWGB0TDYAPCtoHLfTJY12V3KCpim8kUyFeH6peM8sM3cC
LE2dkxLw4c6L943Q+TiV/dUIWcu+MKUcE31guCxMyJwoxobxxKStR11hvhqXpgZE
FZzOpDSXQTRJ//26KyNKF4swv7ah4I2w4w2bi/6VPPimVSxkDiGT8F9jarZK7VVa
wrsYMk1NSu5KCcNJYZGnyV81Fo/ANZG2igc2nsriXIlgKrG5Mt83PfJ5G6SRdGo2
DdpyYWzCOeHvstv3nFjhnl/1FfaRAX6R0HLYrAZhWwf6EvCNlQiNtJ2uphlhcSiS
1QsrMu+ZQqajznrNaWLo8Hj2h5vdpnUAagRvJ9/dR4Jy5AmRxR7hvnWT0tfZsDO9
btbkev8TNxLV7ZMEgi7BlSgIgvFVpiIB4uV3iBOmzbzF1xlLk0zygtvILBNDvDAV
7h7C+zQvYtF6seBWgibgceZlkx3f4hRFR+Z+bDBW5N0KtnSr2bag2c4E0FIecm1z
chYFLG89JUVjIJBgk/SEQtnZz1y1APQrt4IeBN7ubMsDjvllSPFsIVLSibzpFVEp
q+VpmMmKz2m0sf+V61ykTCz5wxEDjLfwlovT2CWA2BAKofp7H6zrjeQNrWxkEb9X
a0c12JVYbuV28wy84o+Q6jU1L1SXG5a2pGbwnfiT+r+h2E7wgk/u3RzEUkvlE1ne
N5zmCieVQPuq7fl0/CNEOVbJ9jx1FprNlpk4Bzm//wQNzNIQoC1W7isQoJUENBKe
iWITwtoh0QcK/HfDi6x8T/MqMvgvdtsWjJ5t4C2FB6EcmhtaEyanPG50J4AJRmxT
HbuMOzziMZAJWHPS1ZDnMa4yb5/+qH06090tnyGAVmHE8m6omE4mZ744zQZP8Q7F
2o416cAMcXzFMlzyxhHqzVdIvFHGOKwFvhLKwdrxyu15pxrM2ql3Eg6dEQptY8/z
NJ5dbBsnLgfZHWZwA1isd3q5iqZl3kztoCdBnAxUtYHdH+FHg5UlocW53t96NIYY
vBKah3lSbNJt86ivMkMYJOZxbLxBgFbwAoPg0EOlAY4LFC2vSOCHgZzklDsS0ejE
AZDV8INbr56xkTy2bVzq95tgZfWNv2gF4iSqfeQdHdJ/2ku10CVdHQl6gSgqi0w6
xctduuXJLS/eKOuc1qHNcDPmv4VA/c61KDAj6yCAZTy3saSGnOTFmcBfEAPD8FfL
1wDCtdWfBXq8caMbM/Ib6UHy1Lz8NMx9htz1yLb1Ip4W7yU9YkSepQYkT9fvwutS
fhfEB4/LlRFxHcfizB4wwOzqeX5xXNN2qS7TlFPTR0iteSwq9qL/W7Y16JghcR6w
XAJML+KKOAYsl3TjpaLW5B4ql6Ox7SaIAplVZKTVchKfGg42RUaft1I6t11RqDp/
EdBXhuR4w+/KWcI1Z0YIQZMuGkdlyU+u7YYftMpuMkjMgluh9sP9Inn2lJ8gXEme
UOaJIAoM17NOyuosnud2gE2OEcbzUL5BvgI4bJ5T32UCx/cpnLHCCiWN2JVR6og/
iPA+dwNlDnIDmJ8XrbF3GjvEdRHuk0H4vcYDkfuUYcSNB3/pRRQaHPPyOu5s3yKT
ehWlFO3Y/qa1Gpc7xza7UyxQyTNtx2u/w81H4gh/Dlh1T57YDZeYcjrRwvQZPbcF
SHMyewvYMilSFPam9MeTTJPYQEtBIkTlGwu1V/qmr6o1C+OUwquoGFo+Fk088z1s
XgNO7a/nz5/m/BitaKSd8eSlHFIFL0g7WD85v0bPutUaMaYSYM5ahb3wyXiG2X5z
pobOj6MxRy70doadzFwwpjpRieJ8YtpVP1MApYB5YEcu9Y3285fHUDeWJPELwwVt
kbXyaAkmhXrSLu8BfXOXrA==
`protect END_PROTECTED
