`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4JQ8nwPOyDY/4tLHYrhe6Zuof/mzQBdSIA+r6jBu8N4SF3jdYdUsmub707zuvxR
p+phbXK+X8b93FrMX8I0ZIAF7TIMqcvadLzBO3m6NoNyckUh/NqvEyu5xO+SOBmh
qfiEx8UTQ2ezrGXGzdMp9c1to6PYQrfYn2df0gpQ0mjq+JmwGojfQ3z+WFuhicD/
8bUgOmp/MNXTTIk73bxT/rA951twFmGh/iTHQaubyYszTSZK4+TGJi3dTNiTCAMv
Bb6bhFykCr6LBd04W7PIfrTjVx98sGsObvWInJB/oKhtL3gtVGx14icYpYlbweWy
PUkWcAB3j8geU0fBSOXnA+0isrwdfmfa8XOXRKvRpBAHpsp11KNqH6MAbFkuPHr7
nlQWKP7quZSZmDF3enGJPR01IWHHdwiijyIx9smKvHrZZxVrwqTP3zoMiFerB1N/
FppBzHW0/2kRR08PKE1h1KjcfHYgDHoSAZb3TfEPECwAz6zImiaYKDjRoNmMVrnv
if+gvLgITKpNmosKW+PalA==
`protect END_PROTECTED
