`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOd5OkkUbVgJMLsYNRZgSuNHrKDjrnzXBlqkuMOo1Rw9NtFMAaIbfP+VZOoBmmJJ
Imnz12ZFA5YxUlG3Vs1GnM9Df9Osq3RVFH9Pa+ZyJYwU9qLAdAsunXiEVw5KvjdF
9GwyCJ+tzKDtzK9DMzU/RqV1EIe4U9SsEX/1Mp3Qo5A1O12KjLVScFy/MVsKByCv
OhZBk44jzz5dq8Nys/A2Tu0Wsoq4mh6K6bn934gRtTjs1wYQggacDB1firyBPLtB
owOVsFNYCHv2Z2Zkd+AUdPlhiaA5r00EqjNg+jNckHfnysb7btHhtFJk3hAAoe8C
rlCiWglhGi6W0beEoRdU3RAlNiNDTp1vvMPdM3QLh+cZxEItimRq/AUKvZkLQkuj
TRjSGU4vUGjz9OVRaoz3x+YTa/4/N7G+Q7UkV/6FZ4PWsX1xqmgCZu5XHyzshjkA
TgBaD72B8YBWyItNIverFj9/ovnq5JOpIYQOO60N8jDVQdgzttD/nFSmV6ALJcZy
rIg4xoogN+3zXHDe/GxjDLlWztmSYM3buX35HM7ZdDqZDvro1vIHsDizq2AZtM72
tN4T7twzxlRjNFO29vZ+rQWA3gWG0FZU/JZ9q9Ie8MPwzf2qA8lumzSMng6IMb1Z
vtf6yJwSWCwvMBn3Lj823GodkYxdMaKwZ7ukfMeNuZkGRjLoXJ/wDAxmCmHLWUrb
NGlqEkqiwUzWW+2S3c0zr6RoTQaIG1Do1IZJZXDQvRp18lOphn6EEa8weyc+Dc2+
+cro5Y519BksxDrdrH6Ooba2OiLc+YaQqndwfQ+0GhDcDcU9HwkrSsEKrU0CLqLc
3LVoYsR8yx3maSb7g2XhVqopIhyD++RcAIv/+Gq726A44MCo7WIUK+TLpdDhmWFT
EpUyesD5XLu9Nif0qxydYTwWIr8/R+oahThWeIBpACIVsTcya3oYAilEcI4JeErG
NeNFsznHRzhuDRwPd2YDSHtayCd4kUYf1hyyCooAqy+0V2CccS1YFmRfHM2AqZRs
GCW6EblRKkTVfm8tWYjvzNVejILhb8DZSPzU0igQwlq3XkneOxctAI8DFHeJqcWv
44FMz54ggEZELyCaxtOcpii1EycRUrK2iQbm8b6Qzh8mzK37VIowtMLd3FmmB6mC
6AjFBnO7vQRDPTznXXyAg1HTN+rIsPq5my1SRVe5rfko9VhIyZtWncxXGV8XRg9N
hcc1c0GGAdgMTbo5qtUdZqxccOEgf7Z0iZH0aLhEpej9Ox4K/HMNjfZHVuN72ult
szdonGI5DvRsD0uWgssEA531RgI8oNPuGWojuL0zRLFhHaJJmovC94cEmg7T0rrW
Gr5EvHrgNJKU1IcLy/ov+OrIbEfb/1MgXoHVfYY7IAV0kG0XPliWofi3B9cjp89v
23sU4gbHFz5HGOaXjkgIlLtCRd4QlQpHHJFitEm3SXjYczqYvObUt1zmvpXABER6
VjrYK0NvTe5Xt8UGi6Vixfw9r9d5Bw3OjqoD27QTDtFDobDAJL+BuEBadlt58KP2
I9gSw2gI0FJtv28rbbo2kj8p8KN3m+6s/h4ysoIQ0TBzTpa7kKrILogZ9FhB7bi9
e+1wE/el1Zx0+jzNPfMq+ni/7FDO5kIvxLYEn8/eN0EMknI9P2G3GXfJ+7g8AzVU
9bdwDDxIJlYbbJfd9R8kN05ZgCfuax335uwUS3G08Hd40fjVvMEj9hO40Ky1jVzl
SKAIe8OjNqXz3zyAEB0YxzDK19xeiBNl2GJPKCj9PFs4w3UNESih0VvK/ivD8NA7
WMy+qMPf22qMNyqX3VjpQ05VUsPXEm7L1KWzKtQzo7+0lSwoJSQKqH4qnfzSkKCX
3mDW8zfqEB3bp01EIY5MrLrYs7F3wbt0NPXliyn3vRk=
`protect END_PROTECTED
