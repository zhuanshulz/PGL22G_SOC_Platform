`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QbCFjUZO16Od4ken99cro+ZmAf9Y3nM8KZcm3tz1LSn1y3R53w5uTAHZPJlxPtxz
JEWbLhAoGTmPTWfTSg3+3ZEbZ0WhXZVYfkFpKsYXs163eByrJYaTLHFCB2siQ91G
ksx+45vKn0kLO90vwkUffiG+1arWlkvTxhYDSrcDwEFhb3P0di3OzxZRpcPDkrxV
kKQhKgzkjiuMLiQupra0ooNk61lRva2uAIIk5Y3pkSNcBEnwUHXaDEpd3d0Td0IM
LoHkSj4j/Dxnx2V9Ga/KNxapzEP6Haf+7QE32xeMwr0A00yAuiZQ4gl9gmbIXXnl
sT1wAen0D20eDGNyPNN090gP+98lfpWtkkMg9JUXqZFXv/7AFoBHEqoU2oFSaMHK
X3otLIC8ncoWJhNRn61ZtQ==
`protect END_PROTECTED
