`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPEU4CWe8gOcXnAsfJCE05FwEBugG6cItt824zrCs1kUKQ0Emoqo0jY/qUaenHcV
MUlA48iI6oToB2K8JiHFarQYEoyRLVUcO47LjZwJeXADqW4Vld8Dxu1GgZQk6kUk
IMhsZPqPPsl2W/2etupVQyJ5w8gkAiZzCUGRBMMheTGTC8n2+pWRqtli4vwG07+J
5TGW3tL7DJ2gOI4pbA4t4eM0u2wL29icHdOkdvaYrWHEG7znlnbETxbdyamEfGfb
h73/KTPw4923NhdzCwMm0QPG6HjuuR1MDRIO966ou7awQKhpgu5HeUfChJH/9pYW
/6iIK1JR/lc84yiHDo6ZvIhS+Iq71ZoFkJrYFE2cxNaYr9fy0CkSrKgzaLXWzDQr
j7O0wozK+QvbYqvV9mKQYZy03B2/GF4sqCBBlL69J65vt7WqdOmdkCxJVFWQHhfb
+NukAu7cTLCxQ4Vq1R/soQIm5bPmHKKnVz/6qOIZsVzdlgsR0XLJMQKmaR6Kuo0T
nL0GTLRCEek43ZO5mPhiaLVwqVN6i+W4bF9VM11QFAxIPOhspCaPjn1bOo6hJMi1
VD+K7HC7XGyG8Dn+WX7WWAyWPtRmaFNsmibulDWmy/cgl4DPa2X5rUjP/NK3L/HJ
`protect END_PROTECTED
