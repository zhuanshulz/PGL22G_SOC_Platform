`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lVpY33cOjS9BzZq3A5IbfpUWHYgEJ3rUGJ45CpKfJL1uUy/lKj5PWZdi+IXdumMT
UmJgDBmp52VfeDDbx3teLhoIQ+Ly84Z//kHuf4OSFMaCwKvtfPB8pmwcSMLe5GEQ
XP4EZeYydc1irQe81smOeR4Go/mg2Lv0p+S0lZRZfJLaTBV5KD9F5WBHzyT4GknJ
8gZEuMOblPujMc9BQMDALbKfBwBi1PFvJiZauadOYH0D5GrV9I/jDpkIxnwaGhkt
4OA79iS2hHgTe3ClDRW+FXq/c3Fbh1tQfFdXpZ0TB/Hbesf1I+Gr0o1AZRTgyjgX
/2ZJgbl2ibrgVi2Az+G7C8deYkvvT6kF+L0eSuQ/0asqGLnQEsGpD4hkop4Fa0vU
Qd5E0muFkitn1zHPFOx0QiBl5MIPRF4qc4JEPX+NjNGneb9r1T8dbDtBjS+uQcYo
yAL72amKtRrNmSzxC2BxG4WQvAQtvMIl8KKTqnD+ZPjxtefybVI43CEAAIonmUOK
6rKDyndGn4UDMuHl0M7R8XsLQd699FFYlU3Scz0ZIwyZkqGdVRmrF6lTKBVeI0aE
00TklPyZ8u79sn8WLlb4uowohzrBT+b2bxHJxNDU7GjcrfUNMp5Y/yZNeDqJjFnb
8DhBRSo/7L80PmOYL7DhCJEw4kDvneR7rudPI05jfiaQrPISu/iv8S61n7COZNau
AWH9DuWWyHecIN/vizFDojtgce/MgXwi17CKUn9zNbCKpyWzGXsQ/kB5RE+W/Emi
o2Mp4v030N1m5pGfZRssT66r5v9dfuL532Wjry+u2dSI/4R5pxbJN38JPJoqaSMV
Hu6MTQKjqJLJ3+ggjIH1s6xuI5OvFfia7vRiXykYMzKboc/vxiMUZBWLo6d35Vsn
kRjHDzbkefflswGwPAQhg46IOKjrQdg/7UplU2g9xE+vRJYFrQlvy2qZ8mU7AiXa
Ue3kh8VUOLsTwVkuhJBld94hzclhHKATHMN/jj8TXvuCf1gmI7EgwLGoBXt5Ct9S
zoB0LVH/YoWAw44IUMcYNxpXuUjdQPfxMpX3SeLXSAGCFmsKMUIkcAlilDwcivnE
uQ4Vrm1NrTHuXzX8RsMwAVOjPEImVPt+e5m2Fr6IDR7FfbuInJLbBbj4wiEsX+2p
L47Nsx71hnREb+p24/jG0ZfpKtpcEh0v3sYMX+HasxbnhKNs5ddbFiBnWDWaPrAW
DMV1vgPoghF1Qqkv74vPDPnptuCzXdH6bUS7ELvFgQ5E7vbwLHw2uSJbroQiYNoV
Rt5UovOzs/nJbYScP3NUVdVBDg2Qm8u4HmDJNHju6hfd5pI3sx6g4VguOcdM4qLk
vJ1SY2Gs9hyVgYDUcTSFlVhge9g3YchBrjuL4b4lJy1rxQ23cqjsHxeth+t4/TWX
bbthcVAdoLFzk6kNRvnpzYh+X2BvgmrctigXRufWaCYA35zdHWfJifKkKEI+o2e8
4+8B8gPupomDEmCzMpcKJHdqVo0VeuCVCMfA+jGfOS01IbSC2E+NceRf2cH62zfq
w510KQOXFPq6nh8b5jgXc5LwpA41d/XQlctFazyozFuBwOkUzZzyuJz7pphMOXty
C9NjRqrvpr9vI3RtE/+Hw82wq9l8Ht8z7+rI1HCiJ7Vp9fKE/m6GOz6gJhFB1sPJ
afvi+fyck0Py/sk2nZrsaCrzDZNk0WiK6PBlpANDAe8=
`protect END_PROTECTED
