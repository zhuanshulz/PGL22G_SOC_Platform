`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NrpvvKfdM1KhZfEpi1eiM8PtUoXNRrR0IkzMq6nfBx4R+8DDXyr5k/BZKuOmHCOh
/sMAWaxOo1iRCo+ErXL3+EHHA7GeFaxEhxTRPtXdrfrYHbmuc94UDQRPejSYhu4Z
z4I2pNVN1G5fuxrNOyYrtm+xRido7uXKPTujtMPTNe+nKzGTbCm15Duy1U1gAUE8
13J06Iwx93r5yPOlykpd9bWD6L2kHSS+zfyBlnn8pSJf4yw9sU8UQ3nHbw/R8NmN
8xODnE7g8ORDjAAFJpc/H6HyCfoYmZVP/S9mmmYu7cA=
`protect END_PROTECTED
