`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tt/r0WlAIPODub2M+SWAadjB4vWBB7Bu6zjW2P2a5EltFdPY7kj8PMEoNRiRTAhh
6foRnWvDkUU01PzLzq9nWh5JZwp59BkNGIP6t15lSVxmXcT1tRvjF+YzIW8Z4OgS
8aWCwLx8erg3R2QYNbx6PoiBWiJCJ6PqkN+kbKP76gSaVO64jtV9J90bmgn3/amg
IFAR1otd5XesXUhH7YAzHKTqdx4Cwqc6z43wbZ3+J7EdmNCp8hXhaSwZQWFEaV+v
0HkVcHcLuysco7dvzVDebyA9ZfvOw+/9uBRGQIUstm+YgUrwqA9cS3k0eixIYyv6
iefwgppDYDp29h9Nu/d7cCD0LDGrXNFnttVPNdp+Q4SqkAUNL/5UT2cZiIIpYmRx
gFKyBCl+1riFHhjGfrqsq7H+MvjNoQqF0/Ytbz92JJiYGDahmUBcFVXjfSAXoX+d
CZ03Vjp+VAVfbqm/Xvu/XjBMm/o68QmUTTkyLNIgsTuguPZt5pVcFoFXk2bFxdcA
bKgCQNz6t2SSLncycKh2wIkafokdOUH2wSRTePvmYC1J0HMSGeF4b4DiVq46lqMb
MHrEEgS+8ZsJAfsrTPF+7Pr8RHFArE12bhYMfeGM1JqLre+HPRzBpWuC/u6zFFqr
yPyJgUo8qGV115J3bZNowMR868plk8iUcEISjgkINUvJ1qIp4AD0kLbvsHP4qd8H
AmIjIJ4Ng/WCyHS5LfoNrl2AydSBqL6pgNjObIb0w3xEAIB3IBm5vY3d7ws6Wn4H
q3z8vEAjvPXjcN/tTiSacolAQm8Bsp3KKVTAZEGweqh98Y/U8clv15H75AEmv/xY
lMkenDNG7Ee/tLVvC9E3O2o2pk5cOFWwCw6L+j/anvNtV/1d0QyXqCF1Ly9+N3rW
2lvSggSqeY3YeDq2oWrzJ+SfHy3vxSq6C9ZGjFz6zWqykuKsbOI3BbGuo+9/VHpn
DbBXC5bncw2I0zBlgjqafPZh9xdTaaQa2adH5qiZaTflTck02GZBLTnEhMIYe9Jh
XzjQQ3o+Kj+KcxOmigwQW01MhBDJ9oQiErJWRTja7OeSWOULDAPmqjWzD6T+yrkp
3HcZX2b0Lz4nwPjr95wO9pK6/ZwUmOqjTJ+8XtXv2wOQO115KFrupDVSK8McUlCX
Ky9ps4ImSpKEMtW6YLTYZQBgKsFao+UnwNPqb4cfTUn5UUphQ5tcjsVEz1Iqw6oD
bpFhDA89nfbz2NQLyqR4vQtoWFvcWjp6EqYTp9nXfFrpUTyxUToZMy+zY+sCgzkO
7DbZUrG1tnX4LDcICxEI8q1hnjbtIdKuiIJ25MhSoR2VsqJLA/NEaN/sgMtRIC2c
RaiYT1PRQpmGYWMP4zUcLD0GwL964hdKsBYxpRx/2mXO9sWv6V2WDnZjGtcuZSee
MsGbkUIVi+A7RVWUvLi6LgMLOFTKorucVQzQyMZtp+jKmm6zN4/5KYNbyXGNhwqP
IF8Se2zagQHnSNTxczdoUOQ27fXt65UNyCyW3tjuBkioEoNVQJl9g2cVvKhDIg0e
LPbI3v95DP/Z+aRUFu0DZNbxonqpg4/iuQjhqjyMaN/Ds6riH9UTd0qKj3x0bjiL
SA4YpWaGTxDZZciLygaW0IakVBySmihfUlJt98mbQ4qGAy+hmDibYYEK6+1SsqH2
TeA65fqerM2ER84jPFlTxbx7XWXWQlPg/H+hKJOVogdHXGVjtemw/0gZp2p2Ywml
DevYrScb9EfijN1+owpXGjvDdLv6B2wt22E1OU2+6JHUKh2stIMkffisD8O8RIo4
67JwNsIXcTAcrivTCzaFl+n99U2vHAbgksKpJ6aUWHZ1KTHmjWBL31I/Zffh9jmE
axAqqRO3ljt35kOMg+nUMILVTgDoCXpD7iHtEfnEqJNo1gnECVYIoedPTA7vpxul
x66s9Kxccrh9cfQKROjoDoDnEybMt0bWgzRDshQ9SNAr7j5TIdt5IlnYBQmzuHt/
MZJnG1gvc0ePFbbdO82E49QZ3cx7c5sJOFvrhD0FB6WQ8kwZSWuSJvmMqXtr0+HU
F2rgpL5Zwcvay4ZTUQqmqOfDphzl4x0f1+zxpyYHWHrsKue7M83UjAs4W5CUlfKg
oYUtKGMmmo9K4obOB09JmXRXHFmhvo64URBI5a+vbW3h9EadBZ0fotrhZGXbbJ9t
SzVlaL3Dp7D92K4Cmj3WTEVx7gy9lzXxOMhNd47+jG5qXEs2unssCYEvGtD4lNGi
qx4mR2gX3Lg2iqKCfjHxedaULq/MrYUlaU4W0j+d5Pe2FqRBOgAkRUjFWrahS3Kb
Kz46BjK891DKCl+yF7SJxQSL5IKstTz90KWaVd7eWDEiAZxfpKL7rpIulM9Aqq/D
Gjy3l6MBIdGuYoYpQyzarEO0QoamePbr8s+z/Q8GImivsLCzBFDtSc/rkeBwiN9o
ULTSgGHTErFd3XOWrd3jF4s7E9nYjc4QeurxKCy0PXpGMB1ZRiG1fTfgqOgw0Rx4
QfR8zhKtLFSQqBwnLwlfdRQ6ZrezYr9HwaNhp2bmZYBCOt/uqn6tj+1z6FNccMue
juWbBn6rghaozjIxx/f1Mfw1hKatnP1qLAU7FSc+3qVDvGJ7izMN0VCBeX1bJIGD
5cgSVes2pN4asqwJlA0o9TmENM9CSGTQQhI0l2J+J5jG6djDwIysDKBTxW5d2V6o
OiOaY9GzM3CZ8r8axGTL6PgSthVfB1GHU8ULlpUiq3+RKmJ0PRXkAFxdbZ+syGWQ
zCzP6R0noBzN0wxgjCND6Jom102Agl6c8PQMRM8R6kC8aUioxfFq0RW/pW6fV5un
sKv3UoZuPnIoTcwXWD5QvUZF6TFuFQg1RKxQ5FIcib8GCdxM2IAw2AnpQRlq8AEp
rNiPcp/ULxRUr7ddw4hEFgY2eYiZqzb0L+9zOSITY7LJB7QDO6XACP2R6qy1ARLd
cKRzEkXj8loSg6K6PcJjFAJ9aFkx6mK8s4YgOc98/bodHayj3IEitxcbAGzpq2UA
6/vId30MOAWrjwrKZZkSLBMpxRVHRFwuQAI/IlHblph+7ILiYVwQstRa8xAZpjfu
lmNdd2DBLEGkTROsyK8olRtOjnQ6uLfVQXoWDXbi5GF+n4kKCUt9gu/n1VDOnf0R
bWElc2MtK8QVG5VcyGhpGTZrxtmmhJXZRnwnXpFyBBtTAKI3SvdIT1rYnAhgeKeF
RpaaTyNq1wQ11TFrGrBL2ENT0jk+fAmjZ1zhM6jwEv1t88SYEyRQYfCMHp15XILe
PXZWB2Ko4b2ErAp/5tGuf7lgtdndBTL+zzn9N5rS0x2YjsU9ajdsBUA1Xkp144MU
TNkGZLaRcx5YOwRMHsexdvApPxZbP9gn8NnUKyJmzk5ggEBBTeuDQakux1WVadLt
zGaEOkLM8pxeWcwIyJxOm9b/tt+2WEOUsCkjXlwi4bz/u53OX4rJPyeGKPk781M0
5m3+K0UbKUSCdmPeOT9ZBNSGc7id1ErplX05TnUnK0339DvQyWGdwtBGW+NZU4Th
r93z9MbKB0+Bs749aEo044OqlQMLUe76d0MwXBz/q6R0/wt+Te6XVrGNw7/knnda
DbWcCX/YKaHVyFpvzqBMUFsilZ9EQTKwq4Vl9/kKRM3M8Fz7/GIvqnc3QO3bslTU
K7pvIvZLNe/DD/spGasS7zt2Yo+wM66JFA3aP6q1ZJO65lNIDUBBBb6Ho7T+cCuz
nPXxSXvXEpVJWHCXW3TClcqa53qlU12sy04136oYOUyqENSAGkXIMAyFYdYIIqJB
GoqUDezd5daa3bgl/wkeSI9ZqSYS6ZWfbtxUVz19RS8HX0Hz3HlOT5/b4W5Z40l8
nMacEdrk5ouR5ufRil2XH12mnEIslnGcYxbwaUcrF73ryuVnFCuJrl9G7jSq7sl3
hpU6R0gNefunOy9s5y3BJZcU4+K+WvXH+6bryYyFDM/c3rFHb+9nYPNVSbMTgKzN
EjpsGXbxJIf+HJ4I+Wu29IOGiSVvwb449y5yvwPAMbwmgqScNGCrFdbqjP/fxAsh
A7ctPnQAIv2c8XBz8iEwzio7xsqsPHtObrZcks4xd8T9qiHNsqddy0+568zGwgA+
x/wh5B35xUYCk3JRL/u6h4TTwGR7cXjiVYcMuGSH6Nvhvx/2wf/c6uaJvSc1YJY+
Y/gl0GAxJIMsH0o1TswIftKzJEG9hdmSaD0N9MZ/WjfNLvS6F/pHKUXk5EhTYfSQ
UL6SP8lTPA9oBbW9xz4THpfDCV3Kr1+6Z1z40RG9Qqfgubl2w4jlFgCdTlIaaSMJ
EBoFdSJijukJHp7BA0w3D5pSobkIgx2J9PDkRMMRlmUQ4GQVvWHg1bcE8nqmfF7K
vzeKH6i4NzicROK1dF+SnxET908FeNH0wbvN8dzX1kI5qQDWwkqczElxlAqKbbfx
jYz2G4rcFLm0jVlukw7LJdlXJfvhUn2AGxXoI416xxVzjdtckijz64vPiOd6Mopi
HrPG67xZrhXCPCyMelJ/i2IpE1J24nCBl25zMq8MlGr6wA2CEIyXYSEE4KIvWwc5
hr2RKWZVRd3aULrYUhrWUq1l5Zve54ZtCuA+xXkJnDKcrh2mSYTqytdgHVkL+gDn
2AVVv7YREbeRyMrSD6q2PBOmYqVdD9gkgxxThnfQjQfrRB6d4/G7jPDNmdoe1fSw
otRSq1JcLu0hJoaHqTvGhLO/4T7g4AkZcvK02mhSjSGBSWESi54o80xsObBb8qtk
qQgSwbthvyOzb3PBjHQlkKU4rr0bn5aRxln6ZLiTuEoCb63NqmedR3ZAKwhobtVH
P0JvP0dEEK5/+/IXEI3u5N0JWzKoYRl7ZHvMh7ekPQiWrNMdmQexprX5TGRP5XvD
grJzuOSHaNPZZ9zoMFr5FLlsbQ5M2Pmq7Ik2ULMAAa4s0ZBPHqhYqHvIt87dukwR
4SuYatzaC7p1GA/ke+7rldDyhXDiAXSM90oZgqSSog28rr1ItchcS3wgyg97iEIW
JmsDDrvFLr+rg7eGbqP6/UM2amjoD2BCHOmpmCRobfzxOkiN6y5RH2Aeshtq3nQg
2IIg4n6tCRxC24a1HlGHm7aSmiw4QNN7cRSv6CKvfGy+S0aKwmBQIXI4aGZMfMxd
m6V3b8bECyZX2z05itiKPJus9FETAy9DqQWAJ6OGE8LVDJS8aXS7kZewC0xVQAM4
JlVcbGqbt+CD/P7a9eL/d9t43ZkpiNNS4IVSYIPODA+8SC4xGSZlC02dz2nKHVLt
rWY2ZcKdxWhv/RxylVq2idZ8eWfrRqpnHOa3T58CfxGQrR5OD541EA0hVpI8MxWi
23qBndJVUwrf63QUrSwv9mFCkxS1VeutEstpibnep0KIxXHNEaSVMkjDDJDOQVjE
dYQ8T4nBYjkVWj99KGebf7fNJi4Tv57o0tQY9Z1xF1FYIJoarXy1ZJZ5vI0YVsOr
jPcpti+H9TOjB5wryqh/89KHtmA3Jj0ETkkdb6ANa5VnhICj6CEmIoDwmRwf5enz
IKhjtyDf35hLJj+mRq9zkUYTE8yzM5ygX0iVOddN9Yw7zJHAOl9e7+CB12v5/zQe
gdKq4JzUZXmA+jGWWh7kMD3/c7m2/A3eaRlyZuRXWgZTS2JlL0+Iu2pKOhstryAu
/HFveo/lY0xj5mA6NuplBJ8dEt4LcFYT3rlzMo+Z6ErLJdByAOhcZRr1EcF/zAON
DEWkZaC178cNaRmqM+JaeFLdx4UeQitXVDo5LG8kgQHzsnzDGL2C9FBO0myBK4Fi
peHLaEjeRQOszd/lR8q/Fz4ree+hXE2k51ryXYXbxtfuzsbCANaPW6mnQeWXvjAC
H+vXspAELIpu0oy5o4OlDDvbe9xB/1CyKfTZndTDS8NWtihI0BF5Vc3kWy8YtRaY
xYlOQ8uiZAkLza8VEm49XOaJF5tv6hA1378qH5PJgFf5pt9cRXbd1tXjYdDefWTO
jiba3au1SAwbkKFpGXtdTSZJeCj2MTIY6CZssJvV+bqEYtiqRIMEzB8CZuK08WUC
9nwFvlBS5y7NrIkleXUlvcQ0V2ee4Z3N1Tq51eRL8g5iI3hXZfmc6JJ2/yAWOlJo
H4ixNYND0a8jYzj/2BWtjD5Wf2/XcmWKlFVX7pxPwHjlETMIvBb7mCvzhR1/nMCz
MfXGpntQVZTrmFkooT6ItwNk8rhn01BdaFDYOcjNxCayHB+GBk+PK72rxD3xR2dx
ZbqMiSBhUo48/QK/MWNMZYOwPDsHVVbjPWHNa11d8A2upEoNNwzuyMiVzl9t/Fyg
fF6vfcJwQK+xrMXWiunKEyHe8iEeJLV8LFJ658CY5WmHbGZeYit2udg7dH85PpOY
FR6F4dKa3awrwQZQJdExdKuWFMfmEdEX8BIXFk5D6ANxY/1XetffwoQ5ssy/8EIT
3WOkKTBP8fN1HmD52nlQEEkMBCFID4sQm5+PHfU7uxoqy3+Kf9/KpIEUWognvGIg
JxAvjIQtLpoN70bRgJE7v2wSw+u7npD6bpex4SWAnuko2jg292sWbnScpwaR4v8Q
AH0eQtTjpyR+quj9galifyncQT8lpxbftwi95ACQSYWxinRHlgkLR8Z9GSGQwAhW
bJpfmNevAX1mBkoJTYPHnooUGrXUcrsbGM0anrpLOjL/X4ZgmadrQVlwdymqnSE4
fvjyEqNHDU6JPyF0F4IN9/quBFhct0HvMvH8XM5i0dx3JUBY7BFCInzBG6XCZzla
BJygwzvPYoLsur4KohVy/Ly+SlzqI4OZSikeQg8flsutpYSdqIr3XtIFJHSNhANg
RC3FjgtXEaV87rhYnG4rtXX7LJgrJnFZGNd2BfVON+vaK5ueaGUWlxWaGrtiN5BN
xbJTTuMVLVIOIkqdDOGMN5NDdZIP9NzvvTMh1jN53feO9QolbYEJ30EavRefRTEu
u53gHCYm/rhs1GcHE2JKQRbY2PL+OhpP/UB6r9esTru5QdD7/PAFO6HOJS7UOaAE
StvIkxwBzYV4p0Lrjwt0w/Wgj323q0IqiE6LNLBlq7eUROvugb61Lw+Mi5Tnu+g1
zn1CNdQLigXi/hgIIT9LGbcz07DFKZN95Zqouo7OXQiGFXo3HzNwI2zaiUyHd87O
vdIYG4ApDcZ785nwk6UI+gsq3qqnzRBH8lZuWc5i6yjvbsGP5g1qgkK006Zsft0A
y4fpvg/sgTOIRBlrtnViIVdUDQtSoijoK93q0Q4vQuKTcmpppESsfoNVXi2gBqKR
3GW8RlqpfGxRpJ+2Ryp/iZ/kP7dx9G0/gNLthrcPaGc65YW+2v9CF+x+eci6nVPx
bUkGzECP5nNDgsiWPeTMwgPVdZt3gxrMgXdVxoxYHQY=
`protect END_PROTECTED
