`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pX35utsf92gqMRwOWkm5txaxoRrXwyMEIiE4WBkyKG+OaNl9QWU2+RGnaWuKk/zw
IjqJUTtMNKxfdLVjlL/caflvgZWzBoRKS6VRuxFN5CtjD0Co5D/P98OC/HAPmkJu
BlkbXxBh+kRTBrKwO+Oo0V8YqSskpkrWR3Wombh4Ds1tO7JhHMn8rnl3bWzLWHde
hLHZx7fOW8CNPlVVNeC28sCKYJjOLSQ9qICi3zL1d2BIe79nDO7VRo5cqeHQkuvr
7fjY+/cDzjiNU9U4vdFid46jbdGk1XcPUfGHXyFNNQOelYctQv/5u8Tn1D+2IuNC
U+A9VyiEbYLaUZiiR+EkxW2UXuk+z3VdTorZc48D0WlSVypOWh0gFCw/G5jsOaxH
QM97cYwqaMW1bJuVmUmHbQ==
`protect END_PROTECTED
