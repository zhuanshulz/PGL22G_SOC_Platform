`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NkBsGrH3+KQWlIpMWmcAnqkLM9PJKHkl9gXQUpSUfp8rKhmpy+/S7BMTBVuX8O8W
3pMlOybERjwfxxZACVEjiRdY/tUT5vx/RVN5uE2UiXerkUPbqRHgagFJZWMfm9bq
C+AXv8r2Dw7dFuRX3qHLPQuaGpEtmgut/So/khsnqs6r/WoKWL1wwhH6yPQVe62S
zBAsjGWY9FbtGFzIk9Jkm1HLw0WEyFVv+kcLM8wmlNYNoh7PhYTcp585gkeoe0uZ
Kdidqgdq33RK7PoCpWNo3xKay0YZTnlz6Qwqv+Sv0gIbDUktbyKHqVSVCdV9fyvo
5pGi5ZSKeAB9GBo8sBEFoitfxXeann/9cusJU/utzklgB3obGjcKyxOoIrGFO5tk
T6Nj7osVnCvzv5DShy9rqQ==
`protect END_PROTECTED
