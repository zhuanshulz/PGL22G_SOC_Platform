`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CT9p/hJEdUIHnoY6kqhImGxU0EDZ7z7OUsqL8Q3OGSstFSdpSpLuDsCZKwCYcY3P
Co2aF+C3GAucVTkMLc2osDKe0+QEJPcwZFO8Aq0AmGE9LMVY5IEYUx3I+9VqznnG
WGZ5kqcJAbOQvd/zvaLGx1Yw7bSPbqT91hXeolH9HHEd/97mVP8Fj4/K2qGgzrT0
M1UeK/2oa422m6ikpqacEaBBdDik7+PFoMq16Ku5lNJJccDGgsfheD/420z0zRbk
64AWeCCUt5+k++3MwFGejoOLE8em7kNEKw1cTzgsJko8LVmPXIIn/i165loAaiuo
gFh7sXuqZ4VVLenyUcRVfMsaCRRvY15N/6Ew/fgudn6ovj2tK/P/e1f4nSWtsF3L
ZhdMwfxt8bCZOq0de3f5T3rCZGbwXcHvtvf9vAvcU8PV6dRN0q9iwL6K4T8usal6
W+TNnj3IObTVlwbqPMC+jfJI81mzycboYBebOqBGR4zVsSd/dbX1kEMN5N73BdFe
3B3RuH6sUFMyb/vuA5kxbvHwBJ1cTBgeGQ7/GEkDj8C5Y4SICa2sdUHMS8x4vwMC
aRDbWjh2JMK9eoRYuW5tvk70L6G/OjPndkqzIXu6arNSiRyYCRNR9wUh8tzUPx1E
qPAZPXFfpvJTrhp/F6vFr4loBJL1A5keZKGtyio9F3uiGYUEBd4uAw0xpO023bsc
s1aBOf5WY2M58OO7C6xkzame7bST0/YJW5mRfTU02tOL/E0tn278cjMSm93Gx2l2
VHGqf+Z3taZkXi3qe5dhXCz4D00U0O7gmUPGzkCAVCnsnJgUl0urucDxJMuuYmsF
IFt7bKJQk73syp2v3tk/avixhbwAVXiYKdbojsw2kIsX68voLH37YCOXtUMXKePD
IOPr+dgbsny6rEnh95G33mzpMMH02WtJyumgxgtr7+nxqHu2rzN0rMh4jE1C36Vh
SSeoUzeZyNKD/U+euGBF76VgucOMRrVwHbHWoB9jJDdoK4q3Euhg2LY9fmgSuYUT
KOHJfnJBlEkxtsNkSA00D2SR7nIheA3cB5iQ/9kDCLCRcCb7/bSIWXFA8HN9+ERn
aDLbyG7NtH9qXbbJ21bcsMekgDRTMPgmAJfNI0Q01hmmDJCKXd+50RC3TRbDYCxI
8Azq0TZGJ8SB46hzF60lHozkIJrAwiBiyMKRKOtuMkI=
`protect END_PROTECTED
