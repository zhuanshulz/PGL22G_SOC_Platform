`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7z/fdbqofITmH+OCJQtWt15SinPN1Mm+FovCm7TQd+NqMjyve3rx/Tb7HX2wbx3C
6lBxXUSuktliAzJyZl8nfuDf+KCuSrC4oqraIdobfijgv4wJcoZHlC5iV55ASRVQ
Hv9xBiSFKTTdPSnzbDU8BR7v7qzV4ZeO73OSnGudjDGSgebkl3jGKTWr6y37K4L9
HhH8DgbRGswFxoHBCLnzVjbL++Zd6ONfSQJ9MRiL2cmliKZiRHz0Sv3arWGmNDmT
vQ13Ed9FKrILjyoBIfIqb+rn64QAYxC26RFNHe0+PwtkeMw34KdHii9WsQL4/3zJ
8QXabU82PwPyz/3vmFghrZ3Ypm/8jwew86osNlSQ2zTNUByLbscccbP3Pi1ETGIX
HDRVq5b+vRhpeB/V2Gt/n3Hq2aiqYaL/n8weGYZ9JCzKm+kQc4YzPM8hSQ22ThWM
GnHqzt5L/ELj79ErD4LRefloaHeP4/6hqJSM1zOiYl8r7PPTP7ly+bFPuj7Qu4nP
8Q32jNtVFRYdnH8TvD9ymA2Xm9eBBOKnkxjzM1JAFsSVTS6sX35L1svzyAx8K85c
YWdQS5U9vtQk9yQ49g7soDhzEDlr4wUgOxRwDwmj5A4QJFvVmn+z+qyHCm0lDXB7
a5UIiu+TtYZWUr4rtF4ui43ANVqKLQHUlqoIHc+dKHPNmxzJdWbN1WOafNgVb7qm
VnkKJveNwCKEkTYyBji7s0UZbJUbq5q07mEK+p/XojZNldO/Ahyp4Hum2oXL2xEX
2Xbk8qCDjxZfQaqeRL+bVlXfk86Z5loJKZ3TykD+OPLOT196tu5uQw3ycsCRNb0P
AQ2+SK7SAzfUKAErN6wc0m1l4+YBNaNGsAzQeEEi0Y4z9TCQIQeeN4TA9rKJsxSt
xCQhFLsZdPGrxiYOsM8gu+YrrFtkjncfZzB6LAr2wKRERVngHEM2xQIOc0inb/Fv
npOAfFcse95/F/5J6wnWTarnceY4sYyANrgG7eyaz7QRNOOZwHe7ny5KI1ZroH50
tKIv3WDY8X3mJKFsq3EvvWM0Cqu02sq97FmYY3RQMUBxnzKHsFNKWQhKsckFbAoF
s1Y/HUMyEWJd7sEq+Ou5lnA7JdjSNg7tQ46cwMoc5x+M3LCVDQcQDkGPgFFhqIem
aXQJqBCf6PrTJurYDBb+IoH++sErvred6kEvjMHAoWUiQkosQLCutQRgzq5czxiG
eBLyEKVMdE12HpUMGlGXDXCrFX88qMHqT8OSZ8cqmZ7kMpwE9jUrsr/ez5hLPLsy
z5c/bbqtoPtpm9sZN+sYGJq5I0aAMcSifnqfkWqZx/Xl7JuaD5Q3WOlv+l+/egMv
JNUGgYnv3OlEKue3MbGRQYvfDLyg8aVtT8W0ZCtpuZfucivD4lf41iHe34Hqk3Do
RCuZp//IRiNGoV7ZFdZBp0yrSiqngI21iEOQe/Oq10oxA+LC9W88slZqQmK3skeI
1JbT1WYxBejRQoreaZeFcBEeSSUeT2sjIkclDot7UhFt053FJpd7ZtT/ilyGkvc4
1TN19aN1jQ8PE9biT8zNl2bnlafmhM9gjfPOXeRwVgSfYVLfZzMU3C6VxXpyQppn
8M4pdVmpEbbZuzrUdf/OlMTX9QPJSn/0A2ZfHSGxJ8/axvsCpcxq/gm4MThQxPEX
PdC1VZvxax/om+CD0HrnU+oVYsNeEH5lpCFur4Lfg5TWwqXYzTQVgGEf5HbhERLd
J+JuSv89y8YaheDpY87BTI4iL+kfotCM5hO9eN5O6cBaFj/mgcdc/lLZy+7pNKkF
ohLZ4j9y59gWWOebTJiLbsKsIFI/RIxiYlKNvysr3kTt69IW+mYteoNWPXWC8joc
cnzSUz2aCynf0L2re63XPtk4cdfIpocF5xJjIVQ3OYMiU6eHp/6gF2UAvm4M/4DE
qAqHosmBFkKH9u7QJZtS9xMIudI+di45UWSpOu022gMsdZX224F04OeQmIdy4L7W
pNxZPFCIcZct6ilMAfqCDmFNhXyQIXPQDTvRSuPMpVIylxzJm88o+WRFsjjLrbno
qvFuibxlJrCXJIElEhJ1cNr5WcdEqbqK1hC/mHbLW+zxrrOjnoOAPJ/7fNQXyvkv
dIehMulLYkrJLjamrLqkGzqyEYIex82HhsBftFtu34Dfzv83L8McLFN5uAGAHsmY
TkjCchgo8acGc5MXZA4hCBzEo0dqQ0fhx5OYqYPBrb9kBhd4EVzUQbqe3eudlFwY
CrUce5CGjbOe5MqW1GD6MbJuLe2eYSwiCvsjayRvkmwmWEAfwfe1bZ2tYXCVaKHN
SmqbmZjn0rOg0nB1Zy/hF389WWSsO1bDBzr92CU2XCwc74hSFlyrH5nipiXpSvOC
ZOa3/MUwD8wdUT/IbacEtm2luHF80HEZekHWXXZXCXIVblV3JaTw5AYG7nB5jBZ6
ZsRUfj8VIIXSrWh4YS3X+Zdied7fynmHUY2WX6imd6r9iEeCiwpYltWBqz+0ruDX
0jGBhnasJbMkv+eozNXT7LPEzWoF0dlx4SXJCH/cDPKPMQNK6cA7sxhCsDcwi4I/
MUR8nkBJw/uIn0AYoYL2ea9VTCQ5DrGb2Q/RuRDPecnh1bGBTGvwENISgET7gRAM
6I0l9Rc579qAtfr2tN/RJMoMNUo93AuNjSlMw4iNbs7dwzk2/p8RdcbhKB/PPBIL
xPBiJoimNqPfogK8LP5qMpxx9KpPUdIJDcUEzrDnkwl5EbVx+EvuXrFfWyRo/tPd
KyPDuDOF2IqH4V/YgpEsjKdAlZv1qarkEtP2pMF/QR4jkWEyudqG3mfS3tRrmsf1
XeeRa59a1xTty9HyyMcS7NPTjvzMwE7pd2EvfRfEwAIg+GvzAlktKzAgem4YVxIR
s5FhIcUJH2fwD1/SqXgD81A88mUm68/lg/84DqCxkEuSRbgow8lV+Dt4WGHeuv/F
ulrWKPQ6g+QkL0RxbWhZQnq4wHm6lYpxW+i8D44yoeU4/WE5Wvo65ESMz2wlMFBZ
ljTZOtJVtfRxdE/1ydbSZm60fn+818ANnIs03FxhsIEmO5BCzo8t7zHPt1rmQQhv
z8XXuHLmDIoGIQGTF+RJkAste+aNCKNs3XIBzZ47xGKrl37nbhKJtHR8o1gqQUUT
71+zyvPkhxQz0KjPt3l+f/TupsPjKLJ9TK9UbiO7jgLFDBSLtTJODH1v16FEFe44
C9MxAOPSUxhstPOaLTwUm0inR28Fm+qm/b+imgsTuDKfmQsda/og2va9Fn8gg9Yk
9CjHbMQ9RSbpH0vp2kT76/HPWESBFaPj+0aR7/+tqI/W1V36hTeADjZVDf7URNpc
anKb4TV6CF20lAYuxqjQjxxHS/B0k4otEsTisfS9cmh+8543wwEHnbW1335vNyU5
Oe3AkYVnoiRoME165qmZeS3N9Oz7Eqo1WjmNGLz/pKXFcg3RkC78GcxqxxYAiE47
hYdYZyhGnkI+VMqueBmmW+uog8B6uaq6Dh3KssLwG/MS7fAAMYm3dGkrTcJ5Pejs
Vjb2LdpFxjYNsqViW+hCYP6fXoV9ekweVJ+tTo1POn9BQiOooAsVaLC1Ds/qa7oU
Fk0Pcav0X6fFY8mOrnLe56mwcfw0MNYecLYJly7FKowZcdL1lw98SZiRLZEYPq24
Buru7H+p42HdqA73SHZynv6VqDT3QESafcDmvld6yg3dH6RwzqyzeO8IOEh/QY8u
QifEYyofH5pNAubmG+k3TRRBahmWpo/Gi+i0me0rzrllYajp/JUXLmvT0LXL+xlu
mlIVAmEfBgHQkNshmneEDaGwTp3Wy4w2dugeNvmw7Dwq87uHL4ekXNsZoOK/7ea0
AvjJFeQvakZsQumnB+mstVVcFrceM3yvVrRVnMOzVGSS+DsH9E00SJ3qejsp1Quq
7mOipq4BHfAORneXYWPtmdr+MCgpINw/t8nGpBW6WrxIXXtHZXnjbpVjTxrXmjf2
82rD84Ozhoo24hcz+7mGlxS/MG/X5Pn9WxM3eUjzrnmvr0vOXMdB5BNZvmIUIgkZ
28bqeTkpRIbmmeJAgz46e/WL+zj5Aj+5ygE6JEs/KloF06hy6uPNZvsrJJKA7mbr
/67IslK97Rwe9pHQsEXrEkOA/C1pX2QiX5+TJzqkfpiiJGR5hn6JZm34qcsFSiEs
nafwiv1Iy2iD6j0bFi6ZZ6nkMiw5wQYkFlhC90lRgQ2kFdWtCqDZztCx/DeCyAN0
T5VQw91SwGrDj70jHP40ZnCDE9CT7h7dbulxH3LAHrVbHU0ndRXZzMf1FgwmhjnY
S9HWYyERm5l5BvnE/mY2RfS/XBnOFiuisLbFku+du04Kal8XR4pGK8v/ucWFj9tU
Ibpproh/t08+efCb9O2X8xnJnLZLxDgukvnjkiiVjOT8BXu4jwYx3a7tNIazrJp1
tnhNtHVY2x93bqO2/KcJ3xND7rOL6vOCIki00lMzNa+P90sykzqdRhC1T0OvlqQ4
6xG5Djl087FImHx/9+p0XQPctoTfFwSFRHvRT391sSjl7P68Zmatl2SWFuUsu4Z8
Kj4VzpV59uoM8UHQS7QCB3cnOh3upkZkDfP5MKz8CFByUbH9Yb0NDzA4+fDGXOmz
X4JyX2bjBy5UppXz3MigMk9pzoaxeXlK2bGSDnD6pJaWspX+6EwnVCnqUoByvMJk
mQH0C1Ut02lKeVxsv7x9wM6RGmiZRxOZ/dC6FN1xqDLR8Ej/KfKvg6GwzvqRiRW1
MVU8n4e2+o7RW7NvOTgp57G/BJGImI0B8uYVN3m+iBiwtR6YHl1PeuKyeVfhxdsl
mtY6iDjamGOHKnkHyruAq7I63S/NlP6OZXNYNMoWKf52OnFt/E7cHHmsHccYVBmI
+ZsP64jNLolTBDZkRup33v7SeqnHNJqMJhRo760XXthpNHn0vr1Hr1BhO2IdicsY
k6QEynlTSFu71LjXSHpVmBq83XsXltDcEL8I9CbqgDzFqEzF3RzQgPIkp0Acavqv
wrjIdoZankQddLtggQc4FAEuRzkMJNvqJluxH/3qj3LyaQqu9UqvHUiorKf2YCdQ
fKhLQigcvlJenNDg7G4xlvg0sb87sQg2GxEgspsfPJEARvcYErcMS5uJboWsUCrs
FwNax1BwFYwBHd00F6y5IcpRGgEG3ST3SfC3gqw5BABhMISfMvH47RE0DhcUIjOg
fdPIALhoJlhWAsK+RFe68jnmWDD6dtX+m7ayUgo5RiTgph5MTYlwfOV6usL0uCe8
rnGnk5O0Rq//RnfDT+VzuJK1F/Zhsl95j9VSPJX5hvdwfjYzzpKI0OHJ2UEo1yJj
AmZLZmT65qNzPYhOg3Yfjdu8t4A27Vzksc/LitOCtfjgFdTaPIHmmQOEAmd88sDm
Jp1pcCZz/FjTkWo+PMza/nfdGBLCEH74pcFI6HVxNspXZ82o270PMztYu6KqTdzO
n2MAATcmLQgzZqujAzBTj4fmqM74prKmYyBVfV2UD4+7v0EaDL+JvDtcsd6dreTg
eEB46mcP15I1Hvky5vwPCVMKxdd5oOz3f+/XoeMnxu3PV6q4CMeVcJ8YMan/gWr1
cNXHc6ztFpDfMrcsB+GS4jTSDB/xX83HoUFEduV8N2/8Du2VEUcO8U6/McSGpfAD
QefZSE1CWoqEn1flECSolfMd1RyV4gGZM25xh64Mkp/gTsZGMHYSARPxUuiCUL6D
+r87E4uAwUK3U6WXvYHtidCD17qX29ztu+LJv3o33hV+twhRmntbHa4oAvsOk6Jp
/ln73LhLLJpKSK5R2SDiXaitE6OWsH4Q9rRkJJcXXOLiDmFHdpsynA1ioMmqV6Kl
78QwfJGOK4nIPc1xAVCksf/ubIuMG5zJEc97FZD1E4vvrs4fui5DLkMeP9rLjZWU
qVC9zw6XjpI0jAwJpzx8ZnWwcui+jobNGLmDXj3lusR21ElIXxjSYfTCYeS2eAOF
b6AWD9WZW65Qi7bcBzfj4nbk0xVfAzvP4k7esQWKvZhAiV7FClwomIZ0SwKk3Bu4
9yBhvSuMJHsuuoSB9iwzUCt1VLCNQtdE+pM8Vr4y/JbjcnvTet7WJWEqCbfi5TKu
fRE4fwgScsXYWKiRriDhB4D03n3/iMY1Dtnfmc+BC2pJ7ZbnnlFGvVX4eXfEx4Ik
CptfUIqRavWbdN3mvOjR5SJ2jeaXkXvYG9m+plgjExHgvSTV3YqerGDSuH1ASrPy
s+JBqv2G6nhdrXTfnUaWYQDqJPIJTLHbN65Akyd5jUVQjfWD4qO2zrqSKTfkHA0i
3bQImjx5RayXKhsaCI7KN7gGb0PLxSE9SZ9/CRB+afwfVIxoafYy/QOUBOKFtuye
ldS+pyefiWxyczfTNzO3FAwGbcZ2tSa+ZkoShiKPXgQdSo1gFy4SpUVs6lVbJEva
ONvJJY+HPyoMPmkEe0Rm1Nk9/HpycP6bEgKZik8P8WJfFVdvZCA1hRdBKfQuwknu
9lkHbC7rtwJr+2gQK6o21ZO++AYRnTlWyT0yg6+/2ReeA/8gwZWVqFJSEZcs5cz7
CME3jqee6CA4t8NexEecatKIROjdHAsyBVCtPmDium+i7vyW+/PWIS1S0TPIxBuT
za0NacEfgwmuqMQeQAeBcnC01ETxz3Z3HzYoN314gFuUIzyMNLJTvtLguK9FQVe9
SOf84BZMWOF1/s/xm7jAnYUlaCpWVAldlEMp59Zx0jra3Qc3pJ/Cxc+NT8Q+73sX
4ryLm3GZ2B/Zm5mk3PBM3nEj0iR9Zw/2Qjnid8TNKUW7PhKck6qZVTHDdvFwMSrJ
+ZQ2XvwhGMAKvmV1SyvgeH/UbjeUOEE9d8cKGvmeUOLBGNzsDGbC6qpkcmUSaOEn
7JPfTgYNRTBUX6OBQCyNZv+vbG8Ni3XXOLw4p4JKMYuXALbLwBNPpc/NNOZc99Hd
4oQQFHS0aU174pJxibyNRUXvvvLGZsommivQ+XI5oNlfn+loy41keoOlQnPMWicS
Mld5hrWee3pR25VpCnB6BIE18MtxXh+xvALy6CKmuZ1pOHVBmF6dHFHRozTOANBW
HESq65cjJZxX9Jr4qaR2lg94jGIHVaX8BLekQ2MW6ec4NhJ/MFo8w4Y7FM7GYKrg
PAP2vJBsFTq5op/oLTw3uwVBC0qbz2yYIT2ZWheN9/rzfLfYk5Z5RNth+6tY6aO2
WC2bMfq8/S5+92Ph5jLh4bmuTY93dW0fCSsTMFno6DsxjpMqLjbLIJkq2iBQ67D/
1lz11ajKEPw4x2sRxw1/xjrBEgTebsJ/sqlpYbhfGC52jusa0BgTKUplSN48nB/T
XbF80eSZ2fmjJ4kBtLE1G6NicQ/7SAWwD9+Vw7kfdvT7eWard5duJpRXcIXYjaeL
ZXQq96JM6NTyhDIRCQ+l03gjRj5cdKRnGke7EyLnJw3OblcQs9xTzXLoWRDrigEa
dSxhe+7769G6EFfB0jE+ZMUt9FqRZXHRMgt3jbXJaWVGVp5NXbzIM+nbs+bmsbTw
9enE1yQXSzoW38xo5meEdYSAyNBM2LR8/0VpCgk6BLAqt48p0FBXr5j3mL2WnIaG
1+LcljPW4NdGDEk1IQjOWzQqrL4yKPnBy7s1j3ssxsR0sAIGh2wV6gKTeNsOHr+v
pLCjX4ObVReN3bJfwc7GnwQicFh9qo+MuAXUo90zaeIC7u8ie791phKIBX63PBrI
nL5u9LV3XUxA9iO0y+c+Ohl4th/jZNdYyef/+UHWN7rdjCgAcubNgRyp0CRnc/w3
bX69jYvv7H/q1pvNJOySQICptROp+b+rBvGKGXm6eAPaguO6bZNy435cz22znFVM
607gY9pslTzEun3/bnNLJdrLbqGXAID8J4BQ83g/TwWQBmM0BFx2EJ6y6cDtZAHg
VEO88P0x5J9QkbkK9Nhn51p3W7GnWcNJxjnj+EohjJrPuly1dDFFPh37qSNbbbRa
DBTwg0//GB0/OZEUQq3UfRmp8P6dkJCCnOGNNfsJa32enloUx9IQN+yckeVj4KAB
2ThzKrfeTnLiXn5emWgHTh4c+7SVYAIO0rkVgLqx6XER3Qs09ueyx/DHCG9LYzoc
nxfPqSoUiVMznyHov1f3RZOIPcjs0ltUxUfOS8KJyPwNUDbxuhES6jlc3Tk0D5iX
tkoFf2RaiHJsxuVb0Ga53PfZsT5Fr3GY4+y5MDl16U4oDRQDru0ZY4ySP4J/FkRM
XmGIBJcuCNjz+gjmZU5+8SpF8VKoS3dkIhKngKqZLhuDcKt2LwMD98h8nZjAIAJY
MATqXYec3j6Oi2awpNEWRHd3PSxuD/N/k2s+le+h5u7K6jZ+Jn0FrfKvmE/5hJA0
F2MIvy1wqeb+6bwSpszJyzOxaMnOHlLOjHR9hECy3GismnUSybeQ2HxZVqX2qtAD
mDRDSMr39/JJciEdeEPeVr7quPV0hEOypp+QYhN7dUN4IFLPVmdoTSyUZHrYn6lN
JQgOtn+afEly5bJUnvyFb/a1OhgSsfIFt29EQbpNXh19mJSM9VKz1JEGg/n409kX
0MUgvmHksNo/AtBehyHIJywmW2l2OEbbazaMOh5/eMKVPHzfClcKaakCmye9ytOH
eR9zdMbhE2I7Zc1GdHwYHVliIue7xZ7uA/vMwNwZ5Z/K/EbjqEUXsNdLDVFHQLqM
5vf1TLrntQEJP8pu33powDL0PYsmDyLnTIXg0X/uU18BWgM9axdA3WYOT3mk3QwL
U6r214M8wbyyLKrpj96GDWuQVchNal8SVYqt8oogwFk9vLvU3S/qWnJKF2WXFGGl
gq/NHloYMYfL1uGlxJevv8slGcTEKdmzS4wGjHe0PlsuMgTZ+egXF0E8trMHBNws
dOBvSPKWQxudR4HqcxSOxs6Wgn6A6TIs9hYQNm1ya1+kHXGTTGJmpNNYoGjsm18U
44GAurzdSgbh47Z/sHXAv3L8wAgZDLk43siVDwAm2Dbp6dHjYqH6+3Q2pb5ZRr4e
3lWL7hmt8rRFkZtUQvRH+QpK4oBBTA3k1nQWY/6fiJ0JqiXTgpGAyceCnhSaIgik
oPJCJClh3i3FZwvEQ4Rc8WqPGLIjv4zgGrSrRwNEhbSEJOaPpjRGoqUGkgJVNw5x
H8qE2HgPvAXV/klYejEbPgEDbU2ExIBc1tiC4t/3nry9ijx3yUjhYuNR/bx9bkIf
8JUOADF9MXRdGnqaN40HaL2BOIlEx3NoQ+sMaUF3c8DOp942cyX5nX/DtZ5Is+sh
UojXstK7YmELPXVZWZclXd66TZ0bf09FIV7RHhnxM+v0T+urcDJZMwCZ0S0xCSLu
lINrIy3dK6Zke9be1+7x/evD9436h/9VI/pEnMgDt2983MB8BAWn6w0VmvyJx/tJ
CoGtzcn90Nmw3exhIK9ynRSSFYWmsvtX1xbi9ZQdGxoQFv5fIV/cVvqlnWPz9EeZ
mdnkXBEMzTgAVxWfwGM4jKQwOfFW8IbWCcy1fLKvrx9bJwxJzqf/C0WJ/c5WW9P8
RdAE1veMYLA6/t7ov09urEt0gPQgxgG7ml5OfNvXsLUGjaDGum/4yHIerY++PFO6
9fPvW4mMeVuGVFF4a8FhuzMy6c9x3P8rSRAkiteXgouM4fjGR+X1yqotGbf9H3g6
FMX6klJJaAGZ120TEE1v27HaIy0+8qBynCdBMDM3B7ZPxuslJZ9VKzb5A/xRRIGS
Yryg9dYWK8k5LwCJOJKWRj6l8/Jx2pj8WGfpksv6+AunLjGm3shdtz0X76ICozk/
zNbJR7G3Js4oG2gnj3KNIoSnegub7cNpqDf0EuHlrCz/7MuEyF0JmRn8/F9/hi3k
zfZ0FWYzmcg+SP0pkeuRC6PGbKAJYMA3cwTDO9xg4O/EpzGRa3SZdfEM9b8I16WJ
rr0y/lnLei0D/q0KlTlDsAgFiCagc0/KTAHJ/hfCGn9n25MauDP52p+JATbCXI5A
uFWSzIPXjT0AkJTsUJmtMkLCmuxhxKE8rhtQ+SXIDLiczy0yfcskFPXQcwd6NhrB
jhFoQkV7ZsP2b3bnpp8Payyqd1UJr5txeqX0wl9MjXhFeEboGSp1HmZSR//FXXZy
Do6VPWgMrDWxmM4ttKP51NcQK22SyheYMazN0CEeEwHy13QbFkXD9IcB4mNMlKmC
ACv4Y9LM7SMq5yNGRKMZc/Xskx6RePGNcLjD9cg3N35LwJk5q4WJnQKhF7OXfmYl
EeYcBsqsOI1b8Af2zlwuJouPO7EZeq6SWSgL+NsbvSyFhErNMlOcVoeOtke9gVG0
ZtfSe30JficD1isYjY357DIwtKo/7Bzgh6HBrKB1UIh0vqV9msykG4tDk+2ZVQZM
kp9MSOq9rvN2ymUn7l0DSnN0BOvMnFHgLCB8Prtnm/Xwwe4LRgFvXMswIJqti5ZU
8D5dsehTuB2dbZ4XoiG6dQjczlQdaS+12TgVOlvpnWicLdGx/kR2FCh+k01o04Mf
y4+gfeKTsEENNUQUHAdWxZokmekNqAD3L3Xm0c2gRMlgYg3vYpJHj0m6lgrboZyo
y9oyoovmmHKCOgOiXmnVGDgePIbSDmk4M1deiBnqiQFbqjIVpX7CfRRvawqk8ly1
m8HYK9Df3O5LFe2RGDij3vDnxTdc018po8PN93B1shil1ifjz6TU9EI2v3crC3sr
DhHu/g4lfRrUSJoLfZKBPGfluO244ZFxFGFcOtUiGtuuEKsxhD1qO7zuAQCHfR+Q
nGW1Y9k9d5qxEcOfZr0GgfM2xEJEORMjPYWk/ZK16tWlEBZzz9r4RTPgYrm/Fot0
JHfgX1kXDjqhQDZEwttm8ez0lcn7YWj4c+mE3PldBxvWINk9dBIM7UzNMYyfj1AT
XkfJWrRVXC0OcXoHEYi1sv9phmL5Zrxl3ffWhDwFAYTdlqZ2A/Nq8+BOlZbbrilm
hwRKYnPPzT/IyRHl5ODvrNXqKcHvR9BkZYL30nK4yZAO0uIk/9gEReNGTQqTI44l
dCEEy5bAJDPtzBZMvc7RjoxYin/2YGc28UcevOHaEA0JSTyzRSmeUUrmNUhZA9xv
iiQpX7GKtK4KiwiAs2oGEx7PClBbWcGfWXJMpusXkosSwbXvUfor1UQbJpj7w78F
xVGn4//n0yPhASbwvla7WwCOpvT9kB+QFlxEYTjjhvFdN76NSczaghfIUn6FE4T0
19U+vvZ3TPX18djXTH4YtV2n9y5hsnq6WuBVqPSkVW7vlhtRQVWIhVq6MQRvCLPF
F9eygSNQ6lJFx4GBZy99gIaRhw0fzU2glKkYDsCzKqvQAdEh4jhIsikLItjGzjzG
WFy5OZXzaRq2j77UaVxi0l/ziHxrxQ95DXxIU2IgRvzfQZc/+mwx6NnWZXGxSKne
nEcVVdGs2ZT26xOrSXkLkaKkQIh4y7Nbzxu3usC1gN4uHcZRJyUxiVmey/qwjcC7
XThosEUDhsjm8sHIE4TH1jVuVpN7NIQxlQImqCjIbby2wd20wgThRwrsw23nnPs+
rmLJmodasl/0iQW13w8zW7ZzEzU0iiiQnbuD6c25sZBoJdnBrajeZ/8LiQvXtUu6
NVRbsdWQ0EyfAfxIexggVND6999UrhKnas0F8BOkeY6Oi38NFgyCXL77/OKu0+qJ
6Rw6kK5+Cr6KcmWGwZk7SE2rnZ6NlTmKUE7Fbhh4AcaOj3lIeWpnZg4esAkOUz92
ERSGgyp1dlsxoen5o8dcvZlulceib8h4R8vOY1a1aej4y3EgvOil61DeTF+qn+6g
y1nIq9iJdQx7uOijVvtHfwmC1uESggVUkJtGXM8DDQFyb5YVxPN7vDbYWNIeA6zP
6p8iGuuOo2QNLC4swg70UJiZnQJ8rzkOh2GBHK8JbdOcvl1Ex9XDGa/WxHVt2YHD
iTxNY3r6J1cjPh81CGHduhM9d9PoWJWphSW4t3mS4k+TacZUhdREY2+6xDmz7AjO
2ZNBCkbPHKebVptQaoP40snMIxFWBfiITa2gg+og7vmVaHlafCr0mUGDa0mGYzAr
jzAI35iYnT2mnOmcLmtVgw==
`protect END_PROTECTED
