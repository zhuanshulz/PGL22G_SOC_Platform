`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A48H5bneKWRWlqI31A7klOPZ436jknWFPUARZ0awWUMULkcnUkbr1HhF739+QmBJ
/sdWYoL5DJXQwhgfvTxvCNZ32X9pG4VkB+K9N/ihiIng2beQaNrt9thEaP60aqLe
aNOFdy5iTvrVTuw8lIBbs1Q+Yk3/5gkxaKJDBCnDXLNR98jvqOGgD9H8ckULgmHp
psLKjVfC4hO6CMPHv8BW2Fv4ahqtvZ2iIzBa+WEb1qB9cQ5Jkg0HdjGET0Mu6lJe
HEzK7CAQXBdtj0Ve3Dmpi0uf+c9gaBQbk+MKN+SLaPCt6udFjzdVFes/1Qeq14jg
CO/dd7HELaoSqRGIuTCu6flC9FMfUz0sPA8+ki2P7zX3KhMCjny0w0ORaRob8mcn
AWeeJt+vsOG/9OjF+1fUqa6hEerEtSHxdPz2BcNqLlsZuUhdOEdPLVvbMryUBSdy
U85IMLS4qfDSdnKZPBT4PybK7TCkinSbOXMJzXM4w4AQAqU+A/ZrbgERQy52HkTS
DDlCEMXb1IxI8bSX9xtvHT1PlLc5aSP18nr3ThDgmHVwz7mgahbCHZA2zd5nRJ0g
OQFI75ubNqWmjz9+koZRaaxt6o1Pii12wra6IZRDrIU=
`protect END_PROTECTED
