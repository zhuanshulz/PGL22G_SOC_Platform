`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEU81NTczzSaITSvWjHrWl0J4Fe9jG7NhVjvwJajw4uSBdaLWx5PqS60V2WKQWE2
BxWJo9rPYuhCWzQ3OgCcwvmEBxsFuNdP42Geor9hRKlLr78QABcBIucphbiyUJhG
h2AX3HV0UfET0dUM5j5vMfb/axzSchsyoBKMiGRa2vtBZjtXjNXIfq1feKX0dgU6
dTkrooeQ6WcxEE2Qrm0uwHv9n2s1Vk6SctSejdlO85mNuOjMPIG2eN+WY6hCf9sA
vc0dyHunAi31mODT+ReMB4GKXguAhvnjyP5mUs4U7b3tPILoQRe5Tlx8kNTnXoey
u+HenDK2mAkGvGcB5HVL2fCAr/JTbQ4UdAHncsNY+MH7I1Xyco9d7JOl+r9czwtR
ejA/V3B8gujAaLMEBz0Gn2Rh7mjpW7gzZojIz6F6KJ7hlOFVaYMNF9439lfwiKGS
FrSZwMZSZsAsO8+Cz+x+ycpimxt8m2HJYbpe/kyLcowdG04zmNcy0VyZaXBoz662
r+ww9U9OdTwB9tyBzUBAEKyoVGJl7GfvTi6Kr0MRLN3nGll/I4y/9C3UtSKeC5ON
f9gg7E1n0k3Ixg0O/c6bealJTPbK2FqHGW3nmjm0xJD26+SqmMIXAi7Pe/jL7cNT
tXpLcKY752FH7TmBZdrnAGa0+h+lXEdv/M7WVW9osikVGhmPb0tF+RRQl/Sou70k
sLvV61eJrX5TnH0aYbfIzBffvu2EPEHKagtu2P/OPATZxCu57bj8Zp3laYcfyvPS
cX7h7vMnOdTGaCHIq+G1S3pOWLsjRATrwT7gK3/FjgKguengnIFObw8chxmM083/
B5dwC5xjn1xq5h/jOyl4WPRVaQCeHyZ50a/cN4+xK+uB3KG5g8AgKY28uckitFKc
/U7jHOaY6zzX6f5Z91/zTuUzj1k1+Li6I4dhat3hEPTdLQ/Nm5PIHJGlmC7svPQd
bJ+C+Lyda7xg3De3TD6ZV9RJlHCHI4TrUXM7rpN5uLKBJnx9xZHjv+K/crofZhXZ
7sCQ58xUlQ4WQwBziSaySkOOdVfb8O3LSj+dkqQ9njri/OrRkILYwxgHxxvXBImh
TQRt66+B3ytvZtYb89ggXimfMoALLBsrbso9HEiOPbrtSNxUpMF0KU2o6GK8QJDT
WYg8r3E4qaJxSfrDpoza2jl1zVNtlQz3zFMEB52iJ6Ltx5VlulkwxGEn4o3hr5jd
UwCc32o0VTf6yTfoG1xZqSHzZ39LXfklPYqj5BF0qRQZYmmAraEF4XpOJVVO9Lpf
DCoeVGnnoZT3wz4eQl8v/rpwEtQ7EyYYFsODGbcXRuARCAOSuLQcXlGELESaRKTF
zlDjFZRmGoLTSDWsSAAWSNgmVUtZtMqnjHi8tBuzfsCVm8S8d00gxbacoHl/pamU
keg/5elc9OfJP2YVEzjJORIxjn18ws79v4mlxHIqUdu96+kFfgUPrFmWCcd8J9Ta
YhnJIx2dbHrjDruvV7EXKsZusWT/rcUocQjAZBpVGZExUDzOQWVli7/tzorMfZRh
ILBwQIGKgSBZHFD5UOhMjqYZq2DbKHD3U3Ckn45jh/RLRYvlQMJQJh6kzp8UryfJ
5b8zf6p2THAJDVg2vtlvt2PW4ylIBOwx1VmK+BWNpKIKh8ItJNg70wJAlg2CTrZa
+RNVaWxcikpOoNkqKZxnXywwPygz4LsZG1N0MO+I78Jx/WURNd9Eb6YTRrRk+v40
ShLyX1Y0giJHcWtVkw3wiSPO15lV+KoULjYDFk72dX1P8/+6n3FuNab6eRXvZmzE
TgJqfasiNMda5ojRDXemN5eCtKuWoIbhPd73QxfEYPhkRwPchf/pViExr15FRqNM
649T1HIGs4n91Wu5CUwVlP9W29sFTg6SPJOk9IzZvOdE7x5TvJvEwyi5xWsYySgq
QSGPJkE2dtnheinggZ/hiHU23GaQKn1cBR9AEI2ZU1Cf44Crou1hCJ/K10JywJhy
7btcE+V3DqQuExPKt7aC6z+T+3dlmO+DK3mEkifTSxkUXGfPIGY2lHYapFchqVmC
hXGsgsuzqypqP/CbPH7tX7IkrHJ3JT1H0I8v34nVME4tqlkfANj2EH1GShfd+Uzz
96+J8t+PuOabuXDO29xznnppxxoAA8bCUDx+nTai5Soqxm372l26SpL7FvwQB7iN
+1k4V9pHupUkXUi2zJkxhNyvEFJr2JsmT7wwl0A7QMfRN8esqWiFFi3tNsPRPlJO
p06yQeLE9PyTFE8IJjydWYVjIMy/B5ih501nSl7pxG6RKvVwyzUL32d8xfkYRtqI
8raad9QM7Lbo+F5Ulw2HQFh8ZJ2StPAqK6ylnGpJSV8E2iDmOame/i6DVGIpUsM0
3ZCQMSvabBRMj3Ltet+yljnuhrdDOpwPKV3TPiCEdY9YCMeCN48svzLCgWnFL3SC
y+9TtpV1Gr+T50wvEydSWAX3RtBDwp/itGFA4gLW81o9jMbh0ciw+WA745QG3+g1
yMz04hWMow5mFrNas9tsbz0Pp/+ZpiHTiezd2Kibmb0spZsvfAsPlYAEQkGHaGPU
FWXPqWogmhLr+se3tQFoPwvXCWp0/fW8br/7WU5LKn9Wh0lTeLpY1AhG+KZ8N8Og
D6/+92dLQ94FqWR9KVeBPQbg8LSByM0eXItRTIRTLXu9z7pQvB94ZDeF5Qk+UtCN
PrFrvw5sGH+we3MRxthtVaWkwcGCPVZ4I1UwfwqIw8uj4gqvBj73ZHJ1NJDIFZQB
3AIjfh20GpGe+sW4oWVWgpK2A7RN8w0Ymx0R++BGEiGI5r3XNSz23XfppR1m3QNa
DBbxm+YBzG6asd3SHVpvI+8vOJJj4FNpUoa3HCEqM478B6a8lHquuCiIUnG+3Pjt
ZhnMKifQveJ2IMd/Awih7Dm8DVzCZiH+g/Ltjc4MoVEBEFCesdHKUB7g0AqTmF9P
DKojxEovrgTjvGf7DEPSGiDatjbdca6ZGA/If2SWG5CYbQ55v6rdsyCWicjUmoOu
PC2ktzG5PvApZWk1rK7YbIVPEllf92RV1WhEy/nmWpat0kws1gXP3SvwouXlIrQY
/qebIMBWMVEnjOfXoqAYrJwe9aCFPAk+Ob8Dz6o8zVIfNwkZWb1DjyYzN6miGCM8
obZks+9I6xSyvseI/LMk49nGliSNRbXQUgaV7FKmk47rhO1l2uGQOBQgxTE9FqL9
c/Ds5zwkyQtizgms1p2ra0t1mrSKC0r3GUdFsxHRGecx9KClSnXKRWXJO0ApjlEv
DmFU7XrG/JWei2yH3wmLREP6hV18G8Nt0t5NQZEEVJD1WGuWheKqytc4fB2dxsQn
sVlxELCY2262amnz4U49jxMKVD9ET66smZmF7F6JfSqlaFnkyD67ZHuoX9w+rTVO
srQpA/cr5wwMIWZVoh8rCBpZFJ/4bOxI4HXJ+UAC1IL2nL0Ty7Cabe/ViZ9rIxVL
YE7vbpzuYTl6zPW0GlJvUizQeR9dlpRBaJJ/GQJB+wwPaqMgZU3CMoaPSkA+GuYK
iVSRsS8ia7svh72HcQeBqxGcxXxU+Pmxkt5LSp925bf7StcAFAzwaO+2cogNxSjR
VGBBJ2sm+yWzTRQq8b0a6cBeo1wOR0QodtZ0xvBIwL+kx+ZYbEmiuHDR+ZvoV6dN
btwnOqdGU34Qkp9f5gHRHJkPzhJXbusB7ld0FVZvep+Tqo/eJLVw1DAjS6tSlGLh
gfdAJ9OJnoItQOcyYeYZfTLRCV5CoGlkQeQsW5RCKO2+4foXO0RuYCe6DP3UCZXQ
jv7Guc1Rc/+u88NLPiiyW32TgrLYQ5yA9wWFNO45/NC8E8OKqKp4b0vCiHTwl5+L
0idqYI9qarN+WcBDQ7M/FaN8BDIjS9D7liUIbafEZBayg55pAwCKCg4Y3ijYGeyw
qbmWI896sevmJjMUWHBAj2jkCwLTflJnqiVMgw1Di6Vj6+mKHk029jv7DGt5T/x+
057d+pVnwtMMTn+r+/zA9RzwqViUj9c5dVzTYXYNTmPhOXdMPLjsDBJIyevUUx+J
pvfl2fg74IVeBj48AC02zZ5OGR8MeN8v/EcVjrh2dGYmkMSToyg7//YpKly81EPz
2CpJCV1BWA1nv1Isp4l4NOq4YlDFTGDBrY2mJQXqIhPhpoFKuCIwCm9tT/k/ns8p
mUOqgWH5iax/6P0cvNrpLKkf+UWJqWFrQmMWYpZgmknhMe/HsZ5JcbnNEbejBTQ0
3mDCbnLT78uWznS4LMQHmUWmlY3scoNtMk1wiZEFSmtUaksQ2mlZd+aulUk7WcqY
P4GNk5gwEyd2vZN0ArZNXlH46Y1nczT5ghI92gXRPvyfin2e90aS4jXTCxhwwwlX
tAR7sxsGkQVEwhL46L9MO/3s9O1lfHgy5LlssIQJLIXw3hksF/2cx6AkaGhEUMts
axrLMRX5QettrQjD3AOSOwuhU/qEjtoR1+EdBIqk40PxKhcKYfF2N3C3xWcrs/44
mZEDMjvd8gj+xx0s9m/7rO5I0kD8sM4HecyLB1yg1f9e/ebOzkou+wj1pdGzsuto
gC345ygi/O/sHKy7/xr+FpvSH6VldFFFODQsdjk7YT6kUzRwzqNwZv7VBz4WswSH
6ARbW+5Pj8PxGcrP8avCDroQhiA/8Dc2HM13IKIz4YFoDak4jLRdns+i2EZwvYxK
gzWKbLH+QvtlskwvAfXzBD7o/zIbNJUIUjL5G5Uq9y+MesYKW/kfSBceyyPtq5va
xekoN3OZZpQlbBc6/C1PQQE0RkEeZGWEZTdFpmyJl760lAbUOmOmc7X85GpT6Y6p
mwMZCl8VmnYtfyes+M+IPuxfnR4JjARZtgVr3SwP+a/OOO70xPU6MmoruHtXZAkO
I5u0fD4b0JKV/yLME5VyzG/r4yAKfAyJ+0HA7Jbk3isRgLeMaXZKOPDpZwNGHq8i
wq4i7muxwEot0bXfaLdS86qeSOI2GNxuEUpojx35dg9qaeVWlbf0TQ6D6rIEcX0a
5doAGt3kA/b92/4MA9HChIwxUPBz6acWAtvvCJtbMwPcuQYTmaIJ8oVA/S8j69fy
PG9epKfqeaXC2rRf47aBUw+A0FFu8BLn0Ig1PL6HVjaITCRH4Y3Bwah2UAeC/ZTx
F6E8cMbpu3X1o9gPIXNCeKYxX2usCxGhHksVQ33Ch1l5ABizOPlghUnonTDz/rDL
hlNm7L72QICjGX2fGuVdd/aicNIVTBDmrd9NGiuph/IIX9OZMW/6806VQfVwgcls
/joz9TT2m55tCWrHNgXzpAhzgCjLDty4XBa88KNHphad9g6UZaT/B2EUqQ9kvcGN
fMIrxADVXeRN75/WCRS0dqe89Zn8OfUnvbW8TTE/yFv9JPrAyC9X40+leVQafewg
hYJSdYYlEDkKwITOllu61MKdsxDyKl18F4/BfSTMKtbWpBaI97m/9XBAGxbyOEYH
vPYgRUlSBvdgkrNE8amSWfkY6w9/UP6v0DigUCYV3OTSkMx99sgXdOjJeQbu4MVX
r6m8Ok/aL5t/2BaXn2mpLPD2zo4RMd+zBwN2G/Ev281g4hcIC1AHvp7vl8D1gTAy
o1kckzSqoLGXynC1FOAyurZ5Dt3IFt+VCH3r3dIjSXKjf90lbOjypKMpChNiP7EE
LSwLsyL3g5h5tro4g77JDqVxQebLPE19wiSZ+NtSZZG4T6gqGNRe1dEnh8dNpOP4
hSrSjnFeIGjviS2I5uWK8i3jPPHKB1R5DRcY5dFHCYnChJ1Up2WDsHwrTshVBJYc
HUpa7Wqlm8hUVqGa5DqM1d6gNWI+dyit1TZmHQsSqjbQznXA5Ds0kvkk4yz3aFva
XcfkrRouAzB1+ajg/npmbYGQ4ch2Q/QEe5bmIVaQS8xWFbJom3AJrdDsSiJshHml
vvjruX4uOYDYTo7QMKWUjtfyMUx1wxNeipkmHXfS5iC7xkjmiHoUJQ3p5np2avob
XCXZtFilw6GWYIQ4FP4Lkv37S5dreAtGbgBsnTNUpJdL/TPlfYRg6U6ubVdKkw5Q
8WekVx+ZBPd9xUF+IpJ8bjlT3SYTZnhVeQ6U2p1M+3PMpUMqFHvikgS41xgLWiBe
SXZV/08LRlCOWraLfUBzWYozT8poI9Zxj9ce08WmhIcgVwx9XyY/sIzSaGLBGJkV
`protect END_PROTECTED
