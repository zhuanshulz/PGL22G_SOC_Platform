`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k9XE4JaWSm/iRvKXcL0LeX6hGvD8cjSDFaCoV4DuCytTUQ/HznSN0cwtdTLH9TR6
lFXVJF5xw30Jbvi5s1F3nNmdP4ElO060lvp9/6Z4Os+Se2tvAI2W6P4y2IM1FoXR
CNM8fVJNyqgqZBJ/zLKHKyf22a/HpDBDHKThMqmpaFxYAe36gJiw8NdZw17YwAI6
0mFFmM5+0JJi/CnGlJj26YER/30+1ehU7+YqC6wMDIcokSQkJeadAILcRtBupaV6
W8H9vpY3GLhuIg7Yp85i5B6Gv4UTPXy+w2Ta4UUNsUAWdqxWK3DmPtcOCHNDm9+8
S035Sel6mO8qlfZGCdR9ZgSDyAa2ACHMo1OoZ48mOcS1dSfj/b+6lfk2Udr8j4m0
qEve40lr0gpHcTYWHArzNFI2ilTPUU4tKhwe9MkamE52L3rygztH4sPodDFb0zf9
P2/pulUJaD01MzHADucaPJZh6OvOfUO3mFNv9JExbA3ZNzyeIz0HAa62RrTxR5Et
XMdz/eJxkv0zjm1FXPwgdMr7oWqkdtsqZRNCH/JNo+jSyRUlgg+0EJ640Ma5Ho54
jSGnPGHsQ6a99hfMwV9Sqs2sWBsZYYukutNTIfieb4RvlwN71ZrTTcyqLBL4D14V
70TcAwhgGQIUeERyGbXdW9WFRychGt7bAKlcHTAJBD3ey0Flz/riuXsLhhMzXNyD
/k96TaRhewEUSkVvJm0uPOS9P9Zb6lkmnA228RyNTa+Q0skKM9kOJBdISAZ1N7+/
PmgRQflAGx4JFESxqYFpToH+u1nBV1SI5evBJfVq6OmFuQcK9ZrovXkU69h8O8n8
02M0krTn8aZdLicIDGQB4O728koGqWkEsy6oNgzW3+Aal38J6zhCnwwFnkKY0k44
LjkDee/5F1OkJ1xbY3GjvYR5B1hqJCDo1kKZTL8KSut8rmi58InQ7Q9t1Fsd6xdW
IsRQ4XK+pQM9u3eg7lOXLeyypvzSojAB8R1KfaYHx2NiU43uAqqfnCeRRrxaT+dK
Vk1whMfIYJVE5Gtocs2snKKPjj9oXvMevyPRlILBgvuxUZ8XEyG2+U7P9nhN7Zwu
TYAHgFoYHWkoxH7zUKLg85zedyjbP2Y41W4Rsob7ujwwhZb6ZTTQWCnyK+4Cfgo0
NOVZTZspZHOitisaxg1clgsz6QilxhF0xFV7oDbHgUw82E49oF2Zm/QHDv0W9YPN
BOKKbyWeI8p/VcsZytx3HnuXKMcIdGeu6sexL3P8itVzhA6QoX6gMLuOHaqgeeYB
ov4N1QqHlCE/zenba+6p2efJvptR0QgrU1XtjswcFNCDnBTrzQFwiiLwpRTQDn6w
v9mVW946GDVQqGCKKpOMfgwNoHwMT91KyyWo8ClqtYE4XzMH6MYglyKSysYWqY3p
RuRwPVHsfWLbxL39X5CI1gvdH4P6eeqQwi4iBn5140gdh2Z7Smyb7MQFSBRfiN+C
9bftcxCfEt0AF8mTazSWCWDWc6tte1UpPdMZINGYcu9OskF8r6AF/rvsZ/wl1q2A
5ygNEBUeZqZpgb2FWo1YKX0X5Vj40d1d+voz520jxgPuUFraOEdXx+Y/de/w05iz
OQN84A+Xh0Cng3O21lvJKW80kobxYLzpDGOAy3N4whN1W8MsqFP22pz1LBjm2XnX
sPsIG6/TIm1PXDHSi15653BfX2/fPCrl9SQJoFDXcXnJ58uZlzO7koaIFw4cWbzV
y3KeBVltF0MKr/FN5wPTPOd/ovuavz3GPt6ZiyOSgBzxpW+iO2aFlIFj6nfD7Yrm
hWh0EupyH/4+kliodwqQUXuUcz+OdvD2GdJAX8YyDQFVyWiRb/I+Ndk0Zjbj5HC7
m7bmwRodNY3OYms00lg1sqi0op+5MZVTyW5Kupsj16SjLdQ95JGWItVT9f7rRNrI
qbx3oePKlFIz1jYziwPreZus552Mh5nm28lMw8l5C7/JrrkV7tZHaI/Xh1uRfg5/
Irqu2JbOYVTwtHWz8oNFp2ghMhCBjNRqTxy45jAkkHBoMfj2zXzP9ytnPc1z+YWS
cTU4/QmnuPCcsmSSgQfd357Wl5bsguGUdxh/9QXaAcExe6wVO77wgK96ly9cPu19
lskiY8Iaxw4XP8FqBuk4CmMFiPYjn4/EHhUOiWe5UxEdaWpZ+PwbZ4slsOIa7WE7
aCzrr8K1/fYwMJzWBmpahC3m53LZJfQs4h7W9SiDl5rnR8Hi4e3jjMhI5NhmhXCO
rid2+WBrFcuLBXYJ7G208NW2fbwj/0bd+sn34xkl9r6NQe9/1U7jqWJ6qAE37xmR
9ZRfyHdU+oGNUBswfyz3fwVsEmWv5O8QEjOQ49NH0DUewt9SAUXOWlx3N0dYXmsE
nUBLzAqQy385f1/N+xh2cpcq4HKjBG8kST94eBP9BRBYtvfae3LCPCNt9sVI8XOx
vfY5WYJE2I/FXj3PdKzsfJ7CeAN94u1Y2rXGpNQrRU7alMBCJgL6oEk+0M6WsnOq
xESs7/J5fJDTuoyFpc7g7OqjJ7z72/v4xPh2z3qZe0o7rcLNp0D1oAtwkEHKQ4DW
mH59IucvDA7Wludx9nKvlpZTi3im9M3UxbHlsQ6N0cG2+iSQRH6r6+rmOiH4eNrp
q9VXxuvcQ40spLKtutxZXq0/olW7nvcwwV4ubtECPlAfhDynonikBcwMRBRwBEjP
ZMzqrAJwd8I0DQ1rTT2iK/DM8JkgwWBDIlybD1rpmZAwofyKCZst1cNWe/RANyx0
3egAMkmNI68ZFDPUE7KeSGl18WAWlMdNJN2QJvxCMi4HYvQqU7X5l8larIusetFm
2hktzVRFe9rE+GwwAsw/Ow==
`protect END_PROTECTED
