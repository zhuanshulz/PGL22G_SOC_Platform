`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mQU0gJLc8jPAYIPVXldNaWLKVuLaPV5IIhzj+utA4pv2YYAMmotIDDHqxV9t1sr4
9UfeaLVWpYCFg1uVcmIyWn/8abiWzsjD2bim8amGuVt7tC3lJghTfQSvrkXNE8Z5
8KYevNXBO+jdhQYtnyZRfOrNob9+7afK/0OITlrdgCXe8XTI23dJa7DLsZCwLIZq
My7zlCMbvUSJo49i6HtBtmxEfvbboCpZnoB7iw8KPf9eX0oqU3xco/qLUN2TIhvq
b58udtw49maGtHWxUGm9pqCosFn+HXI9FM8EDHBRGAPB0YclzTYuuc4/ma6llj9Z
/9taPEp3DqF5kc6S7Mn6e2THsVqDEL/2rQe9D10pVS1Q+2Rt9SYcOpnEiVHi6los
zQ+R1aMfL7QnBUWWc/JE/r6ZaFyrjFi8evAblgcZghSDgz9+t0M8Ne5KofL8wxU6
a4L1shKmMQpmvdQMPD5DWe0TGyVZE2Bcm1gKFxHkGhrR4SWrMWNcZhqsKatTkWnk
EOLne41MSxVTgVMC9BwhwW9gdUa7ok+2K0jmvK0ScS9vY2hwKHj61Z4Qv/kBzT4s
m5mb75RKc/ZrB7GqasqBas7VEMbC9cAV2nlTIvMIoS7/EOuCJuzxn08pcLsQChvr
vbd0pjRagfb10Vpie+q/uz4IintqFkBTmj3+Je3rYj+BB2sCWPIv5Q8kR/J85F6X
lAF+ykuY4u+jk0IvyNH7HK+8+WsnDWBkwauIKfnjDZa2O3g3uyEspzXtOkDhiqJy
Tgktd4Wj3qBvzwzZvGeUl2wUCsk2SSdpo9+SEkz2U+tXUkTlebQo75js2lV56z6i
NzlDFTcN/TOMZpNDYQECZ04EyuxHsQz70NnCt0nxuTDoQ+jNfWM9Qumn8GZsLMRE
`protect END_PROTECTED
