`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPqaBw4SNLtp580EyycblETDYX9bc5iVeVh+M0r9eAyUezzbrR83iXJBWadz2u92
KJc4Tj9UTJ8G5hFoxfA5OpvU6RMBCR0y1+iyLBKdlPEVQOm06vhTGp4gid32C/CN
6RSSEscKEiqQA+qpZhYgME+QFatkup5s+3VbmuzeEeBNKxpQDE7iUSXYNYMzSt2T
pRsy2BXPMkarwtF/28g+2c66wnBfgaHhHsHcRe5sBZwHgWHXS1oLllm4DDMk0ut2
BkWPA0NAxJr3yy6WNwvTePIyZuLaBHeCTj0x/D552+8yH+8iOOUTgmd6Ro+Trr/F
eyKGO/PF199qOsB2TTupsvR/JmqECDslhZ5/9INAHpzhuPS8oyDrOX5h3M11Lwzj
xZCNSQtGtbXlyk1dm83A5QoxPmEZdBMDBP6nvYQVk35+DtW9DPeBQx62Fnw5v2RH
0yL9p6KQkfJw1vaz7Nr4b2he6dT00bD7zUVDpJbMJeQ/famnNFAwDlRsPIXkGk5d
oZinTC2I1+aMh0qqOCKE/AofFrMsNsAaYncKOiuNef27qPj2sGYHPV8Nd5GIJzKf
iODr6X5FnJj9otm330tnkUvQHipGsobLNq6KFxDVn0guU+o5kM+q38PKfFqLBLU4
bAdLbcWBAHEdtBRUpoKSNRDnS1vH+umKP2/c7BCcsp7kXrX0uK51W37ioYv4ANFL
OKsNAfc030ZkSaWpfzFBsvd0GMqy5eqrRJNacv6aJeDN0mJVz/gAK2jGBxFNRX59
X7xdp+W4exTQmF+Y1bCLXdbNQ4vNrz/1UWohofZll/nXdmb3ojQnffXHqmpgMvuI
tUwyLXeqwgsx74YZn2USECRutCb+dsjqVdHYS/zURYTRuA94EChJHIbz5jcSHzB7
Bj38hvsaHqkmg2s/5Qpnfgyi8YM+cqCmF0Y6jFwEIMp+9BcCut6dx2wRdI2GScB/
hUTrvEHk0QCqrYoBQgkZ2Ld2Whw/DqC5kzcPONVW+/PD+MPtTe+mzuHCRuXQzAmD
rGlLLJdatA++OKsUHtWIqCAnzJ8Kt6knuayk8lT/7w8i43rYE75Ozs6S9JmG/sFN
IggGGQ3qUATUUYY51kuFTiTodjgZG9i3fy7S45ImwotT7OB6Rg9FGR6oNxTEM12H
gfiCw3G13FJG7YfnAmOGMGy33qdW39YLAXLpYMHOj9PndkA84FqHm7iJYtOZ6iui
sQsHOP81xsYq9s4a14UUj9STrfFnH4d+7iaHriN7viMUi+qhyO/Eg9XvQQV80roG
p0Rj+tzoaJBznCrnvpwuLJD6yQwp4AzHqX3V80ximr6K8EVB06lfg5qTcsktR5Xn
BnIZSESYmIXPHqZpn69L5p4PAnLFiYdF9GJvslQxoW0lRr2XkAWgcUmSCbK0Mev1
gnmZmXxemaEPPvFnsVQf+2zojEr5N5GrNd/uTkryjmDyjMovN0HMmznHA39LVib4
H9Z6hXN5jbR06rkHmAwhouOLWXP68MhaN9RHgIkvh5fhUuljs0Icu0OLy+XiS1Em
lVGJeleeqA6GQkMkQafx94Lv9U0rkbPGYYWKgE308Adi2FBx/b5VZUwx7xmEpa/6
uGpirmkV1DVfMIFAbAT1tSWVbNxu8vs1jGtuPcTJVZ35OpCQ9OZ/CnblxuahHX4T
/o8vYlTtjM8sUOFv0OF1dLxkfc3XSRF+6UjbxtVfA+O51DCYEP4EWg/TXFKVOCOi
LOKuGMp2uN/KIf+WSYxt83pZwGXo5N3W6PiionRWRmvaWKn1FKmDr6/TXHBVektI
6kGcJz0/1zMU/STguPq1jzZUtJCcRi2p5PhLRxPbclF3uIGP6/qemPC4n05RsXwB
PztA2SM6fojBUejhy+ufRagHcxhwtIQHNhUiIs8mwE9GBnnQZ061nlsBU6OykE7X
6T4bwq7uaXu2hdT7+dzR/8mlkHFuwHYELzUQQo+EjAoGZYljKB9h5p6dFyNj3O6I
FBBrxufD8A8mlVGfVc2xAyFCzltttFWWRxf35urgP43tTfcBqNx/PdtVkDGpq4oy
Vyn3b6527xpaPbfa5nTXoZm0pvo3ONuYzJF6CIH8fOanEFz0SQlcOufiqNtHlIYr
J+a7CydwENqqmTznryo2eS/tPSQL+wqaRmcu6RAdjFUs4U278jh3wJfjQUC5FOYK
lFXoXFGf9sV4z3zUYivhq/YHa+57vY0cuXtlTTkti30DIJ2qNp8JrMmtkYvjusE5
05/DUDwehB0XIehgWbpXqgpZcUjk2XjKWopv5LxykQjUJgiMj6CoHrAMscq8HWMs
9IAfPstiyhAeOxkQW9hj3VGIG1nTCfmEidPLfxh4DgBIqclYpIexPagpl4TRygdS
E0ZEOApFR1wb+strVg3PP6g4UnvZdQurF1yim4kUSZDIYus8UKCq4y8gcj47ZHB0
+98zYEZJiN+cXm5LLX81VcxGvwjPUMwVE2kIv0hsJ/JW/cfPRAj+VddGwvK7pOTn
7rCSzGkazHkzukmBGqxyyhJaTl8Zr2bXZx3ZgPK2j6v9IwwbPMrfrXJ/08wSlN81
pdcU/rhFnKLV3Io7d0BrKBzOMzUxcJkPo+p0rbbOf77+SykAezUNObBrtLqLhNCX
uvCbiBQ1xQi5mImaNSUJMwAVAa0zQoeIfDycZ/HaMmJvLK4hQcxOBJe/f5EvLy2v
tEfQTaQb+Bd3QYaXsGiG+g1aZFFFmCRo2t8Ibs2zhl11ovAj+bpJ64R4dbaMooxL
aLhnsNE4tiKq1bb3oEYOAZagXTpP/+5jD6vXWYyqzrdB6QGCtLBolGebk3Rvb4LQ
cMRcI4H4b1uKsRoqFXZYMYidI6CSkQFKIdBYAIxcBklGwAOYg8gF95jrGz09VTXK
n3gZxz2LySjbSWpoCdLShrOBomXHQYMf6Up+JnJtTvbFw9I73I/hG7mxcNbldERY
+4slaO9A8GF4Qktl7qUEMc7Vi0L4p9QzK0Sh0ZPArhR/WxKJ8IRweEW5p1t358Z3
uOFM4A1cXEJG3iuIjc6DEz8S68/vCZInboEOuFm91VkDq//JB9vTio3xj0mvIySk
ZNJUa4I/nb3zcZgbi6hoEwWAPp0nJeTodfGSEWuiInO8jjEls0bVCVvM52GOYVQN
6x7W2N5O7PESrzbD6IlA51e8oDPOgEYeBU5exwuGwp4tlKsflcTkFywX9Fd9aGV8
nr7Az2l2XcSZfqn18moOWFD0y2l43tZkpMwZrWOqmrIcGhOBnhmyY7rK/P2k+0b1
6zHcSubPQUoSPqiN3pIzqg==
`protect END_PROTECTED
