`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VpH0iMQKQfrE/QiipdNesqZBltJpi5FiAJt5j5MpZh7Dhz0/KqLyOfBTPpnwSdy8
yElpq8e/ANldlFowXF2pKF4MB5mQIDsFfjzER2+8dxAUXTgv2rL2kjPkzSPLBJQz
RrDuj1hakd6aQiZck9w7ekfbAq5R6C7uyBrcFGAQsjVWVUREOvZwT7CNLt9mUtOm
yg6GnSjNSPTZ0toIZkJXnZmA3gMww9/hPDYZ8D8bhhiBocnLKsQzrLkS98oButjk
dS71u53jJrg0+tjiPQ2g4XUE+CYqDvEpUndyk/PogWKNHkBZuvDSj/ic77vkR37o
vnilVaJ/Hb6MoSSH73tl/pbt1mfUF7SZixg3o31pbGNl5saQsMwvrRbHBUA1Nmv3
qeYpQU43FYubeWVtZmCvDC9ni4YZoYpgyGDHX0WUO9heEtf6gxroCzL5EbFN4D97
`protect END_PROTECTED
