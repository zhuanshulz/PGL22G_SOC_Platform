`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGUFPGYp5j1ybAfCCdV9vZ/lQSsWvDS32wLLvl8zYN2PkcNuB3nN5kQLyt1586Ml
NCDAPW5LHM5j8ML1dhCXrUYkmchfOPLr611CRYDlXNdZSxEsOJ6TcpfjktQlXF2T
XxDXu+mVCwzl2u9AtpX02LEfKxa/rxPU0GJqSNQWpjpqbwRQ/6dczaUNwMaInoaG
VW0qFYKZxLt0Tcm44P/0TQljus6rd6N48WkAcfx4FJ5HxvM5MgR7uhL2frbBh0ne
3LYs949rx3r557vbUzkVNzHlhQ6CLMeBuCRmy+mNL4jPy0NjqdsvQRnNGT1bRdAB
iDyfVkeQ6/GOtgsrRy3HTJbGmJSkJ8cv/639Ua+bvNR59i03HDgthnvSGGvx0Hv3
2iSlHyZLEyMbMMYAYEZk7g==
`protect END_PROTECTED
