`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q++o3BNZXhOt+SeUxEI2xmJvVVqDMTbYHU3yM5OOCgdLV1pfurZYXRuYoY5jbiaC
WZ3gxMsByBM9qmy5cBmlv4FkiUrbPE9hDiEcU1L4i4UoTh4yLC+JD4TWmF93mRaq
i3/GePcQxep5mR6UcAm+B251G5sOAgLCkcfvbMnCjxjHW5IUnDuLQfdPnWvJHXbX
qXlEWsLwGKNe7nuMHLettn2SOC1Mnp3Bvf40tKGZs6aK9VsENrM97OpyfJFff5DK
XuSeylvjHRuNP7gGn77Gw1YTfVY+KE9lJzrrSF2P3EByf0/X92WsDhrfeJyffqgq
4tHS9M5IybriYm3JC6GJgsaQ26OlCCuJPzstQq0064FqO+4fFnFiVk9ua+76qppv
jhh5BWyp5yREuXrhGT2vmIDZTJqu6MJYGAdbIvKNxc05r8K+LKbnO2ImgBrw3U2X
SdEpvGQj0jd0pJ6EeoAF0D3bGsLNMfvwprejuTYsg8bZIr/n8irpLj8H/SpFyuTF
mlGqEFMGDku2u5gzriVPHStsb5Cj7Pne4C+pEpgFrtgqks4w7VUhgJXL8iJ/bNua
0VD88OVAv2EyTob8yTEobf28U3wjr08g+c9WjdpX3p6UAv3IhF2Lh2w4UKrb/aUi
IMoshsftxCuyvZod5/5nX+qWoBdGAljrKOZpCWouMevQBCzSvWVoVfNjPz3zly2B
BZ29BRDyJ5sUVHK8MKHJHcwx6Ah9Ta9dQUulk1wpH+lYvKr5b+BmAM4HJ/eZPsC5
CGcIyK650TJoeoypstjeIznU+hVguA+tyKQS4xU6eF3CNsBGLK7DvWEnLlt3R3tf
7mxT4Ugnjz1gnc2QFNPk30iOdEoF7vSO4O/HQFRXTaxkaPo5KZKKJeCCj1xNCBE1
Ey+feuo2eBLHVrR8bvta66546Vn4HDW606vFQqJSt13HozrmiEsVKm3sSvfYj8mM
HqsWdq4jJVuM1+NDfJn3vRyd1S9AgaM/b2LVD4pY1uN3xywN8d4KD+b+mdDnQw3A
zYb7aP+yyYpSzqEUtXn2Z8+SPxzTgtMEzsn0qgPLU2qzXRtbzyf4Cn8RHdWAaOST
XgQ7SKreCnb8HlEB1Pm8GyuYj+FGhDjijMwcfFM+Oqxe/YJK0WmwfGpjcHuK/fSh
Bh4zBkhJTvLsQr/qbIGRe+H3J4u9JyR1puvakmx6ETolwLDYHYLmAyXvIS58A/mr
ybiT0KsLtiSL2T4mczUO7vOZZZ/d0eT1FCd32sCUdeUVX75eN01QrG1vaJxZO1aX
OmplWXJA5bMCNgCsJYKCD8W/3W2gKFC1CwODEgd+mHDm7IF1ZfmInAMeHkgCeCfV
UpJapNFhOfKZue6Vp/cb6aqVp9Dz+xJr6+wpzqq6ok439WZe6WGzzc9jbGGHwcRV
JMuINF/usCrv1LLMRmUclooseo6dVdyCvJQeKHSJ/u3EkGAJGsO6pZKNOu4Cn/CL
wNz80a5+YhKXPmKkP966pnxwSwHfd6uFGFrzm9wcFDCwhFXygi5yeDmJbjWO4e8b
PRPlkKcy+QW4Znno/L5JskD8R49nNsRG4diZUhZao1yRjfRYZJCFze79Pkq+Bf5N
BpBeaxbbBCpEUqRrMti/3vv7JMamJh3HwylcpVnXRL/KV50WcC98VXnGMUgiHK8S
r3vs4HJN37LEuLmAdpHOYqvZfpaX8thM5jSsBDktCA7kmzC4iPjIVAx4rHYqvbxm
tgEq7hEiV+pPX7mXWhwUGD97KKIFd66q9OcVPUxsj87dC7ZpiZkAqywDRZX15HUO
DqVX/EmyF5sbien5d2WQzPrJW/7Mx209Dadvx07+GMTazbmn9dJ7SRR1oYUxXucv
X8AhJlyaNeZEWQgAqIoljUGqzecNrTu8mwRdOjYF38dyKnkEV9Uv1LDU0Kf2F75o
wrguU5QcaLqCkTwJ/XExMHBm9rjg2XtNysjf773M16s=
`protect END_PROTECTED
