`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCTSp/69NZofqqM5WpPgBd4MvIVme4jssV7ATatSfMuZWcQXUk44CaKYiG3tGefm
1QoS4IngFPH9k+GXrcSaGXpPxJSg9ZYAGsuS7alIpl0e7b4C8T3ZrXsxIDmXZ0+/
kBC3SRhS/ra/KYRmsotZBmwJt7jF2zX1Zc2IM7iSdcolq3vopU8bzIOvNLX+VrRC
k+lv0p/g6Q8ruFXAqgXJFtoUNpKSpJ7xu3yeCvxAT+y+Vkp6E7mnZOViRJUanfEp
ZTNmGtn8Fvv08fE6uR3HdMIVjRqZ/U3MSIy4SeHTCPpwF95peI83QR9g76k5EZ46
TBE5F4iDSMjsDXrcqLcEA2iNyxU6+al85U0UknI0Iu+8wgZX0TtwjUC2+1yWjy4w
EAmPQslUC1P+iYLOZ4X9wIU0emrdu6MFOTfa8DBewgwxdPGfzfeDmO9aRbFqSlC1
3WOFVD+iJ7bAvzhkGIRx2bOBKh0tZfiroyrX61o7kwFRbTeGxtYwmn1C4DOOFic6
2z84xbzkfbpT187+H69uy8nSpx1xlDelrBRdMn4dsWzzn51zhQDNMGw18b0v67dG
eMhIPBLpHF7uJgifibjG8tOwbqJ2KUTc1+a7j+Q+kfEPB0kJm4PzjPd1DT7JUC9P
MXrYe59JtJcI05Pjh7XvAjuqrwwPXDm7Lr3+YPcgcR1taWu9cq3i23kBFNW5W7n1
GJQyNv3jqo0BmicH3TCYGwirgpTi45ds2jx2qVFM4tXEgpnD6LOnzPLVU0uQNFRh
RXhZmXjmy4d52TLhg6YfLZqIMokuor+MkEQQjUYgwh+UN5WsOGKW91CMOcS7Q5yV
FDuLEZJNkfneh4zriTz9jEJ48AfFKH8AuPnWvZBuQNgthJHuwT1WUexBXwS/NHro
sG+OM9ZOva6e1JBT1G4lBfe0xWfujdVL4nRG0ybL8SFeDbRB4oeD7yT1dkhSVVIb
8DoHHzqyUqzhcIt/+4M/55bowiUYcmty5VP8YdONMmHF1DEXoBio6BSEwG4eq/R9
vv8K4UtylSABsFSMKhirYSTLsoThaDKO0jkjJiPvlmGeH2LvjY8ncBDU+LmBJXMx
FTcWsa8LouVrwiSuXA7LX9s6h7yA7KqBnYX1gX/GY1Rb0CPE4c9p03s0QRBf40/4
rAjcuBFwrLRfJMwwmhIYNNd6gIN3pP7bPFYzGU3znwF5m/1m2ctXu69IYrQrCcpU
7fr4PCHkMjFptjoyguy50P02edrNQu9ajjD6lH/PMNadfqJ4lCqcnzxhHBR/rge6
FvCpEkUZ6zI4EB+3QQ8dxUfckjBqBYpIMxc+q+dAesNqITgPoMva+QBHJB/m6+g6
qTq6zNss7x37nIWSs8Pe8otCiAcZtpCwVgKQWkc4lMQs2Xf3lVaCxVpP20ASOszh
VD2/h5fr4s2vBYWXrmhrL73VzTJctxB2HaUe5sIpHc+Gu/tFd+mRzpQMBAcWWRba
2hsU8U0LxscuOgnp0+YkXHBZY1kU4k0Z/yOpTC9WQfTYFOL0chxGAJCjW2R+ot6N
CuUvWG5FlUUq+YRK7JrJ+R16Frz3VVTTe5LYAiXfWcV6gcGB64uEpjr6a9OY+NXT
O0ReneCgoi4+eypOjvy3IsE0tDNs/gNJJVCKyE8JRzOOSLbIxEaU0mh6KNi3rUgx
+tHaZc2u7UkoWr6Kx6RufcjkVcYXasS0eEJdvKo6WhWGgDdkZmalkHnG23Q3G91F
fGd4XgpaZ8ieSxtFtKxeSjqzToJvkJJ7uc7gw83ISyStD6s3VPJa4OfJZYD3/NMD
0uv24t2gd+Cgiq/I/jemruknCrygYd2diPPkch5Owt650RuHXe0CVT2ZCv4MgYc1
QZqdSgxk7+vna0simDyPfxqDJJ1dqcitgME+HVBiG3afM+Ir82o/17gpRj7xgt2H
RYxp4pOAhhbt/hIwWd2sX9OWJZ8dCOoGf+Uwu4PnLheEcnSURcl/eI3pF0LI4cg3
Bx7/EPFoz6exOPwu4nX7AKEPpWJpL1MBeTxRiRTGEB+fuzrs5Cam0tJoNL6/JQGv
gj1MQjTzMfFBOtJvbterv38fHAaoVfeoHaBLinNdeBQ2QDuaz4jkDjw3WuaEISIg
JPqhBBODOs58+Jtzk8qDYFoF9AqmL5e+GTHzmyPNF04BQDVihUXxwsAmzXhGhucS
cQTUpIWos00mpJuGewQ76wZ69qZFsEefstZ2QXzxehg19y4eOibH/KcW6vrWhlKS
HBC+9juGfYqVOY1iER88pCNLaPpBq5Y8i+BYjujnhiJJVjI9tNHZKDF5WHxeVDur
woXn57f5P4HPd8g7mz09F/K9mPnU1SpQXKKswn8OlusQ0rIf2zQ3ziq1y0JKYFny
8Aq4H2EDXb1UtNnCuwCsdSO+0cvp41JWHJHcT7UovF+CbaxQb1uIq6T4t1lBHn3I
O7Z5FPdcCbf9o1RE1wAh9zJcGCW+UCrYqauY1jV9tJ3Dm5kP5JVgy4WhYbEXKlG2
Lq6O9SzOlWtkLXiSt/8E4dr0QRf0ZtBn2UYwbFS/le7RNSSMSsfFEu6/Rk/E8716
MrfEi7VJ64o4a5W+71K+MEqs9fQGHze+YQ5Il+rj+IDIWbd1FGBLPmwE24qY7ix8
Dzpqokyi7FUpFyaHlK+JFqQ9/gGhP7AC+YQQmBvnaDMQjJ687YHFch82uBl1hcOG
WSJLktIUhkaxUCuCXE3XIltJi6/BeV+uAYc890PYE4rKa64W3BAsJqMHzEzt5QMx
a4e4CrSzZfxZQe96FB1SdGwXuDELUwnqn1jHMqCt+WMBarbEjJIE43ejBEGBr9vL
rmJ6U/+Ot/yGNcpMRoH2AB2mr8JZXciw2k7cZQIeX8qsuMRQTCbSYHnD1LdVspZI
ZxWMKz8wXoNfKB/fICuu1H1QbrcW/h5C4IvYfOUQzMrXq/EY83Sol48Z7qVNgZB2
fWzDmMskZfgjb3r7fX8ghipqzIf/OWdj3jHm29SO13YX6qHJY3a5CzESqMco8m/d
0L1ZPo26Mf+JVgfdNnJyXKdBPZcZdo7eF9rjAH8i7WmdiA7m9qwZhEOFMLYmZbV7
UFGaBvOs76Jg3I68wDUPSjfNWJYvl+rrA5Ec7ubRANThlY/b6aAXoPxK0dQowHcF
mNRFMnH2Nx9yrZAlbKRZQCNaDFA4vpOuR4lGDkuUhF1LIxynOHNoaAiC68K0k6Fk
UaPdjBk2AWBjFxoOyhRsFOYuUk5tIbEWonld/P2rWtkIqF++uJavwSWo5fPtlDEH
Fk3I7LERRh3uUfmc7WgQoYa0PfzrP+uWpap/qaya2F+F81BWLXSGKnx/33W5+f+8
Yx0wZFj8YcwoC8OVKMoh9tMD3um5i4zA6cDXOd3c7V2vGp6Aoycgs6qoLeVaMZN3
JD/VIzyb/clq0K7C+dRLxLyICOk4d/S3+pnsoscktN/qo8uH7BnLgHm1qTevgqQ8
mPfF0VXT1hAEAJlV5p+SCtSRMsowrayU9nklrrUZnf19SNClcIRxnYbBKXZ2bd8X
JONZgFv9bJyphgWPHksOhiFkaPjJbOAFuzA/Yr8A/pdYWimjh/T5UNPo3ZsOALiL
+De34KQpkY/TnM+lZ64gHCC5RcMqM89aRsbYqT+OgkUMc9QKDzu0lgNWZ1cBdJ87
3p4xKgSuD6cwhSGIYee93DC/nTWPBoDOcNb+S63UFoNf1Z+fnZJuH5gzt+tswPzt
D/mvy6UQ38llRTTrfyXv6CPQz/LAGDP7QzDdDYrmIu/dBoVLyVmPRjIOv+6RdL8L
Z4kDUyuVlV/+GlvK2J8yyTSQEzB/S/yS3Xdkx9sRTnhdQtHMw0gVlbo1EOj90gq3
Oa2+BbG3f3vQdcUskrgACU84neIENASTUEUEyI5DsWYssczlJiYuIkysKikTKVmA
3Z7J2la0bpQOf9E2uk5aQsvCjML7pXWrmM8Tf74SzopyiwUvqifAu7HB7IyWo8hl
2nxnRFzGoIFP7ouNGLmegFIxPRCvuzNmse2ugbJ+fAAFRFIvvj86zcsnNhu5Vokm
oe+ZaRTlRdaXGo5XLhQRC+A9ohJdDelDnRbmFsRNxORV89BquvuXkSTKv2rvQv68
/cxi2HBVEvZ4uEHi0PvmJngQMrlzp68gg5EABi/GT/tn37Poe/Ry24EV6Gb0phr9
+xJhFTsAcXMVfbfqJ7W1xvPsrso5TZPOaAphbokzK4E+b/lElq7+6fxGF9xjEexg
pXAV8wzB1pe5by0WjGNx0OPCDLvdmT1+pkuvCryUODMf6Hfq3xLJQbetHyt/kTpC
WMkFuG0PVsmGUghLZH8Dv8yPyHA9A7SbVhtAK9kcd9MqfqIpVbEJSlLbFyXxqS0l
NSTt26gSOymETOT0U0VwOTajQQ57SaqQh3G38IZ/Kzq+R1K1vUsDcBwjY7nx2OnP
P2Vfigv+CL/djzdQzYKjqhCg0X8g22DCLzDPpkpvEqqzhDD6Icv6wl6YorFf2226
K4Y18Zn3Tcud7bx69FYPZgxdWHH0VXM7FdW91ZgTaj5Nd6G3FB8VhS9nBvNIGbrv
IC0pdbseAF1UVfWKahNT/k+cO9HjLFxAY2cWV3ZqhUzRORwWhNfnWDYirseh8y+8
WTKRMIHCwDSKJZHyJFqFWsxHnPYzFAjcSWmNyg+ozHSy2sKzBIo0b2f/DFDoO+yl
7CUo7yMHAwXMmpNVcZhgvIf+ffl6IO2JITnRemvR0pZb7dD1VK0Y6FGgcO8dtNva
IY9tYouSAZqCWt4YKeOriKWbjxLpY2gVTc+3Rq7cmm6dRXYy+qGR4pOSeowJ0652
Sgcqdwhx+7IGXwgm33IN/uYTl8ANWWgyJcXOOALwKspfEF7Fl2FQq+qIWJ3MDsf5
GqNQR4kzyv/2jPhvJ2sAtKCv4bYYb7TBYjMsRuM6U2EEjsPskRswI3wRbKUoHHbN
cazC4KIIepXBsam5k0UxxZd1VoXqcDxFLd8QfJKKr0gb/1G+VLT5IPSaL0EF2Xyp
KNOyKNbcB2HntNtHxwDNdMETvaEzuwCEQS61NUWX2FlHLSJd7+ooM3E3AJwAwu+O
/xWcpaT4aP3S5VB/U9whbbaJ5KN6t2fChVoh4AaeYPSuXwlT4ugQZzwMQBnc5PHU
Zt2EIHSYH2PpXSOnbJ1AE+9rVNScGy5BDOZ4ONyYXr86iodw08seotk+zSxj79zz
XH689LYNf/F3i0VkW15+ffKrgor0YxvAWpaVr08YecHn1F1Zhg2evfeSOuNdWeVM
rayb0E6MoICCMBitzRlFgNIKtet77H1K09aO6nMtqXgfbcs85hxFbtNQQdAyhC/k
XiSfAi3dNcLMImKAAg4K8tk3Sjvuq3zAJOjixvz2bBeacpgOVwhw87Fm/pZvdi8B
ug/qaKpF6FlBZE0cLMxJ4OShqFpWTJrJImmSBpJj1j9mUMmluwYerUgC9E9eByj4
+1ynMigEzTeaWiH0HDNxFqjbQlZyC2JvKeaV2N2oy+9+HXSXEoeNxHQ4GtFlw+CW
IOUbZ8QlgXA79eaXh9kg9SFKTltdReZVSWvLKWaml71ej6v0d+/ur5Vv7Uraizga
YFnLm6rui1mmEXhWFJR8Lh0FWLWhjyiJcSENvj8zielWbyMmes0u36Kj7v8z3209
88TKuTAafSmMsG17/+2rRPT+GNvjs7Df7xK2OvweSxoskJsdEu3vHaBr/yEKTBqs
79zUd4oOk5pgj7NHfFo/wyp1klbxmWdQcchm6GLfE15Gi7sgvh6usq4fcl/2l2GG
83Y1oFpkEOwoqZlF5HvG9xSdri9WCO/LqBHqhhkuLO2NlSkodezGRFMEhvexZXF2
Ien4gTxhWZsKVPcOYpXPHh++D1Zh2e/fTbZ+NFbJTP05hwSIJKkTU/VB34pKZKsX
+k67OrlZhc2WuHb5zaOaKtXkOxADmp6pgsIjAmY7J2InLtC6w9yTwK2mP08rJX9W
uPZj/T6ELlau4CSPo6qrCn0tSA9rB2/iOawHKVLIxaj6GtyjTBHv6SHT+NX2dXwQ
gVWxTj7iQ+PhrgI2zBoWx+AyaIcRR5A72zuc6fZCMkizZ/OOXUy9m+6uNPYInerx
VtOD7SujFBSbtFU7f++ZPYHAZLNn1l8vYeHigDEtr621Mevc6M3/AdfHHB15nMi4
CbwpYHHQX/aTl9+2IMBkUw4pDSWPCXJ7rV8UG5P2PZqvFCpE14o1A8scY00+RD3O
MPHfU5wR4YsWmK9ODYT9clBhbZfIze4YVJdmh08kV/gMBec2w+MFmpAgViPtptpS
usPRb4Y2A30P8Xh+4FggEBqWul1K+hLsWF0d8LvR3dRi6Q0VQEvR927kt0qVL47R
Fmsi6rZ7AWubCkNp53iQgd1hFmkEu2AF2i0BLmZrRRAmj1g4YsWkljhAJFRicftd
tHbJewnIgmJH7NZwYqUm+Zx9zyLhb8Vi0x31lmG+QAoP19p1RPZBBNRZ+OxL3AJK
ka6+Gr8N30O+1hW5BruddmJr3/zYz+bREU2f6kI/+Vwo22zZ0mh3w7H0u3bwam3x
vIOpeGtj66UrLv/Jmft+QMpxcpkbD9FA3xBodK20Qe8taHyLYAVWcXs+tJJpwL3b
gKYr43ZiF/6cIsxWD/kcK7XpOvgyxeAyPuUPM5vc0PDRumThSvJiF6rZEHpHErxO
LWZ9bka5E6BZ88mTwmNhJxKpdW7a+4Vxy8TfsHldpvrjRVBcTEE8/6gcmtLMwuZx
SO3o99j7TEpN8kLljrPHIA02RCCgs+DARC9yB47ybWRYucWAiyH2Bv0CYvORiOWg
cHlduuKbjAf2hviwzOVbYWrp/xiDsKhnr7/IRsUvIY6C1OoHUcxuPxT2crt9oFYi
Zqyko4EFrjM4fLyKvfNqPfP9GyglZeIrNmR8n6MSMyrnJ/Q/LOCAhxZidPNux6Xq
36SGuP7FLsaSy9QWVbW60bB1MNw4OjAOyCeSqlfbRW8SP+d0tpRcqFXs9w2HK5qo
FDx+kCXQ6/BrLGgaByk0lcyqzQWNRLlydkgsfviM2ZSMPT6tKzf7pxnzSpMWmiTF
7a9M9gpqch5df4Xd7ZO5tRvgjh7i88wHdNIfy++5dGuN8JBmxqSCgNN/2oNowjNj
u4aXDXUEo4Ct83gb4uF0umlHNGm7xJuSzaOfPhiSUSYaKxbiH1zNam7vjK1e1mVV
3lQJNnq2cDZqlNKJbTcP235dxfs+85zllNL3pTJ8rIk6fQAz7GoeM0JOZ/SCWVMm
Nr5ej7zVkW/vu6tgR40LIP6T7d7T9OgfBAQBSQmm4I7rR0F0YlaR86v2QXoF29dM
2RuskPxDeDqJ+DEueaQ6CE9IGioNomR8ZllZ5DnlKOXnqarDCXJaKNh6r2WQkm8k
DxVQdG/OkTNM5Iw6sjjWxk19AOAoEcRlKggLUkkWopC7PTb+0SJZqQVYmXU76zbe
l6TxTqY18Sy4f+crWGK+jEGuD1DcxTNU2h3EtvdYzWhH+/5+KR+UUjVQuig8+Hsg
F0Ppm/4xvguzKNbsLk3Gr55gYI2g6N32wOMn96bpM3j7ojmHgLenzvYxbXP6JHJB
hKTVXhqQAppxQu0v9iXloEkxFBzhXi1ndp5GPCAvL3pSj4ZyIcVe2hROl8AE+P2Y
KZgFOQeT7EunsmP1DL1BEA==
`protect END_PROTECTED
