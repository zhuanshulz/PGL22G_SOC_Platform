`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fw+6u3sHHU+RNS1DtHsQSCoOdXWK0untZorWHUaiRauqqQ6uldW6yj18ISqVvEq5
OqIeonEQW1GjIoirRJksS8MtJulqoL1gg3U9PlljD+tJ1cQlgrMoonk8KdM/e4dI
Gk8E96zQp+gtxbVXjEDlO9T5wabteP+OiRuFkvmlJ0r0kB88Ixc2yUB6HQIWbePc
jODG1sAKxTJoHWyIh0f3MdSlftE2xoCUZycQUPYzI0VKzUHx3tgbotk3pdF1veTi
uUzvkIkY5fHcW+VTz+FqdHVo9qacgck4+WzF8OanM0/Ix361fePVgzdD9vE3uH7j
3XpR6Rcbv5SwY2dCETYputPm/qJYjGATK7NhpRpNDgBwCgvocdt7CdwfzB6cDN8X
+VhLmx892cHKGNpP3qRBKNA4p0XFD1ihvOsm2ryoB45Vybg59EMWiLfvW/ZqOLQI
m6N/dLfE5GLCmR2VDAXShLaasGaIJoRJU1u5yY+Qe4eSHvOoNWbppQComoAbexUx
DP0kB0Whwk4Dk0bJ2l1TVw==
`protect END_PROTECTED
