`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wW9zl++egJTU/QD6CzXAt6y/TmEbs1n36nOMHQi/K2CuFlTsIlBLKW/EkQuTlUd8
iR7A0fBx+EQnPoqjQjIpoOnKUdWBM73PpoECDPu24y4IiKeX+iJBlu6TATpxxZ6u
xIDEGCkx6cm8tvs/xG7JAWaRbdSBSFwUW2sKQ7zQ50ZTMWVGsiFwt0lKQ3EBn9H1
rmQcYiwC7raXgGOJO1owf12/PBI1RLEdifFqK9wC1elsC1C4Jo7isuybsBM3u3sQ
OT03PI9UQfYaDoWoamfAnW+rLKtl3RcB7lSR15FbS0FzlD4I6IZ+3wynvRpPYS/S
S6YR9W8eLpefqeT98e0gt75SqKAdQtXE5UI6G4MWlwUNPngkfIOZsttQKHz+ZHle
dZUeiqXKQauNQJzyokJWMOtG466F0BJZ0//HaAclcBppX09QqgAsHbhSUZYz3I86
iL5AcG7CzFZGvblgLfRBdriTZHLO01xnM0huZwLDJ8hBOE46GyruDs1cebNV9igC
5VUXC263kVy/mIRs5ASkltK2lqxxyZuKk9utxMJOLyNmXMtuWzoxpAMwtSjkq3vC
lUz0ia2CmgyfUsgpxckREQ==
`protect END_PROTECTED
