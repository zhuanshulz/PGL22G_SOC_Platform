`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYNkzcHFoIO7EO62BnuPfrdwed62fwDPnJCA2tl/Zvmk9h3GLOb2+GlYNubfTgKU
LSq6Tb1aXQ2cZ2nz9+az+759qrtsA2VjlWJbi/xldeANpzYohnQs53fcWKzf5Dwh
uEpUoPamfoqV47J0kznpy/moGzp3H6MjKLAus1QNbkGH5gUhvGwpDRgIAgoo26bV
5XoCm8uj5gki4FufYU2vECqjktEnjRmmRITuuV5MOHxIGkJRNNe3qZzkn0T6w1ZQ
WWET8xrrwbzpB5gaUta7QuftX5/i8/a+NwHgU+Vc+RDaqV5ionkg3c1YFXVAwT+U
6er6aZ7XfX6T8wqVAe7HvLVw/qd3AWnNz/+C/uiqUzMZhF7c2KL5cfOMPSsdeC2o
XqkqIuSlb6Vni9XvEGx6/npI87BuUfvZCxvTgV8068btu5gNbS9BfVBPBhCjn/3H
`protect END_PROTECTED
