`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8I48h7/RQPK65tvieUvDoU1dE6VCrkz/SKbYNEMCYWIDmNpCTaydipMcBPVWBiw
F8mWRPj1iBfg/nQDMUbjG9+TlabS1Mqd6lmOqFZ8/ibqJZcqzJvU/gOxe0SXV1XQ
+3+zqt4dCpHEaskctkQTQWfsCG3E7UqrlQsNJZuxR4fiVXt75uMlqIxeYm2tqkwU
Ay6ioJtv2sV8hdlXuWqxit3Jst7+t519ZpufMbtlinLVj+8jWaPCiNEIy4Qr7B2w
GWcKkYZOW64PMkrpjN3WtBUMA6MIrZN1aFljGjvb6gTw9FYeIlqTkoTdIyVDk05E
z/1zu1R45Nm+qxMLg2yTCHrKkW4e6d2IFo6nNqi3OlnVXy8hBTSuo5TWGx7n/ZW3
`protect END_PROTECTED
