`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FmEimZxA9+l6LSV1now3S4I7BCVp34xPahoxR0g8iLi3bhFBd/SaMpH0SxBIxugP
//BphHmr0ohaGdWHr4rDZd2Pu+MS51/GVo1xVipCHTyGsMgAsyctJblqIw8d697F
L3AXTa8YdMF07Xw8CIuA6477MYhjpAoE7CX4wenmtHqq2BHEroKX59dUdTnIvGVh
yblNYW8P2JnHNeA6apCv4+anVLByWaZF4qb/GsuKfXMh01LJNXzuFatPd9Ur+zan
j6G4eEIOutZHqCsS+LR8GhTuexlGCcynpP6FNEQFf2W5G6+u/d6Mu8Zdkt68BbfW
kqrAkaZMwbtybmgPEQDdNpuXljrmv1khMzOAM8GAwTA36v0PpSGbwqApRaQ73JrL
klZW+uJgmXqIyHuSnBjXtznZMLPgil/rZviSgZIxhhGW84tigCf33p0QeU3CRXbG
IntvT1NC1kSjqDSILoH8Wc7urWuipUKb/ZH/lVAxWorsy1jpF7c4q5rMbQ2DEbSa
8gb/9k9Kg/JniazkRP7uOpLApU4MzHwZMCvDBGHRKeRe2dJbkA5+d0dcH8SI2yYj
5HGd3FFKeVYr1JpF9raBY1ezrzNIlQY+Rcya+4A7z+I5omFYzXj7ehZ3JLrAdVvc
Wy+4OeFL1Cmrvgk7IAUFZ3xZT9iIQH2+LFeo9HGNXeMDH1mG5enZsV3mYpna3UBd
zLBZ0iqCl6bI1XSREyuQr4pRK0ulqAm/d9c5ZrkLXlN0n5TkctvsQi/+JlFpZcA8
6Ltor/gg629tJUUBqQAwUsl0PW4t00cq60RB4jFaOown6BRfsrKr5zyEcNT0i995
5+QEj5dQr+aqlZtpTtbOKl5zQ+KwiT5RGQjnu+HMe7gkKE9lSOUK7MZ2VRtfMv5t
ilIpudQO8+nR2i41fcfRuOrfoNAYmnpyrbipN9pZW2LJf+fuYsjAmCJxqXAafFtH
09VPQyyodcCNHwMmxc8zAd8xnZ+I1sr6z+N0CgmIej8HDnPFus/oyWz2rj3ntDU5
epw6vWnd/rlXz09/DBnfEYeJ9uMmsVQx8kC/31NIwLPOd6shc6TzWIkkXI1oOrlX
WUuAbO83eClKtJIEjov5XjBRRNWq/e/oq9mxv5GvgLiL8WEJGBXzkUd04rrdPmMc
nKyOXBXhI02UkXfddxnyDxbDsGoHCBHoTJ7seACM2yFuJWkwchCaqMOD6yv6mj42
YfDzxC2Y2dpWnPU+MDj19OWk2MdR4Ts8A9NcJ+56+ZajKcKErd8JRBcMxVIm6aKq
2M/6XV+u/3Ma2UZsrVEREwFSseyWniyXS2drZBG00qL+a9SmSp9OrCY/UKI02/JH
`protect END_PROTECTED
