`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4AKvMSTvPAuWtqh0e/JOrlzG9d1eDvqe/a81o2pb9g1YnJZD2FdGamfviGYBSiCp
xKgn4f+IWVy0Yje8GBACY1cUZ4pN/cvAVz2IcX11ts0M65kAxzb7VX/aMTSEG9J2
B01ECLmXN2rUvR+qy/7q/CS50Mfbsor5mUv2j1d8XV1bzhIaxoJTrUTcVpsWRXYQ
mohf4yNqWQRp5Q4cIF0A46VH+mbwxumV1iZGkslWFIm3y3YtvxziZHmjHNjb25Zs
VLb+fI80Ki69IB7mVYDX3bBX+G3tXST1z/FwkGIlDGSYN46QFmmD0zpGAT0A+27P
oTuPfshtvSO1twn3LND4tSmNteA+cvdoDLumWCzva3wnIdEPrG1qnyqFF2JIBdQe
wf+Bj1iyj2dw6IaSXdlaHBoCUoPTH1PC6w5icucFeAyVgGUWIUJma3aZ/I/6Yz2X
D3hO82tLRkjBC4dT88d5jO9xv2TVpc9D1uQ0JsRd9pxM+XKUyuXO5Hm45U6N1ER/
6wZaU+koQGYrVQQ5GioUAFOad1lDBIBefpiPM60fr/hgcDfeV4tqz8WhhfBDm1BS
Z7U4bWdtOiA0/qm7mTVXasfqxoKlEbLIwFXczmym+5gkBBqzbqa9sCPXfsSI8D5x
32lMXUsvjbXtHvQlGzSXK+5dUkJcYNIZP9PhJG5mXkHrHZxeHU0CIujYzfu3PeXo
6V+va0BA2GIPXX11v79IGAxZHwyz5Qg1mC+ZsY2z9o/Q/FvRLinys9ad/A/hFrrm
f7egT5t9UwwOwXtFrLtF57kFOcJ3DLMkQCHDSY9xEOZd8RqmbS74JFwmAHTE7qho
t0e/FWQ+CKg47wUnmLX/MvesE3kYUqeJZe5UQpWXhUB0QBWc2Mj3RjOleOat3h69
gPUB/4puXGiHtIM8jcZCRUb1cjhVV2ebSFKzwe/SNNLgD0jSp9WknItV0qe73B5b
m/+5WeHTmzhj50OCKWp3nsstno9OZU3SToBhkfQqnL/CiL1PN9ri2Rslvrk2oIBR
6MtO5fzvx8qX/9tP0I0+JkieHNhOm3sEOpgxjt30f79Xni8WSckHEbawUqjgsy/s
RyX4jJbRB1o7s4oklWhaUshcVPzxH+Qs+xfEkp4HfXCjvXNC7CrUfa+s4NLqezdd
mGbk15EILPxIWj6WM2/6NhqDxTuXs5nzJMuDtNyVR3UVLKNvfNIWX0YxtVLFM7PK
hP0JGWA1a0Y+5IbS15AO55D8g3Flo04dxgUrO3VD/gBG8oqTbdyh8unLwYsNfUui
IfracTOFaC1ttiAtHvbL9ZCfstwEU2xjFQCkiFcKk3EZ+JU8b62HNsOV4sjAN2pF
QnINTtQO41VCoLeLe8FGTKKKFec5rmgLuPYYx1ztQmygF/8enul/20h9EbvBRO4E
x4sYn14a655pvVid6RJ2XZUGA7RWxUNTrlwbIgexx+RTGJBO49iyfb0p+ERYHTN5
8ivmLHLftHGsehHVtoDIX/4+imR4WC/NProVKaCTZylzbNX+4mEHDqxo3RymYpOy
99HSdFRoHtASMaiQKZY2i57EGo0NfXms4+L1KIpLzPBGCtAN2IdO4EGIZ7gwiDqW
QVuYnOHvrZuVdUVOVrJuMnxfgJfB8N1Mj8TZRcew1RPlE/MUA4/LRrxXcRP44u7y
gLgIXqAvjQ/oCRWwR9B4iqj+rali0f7zt81XA6Kj7IYOECqZN16EImFnyUl/t080
C6XMeU8ZZXPIjIcJA1chOykL89AL9sW1qo6Ktb+gqctc8SCCi4NlC4nW3J19BSag
AwgthefBC3WpkmTJCWVuqcRovunQ6veG3bWL2GZmo0a6WH3KhoKIEfHgVRNI/Oc0
8xScaViZV9wGswmb9gglTaE1W7+hbh7lcwMKchMKkSMU6p+82MFwYa7fHIm6YLzI
7C+YVjLNXdj+d2NhyV54aP9rAgVLuMGtgX2r9b1a55uRZ4yvU9ALFquO8pMYDnoi
WeKaWKrw0MG6CxQdDv22H9HbNpwWlwRoa1qkoyM/vc5XE30lf4CZi6LwFywum9bJ
MyiMs9dNyoW6hcsgkbJA9Q4ZeNatTKLd45Ei+UlfMX1V+y6QAyy9aJv8/FWlDgxs
AWmVnWbeUQixdYO16qgHqpAVrZB15cAkEuwh6GizI07+m1uSLdaAS6b5jX/FK/mA
GXdz8henvnAPpTjBt5hp/zs2kxmB32zv1AJpqlSjc51+RBvzT+AmfHYkon8W47VR
3jNjl3urTU7pNmLERRCh34dhdEJ8g/luwcE26hqauTvmDooJnXziPRpC27Z6k+ua
1exiP8joud6qruBvjVbrDmwuSMcXVSsd5Z3viMLmU91XYwRDWkotbKQcR69aBacQ
aKebNPPj2xg5/YIqjni2MOTz/zTYodM5GpmljE39u7o=
`protect END_PROTECTED
