`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/yFDRd5z++qPfFwj27zT6d9M3gcK02OaoXWVw1aZl1nUsROPtYcW2i25R1dH34X
h5nrAESE/JB2yx8FlkR0ZeS0+Czr7vW1J4TOI0QG4rFk3vlNsDhkePoiVZ95QQmg
vadY2YyLMH14MqpDT2rfVl+0IanpNBV+clDzanj6NoQTHDdzdg7i4MKxV+Ra4y1Y
GQbhLtKAp9AmI/ZKZLm1M3MIi0OO7xQVGor9Uw9HDRv/kDPwkZ3V/oAZzNHtzPG5
Nq6swO2LJ1DQmcHIubLNmZ7VADAjBPxFoGuN3dNR5g96bMHkuBKRwVtPACDb7g6a
DB4qCAHxoMc64On9sGD1rEFoRC3deXCSmppZfxJ2+oj+43xnBh3uCM4+FXH9lR0n
Jne+tb9mC3X3AxnWZAQCqCphmrsdAceZHg7cCXyvgGcSmflfEZbk60+ivLR7Ow0w
903PE3iRIa9sLOKy5aEvu5tZAmbEocv4PBwEtuiVUJyJdPSuQBrTbIVITGqHhxDj
ve0dM/6GC4VV4WuO77eg3Ee1WM1OLEnrzFTwwzNWKW9bK1iZmsx/Vo5wX8pkgJbU
IEBsFQCXUeoy5fRDkBHR8dB+bwi/FSHbH7SO1BTt5aD6rR1KCVRDMM6Hx4rVIfqj
WO2oHkT/nJjCurS65Wb5N9O8AnjoyNmDxcKi0rxQoVH/pG9vrf0mRNm5pzVPXQq/
kyY6nZPjk5ZTXxvfMj4lDVerCEGMysqUQKqebYdcRsGXS1Aa+SENM1CHgnpP4mAC
zEy30hMRzo1YM5tdTQVe47FZ3Bu8MEqcEWN0h2fbcYe/5KKpxDbcnyDslsJVY19c
GTgVnEWv3m9acb9jhgYEpHLtOLSek9vBsGw8Hmbcb855u/gdWoZbkoTVcJ/lUDjX
+S/TZRyl4R1O0+q3xyIEbZY7iszBGQEVpeMg+8gI0xabnID7mIKnyZrOl2TP/zAu
X9zSIFBfmSqHWG4P6ZSrUuAJIFL1dZS15JkNrVx/dqOm8RUPWNZPuAKiO83V9gJD
6xy5F6V/Sx/EP5i6ITo5lhMQFCqJ88joZ2ceZvn8s5CO86VEwqcZhkw2lv0ZtmoY
8ZD7a4VjnJ6RhPzLn/PYmAnre61vBZ71RsiVT025M5i47ob7RvhvfqKJYkk4Lw9z
tBzagHWDSIvciMiwggs3oTCtdxWdSFbLm0SSvhjvnHSGhx3v3W5Cg06glwOhjWqz
zibe0cawzSvkPb2/PzKyox+Qbrf9fe3o838AiRAHgBF0QgTTeC4wkg6I/Y6klw/3
kzMk1F1Kuy3IpVrfDYFkCx3zudYej2Mv+j4wnHpWO3QT0Jgo1QkfIHP4V87RQPjs
tjK3rP4E4nJnSREI6HpxdXp9s1fBBYASPu0z88L6K+aSA5amtj0SjDoozlJ69CCJ
jkq2rlPXxWUotpYFKicVrCW1UFfcUDVJVHvewkBd98xjVlTER3R1Tr3C/BvYIgJA
lEF4GoXCauhpV6xIF/U2fiLwZN+mW14T3GaygsQHfI8UFznjetMU3IkxCM/y3/Gd
ErFO/f2u5fzBTir8+RjK9Tuy5L868qs3bJnoX82Q/uh8SFp73rNIcGSx8LwrJ5hL
b/ZhuOU/WLn4/WdOgSLoQzscKjbfgblSd1wPm6gsZC65fswgolUJNXEzz9SVv3bn
1ggImvPI3QXqUPr7FihoJxPOLLR/FiQ8m9LiDtVCvW20rugtzDDRWDE3C7TEG5aM
D0WBqKjYmeB/PrKPWJATcbk55oHITiIaZkfnj5WX7UdtCPCn5Lgll+JU4C8PYNkS
FYs3XIUj3MpoIprXWl7cPsGsWEpoSXs/+sFfXkWM75B42a02GxSWg/DCkTpMdVG0
HNHry3yiHTYsWJ/EqWSll7tmNRvt7/UulmBz+X7mtHyswC7i/76ZwZMI6yLr0I0g
DWobM/45103879ZgTld3CdwjHJucHuS4/ooqPvBp5+BWc6A6HrSe8DqqU785/tmS
hJIB+citwFq7oJMoFm/FToWLyeLBG4BIBEE51TINyXgGryq3ee0rcecH95jplYAc
79V1pOCOBlSUms5Sn99iZYQTRQ9naTAieBDID5MPVuf08IMr813VNdSTmWa1npic
vtcFX6pTkkThUjLsx8wtQ3zpIhwOTfLaHB996hRUnBxhgN4Sl9MiIluPJJx6kCIS
suFBqxBuLSKvdKDyvGzDzIVS9IWdEPCum4PVTSUTc+v9VqmCCLDUmS59t0xZIkzb
Ddq9zpYfKu19a3NisI48ztKpTYeAOxij0SAJ9eeI6dyZJLPx2HK6obg4/4mOO7vF
53UScpsoB9cmB5XubwqIeQiTbcvbbIgya5ESs9b5Iu/FbtQKI007Nm8H8a12KihC
ph7FojIHJ86o00r89AIsBn6vbpNE7fjke3eP1cAe4pY0RpdsQArYLmafuJZgNs8j
pow40/OczGLnze/CNGEvsAHHx+3p0NRHMCvcZ5sM9xWoQEMrn4NKRlkHEWuko+1s
RW1ZPJmnCCqYS0Rp405PF0E6Kcx8EypBKRlngizogwGFEYlhHmHg5fjRPesdXuUs
NfOwuvSikXkQ3r8LqYBaM97rHEgnKPVByuhqXy5cYx/z9fxEZDTqxEEJ5R1C3nOo
mZ/3UocTDYfY8VweXz5Khsx5Ph68PLz/oulPpaI50q0hjI1Z4kTaA00LtXPW7qY2
04AhisSbiJnfK7kUKA3ClwS52sL+9v4dgWrqvZjSQJBy06x83XzsZTEdhgkwXwb3
HfMUI0syOpfWysmLlQiF0mfJ3Z63kpuzWFuwkPXUkZcbwjd8E3i1ai1aZQQL60FK
MEhTU8erAZbWDl46X6rXEo/P98KQj96yI7UV5Hw/Bn9Rzw5wgCTu81Vf2TVriyqo
Ip8zlso3Dx6gikmju59YASYWgPBgR2vAp2odLGLSIHKXpsZIfz47V2MysMCuNVI+
P4/Ja1FQFgAmK/BwCS1nvP4AcRFBhhYnmKv84Bjws96pHpH0z0sxRenOMXU8rbyo
m5tnnXEJTCe/V6/zJ2ESGtSnQPSivAExkrbbaIjo8Dctuz/E6RHPHx8oTzgCyyXF
PT+IAcPfJs1mr2YLm/vPK/8hfroCOPJSah9S7X9JbG560w6CKp3CYtP3KE0p7Mi3
sxAunwwrSi8QsYi+jV90/vJm2T6eNybC6t+iWIxs/bWTz6sCagEGfMc6wOUpVQGH
ruldEPZsP43TeiDuK0X77RV5Jm2XzgMAUujMVoDe9eC65HS5/FTXWeGdHXnDerPM
VVTM3N8tPPWv3+C6/IlJveXQKKKhHNuE4GWZvgA8RSqZqNAWH1RTziRRPfYmPtTx
HLaPfB6S09V2h9YDzwyJW7QT0BfGC1xNn/14bKujDPlBb9QohyN78kcVvoX08rF0
62o/TqyF5vDgzbbphGjfE0sEypz7fngocLOcyezZamsKyzfGrrpbsN9V0XFw9+K/
DTHZ8CidYni57YKA6AeLOKaDzYvlibsqhQzzUdEMHRmlBGwaa8piJamFlP+Xw5Fh
Xc+8jSBSugyHGP2NpcNfS2AmarZQgIBqH5mhEGbaB5UDHb/uMsrJ2A8HOd6lrWY6
7MxcpqHbfhEn9KhVCupfi0NStv0dwUoQs2/exRV6NEfilaMd8q10+okdQ65avwPU
CI9dy9RaTsmkBRTQNPMm98M+8YPHRztrCNMhfPRSLlGsHNezJRSfxt7kNhDSCOEj
sXPI34lHJk44/KEB3xwUpnXVhpxtyG69UEDvu+J9w7ogF4LzUR/kHpNlPA4XEs8b
VTZRwAaMv+R8LlGsYoYrjCXJz1cDXDxXPY5grrdbxYctqeej9HXTNbsN6f2ojhyX
o0+WEBiQo1fpsgreePL6DqrV0zs0xEXMjlb+ooG34jsSPyknK6/54Zi4/Ch3/Dvt
Syso+JUIHpK4wfcGqqPzZkX5p3rQmGl+DJ1I8cwrsAgLmHO9LyZXd7ILBCJM2UCk
xPZc9j3NjZNeo9GmOZyP1IoMrJFWxR9mn/mFsDuS5xVAPPprx+S9RqUTzHeSE3FV
kJVjQs4paSTobkn/9XMQFrH4jPM72E9BnrGdMZlAuCEJ8S1C8i/jI2MrUSLEys8i
TCZFir8tpNDj1jNrP0BfXFJ6exT/wPzz8Wz+0JQw8E62v/1UA9tTM9uAYf4psH1/
o8kLUupeUCRlmuMVu0QMm+aUePuS7iQLoBDxQkSftXy5gq9oTTQXdLrmnYkPZSLr
CMoqC55PqNa8a2a6shUa4HnKz63K07b2gx0WS2YVjZw/uZU5m7AP8J0BJBmf8JHq
i6Z4dbqwyGCZ30E5RYY+ItsArpi+vQMIFGqOibBWPV/ScohtCn+hht1JjEgetweC
HpFflqfaAVQiQkPetD4VPwwqVykaSKdC7PYYMPSgj8Iw26cXJqhtONUIylgukmKy
KrzgKDY/wBdUEP5m9xgz5t48AYfpXlkDyApqbH2GIGd/QhgqIJBssa/vym4OXqnZ
sUUcVvwoenIvSZZ5Wl+2ICT0oHAgVeQZiL/V4TvNMDczxVrVgoFgT4VFDo7cFsdQ
apjrtT8KQl+1vXybw1A6Ztyd31YYXSKhBjKfHKR1MHr2D3qbppMDoCDG2m/bTqhH
t7yAn58aVgsMAfRxD2Gk1CfmWMK03HxoKLGZsYenEsaSLSEQf9H7ngaSN17Iu5H6
IRI+RbSObv6RFt89wVzLTlHfmBfYidqh5XzK0CzJtnVoYQNJ5aRK7nfQ+EutjH+B
6p6vZ9X3CHzXFgU/KsOcsjdaAweFZARWfyh7yv2xd+cFwNk+FmfP9byrS3IyiFvw
mNfRlqQRVb+yeABpUkEOU/+z3ghQ/B/GfLDASOMWrYk4Bfeq4kIgYH/0Pv7MhVx6
v56s0v64mZ2w76OUPyo0EiIRNUtNLeWgS3VGGxqpEuS+OB57BLoa6Gde2zWXoO8t
oX7fNQtk5RNVwO+ObogBSayr1jiaSFgLSQPMu9IbT7bxcZWvsibfKKSJlQ/qoTlF
LLl7Xebjgxr24MLi6O2M3ATwIIwJc+mn+cmVArGqCvVhy9mS4cPJQ+RwK4fhM+9o
`protect END_PROTECTED
