`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nK8PhyYTh3pLtCCvhIyy5i9nSg0soLssp5tJezGdrGHTLwjNYDpZQT0idh/Edw4w
06iUvs16+jr2wLSIPW/D/yz4Pxvq7SLwXaXH7k/Em4KshYIkz2ldRGd60i1t4K3k
fRDyofR5zCwrwnQcCihYe3AtkrFr+cmbwEc6kxBow6wKkz3i9TnCivPRsh2rSDRb
L6CKGav+qcxRHo+kJlWarY6kvoDY5bbLDe2H4HrlkQlvsXzbjeW5ZbXFWuFRJZyx
hWByhzGFYQilFwc/lfIF/miBBL/sh0bULtHDudhJ/cn0Dmhd4C4By8dI3/UjzXFr
9IfaZkJLWfPk7YjvacOvao+l+K0DHTkLhViQdUFtjFOUyqZec/uFL5xhJ6t70kwR
PEdiQ53ea4x5VarSBs2y57GMblYZhGu64bmiVZNMU468eTpIkat1e3eW/YGPmIqL
8/W2QDN85HuHNcLYe8u/fnFVtLXzRkTRF/KT2UqglVjMjluC6A9ma4+Tpv+7b14t
OUH+NBTsvM8scQnEcdb9LIwYttjDK+ExgffeWCHTtKzBf53zV8oSKPqMdVAwX5zp
jCvVuKfVGWKAyTIrAVbAM5WzN9/qUIyflbkqrDeGjeuyPVIQTDiy7swhxc7wQs5j
gsLjHljM1xUMv678y0sdfC7j8aIL/uaBHafyUey8DVS80SsYDNQ8fotoGtF/GZ3C
KuCRz57jipkCJ7iiqzvLL77NspOCxN56InXtAS2muMskkVelXX/we4pea8HogLHP
nH8yDO6oJLHTeGMR2rk1jOlVyeGYIOtxWfhzMJ/aBCWPXJjsc5HaGkU9ugMsDxE0
5pNBgm5ySyuUlYhhPJdOWcpHZPKAVVmbMsQVmfBnJsN7xVX8pU9Bi6WNqPGDfj0C
RQVmtzmvmHEoQc8/JCNT3EZ+SxTcHEgUII04C5PRbp4M60/p/wX8OjpPTe9gW+T0
ooDKJapSTO6tdFLtL3ZjhM3KKr0EirJZiDDrsTjcNMP0/Yg1kmkclrfNGHISx+Tp
2km+harI93X0iTLofLoto2C28JS/Xj+hndUUMOKko8+8mTU71MJ7D1vNkwMTLW+/
530H6bYlhoaN7K91mgkfqKqse4CDm+2m3gLadxhI3ay3cuc2WAS7+7yrjsygn7N6
ZlnWB3wCX5shchN1NICnDdWIR9dEFaPaJBAhZYO3RvNFpSU668ypaHd/OuIzZhK5
n2gAxE4TJ0CpQdMhV+hNY0u5a+PPUfuPfKlb8He+ajWFjEzDdwJuRlICsvuW+qIv
yqdx2xIgbOEEk29iE4n2EQUr036xYO4g+RelFmFS0nAGV0hQcZXRlczkzddrdYsA
TcaNGaBU3C+3TAyled9egilqBm+ipHDmlDgNHF/AVHnFX9gHmNhcmd73ax+CcxgN
hJGmsLN2YUmZj0KT4d+hDgoc9sLoYZftBENb8XMIxFQKM7ASRYzG8BmNLyifwoXR
bYeJysLyH1cbUg3rkQgjC1iqo9nxm4hlw58kcPodSmDaLjaR5w31YN4uJ91Gn/9X
9Uw/8Hby2Tf7rl4n+oCjPfq23GBbyUp3+fMhA308XPjICvamHdr97zHm7EYT+nIT
8et7nbGS0ICzgKqMb4ZDHQ==
`protect END_PROTECTED
