`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PV5csyfOwfhj3YvR1TUSgGer8wp4SxL+/NTHgepAFvPM7TZFMIqms8ku3UFxgCJW
8Ck/Tb4w65d6SAtYGvbJvJVKobwtLFH6ueVWADoxZY1aqvmHocj429zEWqcRDqHV
eeokLp83T2ScLnvvs7d8Z7nlRDZRUHa+cQW5MY6jMwujHfL0hlN6C4qG+PiyA3wr
jxrmlgYe+TC3vkMZaZZYNZJFwy/O9+lw5bbCjzPRSid6WdDCDJyPhhrcuJybHGN9
yILjELhdGxLUEDYgsia/sIur/0rKfhW8dC6ebo1h3cov35JLAx/JEAIR1HpoDL19
wVG0opUAHi1YckcKnPLsxxH/ds+GrxQ6IAEz516nmQ5+E7UqI6+U9R8zvDTdqbsz
/592/VYTGqey3K2F/G5qZA==
`protect END_PROTECTED
