`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qQIThGtbRkK6Kor2rKevS8ESy35ZAsrwsflmFo5f44suYTEHqQcahipoWknCYP67
4wULzLAA5dA+WNrxpb8igFO5OfjUfx4DM4X+5+NGgzI3zyN1TALpM2nk6+MwZfal
92oJPJ2ggu5My0gjeZNwHTnHE9S1dRpVtIZfAwHwQ9kY15/HGliQex4ASsbgkTCT
moniarm9tePQ9je3Op6Upd+CHiM0E7hSP+HFzM3C0f0cl1unkEQLsXt25V1zOlbh
Aq6m3RIW8p8RQ/Y+bNfYHIxLyg/8ns6tXTGooiVCuFVaWOtPzO9PUFHB0hv4sOUc
Az37IqSm3ip6ocyV4/QLOdsT21EQYGCvknS3qfZhgoroDey/ZBpfFsF4SM2cMtSy
IDIjYdR82EnO1juG3ETBslUVgVMqgWJO8+YO93eJKOV3d2+LVWJaCKwdUujMGCbl
hsTT1M5YZnv1I/glQeBkvyIyDqmFGnJ7josvXOjKKyWJ63SxaWWMF6CnzAmKyij9
fkcUSmrWakQmu97RMiXPBJ/Jkc9SQPrzQ57Mk7Uvt0cyn6dpGq2/ru9AAuB+At4c
NA1WUCLPfRWe5VR0vuwc6w==
`protect END_PROTECTED
