`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
teb9Jc8iZqTPiC4PG0pCJeEGK6nHlUE0Cc4vLZCageD02kMtif42B8F+hWMwqjA8
1lNQ6urGX5IaasMHMFf5sXAF9HwndztPHDwJ8EKy3cB8T2fvfLQwlHLdAXUyTsa0
UnNhdvXqNb5t2yzuV/JLARSWdm77lomx96qpdKbA70i6S6oXgkB/R/Mht5aajCMH
Qpah1r0lSPceVmHTARO74d1z8VbdvzL8L8vo9pftk463C8pOZLjC04AENvtZFRka
Xugz7twEwxPefM8TMIrrXAGoC6AVK65wocOTKB17QdQaS9INELm1tW5dyvo7lK+W
p3n1mtreZFtNjr8hovAeadV0lNMz4WYAJFD2L7wHH3IVkNy5vZzmDTli2glXprki
It4nEvqOB6sRsEOvNaufUGYD/OOdtATBY0JG4a/5P0zMm/vf0xjzcb9ESC+gVlBg
`protect END_PROTECTED
