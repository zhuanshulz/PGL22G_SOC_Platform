`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCJ86nwzi33uIX279quOqr+BZrZpiXpPQ6jRa0BkhJdhJXou/1ugk314hxz5r58E
usR9FktcgmlOC6T1bNOxBuBkgo3vQbffomoZ7GGtJXstAk1JElsPCgknwkPC8ePM
MdghTT1nx9cGJeSGrrNCinLEb4PalIPTGDcejBO5Fc7RRtYcinVxUDbbkk/mNn9b
i6Mh0ryjTRV8469L5n7X6XtTnrhLKJtU7bMrOnBheT2QDMtt25AUySVyP7F61FuA
SZ4JWH/Kuiz9qLBVKGqh8OBS3UdCnrxXiEjVJbp1Cl2FKNW/oowB+nvOFhZZ5Z09
P0oUKdEEJmiNwv+DrW4FQyq21TywSC8eoXb4mZFW3XgZR8a5NNQRE5VSJ4+i8F0r
x4WhNu3Pfa+s5RAjLE9Bz/ZNMG3noRkgJAAy1eY1oQ85I5RrmO0G8Evn8INdlStV
3BcClXrrMsMM4neIcYkdjPcl+Qsxv8SF1kZLLMSgcSuHoH1b1LLzvSx6quw7QHkG
0x6J2KxCHt4c2o4ba+0/OSErYjRyBSUU8c9TLAYPvCEnKwwglLRsS3lF8dtKCOIq
dixSIWtOnF5XrVbW/yEbaYmNlyN8GSe7Aj5Meo313Ew5lwQIPKVLrOkMJPmrY1jr
9tF6eDSD18pGxQUJpJ/mA4MfibwK/qO36F0gBkKksWZ1i/Fzn1UTkIyUVfn6o/C9
4XAGIhwZpqrN4NPtOPBLZ/NtC1CIx/eZv7fuJ5R3No8KVQWxy3IzmZGrec6ftXFi
eQQ/9i6K5rYlLKyF1pDOv7mDCIxCx2pRr3EpQA0D7QGFaEQI1or96ZiUETRUG7xs
wz+7sEtwBJ/fHcmWm2caLonQKkubkpUkgSK4UdZtqyi1Yb9+LFiDXy9SY0cST2K7
8mmE9B7k8EvuRvIGTQodXKx5FYSHcMzBtJDFaj/8U564CUrZxxuxTrEQBVGWKQle
F6uhnSfamklWlpJfSPH0VuDQCn9Z6Xa83W2HZvUe55sL2WaoDelr5+zAmIU/sSxj
kIF3zcMM5PaUyS5mCUIPP0dSvdemM/o50lcNmdyz/1I/kgTe0uNd1z0GQ11nOssd
Htu4RB+ll77kecpJ2jYUod6ivyxcM/gZ/uUsnTloRZyTYe4scEbPqph18zyKrRwv
QbxeGf+1LjpuTLjBJW9qD9CFQvNePgjXRvtc9nVFiWNewYCwFOq5HkUtEV4tn+32
x8Rn9SBgPtIUlEXoKCxxaERiAvCMOZ3MplOhtNQuUxnLfjhkcqu4CBQefFz8i+qq
9cYS3ymAULDsoyZcBshTrQXw1b4Qa+OiMwKJnLzq/5c+75Fx6s7Pqt/Xuk9cMRhT
d+wv66E8lEA4gI5S65ma0Y7r7Q4YBhyYaCUym4KG/midg6/j0C3Yqu8ENRWZvMg3
YAs15swizB3NaXtYYpZXYUbAJB35Xwh25dx02tTqJPKkdhHSmXe4uVcUQPrklkqF
hxuKYuCZ8ZxKJZR/wD1MZFCg+gRn93f3EsEIELY3UmvYRAdUJ+hLcUOkF1eE5qWg
M+0f9Pec3bneeiB4mVfT/53mbJpDrYRT4PXbbGqzhLMvLJqbirXloyKA7f3yikIr
BOtfwZRK9WpbKbK21IWpD3364dCYsHFubHKfubB/ck2YleGl0kMF6ia7M4amoYni
aBxxlJCmMmW+cYAkF5iodD4OjEqYRge1yD5TPb046v/7WFSZgTHAwWB7gFSYhhb8
3XIcWpNOXVJa8xNsnv9HRJWND5hGbp5sA2yqoP/wnskqgAJIDGQJI5KOGI67NC6m
z2vU5dni7jg1Bsew06KdL7H3AWqy/AJhuKscRXFVp9NLuAakoB9dBycF6sFwayq9
BVQxin9TPtNxnqWRAJH3WmzkrgxRKx7AJ1dG/ILyFAuti8LBDe2LvwcaIu+aYfcw
oy5JvPh7U2CNLubw0h8i9tpFM99V1tl+Lj1gzHlla3H2Pz/B/0m93FYvP9Ce7Z0c
dTdTlZCbBBK3Hzvd8eplpFUhvW/e1diB8m70GzjhkkRS88Xwy2G5ewpJPwIVA9dd
yNIvPR7X/kSE7TCbFBS8HxcyPwcRwIlP9UFzVmsy2cFvyj7C72NU6l4hi9jD5YWj
PVlZLo5naGbHnfkKphxBBvQf4oHFh+Tahe9sO8Vlq6+nPAgPZJXBJUXtkNEiIEdH
nHUCD99YJAkiqCsPEDnTcow86sSKHbilBG1ASHXRNe6/UFLFQcbsHgA1F6BN2BYh
hFcigvWJ7FDn3cjhlbzQPAKKe4kK3FkRAoh643uZgacxHLHNPPXguBZrhZqhmk24
jXzcqIf+Is/cqbq3BhK5I/xwOabR7JtACCBQZmoavmk1YQt8Kyi1ywp+Gz5zU3LB
SlUBGKHUdUdl+df2U0Q+wYF5Q5+D0vXj/za/4RDYQYIYfa24nVywEkQC/XxvXYnb
9obWwQifGdRntjENYkyHw0RBgujx7ymgSxxtIAy7SPiEYgoj2t1vJXnt/GsjV2AX
NdSJiRJj7Peva5mQQugoXwuh5Y9a6CmlX7OH8ydC0A+kINxFskCnGPzAcYLft5AY
6Pa6NpgJBZxt0YfmYBxoMO/0wrTbvejPp82okI28AQUX0YdgB3x9zYscnTLwxmzf
WF8ggNTYwbyU0nfUGD/zKMVsEG/E8Cu7GDkMS8a6x0QTmbMo0YAE7D10fZ+Fqw0j
zhwxi3xxujQJZX/+6zN3vRHywb4KdvNtC/7RbXb6Pt3yP0cE4psyemGtIi9UY/Uh
h0hIoLIdEt07++QdeXfjNCMJOPE7M53N/CDC/Y5y/xsN1kg/la9FGljd+6oASZ7J
fy+oMM3U6A6cFXH3ZPLO2DV/QBn4OhApjls5GOaJu2lJpaNm4yv9sOCMYrTPWiwc
lKGScpXa01rb7N9gB3T61Z4ixNU+jwAnoyCDWwXsRGrO6JYOErx5Phw9ZKoRaM9H
XQRsCBaUQOLVwl/4XSkUo9HTpFlo5bbQ2haMFh9a5ydUeYgOCoSd/dyRFpPOK4Hh
gbEfQ9YP2+iPCm7OzMBcFhY4C9LWy+gifE/s99f/14EriTNTlgMaaco19s7/oCth
OBEQSlbMEmoVBwjuDJAAi1GZYCota0ailq7g9FJu1/xTpjG9EtOLWFiw+Ogyc0oH
nsdpQeQ7itIggcKgYw+1lRD/CfVM2JWC1AF99LubRLzgVkzgU/InUpSU16/eQLFL
+qDO3FKSk+q8fWK6cMEU88q8g0pX6d+b5+IJ70op2aJ/4etCgErjOrgoQGvkIH4d
Ncr0ySrp4kgB/GJ9chi754ICIcybSR1UGNIXdk2dT2FHApnv6nPa7s6WxxR5jmJ8
AJgGUZbE3w9U2Lfqb5bn7dqjJ66CN6JHF8vpIpzz+UKMgRQDoGvb3nhuQlTRToAc
sJ+ucZaNoqhisYnfXuFRr22EzbVRC9QQNmdQwKCbF6uabttq3lyQtNdFHbTVXLO+
YNP7M0TO3BBVbkPQh7q/XJILDpY6FaMftbLrqnp8j6whAd2TsWHwt8uXL7tLFGcG
Pbz6+U3LnuVrmuz08um6a+PqdAzS5PFBKF16Y4Bkg/a96b8kvzuxxfm+Z7cFHjeN
3QVvLT+z72Ks3ufyd7LhGwuZhiJAfJwx6fYXe+fqLVyHkj3ds7VhJmgANepdt7dx
fN5mqTlo48PAdIuwCLuifU9Xqh3Nv6hfhts2XvywC8FVRaLHwAIIkdHzYXrcveeC
ntbee/GAuJiIg4a91y89sEgVY8w5pdyk2GHc36bYAUw7G/2kKMqY+93WTqAzVBNM
VLwDh297A09zF+F5qSq3v9b5S2M+Dn6DmfWY+7lf98EElcksVz+ND8nVbyI/b13Q
nk217A0iSfuTfUyD5e22gY3b9XaN3uy5g666OsgdhHtaKQCtRu7fpUIbwINaxYjM
kEPbZ5yQ+mkJ4xf1SkcGhCgcz64BingHpCM0+7b2IVqZd7HauCOiapUHjv8DZvoI
FaqZwwJ/U/bQSU6ColR9N3eL9bwue2SJTfy8twY5UI1i56w+UCT8uhUTn4cpC36j
PhY8sS2Y7T4Mmy32hrHathK/l+NtljAlJi7eQgX62/DMK/nk+RGuaK190PowTYlV
6c8CG8EaOOeife+AA38lNYaMlu5d1LczCg3Cg0Kz8zRK9QXLyvogyWZ0KCk1Y3os
OM1ylzlK8E7IdpQReFWotbEsZMNNjFfUyNs6wnPRo+j7Si+uZ1Ua3LvrlcLjKLBR
HJ8GKLeemwEBCTgFe7WwNGO1S4xd5WbjrrA0FdZwpE3zeviJVjOsyV+NvmjWLE88
SUU6Ewz1BLaYmN2AF3A4vXb5ruskAlpMJOfAT8fbVyk6gBH5EvyST/Mc2JqYR5+S
xOIwYz5f1U+t0fgBg5uWSva+Lht4EM0qARJc838PkN7VJfVG/MRGXuWYnnDJgSYz
bat/JYGAPv4KjjdMpy3AAC35O+sXZZCv4L/rtR3wZ799PODL5UFXzB2c5ch/pshP
4R5MXtyIGXaG5h/fDJqE8I1MOJ6e07iF3OfiRksd6k8gBg8PslZeK2uCwW6j7Kii
VqHeYFnH+gW/nV836mc9pqEIq44Dea+gclH5pho0jCmGObqmkIOzJj9wtEac3AT3
hqGf6+SVxB5/Aj+ZIO98PkCuvJBELxdhOLHaSTq7mI1ZDf2OWybc3I3IWPHoZyr+
kuYJnXLWfhwVu7Y7p+Yhxj46FwdEKJJ1re6fCe0smIM2HmrpS93Krb5yqynUO+Sj
9FcSBu//v04LqLRrGNk/f1+fSSz/SUtP/hvoXL4DQEP8wj9hgdSf79BWXHBPftxy
4sji1pHM7aj2W4Vq8MvAVtqI5/EjZpAX2EPqZxziIAAzMNOEyWv9H7sTNJfx9xEC
yOl+2n2Fr6X0pX2eA/D4uky96BZ7uR+x081DeK0TBteKgTUZRt7nbtDksp6qERZt
VZxwU1ThWDHZ8KDVxKoan3NAQq16i+QulOjbM4jygX2oEW2u1rPvH/Q2CESTRhyy
nRgDvC3b8ezASOqW2YEQwCP4gWS/QKJEfuHxK+WnVKwZV37aIZkRtcdff2r6csuT
+VNdgyWFu28QyW+st+Q7eKaxIXtuEgzXcLqHXD3RYNQkZHUw/7ZF6FGgZ1JbrgbI
PHRm43UXmHml2IqNQbF5DmSjKdmGRAQMCuQ4q8ep8BcMfPCuSQ54e8hIaNc/oZzR
SOw9WB81qOloCadRTR/L8ZyokEagradGVzHAqIiOj2MwUzuSDBf3Vw7O0rmygsEV
HslAE1w+46iyrqjOEmRNOZZYr6LsPcfk/+kaLNGpNB30OnXambePpJWFbD6cFUb+
DtTaMfIw/l4yKKOQ+Fmg1zWSiJziPQFUBajnda2KTxHyzI9wC7X6ZFhGPaKvHE2E
EkkVxRxL2KVw9K7jsZsEFs9AlPsspxA7EH8jr+J0lbS6e82ihzsPjx0vilA21OE5
n/TNiVCDoqMFKLhsGdHUHdQOPjmwxRfUNcSObg9IMK3+1R1G0p0l3yN3seIw3dWf
g3Hml/U7hrxcpDfDC1Yz9C+9IwInUxNBlaH5sgp87FtzpCSi28m5SDP75/d4NNhM
XRIBTXDmdHv7wlqixb+//NItLBBSTuRF868enuF38Ta3xW8iZR1C0Alc6rD3dFkA
sd8fxS1sqB6XUljeJu0PASMy3w5oz9qzG7yQss7/JF7DCynW81kGeFC6gLCQP9lt
g13MrDzqM9x1qVH+EKRsNJ9OGDvBcN9ark+o/6q+J9Ty37UaWO8qydSswfG1RXia
MO/gXcKNY03CQ1TdomuK5MDefL706lFxSXiJ/vk1KRVRO3mptOB0mbZXx1GJCG7Y
srAdb1k87pJIKW/J6dtv0VIyIz0yO9woWsfhZNT4KlJID61Q60DE6QCVQ7zMxhjS
M6W4lQ6HgEzdxJzoWN9VctTlWvS2tQjnupvmOV8O3qhpQI7/MH3M7DKWiXfqktu+
YNmbhH49bYM80u1Zo7xrVJ1Lv91OTWaP5B17RoK3mg920BzhBSZjCtLYDc8PcWl+
EMf7Lu1aBC6HBsb+loCAwkUE2dyqkz75XaW/ylGvzih7fFoVjqXlIxsMjYQOSLMS
hJWwiFUQyQmkgUcsZWbn0NfeTEeDmIWsuRuFRMgiSxWRgYmP5D6aflW3D2vBhaWx
S68HiHeLzzYvnqSzcVuDIX73KlOofA/JpfnW5noEFHeX0f8mVd/V4LDlS7J2BmRp
hMUImdotGhAwjwZgv/oKA4yU3PW0QH7Nx+nHyuD8IXCrQOPCY9uSVu8WeycEB5e0
vd6jqUpDJmf5wBaLxSUefJTav4XI5/D3YT33lHKzQ9rFrd24LFZ0uvgNIjFaRzzz
JjFt+PfFfcQS0pPpoE0adjuVC3XddlH+5a9iOZ9VAXQYwyQpJtBi2K9z8b4RbH4L
zqVmDSJCtxxF/+8n68ubfAlpX6AZSRJBRZyG4eUlZBmkvrjX7i5LKIpJKtVAEkSW
0jx8BHgB2tg4/tvl4/jByuv3y0R8XlfKlJWFmyX+g0ZOGM4lPMSxwX8cU/eF/kD1
zFgUsaYDgrxffgJORZDfUyDyDl/LGxsEIh2RJwnkz5oH1F6/B2s1yHr+IkZXzha4
HdJ96pqjvvxsx66h0lzAKFjW5jURLssFi9w6VyE2fT52l23GFqKjSNJKj0jLC92e
2utzL0dAzUEo5SuSSVPWhsIKPulljeWGrvZcKPsDQMAUNQ8UsZ/JgCPWZz6nhIRh
WtEuTIHPG7cAx2ro1PhRsYvIG1qhkKtivk+1jnu7wUfsXK3Fd/4i4jFx4vju4KDa
U5D0FcXEpSL0ycwjgC9GCHidCYtkmTXJusKsy740IM2rEDdvo0BAQSGR0KKsFsuC
ItaXjMysm1hMuAy1CK+2LMgurTYhjMjoZ6cf2KP1omrkg93Ns00OA1AzB4C4In9y
gbJpGb9qwnLM9fC6ZqxW6JPpnDZhgi3gjbdRjkbH+0ztRRx4319GdmQL4W+4MLnA
9dQH9u4ICZJasCVBPTfpNjyu1S0o/nJkzikUm39yhQ0=
`protect END_PROTECTED
