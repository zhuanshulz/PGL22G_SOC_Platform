`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6z1KgsCtgnzry5lbxnfwj93psm9cz8qKRPXNll4t73So60hID9M1T1uOUWaV0Zs8
Zgo/vBkIyM4CGJAKUNBoocIm6HVc5jnQaXofLEJoP1qPXavEdu6FHnWD3xuE6M5b
SzMBRJLcbGfdQtrMSCYQ8eabQRsGd3KWuPpZKFUJBWdLO1AU3ZSLH6OIvDCHK1YD
KigVdF4j2KLA+eD6k3E74G1AxOYtCnvIqLKd/FE23MycM6cwL/t380eo4h6Y4RAt
tA60y5U1wViZnfnGiv/9SxpfNZpBo0kDey7iiRjc4y4DHnJTLg8zkhKLVSnZddVo
AMSoiTl3fl5wZd1Eg+VtMyvMyBpdsRLTumU0/FYFkCoPpn2YRP+Y2Ph/UzaW4WfO
55adsoCURwmIWKNCZm/U6awyCgS/4kY9CXd+92XnIxuq+lX+k6cqgaa3NUm0tf2H
VSdF5RMPdo8UturfKEvboeRwGjoMetkrAIvYisF9tGx248zNVjEBdd2MHB8xMvaq
O6Hm4eeuAO3FpVxWOuOJJeDxKMvY/Sgt2OIYjAxOg6//Se8erj89NMx5+zBrY+Qw
yxUwTV3p6Bxrlqf7wBjlSvO34kzAJmuKxA41hoLOD9Q8H5F3k47o8XTY17AxSbar
WCRWjYjQB6jfbX9ylhoP965sE2BulxlNxz2BJs1lNqaO4hW13AW9PN/W04v3R9Tt
en5fxNKErdsNKTvAfXk+A2xWJYjx8qm4OfYza8rfmUQiuYK+NPnegeQKBv2cpidA
i7/voT8fuWo/bnYzQq/ZG+XfN4gk9UdJXxrQHWv/l+ROnLLPTJFnlWI/soh1UOSg
uEFNItk8fyFmb23RIaFHlPedH1xkxX/b0Cv4aUYj5Ph/qcAkfPc07o0HaAbIPa5W
C6DGqtRrsZTvLMSaCITAoRaZ2nGBxVW4oJ2/Q8BHfYKG8oO1AaIi3kbyBTQs2du5
hMJlBf6xSThJTJnJtoUN32OcruzzeCOznWs+CG+K3FzOo7ogiW0eMJPATqvRhsXw
aTSgqItXoT2Ik1JDWr+ZIWCZo7GOxirJ3qXQBF1VkWLPSl1vJHnzT61foBr4GriI
88KteIS2BRjCwe+T+tvpeD/hZGMnX7LtjQhF+17GUj3WnpeyjMhLm9WaQDKE7Kgg
AQp+42137a7qGYWqr07XY7uJianaQWDavBQdjRnTnUoiaGQSHpR5tTLXIAjSJcAI
SFyWxWtq1hGQiBCDOkIGNyfCvxvgkkGWB6F39Beaic4yXygqGB+/djOCXoKY5/+2
oK8Pj0DY9URfLC491hpnbY49i/UuSqpZpGQMjHOyT92QJQUwDgCMdKnegkMJOmOG
CodVwjbOP2REKGchEy+p4ogMqjbSGoDCBRiC3O1ArDqiynei43p3fh3jhGkuvB04
mLISkMJUwcX1Tuxe2QxCYoQBZJfHGtdoa1M5xx1wRHeCdBqGFCOvhLdoJJydUc/O
m3zkj3lgfr51sm7yfTO6e8V1ADTOmAnJPdkQ2CFgsfqS60XEU2H+XxOGxwb6Qih+
BNwLJzilZrBZQw7q5CkNLx68H3wHHD+6m/EaEte6HhyyFIaKSLYc2gIYVDOZF8Ne
jljb/JMXDZWNCwtUrERRBxjDM+QNbDki8/TMxsFXYQi9/LIKEFZljZEIB7qcfYNj
5aTTy+qyhK6b8IWAMOOu0VJ+2hhkP5HIeRhbpVI5Byz4O2gCKliCQu6PVeCAXzQX
Xu3O/jCWb7/DsfFpjxlDbugANsSqG5sfniysbZJoSdF7qi1sz3j4ShmeOJxKccZV
fIppWR1zyDfe5x2SElzQO1flj4UC/7D1D9TpcNeTy/A2+9M0hrCeFNvD81bmepIt
qefDhJnkKdHuB1IKJc2e4XCd4OH7MZkFmTbbqYb6R+r7kBzlz/M+fpHcV2DBlbUw
f1OF/T0RVz8IYZBcEFY+QocHQWSZw6sT4Dc9z30LWZzKkDthY9ptwoSWkcPv3lWU
Sj9N1tGTp2svZx8IFHBqr73U+4+Z6KdlqEHJtaJmZvM7i9JhbS7O06KqYPMSNMl7
IYt3AAbsAN7dMJs2UL+GQ5IcqBdkQd36Rj2oXBKBsRkfNv59yHqety5rNXdOyOUK
GP9lVzbc9QbAe4pb7dilVoB9H5i+9azWURvvALLmUJkmzkLAtlyfWxTcXkAEe/5t
SSU9a9OVD677zin6yWSetdYEryZ9coJr1Jc14S7OAAIz27p/h6oAS6HrwqeBlf2g
zJepteY6I5+XfZtalVQzQwg1qWuJAgex3woxCHFemwokck6ULvHrMak+nmVOuMHK
yTdWjtNLtRTrIcgkj0hfsGOYT7nc065H2Oj/myf8uqe4fyreUS1a7D476kY3/YU0
mpT16LokGTF+z961wvWx7M+LhdUjhZjhkPSMdDWBR+VJINdNBfRX95pQ3NqRr7rj
ZYc5ufYkb0NM0mmPYcldXM4gtflCgl47oX/gBRna1mDw1Snd23g8XZ4y7idI2zE4
ORFFaHy//bfe9SQXKF2LQBqbTTDwM2pdLjaOu2fB+E1EStrEw6qRBvyuxmwvEqJh
YgPAVZvVMo6tBvi9Ntu9fBF6be+0+Y/xcJw6AQ1ROlC9Eyx7VSkEFgZ8fGLbeqLs
Iq8lGSkrw/90bCTonWYauAQRSDHkQXLKvIroy6IwoQXAREPmjpGIjMT4N0JZ6xVl
gSznNhfSrLeq7HBWI2sUgB6C+amAGL/u2P4bv+rhcTB/P9OmDCdTpxsl1f7ZtnN3
Scy25fYRkyUtVj8b+X0WbzxCC5c7Ak8X3uW/5QJjFfwlwL4gXrzGwI1YX1YHoVVv
klsrqjWdUErokehHAbU+g/6SpaCSIF8djzbI4dbjBXbp5HQRQCNW90VR/SG1DRGT
0p9r/wz5Jm8OyhfHqARZiG5sDoaEncAI/g0vca52HSBIURmw5lBRhQ7MfnEXPmmm
d9iJAxpZO0e/Fp3lMu04m/WVa4eWTgSkiXeoPyGBlzrBv5p/3ogBTD+6bHFtU9Nm
C0neqXzVN9z4GGG4M1w14yUbIGdfqPXI41t0KcH+CDVheDekNHnLROgneFFQpKhi
CQMonA7m/wA7fXGkqqSYDR5XrKSlNiWJ6IzbBXA+9dDdRIMum42w+YcCe2o2xOqI
TQwSzfCFHN93LO2GgZnBJRVG1rGRGXZEmTaT9Z1jdDQnOhTpD/GoddOEmHh3YrNm
9LbtZVEUnrPSBZ9axBMWBL8t/WIwcqW9EQLCty6rfwCE6u+WDvFv/YuPZ6+c8e/q
3FFJidfR/iu88hMqpK5SwbOnNYbRcYKpDtaGUy6hz43AzAk+QpT4Fjk7kCSG5GCv
IXx+PJBci/RhSRRRRa2ajpmP3w4Y5ZxZswjXmWbEHGEVxt9C3mqbld8q0N07Jp8L
JCojZlRzyqMPVsY7Pbnic7GEhNuc84eP/+JslNNceCOAZQ/bCoun7CadpyCCPqZX
kpX708dNNy2gjNHLyt0ygK7xjGbKz+UtZ3ZT5ZbQEinVOlrvpwAT8QjAqt35YGWO
EwKIHNDvbARuL77cRTHDPpQ3aUcpOAq7u4F2SO+GpXx+XLYpaXaOowBxl6KSR8yz
Z7Mpx7CSCiiZhFnzTs4W/yH0HVio7BfqC0u8Jow1Z+ToNkxjEdKvLmgeuVVuJHDh
SjPccISRgqayPFY3I4x0Qb+hDGGRt++uJdJ3Y8yDcOp/to5aWF5RZ2C1eA9Utjq/
25uqjY5c4dxcEp9x+QYV5sotsJrT+pEb24CiddkZIE1pZxeL10cAXqlUmVy6njy7
Jl6LzWbWku3kmqJveZcm85pfHV5KhELVTJ4Dg2bETUcEtO6gJjB96MNYpVUjpB7S
Qvzo2ZMtOISG9HvfzMaVyPewVVWQPVDW85cdyfVO7GsFcFAoNAKOKc5FOCbmI7gm
p71w4N7uj4KSwIk1TSBvUhOcMGQSFbWrIHPtsyGoIwu9JgbD904tVoAAcJZpysuI
8D8B5BJPjRPlfgepWdzv4GfFlpf8JdDclB+5NJY0XuR17s6Q0PHOBsqFyN35QRu/
J5smKv8n7K2VBFfPajzgjqhgeiYqAfoJ07wydGeWyMSXfpkbN8QBc7ZurM3ppbkb
iSy49fTuPXv4CPHW5pcpGKK7EDz/z0uqZO6wKgNi5hTVK0Ue6d1wJAjPCzGbpQpd
CLOAy5ASOBjNckWZdYHZftLncpz8Xl+SdLkidPP2PDRMQIjmF+sq1fvGHl8W/M6K
KK7FAtHv4lpqMGGR4ipk421D1651358ttzMqaowob3Y1dT1xf8bRkkS1k0ceKHpy
G1Uwz4tXpJ0/zBrk9bQd6FYLOmMRaer6nwjr8Z4k35O8n72+dCjhoejziKpgosmu
Ln9Sn1XPbgnydT1suAEqNTykmJ/wtqNoe5HAUnPEwubeSjwBK2j8Q69x+CUdYLKH
7Q+cyYeFe01vkyQFD43UP+1Za+K1eF39Dni+Wya98mFxje8/JC3/Ps+T2bUG7PVX
V5BAy/X3gHImSomTfdRtbdzoVzTU70leWx/woWwhbjgQ3SBw5hutaz9upwpGNVhp
iXToUV76YpKBvswi3fdwX4i9w8DUOZAmeDXHGQEuz4OY7ZNlX1YsRsVM6cFPPYGQ
jqVYSg2D/0KJ3YHVlA4AfFS6+39MHe0KwXWYpmhmpPDzYz03DsvbC/6uqL6ZjDtv
Nw8dGXOLTutwXy4TeRzBhYXVJMi6vMM591juFYtGcKDvh0awx9iGVc3O/JirII21
hFr1fpg5Ivi6Cq2vOK6Lrgqh1sOnbXEOx7zBF+aykefWm4YcuZz23l9hHmb9uk6c
eUYwtLv3UE4/7bQfynQ0BSegL8z7rpj/NLvT/vf/uEL3hNAJg/oI7xMvCOXEa69G
euyDgHeVIj+hUzDy/15VyToTyaYhyOtwtFpdfBx0g08JA7KI0nBCe0eXMI5DXf1Y
KjLhMQtb1SB9B53hmXmZZjPsdJ5Fqf2lSW2B+oFAucc2Ask8q6tlZEPEgFWpFeie
7289r2pM8K1c8QaujzbRtfV3I0pa6vg6PPONhYGWp5buptIdIuWYYv6w+pWQWo3U
IEuFs0sWEIl2vBN0gcQVBnayN5Ehv5nvrHJfQxBpYIbmHUp5xNovMAW28LDIPBld
0uDrV0S05NPTHWwRPsECi7hlEGaeSaeC6SKM/hmaVEXdWyEeFjqILVo0s/b1/9rF
Lt/WTkY3G+BC48KbUUeTgYYYKymYfdN6VaVM0VBaNyOY2VBdtkl9pWlBc8UcssPY
dahttDHFdrowB+Ht2XyfYCFwgEaP4de4bpct976TDcd4cjw2ZXSaylDtrF3JVZct
5B4hZcU851VZecVH7M+3IzbLakG/RYAYJhs2CqZJYoQOxxATH1DoO22fwIvHWEXi
heOBiBp29wLLRJlsJEELIFg4BWZfFFhwBZh7QoBWhx5dkwcgIn2fGCIvP9zYcW1T
1FjQWhWMjnup/pkbj6cZ6g0hokq+cGznN2MDh9SZ4EQZsN7bbkvAPZ4H5jzl9lIh
5S2WXUpLlWNDxdU3vU+Q9W7IWVx8R4FRG6SUqKMMHCsMJ//nO0coH9TGLDwfT+D2
JxYwFKpJzgh9PGbFqMXC7a1Axcjq/jYyrKpMlrpGD7BX7jM0ROqMG0tQxxqW9mc7
tDhyYFdZrCg/7Y2x0+Hhgx+qlBRZCzbER+eXLZvKA0PoLWUfOXxss54yUcW4J85z
pjZtqdShCRt14CMWySiDddrLHAkN2pqnXtvOlNcWNX+fVaF7zJZB37AtRCplCl+r
NZtrK/RfyPGu+/UlbmaVFdKhZ/QzUdzgA4gT2E8TCSOAF1c5VnUDaMojclmNhsi7
xKA644bdJ7U+weQIQSmqD4Np1uANHxtZkI+aWHbB6Y9K+tP/UKUFQyaWr1o2Lz7o
7WH5o7vOa5B7eCNt+NeLw5XKRklIae4YLeJDpM3f/nV8knBLJFxPQDWXBDxGSy1e
yUxkaCNcwtIr6iKL1ocUYLTIqVf4epi9+cWG4wRkQ+mthKx3PxfGEakSztdwPja4
j9CBMzwtTkjFlmToUXKmq6+wiPoHLNynCO7D3jhLtRCdu3PRY20motQpocGZ+4/w
jqS8Dp79H9ZVtnAL+ZFdXkbLeqAIZg6uWaXa3F04SuUiqJs57EZSOvslosnGTzQH
dtnMZDNzzWgO+c5xqHLzeMuU8VzAd8JapXPIM3o9CRz69FJp33cUvmitbxo81jCA
zplG6hkz4S3jrBjdKMeXABbwI3DY/FGqPX5tRD+h7x4egxF5T4nDZTaIhMjvqopK
HEfpAqQSQaEUyIgF46dHgBHzQ6fgt79aTEzINK/TWnfGohseteiImRsnV2Njc2pS
Hd6OaQNpKkF3EGNNFTCALo6B3MzQN7/mE30yRSwSPhcw3WsrWjFqG5/LXUFYU5X1
AB5sCOtmCTnkcK+ocT6xBp9YC+l7a3qcbHA3xoO2cODpZnL219pl4CT8TT9FOIsP
V7wUA2TOl+cH9qzVt61etC3s7BKevqCyDS/0efghCBzhCxaDcvTDHReiYY/zo+QG
MU7+83M/MJl1V4czHLj/dSoYw0WQjmWVZco3RUPLD3h8q0tjo+FzDMB9kljz2MB6
GZVpOOCy6x90aSTbCFbUlHIZhwvWdIJMS+MV1YEprF0SnHpDmxWmYomceluYuHO7
21SScJAosbVW6SDtewIEWW4Q27y5hWeJo6LEXEjsvOR8YMBkjNIEPYXQbZRs3WuK
IKWlf9NKmRuHBD3pWxkG7UiXede6LMtj8Xa9FZ7XBmwXRZ/GK/JNA9XDBhlef/0i
kG7JrbuWWxA60Q0PYtRwI1axmkWJjYR0QG2PSvum4RX0c4jZtflm4qYYjl3IOQZN
UGO7wa1C6Fqrx8p4oK+5Yn/r4zw04cENVMxeYp1fbHkZyARdK4N0Mg/y4f2PjpA7
wiQoIg9BLN/j4N1mL4tCvXtouVgLkvxLtKxHFTBz0/UHYaRhvRyFwMU+1SS4aft7
oI3JghwQxHIoPihdy3K2Rz4vctpMJxGEPslDQ4kPFyRUD+PLdQamWd0OGQpaZ++B
YOgwm36aBd2prItWgpdTS8j9LPjiJ7n1i/GY5E9JNPwV6NB7gKdePs8ia8cknWFy
qhHlusJVmgvGoWR59kSfjSDvS83nUQxG27EO5Uuy2ZPJwtdvwBZ/8PEPZkSReOLI
GxZvoN2tM2LqbOqJMSWg/Y9ATAYsY/DvaEWyt2uTk2wdJ3nuEbNuPf7dtRHTelAq
cPupPBnlYkt3lWZIDyZ87PrA0tU4Cs8Quyqw7r0HgTPCVDYBWZD5Z87yiO9u3cvt
/8Oja3W/1jxXThOUd5uax5xapRMZoRteOgta+kgHAxGRrKM9Ik3ar+yeCoc5L6am
wcVwj9Wqfo+CsBPecPHVF4kbvDf5U8x4bTkF9jh/c2LK2n2zvBVwb12Gk50zKRoT
FWcbGtmPiYe3DR/rWxie37pqBewZjYNE8S/G8iZHAoL66sEgE6ZxnkxTWCdwBsbu
VCzsHMVDprfPvRUMoQW9Avqs4Ifq3FMLOc0YK32WDl9yf/XxKEJw1DslyE11DrxN
OEd5I6V6U+z6c4lwqXOyFhe0wsr2LbOH6WaHseZmFxBcYHcQwzwSSe/qkLaxOTXB
ivo7fxG5k1pI9wSeKO43AgjbPIz4a1fK0Unnm/KIzQiBtXJACLEMTd94KHHGCAmS
lP8SOt03sGxQBAZw6wZnmRrtMUb5cpxnLO+YutSPUJuVKFrEgGVt2thpdZrEJlSp
Xt5SuAhSdJqunz48p7RkK1NMIty3obp+TqxNYGRR9g6LcBH4GdgFtwanDHcUvgjn
eEpNdU4/N2GO1McE2l3q5kDZdBb1lRaQsD/69IqOrdD7N02eMasEfknlo2ZHDHXa
HZan8u9hylDto8wg4oKqG/649aJQjqBxiCCDGljOM/BVY9futtqAzbRN1mu5GtNx
mYOq+0jTeftAF4Pyua5udXKvIm+8SSwjzVFGKDKaCELk7JDpgqNLzhemasElGWoO
bn/sEcHNlnXdIwVhKpqPKD6bKQfZc88qD5J/9Z+IpUOvjrvWIjz6QmUMHz51BojF
wM14l8G8SjtQRhdf4squdFIg+0/NKkDkLJhv3xednIq8+K4Uq733V6fHdvatlK0U
fM/MmVsJRz0NCwTcJDSutUVmz1T0dYEUC8MBl7iZmIo6K/WIydfUL8qRVdxmjw5t
3RZiP972sxoYBKg2WTQhTJDjRo8itUpWLeksMBz85daCXDPX8uHbpVdq4n18My3K
i/tMCzktWdB5QfJiba6MrGCE6XXbDaA5khdEK40mbucE9Aj3mStLqytYLOI6pT6r
t2TGMccRXw0ybuHHJF08gLb+4OxEPzxXpJ0kEW8nfuSmxsAYkgkNEQ1drQkbP5++
B5msMRuUi92fAmaP7rOEc0hMrkPHzrGKKnTxh95tsYEu+rlrBr5vEj5O6fU57Usc
sf0HiloBv26bZ6Y8ySlQ3hKOBBz4FrfaAudOgoehq7Uqb6YAkGdf0Y+hRUb2b9D6
kWydZ3LzkwGMsZHUqu1D61FMjdBuVAB0PEoSqAcJwCPyqGfXTmdGIjMRWVpKHf/t
stbSe/RXXg4iuox44TaMFy+fih7Zs6+yN03qzBSXjuc0LTQxnhbGij9EApuH1iX2
OCQ6/qh/Z1kcOBdzwT0mTZUjbZD7DzUTstxRypxuK4CGFb4gg7DbbuMEB6Ph6/iF
qg8O/9IT08MvWg5fV1dVMCzjVMZ6sqdaAS19FMt5FAAngUIQxldYlZOx/OWZqoyB
a0v6wCKaPJSdlnwWjBkAWPf5G57hsg/xbUjG6dkLmklqvexqI5P8AvVaAQ7w+Y42
zLfvwH5WDG8FWQm8tZIkUeuE6+zTvMYTNOVB28EGvpLt66fEPWeYMe6v4Tm2V0/7
qeCFv27bA4HAGin/TbaalJIXamiOirkxVv6GqWwwq7LMDXwqMRAX8UYzVr9rs6XT
zZkC1T+3ELnmfPV68OJjuJb+BQ//D42cDOM4owuVMEby1Nycz+2YvFTkGdPdjNeC
kHI06D+4uBmeBcNXU0/t5jlaySAmx+4LWVCv9QmMbnTpzepk+P3KR1BvRcOSKfkl
Gpmv05ew6cF/BWt+QSUD/IhYHom3PLS84Qknx0Mx3NlBqb9qQZEnd8R3PnuMWZZR
HGTnr2jLzuy3NdivJWUQ3hfPxJWPLKFNhsPGSvTCBLYnUeTh71I7qxDr3tsM63Mp
k9azj4jmOXkqVcs00tA2luF2L8ugTshIaR5OeNQqqla29qmhd9oGawfs2cPEqCtI
M29mdKdRXIzfefVGmEVGOFmQzod85cq/oIjh9LOt4o7xQQtdX/bCCdutMaOSCM47
Aqtv8gEFbHIp0tw2Vg5egvMhItqFs5BLQS8Wp9lhh9ao3XxpEe5Cj39F/tQaXh25
Ls+DZO4OiT5TAu6xEw7WbX/4koWgJ7DfcXMCZJrsxV86R1ADxGEoTWjGdWliFvGo
YjEz8dahbVGYZ7HKIoTO6cXDxpdUbnSVVZxweAQpZNe1zdaG9KicVKMV1fG5R45Q
MnYMVrH0DA+NFdLEkpTEY6R/uQ4YDaYovQcPrn1HotjjjPjo0oS9HMQLCHYr0H8U
8lIxhUqtIporqvJkuWOXlynM2nzpt1pbXDko5wYcd96R89XoM6udb7rIWfb0W31e
GORznAfCElApxYJI8zu8TFiJw/CtskjegjEgMkiRVigwkCuC2d+ONLxYkF8XR6tD
ooSmXhhVTKM+3UlAPOFnVKAtx9/oUR6Jnr/lnSzleIVT0FPgcHSZ9EkQqP0pQ0tJ
Jk0SpM64FTm2/YAiAfbMobE4XCmTPiaL3bNisV0byr9wnVBO41oxKntdufRv3cJE
l5udWMOQiTu63sEu3E8ZA9VQFZFI/ad+K8KGRMnDvyHBXin3YSbhNgeiVV9f5noZ
EEoZ+oh27VEbJSV/BQJgkL3Y+VFtkgosAyghivHaOXueLW8kMo1XvxIyL7Jzmn4R
XlW8Xh11vtfcsZbSbVQ3pXQ45+9G3S8e3BefaoRetCVyL6cgExdcCZDkCsKFBlCH
Zhgfo7XIkKWcdpQzRuQuzcgeXve1/mIRjDaK9+cq97py5e63F0v+45DwB7ewA1uT
Kw+e/+kBbRqL8VlimNvlUeGFb/FF88hXQV3wjLHoJqOUiTH8zwxfQV1TopibXpQV
WB2WgXJT4KLyAtsVoCMo3yEZHTVhFHjTV+Oq7NAbZvTcat8BzKMv7CkxIEpKRFwq
bIwBKovWiY2ALI00QN7zcTZpEg3VBQtETGarAo8xVrR2CVpDYn+u9QTquI9LwIhG
/Qo7Vz3tq3PJBHnHAcPNZeqTQPzb5izNEhjePKp43kb1IXktCacjl3mBYg2e7Nr3
QozGdyBF4QbkZDNrBRovuYBhV37P/0qo+2wSLOS4wgafhUx9LVXPud+jpP0bfJSU
J6THYTJ1BpCtr5i2eTOiqt5PYoKIOzk0YJUFdicMB8RF8KuXlutZYqFJoSOTaBu9
cfo5FIh/0vbVNtjdUDNI2VMJE8bvC+7fztvtlslD1ak0SW/UUQIT+pIkHoFmUGVP
HEiDsBVrtzYv9kkkt8jCBSMjdQkygqSo8e1qpyR00S+jBMzVf36LRyse1S31PU8L
D8EfCqr7ZmXv9UQl0Yjuh84rHwOkGbxdJ8X+niuqt0JMo4W3OCdma2xFflBLS3xb
/yFZot0ED+/RMpfuYPOpbyDr2FOVC4QpgC1dXr2qkDbiYPv0YjOPWiXNL8wIzqcR
/Vj4TfKGumIkeolfkp/2rp0cEtkpmtqXtU2QaU52b0CZmf33q+ZSC/w2qPSn5g2v
F7h5AuJSYBSiMxnGgVNlqgxUNBwis0gfnJT0eNfOQW1eHuvgnf6v2G+FT06USAHw
jshn+VWSowAC4u+Nr51B0XIFXa1LzFMw2D8ngv7VRk1IpOSQLXCaQH2/DbGANn7c
l6zd6TD2mQIebM5DDKwkO4LHhy3MDgGkjrL0IPRqzwDPfgMs45CoF++kmcezhfPz
iADwJ95SZEwAot3cscWmyXvKy3t2QndF6JBdnme3LMEO1oI/oXcdcDFq90iOAoTw
MbcixmkjFzJez7Egrxcw2rdXQIPNh88pvb4337xLVfpiiR4J+fz8oJBjJ7r0eaOy
Odgjrf1dEgDcC8uQ1cWQv7p0UVT9qyIrBkpX3lYgUcWZMdyinLf07gMYLLUOpvmq
IsFxBpHtltXZ7Vd+JYN8Uu7sM/z2jv6FZGfXOjgNtyaqT92p+ztLdpJECd/tQGIH
Dq/IBliBMl8xiD5uPlsXgXAUwBTTMFW9M7F/8zn6SKf6gaP2jP2qT+d8VOz/BRZF
a/GbAJONve2zzwDrsR/zUh0pAgYe9tHt5sAEu9YLnUMYEA42bMsmtla3AMiieBPV
7xE8WCTpuLQ/CbtsiIwy7XQKD0hssxIzuSQtHXS+9+oLSySoexF4r0uKtokRQWLm
upHgLV7BIq2m4NkfyBiEmowUjQVYp3nTj+Pv3wOZ5igAkwJxyjhxW3Xt2FNNhu4h
aLb1TGELeww9RpM5MCqwApO3F9yRWZLs/uKpAu0C68AwRFAw11JLk2+JieGYo4Cs
amNT0nAAvCzz3z51Nw09lIyLo2cOFvtaBYWH0dKWMlqdYHHNtjvcwFwEbAXGzgvf
FkoQEitzeajhXprrPt8JU2ax006/dAasupYxskLPiesmwjdHYGhTz6h4UMglUPS8
a9AqbjOenYzOHRrGeEwfusXEtxtuXMgeGkAGrmRFlJng5+AeAYKr5+9pfQHt/GBb
A2jsABIpIwov0SXQ3jeHkWGdRFgDA04QYEZGUA1NjVGsYCyT+GJ8bbgpP3mohsy3
pRAVFceDm70UQF/s+zRqhpX7R0UrH7aUjUkGFm4+ewLbPnRS8v+wsktqoPKPthD9
W7+aQVKr5XNHAwn+N5doVIio60GB3htl1cpLQ70JeHbGkanIW+Ph7weMMTKHT4pG
xxx4SWBS2mVFC7GNCrp9ssM2KzHKbk7yOZ9nIA2DDVXKijEO5nIanCHiTOTyeYH2
CehZ8iU2bHNeWH76wQ0ESb1GTc71yejk58x/KHz2aJg9aAqDwk33E8l/Dv4KjPc6
re0UM/9JkOgCfDwapVxgAoE66erZ/sVWABXvLInIDLq+k9ta2jQljXXZsdlyX109
reNQ1eZddefw+mkNe1cnKUA7SJozstDPEz2B0xzZI8Fp05UJ3oyR/pjbkd2oYezn
zXd791dH656BX/Dfg6zLDcCUdWKRbYMSkzbVFAMGSoaEEMKAvvi1zQHFhNnBJ/Jc
npbXRXalA+e4nfULFVTXE6psfGZHDuwVxqDcryo4CiYAjo0eHr+4TxXRWjdn8O0j
gQDDYBFofWZqgZQa8RjScfXTN8D7CAmEy0/gifrwiQ5yvqEV+1OSVB3NGTY7obg4
/sTWn9U0yvSEIHSBVPRsu5oNN6W29CvyU5Y0mKMAMPTay9El+p+Q7QOSiucbEZhv
NCxylo1p/VBwf8dDXTI1oj1/vfPslNe7CEUQ4pnTXrs6wi776Sxfl3O4AUmC2ldf
AVrZuxci5/l3X3QeSN2cLxSLJH8EXRGYy4yoqTpcbVFroQliNC9TMUCLNOvtIQj5
+kNvIpDN34pUn8qlwswQThjuzdqq8iON3y323jTt+yLIgs+ccqeihPkdmPK7Ey6e
2meEPfJfoaSR0+gGserEMsUjLJQeMBuvtNh3yxkVd4Bv7VKVZQdfr/nLVee1uU6B
9M3YIxKITsmbS/9D1Eco5f75gKZUHuSsqcjsz4iK91tyDTYiQGcK2R741H1baiSr
NmLsaAoeoKL/ZxYeUDfk4E+0f2NEaWx878rbMAexznfNKc8n7vKhzgLQqjnzWNc4
0TP/WePT/cgVPYsUsUOgnSGhztUOBZAfl5P3qB01Ro+bROccLj8mfhD4RBLLcdB8
K/kqi/aPP84u/RYhRFz7mtx5X0vO34FavJNNr3GURVEeTXD5pS0R1McGeZstUNJb
nmyGBiQcI7kclExBOiAf71D1t8iC1AkrfWekDE6sYhT14kos4z9zFiSKdUXVo4fK
BLDD6hUUOm9LTrMPvxkTOpLTJTvEv7+hz7oIaLBPaiWb2cOqSDZm543kcqgsNvwu
hpDP3Rh/KLjYByMFYRZepYxnVfyxDnPggrMeNui44Nb16W/runYnymhfmD7RfnYP
NcVodmyLWokLKg8bw2XAhCrItSMtCUObYdELoEIIXvqJ/nD9O8G1FcRXo6tjWwdM
4Qe9cQwg7CYG5tlt5S7SNXq80R695vUm3+xX9YtjEOBeG9ApH+OWQy1nlhFRRa8+
kyGOYuoebSHh7TU/oTTTZSmIFacrIBINWpPpkkXW5QmWc0+dTxCV8/KRSkke0uQu
cFisBlPLXdZk00ZvXrlXx1LUJTfdgoA99rUuLG5EpliwSOfQHWgEf1Xp0GIjn3mD
ZQxOIpcy2tgjmrxOXX6Xloy3bMFpLYeUoXP1G2rxhaegZPgBxeM+sWN3a2DujvKi
D64I2dBj+yd2IX/R4kRVNxZ3BS+PnKrsIw0xDW7ykV3NKsHRosRSpylUeFiET49e
s4Zhrhiw36tMYbjaodyWT/Ddose0Ej+r1b2uX7zJHmzxdMquQOst8c1gF4H0aUud
/gkTPSSPSvQB1DI3TZ8gMzcBWIx605CTQKI2Zr6FM5RlZW6lgvThXZT8bfj+wBw3
G/boYeY4pmTzL60xaV1LKApUlR81V1cJjyDvSy9RRM0fMNDU1F2kaWdIQRXxewZk
MH0BEIJm5y/kXG1SiU/uTKhSRv+g55OR9iSbLwEwQrPKv01hzsmJgPS+CCahZj/j
IMK7zhRJzPd476oN8AqrH22Pq9VzmKyyFW/wZtK1iIQ1kDY0OgHqX1qQlHvEAgbI
PsJi1nEDR+SZC53EJS6h0UnxNf4sc4xPq3FG6la1tyNdZAAF9rMve3+oxT84FGTk
ejG7j3qTacZ6/Z4vXzDvEQhbfag5OHpjp+ZkVJ5ELU8CcYqLXPBADmrOwiJvGTP8
r2ebtZ7OPvYgfEJT/wgkoGg1czTg3bBosyCrssAPYbbxcBaY5aT2TqK4BFQcNlSs
ZWxQzM0IMKZfVxJkLRGCTAVMMrkHnS4SU1igZuDAiKKfMWDsPVcSQygM3hckncNQ
1DNHzN/KYnVu2YUZVWb5+z7ZrAKtXZqye2+H+HNm24KduAFjog6GGv3j1b2o6jra
UKmtqaq17qBDy7XPLv9/P1ejLokPrcls8zwexep8fVcpVJaEZCjnvtVABWEJQnmM
FIn2kNxELD/LJtDEQ1YK6vV9yd4Nl/nZChPZcb9z9khT1b/yTEt065/MMXssXOmx
5k7ZlPYiw7U1r0XQQ59zGp75rjowwPjJkARJfku/qbExjJWFM7ZysmNbHUnIxBMn
omx1biz+lfGEIveAARBYsGsz9EpmoXuVT43Sqqi69BGNvXrDgsZTg7zjYV6+h6gx
8uDfPrvoFwKrzZOS5ykVe14DLAgSlrPd75jZqc0a6h9Pe+kImX6nOW+W0DXSY/py
iIp1Rxo4X3cAvFqKfNoBRHgL/4RxhIbJ5sX4+udJBRKSI60NHlSNwgiuq30NJ/oW
zlEisH/sVTF5nwtEPSInsTCnNVHDHPKW8RcqaM5jlsrJ8CTxM/XSFE+TZHEidXtG
4qH+4i5rrkjjDOH1rPOgB/xvfJA3x3vWUdMPd5E/Pk74w0e2GNK6BvTCkjT/mhBb
1MCfdGE3rg6PIsxDa3W+B25FmAOvZSWKqUgJk+ovlf2PqvGQnGKDwdcr6akLsp1L
c4wamiNKWiC57YyYeudvKkUa75koqo4o4AEcA5PNftckuYA7MUmk2HVgxLVAfBrL
1ObkKI+zUgb7Gc0iyUg/W5bPV2Ys+KA3MtU6Ih96tj/6JQaUtK8fUSkocPN1m7hb
k5LaLrZgzImuK8bBYvsGqLMLu7AjctNug14hADj7TcXcxAaaObR+6mSI97dwOFOH
aa60UUaF5JE/xlFk01yDSBYTL18NcEwhp9lqDCAiR3HTLotTRLH4fWoO+uCjnfR0
56XUWBl7b/d5lBNP3lDiLHW2CTIJQ5BuLhwwXnNcuAf0xy2lFaNGiw/zq2QaflpQ
MG+3ur8/b9SzuMIHnFcONFZ/hSNA+g34rl3N86X9soC0UKvJ33NdelfbB7zUspFP
NmYXdS7xbiLFJCVJ5jKqMwCl4WZBZzb1BmkIPSUJmZnVI1fYDJ8KYEoQVvqI8pkk
A3mnQGoQkpxUgYmVHGSOAmfxMaPN9KFzmx0FT4NS3XSjc+D9MsFigl2n4IiDthZ7
Z2L8ip62qFRA78nVA6mOQT+3w6vilyu9xEt1GlCpP0XbqGELc/24//m1LzDefzQN
eEbMkRS8MjBrDv6kFhtt3IZVyseWPC+UFa7lgBOtyBIcz33NNo8e4B5Q4kRptBHa
prtPwfXfiB3qS0fiR4qTT1CWmHe8H7Ntu3L57XIGfZpGsmbZRzIiouD7cxqIR0sj
P1ZqZ54sXfOYKEy1YZFCxvNQBgV9HK95quWIijmZXphg19h10R/lNn4mV2GvsTUm
93vZ2zMrFumi3TCDLNUP8zb11G0yyi4Oai3D84uk8/BM83hgn5kE5yvBms49Lv/H
LhntWcfcKMUNksgZkU4/WyCgZaFbo57+aIM/qh5S3ejzUBc01H+0gTu3KSIjYLuR
pXLO/xxqZs6u6Jq+jONAd1Leyw8A8YC+8Uh4smD9VgONTrXzE7M4lKKQeCXnfTII
LrOuqpF0TAizum+wtZnric4ykLWQOsbg+X10nfTHjUrq7WTKUh17jDHpz9xHpIWB
cppXpWYYHbxIqDUIUNAnM9RSFQZZ/QMb3Gt7TeL6TzI+islVSYr7rpexzCyFI+AJ
fcI7kMT7y8lDj/Av+mVI/J2TOjYOzoIFcCl/vSzsknj+F1qAxUjDNMRx9OJaIwWv
jE3skv6uVlhiVuFAAxVukRyNz1/GKn7BlEIrLaf9rTEDyXPiRQT9wXEWoRjGEkZ2
NvZR2ZpDsahix/jdevrU/O5CNSCdxXoPMecUxU+4DJKqryEoEX7Y6H60vonFfffM
+BiPkbYC0e72QPi2n+LwZnGGXoNJXW24vG0tj2HQ00MhKgilMCJ27Ij//3Q00SEY
FQbPOmIprwgGcj5i2wRhiJA9mHzZwMUsFI0wOYLDOV1c2bzkq7P+eXpIMLrhHtPZ
IaaP1JRF7h5z2oNhId+AUyj02cXMiI+cEyZn6n1zGgcAQ29lJeTSqAtC6H6JBUSy
LnEsM2VB03QMhMjpeytbaRKq6P+euAMaNpF+JU4cFNT/F+AJt7a0b0wlnLdpAAsu
BB164w+Vbv9dOsjMFrNOWh2t0Vg3HqpZ3IMl1IyMMluguJo7mLPfoHJOufbnXIiR
3+f0JX1at5f5mbzlk8Uglz3JsWaac2PwzBqUR2hleeWitJscSWVMcixPl0kgRbQe
97DwBIAMU6tMdotB8iZ2cwd9tlyPGI9iCqnmuN7vGrCVeWhH8bEHycia/Qeo9BgD
D6BlDQeyuGed0IpfUpOK3yVvlewkdah5DG+5MpGFj/l3NNn1dQmGR9Adc49eyYBU
/1aN+IfjQy0bDwp1ln5D/qQmGizV6xXhuEqBnmAipivQyqvMNniaCXbjF7FiUCFc
BQ9t6en18D9czAPSfqoNw9PE5h0iNV05xy51ZzYjm+sp/kpWgzDbIoEitk+W6L+v
cl/sevo5b05ne7b3SIC90YDv4Z5NJKrZgrZRd5Xj5+L06XS0P2n28sQznyWvCHOn
P+8Gg5+2GWoWf6J31ZAzCKu2ZaR2ijcMSQtJu/u/x/2c3dtYDb7SZ7zdaXx7Fc8R
R7NTALIEy0qgQy2Wj3qaTQiN2z6XEZd3r1weBGLstSQ98edIJi9kjXEA3K1PL/rI
npKuG7Z+P/d+DQ2U+qhfXf9wv+D0BakzMkuSoree1HUYEYPY8hIYpi3YKN6tPxOC
Mj4XDv1qWu+GeqpdUZ3YSmhFjteWh5V4jzb7wM63/VbAlinrRF+0pjzAXNHnRwhR
v2Z3FcOCY9Y8cUwKlZaP5ITzrvkL+sHG9nL61tyYnPEo1unX8VdjhQDAjyzLzs/V
ylwQ+FngAZ8hK58UyGSl9QSe+CZt4DhQPlAkHqzxBRuyiIUnQTk5dEeRODeyy2nk
PE64Igiz+RmoKnkFH3S80v0AIDDK4GQSu1QdclHpThRTly8h8bilWB8QhErdw9LH
N7QwUiSWlmYwTWTYlSnLNZ+jMk8s6l8tJeJQdZwdCKF2WzXeMqKFJ5nKBzP1mxOA
kKgwuMRamBhhU3St6FP/IG2EBo+V9Ak/b8YLplNOwt/Mb3xKnliNrlyQvGgzrsLV
jmq7c8vQICCpwOP0nk+V9Z5S29iz6JuomPvguafNRObO4ZIPCrnFzhjiQ2AEhjua
Y7LHDZmi9FAhtefZMjs62/rnmAXaXUBISEtLBK9bqmbzE5Qq6tGp7ycDSOTKSdDN
08RUKLfkq025bTkKWjtfiHvzNav8n/1eU86haG1L4XmX0+sDRRnl2Y8sG1kmEH5j
eiixSTy4jDjRLTUkIA/RHfiwGPZqojawnGoNgrP3Xe7mLJxAFYxhWZzJ0B+LJ5fr
dloQGSyaGyEdtj+J1EQjL5lcNLJywPj2WiQ9JeXqIWfXR+rResA1qOdVPZiw0ZTH
SLfeqgmJ0k11KbXZpqvwXUZQYpCJ/6C4A0BPeGi6NYy5F102AG+RSUbAuW5i6Hmg
0uzMdd0zpAzNzVKuLSFZ23c7W7dqabOXL/J8EIwL0oxpTMq4SasViPN62eBtCye/
/pzFucsVJrJfqIdHs8RaMiZPaU/ZkJZPAFKsuz+YIsbHdhvXg6TXTM5YgGEM96wE
pAMpDhho10X8l34F70Kp1nP3Rt1vuOcZyat7IENDNj4yQ+TFnxdueTdqDipj/SGs
Twbc2PZP7EZENpvfs9fhbOWlVH0bX5a6jSseuR0Ey3zE/EYNmrbR+/gc2W+I1jDA
j57G/vA4Ml5NntN14UjlwGX6S9QVBIbrgL++ezlrcMcTRmsXqNHlwGS4nBM3UKSP
n5pKEgbGHTxMYygErUZjr1DLVNsBAhafH1HffEeqIbSCm/ik49c4sZMy8RsCcrWe
Zvwf9VU9TW0rOwkl3lcvRjvIIBVrzCDHeJOsWuzWJMQzfRFzhZpGl+bkwfJbemZq
49kpFFP90Ilkozbtu4b9L1qMZUVIO8qp2zdZtMS2/tSkVn3B8wec75e7zmWlXFMc
Ho3XwbI/44he1cs2O3xLtaULP4qdYNt3Budl+F2SNXCSC8IyH8kjILgXNcuCmJ31
6CH/mg6GfF3RBcBBbfZvIz7IqwkKMqvsEnczXLVIIOhMgYPG6/I7SWpTUuMRUASQ
aYlpCOXcHRWQ3hAxiOYWDNNuMyouMZ+T3K5t9EJMBvwCf2Y+5qORR5fjjtomoxqj
HxflgTjOvm1lfBHxKpnWgEUmuC3+7MITWwlRol1PVjuX/76fwoQMAPJTyyoej1bG
S3uN3bo//edhnunNEO3P+yyoHCvBchPEpEyHcOQ39rmqujzg1lKcnxu9I21iNzd2
Ca4FLJGXK7QK0Pe7mMlatr5aaVTu4LMuBcguOqqfKqxbmit4kBVkFJreIlVtbVRL
gYMZtrPKIqDs3884zQJytwkGdpLGH1NjqNTS/BRiKCX07NJXUe4/sIE9U1a4+M/D
t8L/ZfI95jD+6FbHPvtUzXkBwp2yGoS+uPyMZgssVETrg5SxD0EmtGsJWfXJfaZp
+mRBgF+uPrJrGKf9/RkANJ4bVAsURzB4g9jvqvg/Xpts0Sr1Ua9yV43freprlfIh
0+UlCzzieeVp8ObI3GTpkfC+jlbOD9XngflCrTAStqnLrRn92izVA9XDafCWMXGF
HIJlL7Ql9MbXR/J8ZKB5psjJJk6mO4xT9NRTUQr2zjbTgTHDwL83UKE/wGRU6iMM
3wcnqMNA0Mx0PkMs5Qc2jxBOnYSLihf7F9nGnh+IKl2jfFOF7+xEVF0HsYeELgA9
voihzy//UzHyFKPejC23L65QwrUuVsGY9tllmq8UL8U3d0X91mhXEaXCkF8GRudB
Ui8gw813mwi4RqL/1iu+lpOQlg5w+qpk5opLCT32O5BWJxtOcehn+6NaKvnQBS9u
8LkhKuTBRjPHucruqrfxUze0vK+nkKwKcrTQ1RwM/5qChWBlazfe/1PgkSuKAVvg
f4ZmTT1CynmiVzg60Ww7R/jST8Tz3KAGEiLxHlbeG91GLS+k1ePRW+6FDAIBfSHj
3JjRL1udapFNe45DzJ7hd/uPcVlnmflyKUfnP8YK8x96hl2CBcWGhrEs8nRLbfrS
fKUw8V3GHiCoVzwvxKumsqMO7kuUHnlqXONoPfD6LZEMd5UUrdHvf8X6lvUXqTLx
yueC7fm470xA6FtzvMsfFzEhoRWFK3h6XhjUIY+RrMVw6u+tBa5U8oTSY8Oh9/r6
KsOChM2MfSMXQ8uI8mz3oS1Vnk31xA1EJ6YG71F06IgwVY50UyY39XYp4TjqTxaJ
oNbPXD3u8uFwc3IH3rhHZ2ACE+F1A0mxdPnwSbJ0zno7FalkvH2ZEN29ZOwYb2hC
5NKRBGeweTh0xXSTTB/u75wud15nLIfh+zsiavS0lxYGvBkjY3XHgENEwPfr0ycp
4xTkU3QtKx2j35bdMDSqxlp6jPTx5V7dPUxO3/V/DS6ohw5q4COCMHq6AdINuH+M
aDWipf1eu4MiDQP0LPkyRuQi2q2CL3aRSQve2L35d0Ul7et36bYXpiiIk/MkOlkq
IM74xR5JeWBf6QK6YZpl5XX7PavwYnnNK/87krxAl2lVs8OeEQiPcp3jy+sO4Z1i
eYFUKrwEZfT6a+Sl4xnwhR7XZdjWP/TTF1VzlxHwuzNram5RQdVnYZX8rgqahNyb
dcYlGDXVVPlO23LfszzDSsgF+G2lKsNAb/yBmpkX6S5kdLtymJk0UkDOF5ikjqWL
OxES+Y6nra97pUReH7yTf0yi7GBc6zgz321lZDRFgsQZ5AThVCatX5CqbzPFGs0f
5iS1k/5iSqCHO4xbHHlagcyBnP1YtRiaz50MvTRkqgbd7kwHHwLAlEbSv0o6ag7i
JtEUgOipyBBW6imt17V645Rp3DP78aQjja8r+aIRRLWx3nthxb9eJ2FKPQcHvWX5
fxJnOwLKDzwmE+1wgRbTL2lacxrCslVsVfe+LbkNMExHEDSE7F6Mw4eahlz9HAzX
WXSXoVMg+alhpkLD4plhpeEmN2TmgbkTtZmfHQ6ya4qtvSNgWn+oNo5czv3mtBwS
GLZGSLrXoZ1LDulSg7InUGEq1rBcAjUF6NstF9Jn5pfVILsF89+bBY7azUjYba3+
SMMUUFbsR+9Y/mGvee2l5lvBJDT9lC/8exWaxlDcJ4l65OYNNWpe1f+H9WrWCcWe
kDZgo8m2cVZxEq82Hl5d//5QC8VkrDg0Pz9VWkX3ITrOGF3fK5AB0Lidqo3P/kSy
obepyRYR6io4VRHCIwXQ7ICA3lgW9fAhr6wZ5jlSqdMsyDpsh+JyiX/K67BwoAE0
QTY05zk1mW5n6Lt8uD4Y1pvFkOE/5qCGzKrPdiEkjvo=
`protect END_PROTECTED
