`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xL3H/P4jzozyQ6jjdlNz7nl4MMWak7kp4VJWaF45zS44jSIeqO+UHrPn+HjcChB5
09AExblAPB9Mljo8AtzVcfftbKtNi5G41ldSZnjCdZvKzl3TXFl+x2UwySQbSnIg
6FkbwnOsDt6p7kJKA2Wek4VCNRSkkd5UN+59YaJMHUm4AZuZ9PuEvjdY7lU98b5t
RimK153yrurduw/3ljQKbwbmdQuhE8wSzdKU2Diaz/FtPne5nvvwsomrSqNsZ41E
WIwNYq1E25rLamqSSLKNDVhEgj8x2C7l/r+ba/oUkila1qvdXSbQS89XJ2vi9GQu
uxHVg2FIVvvmz7qKlzHT1cHgv/kJNVOoFZCy0BqdCiht0C0ErJJVkAnzB3selREt
CRis5BZU3AARDRLtNxKDFHm7ARuViI8Oe66elAzuLjDeN8yhyERKiQDJV4FjbSJM
TEX/kxlZmaeiDyu8/idI03nDmXppUMX1w/z8412SmJswiBfDVqj3RTUlMw8IXkyv
lsMezS9zZP7xsiSSPTu5/sfhWSvYD0PMFTLkfXP0RwmA4bFJMmbVBLlv2ACVmWi5
UtR0DuXPYkeU0W+OiMtlLQ==
`protect END_PROTECTED
