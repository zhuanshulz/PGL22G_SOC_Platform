`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ypViotNR1Bk0JVrmC9sbh7zz2KVsxXJNkGNRdzt6Nz4jNy15iZtFatKgKmVGfiX
3m6fP98pCudNWttJy0Bwpw1ephWgtE7z5gkUZcgoiwJFEIHRGSDgH1ArnF/YZ2LB
O/EDECTDMSty5MjX5Vpwj/u8/lO2UR14FxQkvS/9mbDUuP+JwtF859bCCFr9YKai
rep9VzgOOe1I1PquvdMbTR77Emc3JpL0s7twqqSpedL/ahUKVEtkqGl12EiI3AFz
sMtEJTgETwwJ5IkulZH1u+dvGKrMbT7Q01shx2T5jTVnj3KLEIsDblW6hRflObYX
WWuuhMlDRvegRQqfaq4sII55j+m4nfqyv06eYWG2YYY/9IzGgZu2C5vMGVKGQnhM
3jApxF0bEEmD+QEuC6B8q0YWGxznMCwAzw7XJfCcQ1++OvXnuls2QVnDhqqcaZlA
yJ/7oNT92GkKXFN0R41d9W1kv7VGw5wkfOWN9nCoMnWcben6lXxORjBZ7Frdwt+j
hrGEdM0IMDtXFoPhW4hSpgGqrHBAfoADxNrPAYbXcui1klQJOBc61hvgkPDZj7Gt
ibWR4K0a2gLEI01JjMubzvs/6c0QCoMO27YRXcr2t01puZKq35uYD7hc8KFj8Kn3
GCJRWQ9UOv4HPZ/RwQCVSMBoZC9Jgrf2oARXpmLcUYCoMaGswUOV4Xj7mWSelrTZ
EBXTIym3LvDkpJp9VNqzDcWCPNDeyLJOU03SUFJ71kTAfimemhMPMAs2SgW5aBjB
PO6LljgYoSCGRusMs95hqay4qJoGgCdtnV1oIJuvwqpbCNeTlXrBkDRfoyzNDNXE
/K4rPVdpQcsIwRlAhpmjWetnaP8XIbThaZZxsC72VQxwdUH2Wj98aF8L8jdjjZvL
Ovtvnytsic5gc21DhH+uD1g9O74FY832EHA3+tqOyw/rwDYJWDyCqR4jgtU9wtml
1Dx7myL8fUdH0eRK4axYoXCHyLPqm3xwonj/0+iUOUhtmQ798EfHMiC5mQbquQHP
dRIQp7OYaWR1LKUG6ohfDn2nGLWEP6DB9HSb3VALDYlFzpZHMDT4UqEQxmQK9rZO
7K5obQaiuGZRaIYsmklL0IR7Q/WxmcgdcagS911nOBc8o6NWroYwHvTpZ6dBA+Vl
o+rZXJcsKY3D9A9Ja1jLhzFvyE6cJ7SOa2lKuM581ezZwbWYtKhkJyRPa/IMr1nB
v2ICdFf5rD4GfDEn5uvzSldX1wumETkrj7Sf7WryeJ3lGEPWE2/Hn79aExojbzmW
Ri2De+MVADgxu9nSJaF+8HmYSFvtBe6C219NMzSkDetVXF42IXh/M0RxkRj/EY9G
UWyZ16IpDg+qCP6U8Hzf4ejgw9C187IB2yix9X+dlknEb5hn+lMmqISJZWTaMAl5
ewk10yX81oljzsEzKn75sxkvUX3lM4zM2Q5TnTWU8GthgWpVhnGBtXKHxM8Uzid7
SRbQ5jW+HcMXcaEd3k5N4kqsKh6HBTxb18NuMbS473eXVoAXy7aMiVY4r0d+ColD
RzDzvZKle95xiJ0Pl92ZzxDgKy+PxXcyhLqwrl6JPDDDX0woe33DzB3qAfDUufAD
U4l3sFViLMuqc9H7L/MEi1/cqRshP9u2COvMAqeJ4nYIQqBYaUh9n074ujGppmRg
/eUSFth6duK72o5ByoNaNZv/9zRheq5CV9aqdmK1MuLfZia1SqjS5xn5mYScUMLr
AQDvAXgf5JcfIrzPq0h1586qmnVGWz86DxJ3SsfNaPDNS1pPUH1NOF2EObnt/V2c
C4EXVXlulmow7HdSt2eI0JpSi10aF3uPoWHqrJCCtr22Nmxwnc/atID2IwCbXEhP
ph0sBK4W+kam/lGhUlighTsVVDUBb08yb8K8lbQbF+Il9SElAgJkFrTmIyd+w9kl
8ngqe+GUaO+6+y2MUreddxwiHQltoqQ3klej3TrJlD8oxVZfmtBXw2ax29mnlfyV
Wm3pMFLR9GB+58RvKOHIMtRRljKG7s2T++2Hz6MFm41ONBYlyJeuKjOGcMKufyJh
kFQ75Kwv2vbVU3NhmyRLql+VloHg1aHPxa3VJCWbivWgwCinB31NIUOHKTsDwVDe
HDhrbr6DP0On6tmIzHDHKJJM8pLw3mD98q09i/MSANTA0paqHZFcwJPXcIk+U7lr
fGbyWetsFlp+14CutmgzMt9a7p467LAAX9D2bpjDuZufOPkKlOo+Tu6Wk+IVWNan
WJYTCgf9DVJNQekMfWdblo6YD8+d8eC+D1RQr4xTvXCQYEPunHtAuAvxK7EEML6f
gw1S03EECOup+UZ4IdnkBs8ErlcRzMm739v6Woq20yudE5CIosk0DLrhox17oIZ7
Q9XMAKs20cpfku2RoF5Z1F7/XNP3kBfkgdQZOrxjMNF+vvdetcyXZVnb+36XFsN1
hAAtJAUEgpDbxS5CPsbJ4E9sQKkI7qBpAsPy/qyQiVPBTrysGiYAgmhufGiqZUMQ
hUGglz9Q8uJmyC1kRApxiKaITN+i8gtNFkFrutxwATRJolke4qlUvETWfGLdpyiG
40ZPFWDfGjJYEYu/f0qJGQkRcwIlYTgdeOZ+hIqU/eysijnQJeXupEGsJEQl2tA4
/LU9vWaMMeNaLg/ZRP0yrsmbJAFUE6scPsBfRClSHlKEgPTkzz2Rks7gL3Psk+X1
OAX3AHnODOPuOiRbARxVduuXwdf3eXaP0OttRB5ujwKbbvgWGKwCmoY9guJvD8Qt
SSaPA4np7tgoxQdM3wxXdqPfTiqCEmMAt8ooGBMsmz1Enn2fuYI+bwzcjUAC033i
04A10FN3P6pcRHA3YPeCuMf3TRk2cOJow/YCLe8YDiUFx5Vo+iIL7k/a2MZ7bPik
CXIdWdE7Ojs3/tVIPYT5ea8yhzGEUGEBqX5teaE8WoYL7+rhXKMYNsKOj65Ic1uH
ImQXEbtd0JjON51/ymkGoWB6jKhUsOenVGvdyYnMvZwSI0yZXFJkL3UYk63zB0VX
O2xybPbvUafGdzGeYjsNrR/BeOk+fX5fnXCEhk1HP/GTapODNzTto2KIc0tyYuz/
9KpWjEpqSAJbkK4wQm807HAHSOBx2G/TYDCKfwAT5vnqt7ttEw66YSuSKfRcOACT
CD8LZnnKCooPpkibJRLkUI/KlJYbPuLreURUEW/I3JhEdjnPC4yjzJFYB/Vp8YFC
bNWM4bIFh+/VZhBXNRqFPKs1k2nlDO1dp6vr/tQON1a0gEwsErRFjFI02WFjJAM2
pcOaR2Pw07hWbEI9hZw04JEzokoBpxFRotwwtOT33vTcORrscoJC1uxa5sXboyRh
mAxltVGDSYCFA815eou8eeCIQ25a36cDxTgx8yJXgZoLDxiNHvuOvkjbVl1vg9qE
52R4WJDFxGTsH0eiIqoh/0/wD2Myg7MwE1Z76xtu+6jFy9jScM3lpAPTd4DaV4h6
hqjJ/cEr0hLFM33QsUJL1DskUzVJ0Mv67i4Th0viWNuTVmcvlORm2OYC/IA8OkFd
sLmQ4VSgztSFUuCwa0S+kQebmyPpLBZS+vruvQZ0Foo5gTAVc4ecgrCQGb7eH2ax
9e1r4HhsmUKx+SwwwbqDDyC8bOz2WwN+AV3mEqLUYLa9FpJfPTOSBkFl57pbbmI4
pvXBC5qOJXqrsHTknbMGhyFe0k4vji6Vp1k6xYU0Gd3Zo9NldjXwl2hFpuX02VDW
o6kPQ++KW8JZR6q7mTbDeXc3riuYM2TKnsrs4kXM6+o0Lo4aLxHTPNRcUGxWJuT3
vaGsxW1IaQy1eoARv5mVPHpjtIIKsf8/U84Ao05+4g7ssJholegZdtTmy+9Hh4y9
Z1KYsCmyKo989HxM8tjecNHw1jucwfIz2qFF4Irlg8O0gWxY5c17aiNyLSRU4lCI
`protect END_PROTECTED
