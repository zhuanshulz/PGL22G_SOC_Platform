`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spqO5y3UrZwEMhrXFkFnfGmxvhiyRvHO70ksOSLFCNZuhO463oeInbAEly0H9kkx
tjUmR/bE+eS8sLdr5XqUARAflBgU0DMt4czYqwpqLlCsCghoEC1C4wU89USseP3g
HZlRRs/1N2FSyZdoVQuSfvis7kXagTk8cDzbtV6jszo2FCbCT/qas+9/AHx4c5NF
MfagNw3Qfk9ZR4SBaeS1q948Vpm7h3rjKOzOUPPHBWz9hzBEfY3d3wDX6zKG82Aw
s/YM5gglsPRNg81z1iq+hcMNHzUaCHI2LXnpKZ53tiMIFFeoucrpL/ZntTeabuD6
WX1OwCT2Vut5WXhRtwZyuMu09SRHKEqufiUGkFoqpaLkHYlUS/T756+AC/4ualmF
5xNDbgdv/z/hkbor9I+4g19eGGI+FkIDywkRkm11s3qjrL2F0kHJVDReDYAncgnU
/LV0DBsPdmpEEDAwDjgeY5AE6XGLnpVuMi3DNHw+wny65MRmfhdpi82Cp9OhTKvJ
y19TAKF4y/cf9OzC0c+wj9lacWyenqP2GkfSr2oQIZVr29Cov8M44BQyozjBDu+7
aI4o6r0hziomzRGrC8YWmRUqDB2m9wCsfqnGOWnsLg7XcBvkDDQe+SF2CKYMtT0/
iXHpW74xRC3ChLMc1j1YGUGT/MV1rH2BwZz4OVne4J7o5sLVHBvAiqBQatKicOUd
qQGkO2CBgOzNNZBxyY+nZwxTjlmgvI6QZ2qTpIBSRvT8q/1pTsXXZqjaJGCsDRD1
B4p9uzKd23wlt4AcrfQx5AlfroWqE3SfnC8N31RGO+a5dJixleThFPpQlZnU2m5v
IGpU93vXsSXzKehqmEEm4VMEWPU+OJi1uxUQp//AakVkSV6prgy9YEywirS5/WPs
gtAET+5YSVbJYEpk8sKc4Tllnsv2MXwHRvdxHSQQ4tK9yaZDWkSIw0/LMBM2qRNs
Uw9Paob5MeUT/enRxlpPt+bbrVwonCv468e33dPMdv2DcpbWfp/47Z/8nwY6itsR
zmAX/75P4S8kcoi9MFniS8Qmbqnmm0B75WdsDcip1jyli+ea8i9ZGq3yaEuZBCh6
C5IDqZGGBKz1ybOTFS76/54+lVrf/3aMlfjkDtK8WycXI7gEhtYXS89ZOpj4Ondm
rGdXsZgEpM+RmE9lc3Rry8/vR/8/GvI2n2eIVjCt2z0Df68Okj/TUV/R3kEJcyal
JOxftgdor0bEz7CccAuZ7zk/4Wf6RmpWxe1vlPtqRaEqwTC6a15aoHRPWrAC1vMz
`protect END_PROTECTED
