`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJwkxCONCYjP9QvO/84SFszI83HbhRhn+pmMev7Xg32nH8G1Pd5rrrbsPiKuop4C
Zs5o84jvEc1QiYoHVkiB3pQA7r5sAw7UJX8Z21jZ4MXrqRZcliDwA8B25tUqt+Ik
V1Yb3h6ur4rhT4xyIvzk7RbH98VqmXjEDS6CTKdq4guHIVr9ceVwadODMoOnOWbM
9VvbM3BdkBB9HKAymcmOVIrtEnNh/Q1sxgN8qmgrvQk7dNWRlso6y9bEb5pG2v7s
HlTOkk0SgTspaaIBdgpTARKhDk6n0lMXa7ZCQSdgqHhqhjfMx/cBAe573j3wlFJb
+Gh9jv8Nu5fybWpGSTGN5GA6QXUgv8kWzg9AH5GwW12X1ufzJ+JYQ5cOF56mzfkr
zTmwzyjqxJLhrgcGo5UljGGhWBOI5XIXHClPQvlPMrXxaLI/kuHFSqRlwr/nVQM7
`protect END_PROTECTED
