`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWzq3x6M8gWBbW6d59mGmQRyNjSwqoKREs/LoR0UwdLuEKR2v1YbQXd0BxDs1TMZ
vsCM30d4rcdaWSFdnv7mr5ITNvf+mdmsUwHvogXZ5fHDZADAcpQGTW9RCdtk+If2
m4Gf0ZKCjbLokft/GwlIWWGuiYXNfpI+YCe++TIUeNC/rvZvn4fc0RhRs8Vyi8AF
vxP5H3GnrSWG7QUo7fl5bJYm16ZuDy11vahn2HNMfKmF9x9ZIm4QlDOn0dqGW/WZ
bScVDJjBLqGXGeWKVkMnGwZRvCCZzsi+MeWy2JYFGnG0PRlDGxkYZr+Ee9Tn+fV+
c2RQTYvdcG9uRFKHxaHuQxtIJMm3zi0Su5LkDWiiyvIbp9TZG34P7OCUhhKxXpJ8
N+rrT5993YUy6gdqpioQPPmgdevSkzPtXoIWZ3fX9c1CM8NSZeCJmF1cJ+8Hnum/
mBxQGXzZ64HtBVXXdgQOea6jhe+x0AaK4TuyimKXC7NwuE4OcAkOU9KeXl42LlAJ
qXKt9wNCH/6f7E4nAduuuFtr+PC2jyF/j3BUL3C2Er4/aDbkUYzISU8IcM+V+P1G
G0eOAkEkTJZP5afZz3Y/+KruRgXb1I0xpUiw1tT7CgxwuCxoUUvsTQwSK8v1hpey
gkJHf/kRXRG1Hu0tbdVVNgBXADfr3+C911VVPhRWj533TNNcmyNdUbVhFAznFjAe
7KraIYCR7WUQLREWFxPZSJUpw7k9O+SveQceZ+EtE3bTqWMYP9xbN3C1y1MjwGfv
WokBriROsQMkczjNz7yTB9a+0gy6ZYi01gGq37pDUwfoeg93hAPc11DUJ0FuM1iR
Uo9XwKgaeN406CuvfBxZR+0T2+IC86R0YNFjYsrAHQiuyVAa9SMU9wHYrWcZd+C7
`protect END_PROTECTED
