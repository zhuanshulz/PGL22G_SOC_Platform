`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oh1sfTB6GjnM6t6NxrXDUsp0VM3bfo0JFON3vOR86JW8EDVYdfL5+ExYWuSdMDUj
f1wN71WtoTfDVjNf2Gr916jFu0sDCTU7su7ewEO5F2lfMyQch2qlpaG6DZnLClZC
k0JRoXAaU4fc8z14ysMIxHNxhkQObHvdpdbRdmwjXnPjtl11ntbE5k3OBa/PEi2v
7CR2vpvBkcgZT8bmT0jyYBD7bmRO5HNZwkLWr81/P5UAnMoV+VSqW7bFY7N/g/id
tgUIogZmH5j1CfATMsGXqo+YX2x5zPMcuvFvzxFAzKEZFxtnfB2Li/NnR98zSmha
QDIbVg57KlGvfntv33e1mo/3Ha8WzSCTGhlGcFVqyjXYiEMD9OKLuKojHOSlktj1
qK1LvBuBmIS7hVHg3zeJWySLVFSenvel4WAmUM7wlwLh6CSkT946RUVOb9I3nclX
z6gc5m/MpxPH1MZ9DxVKCuHMPoefQnmOxdMb7LQxPw2ShNtQ7GTMrNKI6u8ZuTZ+
YObUQxQ8gFm/wgJH+egH9MSXdJvfBu0mAPT3dG0RL4IreNA9JJi9UZ8tmV3VpJMK
vxQDu9zVCtkoTMYACZfZWBjsMrWz5CssLn993pvEg3rHQ61DkHyaHkJKQ/VSFAN2
QwP9sjiAjJ57V/zTdKZg2T+5QmQbxqq3CtAhz/Pq/ousqUYSZ0bXK6wYp2PAsKJ6
Hs7FjKFIzirAwxDv5lzzZMbuaqfqCKMvh81lFSUDVc0wDky2X2HAYtXjwhdEhZ64
rHq2LxyxG02upV1WCQVu8MrjKEzfJWgfAXL5ghLYiRTVkOrsLTNBGkrv04JFOx1T
CKhVKW4RM2/+GI3cj2SV0hGFqw6G87rWM0iz6T+Qdiu4HVeR/uz4fLcJepXH2fme
TmbiG0DssnIZHo87FStL9j4bHX/g3eZsRyTwW6sl/z2xA4mIXi5EoyEOybKGyo0c
qxbAMILULNVmZlmHguN4ldLfepTNp8hszaJjdBEzigigRxCJuDq/b79j9Fcq2d3b
mF9buF3sJKTR89jTLgmSMoilH0f7l7aSS5+SA5Pxbh3NSBVIEO/4G/yp2OlgD/+V
lq2hNCI66maiveSsjekhcfq9P6cRgdcOH7nRr9PzAel0NpLuCrjC0wEanJI+z6G9
YIdhnTPEj2KMmsPhnnRIufN/StSPuue4LJ1+X4lLgb0nWXzMCLLqNUVO9tavsHLK
uPy+Aj0yPh2LgJ6hEzbvYBJ84wPS0/03G6DJP7HSjvZEVVH7FD+Fb4riCJCdBbaz
mNH/64utA1Zi7nIChyAO17LSMjKXeWpnLHfNWvYCYPcqvmaeA5C+FVCUP5CS3kAb
Pp+vTJrwV3p0Stsfk3SVRWAxr20l++6+B8dOKxl3v3G7iwQkFblouOIoRonL4G3U
Guh+m7r2hMv7FA2JeLKAZpaQ6qpKa/kk+hhnYBt21X/EEPEPqstb9U1wX+krUQ34
`protect END_PROTECTED
