`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qaeBRE5G+iTsIiDDLIEbN3hJ9YO8wM4sDSSHi8Giw2eQCFw1Z7EynmzFqRuOhF9
PyxeC4Je0oca4cl+QMUoISVd076bMV6pLwu6dIWue9nZc/H8NbE4gyC82I5u6FG+
a9ibJqbaiFMOlujzUWyOMgUZLl2nC4DO1rbsi6HJtpq5qEIPjrAr38cO3wVxL+0c
fIv7Ri8tc1EkZasRCVKtUFSTP6G/VK4Q/tt8OAxtqDDVJkykVxckCWQ/2C1uBw6J
mX5ahhdQkCxQAfpEobZqhXIRGD+aJaG3OyqD8xuvp13tn6SDrrz93387xy0ozNGA
JK3r4q74eKEf5CLKpBuJB1SkkgCzIyXBZiKGsg544SEbNZOoGMJyEyIuut4LJxeb
YqaY45wR5SM9K38OMsCrnogadjrc6ucgo3QjnL9lcIqt5BZIwIrc+q3gA6s8hl3D
fwoW4jj4I+d0FXlZ0Pucsmm15n0JYBwNc9aZFFfav73bgzv0KdGfrrLJI15z6ih9
njpm8Rl5zzr9VknUxZkzn5mD+oQyOdLB42qGztG839OVWLjMIme+IUo7PL8mf3is
byX3pKpjFIi8NBngRi+0ugyhMKKwEXaTgX4kFD6/J8gAIVQy3BveLXycZzVsoORx
Tkz63ag280eZn/X/hbM5hIMEigOtFMBrKQIkqQ51jXkti9XoJ5BJETK/m4wqdN7B
p+9fA+796+ziAXE2uQWvpSQICsL1GjYVmiMmGavtJABfFAFFWU5sE1q99IoISGkn
ZPyLbGAUFKY0b+y6IVgnKjSH9XHbY3Rw4ZmAtmdNp59FBzZ5rocyMQB4eQ0w76Hk
yhFlLsvZYVtSU4RznYAcrD2wDgDbskYq7qwBd8lArsfypqNaVM2RgiicsZr9NmsX
xvero4tbgdH60qPejoX+ktdqHxwZk/SuvkX9TyNzc2kOtpnYQtQs9wgjCDJ+ul9q
dj1HwRv+5uWZDbLelWSZm9xof02aqSU1BiyeSSfKu9fF7CByZ0JIVGIBDPWSH+5z
/sDHpPE8EwwM43LglYlMC715JYb7BeN4jNvl7uZLce/89ktXoet8AHA1+qmbziww
uOmGqCswGpiXBaL7KZW3w/BrMEBrv2UcE+PbnRw87DZuPTwhfW+M1k+DThv6qn2K
NxzxRpEp2BUTtSd9s9JUhVQhqjTPY87mCz5whX0LHAt0JNUV+cxwUFkg6c7avmM6
vTfJLJhhbA+bpqlC1xmGVegtI6//hq2JW2lnACpmrXRC6ztRlsKfE1rMj0FNLj1A
JmLUGV8i+T+/uun65OYUPGMPygFpiHxRy+REkmwUhlmPMnHKnue7UNI2Lc9TA4tR
bbDmC6h+jHzRlg5S6kqLbgfCpON08vJlqM6+AXF4QXZzpZkkjv3ntyMVvy2mhNQT
Md5kFXKASinbsYGJLKrHvlEry0LE5BOLKn7x3n8stk7SDNe6NxtOP7oVMYS0GIlH
+Qy3uPAWu8W8UZSOzeibk/xDlQqp6PiRGNYcpRoMq8RbnDkzRlwJe0d7YAdG9nWz
ekX8Dgk3hDTdFig3j5HH+LDgoiVk6+zVVmsM9PWz4Dj5ceoj0P6IvIUiblAGXWUV
HRoG8wCHVf1TRgt1jzjnGnhqhW8DQaRUen/CJKOMYrOX9sVHW8MTNvKuYheYQFIZ
vP27RwXM7n756zGnLOk1r9gZr3NQbMP1O65i1ofn7U13X+t+2w5qBs/YLhjZzmnu
BbgrxLtSY7hcN8O3ISwdGCyGcXkV2bR5gyrI5felMr1aGd9T66ifFtjX72L2w3xr
QjmvmjC1VOGvRuvH3aoX2+yAHB1pkMGDpYv2rqZqYfQiVZTT7ED51KO7LilQXY4f
KuQgiGqTFESGIbvMMVHfioe82Iz3piLAWGQK3BES8ryZgVnIqSmvy1i8SwtLQ4h0
XfnYkFP7cppwPi9blhaudtTIELAjA+ipl4NTm4lhp4UFr3EmrjpnHs1METWHGRZj
bPvhojKT6m4nk5djlZc7azFAxoBLAY7ZgGPRKhmR9OGN/hTxTg/lmukv2OVOpsIy
JtFhjoA48MUObdqmSwPZrQeId1pxZkd3lTfITJaqRmIZb8e2mK+wwCiNOpSFrD9m
oAMNvU5ve5u6cjWb2/OJccyB23E5MIa6ALdV9vMFp85C5/efXjc1B9/gjBjswzbA
ocgu7rpUZpzUIuw6vDrKQ7Zw/SlWG2RfjVbR5t2S5zD0gaMluL/WvonitkcHnfqG
fZvNDUtDhQQrj9oMF3OO8dRlRI/cz2Dzsl16keuUj8mF7J5L7foTLD1zVpC4tgeq
nJXhCFc8026rK7quh0D3GK/PMgoqgn63UOTj7i3DR448E79RIIq2SpilogDVZfXf
v9CU7CtjWkMeOUmL5G4pbW+AMYdrXV57VGz8Ew4tGI1xL7c2Cj5jhWOkjXRqfvCz
CQ0g7VB6aO9eTst4jLIU68SfDRw+sCl9aFKQk5iaQ3azyU9ABlXYBp4B9EvNqOX0
HvyuND/SgUkOj2ka6YuOzXSAIKkvoSg/LuYPyqbxi/msIl4T5WxJ9byyY0+ojHi5
YRonUtt/cuCKh9kxaSrYU+9vefDG8GMPyH4WdI7MRVC/I5amv1e+ODEC2BrVmIKS
OzZJ9eS1v752+MGKQvCCU/qsOknuVUS4o7W2Rkh0wjFlj0iJmT/wcEyBLBq2aqHX
Afo+JUjkfWTFlQOn4lr0qLBUSUJbw0rtDO6eW+joamLFvMNdEbH5zAqi9J2DWIZF
Bf8wkuwiYJXoeDI7KYq20UAZIVH+ZER0E8GPtDDnMT3KJTYCV4TpR46IFBCNcfda
qYu98qLo9PhDWDoUl9o3JPnwjOjew6G2FLqM5r7aryOzuLDcI2gmydNjvOR3zPz1
`protect END_PROTECTED
