`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
heQNGQEg5c/CLADY3G+OacacMQQy4X3/oCvkDV11HL5FaoNvOtXzVOhm/IsWC7XJ
Xf12NCmrbfi/aeDmhVVxQ817wlMfQbw83W+U87k7mRA3n23K1RlWZE1/lJdc7XAL
a12P000hh8XFuODyAXwxYBz9bSME//9k9ELI0vDEA5a3STCwIHut95nr3cJiQ3ps
r0+sspN8SG/VpLkuyIsN1scpXs0zezRUJCIC+mTw+pu1nB5YjPsWRA4kBD/4JgU+
VJTOyb50uw2C847ttAp+XpMltQKs7Ho0EJX1SCf10a9h6B9tDOzf9ew6fUjbBUjy
Z5BTPa9aE9+Xh9VslD3RH0GaRaVapczmijI4g56xnrwXdFVRZh1Y7A6E5qNX5oFH
/EaM6EY0iN/BmHyO+Gs4EatKxkRNXSdfpJGhONXMedRlNhh7iZ0g8JjNyf+ZMLFP
6bh4ZR+jYJgAH9j6zO1KCuKb5k7Pj3knysuA0Nwz8ka90+QBWeaUvEuOUQ20h8ZB
CLZmTZCgipkDhZ95m1A4uw==
`protect END_PROTECTED
