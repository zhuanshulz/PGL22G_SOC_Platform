`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jbKoHR9efWRT5xrQBpr2Ecaj+Q5MROqOqHGN0mXGtKNKOsOO+sm4WATTRqV+XDqB
GdR06/PzxP/+J0m0jUxFAmaUv9nyshWMdvy3hh5H43SUm80YzJ5erkQ6mQVwUJiB
H+NGrkBXZfwKI+PFCfn14bu22cv7abn58gAvYKwgI0vo7PWZSZvGG7d3LsMyUSBo
AjIW0WEzpmp38lGetxET5olJDEl90hqMYrYFXWkdLMmx3x0UIX8773hbG9bSF1Ks
pth62KlD398XuoVKLK9Kz4uet4Hwb5KKwjEw+/bNpVL3XrJKgKBsUun7Vyu7/8hy
t3xAMq/dQZQbRA0QSvyT1EvmsPKCEdXgnN3hHhf1Xh6UPLwjgo77TvZaiNWZgl8a
`protect END_PROTECTED
