`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bvT0ggUIectTa6QinhH0tyjW1z75OjVOlzVmC4rv8eTFZPPZ7WHYOhuwzPWtqFh
Jl3E+Q7FUCT4HS6E/iTufv9qwet6WBnU8noZKrrMGt6h/F3vQmu678eHvXAVGzbE
rRAVvwcZQS16hJzputdC0qdU7qszjczs5Ur1OlW8U3qhkljysQONf5M6gUiiBFt/
OB1yOTmlUpePwCqJWrdae61JtviksT8CqUP3uFKMBxZH68tHBhbVy8yLZqhq2fPR
xL5Jg6+Cl8Y2Eu4s+YZM9jpcIUWZT+m9gqpLnfaNjLv79RXTwfKGDLWXe9cfIbbL
Jxt+pGgSC+UD+Z3dH4d30rWvyeaQnG0Ny5KIXiQs8YUawZZbxy07/LYWJtCpLIvJ
1WNyP3XQI+FAsNop13PNbLbNPx/nT8JpE+xB+U9gakXcry56WhcjZrJFbp9fTGuY
+07QfBzjq7naLnmIbu35p52cPpToznjMYzFdoOuUxX3Iak1bhMtB+XUYXVnsaFLb
9jzJ5VroTIU4Xw5OFfdmPUwqpXCd7gYZgQghTHu4IQlDRX9mnndjLWa/+3gDuJ1S
D83SFRt9YgUdvRzOlShYBleeELMSaP/naaL1LCmxBS1OAQF4wBYyVBMxihXkkMHe
bKM7XLIYjuM+tabU84/FxC1BNimIhuvLDb1Vb9LqL5m+AehqsGnHYQxb8TKfNAm7
jcJFiiEDqCAa8tYyZFiQUWyTCRZxOMn1i0kGCwC+NgXSSxOHu/qLWjaKhk62qetz
oPWBY7zZZJ4viWe6DIuzz/6H3NvjV8s7ISfhyUHJhvlpv7tdNL6DAsk0/8l444cW
OES4sg5dYo9BWw48E1klZMGT1OTat66Aaq6w9b0RdAV9T9+TBsOqMj6+lzTU5IbZ
r2A3qSKHrZOpIb2aVMvMAd9HjvnAYLF5Peicj80f5Q8mL5TJ1k+b7HX85Kvrus6A
SLr/QSkfGyl0wVXEkMmEWXS2mLKgOLFT2y7AdSOOoKMEGK+ppv1TnzwBwwz25RYR
UGx8NHASqaWNJ29AwEdoKJXdIX+Funv1Lq5d2tCmk0Ns0EpqfWf3g61PxjAaSL7l
vzjBXTekipTs+iwvPzrwzmuaYe7mS7zDVhDKeOcccaak4kl+wgWRsQAdtJ5tuDC6
7z/GpKSpreZvfqwMBQHyqcaZbsVWM8/y4YZiy40isEdZ/p5CeiaBPhjE2zgzW6A7
ySDvytX9rrkD5Q8aOIYMn9OQeR8jSG9IEoMynwUF5AvUus9voF8tnXM7EP35Ex/0
BRI/DypgQkEth4LvuAG+89znKorJtqASKzycA3XFWSdNkEmrmKDS1lGQ920tlcIp
gEFFhbwqZ7EqrWLSWTdgRfUq2QZXUf4FUecl8LAUDVGQbV13azIqMvOwtbHLPQ+C
F58G6QginDJlof/Pu58L+4l9a5P6iuj+utmTpIvbbAq03uKerJQyL2r5dkLAK/UR
uigTQhb1jbnTjESKJtE/8j5TD7hwJYG0umq4twXLlf8/UvYApV4mfu6qVtmcgt7M
YlByLHAlzXqhouyKBUOt26EicV73vtMhuOB233U7TZdwQZszGuxVTVyizI+Sfd9R
/pNlLbU/IAZLYxr+4ix8mDPUyZNNb/iXFoffkrCnvXdeMkwarvh78X2dOrerqnXI
2nNyxLu/feW9jQAdVkPgHnfBy8AViDbPfT9cZEIdWVp9kKjUtWjcH+u74SWFcPGc
hotXNQGhLe6b/Nvn8rfJttU01gcQiXzeQxfuVUMLON+Nt3StyKfcbZXzBYSBMZoW
CETL9FjrcmZZDQKOzlwW2bBI3vKBo3+3tnmrG6YjFxx3qXPuNBONJ78JnsEXzvIS
BJHxOAAwD6LmxxrdTEwRs2DLFdp7TpT5TGANNN8HxOiebXb7r7yP++XTC65BsOWx
Gud/Qf7+xbF79xk9WW/+q7QbyamVL0m2Q+fvXNCA3Z5Erjftjyxf5NRsy3h6dGPk
m2SQ2jkZjtXwS1//q7vEadisPQEag0Jwd0xS2W3i/g57qqtDg4GqJRd9zx7ye2oW
11QYT5lo/hotGhV5i5D+UrXWAbexQAmDQ4hQqdf/O1MNrOzv+1NcwotL3KdvFHf4
Z4JFO1P+No/GNrPJznMFKP2RByFwNb7h/bNmjPVlK0Hbl5SKDKMiFJD0kaPofkbj
SVRsGLbit3WW0hY0h1IJT7h10W/genon2KI8+Wor983ITLLtMJ739XcY2h3/cp4C
JhNeNM5SnDHfDx1bPP3x5KWAKqjLPuJflKt4yJyuBijSVZFX1OeJ+fY/AGzQTmXZ
t6SPfhHcmc1pq514Gh6YFTI++5HrdJC3NBbmSVz8b9cs2hAXgYmNQi0HikSDVbM1
qQYZfflYOnPH6Y/SoT0wyf5HSNOYEGMMztGodJyYs/WQ/zFT6F/aRBOw5hDrksLH
Z79hp3MMklEPFv5xzv3q7e6yyjb2wOlHYU6f8gg7oXZe08BBD8UoNmjkjf0SWchP
aDxu9HnI8UYBHilo+9Hz1yY9H8Swg1JX2+4ilIu93OhBQcqAYGRMLP1ydAfk89mR
I5r6Co9QxXZijruOnyjm6z2ocqX9LPL2a/PXOoIcwtxHqwpGVuWSd5wxsJ9FwZuU
ZzdMXg8nmSEBsImCFv1GWaShT+qHClntjRpdJDp2F9rDQaw572dOyD5QkvI+5ZUU
4Ox1wcY2HQJphYDC4BEdNKEvH3T6jAuR7hyYBw0Kt5YU9+a8rlvAdSM3LUb4UGmp
vTiokExUJUCM1nUoEWV6olDukxl/0YZ+pwT3p1y/Lo+3MJOBnEeWI/TyU0Rxlas/
Wi71FF2dNBxSuAkC/PWpuOsrGUaosJzBbECQZbetUtbB4J5KwotNfxIzETANTK+5
bs6Cpz53Pp47sx+D6Qi290xNWloPXX0xC6qOWWnAGqI1JXQTqp/aTLnhTfvP4Y1q
/DTi1K+QR20XtThoBg9Mo8Yt6/kE0YlQO+7okqAg6Wy7ktzZSj3ZLSAKX3OBJB3v
zi2I/Owc6n9EslYyEApD2fJMb+Cm80IGARUSxaR1bEttlBJRmxhj2pE10HtNGS6K
iQAKdit1fTpIpNx/thiiXY3mKYfZmwZN5uFTjq+zePfD3XHvBvbYkgvgAlTROzKY
GShVyNFXSRi29TP/hrPImOWUWSdi4Jt7FzXd5gaTWqIB78M65IpyralOTXjLaRu9
CBHwcTrBgq2uZdvcP9M6PHsJY0qUKg1DE1LLMry4DC4RDqat27LRiBxoRPsLLh5Y
evRpoB98VL5HzwSPrefH1JPf5wJLGSQf8fE28ViWv6cqSDN1GLJMx2oOwLAFlIvS
kvEzgcHGC7YDklWRkVbSugQyvrrSYbM+KYJW9i33Pe+mBRjn+Lxt+Dn5A9uWDjjX
Uf7QAr6LVqAZJ2M1QJYqCEnL75JTQAqv0ligZB1ETHbnggbDEX53UbMxanRsXpGx
EW1/XkoJOqK5LpHNiwsr3kNaqEKgPjgrqsxDg3Mlh9YnkInqEV9e1jJUMl43XPQ5
WIkG0NfaY4AQ4g7kuvzNklbw63B7WjKJbbpwz5RxoGAFnu40kjBMYm+kbOn6t4b1
Hpy4tvbN0UYHNMQbioM0UL5GIqM6CNSbU50jb8go6Mc8Pp8HHI3TtcBtbBVfJZSK
GnPO1aJQmGBJiJxTEodxnDnQdBsZ7P6gFefv+16fiQ4vwCM9Q3IQV2uutJN9wd/U
ne69LTC/CiZTccaBG+AWUxuFZjRjXcSkz51HxxutyWi6yOvY6Lg8kFD7eWHtLgSx
PQWSb5YLjiSdItC3ub5sSNuf4NFvFsRX+QtYd0ZJRvj6uYlui7PuQvypFDmfN9if
2eayt94257vDoLdcJ8sugsPkM4lPyeZF/eVFMLWj9CrM0p6gKnYj2gXOZhQSjbiX
vpgvK8CoMxtPdOFlJ9V7Snl/0EtiNgJmVsUwvc/vyiZVXMCF4ugVXi974DFSJ79h
oco1pDwEOUTcN+xWUSFO9b4ojofid4Hi6kggYIBYBkEXL2EVdv6x31nXxjKI+jjZ
eVynaVICsu1VfKK9BAwyaNu60tAJ4K/VhSPklJ4VpkduhrnXm6t7qVMsOSjDaNnT
SuglCxqcswkvh0MZohTPNB7prsxDVKV1CX+fXjMSrcRUal1yTCftkgRbmavMPpx5
xY48XLKC3z5f4HFMgPv+kUshVv6lzSGoDH1I8OZZdCCGBIYWMpGEylFdPHvVqLll
X4K/WnPeJRVB9/9kH13uoyJWgC+MiZKnZKjYBtZ45NMClGHpKXvZ3GyqvzeEC9Kf
BRKpETKu+fdFD2ZGu/rrUS7/f/8figkVM0qQuzup15XYzifk92ciGFgBjlbYqg+o
tqYUlyTvuGgSEaNdkRDuGc3g01ZvqSwkcJ9STD4wZR9dw36KN5oCoLZc5dFvuJI2
lF0sT/alcyKYBzb4BvE9lJbhbmL1saPT0eJhJ4rN5mRuRpyOs0PAenRogDvWPJ7e
yheFphEbf5yW/qXzGp+YY2E2tp9QtJNuKkpPp98JdARTdoNDyQl6E+809AtSeOxo
9l3ExeFM7dg0n5c659Z+siqSo2LEMYgqxRtvvdkX2/YkykrXnEISY3TEgIJ1TnR9
r0Jm3KXD+OiX694XMxQPsKH0VtAFO3I3MQwsmJXkttGuPUXzyvESyKDRDS0qbQl+
m5iOu/u/oPGGiCHIdRyXWzicluIEXus7azvmt3dZLeel1XX98XDGtO52aIz+QND2
O+voPulcr+n4USOoCEBMn+yQMCLT32ldLwTuKEGdupMAAbotjqpZ6W4HN/1Q3eg7
09uFkM9Wb9Hsqjwqj2CAjbsR2ZOVqd3sl7kh2QxlLIINGYukA/06AbSefVTR97WV
lKeiYPPD6Xk9wEkHoB3z4MR3rsRsFtd5E5dyAFVLTrpgfUmrOk6dAre9jQ0eVGXc
YzQfmbZDSPdZCqgCW3fup+1/+lv6NC1JMK4shCI3SFgDwyRs0o2XH1B2maEhf5V0
0h0PA/7XMrhW+33WGjJ/aU15D+lvWfe/dtPYkfg77k7rJ3S7dwwIaXBdoYea0h0U
FCjoe3m+FMjqXNIyBcb5VH7YcVdUz/Tb2G+LSAywoTTubmAjhzYSlyYRbNbUezJu
qfi/w3W8Tjoy87ZmpNXreYu/F3dDzk8JfAuvUHg8Do/oSwe5OjQxOdFhxd0Gm8QT
hAzIIMiFbrMtxexpQjXA1PR/oO4E2AH+Nm+PagSgQu3MDLQc6YVMV+dj9Dwv88FY
2uv7o31ceEQb2W3c0tnqwS+L/ye4K7d/nZmkBoHNaCRYyHW0pdFI3TrxmJYiLK/D
FAMi/X3gqReXvzPEcG7rt91jCWLIbI+gth7YUpNt9HwXGZZUZ4cW8fIhs9gDm68w
Omfd4cpXGXpC2vgwc13wSJTYegUbFwvsT4/enzc0Hb+l9Ea0EcgnuF3czgj8ly5g
MoImcLoTTqVq4U4J5xGWmvp0EMose9pTVCuguh5uZv/wMMkzfRogDDwnLR9jK8xc
RT30GGUAiYg75qCn1sndCJrhs+hgN4DKui7V8cpc4V3HK+sqONT/iLsYsECHirCF
Cvc8CyCE9eTRv3mB6xHl+moLDhWtB9oz4KzISd4CYirumAAlv1EgyDYydyc4QrHr
X+ODVgKoxlBfvXOatuysFE87W7/qEECx9HQvquNlHdspynSVpY5yLbPUMZegypTi
lqFsjWEXpHzIXNs1DR30CZIsgOEg0ooIokiuVx7bCrauhPplQfsurSrFFURrJlN2
RJoQ8IZ7aKxMyOHISmGtRAKhEsP6ZJkz8Kn7mD2MjDu0UkfXVrtIjXzKnb/ld7eT
Z3SnCWAKAtm2lGm2/eEVVdbNENm69Jkd3k6J5ePAq9RkQ2fL9/I0S2rLDAtqjpPL
Vf7vlS+BPuXTKAPf5QmSjsI2qx5+RdQBgo1frKLbsV39ALd9uxPh7U3gjk76FDlf
8O5kS9mGz5QwZYmgqhiwi96dgVkmKH6fGSqQuiejXJVe8whOhNjA16vGgioQSrz+
xx138u71Xv7m0FvCziH6kEjCIfG6uaqVE4Vt7eu1yWSlKQQfZ95aFTgawPbLddPa
6/X8dkUhITcFJ58qy99m6+yZs8LbV27jFLJXpWCRoHhGf0ip1BKX08KtOMraq6Jt
qq7tMqyjq5Orhl2n21GP2Ek4ySJEyjPNcxUtI63KTnZhtMCHDf26has8tt9XEWam
su79/zK4XtXwGuzFMArAgxkExS3QH1P1rit3RVdusRbYgGH+vQrboa2pKxc5fqig
n6M54cZxUzF9xsUq6xTiEa0CzRDqf30dfIhJB4uhGapBlDcOtplI7L55sWeK0PDf
kYubkVVaTtYkn6A+goLFFRcrELTqF1Fd0EUuUDPU+5sVYJenr5AsXy69cpw8Fikh
fucKDIMF6AIiKVRzcsIw2Gln2oljlvILBnNhz2WdHY0vOoLqZPKmQ7UDyHnQpquB
Y1tJ6KYgps8R8yfcD1cooPeB3OibvtZFG8DhCte/sfqu49r1SnmpNA83681eADy9
m7SfxXzSjo0TX1qguTKSSOtSIbtyqMuMSVciJGhBdxUg5KpUyBezQyWis0srh7Pc
6UtbDyTjFBds+HgYpDVEhiEgBf2jufriM/S4Va7YO+Ru3qarVRQqA/lhcPdWm72i
CltEU/uFevvV78y1Onk15bcX7rk1E9PJYjpaSB51sW0jxz1dWd4wH+AIl2gNZFan
ZJ2KPti5p651wrzBOfVtgLdS2eg+IGQaY5FviRKO24cEYqKq5ZRmmYNTSAmE8A/o
bUE79QDCb8lUNoSftPQmjff9knHsSSIsxsR5OoIlNUpUFrSjaUPFgb8jKwwaiA94
aIrNhCZn+FkQI6VrrjF8IkfL26MwXXYJY23TS8cqe8JLJKamFLHRr3ziDz3j9q8v
2CMqetoqXzxcz3yZoYUtdxfTmT8AIAYAkZB69ahDEQNgJ9GXokYBgF6Mp8Z6eZtm
w9wttnCMiizU3JCTCd0aZk7VLB+S7q810cpvFSixdWEdsheFkhd1+Y+5DyoW4f/q
cF161/QHaOscuqSEY4nlrV6a7mLTkZviaIpiK/Zb503uZaPq2VxnoqsuVmuX2QRF
ZPh8wzj44xvg2UEFsyWWzPxyirhTW0ue665wDL4bSJ1wmNnR1l8jJfZ9SYk1JL8e
GsMI2QiI67Iwhj3NRfsJES+TvSfdYVCpYd89wHEFp6THV/zzCXQumO57XxaF3vr4
qq98Fx7wSYI5q1PH/t0kCeyO1DVDUtDjROR1E3kzf2oZYTwIHJfQB1K0nbOcgoW8
s93akSM9kgpOOiFT7ZH6NIxH5JUINzMazSWjM2EtW0E5ivYdsKnrd3QM9aaZ3Z+/
RlbnEjkSTc7rIoG4DLhpH3cBbysj3apWmzLQIG8rVQ0bevOfu16rf9g6wosdKXbz
30XmaJmAme9Na+3bIGRJ+utzYGwL/npGo8sCKPPMwhfjGSWS/ukXlOttMOnaeP2p
YfA+lzMIa60r6/gms49xiafqZnRXDs7Yrrf2yt4nkZxvfeQGgLuU7YUpx5OJvmNK
96LS7tjPx8xmR5ClKAVQAs3wbmKwRV7EpyzRxP3OOiXZfCeoVRHfjo7y25e6NkxO
+vYjofQ298eEs5HbYrOvsvXy/G4lLOTeHsYZMgEhldd9GtzLJSfeEPZrc5srog3q
uhqMV0iz31BV/Ss+LhJPIFigIIt0pFwYjXXCe4kNcYTqvsTmFA2ptDYrFn6rzR4X
R8cU1iOtC6BFAt9wUyWn6DXlWxkQ0px6/5zAg77yW13+ekciWMu89/HUK/1XM4iK
aOkJcjTGpU7cjdf+ZWNLQSycfODbXw6Y57HUFVU+aGWcYFJc0ZEhIhqKtuSPeZbI
FexOqUxIgU2jtAfwdrsOnW2Nw/XZnRgYD7IHRKGLQlo3B2eM02nrmEkY55ro0Hq9
c9fOhFGaKvHgoURLfPe0PVgVfccJ+OY+bmEnJpuLAuGPdGjuyOeT8kE2JGzq4HRC
+F5QV3PiDZC+a+6KuR5su5ty/QwBmHg82bRhOBRZNTHSZZgEzc1bI2sguY9cM+dY
2jI7aDiFuFacKdRyRYfOlcnjPXZ+ro8ZLewVvRA1sR200ytGQ7EHGofWw0cxVhDu
bQxwieX4ZfKpfoTX1cDbHTeaa+eBu4bCTdWpDD64bgwE7eARdGAeHSgRPh6+zVdm
ekJTckhTrpOTL6OIh4z5yZCkQ3dUgG+oCWsbGd/3uJwyxZWoM2zklrRn8+hsthwo
qjFnuRv9edaZ63ZV4KPldU5/l8Uc0UWr0fmRCvxBKB5gTktPL44TFiWpaiDH5fVd
cGIHnza0iLu5xSv/SjhkzK0SVz7nwvxc2X9vz3YcaUmwgnRfssofUhD2/sYDBET7
i+ESRR4r87z7cbz/n0OTFArMcvAcA3suFyIiOdbkSsQ7D96ERR0xUHTFaK+CLqVe
4egoYTGEGWeI8vM1Kw10EJw4tGA56KFq6Irc7RJkFumpF763WPgyxxsAVLYYxfRF
JNslB0FAotJPh5SxT6eoVxhFO0b2iQmw9CqV5UzqP7pGsGVOK8kuhG4Q9kxDHld3
HUS9A1xZIAGI/YF+sP8Tqf1rEtQvYARVovWkHQ4DG4Dxe7s5kQbQ+xgDlyNEbPvJ
o+r4HgfoIt6yzFQYnwUBzFaAhmH6JvLNgjzJKZgYMtAlhCkgf4ERyykHepgi/2L7
bC3fa9GVgvvsG4BWqxle733EMccggSb860MCyf/1e0opPFrwKTp+ISwXsc99STK+
EiKvInGZPWb6UNoJmk3PS8ahC8+8OdElTainQtDwH7/YOKyviZ2ILizBeL7xpEab
cy3WlVDwBdN2LBRPA7B/KYW/7d6M+pqQDfWf7FU3R38pLdKbx+ACJtr4O7V1oCMC
6cHsl1w55WVji2Kug2cAgOtDXcg/l0SVuLz08Go8RANKTZNQzGyyZH5wTP781Cyn
D5fiEfkqEr3iXY7++fkFMiWag5iEOYkwy0EdWJOQYAuuDSfsUr7OsxJWiYh6VUAI
T76d08U1xQ1bLo+Zgdk+AB/fPI1r8zDJq/jNDUJgo/a5gIHgRvJxZ0Zq+szNxFiM
NwrTCrBHzM486dMM9/JxCEtDHg6jY64jWhS77JMi035GpLzf30LxkWmD4fxVSECJ
PRQwcBtfVGl2U51XFD453mECTIaEDBIl+4xWcSH4Iix9V2dVTjjlIzYLiFNlRwCc
6WUJEVfbbI/jFXw7cPIIM39GbUr7fSZbG05NgjV/MB+EWIorlrP4+RpcmHYy8v0e
XGKx01CrmxxE4N7awAePu6J6M9C3wbh34M7wJkZxmNHeBvYFGqRUBNF68BmSSMec
ecviEKhHco8QKGM5qjxswUS/zCwmWvIZKxvxphP8x/VejJkHyScUH0OnD/2O+5Ii
AUfWG8mP9tToS7jqrymGmcfLOkSzUuEPqwcnUzQcZMdUiLtml8MBBsS6jKkAdyhX
Yo1n6Yd58cuHn3oD4fBpSzVq3NSMnMNJJ2fA9fJNRIHawmh1InSRc1qKiBNwRhCX
SuNrVIRz3T/Lfx3wQ4fDEQhU/mYp8YvzRD9WI5GOizi0R4zm8fx4USWwMNhJf3FA
ahtkvnrV7SLuA622Au2LlZiZEON1KBj6jaNWmtcQFp7I14J/SX3bXcs8aghOY3UI
GatwuWqTn5zr1Dthw+LQkqOisI0HqSyIfjwi0ihosDhhu/5wSkm2SWN7P5To4o2J
ztD1OtHA7ru8TayA57lGflfv4gw8onU/POGBM3gbFBlbry/xzaI9WmJCRdAteoLT
4fWlqcsd4iR5dESf5qC/6yGBpFPqA+/BCoEP6hs/RpyYKrHvUOwdFpTZgks83bKP
nss9Stp6oGkfcZ2lTFnHP0g8P4A8gcd9fSaStpTTCKStgxE9P3mBP4WvXdTGeVMt
6JHPvefaz9shJ4dez30xoJiND7MuNyo4LUIatWB8JLmpfTtDpMrU8fFozCMo2c24
pVeRHRvuutgI3FppYuaHUNH4GIIGtqCdBhaWyFiecnRVz7MhEk6oyOJs4lzpU8uf
0nKRm/sFJ0lBcyzkjPvorXSOSMZNtxq1UtryqhreA2Edm+Wus/CRmXKOfveYVyc+
HssGmRjrRa9hL4ME066XXTrViwkMyoV1sq4EBX1UVphFq18wS3D7du22Rozidnei
TTesdrIOl4oTAEKrjNEMs97G6i7jexirEfi7/i9d09J5UtKNeOv/jhPezPaSNbr3
kaaPzPn6ZXcr1JWi33EIduVyYSObjMLeaKjq3xnrbZ+svzhVBRRzMcFZyHR9SXLF
Qx+HjyGrn9o93WuCcDP0flAgRYP1ygJB7x4ktk2uORZth4PPQxnhISve7XPeYVEj
2GQwpn8Qh3EwJKvx9iScThXOLCz2hEPNa9LVsZd+e2QvW4VE3nQuwjiDL5XL8yRR
CHWayGrmitYZMF7EsDK4j6SxW+onwX7KhNYOiO4hGQG0jee21zkcS+g3y8zob1XS
+ipmkaeOTMPdcUYEEKjLupKEGFzxXVS0tX5dp+Xt10e6tJrfqcOi/HCvFvVeEq4/
UcFemlAkvlW2Z2WKGHoQPj5i2q9ct+cU4ZSKEjlCBhsL6X/WISCrqDAjg2lHV+ex
HUhe4F53nfbgX69VA54yiAE13jgFfl/KNFP6WftKN0EwZhgbI9YlwpPCFj1BHiT5
HY8PEs+zM5/+lC/iAxCcCpkZK0VwGzIyYPTZPfI3kZgBXNLTM6M/+7yxYCiMEaKr
0lSbtO0RjL1UYl6vzf/c0VJs967P3j7Uthy5B3z6PjjXB4L0ywrD3PbCEUQPPGfG
hvoVUQ29T1txSxhGK/P0vMNuc6e+R4sQDPVd0fH4qbYXl6iVKxm5fCu71n6J+Fp0
O/EeoBSt8NmxoIi4UalXrvUhtnoEm+Az3KeI6eQrdpTzZxsix5HetlCUbXCPAVj0
bW6kYG+NxlI8yBjjS1dc5hwv5o02/SlpfpWnRFrDXPmD4QmGOVsKCddIVedg9R34
OVb3FlH6uccUIF9NMl4XZcZx9Oynr8qu3FJs3p7tat9p4HJI1uIGJKePOfS4s8OI
AqQ/dka8+a+myF5sRUJ3uDLPDRUkkOwOW2YBDNqFgGIvyj3J3V6bxNx/ZrS/KBJ1
wiviAyNbJ5yKmIB0fE0cEyuzpZaLw+KEWYMa3QMkPZYM7A+Xrq8ByfEf+Pe8KQs4
zPd6p5m4ZNV1kKulo+orwKUfaOwGiz8Hrrz85qkrxahM4N5+bulXEbIgbY18FL7+
G/9F+K+Pla+8gsoWEsVnIjdTx/BNRwqTwJ9Smo6JYddDasImLduTJ5HRHzGM/lyC
DETeSDr6tULez8JUasc3W0DCo7vTXvbtzCyCqg3G6CmF7hos8d/rO2mmDgEp8svX
eXEknbc3gfKv7AiXh0ivwySq6TYbOGgOj1Rve8jyexak8AAyVuC3EBtpCPf8diCj
SE/Z8ZMfTI1evgm8aSjd/42x+s8nfe3ajDAu7ps8t7UwEZalo6f2bAnFDE5Qp+lz
jYOfPmx+NwW1SuIGl0E+CXAqmtHJ5kXkTGjyBIZBz4rAIswL4Do0OVl9mm0xaYUt
BX3aEr9BF7O1jWHuKpnXfgbjW4Aw8u7zmTdvaT96PNtmzEvuGmZY26FW/LayRIOa
H6QV24qy0OPt8Uurs7NmTHSnZ22NyeItzPNHERdQn2+aR7u51QfkTbzpPIcJqXZu
cAzBm1bUNnI1NR19aMTUhp7jTw2NHcuYh40xzzSiGkAszY8WxCfjRWoiEk4k6XVK
M7oV9M8xemrzjzeAmTKqotlnAJuU/whM1hejjzw0YECYt02zTgha29AAlIAFmxh3
cClfMh0HecH9jmwleWc94LMnGtaO/xf//13XZ/oIoIOI7ZQ//rDI6B0jsrVJ1Bf2
vZz8dxB4FRT4EBu16701xpF/GREcX5UsNuClY/Urxafr5rZawLDSr/0LVGxTGuQn
DFuW23W33EOe5foH7BwnZpabFYFHPUTWabO4PZzA8YrKY4aV2yLABfXs1Nt8SF4i
MAEaCCWPFrktpWOpkHm+W1JtjRUlajnkWnjbS7/ASCH6tyE+NIMUVViTk+3bMCaU
N5uGvY1zos8ATJMMt/en6KEiHmm0JNLLhcCtdGN9ugLK3+nuDNlBY5xYZw1kVGLM
2ILlGOsTzzLWCpLyDBdWVeqKUTkIbBs4g00bzrODKYHJsfpYZBpxARJbO6u2Ka9A
HCfs334L6UecmUNOi829iniIT4diK1RJ1YvhBej/8gBub1IOqVtx9WXnRgU0FtXG
McAU6MJv7qZKfiWNs4EC53juP/wruojEFfPG2ynRywgYoYbL2VqSA3/a+Oa+zVIb
euplhsBFE5kver7Mlh/hV8W/t2jzv2lFdJa4rjdQm+JaVH8AU6CxfOST64nwAHBs
CDKu2OdNks1Gc4tyjrH5Olg7UfkEqdnEAjtV2q12cKP2Cril2F2bSoJf7C8XaGNF
/SjbnhrQcFyVO6C56G3yFBIgSzXyv8VtAHd0Xm8voI5d3Z3q7tYKBWRNZLj0QTPD
gYAeQNa3EHkuwugkiGKwZM6vxot6B5/z5zxG1Xw9t+7C6JKjmNowNMttS7COISdC
FtxKWME9HQcOknJlViVvguNC1r9+u3MnknSv4dG/wVQmyLjjJcfTOgiSKH2yJVxU
L750alFvuQJB9mY3qspYfCHIsZL+HfVI52KhWpFMhv2yoj6hsue5T7CxU1s2OMr1
rg5enwyqlz3qQl7X2qKqW0gWD4Rx/N2nGkV5ASiM7iFK17Qv9wKMSpKOhSPFvvQe
lmUc5JZINwEmjHJFHQgU+efxzm7kA+WnbmHCTPROJ03N6YH8AE8f8T9zAt7mrjVb
jtqnNswA3P5Kh6+SyGIEepaeXd1QBAa2qj8h25wd90Bj7Lf6oPsD47Wyfz/ejjjg
PxeWsWbwGqvPaNpaaMPCYmzaJ2XDay+eC4U5NBPRhWHUm8jLFnKTsS8rm5+loZ7c
22R8wAXFIXwSYBp/Y3zgmqQoYQx80SbkXW2l8xi/dWKSHBqLFMP/QEzOK42Y19O6
3BdUQx3r7fgHL6cXyr8yZPJuuyAlI2Bmg4J9qTbeFyeyqFmBsclIbdEW6ryRsB1O
Uo8VJf50u2XPDf5da7REQEA9t7CVh6csNyIOc6i6u37TDQNwdihfMpM2A43TFYGF
1Wjsdj4wvwRAQN2wC8aneIrnADWj7ip4iKOay2LM+b3S4qzLK/BL1mzM/Njrlzmf
odik+90EybIY1GxXjcecJ3wesLk0D5Bln6YbRb+DA5t0nbHBHWsZTxb77nxTQCMc
bL/YfNeQdhtr2wj9pgJChjmEW0NUjs0PLbFutlyyOAkSnRrqKuw6MCmtZ24zwlQ0
4g7645MT2emS33F7pXsfPusy48nzj3n7ferGv9hqGmUxxt3zyNnaiVCheuO7w3vv
IZukB9qds6No21pJAbbEo37m+rAk2Aroqs7o4W0qwfFaKdYlYVoyLsPtfM8jEzAP
QxIF84L9Ka+a8rv5zKE9T/po15Ft5SKlVsht5T2jcy7sHmS9mpkN5mAu9jxKZTBi
JRC1NFz2+F+uiCVWJP4oWbBFTZ6FO8uUzSJPDQxcqH5f61NjQkfUq5mZnzVVtW4+
ZJWZ9s2MErxRbv7I6/X9pEphUgBJ2HCEk9CcmBD9oXHBpmPEwaIN+3JAwCPvmB5y
s6AqqZqAhfd/xgaCwQtHb+ylNy9i0xmu06gtYxg/Pc6rpLWljosRbJcMrytKMSGn
qw3T+0VSjvaH/DuVZ990GNHPjtWGvIr9+kONX4QM+CahKSDBagpGkxO3bCQDUXkZ
kyUficKOPBQE2E2oelX4/JUgtlBumO9HcOpYDBXNeMsKLJRqUC2KxAYc7kCXlpoa
k2ka1I/h7jnQSVTL32zAIczj3i/lN2vZvQQ33WWwc7oEci3atu3p5HJKEv1Y06mt
4ToCO3CfbmtEvoSrbAEF22gWxWl/uaYk+1xGCOoptPJJ0gwAWGk71i7hrKhuyVH0
ICXvWbzJh5ksQJW2B0AOrJV9UnVVLZ+CQRotnQBbPc2au5fEQC9quBBXtS3J0gcK
WZMSbnPRx7pq/hkTYiAZOatQKCimUGW6naaXYnIWWt7orOdeWeHpx4AM4Ei061TB
zMiQhdsMRAE/hyI3K8l/1N2owN7biwreWgRnBoqnFDMe47mmieLltjDlHd+F8Lnu
yctJ2YNDJ4eDmcpsSPnKR5ze66AwvKJ1NWWzASV6Md+DDQUuZVa0yKIdTFOtq/bU
B6HDXVM8LFaUCp0muVEmSShBKrtJ8bKM7915zVjAVyhKR1eg+ASpihG8i1Dptmju
pPU4VF3HmlRggNW6s6aSCDskIlNgFeXMH8e5FlLIkOkI0U6pRddJ07epsM57aqMK
4MErd7vgce98IAVvznZXYxMfdifh5ifI+T1XoX4jfTEpO2WCbh2/NKiFndnUCVJ/
ROwX4/Sf25HIH2PaaqUZGYOeVaB5RtEE2dUugqJgJPiOtmNcBMINW6JJOKbA1Eu8
cbe/Z7lDRNTOgzT79ypAcf7AqSOTJawzO6WQai88qrUaBXSV2OVFw3gt8JmUTci1
SshsneGCv7KMAgSXnYNLrAfCJQlwL8CTBLujQFpf7O4l5ZJbuvWUfQzoQpkaqxEX
upWhngl8NrQuGqkeqw3KhWuFm4jvHjHublAob87GT2qX58fuOjEqIOVgJq+1upGk
45yNfihJqsKi8pGvDshjKL80rrDoah0PUWqKMMJftI0hEExQ63M4QJa7+N03wYE2
vXFLc+P4zt85RkEoIMUz8K+Mf+fxxMHZbWFmj7Uk3Wq7HjiZN9CZ+ieDlH/S/PdH
0UNXiij9X5P7YV3kbI2W/uTqoY4U72curFmXWYJh+kmewpU7IsHsIop8D8bJHji8
I8P6Il0JbeoNVTMw4m7fpAjRrPehuYMbnD1fuKaIXdGy7DchGjYLZkK3xk4cxaA6
zz1/yhpQ3KNcVcQfLQ3HEi9kFlfwJR7l1X4kGNGb0P6XjWYNEqmCtK5jMh3dLBSE
DZkwov54jmZ17mDLrbNIajsGqt7Hr+8+/LZI+b8Aiypc93cG4yiK35eGgF4jaehF
p/dOo3Gs8AiZuxv6tpg53pDtFEbCHL63dfPV7VTbfigd42EBWYySU53Ij7b1zAeH
NDvebVzBNKzLBCRI5IzW5cMJh7OinXfVlNtdn6O5RuiKYdqpRqG9bWQiUpwFVVya
HoVlJYh1RnaaVSLJd0mX8OodXq/voEFgFLKqUQ8FBjN9Ku7eMLL1Hr29wkA7f5Pa
5U+M/QnJ6OxL6Spa23WJXtOchhbu5ClNPg+WswU1DlFQRGnqnt3+2ZmdlMSG69g7
EYM9KTmUPfGMSoWBl7s+MNtJq17EXXhle/BkbbBVlB8blLtgfJEVlyP13sHcxfrp
4nH0QT3dv0ZZjvwWM1qeAwIH2JLKwOkOBnD9COaHiU9wqnhFjtqcyYpE/Ewzl6lC
Ad6HzvH96p7LWvUcsvgdH7jXlJEFc3EMRokU/U0L1bgV0JxbpGNdKsNMKd2Bhdc4
0v5qcH/VW4TscEFJb5HVkTLl8z99A8ZcG61Y6Iq9m+5M/JGrz7lyVwy7fB1aEBS0
OsGJn041EABjiEfgP2DyCWoRuvwVO49/WnLijseaEBwEJ7V/7CKAv3+B/EpkBTuY
oDDOaL1i8qUnSueCYr0js6yJCWRohD3IsYbwF5xgOHc70wVSUbtZublZ0q5zePvZ
GmJuberXZWSQEI4eQxoZwlDtjGJRFBd2p1fYLtJTNym3ZC7jgDeqCouhmbh7Lwsu
W9z1v//rt212H/xFiuKwQNmrG6ot2qloNY0gFlTm/OnO9l6a+nd1j6Po6p9OWGm6
Qsq6RYjrDxadqco4OPCxOPYt+jCFtdoImIXsEd4w4o5ZoULvum0qZyE89Z/kEiYC
nWfWQzN7QL+uMKgW5K4zR3B+WIDgHtiaSLwAPg8+TYwTUU91Ab29GoNdw518UQFe
Z3OTU39JcFFucum8XORn3W/tUxhKvjKThaHdxOOsmfPSN1D7MVpjCgGTncKJRMEJ
kqB+VLZuFQjZKOhyRmzNCNwBGkZeZ+vsfJ5vMFPk5ocHYmGptxaPuwUfjtoCn9e/
a12YwYuqV1sYJbyKrcXPSRt5QiHZi/xYMkmSFFufbQhKd2WyUET/oCkV6YEvQvyh
naSlD9Q9ZQfovzTeVdroDuW3CdCsSxjgCn+e2TmBgslcPdSvb8j1iWAZK5O3Bq/r
G/bV3JfIOA/IQ2/lqzCYdtYqcKNV48s9WwQyJyh1Y6melm6oGy8Q1leK0NxrdU9Q
cSG/zIhLb2ruVt1zlrTS5yAhXEzcc+DwaXJSIPe7meIA0WSEH1PxfFKMMr1O1POE
b/KaFyFuUV1LOpdxmY5HWQha7zKM2F4Op18yx+seWLcw7ruWv/OCuG3wwCTQmd5N
MB27/1LH3PaOf91Dnhyqugp58VpW3n8pQBtFEWu1bpDaIISczZTEP32AT+rzUeyW
6A77QKleV1A/vKltSRo4ndqnAhe8g01S1r6eAmz2ojht//vaekqHx51Dvizc/hOb
yHqKdA8+al6wzz6eDLbm5J6dj/P0vOz/WeIZFKWDGQKr/xDaPmqGCS9b4slZAcgt
Ypm14BA4UbVakkzAh8jy/LWIGWLTdRW797t+/tg3+WK7n2lmPPQsqI5GeGyKxEts
RTXPP6PV0yltLSbBZLQetLmJyh3ZWIoiGieV37+in3JPVTeW9vc778Iy4/cSnp48
YZ3V6B8pxmWCurChfd5Us0pJHA84X3FOx2egkk+WwZ6/B6OVXx9mn8H+fzYikH7D
yByD2VeUVIUR1Ipei23dUfy6kCn5PESptdVZJwE1oq47YeD8HoWzh2r1jhlTu/sb
twqkg64lqxdj6mJE0NwOs+XlXPFHd55OqXz+oLuUSQH/eOLGwOKN/HAmKTJbe7DS
gD/4gh2V5+gZL7DU6bkxiCXC6lF8NCKx324ZxLlTGjid37tqb9ukXMIGS6WeSs74
0Goeu+cjbQzItBPW7JNbKA12mp+VATVzSN7msd6pgJ6Ihf/eutT5VTUqP/Sx1m91
G1le+hRhQgBdNhmiVkP11Ifcod7kBf1MUKO4AIDdtzDJjsy21yZQ91mPnioxFuY5
4mWGyc7DOE0AJgrFwgoQaUMyMFdfgoyIWlf1wT9bI1S2JqnUwcgjECD9+qNt8G4H
E2p4dTPJylc/L9js/osjEIgi2elvfcaspGxruVpFNWjQyJKc7DyxgWRHJRzjlpo5
kfT8QlCwKTsxX1rLgGWYPb6VcuVqjjsgP6U4j557Sb78Dg74nwgeCqeX23Em9sb3
Y64YBp/gwBSCP5O4uTtdaGleL7x7bHvP+hNGoq64LUr0GwhvFHgdN2Z3bb6N7XPb
bf/m44yt75oLQDkYRmpqLlbbNU3OTlRYKwl2bL+p9SWoeu21RL/74y/yh1lK7M1e
jWoAcULowilnUbS19O+WoD59sv7XsHr9V8PZWUj8IEjkPU8yzzws3REZhZ/LM9qP
pe9gqhz3NoB0QMYxObbMbzpFNuPHdbNaFHGSCVO6d97z7surBdLqSc4SpNLl6NRo
HkT8PfEE3rr+RjzQomZyAWLQ4aEoIjhCiO8ApP3TD1wcgCZPLoPICagwvqhroge9
Y+D8HZumZ1bxiulYiA4DmptLhDWqopWm6r7ivZhBHbnGju6DisFRVdj4dBFT/tWY
oQjhhYWum2RTAY0GLxnQw6gnI758y+MhyYprHrfMb1sPf+1d/fQRB6lo7MgbP5ez
J1GQwQkNBc4JMgpE+S5MG6MuLKSF3SC9h7hL06a43+tesWdxk2SSI2ewooxPxvTD
5SlksPGSmcY77iI0znfT9wphRPVsZvjpBNy9yFgTffmVUNpBtswVFGIDGXp7l7Cb
2oB0WqRRx6NiXdASF5XnL0GTT4HvLmaA2owWVJ27y2Gjb9rd+UHGKzjd9BBCeSFA
HU2Ryc+PUaTgxtzPurQxGVe9zoJueroHekHRy3/XjqFX4qgiuWrKLyC2g52ksfCC
9hbhghipPx+J76tOgSzz6cX0+Rmplr3bvfP+24Xe9Jm6RfKu+sdE5aom2Xa+40Cb
epTnp+1EnQApmWe7fuOP78UWVTozSgX7xKLrSxCf5NX4AYYrbwDUNR0M+Z6u8rFN
jq5kt+vVnPT+qssI/s4G+IJ9lZbMdUJNtOs/LmVy9IIcFMuin5yUH/zd+q7Melmm
UxxyGD7EsHuUworp17+tp5AHOoPq1jqWhWqarTqt1/ZWT4pn5L43L4x30/ARRcr8
dfSU1Xt7x0PmtBfqDtWVHIFNBGDunuQliy0z+iD5Q2JrD3VgcbivM5W+qRPcmHGP
Ji4XCIyL83c+hXcQ5dIFyjKL7YgYaUB0sSfspmQjlfqDC9AgEKGD8FSXWVOObyIJ
f+8TbZQ3Xp6tmeplMKhB4hV1rEqfhuMhjaEtHOADGvWhp8pvr7zS9jQ+t/RtHoKx
y5B7Uw1YypSGTzN6aLIkMbM+XuwdjXq6lYonA2iZSJ7oAOf7GRkq57d3T1IIhe9N
gvhYVCfEXS8Xbl5S9pp7BF9UEYJqGC/2fPJn2fiFbBwogWf/MV4Z6iB/VHXlZ/x7
TQj9Jodlk5h6not5W2giq/KgiBZwtQw2MXSJWwYkg9xajPRBUpliYMzZpfdsbS93
k5sNWftUG2sgr2Skz0SrbiFhkzhE7GR4hVXr1yXAQGg+HReiuQ6X4Xpz1oigR5s+
bbMYMHNtiuicVXr5JuScq/yi/RxI229h/5KSM5aqu6lknEGs76TPsEs7KRV65jDV
0T+ToEM+h3D/tserOvBTbgHQebqSqJqyqvUGXUJJs8vi1jXoAzgAwyAlMULDZwzJ
DveTmUiuHACWq2R/lzw4CnEuJmBddsHlas9P9RFZS52OE49I9O1C8U9W4QKlFmSy
omVmIh6F2RDu/Dwx70fSDQoMEnVIAhFC9bJM6cPilyfJcaeskEeitzX3fc5nVhIv
DMGZRCgqPCiTY33XjFDCLS/V6L7X/mWuAXS+yItcf+Gc1EwJrGUtfO1hCKu2Yrde
HCsKV6RNwhxbQpGTyHJ+VUa73NozoXLH3f4e7H99/VcbONaMtbVVUS7YIxekCcBo
+fQqXvJ9iuTFlBIrlCgwh8mPBFVia0yBC4+68L7n+CcJ/YHb02rrzKlczRo82TtP
dYgIeOOMsFlmmaXpH/JTbXgVcnz1S1Oz1BTQQVrnfbUewb/w4CPbiSSh2utsfkE/
4qs7gcml4MwAcsZ7duxLKuTgRcxlWdFbANeLgMK+1VHUHJhBDrKcs3tbraohgq1Z
O8ZO8UoHMxEFwBk1HXyQdf1xVU3NiuTSHjtms2n2t/gie+vvH+E1cx23Z8IEIMee
c6AJcv4RVWkzpUUeJ9TzOk3uYwaNYhV3jIs5UXomjp7fgZgqX4SqzSso9jsy/Szz
8iv8pdsp9LuJl59CiO1Hi9p58x0pddRcu5lwvEbyiNFVdpSfO4nrDkpuyCCsn41b
8yB8u6PaVBrYXWVRw6I0CQF5dxHsWiGlW1Z2cDy7nuA8BMJsGLvqqelv4Ey90g9C
fzcjl2So9VyuigOUm04gGTYiXF0zruWxxJGACMY3ctm5we1LNKvyQF+vgnyPsvD7
E2QQ+z4yF9ULa9QJVwFE28ZQ8csX91mygYA5LH5ZIIZcIqYCpkwxwsz+cC5R1V3t
s7rbCwXxNN48HabE1FC98iolnFJt5kvaWJFydvu4VzLLFx65aG3Mob/pEj+Qg7iZ
41LNCgFz+FUZlhMO9X09BveXjDnSFR6B1nzkzK7LBsLZGA9hhNSLfARNJscjcANF
lY5ZCd06eCBwD7ejG1x+wqtZXb7qoVh+J6iwvI57w47IxL8u9II5r7/8q8QXmu6E
yDzyxplpHRxAZxYIldAnw5T2PCiQXNFeOaPFDR3eOe3XtMag/AF1D4ajGwMTTR3M
yUiJywrXESUgP0CyNStC1trJDjgDfmQ1ovsOKP1OEno2TE/oVZ43yhCRC6kNOH0v
1NZ+nyxpizmWv+66gBCT+qbrV1HT2BJkfd6P6YKMm9Fjwy2qcVkBZVoV5sGegJbQ
PE+w1LfzYqQIXZsUHBEKdr5ShzxgqE1sdvmnCcInQmi+jBS6oUShiNxTWgJu6xWI
ywsElJFL9SGMxzMc6rSkssaYBU2kSSbXKVlyiJ/v3cY/rM50HEBL7kx9Hlk80cGW
lApTQ1i1eCItbd8FL2fQN8fEQWMS/qn5qggjm0Ls1dIq+1alOZZQ2kKhwg+KoLGZ
BoRnaoBpr3hYcd6fpL90zQt1JhS6RneHGWTnRh5DyuhuXp9II78BDSbKtwVUVWFw
wdfXXMPE6WuaB6nf9l1ZxJ4Cb8cpH6K9+qlhJLEeowWRwmDRpBbcykZdWE2ZHNPO
kVkBCNbd5leu2wBEnNPV2ijL8CI9DHapkVJfwuzhXspIYY99D0B4VLaj1lH2yQXb
AQPMzHdAP0UmEcF512QVMX8qxbmUTGaObYa8Qg/5zQep9aGPxNQPB9fODwif2Wzi
+BK9jHtj6sEcKV2z2+sFaI8YSMan3HM1W4Wcd0LWMcaudgiFLwzbMP2PQrti3ODf
ynU/4xHU/FXEIA+W9istwHFB+/vO324zeiXkJSFVaiPOvi/iqEjh7s7w3qLxWDF0
5/HXhswkNibDmsCXnWUvXdL1Bl0C16TfhbIKHzbOsXBhWHEQc+5GO4WqQyviatVx
fHPUgmDVAa7jAf2qDi/9AE4KZUC/4Fu+wyZ1c1YHiNkwadTqWrHxK5X4dTCZyCL/
vOugvG9+5MN7V8MJdLkh69P2x8a0caJPB2PZO/9fuqORa4xxEvqT+VhR/1y76VPY
n/rc5ar5XPvIgmr7gQmUPx2N1cIMJCuArkZamU3j6TIHSrKuLr0DHkDsdLdxdomz
Fsiyqil5Zz+hn4LSyTDhWrHGDhhSDiictSzZGXg/DnihJMy27SoHlkp89hEk4emS
uw8dr9+uD505HIiFxqaeRiRh2bYIyU6vJ+E12Gjewm3mT3BCfKDOsgNIG5EsFO0h
D4+2YeQ8tsUzKf7a4Rl9M2zaveUDeQQ1U887GBr1/mNCct+QXbMGPdw2U3bHYvuM
feCO/uowrefqFy4Ql50kC7B2CDff1J1u2Wp/kt7PrFvSH5th5aDccoVEMkWKKVnb
W14QL3sRV6rEaLQQcS47qVYXFL0S7vtzNl/vz9s8d0/eJUUKR9lIaib5PRW27BbW
8ZSfxfTNYsC5xKes2fBAuI/J+39utPkh/2KDoGVouBaunxpFI8xExLkzLXrFtAmZ
tWVto3b4g2n18qAjVhOzmCQjGc3Dojv2DidIpjnGkc8DozzTgD0t+f671P930jcq
R6kTtRf8u45NFsWsPaxs8Ct+xyaCyHAzTJab9NG5GvHZ4hD4oJwenWlXWwWHRlr4
sBlFHPOwuZUYFicOYGTdkkqb0nahx8OiZQJXn9eZniPBkQlAP0nSzA60Wly7Aoe3
B5kxmmqgy+ZbBbVVTExpgEPN7djMfDbtF4ViM2sYtFipGrnvh6FnMupZiCxvs+Z6
pbCbQKzq14U8VdBA/AhrlDyJ8Gnjf9DWQaRDkO+Jpi7WUeSNtkh+cH4bj0bLiaMN
75A7kEw6KzYZAAQrgBvfWBzDh3LJvmssSEhgbSLQLJLicpLkBpEHk0gztjnemuK0
M2egE1j9GM1k9Y/BLBsx4CAW65ezJaVASeFgKYwoET1phZtvUd+MJH/8ikiAeFhI
Is4opH4kUjcZ3d4XbjIV02o+ccsA+BEUb+1m7pxxFASNqUNRe7dCkmTc0nQS/Wh5
xIA23t1bIZvcqBKZqt5hm+BlUTjubIDKUaGKZsYtJWNmv8vQOF0eeVhYtHcOJADo
DF0zHofC3dwgPWpsC413gh/fKXvFuo/n4hihNCb3y+SwY6x9R9JnnJdjAvYXf9zi
tHxQYUQzWu89UJEAiiyKc9e/Ovcorh5rdvUKoqxq7j0B7xbelgkRfafRsXEVcmNA
d24ET7BjXdypAhEZa3mJmrmH20L5ovUyzdlq95FqQFDWl7P8LohSkE7y5bQEVRUq
07yuMGLvZrWBNR1nXJK4IHI1rmcNt/cm7uSbp+VlVoxOq6ixIy8DDSzMqdfRwnlY
TCXum9FA+Aqm5uWzDuK3GGcoQ/qYPMu4Jc4YmIJez28E6dOYNJUeq9DsfnW0r2T7
IeAtDbhia2v5zY6GXegX/MiE1CYzckZbWJ8gcf9AMm1JnmQDRPDuo71bQgAojMQ7
4zifSBkTo/rmfOf0G0RNF0kloCMWAdENj76XD7bjnmxBpLfQYoUgPBlYWScFS38Q
hGLUVkEQGUOJfOYMFVhzk7IE32ILrG8NFq57zznHtvEJ6ik8hLB84Tyr4Gt8oW9J
ZvnC1s3Hkt99cJlU6W7V2ECiQgwVe7M8brSIo0pQX/3/D1iMXF+nGA7AoozBKEX8
D5nIiH4t3qGo/v03iRHiVsnDeANVu0GV3fAe5cDhNCjB3DbD7SGtK7JfxItnQ7s2
biEhSAaGfJ8jNF9y+hANaCh4JRzKU0RuiRwsn7+kDD7HIfGKf8IHDVUz3ZDrbV4T
6jrxMnHnI7O3P44awT1Qw+4iV+QuAvW2ZJbv3dntZx/TT/aVuWVEc5PRbnfCVcmY
BuM54v6kIqn1Z524GPkUAPYs0EDOTtCvsEM/RiCcW5aHyOkDc/DcHDxzgYxyZ1c+
xyLNx7bmkKZ10teHYwh8koXnOH3foleXGx1tHcqs4AbZABTWPePXh8DCu7r0GQbR
QHIlSMuZ0YuU7osZvxINK73+2ZY2FrVoyMlJZVIs2UaC5yuyGFAKY1uBkSvCeF5c
Hhu+nvZGqYPh4+s2xj2LQxjn5Xsn5M8Yvj11zvXd+CMOFk5cQWAbW/OEelANWOt0
GoGsJsI781qsv9uVU9GcZe82q9GZRtCHDJV55JH61cLJyML7+JLpH9M+tOhZUYWH
md2HQR4rb0FgemMSKkzzojoeKPxagslC2KhxHK/cuXDNKoicbOGrOU6WYtotL49h
3K8eMElYVpjnVYDofE6JH1m47Ijfo7iNUzTb2qPqs5uNrTpD+/xLWE6bk18690OQ
t4rMI1AFKBZQ/3FECuNN9BdnDrVwwpTtyzhOe0/KsFIz69KQNHAlyYw93bUl9pIl
s8EsCYfYrxhIskZ2ptawLd4HABNFxsXuCbEMit7UNlwECjp84+sV2CKgr2lbua2d
xtCG5gWqK+pQ2/uFwHgFkF3z55qOmIaIqwyqr5UYpODUNq+MHFt8clGbFWvGTV/3
bx6cXRSFouQxRdDRbTI0iBF6wImvP8BGTVF/m89Ple+PcAkZ8hSF2SFrhsgNYmGG
aJtgt9pRV3vnlWWIn/JVd0wei5iYWUOD+XgScMeYcPC9FM75wssVjFjSWo8mX4bo
nwbaJANNaowiOge+F8AkreZXB18hW765devPyd1PMr6o3y8+NJbAPpZfagV0/yDp
tY/eit31+91PYReByBYAAfySH8Reib2J8OQJH4jGwYMr+fs5IEB2T9e/FwuQZQ23
Ke9/j0ITlyhV+iNY+ZQc+6bCB9/S8bC1HrBd1aWh7KKi5yUHa0jf7nmUhlgrkYJR
RSpMKcWmzLHqxDzOYZ6prEyw/D41w4hlvlWqucSZQtH2XtIIAzxN3VDoqfOuo6BW
wmuF6j1hEoxkm9Tq9MBkxFry+RBlcOVkX1m1phf4obp9me/44BwXO1WIf+U1aoMB
fzfyldg6nZPuTvEeUYacAPaS6ImGYu542jlopZHhm9yW2GwsSGqiiXtqvBn+S/S+
gmhHAxBJaToXfsQqe6i0hl3KGHsQmpKlO4c2Np1jmvXscIO01P2tshdn9jBGmuUx
zvhnG0hZeXpt2rOeSOAzxgK4jCSQD4XiCAxxXdKVJw1lYoyEaCM6wR16VYGAEAlU
eBP1615pVSgRRsLbuo4SqwZKYK7yyb98xxa8k6aF8zvVAtTFPRSeeRfNLdaw/by7
PhJTo9bOZcmZVNjzmtKzUoyRgRqAGUMRkMDEnFwsabnlsUEmkzLUyhM1uS7f/pQ9
EkkqNR+dVwb0Z0my1eXj9M/MxoTLW4F157R/6CDUngmU6jI6HNoOnlLueuT2k6+J
MdStx2l1GDwDyt8TC7ZkPx/NOU7Wl07n7bbMRlwFA6RHOKpEvLEG8AezJ97NEUZM
iu2alwquDdavVLujmqgD/sDSeO++lesJhl3NQ7TTuUnPkETo3oUXvidHmIwALsRA
3PfqEZNNNwRnf+Jl6qjcFkELHXyt6lz4JzuFNIOHb/Dio+IHxSNXDgYOy50lr3QZ
Yfqaq431xqfJzEaNPRmIUfk2Zfvc0NjEuS79VgRoP1mOQCTEtz/+BlIvLU54hbth
YcOjI9BPnpmwrCpToOk7HWZb25xx+XHpTAuQf/oN049N8iSOqlfjg01CDrnaR5he
blmR2zquaH1vV2yRT+zaxKA/B3s3atKkbqHv5Mnu1oZooAOlxkSKgHpx0mBO945b
tl1/D1wYi7FREdvPKRq9WMSRq6Fh1hX67mW3vMmQTJOth4tbRgTnVr/GvF1IBSxk
nYJQW0mTLoHeolBWgwaCBbBiZUMBAb8WIPjE/zBpJJ5Z/fFfTPlD6GoeZMgENwWg
ZwdJlFbjJkSBjrgBEWDD6Ba2H2BW1+bHknxb8ooVqzrqNTgEa1+cxoJBwBJU5Mmv
H3U6c92cPHDFX53DmjARoLNiT65WSehmwYmeHX9tGBp5KVhF00ghFdg6hrT/4Z6Y
nBSft+Oyf+EfeuunyV529rieG/Gm3GRzhXaSuHiw12Xr9PIOquOmJB+YNNJ+mz2i
YwpgJTBWbhxWlMdW10kfi5NU7IAX6iDKNOMmnIxMoGY4jPkt8kYF/C2SBu9mgmDQ
bDS+c3h5Ydl/XQj7FRDb76mGnZhc4mPkXpVV/JaRWwfOBQCdwdnSFgbtCSGGMEQi
K7AZshF9eNziFBFfuyrIFzpgKyuq26MqEyoxIsd5bX3DBt/C85f/cHISx3fOCJFo
5fAshqoz9zMbyzIsRUO+UnnHCel5F7r2X3mOGliVxCaRY8Q5nsfFJSEzH5+x9ToX
2tyxmjvPOPtQOHNqCl1DYcB97KAozv9RdlOQYLM5jajl+Lr6vAAC6ajNd0IDsMIW
sKllXRGXi0SJP+TRHeVTCRmjo1eZRHtvUC0VNb0jd19FI3P536JS0PkE4TYa89HQ
KFa/aUlFi+lb+OtCaL4sxo4r9QgM6AzAF/qJBOsHFRC4o87DJJKMJ+pZ1fa9+4bw
88LscTz5Mc7Axht/cvjhMREW2ZcxO/prdK8MSh/PDc8xT/M/tuh+8sTZQdmXdJ3g
CEBGN5tFFL1qvOHlIh/cupfb8xTxkZByeSY0aAJVv451xsPwXD+4rm+7QT+GPjRA
BfgA/cxDcEtwx7fMxFB7wpDfyns2IWYcOCGfttjJOAew/aeCSQfL1fnAKgCiF4BH
K+lnnw95UiPHGI/GJRjfsGbagbQh9F6gR2Z1ooSFJEdRcme5o7v9pH7I2jIB06XG
6QjwvmGluzTJipOAoedz7IoweYkdBb7PLHdtw+p7AYKTwmtis5CJ8c+5RZWHyZFt
hosele5K+baM/U8On5jq2QkigVLYMB9Guyzfun/4dnTd0WIS3dk9FfcEyNCblg2H
yzm1P3Izs+Ex6wA4G77HKjkfRJ4xJg2G4NN1gy6ViFlull/qKdnH7D27mncffF5X
IO6l5nUKCkOGUlfhu5IWQ5CfXNAVHS7b3zOQU8xJkhlMjrMhheynFH1g58Z5ju4J
eulUiUlwM0FO/Ca6kWzsiRda7QR0G56R+ZKBN8Ns39MsNJ/HOgufR86/HQMxqSAB
V8ZSepyipUmTkWtCdK4qeA9w8/FgaiD1ztmK+WhrtaubA7hpt2qIGJfDWVbz8jAH
S31QOP9iGDp2mqZhkmP6ithfm/NtX5qWPg8PWG5j7JGK7BpIolQQiUwPRxvL4rhJ
iMwcYzv/62RzRflqKA3+7GmR8efhbv94UCnG8Heanlobaoqh6MM1EmTJUij1tA5P
0T8Z2hfZoif/udetU4n/Tu8NTCsJUqSAXmG71hBdA4N/SzCU0t9LQrKBWGPnGxIk
68UhqAzCsCncK1AJIkFTu8HfD+cMxog8nHmbHVSUN/2bwGoGpKwe7Nmt2IGs1+xu
7n6gjcdaAaJPpMH4wQu1+Sn9eAgJM3/R5f1brwKP4VToR0zqaFlah6d+OpvaI/yV
R1xlh9589bOsN5d0o8oAmoSbkkprE6jf+/4BxC9ZeCyqvPTSBaVCdLVRJctJc/ZZ
vFx0LVjwLXYMAsWJiv8ETz1nHMPd1H7krkHbtzLG5PIKQ/k1hy4J4N8mmSeEezrZ
cvf2DaGq3C0cMgIk2cJqfHPWAMPvDz8KWGaAmhr9FxBHY/x9GfHISHlu806KrP8z
AbYVHCpjk+9jbpdEkkBKRJeHXjSBqyBPsjyxRBlu7apsgL2tJ5NNzqawruCkwkZM
9Wf1mr0/F/Mxy5gdXQonQNBR0+uc1pIO31QBC9ApJh4WEBy5F90d6mEQjwMqDEli
KyXkWgNlitztRYTYKKC3VQSCHJPAFr5J0kB7cGvwHNUugkW2JWJdgCQ7hP9H9oMp
2u6T/hqi3WnlexaSPa6WtFGnzwXEchpRwQz/hFndDQnq9zg1ADN05/wycNglf79t
Wv8RfqklQVm3fHzhw6tYeJEVJcSVg6WsZ7Tjztdfo/ABFgqvN6jE4dT1MBaHmfLy
5+fymvl6Tp4Waum4p4Yd+DKrhOQBB7XXysE6rRMjpFW0+hANPn7m7B2JgWsxs7qE
aXyzL+kdhFTOLq3EAjmoyN427cBcWJQvUgEdz77C3YOUV6bbXcXaj7gZ0YabScRy
InphoayNOg7PMqQIeZYk4AUUYQkd017Bk5PbA2ZZTPG38oe+m5PlhSQuHBZTb3FT
jwy0mAwVn+e4elKBtm00JnrYX6njO5rDdWCHORER9u/MQ9V+ylK7YhvFL8ZQTqfz
rRRpGCTo4lsDm7lM5FFqIpxuhpyjtOYd5Gkkn1AJeRMpTkUZLTeIN0TlHZZzIRv+
sPWT/2PX3ANFtDt6/IwyQDyCQBYKZLuOVzSoJRx2HJfScNIHevyW+ggxKTL14bdX
7WZ+hB/IaVYUOOSTrXi/vwUcpKGxZFdsOShcvNpuDc6el9UjPDi8zCd135Qa9HfQ
Hfx5Nq5Yfb6iMEK/N0dPWOocHOIDfSVGZxFVZiIh0sKtsGehS96xeROSTeTl2FI2
wSE1TuY6Yq+WmPjMLCN7jQGPP+a9Hat9Jzhm1eQ5UWU4+y+5M6hIDZk8UtuGSwUM
lM0Ck2FhXRIBdQ9lijKgiQnD+Eo87Mq4Yqx6Y9kyPyMFKRlDSa3M/8FXvhhObuSq
BLrMVaHT6DX8bP3Cnv6slP2SXdSiNB7kbvdDwpdxSvdo1DnU7kJB5MVKXzAsGb5S
/ycxlRvgzSN8nTbDHQHo477sS87C1BEzYFKey2xy1ZF6HI1WQDNJRJ8xvhkJ54dK
+UNCJhmHJe4ccjfvTHSm6mn0OQhlO4iQnKUu8rNsIkjasgjZUej70bbc+raEgggD
hGOUyU40zwLUaQUpA4+MhSYtAetOWtr97KwegyCRudHsQ+PVGJIGjl2mzkfHNV3V
y3/LzbtTcQf/MPx3bkOZ5ENrqZWbD2S55u1CPlttlu6TmNAkx2MKXjtvyI6vzRXJ
WwmaoXGwiNccOY/KQ/0UlCTtyiF8vydPpbnhrqCRLTke58LdSfd22YeE10bSUWpu
vVPsOJQmH8uHcvOJSeCQgSBT+nOY5vjMgDJ+AyngRO6pBYgPqhsE7DAmJZTkB7hj
cs+/yd4bEuCy2s4oXqanUIu+cXrCRi0FwKr0Ok3nf4UDQbZKEC3kAxbdZHmO+Xry
DMtkkPt0+2/cNf2YhpNfxp61ea12y8wc0Zg6ZBuuBrdlxMpsR19BgS5UgdEdQQyO
71EXiM92TJaeir6DDzkLyH+gpdn/ykpKK+azZPbY1HvfXZYyMWd9hesXm0XHkDo3
cFCAOhbuqqT9qqw9b+LtDaMAGcz/XJIDzl6iBM4UlADTwBoFLjUqtD41MtlfDb1q
/mdENJ1pwDMuGTMkq1Uvzeol1QYN9l6PzqaOH/eSp7EkrQe7HUALcDWJTPGFmSXm
3WbdJO6HFATp/Yf9fPHVTeQrbsocC4BbtNtO4q+UFSwpmMgFna3RpP78dtj6KAbU
5Q6ME+khVlf8iKIRncTFZIVk1+DxntuhvrjDs5+M3Su2nyGN29VdHGRjJDjwO5Oz
DoSrfsotqjPoTKMGQLgl8eTIPB3So6FY+E9PXUVs5/hZAnf3CUjOtc+VBo4hDOr3
y6a/Y2RDUtxrrz83xuRMf6LcM3cBAY//MM3wlZxZ1ZdRKIcwD/rwyLWq5I5itYWl
ZhELhI6r1OMJIMK8YbkJRntWwNkgeTyt7x1vjFV2PbC2/cycL2UIDVbARmIlsafE
vjUnO4rziscgkb50IlgYGjj1x3iB0dON6VpXW4DdjtOPKtUFFpDGlAkOvPItO49c
ZxGElM7UJVamHek4VKJj0XhoRWtDZhS2T9o15eQHI6cly/LLbO0i9Jxu7xrESsP6
aDL2Z67mEMhEWeG3wwoDPbunn8Q5jItlbWJ9Mpr66kx3sHNuBxQX67uZDORTY742
tLFh8wHBS3DvOFKiXsv9RU0YbfSTmcglpns9smDcG9o0WrP4ptlSPOg3gYjWK6Rh
Z3G/LsJOQtLUOmvHK1X95sOXDsCMTzr44tyhGMXp7S5wFfxfK555gDhUJbAbvAB+
gc75OWz50aWB8fi2k0xf/5ev28ap+4BkYiPHgDrDydKy56IGYpvIrkbXwNIx1faf
kglFOlUkeI3bQZxp5f4h93bXgSisFkGSKYnGvrxV6zuJxfAYZcmZnsmf9U6OboJ1
M8PCZhqt0nx9yFd08WS/2BM7VAmgl6DwIkr9wEuQgU7pRKTLHbHvLMHv0tKuKL2r
mdpmbHp1KyriYmib4TPt3RPXTKAMBgv1X6rmwPA1GyEsIFlrPg4MP/o8qlQjnBlV
Y2wt3G2MJOYBnRjJY9It+h5osZNVvceXWILykE6nDEei6ObmpUKqPfvwlua8tcct
d8QXnGc5VqZtwToIID98ZT2pjvAgfxpKWseT+ACajXfdo4x92/0wIZ9VNwCk69Cn
hIU2wmZIaZY5AzOTgY+Q8gYqoGd/o/Wo2tLMrsCKuuoWTtUz6t1+6rkMXm/ezvap
ITNKg09VL5c9K+zfq4kk4ae8o1fEySqb6XrYUVuM5F3WMpO/TOfp1H1Lb2wqFbR3
SgTU+52FXtVut3IrQsQ4UHHrVt6GIPv0VwYCgcWz7k27Pur1cuKyggBtb5rFmiGn
aF6vle8Bq2izH7l3Q3AV89yDni/93mQfsVZxTSQWVU8UrSKwQDPdwNC4+oZT57JU
EBtG+kGJUcfhWGMDlBS5OhjTO+ruKRTbtKrj5UKL3pB5DL6Kc56bxNGsaweGVSUq
kO7Spcg/vRq2NO6GfGbcYlCAlrim20OG8fzCL1b7M1bX+qPSgjp5RvSBUjlbbRQT
8Eb8MnCi0D3O2rdN1xAd26+eGCo1q2l/dqjbAnVo6ZsJ8HHQjRKTS148gXDHxUJ+
SSuVC0pz0exwISuYnTDC+10YSn3UdUf29ah4vAchF0+tUQRQv0+/PWpxtcO/ZudB
s1yNdrDHa8s39culF0Aw1PMdiI06WdxWjtFYjCvFY7WdSAXuSq7hQdeNqqePXbe5
a9IwHD10z3ZmbV1bp9rwGFh4QKl+bUyA4EJWCL7ZjU5JuPUEgRntxaEC2P710rY4
QWppLUfOAqBjcUFtR0DMT6774uZ0RHSkC3462K9t2nvrGEJHEppIsIIAChSgfzje
Oc935CuX6ZjabShv4HYxTEpPiNnqQ6JGppuG6s7K1rdWCZ3X789H//w63+/FEtlm
U1nl7CiqE5IMUIMfzTfHyXMQM9fuuGbPiq1hxtx86hMqljGCw1BS7FMa3KMCpBTb
m0jXG4WnTcoykUFNevD0Q69OpYr7mfaii+kCsj3ZwV48x/o9lfUQaA/A5pLenXT8
HDyT9htxijM+iDqUDKjLbqs7FlwCE9hixrUKZpNfjpBUhDeqM9oIxCOgtIUHXE9A
20YYHoWnIIwcJWsShvIxacvleN0N4vC7kYv9BG3ZBc3uyz9TWR3nrn1Lymbo1k1V
HbYwhmDNlSpTBbYoPPNuZ1s+oqlE2XGevqEIDjq5OJwhk8UqxFqc604rC+NwTHXB
KsRmzAEwk8pO3/yholljeTDLz4UQLMiqyT4eadf6jwkaJh89RgbIAcgfSHDvEvOs
yVDvw5ZnJYJ/vZcvSN4wjY+8Kj7q3g6vWQh43AZEzU0U8sS1/IFbyJDyI9pjEuTp
5grVVxpAXFSQhCE3k8AY50uFcKfmzvOhmcYbdbQ15QRfxgz9aIjIlCSy7VhO6rit
HqSRScXXEDgx0lMkVnlu9lRQOFknD0wJVr0TjgavI6RAwl4XEu5rH9LJRQMjn9+x
mdlAYec0eTP6dPASDuPACz/iROQX7hTGZu42fuPxOpdVThKXjbFcRyiopSmexbK8
n8Fwjp9Y2lrL4yy/K1yxITqOoUtL10z+QuOplpU11DItBvVJxBfp+2ETUj7PDFgE
0CnnIn1Aiz+MxRX6cQZvTnKaUwewCo0aGEMh+IWefcUesOHB951SynQ9x51Bbro8
hIP1bw48k2CoKXeffy/XJNqxsOzqW5PRTyAB9vl9UfPTl1BjfYkzuy/8+c0got48
Ws5i41Lpi2MH5SHDEasttmUpDkCtT2yryhTolekJWJeA15+6Lk2r3MxzP0aILxke
HhgQiK/tgsGhepnp2nm2zPsl7u5St1S6cQLJs0baPRvE1wGcuxUPHKnpNGlvs+nE
LA1HtjW3mc1hAz0TLs/ak3wU9UjPBE1gt05xLWvin9iMHTIa+gTN9bRil3wKUsAN
g1nAj2VfeI3njhFlEkTl4H7BNLQLzaBVcDTO1y2yPAt5y2X2U8T4mlrNOO3g/MIm
sw4D4GgadZTS03K/3jvbd7ukh7EF0ljAlanJ/w+WAFDSkm23pgOvGBsVRC1G+BZG
0ofzHGpNueaM7ZSRrrMTkxMtSa48UGTq1eeHXrHJZKSTcoMLrFNeH+l5I8n/0mC2
0NNQXVHbBGaO0aPcCdJNhB8iU8DL/aGQbdOHeVaoEZqGyYgpYqJX1UcJOB6Srm2M
ABCtRMfneuZ0+7yeRLYv1TwiBRN5wwiOFlMkW9x4iWwrcuNpf7qTMRiRaQcjwxhc
HCUmXhQ/8PfYjyP7Vxbh3kwRtavDfCJN5Sn1dzrD6ZUOjW6AnE1JnKqJlM+/Aqg9
/K6UBQZzfQTBRiTO8vhu4VwnqqCqCsQEB6h9WVWXSdPtxrbmFgUI9TdVNRmiA+ac
vU0Uw/poZheNXGIb9x4XQvuooiSyzRhcV4E80sW0vw5Dpsu/hq2wILMMkus4SL0Y
sP1Y6Gd7EMjXcIQKTeEP+lwoM8X/0ElwuNSozvmJSCJlfhWTPXBNEHXigTFK6+Cw
PTpVo4/d6DIunb55ty+QF+I36HgJRysbEQz4vVEEVgu2eXuTYDe1ZnBtqYoE2RZj
GCY9akgKJ3LmRjeHyW5W6SDzJGu30AKrakH4CJWDPbFlVaGgh+dLBGC6goCMNuod
3gSHI5HsCuuoMfLEiET7QookRvLbArSnjcT9tIb907v58VVqfr9NS9SB2t4MSQMh
Svht0wy4UAPLNCUbX23+FuPYUR6ry07wxJOCN6JdoUTqsUpsdyvtLkKa5kiU+EA1
i0GW/gafWhZRD3GIfm99zSPCgZP/lq5fxJ9mvlVHgFxERGlP4GcX2WhCnnbI0dYC
4rgKPuqTOZULHoWXfOmzAUa7UjzWqLBetefZutp6UmJyTUlN9x/Nxl7vXpzmAaB0
nkxwVY6rTH3OM20D7Pg/MtL0EuyG6m+rczNukmdXGvw14delRn4rOVH1qaHjuOaX
FUZ/fzV3DGJSQMBO3Rmjr3sSAmS1ips/6KPJcYsmCgFsbUADcoBzBLZTWC76nJFO
/Za4ArTGiRGgiSXsyz+Hp+1nYIxnhFDmoeacHPvediT4JNMBKGAJtYVIFxp70qSA
OuX5O54NBdJ+DFoUxSDiWI4aBn1jTWPvDJXezZ3itW4TdjRm+iKAzH8sHzd3QBij
MSrIgDuqYBap3Bcpq65cVjCj/zfA+dcrLLZpDQGCjgzYkV/SsdVrMKmuRgXFk6xQ
ng07WA0VUhwVrUq56xaQwq6Z0JtOrD/Mt0Ptc99lCDcJPcbRqKzMSt+PjZc8RRAd
H1lDlpOsEm1s90rJLVCC7qawmN64vWtWBqnWxgQxqAmZKl+8nOXCIuGMHWYc/t9q
X4Tsoac2ZDJ013BC5nhS7d4JjyLmmQyUU37kVhvSEVRHOquEHfM1wfU9OMWuycK4
oQXvLLbU0BBR7avL3SHVhKaIMOsJUoXCHy8sv1mwaDrhsKGnnY70hLIb7/anHqcA
Vmn8PEv5sw9HmEZJ6l05GuH3qz5obc6MMaoUOCr+FXCUJ/D98a1rU9dWTiBF3Ax6
hY4OT135KTESQ4eNjYgUbCCIyQA4SEGDK4tc6xczboE/jM5wdwpaZ1rsOO/8YB0O
F3McmMUAtq47owCSLNLtgvcVDxx9M4I/EBngTgTYYWIgq2nRUQvJbtElXk749HO2
rx0QUrxjXxpJDKip/RG14K6s0rUlMmlzxdEi9VhCdT4NQ5thYaQQSyHXBGHUKHyy
W1uL/nTE+A0z+zSCNAT2WrQVJMZseiZCjBbll39snEoLlZjz8nGUXhIdWOhd4i8e
ucbuBELyF0PQ0vIoHdf2KO6qHI3SCbe6mS4o29fiha7j2zx97li/6f4dgC74wqTZ
gg4QT9qUK4kP5Z80UWEMOJ2Qs7NaZfyUghxJ78itN7X/J94UHWvIDUeyc9+hfbWa
lS2/oI8DNeMnUFntvpsCujlbi29vx2xjhoJr+mLriZ6oOjA4f+NYVT4xFYPdLuCH
n9URBNW3iiwmyjU5TrGcw5U7NzWxS4fFvbqcvTKqg94M6mloNdweGvcMm8w0rs0y
rpsSL7MimjmlD2lqByObxa3vNvhcCNFNB9J/NX/SN/8wkc8nmlNcdv6TuIO6tPF6
XKulFnSqudjXRxD2+iqWhr1355744JCoLPS4SF3gQ4v4rOvw4Otc27V8fPYiE8In
35bNFygovJRBFO18lX19tqCTfbyWX09NR7jyjIRbWFDZ2RXg5xjVUDKhKRvCVQkL
PM6wCuiH/+q46GoumLerYelMuRySAK3+oimE+Bic/lrAj3PApY7drfT3JgXQWhHh
N1pvShWp48JxiKfBEOjCnc3zVh9Oc1xtkHi/IwrKmZUmSnnu80kVhm2vPOR4QfAo
gWnLGazUxAcvWiLloTH+6O0vr2jheWYTNf5A3pL9eAHDwsqBIRxeYOBsPo9rVR5b
IqiNb0lIkI5gZ+59s0Dd2p48gRbmmEkma7aGqCUv1tUYUPWkRuRrP9HtvBGUJ+yZ
m8PgZvvoL2nyn8E24rGxR6olTEGcWSre1gPPNkskvke8IlatMClCysXOghQtW701
gAGv+PkW9rhcaZymt5LXXL9hOAqKqi76sjAunshx8ftZf0neT1/WHTEeoXuNkU70
GNEYcuCBJYHeYOdF/jLbp7M8it7mYKBVe3bBLXlSodGPqW1vqdf4QoBuogQ5Frpq
CgleC4pmaMB7eSbgmJ94FOH3l4nx6ScPQimBFAJIYKBkNgO7aYYxn85i76LrSKIZ
nGW99/EEx02wIj7MhUb/zXbk1+Xg8nMo+yahidRO0FHxi3XoL3JlJErGJJmBRyaw
C7nPlFvZ5isvg4sON2AFswWmE4eeueZPFlysxV4Iw90kEk3fqjk2xjV2hRWC91Yr
7pF9auGj2CXBUhPfvyJaN7nHIYvC4e+vS3DDfKZw233HcGj3LDhi0GTXuYNuY5rC
98gczw+g1+p9AqK/YEFreUL0Rhl8d7tEcyCfi4QYxG0ErpUbA7Eup/kjcrL96tWc
d2+C4p/Yve97/huNJrslDLHEyGpF/nHqfDvBtntd20Yk7XLNq4/dIs405GiJpZOz
9vr1Tcgc216ZG7ZDatz6mjgewa+Ddnef9WWmi4eIRpqjINFa1ewbPgIqqCwL/JHs
XVhKw2PRXA5ppNHfW1+QKH3EHyAO7vH2RiBG7zN6v9GXuwGXkezKLI2QJq1VozX1
Hdd9NHznd09oTgurBjrkrvjXYybFjyVwBqLSrf42ngYS4hwwpW8kwtol+tQXXVq2
BH4jS1cg2QLigrGmO5NEvI+BKxNdWG7bP1KIoBfQ8T+LkvLz12ctBj1soEQUYSFe
jJV+0hd9z/JXlC69TSebQKCKN/lI2YMfBE6gBgPTLJM6Ji79fa025ioqPl+6erEK
O1RBfIGJap5WtHIUmSVQOa8R274hjEub7wFL3NfdgxA4DzuuIc6rcmmuUZ92NQ5+
TDyjPUyzo9t0TgWZbYYGpIDPmDLvWP+XdoS+hd0/YzKsFEX3M84qbDg1QTXJh+vO
2CUWYRWxm/lOR56yCVAGOWbHIhXnWKS8p+ebt4P87ay3LUfjBy51TztodkKiwUJ0
V8vMtyg/74oMaXVVrqPZomIrBqfKNLZpmzd6W7AlSsU6PsRucbW/nmWEsBmAi85b
FJMK36Vwv5lOOliUUv1qhaoEjjWfKzDlggiCTKc++fOiiAuIGm4QD5pWaYHjJvC3
eW+4gJbg44MQ5g7sDOdCVa0CNWuEuvB5IttrBvbxv9SjedhqExl8cXd0qs0ZSLGt
14qG7X+z2BJf5FsOFu4tQvyNTpVnliGXmJiKHfmulPgg+8Bt3EsdO6MviXnT1GoN
+pW2hdGCiNvRFzozZS7qSB+fgK2mG89G97CN2s2n3M50ltA5HhyP6xYGVOKVczah
1gpqhnRXUW9WIt4aqsTyySb3Dv/1GK539jC2YvSAt0oK+ze7h/huec3XfBblbLKS
XaIvk9OYHPvTkWQhmOuFTMCJQyUBtHk/FgiDoe9XqTGmeNAbHPxdLhC8b2mQzPzl
UhqNIpL6+6fheA2Bbc+L6dvEB8GM37Q3VAGEKKO8Mc0zh1B0t7GbLNy+KCo4LSfn
u7iE+NQeNPm9jPEbXKYYaqvKpotR6m65QsDvJVarv6AJ82ozOrPwXfk5FzbkV0HF
5Q/9aa7+DZg/ZrHWhm95gOil9VYaDwE7T2iHy2kyqkwNxFftHqTFZNgxKHvAnf9S
FhjUuisWSgoQJRDQiX+ZPJ3FkFzAvPGor25hZbLB6kKvC3yZcjBsHUcmKh7leqwf
LVdmxotwuavQ8QMrkpHJ2Ih8ItIkcnyqbfx3dlqKpbmDMZVpsM3YL2007dMiLSwU
8J6eFmCmdTr7mEhxwQ2RN/aeRr7a+cxXE5OYuJmlCL92Plcc5ciKtIR5wngwqHj0
rSqPrWFkWtoio54wNU8H+5J2SkVBnNl2sGPUBwFG0+QFEfwHg6qA985vR3+v1eh+
jwZOaZXYIb5dxqcPV90uYE4gjjDfbYRbOJUHGsQuHvPyJmkvtb3XZDBPj/ZJsGRq
tnlm2qjDWaiXIzDpZRZycj7zB/T/Oy5RKGk6i6e3N6oZ47R3/hfXKDo/6GCi3c/W
GB3M+ywRLcexNrS1aJlB7qGhS0AB8YZO+Msd7pnrurlMYwlD0f8HZcu9kKs2V9j1
ijCbfMY5e0P4vKZdv9DoOOhWXtL13jtJEp1y3kozpfXpRk0YJdgpk/BgMKbfgRxA
wuHyJVqDOrJxy2k8EOMGbLFehXoUAVHKfsd2JHX23HhXiLy8d7JDKXkGXujwBNyo
TSf8MtnU3qKpTQpikKTynxOiGMHPwJwsn0TrWQkHmNH6Xpurx2u1hUc0thGZe25w
RGnzYKHZnFh/2zNnBhTziy4IVnVol/9T84esNmdZaQxI74FYgtMBW6HbKqLp2nkZ
RtTt5XjEXV02d527HrC4tQQwoyV9HM5UZM3XC+WevhSleHegHNPPrhKvsijLP2iW
Nyn43JvsHtbQtnPbFWzeWYmv0tpUdV3voYFvT5Gocdb4GEiLwCbj2qxZv9EtTd0N
/3p8V7Kr4D6FTlPQcWA9P2vqM1Yl/NjtCudwHmc69j8m28l5U7lUO1Ea2ql5PjZ2
IrSR6dA79S0zOt1PSEpZfYqEDfiUCX+bnsypG+fBIA8+Y8Fuo4C/EZSJWbok3M4r
8u+oi7xE/cbCEk4XU0O5fqXY3hj8ZiPVV52Th6lDr6NrcQros1gOqCddhZfwzBbB
e49znmUtsmP3Ogxm40psOY7LjwqcQo5nsKyVSJ03GqHKSO9hteEp26ndi2lUowJU
v5up0Mr2DrqkIV/PAlKBQs48O4xTRR1vHmNm17gn+TINV5AlqZyDwCbkZDG1RQkO
Biw/VJoDNxTHeaIstQVuMJAQtBAlp0AyK/7F4x6/hMP1EQP5ife86WDWaMSzvJlZ
HVrUnsY5dZnJ01cP/3/5ATFTqAzeBcVi+72+OpD5EwfcGOjq/2pKXxCl75U7BHph
I9MfNFlH5fAE0e2EPKEyRAf1sOwyQMKrX96RLkrA2/o4IBdASbIsvw6XsaEIz5QU
giFWFyOV+hd+Xp0sSqZjoHE21azOicAWnEjQWlq8Dup6bzDXDP23QZLbX4DEXIj/
Qb2EQWOTiKcHc0ygWJ7hc9UUibiU/yUzpAB1GiLwIpBJJ61sTJCqTX/46dM/aLMh
d7mGeu71p4VfACQtUs4e/OkqVGCgpOStYOKM3a9nuPfqAZhK9bydGsiHR2xeGuzR
4F2Ve3dzN/qM95nlOrldMwPEiGDTOcIFz8CqszcwYf+h6LE97F1x4rm+fq92Eal0
yMJDQkotHBTDXzLtdQEbcXwGZhPOHOnzsDPhVXyW/uwNBZguhXKYby3EB5IF8l33
UtMhJK49S0LII0h2PwXYvkL1EdSxitV4jos4JiNfBNm8Re2RZUbzhAqSTjzL5Gzq
X6d2u+/mEqIflNocPQwSlNeCzPxy9FSFEyR2jDQ/P/HSjKep5UQdfaiDQdiTpkhg
lL3Hn1hGe2HCRKfKj1RBk6Ow2PnIhFScGD8b0LIaY/FHa9pM3bmDJUKB+iZVigZx
b1YWCupceXVd5DpTt6g0D7X7kzklRURejUNeGoDnaHf4U33UMQDEft6UzIYe17Lq
aT6fcRtocW0hmBGEHpuk5oE1HqA5fyi5XgXHyO+NG61e4Q3nvKRutZ/SqKQQwD/+
uSdrmPNyyIHIJTAV6y8FoYh+Zmypurwg9y8yQQ77CxDUFyEchyYiWXe/A3kjeygp
Dz2F1WO2K3SKdWfpGAbo+lVg9phmfYh6oIexHm9wCuOUD5nyZkob+go4sgQJrwZS
NldIDhlSK9xizUaJuc5T4EDebSsMJcju2LJv53DPI7lrgB9Rw9ERN+H2L2glMj0r
kmDvhNjn6EYyszZBOZQaz08uHuYbOl7IvSrweBNkC/dBWxM4nQNQsnJdotEblckQ
4UUlQT7Iue9TOfGfk2x1vHNJ0xjWe71UhzhD62a7hglhVTYlMLILxdPwi9U7Di2G
DISzeSiiCp/0DeiMi+i0P7sW3iDc6cS7xnUhijDCwM3OU+v1uRDmgu5vUOmdCnX5
fTkXotLu/PN8ZkzTv4NgVlopwBmJ96dYgJJE7Ta5YvVvM59P1G2PbEk08Mf4TJHz
7R++6Or9UQa80BYJpLiUWbK2ysc40nMKCldiI/9Spj+te5t2glPl4F9jky/DdLQI
w4O4rj+iKv4XFriYkU/el21N9usHAf/dyAKk3XdyZ9hK3Yof/Xl6dboIp7tyy7bM
gLYVDXWnjVOvwlNoWO4spz7F6KdXtUGtvkQv9X7TSU2XxT3MAdCmIrBp9SjBj906
ezO7AX0hJH7vyCp+yXHUa0XkmP3gvNm6ancGlC9upmJjMBXhNv8cNEw9sXYAmgBC
RjcoIOjnEJwGsI6pZgOHIGxlBhW7ey7Bpv769RKtPxnTqmo4911kyW2FzrAeHyU5
T207gRl8/kMJIs8xx+sFdn3IBBVUuQznd3UsIMu8908i12NRaXtCeg8Up3lDAbCK
veKFdBcCP68uBSGNTnTqsqie009gx9cwv2u/i0lKffqit1fAKfH3sVQMmRfVt2lm
ouIcvFz7jEZZb3X5fArx+YnEjsbeECraiEMao7txX5sy/2wUKWnBoJwlTf8ns84u
HIq5890frPlh73r/NvPeXtDt6MrQdHQuiDRMINHSX5pHle1mnm3/D574TEO/km3Q
PXyvlu9JxqYCZSRp56V6Tkj6Vvu7MSEPRvk+Ya8skhpW2asLWFY79vRmleenJOcS
Oz2Mxu3u7hDqdaM8af64GHM7J9xUGR1Vt6zmlL0PqOvFiXr55rYrTEg0cgAa50Rh
ZXJpUYmGRcR9riSOwp7pEh7GmUBEoBk44VaohmK51Vfd8JPBY34ZvcRnrWFKib0q
MMZBSqjj1vHg04bUC1Dvy2diOG8u4FuNYHi309bwAtSfiba9ZfUG7z5P69kvFkJx
EJP/f5mZuGrRyttV+mSlcuYF2R/m01tS0u63ABrmQhfgan8jZ3y6f0AnK27JKOZE
ltg7K0RpzJY4v5ioU6lC+Qy/zW2eCetvM0JIaRZFEF8x1C9tmIpXwfSOS1pQJk8r
XYsNvqOhrEMrqnc5t6ttR36uJrErUY0UGnje3Rt96YFwVT3pN9xZPTqlysYpygbz
nT+U2JYHvD9WP9K9j18gi2YEkhq7eZHu7Tk6zlsVk5IQwkazZaCX5OAEm++yygZe
fpuSOBGzaJfJxWOrC+wBLRNWjC1iJuRgzMeOw10FwduoBYT9F2NqTuH9KObpNlzE
YdedGRJoDiJnXMjKZ7Aqrr6tK1Azf7pYbh2iXcdB/i06D8D3UmK1q+F6w/2zSBdi
ChztB/g+sWFneRcqgnR0Tc/eDKPrWDpcvdqh7xtpbJW53WETjgOeEdf0ph4jamDG
rV0X+RgqZOYJ4dZP8eOUV9MqrvLvKwKGxOCqMyFUSgW/KS+aNCyD45auP55Qx3m0
SEuiS9gslz3m/7s80PGuX7pF5RWpgkIMUppbXCShWqHG15Wp9H96Ix000L8vvYzD
I77DLp9F1HB1KIvTo72iaMtUBKL1aiKuPNrDLh004l1wQdjz6x2T+RA5bMT1Q+J+
J4QzRbpVliVdVDeTyjanUEaw6m2QU8UaiZe0xq2EEOAbxGj72l9DpGY54hsIJEx3
wJ64T50JIF8zZTnX9NBmX/yfbE7SXWIq3jfUXisJOPkdN3JwwKvI6FdgZuKJfM89
RHniqWoLfelg/0F3cLbPyRQgZuMIUW8JO0Ldv8pn1WXUFl+pxh4y7Q3BODuYSTRT
mlQc3CoCbtTfrJGOZ4kPAjWzfilbpLNLGrf8QLpgx0puNDS6qknyY0Ocx6gLDRzg
gbInpMwiMfCLe+ltdLnD9CBJQ3pvRyxk1BeFfxJRWidJMUvRqXVMLAsQYZGm/mkD
JMvYPfvou+eqva6uMcwLydKrULZfxMgg4x/QUKdqZONGEzvWFdFLJZaL21nca4So
//nDR+RcDYVAgBAH3xluaSU4jCMsOlZlH9YUn2FSb+E30rFKv+izmGXHK37u2oPR
oT1B1DAEUuY9XYtJt+UMUDQWjCfMzkGQvxMQlOJRBHwnz/eD65e951KR9TBpQrHP
LMP3HhEb7c1uwS6nB192QDRtjeuNvzXDD3YBYEMwiWLED0FYkvHiLvWTyJa9UcuW
xJE6gzOKcoSye9cFmR5aFifO6q39W7+a6F5pAoK9NirrwrZ60mywpPJ9IET5PEGo
5DXot3fnQwd5nDbyH2Rh8rTlg9pmuHdGvUX5Gkgx/citcrKSc6mn+QAOaqeNJCXm
9leKPMuZb882SrR921Mpl2HA5eFWJKkKkCEY6KUWMh9T2R6ym9ZCEg5YJKzl0c0V
PBvY8RCXKTFJ0xIqLj6/TGJHQQ4+wwQzSsh0y03Z45N2rLMrbqSI3FftcJbUr028
+gzAZq3k/ZcpbD6kV1px3TnMuwKKhWalFWfn4Kj7qJrGyMaqmFmlujv6lyZKgQd6
BlwhrtFAF/Z9EH+XUCiGBDodVKi63Cr1BIYVFw5n/coIGdGxs2azMM8+AHrQElZj
ZIkOH19umaGSVJMAnGTDsovLQbok6ITHGiKaM+yoGb1Tvw7hK3DeM7m1iBGeEIJP
fs7I8lbpdUshbWWvVOgTd7QmPCfIzi/I10xbCNgXcD1xL9LkXASxHcmUj22Xvcsl
uePwxEztl0y60Je6CT8i4owdROGj7JNhIPoc75SEbrvM8avXBh9NRdbeqKumwnJ0
D6RE/Vj8ERxcSEJtcrqUd9uC2QJMLvOL9JdvpXDVHtTssKGKE5fW/9Jvg/r++txt
ZwFoxp7wEQ7FXSHiJBA0Cthw2GKa/dZBEd2NbRtQ1k+6o7Wyf6DTNwRSwfmcNloV
Himg1TIGXiQ3TcGA7/EIta9V2o2rOz4F9Z1BMoQ1gIlZAkGtJXulYR4oXRfjdybU
mB/2BYWFjVRPp86v99DOWads2lOygRg6KXvkDlgaeRr5CaM5sZOjPGjpSy9Q3TQc
a+UzkwPFb4fuYR1RbodGSK5B+YyIRl+t14Jwb4vXBNtTx4EIIoNp8YIyLDJWrEuj
lr4Zq1CCk4c1g3cqCSKOco6e3/JDeIN4gITKzkO60KcQaimHIl+OfsrE+OOc/PnG
dwKuKI2v6WI99IYH8fm7QRkho8WBuzcx1QVQtTy6beVpnsCvrjEgzVD9wBoK0kIw
8AFO5xDYPNTP8dUAa+2WIMYLRekPab7oELzIE4O6Ya11DrRoeKlrTZVnZZ/PpIpH
znWZV1FBPFjO1nIa8Y2JwE1IRo27MIeDkGyQ5QhtC3E05AbDGCgsd8E0jEDPHZXm
qYqxz7IUWQiUoQ3Ogg+yZlfW5o5DaHWdrS9vhPbi+KB87Et4t7BBZ8eq2GEkUYvO
DNSySro3HGUjklQ9OBMtrDvlZKzeZcQJRgz90bnk8D2999BI9rV+NW2VWNG/xPf2
vThSSzXQA0btkaD7YqubWEtL0t3U1U1hZT/B6/frtG6Nfyg02wEfjEfWfGMbxo+o
Ebicc4FAB/BIAVp5CvA+rFINrLPmx9dSaZ/nCdXXcGVUjfAbivu1euDKuEByl9Eg
tmmZXuXe6BC0Skk3rFos7ajPrn0IO4e/b1/EOuZLJ4OohkRnKwFVYrXRrP4qBTxl
BPxNLv35CnhWbEFpoQLnZQhIZ5V7IWlHJKkvXPtc6TJ2hEWGoJT+urgPe5vulkqb
ucGqIpvPswMcJvWWVv/hyWG4atc2q5Hlf8Wtr+ryv7CS1Z/DQolIMOrPSoXkhoad
vWfzNed7frlsO+IG9ZOzyQSdHzCYgvr3NVT8qW3cAza8Xx7G1IXKAhgpvi8qnOKF
KRm64uhx1nCyA7d+Uk2VbhW+ceQEAcm8lEf7eCljSw2zlBESwtrkppdGVrUZF64D
MKmkqSfxcFOQqJrvXFQxKCKa9TQ1T9U6NEEAPhRV2QJbe/O0il7Lam5lHkFnAB7Z
uco7++iJm7ACn1Rf2Imv7tNqy/MXJGr5x56yWyu1EPjlj6bBhWs9KNp7+f0IuY55
X0/Hm6yQjOXm3pzVX3JlJXwy9An5Ckpm/hvZgxZz+8T9yhOpjuuWbkF0ZcML5awL
G+lPLQXWdRYWq7Wf1op2TdiDxnZxwwnrWTXQY6UQPN+t+jUVJCifngwKb/RRFPKa
2kyR0DJ0nvSJpULpRX52sOfUKFpG83JUlfBFYaiXgRMw6UE4YdcmpKWxUCmGixqx
Y8fEwCVD3L38UdxKyx7Iaf5sfnHUZWiIiFAAF0eh2nWzxhllIz73cUdn0Oe97R1I
+WGpFPtnm217f3iHEtKk4ry1eJO/0hzzmqYLMCJPqsunkrAV/VuAtMYTGoa8euzu
BIBEDOzEn5vI/Gm2KleUCK76eSf5S3hUMEXesaC0k43gyiwHEfzOz0lTCMWMqm0v
xu6icBcRsj9LWgecXVCo0BK+Fc3OfJcohf0OajByJmMW9ZTT5k7QGITMhMt8IrRB
QrQkr9bhxOe90fDon21Kq981nMkYhemsNTsshLxoXsMdKDBBddT7WNfjid34N1jA
yrLG0rglPqPT/h0tB4T/38Pjdm9KIg36G6Oth2Z9EdjLDE/kVsTW9SubT2rtRjQD
Pp5B25QRqP8ESuAvqI4UcVoNgwDQBCXhjs5YwTsPpCvnP3JGOYNiSxnX7KTZGON7
WTzAX4RR4qGU1uwci5ITzIks/5F3n4QG/dxqEsfpz9OjchBJzLK4w6IUnGEC3E0I
aqX8PJ1zMuqzbbh386VVBNuhmWfiaL7+nCIKKRUGZB2gi3Z3ctIX3WDLQ7DLGqoq
aQtp9uXCB17WadLWy9CxRNhs/ub+IG19WapJRUrNJ5qM8WdOqZmwb80HIl40i3+s
opCSeM8CQON8yjQLatPOgWbRoNtMAYM3k0mrOOUgS1MzlukD0J2hzGUFCwwKwlvh
jjRA99vDe5r6K5AaDsFe6tsG5d8gb0cpYvwUBOe3UUzrelVyrz8jaQY9tQ61Nw+Z
hjM/gMFuFlhB1aH7keIWvJkZq7GKY7DeoVlHuC9LpWZVjeJkuLBSc+r5cylFgx8l
5DfPPEq/ufP8crpkZOT1T2tV9eW4wUO2tqapnSbwpDCnGExyVZlmT3HvCbvS4XAG
+3pLsPiYTGAO1qjHnQxO6VyimHpue2wUloKgXnJGlYdCXhaPVSaf+hpyvtccj/v8
fkamalTh8Vouq4qfAamGhUeFn6nDKIAIv1y3eJmZwPR6Rh7ipNQnnnpLXUHYabja
mjRICNc21qrzJb5a3qL3f6Y8xPJ2iyfGSpdymi+mOgw6a8MX96p1lYzA74w+AXPO
d7p/jU23zPo+cZfKLwQC9WPlAvNNTOOhPZ7FEKdyXgjGdzxeYRX/0JfXbEd4976d
88p2/sCyQs/iLXVN4f1FIKG6w7YAgSr2iUKg654vXXvvnKzhNoNopbBePSYY3zrx
VkLlr5sTFrrMl8Zml/a7RjLkiS+5Scb3bVoWrzHOU8fhl9vp+oF0avv1uXoqukOp
y++6NH3HNSi0UCood3w4wcFEFQkpRjTbReU7aRpE/84SHO6Mod/Zb+xLJ0Ay09ox
FUnDtnBorPrn5S7GpgbKEHx5LvPoHzgzdHiAdEQ2QdeI5jkQ9uRtZA7EhoiV0l3V
PGBLICyASOhj4Tz4QHgNiRHlQ0hh5DKvkiMuXMQhXcgXQtNtVRb2Cdu7ESscA7i4
EbU/X6+dg7cXWzszFyQWLzUToXgP+fMmwZFxXWMyIfkWYkTfDRaPYGLMhd/PKi/u
OTtQKbF1v1fk1FpDM3ftlFDo84xedNoBY+FzhLl/y9Qqyyw5WfoaRfHMPa3w37x/
H5hz9CHq3OPQkQ8iVjd7LF8CGKNdK4MvV3afPa0QlkSRWdkzgCneq2ELXEF2837K
s7xLlylyYoQxYj4S6ovY+JRzgBs9/TchhjwQtsX+zI9I3+doDDtqjeoSNgSgvRgJ
U6jgVo4R/wd8iS40i3wEh0Dx01rxV97cqN08r9km5MMCuPTUkG+QWtNK6vQaA2Ve
OpiTvx3hb+CYXiwQ4v49+5Sy0cK0cgKzLwBhtU5Wk46jt/hY9I+rf8Jg+vUSjRu2
J6dORF/bINyO6X7LMuYNyoAcumgZ90f5axJ/fVFReHAeQKMgfp+kiKxxlG3hu+d6
1F2E7dNTNEQWcKS5dOq9I5w21WYdBFCPbc5pVMmtVQ04nAkW0CiV6h+wQnvO39M4
yvEOK3pL1h7oAvdf4gyxGZVfObVAspNl4dRfX/Hnr9bkXuTqywo6LgXcBcx+ITXH
7nTe50sHkNl+vcwQsGGmchLElCWiMBwUI3HNym8D+cN8YHWURDBcYGjZ9VeGSG5V
0pp3lh3pq/78YaJ7/Tm11qGCumNFKbDdneEN6pheUesAwrgWEZDgyu4WM6NWXfYw
m+UWtphB0NjIP3gIL3dIQw+kYB5LzeU2iV5fEJXdJ4+K+fzI3NsR0fbsXN6M+kGg
sdjer1GZhDHy0Epg0C/Qp2sjHB3up/ji7XEE5ao0drigc3GMzqR8aPsc5NLUkYfi
4Nmuhrw7J4Y6pnTqp46ndRArejyq+NUkZUu/6Pczf+Uy4AjsUYIpPzCO8A0F6qX0
OxCHvXWQHV6ZbDfKRQ68R0vYmfFJ0UrqiT6Z+sjMQYuOTwyekcVKPd1jaRPcv5x1
Y94OWNwQ/F6seN2N13Yb39ZMQyNqZpi/hoG+voYWktVGH8r8GFhsFVFcyuDs2SUI
faZQWtweOss2lcXMcWhqo+BGR1dPRAnjusI4AX/N9nMKPjEX9oP2cglkrbKPUmbL
jrOjk0HkxTCDkQnUxQk8h88l+ceikjBUlXg8igTtOl0+1dBAff2Nn79pexIQjwuq
nzr5g9e1jyQzWN465tl54JFuuOXWriC3uWg5iNkJdkIFI8n2tlWZ752KC1n5zxaj
oJV0EBYIz+h/6PXUNoERRFfL3wegZvLVlpqYHnyePJiLIhIYdUs9M8YbWs+Nkgdr
jtUWChdexOiBDO7LPqIxEvLRdO1uB9MATAEZuuux8IZk0SYsq/Ha78+s5fcu7ENL
vPsY/yeylMvVPwfFXgJSnPG7mTYeezSUT3S03aJkCaE2mu8dKEBVz80kV/X8sSTl
UDTWEbvfWy1+B/Qcvz1UfWRwTdRtVlUpCMa25ZDAfoC/RYOVtRCYTgGnqgJspRvy
dMv+Er+fXOx2X+l8EfG6vmVrO3GFgipILCVUZhmF8BKromeh/VGusC3UBOEcBA2I
B/S5MrAzV0vVML12miFutqiubvZXmxqs6N8Vxf8IxyHKEsaEqM96vNwujoo0swj4
zOPWmGpHhCFPK14S2OqfxfqBBBeObFRLT5UTZIzfT83FEszFKFBRY+0jbmxFMFuX
8WeAvHczu6k1BI6AbctBhlRKUamUOWpvgHKWfAteeJYU1qY5TR79htc9s9BLJVKw
AKD47TFSML/ZhkWP1UpqMqnQwuwQ0PRxSaOpO09q6glhQNlglk/oxeNtzV4j9k/X
IZT9VtGrpK2vyYORcqbkKX2pDjAy+4Pk6TRPKuWiN74JQQHK5S9F/LVla0BQEU1N
yYJlDjWVZxrVjYRdBB9UCvQl6bjip8C14RZHaiN3jmaWV3QqfDvZCW7QjnL37BbN
nm0UMxh8PvwCCxr3M5mVe8QkOZHKLG+mg6LW0r5t0THQpgThSOB2uIgcTdOfF0RL
d6PUrO3J29RsTt4rtAWYv9pC/PeDsRWx9b62FHT/W2xixddsAg9x28N6MjIu4H2K
Cj0vKSiNP8YEiF0Mi4kbXtqvr+P9nU6Eg3EH+fNyXJPGYJoh7Px2UcSaEdLPDfrC
T2yjqrCO7387VTdbHUPbbuvn1NrupBmuN4nsZkJUhDuusFCKmUaoKI5NVcYUfO1u
fIZs07QHpOs9sQwNZgzt/71Ry0n/AlTKlh8LR23DhUcyt1lzWT2UiEjouhrbSxZF
sXiRJlUpWF1e6I8NSErmNCMfc0CB7r9uhSdINYskKSBVl+Wusbze7Z85OEFQ2bkC
IfyaTl/+sCFnTJmz3NDwPOrCy27RZw7D875N6K8PD5SvG5dQ2OP+3X5Nejj55Jyq
LLgjvFnvKtPLNwc9cwRPHPMDxEtapleL0l/wm0kCl0h1/L/APNKo3ZHL1qrbhe0+
BXmBwTIyhfzMyvqDu+VdkdDS0E3Tl39+LnIKEov9ZJLWRlltYQBRf6AVrQpNPhBq
Ec0iyWwKRXzDigyOGnDFB5+iJgcvAj0iwu8sCP+k6J1O0+uoqBfrhWHOsjGwkHdI
CAU1OcghnNlML6yfmcoGxRRfLrt0q96OewZrx8rxrGgaUudvDF4z9UstfleFGfvj
f5NdMH8jKEcQuQ+GaBPW5iHFXT6TmSdzddejhClodaFvDf/Jot+1NbyWoZhk1IoW
bVUTfcIOnrhlOOurfBncM8alx2VoK0jildH1ZC2yCggoV35NhI5wjuKg5SoFoVXs
CONyU/3Nl/YDGHxwjBgP1jUCqqz7GQHPOG5iNbmMsskSkgcO4xGbL/gaQo4y5Dwh
SUPzBQnhVUJSvpOmabc1WcZLg9gFJFJyMW994KU0DN4EQYoUq8zDVimEW1Tqneht
n0s7ERJmLgcAvXcwtZBz1OfztazyUVbt3seK8a1QndsOH/3AC+6inYduXNuJzFfQ
xiqOEm1mknvJhs0hVmEio8O2SIGXV7lp5S8MmqpNAxFACQ1GQTnmwp5x/fvJSer/
vDMfbEss+75Uq1Xv6OXA6xpKkKmK72d4tblMKOmUwe0W/dP9E6wo1dawdx6CScGS
StSi7n0cWGI6xJ2D55Z+4mIVkVRMv407oqvQSqlSfdSRsb8KFNDhRvIcbJvvBJwx
xWGg/lET+Ey1WEcfuhd7pqRCeK7QhYrG7oKUlDdNyRyUW9QzlsktJ4kgbA3qg0JG
GFpbVdJRIRSeRrRjlsCIkBKuJTKxIqnLsSyxSxyCzXvKIc30XGFYBO4ApO/UbUm6
jFReqhIRx65CXrxUEUHQjWCL7YpXOqhOHoJ2JclnQQ8FDrINy6sDlXfgBtRamENg
XTU9KyzARVo+vN4VDpfInsOq+VzL7l6FQ18+2x1m8BMzs/WLs1p2ygkxUbJ6gpNo
243Ygoiymv5wju4hdbwpOWFDVj9mkldD66jvs6L6NsgOJTnDTbqi9x2ee6CFzc5p
F4LWvR0xUsQ4cVuJ4ZWmHhDg9NhWNUNQCZnXMKvT0cjJJ+rsgqGtFloNyRUcAtzk
1kGO8KAcIrh9t7TzLuVSxg4EhD9uPM8VxAe69ALn6fx0uJtqcuNpU5FipmaeUImi
ajqAK7bjhGYSSc4RvYHrTqqxWtyvvGtPVtJW5gChHmO2ihvt4zPoHLUytZVfNPBs
qM98v7jeXuDRhJF3f2UZmkuopSqpJrenSMcCs5nmKgCyrZ4M2HjlhUTYiJlLyoxG
Uk2DLwlcuA+syXg2GL4gYpAUP6tr2+EEJWJ2DaQalLFU/tSbhd17fcGiTy5gD1iF
xVCRmv9oplVdFsCJ7vbFvKSza4Qm7gANP9IwvhjJdpX6paR0enK8+s5ykudUM1Rq
ASVw662Efe/JkO+YgzUGgXzqAtYVRdi1C4rZEUtMXUfnqHQ9y/AtNR844uT7Hhrp
5+SNr4JYzmKesR+W9IU6ARl+WDa12tJ8LkhAuTEPyIO8rjMSZDPssbzixmctL9Qr
WcEj3TRe36vdxtH/NVMglCMa/c5taSsa9fD2JhSJd+t6ATNLMS1vSIS+Oro/pSUu
lXidBy0wLoVdKlmc9eQQC8D/J73LPEHoM3v7SgnVQoEltYNF6Qq5/aknkTb/b/E8
reOTbJEtq+vb9wJUKSvUU4xQCb+4F2ZdEXxXB8gnJOUd60GPNOdNBjipgcnlCc64
ZzCM6lz8q+fr3+yJjC3ddwHTn/Icn2nKDMBie5/4FG+m4ilMTqv6vuA4WKTnGola
+mR+/7yH5XVkBX1Z3Wf+ByipBQBJeI+6TTGbNREhlUM2FpJvCKb6xwI5Z5D5duOv
XTeTxjMAFX7l0QEvZFujf17yPKR2fnMsv1LAhBaDL19dLBN4c5DFJcL91n2tYfZI
g3jYqf7j5i2MUaXPXKxy/ZY9mrHWIdkL8mTmh/AkMbKB3LsuMFKfEdK0eOUO2N6p
uULu5dH2RdBipfIsgvYiMa0/ofYWcF9kmbbbVnhLariwsOrFVf/rQhVr+rVR5uqr
+nVumEXumRVvPWIYd9yCi2qqnc9dV9ZlKpUcVX/xwYzmX8QqzEFXPGfnaTL+A7Wf
NxMte+RDfuRO+TdFKRClKukK9pea5YWXQlfWtkyfn2TSl4+SXZGu6E/ewgjFeWTi
8C2V2a4EVT9miTwDEwaTi9Rq0T6TrU0jfHSoAToyFwNjRPOXzR94TA9WuiMg98s2
bWiNv9bqrVKdKIPIMJWRQAp+qUWFmk6hPgEVPNyeQY73BdvBW6rTzE0uiYuPVnje
y5OJLYQc149uGq/2SrmdiSjiaxfwSh66uG6od90aypKjS2nKhooSu4h0isxTu8Wk
1EHYvrtHeJTkgIOkF8YJ7x8l9M19fndc0cZflmSkJu1iZ8CJlGYZFtz6gUg6DoMs
2TfM0twB4xoR+e8FZveLFRc3F8FY0nHoby2KNbGx3/HrPkc6aFqte0pVNgLj4y0R
EPRc4GSRWjaGInjJgo8/ACoxOIz+LqOaSLw25aPKxNcJ4isru5pok5heFVB4XeRU
qpl7zV1+59EnBcw8KfzIJLPclQEU8j0mhb1RGg29r1aC6CkRS5QbttzSSDij5CGN
TlVddyWyHbds79mA3FwrcGy8NrF7keevz48luG7p3CtIKZINYN2EF6yMuD5B3h+B
FlBxLxOUIgqGnUxnsE3aJX74dY/aoo4bSMFdY0L8l6AgapsJMwZ/mCf51OLD1XPB
8K5fzedPoFu3MMffbq9RSS1yWn4TufhQLp/wBJvj9Pd5wgfbKWHDUZq97CCg4FAS
fpKMytfLwk3q5K65OpRVsQc5hBmimaPJLzsev6YwJoINUByMYUyOeYGwnSZAT9Vs
AO8VOfUWP6/bb5a0GefTTIEJLd0jC0UHPOVx51JeI5Wx/Y1XlP3s1KR12Dqr+x/J
3cueF/bsCJpzfoMbuptmaOPWM1r6EUeLf/r+ARnduXAOeFN7R+wjGl8olN6WNtw8
xiyOWaVfwaQwQUnjzaab4SL67wAhTAIrwDClUBPInY614Jj2YQrgDbW8kOXecPK5
dAEwOzorzWIIRv9vNeW4L4rqXYif0Edg12UctOWYu2RO+eFk7xogOohn16ih9PN5
gF6NIZPmd3kF2p4A+PQypWrNNZcfJ5mr0cXDDWr5ph2UwJRlBxUtTPqew0O4CDUy
vjOWTFRNgdGAh+575H7cRMoUqskkYxRJBMOwDG+DcDXrcNgfu4Pcwmk46l9lztMa
ZcuOHUIeOEjZQcNsZoKGVd24vjlfFf++ynEy2RQD5fQ8ZhCdB8MRudEHsRxwjyJV
djjca0q9qcF0n8isP0L8/x+pPlIh11O0gFA2MxQc2cqNZydEVQ8+L902DXYRaFL1
Iul+vTdzyDtHizbD9utRB12bKsapSx1CuhGOEclWZmu1kti6iTST2UAcI46aePb6
pvDaW3tm+f2lJT5DOzevH5TCj8nfzQ+TIVgc6tv5Nn76E8s3SHpF0i4UPmQsbZdi
pnVqyr6rv3Hd/tFM5OPW7Cum6JeYFa/6FfIQD5oJgcaPbprroIbr4YeaWfY914aX
tExCCZbtjmWneDOQNrLlDjLvnpBIvAya1J561RPg6V3uc2UVjYs2cE18mLb2D1Rh
IQ7YBV5NqokqHG3J8knYvQJR+nbq+mR1kT3Y+1Sx7dPgYtEIntDezzb4K/dDNezu
BGC09dbdJa46FKq5QdwXuOvGScmxDCdyvMriRAdQswCwCFA/nKxh25QC97hsgEWu
FeQq51SYfQpgQ9hYx4S+dyvV9ixd4wO4JMBfhCOT7qYjl9ufJOinNicb30slfUbW
gtiUFyVetMZcxvh/mhMkOWmk825SsoniTnYbrHXerzkKwDKLQSw41UGwP1s8YuW2
C1ZTfvdErYEuJv291Al0qyFXTXSDW/T6DIiFn4bNNuyj1XwGjEOX7DS5fXEXPmVH
4AGQwMhgvXZ2yRYj1erUAnzwKD36j5l9bdlu3UEgDCrRcGZoFPPF+9/SHF4nbtO0
8HHRGNqG1mVdufidenzD1/lrPtPDdew/7mn2wErY/T+KF3oLYxAP1UGbZvx8EYqW
tFG5H3M+ppqBofuNCso9UYpJq9yP2m1Z532c2vJPuUYrwQSo3QhmPWGDd5rhh3aC
FYdN+133kne+EgD+mwWg4XnNYJzGRbFMVq2HGhKhYJAjmjnlTrpYVNEa5pRrQSrw
LKg8R/JJGh8BTN5RYzocATfJJvyjE2mlSILqijbFa1TcPr7wyJOUGl+fzU3Xipub
2ym7SQZxOi/OUP5H0N/OCuooZTP3Q98TDLms9518ZkStoi1YcmSjtNjuf/MmNfN7
HzibHHoc8F46gXYDczEgPCfXqbpPs3OHV4zoNjhw8TEXKUcWjTYXfpGBXWnJYF6q
a/Gu9yAXZJE5mxa2egJ7E4Okjd3786WoRBuWhdhDmL4YSinvMEIj/f6/7wLRU/jc
InBfcU66e8X5RpH8QEsfx2kB1ZQ+vlNY/1Xw/ERJehdBnbAhGHzWKzn78yFF1pfv
B1RGOkyz/zp49dR9IEF+kky5XsG7rSuEP2KhmZuSLSrUf6BrlZbIA0NqvfORu3by
J14l7Q5UoKG2pDBXLXmIS54kyPPvbH1WYjG0Xe4oK7Jyin8PtrLxa+KGrTbreyzj
gBUi8s5hq/fkb4P0W6P+kxbu7DppkMiC30yJ7gqtcWEdtj6wXLsRFB07h8sS9FoE
GfGvKBlIvjGeLLqiqHFR7rluxaM3XMHz63sbFci0qFI57tTZiEf2ZjQOsTz5mmHs
tOZCF6sPZ2HYWVAh0+v7FMSDDMnj7qRD0EAWSm+I6zG7z+AIviWTS4w9EvxtiL3B
69JeiYRZRtZq1WjxL55rdSm5oXAMN/nDpvm40WGSLp7NnwWGJhQGz1N4pzuKIdur
IRKF8dBFj8rA2hoA8Mbqmyx09zdZqSUVk3LAEIQ9o+gPYI4lZySNPU68AbiMXb/8
HYlhgP06flcFbT5I1AKfgY+5JbJHQR5ojxePzf+swueTgnMZit5L8mRXH7b4X03C
83S9jCdRFAlWOulHPO59/cgMJZGYauydlq1gWPW2iS6misumFR4OVCpmPgFpskpZ
GNFueTBJ0deYKC4u2NkyDJWtLQyh19T3YlOnR2J/LOuOypBS0S6GLAgTyE3lfWNo
jM4e2g3tcN8fIjlA2wN2bP0B4fByecipUaXW1RrbloEgYxdKgtciurwWuLem8nwQ
E2s5kqkp2BO0VmNs+FNxYIG0Yo29I19kRs15GnY33AlYAQc50AErdE8K5nCJY2Gr
QhCWaF0yXeOcB4h4+NZbTP+BIDU/z9mIKIDTMKS2I33cKZDi25rzzENwJ4gaeZNw
u6eCGuv8IF2dcQnBFV80OjCfQ3/Ldr+E0yeC3vKZGKE27BJG46WxsbbpUNsx/r7d
5wd6BWzagzCJbtGXH5mM5H0XcUYedJgFlAnLLwMyKqNxmm7oJWCQTSKbEkJf411+
EPPJ7jVMxSobMgkmtopiy+vywvAEABI+Bf/lI+kwBJL4pvw6c3/QsIercAVQs2Ee
7o5FUXDkp3/Co3unnn5/yUx7Qd32E5h5Oiu+V4HDTLepbBdJDEJybfbLEk/YyFnV
010yRZGaavKV0KOqbYAJ1oh7kSR3HwNOH2uMRYiqS4uVhaJzaOO3m1R0Qdx9BTzZ
XN+zF2lhGWDNbDrbs7Twt3mksEQN/XdjudEkvfQXtEwMxpLSzVV18NHFaXilrNHh
vVISs3AUXDcg1fy2Vr/4G1B7coFpzXh3tkJma4i5uIRHEizTLX8SQczXeo8KQTMe
F0+vvA0xx0qo04MYz7XP2hoZ3q8LfGHdBSCMFhsnQfUzquYBl5Fv0gBZtC5nZU9B
5uC0FuY/qfCR0U6EaY7cM7cBY1DmIC1L1pN+Qxs3IyLO0n77jAjjdFMdABRqrRvQ
Mg9cUEMp0OsCXdGNlgilvKG8jU7v+fTVZml+lQhCPpO38TP7trVus7THJ2AGc+tn
magdrGEkybN/JzwoPLVB+mYN/2olnFqgcsv/Dw4IysP29d3oKY1lU2VCZLyYBs4i
y1QLqYVy2KLUZ3seXYnf4vBU+y5/gFIYvq5JYz1XbvXc7YGCv5rqgaNRaAdtmAuS
gkk3HPoWEgSLUaL15gQOr55mXKgEpOd+KJFPxn3+s4AHtoevv2/aw2ZCFs9esk+5
Bl2fW8sqi4qbTpXg0wKupdmbyUEMtP0IcIn3q7UnM+p0QaI/BZkA1JtP8us5HFbI
KYWfveM949MMngzE7rbozRGu3y3ME9genxeQzxbEGV1O73OZQ5c1lvXn9osdGZHs
NHmoZpKAx4h2liuAIkmO9S6e8YpKLf1U8nwxUWIHpfEnplMzrnqLuwJeseKXDlwz
NhIozI24TO78cH8qWecTzkJComGeFo4jkTmZVbB31m+Lp8twrss9EKuMOUzXgJ13
KDxV9nDSWGVSX9jk7GFwocVZ+9nKjY2R3gbmBAIlnCxeGAB2yCipQJifYGgmk9yj
550dcR+9Gj/orv24IaqTX1N/EHbHheh19zrZUkUbkUK5fYRQ92Jn7fmHTBiqtW7h
La4tMG4yTlnO4URYZrtyStvT4ISO9+e7DXW2FEf2A/JjNhr10XO0YScOE8+H/Me4
1OMpuYWz1cODA23MgSkxmSq83OJ+c+uGWtj/218pIveo2RLVRHai8OGgtgzg7V2f
IYcLuLYMJhzmHXz5hN+65A76H+f6AQZ0cv/NhfTFCduuKx8hzz30GJDCD2VghCXx
LMWggVkBd/+7wJmFAKQnRX7t22h8yIq1hz41yIx/qx3sZaYOCUJ81bjGutuAAbtm
4yxjzNQRFSsAtT09N3naS+U6OxUd07A6BV7FNP14GKwNdx67s3cvCtFPVQpn3vfB
lpRlkhH422qIpa4wSacPp6lidUm0WZ3qxHnQTeqdHj3s1mBU6KvaSVJqiDeLKZFU
3XYyi7YiIoV+FaI8R6P/ZqjyBdr02pyjTuqpLFToH0EnXe2uJdcFUSNff00Y/7N5
voPqHoFGTq9npGo6dqLwYmMzwrNOrGlmSgLurZvAAcmXwK8A+zal/1HUXY/7LIzT
d/xIpsdRlkxXCr780XbzSm6wbc2tPU5RxP1XdCt4PwwF1bn2idZr+f4q2bCpznVt
fMgdQ4mrAkkxbi2JxEkRo6/PGDJO3gy5m6bcxNxKjoiSp42md2qruC++NpfzcjYs
kAkUqFhPt8UTIIeNQpkz0nL9BwRzvXaG/FD02ZMSOWs4xf+dMWHeq9uhhUoYAwdX
ZCZK1GfZsN6/HjbYq1fT6BdGQUVhvB64DYAwXThwwVo=
`protect END_PROTECTED
