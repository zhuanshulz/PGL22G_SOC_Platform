`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kURLWTZTiOw6cGC+wO88SElQK+pD94yG5AwBhyUrBVO2s0C9S9kgG82jCmfcXFPR
/LHj8XCFRDyVUs8ckREhQR4+mkcPOebdEWaHFZn63RPJcFEfSxQbyX6w8XGwVws7
IgfgraNsVKzPnS0VttkX2s0uv+4tOGIsvRxmuZJQD7BX53oOiNDMATfTd63Q94E7
h9Q0JdC5L7LRudc+eS6ebhnnzgRb6EZ1UuO6h0/D5ij8SbRdT9SDnp8G3ssvjXUf
noK53fQOUU8srf50kWxRCqfInStooIw9PFHBtApir2CT6zaekbjl8qP/KBZTkToV
vYQLm3apjPSVJktwikpGT/LS8qlOQRutTPSGOA7GvjFDpKQjAvDh1ZI8M69dkQUd
UunCLPKPSCbVvvaKozwDDsVRfPuKJWN9bKtxm9W5k2zZZPOF+iltZccUBi1aWoxg
3g5X5aHW5fC1inRlhUViP3GiVnhLPTtG4KHIFQK2dFPlgz+NgqpjMZGmvOAZZFND
nHrTEw0d9y0aWRnwoXyUQi+j+6hDMoyFTPq7aT7VPOv4ayPZBKww6U4z5visP1qK
IWL4aqrPnOOPztr3dfRjn/dmm1RnYmvW89G97RRawxqP1OOTf+nTlq5XiyAV/qf9
iYChWo8kJl4BkL6NB8gEUXTa4GDSFOs9mqRg6cTESQXkAHM6VY9ShMB7cyxlxMkB
akmooY/UTluuh8JvY5RXtSMMYpV/6b0/cDWCUgs0EGQB/A/n1u+Z+19Ftc3RpnVq
ncpx5LomgNfKSdlh+T4+63wSE/m4nf14HZNM2MSAqIshbw/uThFSv4lND/9V5Unn
wszTnMLhBNjXFrMxNShdP7UK8BusDUoJr0JLcyFypQhQWrP+vVDp7LSzIK81FXfy
n4rrBAmNkRbYfspi5d8S2vQ6HxYCgas82w+9QjsYzdGQNQ2mILFhKqT5hTSLQi1q
xZBhG4G88C9ZYyCcmgMOdBvpF6pIBQpvMNwi1V6D1k2HM9q+uQbbKZL3N1jwhzAb
`protect END_PROTECTED
