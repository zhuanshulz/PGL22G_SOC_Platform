`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v08OBC35Bk1eUEyTvgoeNJXaEjTpmvYVAz3bVMuFk+u3gdXwRwN4S4El4zSdzSVc
ST5fo5NTPVkORfHG4W9cldnR+EqwxGDlJd7+ksOxtYRdaevFnyBhZUyUda9IZ1cb
NR5lzH0Sf5VUdnmXIqSdoFbuMcfIqRdfbBsLdGWdIcx1Q6WOZazMTOJNdaUDtKF2
E/4IQMpPYDZvtZuW6tk2i6d5RrLLvZJoH8pLKqAxnOXlOSfcM91eVTOB5c5YNIwg
b+49mEjW1MLjZqm3NpB1RUFSRK9Yddz4QKH6y+H/6hS9+h8aiSiRkLDPhtOLV9SN
/K+VssCdnD7fnhsNYdCdC1Qqip+Y0p/T7o5tK1nCoAIJavtIjkCBi0HS0TMwkPFs
KtJtCvG5730hKzaWFsj9yXIaIYpVHhd1w4t46aYe5pay1RPSZZbI2/j/zqvbXi8I
o+B0tbPJvusztCYNtKgLjJG1HTDieO3megjlKz9dEZnJGfwm+8iSBvAGO9/Octxa
2d6xO3VGe3Winx5T20l6ZU4idsMSptO4phyhwgtvjlpzdV/WcPaC6EksTWyUvdH5
5DiicYNoGYzcPmjpJ/hucGfaPHkFINnjA2JtFdMsfpyXC/H8Kf35vW827tRt4t6d
67hrONwN6vUswVdEarFswlyBDs8p+9jce6TdB+xolJVce++HpJUAqAYD0f+lLS0m
TykpEvS0WR0/XKaCwBKo9VC+t2nKT8aQuw9atG418GOfel4PGxk1l20iH66yO7WQ
e2qjyg1YW1cfTtYK3DFp+thu2BMXKW9CrEJeu1yU8c/mM38ZyTwJYliuK5LSOMCQ
HxKqopUfzTrgloMnMm4CYEDooG4H37ANXDXhOlXY8Sw=
`protect END_PROTECTED
