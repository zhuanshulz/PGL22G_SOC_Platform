`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
puD35FxtNT9XSV3gWTusQNsqZ6ZvUSlsgzzozMvbC1NvH17iwp2/F5ZscXiPdSsh
a5pQRaFo8gWv8ajxpbicT0TJlk8PxE8H2WVrLz9kUjFtin2s5JoWSSlooBQrGLAb
RoIhI3Dy/zYA9A1/bBBVKgbpIC2PdhEK+zaE5WZxG1jxBg5Oa5v0YBPmVt6tc3g9
TW6c9wd93FKaOdeKFPBcyrA8M1/Hq0NGLVUdD5ZcKVrjeZHHftMorKM5gDgjrLuX
roy4gckOoz9gq1S8jBuhaX9hhqRtqda3oDmET7bPN4Kus9ABr6tOCqA2rEcz6x8U
oORc8TWbmAr+KXzvDdRUmU182o1NhaWhND8U4C7WkmzDOK7YObjhN7mXPEZh3ecP
VMzbEmxVf0Qis8Kj+b0ihfickgMBDmZvRfLx0ESAJk0nrc4ndE5DctT24y9OK+8f
OJsao79857hqmrkGvzgze85fOyFpisPxfRn6dDG7zNcpNZd41GmTz9u8kkNi+5s2
E0QuXNEoVtcBo6aDRLGkoSDy1QMum70dMBInWOWIxIlvIzasavdYAUL8Ghbg4avw
nNrnABt0VDvwUMFw4hx6Cy8yMd455yz0rldsdSXraBIMRJ15fG9NgvFAypymxtg3
ZBSDeaRM0pv2n3T+uNMXBs52oyouiRn0kRGM15l//L1yvzhlFEDbhMywuSt/7JG8
9HYzoSxoPW7nI7M63eIy3kkwGgBvQ5iNsD+xAhk2H/SSVfC9Nd4KPA0d6dsXu80L
vMD/mKt8Yy9bdwJoxioUKHFp7TO+Oi0V+KlEaYREWk/8EP8wR897w5woBdo3g/px
ULqSRXMbDsOyZc088aUOnXhQVC//FS3urg8vO+AK/+E7LgeNxm+TdNkMPQy7QhKS
wua0oAlLggst4CpRHvr1DrHTYuWApFSS8qFmkppK+XLPgqORV+enn4J89vVAzb77
Itr3T0PbzlPlI4DuDx3u6KFKr+btoWTCcZwsBWRfvhJ1/M6W3zs0Y4W+afz4Xsyl
FYdcDOmAfpxQprKm0npsYCXrVPBZYGsD2UjAZgcgMoyhDP3vUO9lwELXd2SzmZxB
ij3hbdqw3dQO0ytMzcv7bx9yA+kDHJ2pQRerukqHs8vq1jBBnWUKsNmMMCBpps6K
863k+LxvgfBjTGmFwCypKjUqVM9wnR79Vx0f8lMQKH9meCBftIhQf9RLsN4TXY1N
s7kAp2i38XUIHhuPoSpV6jDLSPKHnS8QxMaczZbtX9hmvvUsYeNt3Z99AbYRPuHl
loGtFceQos0237eEvgJ23V1UBlDxBCTNROX1l4nDLK+fHYs8KA1YATWZ3K9wS78N
8YPZgM00wn71N/98qfm8qM5wbKSqxA6Yy9TLgYQRDmrNB4Ld7BrA4O7lV7oZ96kg
p0uorGRLkbshOmsWSsGqW7+4g0peOA5rlVIi7YS/yAwk7oNOT3UvzenvX/wcSsAx
/wdTX2RND2Ymnaf3G1wSOYLTmkQP5W75eOS/dzw2q/JaOOEF8EKsKeVwkXP+OYBo
BXYvTgebCWvUGOzzO69IRYMW1xfRWCBo6zeh4tLsZYAjSYmuP5ouIhjKS7ZGEafK
Abj91eQw7kVKjWvzDQ8pmpeeMOqVen26rKY/4DIknwh83ItLjImsNokD13ERcI9s
DKICQJoP0XQdlXHUbT1iHdz90fekuddJL1NR0l1nlMm8Iccw2DVNxP3swxsGcbQZ
fB/hAoNwazlxoLkQMr3+oItQvFFH8hR1/4Bq07y0+s3ie/aw3DIa/BuKLG/VdJ31
U1UiQitY36EV3svFSWXkGfPvLmIXnyfbyv26q6J+w4ZW8iPZ0VQjK2H6VlnX6zHc
5+ZTF6szD0w9uxb+3mUx9Bz5PIq+NEBT/LzyLlHM2MqQjrBjfxy6zydjWZnzrW9L
Yj0h5SHcFXGJGylcqapJOn3fCtaAaDUpoZbqJuhxcVdZE/zlqN6WVH1zDzEpjGiB
3WkdlMrjszSjJQhM56TDW5qheC9OR+Ayeq+eqr1wcuEMSeaZKMedrhiVLyI8Bvfp
su+FZnSCsnepB9IemuSCtO48ti99wXIIR0B4X5h57oQP/PE4iaSvbtrqWEIdOojy
45xfrA+ET1wxuIK8StZ1MIYEjRnWo/ZAYKuLFwm9evKSWMWRVXZoU54hLBxX+eMZ
N6V5Wo7Zcup4F6M6TwHcRhr64Ksy44ulAS6SZ8Sw4iicUIsm3FERhi+Oqx1DkSPz
Oqg4v87GMq7tbcN9vodU+PpcwIP/TSuIKpF4PFca7WwxlxQC6NTYbq95XuIZbTXp
c3er+TbnhEqUz85Vi4AJrSO3OO/9p+XQqVzsuIjKeGOu+noNu4sffTqCuTkl2K0U
gplgg49GzDZ+W77n0pRUFjrl9VGfXIEuJhTmGuHJidB2oAiE2KXKqEKOLLfk6tSq
Ip3QC06irZvlrnExAjw9xPJQODPBWqvCW7BPhIgcJuqSWhQiSwNPGDvTP18oYT4i
/dloHg7ADOct7PXdkOqcjSQ3v2mXVxOqyqns+yJrstpS5Uvn+9fQnayW0bzpeOiM
n2ZzcU8byPP+VYxbA2envuaEJLYTOVKOIZ5KSv5lhmjeRU3b4OZ/6ohkh14GIcOr
kYqeMEqP2zSMN0nX2CNxefSYstGwxr+ilzLJyRq6VWg8EdftJmi1TApYKxeCEy70
Un+toPIWHYQZOHLs5vrlbUNV2f14+/erIQXqnalQiZG5x+vP/bmM3udQ4PS/JthK
oWz8oBDMIN6dlFE0d1iVxyHPeOt3Q45Nxu5NQSFz5+ruMdcN9sqCzcD/qYjCqCzv
FusAkFEj1pabue+2NH1N50LuKkCr0ByVyusIriL1QQF/R0W8GaoYLCVsVJGVjSzl
K/PcJSHwkxlUXJfA7gD9nmxUYgO986S0NgX6fZyb6OO9hUcXX1v8H2x2zhNhLEXs
JVoA51YFNLajiZVQR7RUkM+tp4wzWkGbBTeK8ci1IvIXKpRy+ArD+bJWvfHyTwSb
jeH5AQ4jqz/SpF6s+0TxaDgPVrDe9Zbta5EgoFRNQg6d9w0O+QaeRJmwbCgltVO8
BiY/UNnvrv/IFLcFB5Kp1v91nT9HtVZ4g75BdvTBvWJFd8dP5EdCEKWJf6eB4Hgt
0Y88LpnyDmCo/hJu6tKck+Btp2pKL19MA795fYB9do7XYO0T14qG63I5QpAaCGCu
TkzoU+FT1Yvuy6wK83E7B2MojL/jRHcf2mQcS+F4Aj/w7dJch1uidn86AO3uROK+
plsiO5O9iEK3BMv6A1rpSQbOU7nghQOKT0dL6W0SqoYstKaEyPBZp3/htAySgmMD
SfX94mXsTdapmRV3rhzvG3yVMcaTgSAIdjCVlxHgVs9FapJaSc7a3iSFbLHOJyfk
V30HOitufktSKbArIHyTZWzXwJsxIrmVy4QhsvhLJ7r6P7UIW5UzaPMrq8wpyahS
8+ODUlKHmohE8WomE5TUsOLz9/uQuD+ebBfEusY0g0g/8EfWaQKnILMkyzAt0Nzy
s4h8PaMraNm1AL/0fNxfUFkoN7/2VxgK10Fdj4JSB6zJNivG8v7TVz8D554DMTRq
EvHnzmrkw9WMMZ7MNqdPRi6F6AKjNIYUbMimtab8CyBmI9jPmSOycwge4np8lZ2h
/TzL6Ywq6eErHKWpbrxrP6hYtP/NNZOT77E0lwc58AqPiQWZWpkMrZdnQJjQ/HnN
ei7CYTP1pom19g7BgRP1OhIfmXoNZ0bXbael3VNMkFlI+9/nh/QYye3Uk29ia8NJ
Y66RkjzGmx+RnEoAVZGo40T7IpqYBhrZYdxFldRmkzTw1TtSSVPhGfW1apOEq42f
RQ9aZLngDzZYvp2EOKkB5s92duwTUOzMyyQABNg+BazsnYWo7pm1fJBocsFk/fce
xzpp7l2M8FtoLU01nNu60I+gkzbzM66fdGSQL9TZvNJmKFsamRNcirtNmX5FCd/g
eh03Z/PlterUkZyfLQMDt+sNA1/0PFnsNdrcqbkTPALm/coBrZLi8RFrh95Fh+tK
mr33e6UmALU2HA4eEdANL3hLJEOHHj+G0XFBx4hgC5qMsHcZg8OhyMS+PqupdgOF
j4800JLSP/Ib5SucY/tEEDJ9fsuLQxQzVwCRFJzxPcv5vAAMv2bGLb5DtXbQz3yD
YNirMeKrce1x8StzFEdkGMMrZgiuT2Hk+pg1X7RUpWhCSysMQg7ldf49dQ3ME5Z+
PGIuaChsRo7r1I8pnt5g3bE4JQLmSmuSuwjYgkJaTuwSvKT3QtQcebr2AU2keAG6
P1kRTQEoC4mRieyyjBzkmFNcQl2Zhd24/bJ94ht1bmvg1UcubPWD1bGfN3UfqBu3
Ch9uLkFbOjkbQOPTBavIj1fVhlnkHvTYRMjnzQxTCkpIxfqsCkppGMGJdoY1GzoU
zxduWXFBA4K5voohU8pSx6d77fFtKJDzfmP92iQufOSZeGJedAF0t9PEh24+KI4g
SrIU7i30hSuBg6d2MjFFt413jcey2nZ9wSlqWuAQihvsWZaoc2tJ7sHJSSYMS4WT
027UA4XIFFxkvHwLoM7OmQC4TkfbZ4wGuhpyCfqOcTahk+bMaE3fVzkndIyPrRL8
lhH7cge/50FtmQrrczDyDVbWpaNnV2yksToae3lfJWSXeXY6FhNatUN9FT4+VMjB
Rs0w9yU6f9MkPrUBsEKrexlSNTa23Ne5zXJs+z5bihilZpwYuCatz3TewdqKuImR
lLdDXDrWMfyRGXezbW3LGPBPb8HLZtdCc9GNc2P+iyUzOx+VUfxJmNf5nmYNhprT
MHWumOxkd2QAzn/go1gem5g0+skz9/q5AO/5U7WJPt7eItuqVtD7QXW2wAu6QzJV
WXKP0YdQ4WgyC1KPjJLKNWjJfGyOMH27r0OcIIxgy4W5q08lwSOnV41DwlO0M/pT
hApY/DwWajKW/JlV+KGysTu8K2sh2Ql7l6Dz6B24Uam0gpZDXhdYzu8HZ8MRmOmj
ZeWRtxqjyDpX6sH75bqPBJvVFd8ocsKEsAq5BBfkEoOjs8IhGlUe2ck7dNoiwO39
Q3feNdkIPsh3d2HIKCIUjRIne2dfDExAYWrdlFymo/NhJtpoBLg3QKuCDPpvW23l
Viv4mW3l0xyzmKgOF/Hnp7lXM5OF+AwbG26ujZ/X6mb45fpL3qD51lRZOOlKmXNm
3q/JhVTuAAHNC9ixGpk/SpQS2oekbBUD3TNicn7InpCkuR00t3ionlsSvwMFKPyz
6ZgdU+pDUYjGa6HbGRpr3BwyZrGJIfruv7e3IGxbS36oKJOr6PRiReyeAiAK7mUj
/MY2hgOuimHM/y2DUYupPdaSac0paDixEKaRump77lCghveHPbC107DaTVoh8Fz8
rzLQEPyndkEzJ9JP/ARqIDDTuPl8GESqWZ0KAULmw4kmJ5L2bMKwQUVMh5/0ctfM
KQCR5CvcoKyZtBLgHU1mNvFlAGCOCF1PC5wrim2ty/ksSH0FQC+ATZx/xw0HxiAl
xsY7Sd4cgQbCn+G1/I70zKv5FLiim1BN1HWk9cXTGIgO4aIJsB+jwwJUo3pw0MSe
SBu44W/dcqUnf/zTvQ4u29/DCJZZK1DRZW013qXl6HyFF6qNyqHAEv9AyJLs/vpb
80YBYTXrM2r/SjgZtXgdXZh56UxgjTodnAuS6VELg7Jpx5mez+eK4iVohbyN52mW
xY//NDIa31vwoj8qfb8UVFuN4E9UiONoAnSEpiLIK53CRU+XyjN/VZlCVawotnUH
VfBavkgQeWwRH9jCIsueDodSz38AtFk2wAt/RaoSRhL6iICvAVZzMl+j9NQBJpWF
bDzNoTWjif+DHNMVzubLRkndQjtBfCG6j22bLiQd1LELmm98Fo1THDGu6fW6vX6q
5vjyozq04q8Yr4SMWkBJM9TTrw++BpnMDiJe47EB/mvvjESwoOP5U6sVZ/AdiOZf
WQGulMaCpHKD409Q1HLXKtbhGJzk9v6y3HKcKnr2n6ug3oBs1xVOhL+H/0qmTVt9
wZ3VpGR1tszuQwe7s3peH+xP0AYMiI6ee+NLeiFpsycY15jmnl9W+RjmDRtJakkJ
khHPS7V7daF94RkzoU7RhsJBf3cl26QxAPPwTC4S5auCK9gj8/3uoormvYsQvWTF
TLkulYzcDZSSuKeEYLfxtt85OxAlsbQDpNOdapbJngmUV41y5ZQBF86hKNyBs/aj
+EutVZ/X5Kal7cIUMCYB3L5p/j8bLES8OV6dMkrvSqCJFep/9Q/bwh3KP9d4TqWH
Umadqbde2sXidquuTod2/MeQtJFAPRpM4HYV8VbmhLLqUaM2jsiYHznaWxgcODky
86hVHS5siKFZrFbY+srtNWQltiKg/TthOTrC/AWZHxJyHc1GbyaLjFtKGA+JAyrG
2qGPyzatnUFAORzwr5XDr/tIrNA3nLpxWjFddkoE01JW2TjFM+gI+WSFjw06zx1W
QeuR32yHxHxdlEJ/hCl+9SD1JfNiR8r0vWji0bxNW/dmPWq2m+D072wKGqXpnsVW
e1Zl9x6HZBH5e4uuZ6Va+0IB8ForNFXvxDAO1RMoJUyw5uxepGkejnkX0lzpZsAm
blCGnCAVScwYd/G1jX3fBtOw51TjYuNSReHte4/oxUG7YTlNoqRcwI+ZA63pz/9r
QS/ayCDt9gTeOKH+/BHaNHiOAhWItNoizXdOYc6R1QDH9nfoF0H30anwatekjRyC
NreuA1gTwIuXyBKY/4jh++a46hRjgFXv9yX6p4Gci7qZ+mnHLMSf16tdTy/6q6qy
Lo2Exc814YnlM22P49mOh0UoSY5xLNiwXf7REf7Mp4Xm6kSKjGyPr7Jy2PnB1xUM
s3tcbDSCOkImVE49KiL24mHEqMiwgpDMtvTnW02wdJnUIyiSQQob1+HIO5tPHQVj
pd+c4w00BcOLPmaT+2chX/F/e1f277isSUkGbqbaT3BB6ax6XOSZG05rI6CDrxK/
0i9fWXY3riQID9B+IqJpTF0eg4ByZm9GNuJo2v6tqlPlexkE4NDuZXIiy099Faa5
KFa2X02HPGgtgC0OlV3qF4QtO/rcGwSJDd4a7d3aHlhENplE4AdeSXbNeuiLI3Wf
6v0Sr8EhQVhswMTbpC6ZLxSU8R5j6L3nEFrpom7ww00X6B4ArWs9+6gsj2/rJv1i
GdWaXh8LQuNCVBYNzPQ3FJ4+o5zP3CpUB3LxQmtJfkkoLKID60SPPDs2Z6BqCqmK
pnm6S7lHeaxQmkxYDbGBruB4EddvYAQ4qAKsx5rlxUKOVcwctIH1zV7nGVdJlYR/
m9Bg94k7BxOFBJLaS7yfZfNURwghOppQGXeNXNuzGZq1XMfep5AZQdlG/z3jHLw9
b4GwBO/+OuCXou237DTeHWHA7TEdf+KQspC7fs+O74th3Bxoym94RPVjkgTTvD0j
L06owDjNLBElzbBGvFCXMJKBAz0yWhak3+by+maZl2hD4br4Lfj6qEBRJyw6zJth
5B+3Xq4rG/vvn1p/VB2wkk9IuMLdB9vxy4SKcc3ioMaxu6m7hr8WOGR7J08Gggtc
lE3MUqTbUy0k6Sk3ZhLd9r6nn4+rZnF1B0M9QK3lh1XAQxIGOln7rbuyrUfI0po0
OcWIZv1P8nEKSfnYvSeGE5wc5ELogZBeN7PL42Vr5Me6gnsCVHTukmpFWTssW2Qk
83O/9Q25uoKMRg3jLcwUFvTnbsynPJ3Q9IFLdjp9R2W/f6XV9sOO6yLws0n+Xz99
n7ZovTJ8mI0aiOZsUMH1p9s8TBFX4qk5M+xV+SWtz2DA+HUYvxqEYyILzaCntnri
/TPANmD1lqY7bi1bvWVsB98QdAQ/WvhGqlje1voUcMH5ZUnF4Z1frp3EdogNkfSe
6iFFcLsydLn0WEKfFmJ7Yqi3EuUHuU3XZ6hVC5uwPmyz8UOO0oEkwgtTf2TjJqfO
geGzXJ9IGmFzqWJT/afx/mTmOMGzF3os8+tTBV/Z5T1x85pZjwy6yBImNOZxZbuj
OtaUDgMBncR/1791og1tFdRTAvcTdZFK5QH0OrrlB3t5Mgc4qdI4yqiFePLmOTlE
m/VRS+kRuBF3Srv54yE58IvXCBHc6WchZsFkyi/4CZtC75H3US5LccXRjwVltljH
XF/NYL9h6HaWGutxW0cMTsaRekVWNsSltGkCGRPTgylB42b62bK+16mjGnO4mQjD
1IYaFazIwo39QMJ3qSnz1x54eoYu0yBXqXJyBLEmIHXB2GBgX5zcZox4KpgM/IKF
9JakUSzYOb+gWrjz/tPy3XQKio7ZMuHXvIv9DFLLNammbVQniTVpqoTEsWVrv37O
2Fip0ciyH9AoEEpDHxAS8Va9W00Hbfieype7gLPiYQflI+UPlB1hrT3I30B8aebU
948ad/Lvu6ArsFVHFgyQFME7+jR8eK7ePTm+/M0GhRty5bWs+taNnyMTWVuGAzUt
DeNtMD0ncR23L/YuoO7HMInRh3bv5R6GPEGpukmrG2GPN1gr8hMsUUn/lBI4ETWL
Wl5DRrkrYe3IiRyTam0dhyL64EBu0H9anZjbOmpIH8KhFoCzxHce4WWpZulxZvS0
RMOYqUfz16WPjwQkJgqtJp4QINHf4qCtXhNiVPGX9pOfcxi1pk9sbIuaqiQfOyys
pDSjbJDjwVGPZLGUAv8qY41z+zRal8xQdFSM9Ryxxqaw67p01TzFZyBoorvctesW
mjvn/LdyfHrnbN73wNTCSPw5+wR/e565uQOyu28uIV2jNFOwXMv0QJgLT/yJUKOv
YB92Ni7/3q0wgiu7dwowQwdusBHmcPvQ8j6vNbcwoTUgNOIhx3BA9pcfF0Z/viBh
pbTLplRBrRAXORtGP1YlES2IlEcbynfh0bgyLDed0O1Jcd3JUplKGiYHrMMxzdVS
1aEoVWhBX8ozgKEzDUUZgoBUfSzqyBRmkrl0J+8+NCUv4vTW+bYz87TActdUEyg/
mO1DkZAIpXHSmoE9PKDV0r3snF+Tmo/Q4Lez3yi6X19YJ8Up9pQm1PWvhjXaSCO0
a9KOjTSKz+8lDgxiCYac0IHV+ZdT50wmxknqdozeJ1vbNX1eGZdeYWKYqgWJXEKT
Qxx3yb5TpkGFkVdn/qe+UdZ5Y1wqq2nykkTSDAbbHu5K4CPtI06OdS6r7wxEbfjl
N6Pa/LOFmP9G0gRFGD6Xk7+uJBcbSiK7HtxcNNA4bodDG/nr+jeRgNvqtNhgA7eI
1kfv2oy2xy7Tdr0sRUruxxrDM5JrGAP0txkcGpG+4I6+i52i5OHW+p93iOnmsSOe
Q7EAMEBu9IiOsrFPfplwjizvgXNb56Bwg3PGJ1F+xq5UNI8RaCDLm0uoCjtsyHHy
+aP8h9EyEprDaTj4rSEBjiEJKuFHiEIZj4WyjaFZoZjUx2sEstWIZ/0X/K3tCN82
+Sb6+f0d3bceMPV0VNAGcNDEqMRM4uqu03IQjzKwdVPZFET4Yfy1vHbn1B9pXIOs
oI9Qh8GPysKLL3wpnT8FTlY60Cq6YtOISXLRam7v92exOmtrl6uoCj2nF2GrNwEQ
fsiipfoJO2eSdsvm3TRn1zfpZ6ECXCnrdjWUUnfsSxyfbVLcgqLnUUNA7vBJzvpY
we+GuG3vZSLmS4fwXk2Ys6kKBO8uNQ/IUBMUjzw9uzMmf0Jz+AOpGIxKSI/PWk87
j8stA2prRQu2YEKk3YAMtNHjA+fY+hWOl81NzabsLnI0DTbeYgasjE8vG1WIIcCd
I3P1QoP5kDN3YsWLMbewjraVPu9SN8IeZ33S/D850OcA7RfQZmfzHSQqpUDXz8+7
vmyO61Q55SCR28SLpCM2Qc0oQYUWep6qx0XPAPiuF6iVi3SNnBw4OtD1uwjnK6xj
2zKZF/EyiNp/XzjXhCJeqtpQkS9rZv8HsBWn2y4yN8bSLioDWNV0BG+t9HQNxZxY
QprkC258OxyGLA5OCp1letmzblIGJJaPgoXZfkV6erXDJLsN153IucNTIQeboXfF
Cwkwsv8Q+8MQ9SSd0/P+fx+ea3t0LkqjURqIrM/q+qzEhfRWdBrO/lFWdHlmpEFJ
NnUwPAsWzvbfyqLlBRgWoqf2Bqt1P7nXkRHwKs+JOk1QAKkKKy9zjMQnX0nUV8fX
bn9rXK6TU/DQWIEEoD/xIH1QDOrDq0UOXaCFpH2WqZjx9enGm6IxqvKKujXTy/bG
W3mbLXfl4Pj2WDVgDVMlBF68cDIzWmsMwyE3zGNx/C90TUFFhriMYZwaG3GBpY14
Se/YnZGKzkVzgaLNRs75mcchFRvfjW3V+8knqvPsy604j166ue+Jf7cKw0ttEjCn
6is/cPTp1HcefYK1NM+8F9avmylPSUWfFIq9FTe/ruDFp1yYgnq1R1toSO96IOFk
avXIC8sazgVx1Zi5CfFayLhn92RI5JZnSqg1zi4lUDge7Q9Y2FK7AgC4OsLWgyn0
tPotSgnRvW4JBvYtGIocrCl42rQnerR8OWWwJDFKDA/P8UyxbQSfgVA/9K5pKEFX
L/02ieyVpw9ravFJ8FPbEKzTzsj3YPy7I0j5kBCNV1uty0KKR4gsgD8RAsTBu9wN
dI1SJPwaspxHTCLlDq21iy6mT36qppmp7YY+qPE3hOhumA2Mcg6R6tyM7vAbInwB
EHJHgFkkjIKjtnK1wdX0NFnNeN17h5boFxqDcbVk6VBIq/c/Kf/Veiqbfyz8zV7s
jG7ukBXmGGz8Ul6e+rHDoPl/SJLsFxDrv3o1YA/KxkUQOo5BEQPTWsKpPNj3wncY
FkSM4fMg5GQsZapdup96Gv2kR6jBO1easNiWFrwl3v7u0EeSY37abpkJR6QiUhG/
SEcXz59952mLd2n0ynB8syiVswyOgLMTkmTPY7lawVYHc/N1QDjEbT/1wwHTzttU
I9Yu9c3yqFDCmsBISGuzYpbvT8UUpxscvBBs6Oe7qBcP9q67eN6h1aWD8IDee5XQ
6X8X8qelxroLBW/6mcWgtepS9I171FwlrHg3Vw6s3cln1NMFXOT/ePGzf6xJnzOn
50hfgawU30G7rNhJJZCR9/Yy8HHMMtsxr4pPH/peGqF1DIkxLKxgoqzkZtRZir6G
YnrAPvH8NQqfKKnVQslUzkkz0/r26PM/7wlhVy5VUKr4xPmj8oGIfH7edAERB0Cf
PKeGnSPl0w3f8YE1biOZn2qveBXWIeMmb+THYNocBQASj1e4GVfYpobiIlznNu+p
bxKPTEmy3u79kr01N79rzpKBwpFF1NmKUqBwZfHSGg+EnCbQR+XRm0H5tjXG+fJn
9Y12/G/s2th1RT9TWv+5fPBi2PCNaffVIXeS2vbHpcLUcoOq/5BZDJJakBtnDeKm
OGIqXWIxflwhecuUI9MY/3p6yQ9NjYGM19g7nS6OTyqSa9CFuwkNkec4fiDHUNPV
u+2uWLVGZ5nAqKiKNk14pgoahLeHas2It1PE5m7I6dRfZI7E0Cw6zCtSS86bBalV
0Yjg4OL3Qv/b3ASa4cZ2MaU+Y7mjPkyAxzOkAtJrPUmcABDTLbh+JwpdkAiJysFx
2jSwv5pUhkxARN2L89NpprwBLNM0NZAaT36XqDdfzNhX19UjDAnqoRwEAw8EdfIj
NM1StgxReQBLqiePzLJMpaAFwbd4zp2pwhbK0VaElkJgtLdTFWSipwbg7vUZa3QK
7l/l0Aif4nuofS/jypYCBay+hg6fAn2Lq/eQdJCH2fBuq2iVylyeblTS9HAhNt7l
cJTRRk7al0yS0x5f/WhlEI2Q/tkQSte3vjE2jMS1r+8PTvPAVuZ8Ww280q8s0g1L
b4daTg0un7cZrf0q8Ywf2L42ghn+8Eqf52JFVmVSFU1tAi5tJ7fp6yJ/zX2L2LPZ
DYo6+oj7Ei7LE3HR7FBjHx147kCjVJT/l7qVlWbtHTE0sPnax/BejtOz79BiYFp+
KycHv4KlEmA8r9D1C4quYO2QfVum+UFHHKN0ht4E2VtShjTfjFl+KnaQERk5kfcY
V4i8fHQQORhtLFTCAcqIMLljvELU10lUAkMkCp5HxNSzXqvVFo69DF2kU90KiVRx
S/VUZDhn4un+WHg5z8O3z8Yt9U+8W42hKS2LM36MEBN48BG42gYLFoXgaeKbLyUI
XlTj53JjqFFnRk7oBg6izXh92pL0jMbgUQPnrPN8XNUSU56lgclYhNCRiY9mI81R
ywWHfpeGyaMtz31LakLlO3OKDenWTzk+v9y30FdnpqC5FSkVv4aZJUiPJDdxSJou
lK0eQlSPmwjHH75eg5Q7xF1HZddIiWLUwF/WnuNTBE90OVcB7Xn39PY+D4vKqxit
0VvyClCM+DOc//eXOcQvfecJ2U9mpt+jziaLntw3d+m74EvXAx9F1Qtq5wwONKK5
q2I9UqkyGiLGrkzizVTGxtI494WWJrzVgBZdkGMtG3fbVsAhIKFTtBF0EQP/6Tr1
Cd7OglPK1FJJVGNxhtvqqu6adFIWPumFSnAkA8oYxSiUE50VhbvvY8PJjvRVtsSf
RCBnOEfUEMqVLzVawXuZRE8G99Z878FTrnOsnciLwLcj54sdYLcPk83pkdqrWxIM
1XoPB7ZCXNI7KMmBARP4KkY7/RGXbkiICKmeNVnOvuOgdfBLM2pDToSKrr/25DR3
AdV5FV34TJ/Y9IJ6I3oAP4CLgygTwza3nc971pil10zQ+UioDUJMGe9DgEZj7VqX
oLHFb294OYUnmfI0ZSmRYUiFlFSii7lbn2iqOipnNB8/zT76sZ8/ywDz3Zx/72be
zqFKJY37fvSUMibsrhYadOJqH/gaEHM5+pPN91Poy2/dY/1oBu9yPcP2/0Jlzlsb
Zzz9uQtoKeDiIjuy4LTXUaqUIrIhX1+Jwj3XbXguo8Jkm6yciJTbtiZtUAQK44LP
ya/C+pGBxSMPSY/dANTSdldQp1gTDauF+EkYijXnew9LwtrRNNzsju7TusgtELSF
boaU9j0VlLE072/bMa4p9y4zeYzGLMswvSUZ5tqjNNY/SvLjOKshRfd7RXH418DN
uTaA+KqtZP75BzLq128KqeTIHHRFAeLx/j/ogNQrzbnGX7rJlYV8DHakUvfGfp3A
NcKT4CLgKs/TZmf77k/9IBN2Efll+qbvQarp2z6x5ucDLZLsicAyrGN8UjiX/JqY
Nobm5WWXw17NvbBwVqnIYPdn5l4xr9rlRP0dKxZOeg3pwz89U9YQbhxtmEwlhXNK
okdG+ABX0dPgBggVOfj5GeC5LElSPa4RgXArwmYKffqnd0aBsBY+7VdtpKGhBwqg
9bKjV5hoOXAVxODBhUgUWHJRIsXoRRtEScti66MYtLVAIaKWWTy4gzB6BX+I4kft
MIEboxMPxvHWT6zmP1zA62HJonhe1uMej8vIA0t7PRcV+5ENlSzgaTErsw46mlDi
sRvBJXbOBgYI0ZFvscihNPBHbRII4SOuLGjh4XCBBydhomNDgp3OXs26/CGmRb7k
dYOFtPj4utz1MqbwYhw+Bkez96rijmJwC6xj6ysPYNdA8f3CxaBoccJgnQliKVDZ
FFNk6d112WaiD4Rlxmwcul/ExwmqLC6XdJsfy/MjRsWXOXIfo9RiRpzTayXCyZlu
0PKt4WZp+BbUfs7C1g3P+k1gMF8NFJ+vzd2v3eA9FpN1IqM5icarCBAT/U+bXBrM
p5cuhHNBQrTGM/+0jNeTwwt2IterqxsLQYe2xlpSQUbzatJMmEywF7vPMzSF69F6
NnCn1d9pXV/7hbd6H19LGyJ+oXAQu8WVyGzCHe7h8lDb0WVB9v741FFdS6Z3l475
swDUTzGReJt9tE+E7s/cS0rqOXI47t+F5dZ9dJ7UdzZ4X9gpykbknLjB/ygQA6Da
xJnhywfd++nV4IM8nXVWuIfs+NkUgd2YJOXqk/6riQryUZveMmpgSFZT5PYEavIN
NqOBPr+hPQeWWrHx4qj55yrYII+l/9ef6LX7KS2Ox8TCs6CrTZydOpFlC8ovUIzA
HxdbOEQxI2oqy83gmSEDxJ25ScMIp4o+TcARNTsrKiNFT49w/sgMuVQct+AMozHm
MrstrWK/LmRQiSSaZJVUPCTrX4VXWdqaqDwM0Utf20a7/5J9R2MOzy+uoCTAZ30e
gSMx6nHe9If2hPmBN6zyXMdbZ61832bBWV6Coxx/MtGS/dRJJB+N9gnuME8kDkXa
Z3kKZLLDFI5uCHuDtFM5V7ppdc36XGOu1TBdEE9UjHCvsGOUNLBtnsuC/K2TAzwG
Eo/UCS961OUQDVgBaLaYwh412Akp4s66gaPEGjRGm/cpa3fzppITmmKD185Q64d+
d23QLxx917wVDZ+L0iLy7Dgsti2aQRG/CcxGcbB5ne/qr8baAq8oUh8LUBMklo1D
CrcKXkKSRS4rN0J1pyM/IhkzO07n8p44taaBta5Nu6hd4Ui4fn0NwohSxs8v+VOx
+V8JN+NIYUtJ5I3Jy7u8On6T3tMoZ8TDTQ72AdCeLzXNaw9SaMuZ9Msd3zxm9vTL
h+zciIzXCe0h335dygB3NBOqhGTlEWFvmHwR+fB3HOpjnXWFA7dCto78SePJLUET
yeYcD7FexZPz5ao5rMFODxKwmKzQ0C+46VbtwoWlCLpWXD+yR0HbK2h07PiSi3aR
y6JO/G7e3Gc42JqgLCd5w4+d57y495DNxfMnrx9aTpljfRM9WDM5GTtPZbZO4ulE
068USunkxbtejhdNmplUr8An2sgy1g1OCf7Zzyt4j83wvcky3fL4Jy5luuyn92rZ
paE+YcKpp6PQjagx40aCWOxr1h2ZOKBojQhdAsrSFjs0ysZHho84sv3mrsWfi0nI
wnEh+edf95/ydf6Fr9Bc1MH5aMaOS6S3Eoh4celLgJCTtoDxot7j3kLOVzOuC5f1
OH3/kmrY8DqjM0rWjXA1yYOrc7nb2X5Dt72aSVAbXMerEAmnYwcULPxhEeQ1cGmz
3t8ScCrmay9DfbTkMuSo8o2IjtVLTKIlozchLvZ2nefv0T9uCbcfzfByRif6hNJr
VK9YvveBvHvPeuv/p0iPTtwxwHsSsKpl9Gtyak2p9bUAVjQ2ieschy+qjmonmyei
JaJsIhITofdTKmLvOekEeCnbQshNna2opGzgK8Ly3FlYGrqzjntdfjvWSlB79J2o
YqgYgKUe36HYQ1USqw0m+CqAYsslSCzPQuZmuxdOkEe+2+DteERhNkkBCJdeEHvp
cFW2V0rn+6XS55X/dOKPZCzdzluLUG9rdGErO8guzQAHAHLadAebLPcYCu5BQwsv
f1JnZQPs+DqGDV1N8tZhiKQxRk7x9TdhNBAtTOOTg5NB2hwPwa8FBLATK6DOCJB1
wOdyV2ZGyTi62hNRx7ZO7d9L2SqVOhRSidw/uZrRstu9pI4HYTfE8mjb/J+V1Hxw
FJEM/LUStf+KzsWz+sl2yorwddyA0NfuJiRwr9/dwVba0vlubetahgDH8b7mUA0Q
zWVPfk+WeRawWzfYE0TGjT1tAVCXcy5o6QNCUJ4UgcVxzYqsIdVwdPfTI+/+NMjF
qs4l4j/Ddn25igz1VWXJRnmx3xwcIQJmTNedQO+NvJpZuDzKmGQVHEDLjAd7Sqc9
/FKpM9v1RgPVkgNx7dVyUjWp8ZpKvvEBR2EM3WUDAhDARQlowf/oO5FMobArTxrE
X+IVn+wBBTMFmdGtaw1lBVN39yIS8al9EaKti4lOQExZW9jvtSYLGXFv5p6df9d8
E5g8edsmLEwUY6XqOkTDsbNiQy1U8O3rPkI5nqbn30sxj3jSxPES/zQadw5WpZlq
60rxHEuhUlyJcbLJbYFXddQVPMKnNbkI2syHnReBBd39PpfROGVcTT1/LV4Ifk1r
3OZpEachdkmAB8lNWMKAnGKm+m2nVjPYbJGNfrkgL8mpW6ZOspMxDLcGMOhInB9z
34siTXSEHkfkd5AD+fosE+qtNxpERHRZ4AcQPGXhVgwS7sFR8QuiRRRdqhCeE1V4
3XntIxPYnIzDx0L8xFbwMeRMtRGd0mFbGNImWQH0eVvDxNO6F0z239sHgqL8DPOV
awViWbiJflOVUUyQ3tFMmVgsxYDPnngYvM+LgUvJzKuYuRlCxb008HnTnWalrni7
dNkGz+9xhIs6ooaZkUSeT/dZ/mU5BjaWtpb2OZLuZrYe5FTSf2L7heFuJq5xCz2m
I27m9Qv37z+6pbu1IGNqFJV1Yy8bewz76t78kUVukSqn5okBRep6xchL4NlSc4s0
JdY0DLj5G8c1/BYiIuunUe9Md2N99aXngO04vVi/G0BgpU/LtkImdIxUTSDTY9m8
rv+ZBWftTwPP8vuv0GKknyVpiyUBcP4pgsR7LH6gtZ4ZphXqv94hMqY5dnctasih
sBMxQCkzX9FXDJtCytTjqkLirziuaxn41bmtqRvdYUG4XFL85sJ3ER9FDS3Vm/0M
7ffu29a7cbinuSUdE5NO9R74UCozF7ctLfn48FcXSR0GQ80uy5tFYZNbGkx8On7j
lotDBVemnl6PM4pRFg8ThuFACt4I066mqne86yTAx0tkUc/iPc+TgnEFl/KgBA9q
/AHPj6tXWoxpChWJOZJ8Q8ifOctP3080gBm7azvQO8YOk86E7K/bdKSZ13QOtbV/
4iXphazYYgLUTFuH5YJxQwCQ0yQ/LgKefHAgugmeBIQ0clUsJhVa941AJ37oV9Ng
jq9z3C/47tb3O0dsmBnX8xFAhcTMqr84DFrm/CZ5KkY5fXHjbERvAaZS5qmKks/d
Fl2yRinzOx9uoB10gRhotsqPN8IJ3fk73WcGCx3L+sUZkzpSEd539ePO9J57Qda3
VIu3mBPJezTKTjnG2XtM8NOFgoek/WEVBqbnN7plzoIys0gdlyzCEY+HkjXW1pXw
VgLCPyZopQWzhKoGleUxyYxOA48ZXUNWQ/Utw2te+/WoEAHHPrfxcbDjmhv6qVi/
Fdl3b5V3/c3ATe2e7e2uaqL4OsiVO7ULLYyxdMvg4mWtOk2cImA9mK9vnET/BKJZ
TwTf6bbaH/0AeW4OYHZ6z1in/hBiOClVOuYHiWdxAXb8sU0/xe3xv5yeESo5IQdY
/0utFXNPCxqQ7DckPvJDliWyEA+j9tGwVHJYo3mPFTr2aAvay7jb5mjjPjpm5tOu
U4AbHEEbN5XdcysdRhYAL/rTPnepMLK45nm9lLrbwLtEs+TQ2GzJZGgekoUUVF6d
gclT//o2PQ2dnqb78WXjqxESw7eGZS1Ct7rQxqHjGi7XEwySavZif+wmG7m3MeMA
QtQYTjc9DOOP/vualNGAQnP+vAmkUeCEgCJl6Gsn+rdVrx2j8YEOADmK0y7WcaIi
W6eMOo72KHz/PIzdMjeSWpxdFzMGoCHNyiCUlXiJS2qw79DAIM/yud46XXteL0yK
a7KpClYabKrkRcuNKU6vAJhKBOSrdhjQgS7LnBAQvyB8t4bwcsMJlgjY2eMYoRfP
GB/N5/qV5Uspwxpdi/P0JuXhURqRskvlaT3WQgC+EQmijjHX3WfJx4NibScy7k6k
U3WacUzDLG+RT6j2IwUGM1ipJ06KaNlctFgSF5kc//Rv7Epkvc580E/aYe1rwm4G
4hymlT8TXlsjrXYRF8ZqzMjDTvG76vLD/VVSydIr7GzqXOo3rXxLLTi5bG5SU3RE
loHWl8vbbfMjLDKwCnGx13mg9xt40FFiGNZXTX8wmuLw0JnMG7Vr3DY3WHGvzurB
OExRsq+5RsB84+AFOlT7MdgfQ3LRYtGgCGjN8+IrxnIZBmW4YpYsWc3kdLVfZ34K
S+BO+PtHLI7ELZdBa6A+S+2PwJoETVcRWzMHbxRLYF/PJQyoyum5FYbGaYUBcaGr
VSyAi5S9eL2yczP0wYOB5YH0r+VjHgV0JV3Ma3RzfydyZBebTAWIm4uojG5zIRrJ
jZvDNaS96N9avQlSS1Sepi2xVNMH77kQith92+f1nWTaHhk67ptLefFKyKiVc7ci
tj3iPeLzNOw0VlHqydWbZjrrhzqCPv+4n8PnZ/867u2Jx8qDpFOo/ybVNU06HUNi
l/K0VNRWKHhPGZfhXM0tSb5urnSJ651JZflaCR89LJky9pAlOPDcECaxK85qsbVr
wnMR6vTT1yDdANv6OfQhwbNc18wkliCBjVMRK7Oy8lsojELqpxn0X4KheCicHzo4
hlCCavc06X8PpzXMQNoowXp7QqSvS5iKHu+UXVxwkWtVswBHIg/AX9fQL+UyLjRY
zy6ebjhpwHYNaZa1GROEZu2biQcdRmaWvmg6iDFYakd0eZ63N9mfAVMfqKTqvQtU
7RSvFi91Ye1nX6/U2/FQX9QFuaKt6zZgL8bK017og6CKQtVYMyAZ5UDC+pOec4/S
5PrGDdtBlK9T1BXBBLrUPpPA6c2QwBSoCIE7XVhT71GVUU4/yjJFKXj+7obHb2yf
pJ2OPgxIPS2N9I4DX83kTMkXML2mj+W8zumTXdW2u1RRpHT1DYyG+EEikFlLJlNi
aXf/QTE0+E6E+MA6BlLxkMPegJyX4vjwFx3MUGoWnIzvnsFvJI6dc7dlXJexJYuX
EzKMqLe8WNbrioh6JooC97faF48gg8YdiJ0PFVP9oMoWpOBS062W4RxBNfPS1oCd
il7gJ7is1sf6OSRYcZf1j/IhrcOzK9QOJz2dk0s26AF4GVb+mCwvZeTGOAhKbvJC
vij26hPpI55f3CUadIiCfmNVMyA4LsH9nionOs6T4JmsIxncS7sBg8j3quZ48w8k
reZxW6i3YszTpiAaBGFfTE0w4nf9gX1w3Pv63WSoB3ZQQqBDdbtI7OTxBDHMH1Ma
ybecHVT/Vum0fC06uQHJPANHvx28HiqA91+CJ8T+AUI/WECC297IIlNidwv53MT7
e6B7TKkqUitkHy23JFdpqRbYCHEbJiZThH4OqSAFv6BsOjDT6It4zjMJqpw9itnJ
C/J7NXfrMHELAtWAPwHiPOoyLJ+XaXUcCRlhyxbCasHIFqpiSp1mVgzfYV5UYJ7d
OHdJ8+L8bl3Q4EivXj5X3ZA+OPxuJLbxFYdc/hyPelIq4gCrGiXxLtqMpvPggg1n
fKurz7xM1jb8w8M0npG8Lk4nLKmcKjP8XORN1vrgQFEzwraMfLztM1aOn1hW1mbe
Y9HLIxrH1nsRwjKKm8U/8wIv4lw2o7d0Wptz0S6tDxluieJQNP8wKarT+KXBCISK
/8cKQ32qJ5tma1QuQ2q4NYda/fpA+MoOPdeB/bjVU0FEMlHwrn9tnG27UThXHcN7
u/vbFari0K4liEnzK8sZtVtlSXqvTCtEud1s7ImVGghfxgolzp8loaqdW/tyU7s5
LGGE2sAeLQe0UUojiHNotuf0/gY91KUYSCcZbMnIakrX4lA1DjoVuRUjJb6yx9FH
u8k0ayZUBlmK0b3Ts8tbwacw3HAgQAjNKQfkCc//RyyfqSn4cjox+patSiey2s+I
f7XBlTo8SufzVbjaP3+bb4GU0GylS2Lpe503p2GXnrs+vTuMbIkQClKX23XTmZmK
F1wOQr5lqiW5Xlqb2hwlzdPd71Gl96Q63qYDYBaDL+Nq721Elv28gRNJGW0/ia7M
wgcShSXeEm9Y6bGvUUxHZYnrJy897c5kfyaDirRTtH4eK5887hJVkriIaXo6QmcL
AHMjOtgOAKBs9uLc3+C5qrC2E63pWg6Mz6otlfYFQ4YHVpt8SABzLdFud6WpwuTc
D3P0kNOKNVqaU5bzzW8wi03kodDo5MnRJ24fW2PUjccwTmDDltUli/8lHPz2W2CW
zkMWnSVOvoTJiLS30JorGKh2JltbDTfkg8gusXMGQ97mVMjoj4fXFZhrLuU5ST0K
9u2IhR3x0xorZvAXcdR8u4zW1Y9gVfhY8gQT3HBywKJ1KdpGHPh5CHjyeHGz5ROx
R4x8L/RjoB/90wz1HtH8Jec0KQ+FpiWah0hQoH6+udjqW0CVFWf4oemV07yh2TAZ
bzTgEebUVlHp9hkbDt41gsvf/MQBUii7YGWGIBIT2ziCi5Eu+7mvDBbGOmhwGVNW
TQ60lxHe3+2co6moTQOrSzEFBDG5NC0xHXDOQCxeEcKyNw3CbnvD0zkxik2VF0QW
wDYo8Wk5XX0AZ5xEqmjWJx6xDhR4hIvmbL/w2APsAdmDzT5f3WrYGqVJ9979UOHM
+ePMj3pmDs8+DkM9VQQoEr656/T9POQZAk73CYCNfpOB8NC7k4APHVBgKOA/DZwY
hDhpBzo70S8mQMb2G1Cboj/xq+jrdzpri5keZephRXCy/vDdTbJSv4+kP0uS1J+A
3Exst2/YvyV9N9kD4ooyGaM/jdAxQyo0YW3UoQNqZ1njLFwXPhbn8ZbaZbnTsfjH
U3LX6heCYA1lBaGdUsnP1QbWzNTud176UnKfsIeReIrcy08MJCQbev17RuZ/yT/g
NNI1OPR3VUAfaAaaXhf63ISVd0Mllu76R9RnEGqs4ndW5XYhq53DPTT55gwlvbCj
o+Z6+Y7jv1jNhNmrCHHtUnO1N10g0z6twWj9p4KsFFTiRt0AMaAyme3BekHMQVYK
zcXNqILlx8M6fMtRKY1hbk2DeufjlrAAHNPH43jNAnbLdVZvu0RPCE3QttnRMYSJ
hN7DYEs4T7q6ofu2haWcEGA6GoX/iVgNzlHlEoCHePK4du1ENsCPksoNYH0H6PD3
53zQ9AR87OlmQmInbk44rbVMdW39DsmBp/EJIM2gM7m5Qp3RxqewK6+EEo6LWLNs
cqxNI01uWX4bhz1Gs90huintKQj0iU91myyJldqEeIFU9AYxKrOxE8ncfkiaF86u
fYn5h+lQWre2SUYourfGmaH0WaxGMeZyKSQzShDqh57YJN0DxljVK886U8ViiMbq
68tAtaQhKFst09PeKXt0QI00KVDQefN5U+uK2aR5iuBXMV45/4qP+59KSlxqRUfv
pWAMojPDce41jB/UKFaSniA7iJT+wTgZy6jOd0ZSH6ucnCo4d/qnBfc2WKKiutvx
JjVPmQZOvDkme4UKHhlBAyOMhMVOossBm1telg4lYDls2ic/E1mEfxLZraqHDcA4
qFV9DYxaAH5cLddOdOC8nSefwGgOXhIvqDWn9PRWU49z52cxhd/+dwKX9ol5GSwH
c4c9CNlHW0UILALwnnP+jfx2f70q5/prtiooO0OUGf48K1lnVQHwJKlqEoN2fOBb
s3UIRdWQ9zGDNhGrnr6bucBiJhJ/N0KsSIS82vY+SHGm3NanaJguEcZcGfTCHyGE
y5d1/u/eKisCLIGCGOzZ2kQ7SOA+ED6f3Ck0dySi1Uz5q0TNDaTpigTAtMkJPrkK
/IbtrAvSud8iRUuwnqIGEPBSOv5surlgICBAECnZIEqTzOCdd+XgE8W165mpTqcM
e4L/hNwbFaNXGAd4Xl6ZN/xjYTWRFUeORJN2oY83Cw6GQD3H42ogcWwM4Vk8Egv8
w/LTXyrsdI9wrFXxCqyCPG9g5Mek4cVFz5GYjbU6HlI12VgsnXUtzmByDjeh88Zh
AQHL06TwB4iJJAAUh67Cn8KdHoFkw6lpyhBQyKXcgBiYUrgSQQJOAIPtM2/8e4Ng
cyyn1VkizPNyS/ToiH0Qfqiekj4LgKAgjYmqSrgzwMzck0Xz2Gb390X0so1/PUXM
iHwcV7lNze5diXPAbXu1lbEdSWOUJBPsInzv5GT91HpZ5cpy/0uohJXCkd7HODFC
71fzWA0+6vdDXeTwMJKRpH/JhG7ASF69DoDBkCgefmtbsLm81+bLPWj+1uMWVBrR
hG8shnz3iBV2UUUXmrJMOog63E1BiWGrnxvI5MsSd7n58/b9YVjjYS+sR+HZJenE
WgwvSj9eJ6baBXTadUuFGJ40rEvUo5GmfDj1qcBz167AbljFBL4qbo/vjm0OJ2/P
j1ZJAiSSRy9T1sfIjl2XjnbjM5oqesm442PpdcLYN7M8CjWjAykhlbyCxK397Lut
8kov/6B010623qMYAG1ILHccd5Bb19LYWjMPY6fulE2eFOu/BAZ9A36vhwrBWPXp
jl3sFr/R3UHqgVzpIxSsjD7zGS/p9VAGxlZ8Kqw80wckOmQsgmvQWZfxATStA8Ny
C9qVgTRiWmMVVCpz0NOGp3PV4/Bjw10S1k7ZGrbe2MzO8pbQeNarwbWUVdPF7rwD
ske2kcqaicIKcxfkjh2/ZQfVgQrKkiWSyORJKNefv1R5mniTi5nBM0X7f5CL1o7Z
yXzVSvt4D91otCoSDOu7HDSa+7tZ+GROUf2aEJCYmUqCFVRRXE/Zzh0AM1fUDzIX
3g17fTHm3FMi5sez4lQNN/Dwa9XxAiEym07fGrZEHk9E97f8uyugay6l9k99HLjl
5V5C90y13ULnOkHG06lXdUg1bWNdR2UDI3zhgz+YHB1qii/x3IABT+aW72+46hW9
JAi/vp1FVLDrHRKKN+yzKUleWRh1+rZ3EEJ2DqLhoWv6sXbkDjNTPInQE/JBGiAI
ODNKksSu4TfemH/jjjB4XiEQ+h4iJCnc6Us5rfOsfJl/g+7Pp9hEjm0Oz1btYqy2
xusqpa+eBncw/dnyqVUPnlr0CuxqL76BztwXjkc+j7axpmf8HMhYpjHoIb6ZziCh
RKR/QJ0YQvrNZCohUicexPqchA+zN3lYPPHgdhu6TswlKfR5PrzTnZKjMfzd9MMn
OhRbt7jyG/21E44icqnW9+eX3QExV2c6Frnygs6DMFuNaRFhTtkNxdV99VNhyYXx
BF89UZAtaHVXLXmhWZ+uhWQnDvd0bNd2CUX5AUuu05A1Vv7NJ4Hmtnax9jeEW4rt
/wK9jameM9MKhNcl0OWKB8BcEifrKO36lhB00db1P9ujImvtMB0bFNZ3qoHgAkEH
dbhvGIWbjtdP7NO9WqKW7evG46Ke+zfK/TN0S1OadiGoHK/4r42pAyTy1n1Nx4BR
U9jIJE6jhTf14VaKdEDKdDRjltFmRIElnEFSBtpDbRFdnYCDbv/JmYWiJGYxV7gA
XU2zfOaUqY7rzA5mcxOnHkm0aHafshcr+1XPWQzDofUPsCRItyzICEQ09Au78f9k
zbseYFA5WfrpLDQcXOVXjKzlBtQl8WHQcSep3ak95BysMUAAYkT82zkzzRz7NPN7
EzXMEohzA9K37iq1v22mieyEKYb1YbsKQt1OPu6ihM36doRU2cwdBDgjmVCvKyBF
oXhcTYXVeqA3U2wUfA/ZS0V8Ur1WcIPaXYBK5uPe3wqPIYgogRsdl8L7uB18rBeh
i2TCMt2CxUUnDg1nUV3h/WaaQkWi6kJaZySEEqrS9CsmVo1wzultn6g/hMfhf8XW
6u/o6PScCX5QxHbRLuVUEnCh+KS239lQqOGJ54y9q1Ep04yhLf9rY7/DZC5lx3TN
CA3MsHg9VZxC9yfc9eNW1Z37lbra12noNsCD+C/sdVA6wIDxmLpOFNDWTa3J2/jQ
S1N1WOMhsg17cXtSiIqXFaOP1XFhKQ5eZHJ5QJ/+sZdI/TE9u+YkgLvGgBsyYDY4
lNmmXFdnTEWfyTre4HK7t7TJJ4wM05x4tvZSWJNmvv/1cvT0yaH2/L3+5VrdSrIq
QvdOkrwRW9lanEQ66fXhjOI3gXZYQBM0XmkiPoFhMfPlh6YEyjID22NuQWJUrAC+
i02g6V+BLWt2TD6UWH/tcIOqDNLtoCg5yKSdmnp4pEvGLD8aefS9L4R6z9LTxQXa
KHlHfdF1Y0kMBkduWRZyGRqbjBZxvLMnOueeYThlo2wfUMrVOJYFkgOWv7VdGVlM
+LWqZqmAkWM7Skx/tuRixKsR+ouXhMP2AipHa/vFxUPcY/avnZEL3ILnTEhMfDaC
5WKHr1Ok4yhwS2xjjSsUB6ubuOtwcYsOtsKZ05qx8oA4l7MD0NrHzuDvpvJwrv/y
E1Pya27s++5sDsGiZlxBY/QQmuT1AbRtwXFRycUGX00I3YXI7bld1ANZ6InWcikZ
AEzTrQH5I1WZN0v4mqBdqjAbS6qh+UlD+lGNooIzgi9deJcSc3lfr5OOrSmYV89d
cUgkwDb7MZR7W454tpFdoDIx4MHATpcj4phpaGYsYtw25pSOaLfANIhlQ/ik579f
TSCph4lS/Zk4zjgyK33CiAaMx9qH8Nlj5RpYNiZ3ZGjFYKo71ALoo/nY9a11Oc/n
PCAadjaZsVz/Jv4C7Xs+NX9xUhNEndejfr6uZNMAN/WUIiKcHZo376V6r4Rdva9B
U7g+0iJcMeA1SSUpub2g8+Ib6OS8QoHfr9aKHofur7Zl+yTQmocC0ymBqioHmq/d
Z9TKTnNXP3iBf8sNn/PdB6KrpFgXxIDGfqsmBh2iLs9XD7WiiQly+X0npqBNPapX
1Uadu4N3RAG/KS6C5COY1G/yr7nX5HMvM+CPuq1tUK0e+ez/YlEZE963g2HURR0M
XXbbUey4nFVka1fq7okymd+F/0tqBB52LB0GCR8C+Yu3S6jtISqRJSRr9OmYajoz
ene+gbyUAzm4LMzOf6vPLXEF9kDGUEmnM2h0Olhb99/a6RNK7QXSnAbkvS0lQ+Zx
K2ng5MW8Gp1qzLieTfYXXWENN01tZ8B3Iy3NPYZmZRWARcmjcsmuxBdAHatAEMHz
nBHevwMVBeyDgZQ5w5krqq4s0+ksTxS9tlJpvB2Fg/qERbADdcybvQMlWrfplm6w
MA/AEfizR2eN+ZA9wVbmL/w7QRJYrZSNLB5qmEfE7Fxfu6sR6uPJUn15kpIt8F6j
QeOVTleQQZoV8DNvh5znBofb3+MijlSwuRD97Nr4llHVWtU8y1VCygeS9llVBwKa
cbxD0P+J+xKW4EBeAKT3LTjbUEK4obSKGNpP/nRE7+IP9BQtfQcmsd6YdZjfkaXs
eJfGyIqoRXBtzPw4+ADp1exlMTpaBCEXTQGgUV0aP8NJSU2Ry9W4ycwtPslw+x8T
P03w0krqrNsbmUgoZrjrhfskcvozgQolkkpKuuwuWB0o38oUl+NIgwZmtvhT9djt
4pG6fIGfbd0b+s52htPDuY31VX1zn/dz7YJDcrslg1VChney0c3/oIA8tYAyT29P
Fh+6bJVPwwf/2Kg1xauZ2Hzs53Dv7wqH5smsMZKBGNxCwbrDsxRrTHzvuiKkGGlc
Rty4wZK0K55Z99aJBYyjN8nJpgnLWHrlwSylvyqCSut1O7X6M+GI78LkddYhd1FK
TL0Ff5BJLd+0p8bzt/Z5L7p3FYTVKWNJ0SFlfJxpMV/3Qs48fKl2sl7DrM6iES9m
0kG65iSAVBzit/0vUvTD4Y5litI1xbmV4ZBne9p+twWxTyniAW/CTFyJo6N6Py3n
I2OU8gxAV8UK6JqyQQjo9NSr/Qu/8AluYfIhfhM9DIMUXfHQy9hD0b+zl63JACPr
tsYOi1fyOblkfNjzH3xJgd90LH3VVoYeBIH2yzVH12yePXX0OxVBoCVgghdlNIvv
7IRPOfU86f8TmJyp/hyaq7ZH0KFMvmfYjvXvQ/1hJUQIRzJPIqHrv6dj3xV2hcYT
j/UqBlFv5pTk8JUZ29Stez30KTu98uh4LdrURACClxqa6eAkIvHP+A+nzdszu1bJ
lJovbhjnzR47snOS1l+VLZ97RdCwJCbzLO5nNg4G/ctUslZzINB7snsI20crlbCc
EeN/qcBV1iUBCTC/uko2M5JpK4qaoEtyHFX80deM5Xt78oGvBGu8KjzJ1y5dMgyP
C5Ga+1rWdVjptxY6bhQtxv9xOAmvWzO9GxyyaUxglxebpMg0M1gX+UUEYCqd9AQT
hW980W3bx1HBN0e/ppwHXAjNVek+gSaoueBwywbDywxyrFFfjRLxowe9Nn1r03/o
iPduohrlM+T0AiTH4+z6731DRrzkOMzVB+oejkW1CdB2ORGcmh9D07VCBN+vusKX
HghG6xtjBRrtiYo/c4pvBoHJY1Ll03pSFOo2KMYwSq1rCbRgTFNJYSoLEfSM5/2T
V3ZMHHc69FWLIIa2gu6ycMrYfBbLmhQ28ZXD9lTYV+ZLGxh6PM8T6ZUYKfk5bP45
1Sb5H+aau+EYpdRv66wyGTjeX6YMLWZ56ote2+R/g03HrzCzx/klryH69voHSPnW
2+y9A3WsD5x5fIqOi6oUq37Tce0OAfB+MgUQdiDe/GqNeYPd/jSVEFLk9nO6sQ7h
SQdWL4an45uLDNeGAJjHYyJ+K6aWlp1C2Y7nKj7PEEvR44KEd+ZtztxlTTg+lp7U
EpQDdaX65xWky+wnqD3fS0rX6PrLE0I3FpxUZ6auQHx6tkcRCQoXEfTyvI48Ip70
nNxPWe3H8BLG4BG4FQdDMlxyDhxDhT1PArBNLjHpKU+RuyXFhQ+j94Q8k8ETL6zO
xbZZ7utsh1mHOfQay4jq9uHIF6ZO2sqAtsrQvvYjsFctiXQIX7AR01dhroKXF5pD
VPSf/v/AdzYMNOV1/hsI5Nn2Dofr3eSOi/m4CuF/99QosQOs3QWqh8rUh8ODRV1Y
LL9qnWjyEIm8dlH5TP78tvYmRycWF02Tm9JEyowDNhPm8a7H4jfJPBletx305sKh
FO/vB0Gxp4v2EuuHsVnRF+KIvRm77Wl/lHrJsuNJJM6OIxrEp7vu6mDS6WZNGiZ2
/h6onggp8lmwOUeTviz1IcPEY4/ZGzs/yI8hqRDa2UmsXFiGpC+kBuL8nVydOeSO
s+JDog2X2NKZsR0usVxSKkE2V/Bfq2PFtIPm7rXWLKsizesh5WhA/kYmJfi4Gn4S
2UDkKOSyV8QVZerrc8o+eoWkKV+ouI3RitqneMiMvAbofjRPP94VGZzAHgLy+9CV
olKo6hmxcFZ1CyI7zAwZVh76xC/1gIoR8DMRThDFy99RnJc/LSvAmft2WkIg2fQP
vinTT2sANzl53D2GEy0WLjSq8LNbbV5g9RN29Tz/TfrGhH5eIFHYFnUZT0tA2wQ5
22ry0dlTrq0S1Xsx5sBchq+JyCA9DvjKJK8DkYF8OjfWqe/+RFI2d+A10k2eVE74
gulJY8JZv9BH7K2bP7eLGA1yYr6BU4kIgneYl53OU9gOjRQqqHzqVXV1Fn8kbXdZ
Ge9qc7N3232+QJY/DoAyw1KUcquabev4ouhiPgELJvjglrKkH8cNc4kyaYJE9h4a
ZJ7xdp/ciS1e56OnNHuP/ToVATiXtxktRL5X7mz9426/T4iGT4M4DN9IEvh945A6
3pbpio7h6eb1+f4vXy+UmANyNtuO3WKq2+GTjAuApE5TALXnPWfZzcwRDyZgeo2/
ocuVgAYnbwCoxSLyGa5q46J7ymMAAxyrC1WnuCpcAoZWL5fKvqoPMAvA+fEQIqEe
/DoiBesn6Rwy6Cn5WolnbOxV3fhG2d8Cunyn0evaOaPIxgiVmKnUMNG9eguBXU6R
wb283rdahrfz0lHDwSKNQiX3++AzcGL7tQbW3oKv4ZU7LzPakUDFgEdP1rtpkecQ
0skL+oQOkPyEpfvCPq89WGJAO6dqOfGbSAvV4wdNwvomeQRxluRWZ/9qaq7oQbsX
hL6ZPC01G5P+ocQPkfow/rH7fb7shjVmKeKZ3eEfJN+A76tDwzhrLRiDn7Chqlnq
jiP2JXpe24aA7LdAfjBbCs/LOPE8+nrHWM3OhDXKfZ9dZZxqLkmcbibYlugji2qJ
wFW6+SPayjmcqpsHOcnWu7aP6Ir//rOxarxq6o3FV30UXxOjvG6T6tW7jEoeyyD+
ow6O2ifAqR1a+ATV0vR7k0sU88r/lAVcN8FGAX6ZIZbJrM4PKf0ncijYkhq1I8PQ
nQF6oeu90bNQn9bOvfooPlDP9Mv8YRHA14b1JcX9OmUakcVWXGOPD8IKW5iPfNRy
18dVbwhFeGUGqt2d5Ln0ZP3otb7XvdI1laOXD/y1B7ThMb07A85KaXDIUu5Bvb88
s+gB6KFxeB6nC1ZSVSJ7Tsgc1fWO4mL2kBq5tqjG+Kbea8X1sOcX8XCPs30sWgyI
14sGjfaZDUoYMPB8RV140HFfSV1zgXsDV6CzTMiLKmq1l5F0dy1GpUmLMWQioXjJ
v/59Hax6bOK9FiXdxmvcAdxMz0WpbziskAkiKDTOkvZWS4lMm51XWgxReaehV28G
Y2/QTGDFHvK6rNsxb0jFawr7hzQaVfrNHgyHFPic+rDoflJ4lJM35S2WZlRFPNsu
1WVWtp/pBZStDU69qquCnb2+rIjik4WkIxBL3NGCCt6CzL44Amuq9StDKv90Zqe5
4LiwlWhq3S6wf6v1SkCvdEnoRWfQvWHoWOwUqnDaZECd0Ij/7TbZ/fIFLtc/3bFM
EYU5NXvhMDQAit40Q/Q+Ywak3nz0O8Mm0Lxks3x82W1FNd1dbdUy/0sto9rD0JvI
m7gnwuWxVGpgpkfiChQRGkKiBAPinpDUQWtV1Reg3WQYhmh9BMeAJUiwdMTCtiMo
SgWD/YJk6jJWEBXcYouC2g3utmuNOXyQcsrKaL1kDFsfDq+tU08g2F3tuwWTXaPE
zB5IN6/rzdpAQKODCQnJLKF3K8clV1iIdaAEoXfmVRsQ/oNMxAJ7CbALjP9q6w3V
kTZHJaNT0IYweN54A3wqypU0oT+Zn/vT7g2qzqH84w3lmmG3x3g7k+MGUL/v1deq
bxzsXg/E5yvqBIvgiRdpOOqH8Na+efjx0it473Kh7PDd0G9/mn2MPQrZFtuZ6h7z
hnzaDrkljp+59YbvqMenbQjSIQAKNRMjoPJTZTTFoM422d7PR4sCV43njaVDHP7y
AbttVYfPmJgUJEdqkIOOXEOOCr94ty+di2LrHE3KiI5jdMggwzWwYU2N0BRReSOf
pb0kBVt6xTUae5oOe9akcKKqxf4sZtup0mcHEVqWrs35pCDiMtuiKw1pRLo/Qm2Y
ZwofAw/rL6yN6AkWxYtX+3CHNILeMGrSgkIPG9NpWnHT94JsJqSqSIE+1yv3peK3
ajnReV5Z1EFjbYtJ7yFFbz7MvdFReb767KR+ODJmxI2YjAWtNHu9ApFbzRPHgZDP
VE1QpEnVD7bpPsSwBtwp21VyMUhXsb+kBi+TaROawIw5uBOGHU4tWuz2Oy/WuR7m
hvcLoGviyKSmISWYGNLED6ue2vpg1CdekRfr11Juf7tkiW4ZpyV8s2PQd8oti8Kr
pGiYr6N3Iim33N40oe/mVV0IPFruZbO2kCbYy0djRuY8+D9IHRg9A+mY0obUvPwg
19XY9mQhBlDO0CGLhiLi6N69oJjAdw1I3EoYEtS2sF/TJzCUjvR7TwDECumOX4zY
Lo330bUuZJuOO0AhgvcBr2wWim7BfQhwebPj/RpMLAG+cawtjzCv7JgWbVuT9Bpg
g3X52PcxgjiBj9cgdK95r/adHCRKl6orH/5NMgj+j3mQNN73WALhgEd6fvOHAiuU
LWVfeWTbac1WGIK0wJC59JmKyeNt8fajud1IdN1vPM58quMad3p30Yo57bqz4vTx
U6GQk4ytM1QAy7/tP+bfKARVPmgZD2O3rLDZaBIQoyxOKcqyhTUmhqZbYXq4mZNC
XCMIq39RL/6tTaeVm9xy6ix8aU4+7yo7ryrs+OZ2Zjk7W6XNmjcesjLnvmwk4yLr
aq3eN7R0Xq2b5kRXR9ylyLsKv+7PTjzbD+oZ3WQbTgQBOOD6t22ASaeI+syJWkHH
JX+j2W00Z7zFqxJkOKc/bK8BTi2jaeq4nbH5ytSgzS29QHC7ptAYUzHBzL3/ODLS
dwtEBFKeVnw71Dir/efITuetWGfz7TdqoiesOzY3Vk9YMKK6PaKUCHlRY3EnxYIL
F3KqOuqYbZW16EbPlRodvsEThvO5hghWAMfJpiBZI9UNeAHXkQAusMZ6CWfOHySV
ewJVRVpXPZmIMVlHcbluxfNHiTamCaDgwPFsFk7FVPzhk1PcOqsMuJPgGV3grAK8
vFrAuZry+OrZKXl1kXB6fI4hDjP2GRKJ4ZmlQ57/7tTHX2j2vOdXwsIYm/zPvhs7
5wsjocegdqaDgqcXUW8r+jH1XIXtjL6nsfX49dCJwnVRKggNcTTcreWxz5E6p7uL
AblUSqncxhWyRGGeF9j8fs1RvGl4n6HxW02lrwqSohsCHWLlk8xzT1XAK6WSc1yo
eG6SMH5rAe0cvsrka/1P25PMlxaBmy9WB/nua1mEFB5+kNIsNrFFpXLDG8QZW5Ju
y2c4Fq2xi80kShzylyXiXRrlB2K/VaVo9cGguAdc+LT6tbNafPzN88PGB2loY+sd
XTAZchPqji66hQU7Tt9T0+t8SomOkJ3bTIFRN+r0N2/Dq4kKaHpKHnzxNcTTQijq
wxEeasm7ddtNTc503D9HaO/zKyZSBuESMMmQWmEvJNHCVwCMJbJT34PXFTSKNV7C
aTjoYXSSO0sTEOSdFDtsR+9GoEQ5GZ/N3smczvtG9YsuwhIiEla1cEq6RqUhSS1W
/jOsfhoc8Gc5fo6iTvBa9xfUUbsI5YUrVI0fvAcrMJ8VVilhHlcHi0QIKD8yTvDN
VC3wgMZniEx0XgEGWxEN7b3ftWJ2ishiEncKcwkpWmbRTtIT6hfPVfZ2QeEVDpAk
luQeTkVy4j0QL1dBZwk9OTtlFQqsFp9FhPJSEf5sOtSkYUwtsxl07Yxf9PhVU1Tm
aJqYjzYxbiXxl64SpChBjiAX94FYWfh8rQrWnE4FdfpEoWyzB8Z46EB5qIfZQznI
ezWV01d8wEU8+7ZYmHmk+xkdHas/jpJX7VHUAjFOcBGjy+avP4ygswjNLy2yX5aZ
pG3qRRsIs9wzYgwpEqBz5Gk8i0s7GG4Ko1pMUi0QrVd4jeyie66m121QSxhFkuBu
x6usLi2sqS1c0MZ/JPaZvVis0DhYDYk7IBlIz8U03O262hPGvBAwBGzAibYBlhJm
wmA3Pmr/sPWO0ehyblcHCOJoI0/iRmS0a7fSpeFLlOx1zqUwXO8ewissrs6c2JU7
qPxa7X5nLblQiueT3Vc8j/CQx+7XL1OMKKAh9/PS0wTKVjrRhUX/m3guY3+txtQm
gqQBLhtHRw0KMyb08+l0lxhnD0W4s8K7B0S2pPkIiw2j5GLbfBzcswIfr7x/ft70
eXxwtcQuWrcm3u3DecVoaf1iNqiz7lU1/FIsz0o2Oi8iyiX89RddUcLxWO5ZRzy8
Elh4Jm5pZ31VN3g4PAomRuKVshk57afmuq0x+GdTIG36UiJx5uBNxv3Qw12UAZYJ
c1kliLb/TwTfASDghk7m+RTIB8jbaD9IvM0z00lNR9c9tfPJ06DFtJv77l/0nVYC
kkRdJqaMlGqytQWbll1glB2ug8vrk0zZcqx4pn4MOKexzWZ+og+qr+SA0H18XQwr
5hPbjBy64bumKokh+wwJXO86QvO865iZJzinHLZJiRn3EKGSw9sktHlOnepK0NK2
+tIivFsHFHJmwtOc1LjMy0XmMd8NOxJmuh+tC2OJMWVcHGgvyzmLLfojM3chMGvB
xBCYBBuPo5xsG0M51+4ZKrPWHZkV12mSeaYyaCUFQCmk7hgNkWOr3bMcazosWd+p
XN9WUKGU9UR1P1G6VDfto6y5Lg8NX0qeqvf8Ygn1+wrOK6YOitFuvccxOVgJBBSA
A0CGpXfZbt9ioYV6NViUOdmF0hTBCFZk1Af13nStq7tav/EsVt3zg8PnBIMDw1W0
6Hy5s8FD//EK7/tARlOiZri7YalPMFzLlgUVFIlVVY/vsejDxx7T4nMJzfgiu5DM
+l8OZRk9RGyltrGXEj94VatTyDYVJ65Ml4ZmPpDUmBv+oVRX+o6VM+q5oxQBML65
0PX4OnF+jlmWA1EmTDyuhkXWFEIzSiiD6ltVX2wCqgs2bJdHIgpJNqQo/ubmA1WU
2WL+hjaYTfAdBK530NDKB9IH5ruzl+CEaViXtE3S7yNgklpDx8G43aus8mBGnGBL
tiofGIuI8tSia18iAZzr0NCfqH6+BOoCafp2o9P+Jbeuz2RG+OVkazUA4zmcc385
tejm6yk6lFurEr4uyoMM/ryCaQrxIkI4db84tZOexqJzbnqIi9RJmVBDGbmP4rCt
68ZVHBY6V2TxHdL6WYcRJqy64v7f9/4zjvaPyGBW4WU2AMtFMJ1rorrfEHWPKy9M
JfyQcZ/Iu3YP0Z8n5tf4bVeF7xrVIdk8q1k1OWanBr+1qKjLOWEg7uqMWhNSiDvx
lvLrbwFV889qLRdtmwa2b83O/UV3+uIF2hm7tEN2UR4WkU3JdbM+oTfbCqgohgK0
x1Np/NxuHUvnbepxIWIdg6p+ajtbNEPR5rwrQNVn3flU7VnDW2DPWWMXOu8sir53
IC+rtzmffiBuz/evj1mga9iZBRF1RIAQLlE1ggotDj9Y34mVxSrwAu6W0R3TRKKN
SG45uYysSXSWwei7OXiIbhFEIoLiz9v4Qs2uyBBfC9qvAJV/extCdFYtOj75VxJS
t9wealPfeEzGJHNRfIhrwCKxYt1CclGgww+Q9+fniWGjqlcCTegbFFNz/ABd+vfV
b5bpigs0s8Wnzem54fI9JN6p2eFFoW6s0QI87gJXx7QbmqHoh0BzX/Lj50FoPfkC
FBd71jIc81o8luT33MYeoUOQln5z7ZFeHkz1aVxnTXCOOOjkc59CZIPfc/HF4JTH
Rzptb2Ae2JHTv3QAEISqfrxJE5cqqxT4uy7CtmpmQHX53jYgrPizrE+LjJ6qQywe
cjE0VVErW2flEtlAqz/lXSxw/NMkkJYEwIToLqcBYawYkWPr0UIFlqasmCpaqAaa
hYLclISG5H2r/V1uxzT9UtYLyqKudP7noVE5vWRcEfaZwuLU0meLLnN6nKJ6Xp7n
eH06r3P3L84LaKG7Q8E65T8dIHGHwMaenbddCGn0PQTPJ1KFXoslxGVPv51UJgf8
O0eroNzFpnwsM8P/ScNGr+oCQvUkdJl8V8Wv08bkVAzao1WVNEvpZL8aAoWTqOJB
pUb0kmdUXBGnVD4y0hdRR01nBDibnKxrq3t8lCoFk0IuhMindg47tE9+/ksy6Spr
4GdQA2Mlg76UCUQW8UglNgp6VxVFVvs/eLd+hQ4VAQOWYt+/TLAcx93lyo6Xl+5N
wLRsBKyXopznYkPsWj+m0j1itoqMcBZybdmh6QgXOlMvwvfAf6zUeJmpBz/busQ5
0puXF+CwZ497/Nn6QaSROFEzO4qdfVlXgfQWmd/NK3wm7++Vz0bN1rSI9WLXPcKm
rJZa7cA4aeABv9JIuhfVgwdSTtpgGTScGSBl400NT/Y7OLLjzIlW2zqjGPHm5eUD
VvFtZuc2S005Yhdu+Hp0puhKvMw/I9M4qxUQiHkw0qyubKxGiSPp0gQIyEahRUF0
dTpSaJx5Ky3dBD10L95CsqdFS7J2ah+aJreSYTlFvP+CC/4YEstWGrJSIutWVu1n
b6QU5ti8qA3P/SvcM6MXI539VCPne9cOx2XpDtdNF32cc6039yjw2LeU0vl+9JXn
RaCtQ2I6lFYBjp5qE6+Yf1ZVtCl3BZ1/zQxLT8IoK9UFz4Lrv6jhHDWStR35rf3r
yq7o1Q0NZtF1Pthidc5dtIZ19Kca0CVdcXnqd7RJgREtCR8c/qhUPnTEKMMrWt9C
z1/87CUmLnY9WET0jVmXTmNv9wnU/HLLjp/OgTiQtU5dmLhO/et0T1byvVefVy3A
QbTIqUL42zi2G0kqypbaBf2NmICFqJqXDIs18B8X7WAYU6EANGorbIT3xmTtgtkf
lNrjhyql/SzV20wlL8stsX/+nmRahwIzrD5kRWUHGIss9/DWvjff6XNG3i4j4Uam
lJ8pvXRdY9xXlQj5rY/WTyWa34LkHPKd/hU7Ca0FDk/iGxVEnqhwNCfwxVrihVrH
iylFpKEoaEeZpqb+GsTTrXL21rP4YbkzUViHtZj4W2oUtX1P6ZPPQEk4e6r0renP
ZKsILRAvlIfQcYvi2SFZycHeExNjXiuIwqt3XG1mSGnpzIibIWB3e/GDm4PWKpb/
lC29Bp+slOFosX0J/UqRX1eX1m+bqknPaDUGjwkiVe+DVnHcc6jeNHdTwUhnO7Su
3cln9I0fA4Blkm/1k/q3BAsVgSdhWfiFsXRDwVVOGbRqAq2WHWBBU8Timl8vmcZa
mdlI1hPbTPZSCUEolzXDf4vBvVU5uwzeGkqWqHxBXZi8EQq0HwZx7NmK/0hG6EI4
hnbjakbCNNst6a3LotdlO0AmSs2lhQZ8X/zXHARam7uy2+m3xkKcpsIhJ+QwkwTv
gI8HdM3JTpHi0/h/064DU7WnBLLeS2PFe7VpAc5S7LCbonqraPvVd8tQ+yTy7zlH
w94moNqjFNMZNriyJLG94WGOFwjS12eYgY4xUC+ZW0Fw6ss6YRwrVkPn2iaGoNrS
ruAyFMTmQBpt17nlGzTQvIynTlYRp5rrYRXqLbrO8fg9Nb29KkkQqs145poPqJgk
wWCEyjxuHSFJWMnDaK8Tzmots7VrBYxwMMNXSqt/DWWg7VhotvLjZkJQahBLiazB
eBPp/7GSqXtvY8s0V0/QrPFEsGbEplQF7P1jhpcMIAqzYzu12kHe9iJVuJt74e8q
IltsUKST5UMgg9X2eQi8oS+J4irW5bzJ860HKj7qW4/rB1Ln1YS2yj26zbJyJkTp
jWLembrR9HzZSglhwmFqzDR3g7hUBar6i8o+mnHXug4X3H6HAW7+al2Uzge1MaCg
93tbpI94+82FBqav8HiHlhwKW7T8arWLZ2Qe4AsdaDriztzwXfAYGnXk1YfRuLe9
PrCi3jub80OWl4ljcu/5b82Te3/BYYkBkbXQVJstm00vZrLOvtRQyYJEqL3gK8xX
kCiJqiQilAEUFBeiIfUY4hRuCl2nhxiHXa7jBBMkALxphLBSgHIc2rwj5Sbe0LMZ
YDf0lkHUeinKjv74dFJ6tkHIwUFEL4QmbaT1CEsX0Vum1jo8dg0q6Kpeif+Ttm1F
3wHNkZMttGj8gmaX9VkWrMKJhtxGbSNANR/wIU3jYFnjhFEdychGGn688AkVpbrG
5ksxRpm232J30W5EGx9rDBOWkj64D6T+2W8T65VDaxeYkSLghxd3A44BBdfrX+5K
JlIK5MhdHo/90ApaJRQTnUARt3pRxbZt8wL8uTjoZ9dccZOZFV6bYJ8h2FESYYyy
ppQ9R9cNSmgu17xLlOLhxbe8zVjGP7/R2Yj+d9cSMAYFXQT2i60fN62el8ULn8ZK
GFQB3wdcsywjyXO/vpoxAqQI1xOYafV1Shl8pH2PtwGG89Rh99Yz+3O2CW9g2Eiw
GSXODvt/Uxrjc+1k0molIzSShytdrVdAS+QzphrCZ7PGc6d3TllGo4EQhhEtRvFz
yxl+RywqWHcneuSLcusWzhy0omOhGDli/Dr87IOgz1Zt+DslF8U7SHSgRRDkwhsW
NXxE0+DfTvDyOo/BrnsmGGv/TgQhFMOYhcANzF9CeHdaEXllNAoP1LMDWlt1pjFv
imUgYc4aVYC+PisjH2cC2Xa9MAfvQkAeD9erRQE9K8SWX9EqQghlQrFd+TeDbN7l
QBUcRciaTmyyVlzhS/7N1AFh4qyCkqddsqILJjyFgU+yjzUmVQAMPJzxI5DtDd0c
aNEKwVxh+o+EBFhxxPwyihLKXNgk5xkAmvC/uqfeM1RMUz/EfVYyFflFJaQDD/0p
nArk5Razqbdl1WgJxE0271CZQkz29Un4Y7ZVerdZv/sldF4Q1xV1UpONP16WJkpY
lYtjCx4G/nAcGw/elWAp2zjQdyVPur96Un+AUQJt4bYy5u2TscKJjTA3fQpF4oo8
2di2Na2g4g19v5fmYynsKLxpX1LYLxmSXecBkYXtG+nz0sR7OBf3wGZe0XIlToWM
agVHLYX8Cu45ofMGV1cGwAOVWmkociJsh+BtnWJ6PDXXeYjBcGQaus+OfShYxLi0
dF09x926IdoqQ/9u2rjGqIolBdoOEJfQstxfc8/eDmgx2oMNEcP9fS2E4gFBh/98
snJHjvluYlPRnebPqgT0/0ZS2hm69F2AByct85t7y4kEhP7FqJAN3z5+o3XZoRIM
pTBEKC+YMcIwEmoV/vX3HQHt5XQzJYW4jIg1QZwFAKWFRcv4zdUgMPOoa10eC7Mg
T6Be3ZQ3V9snOiBqUndm9M83RZgUg+bO76vJpOv9kM2IdwcLz7OEh18X+pc46B8D
GcTWouL15rHVjiJmGWux2UYPrCtM/B/qEuezMs+ThkX9R33WIL/zvXhgJpgdCLaq
A0ywrIXKOJ6uo0rDtnrc7/sIGhy7p1M7VnhC6Leo6lhrEj04DPFEIMEIE72hRsnz
8yv+2N+UuBGSZeZDk1x4X5kUlWLMGP1YUeTEtp/AwP6BkyYbEjwc+CWGGDnjW7Dr
48A0u0nGOIJE2dfW47akJVLqMr/mxGwRqn8mJBdE+78=
`protect END_PROTECTED
