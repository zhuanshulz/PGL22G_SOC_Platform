`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hniwcaox9WLZfAzc3/pC7fMPYh6xw7SEhOUv/sVfcYBfqbH1uFDpQTNafgNMM//c
7UtEqDzj4+ytYBa93JvTDeaxePlRU+PnS3bl4UZ+FzRgqT3y5s6H7I/uuZUac/XI
ZnqQuJAdfyC6BqwAlvz1Dqj4ncBGEIu9RPaE3KeoMSD3smv1mvOqTaXMTDDFKSVG
VDYPBA2xXuwskNkmH6nInXWaFMt7iC6uifyfKlAw69ukgWfQ4ihajJC4/phshkUx
gthSWyy8FjP+RVg+c7qB6JpycnxwUykoid2iyl0xM+J67sPifBUHficXtstXJ+Cb
w5cbyjeNocOLFm7eQp/88XKQNfLirJV2uVtBB+5vOpoBWFWDYLmSB1RVVmWdS+kO
Sj3OFRjMJx7jspOh0Urro7cafmnyXd5pI+SBJwjE57VPDenGLs4G7B7Ckl4ztSrE
RixIGQ55ly6cFro+SmUkwVTu93sPhHQWp2AKz7j3LGnjr6b4AEn1+T1yOcYdL6ON
CufsEBveiByitQctOZTUOYNIDGnI8Y2dgNNY4KvCI9ZBO6RAxVS0S6SHgz394nse
lrgIbIBHB3C7p6+YCE7nxNLubxjF3BZ/RVWXjUkpSIL6byK/ofks8XsDGuAPxvQ1
VDcf0BtkL+DAaLYybR9FjSMLbwPiPl2xk2B6ciLXT6XgewqkJJfQ5Z6gMWt5PKQd
J8u8yz/UinvvSlhR/bzpjmZcTKp80009Xjlp7n6ha9t5zgL/9+yQ122XqE9VhwGE
9uA9yv9/8tMpsKH7bbZapvpFRqgJQeNMW3taZBqUz1JKGwOB0uwqDbqIuVqE5K62
7cadLEi4r7va2nBXLjf/iRM1H3VsrQm6xUibFopGhMuwtWAR74kMoZuf2/CIR4Jk
HWObm/aI17w4QskIIizPIR6d5kFDfDgHq3AtQNIP8fGrDp4WHmYsfWgBZKzVJ+ww
W62Zplc1WmeBv3T6mePVz4OOOR7/5QCo59NsSLd409pH9PKXo18ips+C/lJVO1Fj
iqHtntpI0YdIiM5zsymNWo0Euf6Zpskem2tgQbR9OaeXaFeGsInu+1u2RS9pjc4p
yvYebeoUzNeTxHANmnN8zAT6qdJ4Urx8mhPY6tWnwS9Wh6nQxLqCk8ELduKJbqAl
3Jrlv4j7mXniexBwCK6eg2Modo+Ko1erXRMqMxwIuhkWy3NtdwTCbuE2xmC2lFKu
94tTLVcvwB+dyESWtPwTGrWZcxxMP0Ovho64i9fp0jNRpJ/nDjwTONfMKkuFJlKH
8LFN+/ek9d7ETvaNBFyOatJ8bR7CHfaoJTnIqS4HXdNhB5/g+IdopAThFrqgUstq
dP1CpcgXJPeF+Ihws5bqOMiqSwUdzLiZG3geOlcDpYSvJU5ZO+ElewX+tSs/vcGN
AmHAInQkkSok9/z+WnL+TxQyztjuWwmQxW42sW4XebMXabbYvCLG5wEA5m0vVwUI
cGS6tj9rwhIbKeNYIHCvUcBWkcjWzddG4ZnP6rM6tMNEqliiPEnmLa8q1NAimqCH
cCtSEU2R9qQhLjyjAy1bUiC8PL/UKIzc7WHe0uIjfF9/ysu0E2CzT35FJRrHGAgQ
wGeRY1wgWThgqvmlxKzOlt6rv/nGfBITOH7S85jV4/4cNeUXZ1JKIeLZLJaBECdH
EDu35xTlUDLRJH2UqqoOv677VdjQbmclwkQqJoTSfjs5Lxrq0SdjvH2suXOi602O
YGkIbvDUvqP0LcnR3PBGvI5BRzv486ukCrM5IdbdCSuhF7wO4NFYjsW30LEN9uf3
yIYSuvbQI2/1Yg+zvRA1JYndJX+PNO+qEAx+mKkE/WqfP4xO7vpXNouYttDlFl3D
wCbwE/erwJs2ThJRZe9FPvXDZukDNPsh7QDGB1IJxYnHQds9hqQQejJvumumFw3Q
J6fZCv/V16cwgDJyQXxNJoD21I9/CrjkjEPJ5XXUg71K5uCb4h8Kw1R5cr004BdR
ragEJCPRArSRWSVHCaoa0sF85IoxbYlZ+QAT6jUwDI2UGiTDytQlXBhBJhYvC0rz
wgs1qjrqnMaaWiSoEsetfgwEnMjqh4HbW/BNJCoK7NMZKgQ9dcJxuOWWYGSkQXNP
UOyJphC+h2dqdr6/vbsrbDKR/xTdxBpLhOWnz35BsTZgAQDPH7QG4ySLYu5VMckJ
0r+iaXDHD9xzSWB6F5PbKM+oACOQHPXIh9JsrHMF25qLS/RBRAWqX/ycchYWUOZr
IKsJDG2pQ1XbL5qLLqI+03cllvfO1BSjMeqzDfuQpoCzQynKRe5Hdrssr2HXhQPY
V9HmH5P0F9zlKwJXOSd5gaj1rLfmSHNC41BCDrzjJP86NgXm3RyG/rTjkWVMJkFM
OijpiR342pbcNAn0nH0t2nflImpdxBqR12cJWvSMxSdo1rDPcNQ6TFPcEsBBb0N9
zNgerwj+7c8K24KjJUBJZ7acTXav9WvNtR1a76jd0Ip362VDcYdBicN6Jr0Ah3sr
MJrYwFioCfBPnq/VAKbJYKXkPO37dg1CU0AhnnjIOuO+uQzuetPhDBlPedBURNzn
MiG0fxa13qlN0bCf2niHlvdUHhHHQPa0bIc0/FzFz4g=
`protect END_PROTECTED
