`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pI11W4t62NlhMUU1tAfN7EmIq4RakA2f9j//zASnmOnMIA7SHTd4X41XxKzd9aWZ
7wpEKtV9YpqTmBqkLnSz08fWIe6/LxhvA0YRW9lScL1V5ohy4MOT+TWnfSf4fvkC
Jgo+TCKuzCIHYnKr5kJxe5eE/TFXvj1jMzbroo1y8mWAlyNFc9Jw4GNHwQxvgBEe
VGWNkrHrX0WNmH5IPh/1pAgiAGejSjrQn6eR0zlQe6TPv/apYxL1z5Jx+nbrP9+n
gsjHJWjwkhVDFVPjgJdgQ+ceGgZXwODhSKNZ/0/anQQ3zm1TDNOC/EAzCjKiGbRi
pV8Zasor3huPeM3/4OgVZA==
`protect END_PROTECTED
