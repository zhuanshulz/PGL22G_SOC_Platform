`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fVxurwLTpOH3pUKZYvtBz433yremjy6pTcTfD0ManolTomQebZELKpsKKM1U0zG
/VdAiDilHFJYpE9FY+QKmxWr6yub25LTaaSV2lK4b0tpd8cr1CJVdwqkYp7EkION
MiX3Nq9hSAMLom27izAEhhm2e0fu1MrQveWI6ZdBKDFg4NvtO57X7bfUwql9mxhP
AsTx98VdLNbmCRmLxSIv9Py6y9hqm6VxG9cP8BhCoTfKDizjVeBKugd8on0IXFu9
pemWv+A5vgyYTmOqlkrtqLXBRyghbDQInjtnJU3IPm/dc2nqaQhh449JeLUVzo5N
K57Pqb05N28gVk1hJHnJEpydvaFn42U7yKDJTVwAgjoxExIbzZz+ou+51gMAh8Y0
yJNeTvLFusxuAIzD4ctGkS/ltXkeCzrf3+OAr5+LxcTiGmTvJ5XT/VUUywFZniI9
gf5wWD89vT53tAGTS2miWHqAxJBjJeG0l+Jd7cQTFZG8XVFm+mp297bEH0YJOiXk
8nuXIJJQrlI+VInVE2z+2daoNd3RGmydOALsZQXeyVMPplcBRKb7zIHKerZb/eir
3Mz5w6VZPRpNZ7arWGi0yvbJHMJSh0BoZQT/AwaMePI=
`protect END_PROTECTED
