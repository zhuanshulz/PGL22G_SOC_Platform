`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuNiA3w6hiMx/o2A2Zvve6xbIxJeB1tl5fGZtNCwAXezM2WNy2QptHAIXfxDkJie
YjVImC3sz0XmWwFmCRUgtTKvwIe/v0B329QjXp++i1HAKkAP2MBhgeSOMjtZsZL4
nJsRrlYiHg1DsrI45vwDfi7VnBnil0sjFRjpzCoywU2sHVV2aiDGyOfcStw4yqW0
lUR6MuKgQL7OYQrTrmF4p0/x5cgDqauULXP+IKaTPCeDOploAOjNDIumXe1+LWtj
epBXnVwD9r7gaHEgvTAgRUime2SZBfDguwh5DQmGPhOnLnjB2dW2s44amZT3sTOs
tLtxpZbZbhniIsEqeaqPeHDsc8/rV/BuGyJjly0cEQq9QKUDUFM1N8utZsOKigud
LlM1DQk03ffgyI0e3zb8W2ZmDkPHJU8qqpUQJ/s+Mjr759ovZpcf5iCCRtNZ+QiN
8yyC9lesocywkqHNTSGIYpBmObApxmwzkO6w2FJbvMqMuq9EoxLiR+bU4GjxT0vY
iPzG8O0uZq00aO9wfpJ512Hb38lYJrfWnnBWAtZOAqB/nNVtUYXG+AyKA5XMZP1I
p4lzjNUOpexys9L+K5gNSktMxKSyytIF9E31ucffngydAHiNgpA7lX+mXeZseQwA
2sDhtDJk/yYS5L/Bt/VDBihIP0FN5r58aBbw0rIrbgh+Wl0M2qUH2l9FbEFwAFjC
8DVQYfb9qekqWegtxOFkhEou/Yc1dlJ4oKLfMksH/akztq3NcpHOAEB2osfFDYU7
KQ70P/9E2xaA/JIob4xlS/5NGQ4ss3XOjqdvaAeiGbCeCt5tCNM6MbP+IgU95aEU
uPVI95bxSOe6XSwh7qFlMok/AMNdjVvK2aWCvEcCm4pANG9NgIhRvyZeKD3mJ3aB
QTl0FXcr3FAgZgfBnfd0JXWa+RErZsmPHISQO2nJefvWuRs+WfE1e/xCMWIFF3kI
vjt3nC5dFpol9tn5ZlLcBa/gS1m9h47dRItNjsC2yBkmynR46V1Woy+LF1YJMnaR
dlmIHjX7bjT5P9g8qeinP1PlITmT5Kn04YnxiGcD7wIhowMDWBsZLhPv/7rasWol
c+AOPFqn9uh16rjZYEHqGwIrPzOnOXXMAp+g3a1hGTxhGnWiz7/1j2sFNAWymXSw
HApluxaM8CuOfRbSK+mrKwtRFguGkFulCxO9cD+oKO+VGTIAKCtxE4bFp8NREMso
qu+u2YT88G3x+wM+MHpH0kzoectmE51c9oDVDYXxYHr2wfCYZA/YnYAHcEcRqLvL
8qEguxvd9DQPrhEg83nF/Rz5boRhChiV9bXVK9VO8lWW5YtYl+5c9BXvsKGPgo6U
BblwmmF3flPxgiyuxfy5kO+g0UM24UtFpWmsfvDuKcnpynJNrB8iiBdlpDTxE4A7
ypbDIdSsBA2Ukq90Xt0GuCGId2bARq/Y+M815H21cSv9Y6bYcF0yIY+dUgd2QSzh
xBRd/0ultN72waTWyOumueQiRj67MLbe6WDVIa3KUxOotAPUMzjTrnnH++r/NlKD
fk0J8hTuL30cN7+Mns1+GP68ITNrYsy7GjKUAVjk5iNCK8wPw/OjDYPwWiLmJNqh
qeN2PcvtaREkZgPYaMC3ElcvaB15trPNn5kJ1OHZr9kivl6tFW8/izsxAmr2WnbK
m1OONl5z/J+iC0Cgw1uAIxF3s40RKjROrwzMSA9sWGc+6Nu/u6t7aPK2bGS75A9W
zChw/k5tiW9TUW2mTazzF/jyn0OoyiviSmpBkzZyAXfnweTssIL2/0VgpEG9s3o9
jX8jfkK3tKt0gN5HZPbU5GFscYopH26cJ/A61scQWYbR/fPbkY5zN5hNZfiFCTkm
S5yNwNYklMh2a1E7mrlPJ0CUq7blN1jcoQYa1Xo2wcI7Revb99nYaGX6JtNArHaL
CKthWTWaUBfO+nX6kQh0T0MCR11HyrauCBjg9/cjYmo/ImKYSSEHlBmDn+k1WbzN
TlC7hQGs0MdlacPBY/cABb5/A6d7Vd7N3O4+WoJ1ohORfozAAPkS9r3AccTh3afI
bs+t5lfXgUtILg9zlk64BUj3dh7Axej7/jwIAkbAAoIfabgPFsBy4hUdec2NG+TR
82pY09JpzQXRg45KIIoZ3aX1zJI390Y6LaHJTsuixkbFoE4uUKmXR2ZSsyZuxlbG
72tWpTTAa8oDOoCaMt7I2XX35DhJTkpXjNGNP+Qt9g8spR9JXLerGulIrXif7ICy
cwnzWg4fgqpN2fQ49FgjYzEwiLmUxoQNIrn3Deherefs8a628dDhpPx5sU3YJQvI
TpeX+wDov7dD2vcN1ROBe5UGgIc+fG2PpJJqHgbPyQeQfD9jNqTq8m9+bV0U023f
Fl8J2HnjbMLm8nTu0UFlCSeYB+B/GkTaeDK4N9Yz073agGUHAx5VO12CdbjpeAiM
DWnLGfnPZltpAcePAIVrLPH6hgQJ1LIaqBKFvDwbufDrh6+S+s4wGMt10iroATrW
AMKaMc17AKBIZY/WbuLZWLp4EW4z2MLQo+S/r6hJP+1F8R62nTaQec+mHbg2rQY4
ReHzpCOQdj4IJtcwUK+fexAJZ6Fbr/Vzo5FlJGg4KHpyejFbu25/6t4Lvxk4skY4
zmQl/WHNMsoBPAiJiLN9EQ67YZZBP0ni89rsc0UliOxRFn0zYRO2mbxOaCNbSyxE
YYG/Zb9OXykw7ZhzkfyMJpGYb7HAA6QGO8Wv7f06bE0DwPEOmKAsV9ftyyZYk8vF
7qruGAo0L+ghsyXu+FZ7vzinO511jm2ucwiuBpCjAruwTIrPt6HzegdErYlkul8J
imPpwcPwZHla0lr5qOaFRvdPNXUfijZb1V8FnaYf5tg1bbOEuI7vvnBI9uCXAzO/
OSybvHccwemI45ZPWRxXfBHOZpel48YqMrOyV5KwJw71a8s/OJ7Vfu61/eMlo81c
UMSEnZ1dXhTnIlXnwEtnWTBd054dylg7PQkgLg1vPwUOa8il+kMvejitBv+du3WH
pQ+LfPZDiwfRXM/IwVb9WbiyNo/nZekMSA2zZlUm4+UQV4cYo9W6M9Ae6RHLlgWc
gdk0iyxHi0P4kCqZ/lt61REAlFBwcS9js62/dgWIb8aRqUXlCjr3Suimp1ly2b8k
daIfXZvS69oJlJAYY+vS8nuhtcQiTJOyibqx+wO0aAx3CBEmmUpaH2k3bIyI3kE3
3bLJyyZwB5F9Bv2ph5V5W2qvR1dKGiZUclpXPhzUhtHhASen1mNhbi5FR1rHU7Re
55pyoAWfvVMB/R2fxd9J/feWRl+Wy90SuPgZvJ2S2Bi19GnrHvvYyQQlAUAtAaqR
EiuKtyrqlWjnveyj4i98VrmnxFwKnmRXvJ/pip3v5WoL1OAPQ2rInkqEFgYFcnGq
jEKCnBvlarkhZr1YYiyfqW2NWv0k+24r6AfX+rVOqIJ+09cvIJHFQjLEcn6qoCWk
p5tnYu6hkhZOvEWScwAd9SGYHww5th3HV7h0Qvyq38DLyhhQ3woUq9mcG/CFSCQj
MZcv4v4dHRu5qi1pYk0NmN0tcYvZQTyfkb/M5hnvsBqPQMEIMtKLNaUjGwlcgWx1
tBDsuVRQILlll+pLu8aYJcMzdkY8UL0XBZRzTFD85FnNHICsta4eX5hFj+oU+t4e
t7meim6CHUQ2TIcNCKnK8H3JYV8C/py3y54zynaRGq6XS4pgzvCd2+PbwbB4WbdU
`protect END_PROTECTED
