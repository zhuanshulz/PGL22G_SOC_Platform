`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ofCJzzlFW5+oozhAMmMFW1Atd6ktr1N8RHTWlR1pKD6rta+7hv2AfJUXNcc1PSVV
x6w1+gn+5ld9Ni/KrVGkZlobhSRjRwtdoIb2wrWXSUAzm3xakc94UTJimmiuY2Di
wyakM9zzKwh/w3RlD+7q0R5i3I90MpWVY3C2/AtmUeSHcDgYx7uIpAc1+MbRT48X
9kFQ5HrwykB+8tCc26DGs90gcFoNr1N3aZLeI+kFUNyMui5NEOugCH62BhIAD2/9
1NUn9FRFkDLtS4V2IC72zBrYvlTstUo+SK4WShzpLxgXewlvCNG1CmAhgFE3avvb
OR1Xj4+FcvXLtyVE7Tw46Jqel8dsJ0we/82LjOP9eCE895zxxsgTJZQeMtm9/ewU
seQL2wb3wR4s2G3jjCPeoB5doUo8BHAsCZHWH2EsduU9jVfbWjzhPKrDxlbL1yhO
T0cst73cAnJtyef2pznKxvUKFiwPrN3xumpTmLI0vDFtONlgHgDKSdR6gjREU6Cz
kCc/69M3naEIHu9L9ofy8fgG8J/Hnd1OOSPVQ6qx2aGRvb4SdhlKENVv1PCMZYob
e7bGb3/cOLf8UNUcV5f4geqPn4iHrxzGmQaDt8gK3oWaSW8beUhAzO69T5JVzIH5
UZDF1pPSWODMSb4NdJGX+SU1sX+Le6pVn5++dIBOP+VKV3ABuaKPuRRfKXf2pup5
ZTeTglhK373HTe2AVmBSf1meafdqJ8rmyGCiuXswzDDdqtDfLv1yzCVHBG+mPryg
gcYtCHGw2x78f/N9sD3+j3zx0Si69rEDjwqik1D2Q+iftZTOIiUbvU3MlvNKmnYs
aK1mdjKOBQMNJNJOD6VPEg==
`protect END_PROTECTED
