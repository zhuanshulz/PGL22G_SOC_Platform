`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
inl29qbU7YvGd1M03QX1IiXk7CaoPj/q3oBiDAcjf2kvGETDZ/GY1VloxDbGIqJa
d070XNAhGsg9timexT+RbbWzJDSC6Iyp3OPksFq9hhSS2rzV4DyW9n+TQiqNSJos
OJUl0PR1IVXxKEj+Wnk9bAlOwNiRTFeU79AG6DtiZUtVzBCsLmhkN1zb5d1ZdQrK
hdSnpawACvHn6AW5LCp2ARz0VebEVl8j9hS0xTFz1O6Tc0wIrG/xxOaZ1rYCOoS0
wMrsshl4R/W/2uLSdu77p2dfbcw4/l2jiXP0psWgiCDO7FzORCegP+xRzpPH67nW
Um47QrbcN8aGWns0Oq/1hkl15iIMGzp8Ek+Z+XGzXXt388j++PZn+IUGDQwcqybS
Si/06I8eAQV8h/cYb2Zyubsq8P5kdRW5yBLKEac3d2xyiivTN2rmvanjgHONzP03
vXOgLLMCLiqtsoGqfVJHUdvNtAnIJyQlrcwcCMtEhGmfqpOlsV5Z0PDXgXI/0DfI
DJWJ7UZUMVPfWe7UTO8Gc1s5TL9gZFlkcmLMZe8SaGQ1AezHhDPpSgJQeQBn2IMG
awL1W7sXH0n9eDTxpzKisu00Qf0Id7UHF3LO7LqPcXNbdano18FYIkzUrTKFd+dM
PkXDwl4mX2iIUGKj9vGoYh6LC7LIb0UzGJ8ut82vku11lU+ZXTBkFJH0F/jLBrk4
cFl3kTQHk23dA13bmKO2BnnGm+p6VWnb9fRZtdZAHJ5M2buKT26L8f75GfxH1M2+
SGciigGVR03S3hfi4EUH55N+NuYVKoab/RlB97usKAm8reZLVK7T+UysMtecJuB4
XFzi8kbHYIR0xhcaSiYJA+3aqZnbkxeFCt1p6sIvoF9k2UeXGgPpYhMyaXzLR+bw
V6RDXqw81FK92VWpl64dct/VOWPC9wovbEH0G5985W6fcsDEyOWPLzv5jriiHGZZ
Dr45oUDkAIrIEAVka+kUIc8EIbudI6uOQv9GPVz45Kj/U3ZN2vgWe4TZOmT2jAdj
vaYJiwgm9kN6eCYjw41O2NHe3W/b5PvQtZy++ZgEfvp7ZOK1pVkZoNh2FEtPjQcX
Z9/MUXPFPX7qVDsCW1WW6FatnVRgADhQ3nTvKATilmGvZXNoktKvzpxdXUga6Z0r
bdWNMZKJx2dghgyLM1xURQ==
`protect END_PROTECTED
