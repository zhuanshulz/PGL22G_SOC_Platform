`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l44wPt4VgidFT8/BC9Ckz0PhCgJhB+VPD6xxAiPuNn2C4jhz+UlaKjBniCsUc40b
7TvFrjfLsSEX84MyaPvksm+Aa0FXW7v1bBAi2z8nrbReJTSFGQQb0NOu6suGuxM3
Z36B8nfaymUoz4Vn+wBiPZrqfVFH4MrX/uDj4BHQCe6AOAfEFE/16FietiZix5pn
JbuFa6PoY3TRB3KR/6LG6ZLU6acwBma1CdRLjHqDH+l/rSCKQAkyFzkKSjs8fSnm
Nj09clTHnFmieymABJncydIKwZQHy0/KxHAejYnMKtKskq1a009fa1qRhaZ14jlf
Sf+VnkkXByBXbZ4jbJjc2H+yd3y5Yvkewc023pgEEnfVjF4gAEnSXwHE3SAD1I6c
xxl5DF3qNDcCeAoMdKWKNXBDH6Ei1sYCWmA7GgMgCk5Zhah+1TnX6nqHdu+e264q
yTbpv74VykoctotmscYME62WsCbyiZ+NmzkA+EvTh6Y4hxEk4OzCjiAk4UdpoDfA
tngjde7GR8PDOSIywEoI3pyuWublhHeq9Ry6O2jBSXaCEAWKt7F1egb2sP004S5P
FhfgFVJ9wjj3gBU/YT1zknjBOmGs7U4cZ5ViOB/5eScfLvoyTnLXea+mRws0ZehU
a5pLvmr9p2v4O5ZxdQy5B7te1Kl3v0iMEGg7NjDsrodBPC3Zqs+T4yE5PrqvwkaI
X0m6ndM61+MY1/jMGTCLShJFW7Nb/h5BcCzqrVgvmWVMNnYhme8nuDuC/j9gJzLB
5BiDJKaCCj+o/UV+g93TaA==
`protect END_PROTECTED
