`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RN1Zfm3vNv1gAm8p85xoviXtjGcvRsjrDzqz4srdfAO8E04YbEFOI04doexHEAdh
4+jQGoWfkVxLiDQgSd2MoXUIeMds44QZuiyUHxW8qYuzpipsuAdyWyx2dn1F0bNO
xiIR5vuKry/qad5nrim5gly3ESeOghv4n1TPH1FVwGcZZObcklOvyYIHGYDqxpVX
NQEic0VAArO8PTe4b8WsTonXfOWOhHrU/5U1CHIBIwN4vONm7OpcVAarvdW6oabB
VJsKeXnVd9rFrJyLuCS6XrZQKitdx6zQ3uCG32jUX9n3445aTYFAW+pq3SG5k6cs
vYKgTSex39V6M5YOOW3XXg==
`protect END_PROTECTED
