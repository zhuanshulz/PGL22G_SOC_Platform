`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
api6G3p8Vleny/T5eOCKdpKDOgLhRzPTm1myLjV2ZedHzd1PKvN9dl9RjcNsPmaL
Kbyr7xbylmtC6lU1bhYymfn+oX9qxlUCV32tqQ5rOWwa1N83GpYxd5mcP4BZTumk
LCkacTSK1iCs1C2YW0Hk2PEB64AK9VdODslTq9y59+nxRGZjpmNzz7zdbUZPLDCc
n8OOlc2SPKVBwlf3eV8s7Ki7dDwZnwVZjgAkwqXWS1eSVil4S8ENriew/x/+Awaw
BXMD9zPeErVh0/upiztJXF3UUL3r/GHcwN/9z1kJLrq4WJwyu2eZ9/8/62oimQSv
G53ee3Vdsj0DOEMrshPHUFmQMAQiscvC8Yf7l8pSOno48cmAj0hvXLj70eZla+RU
XkQBkAf29G2lUG/Z9Z4o1hDuSLGrGdjIdkrVztjbdsY/+Bjoc8+k/PSw8U+Xe0yB
3BaJyVSd1jT33sOlvip3X1e+NAuFC3RSI0HS7UsChdLcAblRC0xnfbM69BmaL4/R
4bAtxDLHFP9E+dQEvl6eWXXu7AWRoN1CjYj0vU6ZUoNS/mb2oU3D3pbY+woqGzlT
0N3H0Fnl7eKXEH/hqSICEo1V7a0THSKIFsEXj6vYK1YvGBf1urSFbf63Si2DPjG3
o5OO2dB8ugfyLLp6jlo9v+LmRsBwGM9rGS8NtJVRA0M=
`protect END_PROTECTED
