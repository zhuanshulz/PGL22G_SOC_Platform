`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rh0LbKr8P309r150/tYXYwJKJjeaGH2wWiGJjT40lKPXhmmVNur+/Sx+WLrG1qDs
mTHsZrSg+/6mYNEY9HOKw0sJ+NJqMQPM3FkB6DoB/6iKNvbqser0DnPoWj4kWcg+
JXdmfgPfg+eHvhewJhqBZQOBcMJr5cVmzPQ9tTeYCqYxNnc1N7EeGn201l3NE1qB
YyRICZTe5gFH6sz17iE4t7CWjya/FJuVIv1vvVxWBoDS5F6b9+8xvuZ9hqAPE4bb
2UlR85FBksIC+cQsDjyXqAbc7TA/CQtMKIyjVWo8fs8=
`protect END_PROTECTED
