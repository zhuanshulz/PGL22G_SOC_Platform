`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+dLs5EtWgBskJDNunOLN0+VWP7sI/EemKjhHVuxkpPWIT1LYpfMgzIh0LMiVhCb
bqolEHi2HO++U9myiJntH9xeypT1tON2DGrsSxeJk26YL6KeimROPNXPCUC8o4gD
i4q5A9N3/Qp9F3Kr1fdoEXnYYvalfaBCC32CP2KH/GrAxKBt/Vu81LkJeHKZA/qv
pMtSx3fN/gnMVSvdcocIfIZze7l2alXJf/ts67k6VgRrrIaWIxTcXi87ccCv1QKh
bQ8Xc24kP9355Al/qCA/YLPElsq2OTX1rJNJfBDCqEhiVJmvboEP110YAdVERRyZ
q+wruElTeXggRi3m81jD+tYXFilMHs5gh/FyVPtTLNb9AjMKMMH/hl5hnAZJm+uq
bZhCID0ZDk8B7BOPxZkHlhurWf1UcqnzyjvL+ckKt+NcPaI23qaTtju5PSJlGVpb
6WTXADr+eMB9YBs0lf+nQY0bQZ8m7/3tJmI9Kxmd/A3LDvYeJB1tNBucqlvzFBUo
lWhCosoZjlyzYqqbaoY6fg==
`protect END_PROTECTED
