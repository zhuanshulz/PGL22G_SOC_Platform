`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ch4liC2RMYYvbGMrGoebJnPFazwlWuYl5BW12Gc98+BAxs0bbRRjnpy6gLwOJX4
lWic1YPtnEBtdFABnqvO0AJK5Ae59NMZGqqFDRGC6jPvMloeJWIVkFNk97c7ERWr
H4YgDaz6fgjPeGGO1o8ePuGnnpbwcFDubnzsF/qJgrrqhHjNGoHypW8w+KAuKs8/
vIuUaPq/W/ZjU+dMrGGvcXrB5VXI9sVc7UeyQ7jyOytM5AwvcsLkc10oSOy8Y72c
z5rvlg9Rzpb2fXWMh10mlzYejeeK6fpGiKgeSY+VnviCJDhlK0Zcme4AYLOnwW6X
k6mPXDIM9DJ8Syihljw42hJFSR6w1qZM9EdW4dNo/qwDTIGLw6IcY9Gkb+nNlQa7
d/FHK9sH95e9NuqxnQeWyWhRDuGylE92mGg1P/Ss01mI/qU0uOLhewjy8IHbfM70
0QDqh3xe8sV9pU/WVmDYM8p8ykS3lLGMJ35YV7VmJph2aF3I8hUnf/ETLAhtMXxj
msI5BGNx1pAidIVFDmd6yxrUUaT+nDwHwzivw4esx1fmb4t6RRBHZLjGqt85yc55
hg7cyJbv6H9e4cLhs0prrCsXHP/IDjxfYXkfGArf00Led4FT7kmIXfuAaTR90keK
/k6blyr3vcwOTHUhWhIBczFtbKHZyJWNuU5HTJRi9hIMVD7VvqKVIwCVat/jAksw
yQnb8/w7modHUi6m/fVBKnQIymqN19qm+C9U4NGBgIP9aYZTxlIyyLPxP33Rwduz
nCnubhOj6VRzqhBKmpap8w4KLDr5p1ZdT98cnvtmmxB8CLDA46zgqI9Nl4+iZQJy
IAwFCMvgGwzZP+DstKC3NSqpMeL9RUW0AOpUZDoL16Sq46fyLsEvs2A5Urj9Yp6Y
++tm4NPtW1/OENXBUv2dA0LchKriXL5C04feSgRolihnho1LqVcRCwN9BQCURbFr
Ek2wOgbI9K2GoDqK5x0Xkd/uZc+rzdW7RaLE8QroWnMiVA6bABnfleWYw4p057ys
Lh9LOpqnVVOE5PAxnrL/14sCyRwTw6nmLnB/zsoFhKs3akyGSPdJAko9Q2czfVjb
`protect END_PROTECTED
