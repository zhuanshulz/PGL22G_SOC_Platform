`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glUyb9IVFo6wWayj0Tr1/8kz16k0RPI3J9mSXfsQf+QUcAfe1UHbnEk8YFUO+nkR
hHx38FXQPL/QpxGFSWUOLMIuRh6FQINhrgppANfqH0URdjpAPSrJWUb4o13aPA5T
C+DqhoWV4naU6tQmbPrXfkjxeMz7pKLVlaiEQgHvqvSw/7mVdbeeNotWA7VuRKl4
1KC0rqCj64OTXN92dfNlTrDFYfnx5LMIdYM76W7Rwg7vZZjybYj/5lpo+0ZQ5aOm
mgGwGsrWkEyyJg2Dw4oCC1S39X3qlvuoXFvQQyNvoMs5BxokTEz57lBCKgTcSjlA
YJ7lUrVSobyC2b9aOYZ+xFX73eq0rHW3gQXSHEPW/DFuvBbK+DmRXmMaOD9BcYOz
Y3cwlnc4rrXZ+iRUB+XNh2FaekI/1CiPiAMEfRM/HzTtaCN7o8xx2OYpkSfzwTf2
y8wNzQRSohEbCLIcgQ/9vdxqf7k8PSk/aV+jjBl3BzgRaVZapUch2u95vd8K9fkD
u4tSfILLlNOoQRnOgBPN0AjirFvhIJ+u613q0L9K6ujG5qdAnHCexcXYgD/T7+f9
xPAWqmKdJ1wxnbhGbGSWL+JxCyJEYI9PTNmiJKa51hH7bk/0xffXLnmzS1d6iML6
rG7ofPEtxy6J97I8xWTFVQ+0PGM19D12uT5TaFvsLq1L35MbTMpT0SqSzAACYARR
WOq1dz37XZBJvhLwbeyMhcnbuFvmuWiLtbJ8K8IUjKTt6EJcX5QkGbMp4BBCr6+e
Ynlpd2M8ymF/JACX4fayl2Ley2w7s7op5Se2/X4Zac8WGZzwfa9KU1FU4LMgNCHg
k511SbOYWlM5ZyEiTAHQ08VqqbmZ3ZX9pN08JLiJdXATrIHGlq4RC9rRr0GjFMPK
KfygWI1cUChGl9hvgpJMMm8Rs0a6uPTPzMFB2/u0sr40miyINZwDlexYZTfx7FDJ
9CKr5o8MRy2Wlwrwgc8jr7av9NluQB3NFJNwEfE7NGQfDbDl2lA93FelIyW0YSsC
mr534LJ0NeZPSlVCeFQWohRSe8qnK8yssXlMiRj/rTDTzi8cfPMZEXeEzDP6dYUj
+si5QC/+uWHyhkySbJzXclK1eRt+BvE1fE6tVNhTjmsvhGiNP+oAmrqLUp2AuZ4p
2lyB+oDxqjD3ZCEto/Xc2G2LUIqM6rf36V2+1OB788Np1M+yZxaV1ew731jaPNsq
e+oBw89qB8Unce/Bf5t+L9YG+o9fda7unMuADN+oFMuWWF7lOS98SzxH55eJC3iu
W4qNnjctZTybpbgey3CMENyR8DgFMlTDh3Uphx0XEK0+6WFBlE+7y5CIVR9CNdw2
kqiPMESHlL+5Ff5fMnvofepOtePXmHc0pynbvIPJFLHYcTXmT3KKXuIx4o33dl9j
SrHrzspSJzJv3xFZydJGE7Ytud9YR6ujM95SihUbwHk8mFgYKdhcqrpoDY1XzH99
N0V93IbJgNZBCTWfGI8MV4aHkn40m9QbrX2hoUe24rMX2bTWgrkJOOOetmxMHTLF
DjvpHYCrKnUafYQI12MOnIcXILAv6gmPEnt1Xb4ncfZefRkZWJiEgIpLayDcyE8t
jQHTvB+NRaSN2mPs6bZDqw6TcE1VSnvQ0gRRhIfZ7fGktQKFn7kzJecCxrK9B3PI
Srwu6+LWBPDhH1+udpRouzQ88qCTnz+kgccIOkv0gmW1bMfTkT4oN/Z5oj6XFU15
l5Z1Kt1s69BEuhyGPiikA8cAMcdpMpiHKtGvI0HRabfjEhDp+20EJZD4314JkeYH
bT4FeGDd0hx2OPdTPH4S8Kr2B78zU0A8Ejsqn00wRupEIEfvpULM9jbx8wo9UYjx
I4l9spXU5NPeopNxmDyVARv1VE4UxmF3H7+j7wufeFrjwJFoMVkLLyPislcImsiC
pBJtofvuAgnQ9NbW3GSJDzIP8cO5lasRV+v3xnmmZceBCbdjda1H6ePm1Xph3Gpo
Jb38oSwBihhwtcRi/9vFVio3bwg27jXSJ14gvXzLxm08bqqkY/zByaRvQkUZTSLp
PPDIwVN5kWcHkoNbE51rHQ7uB3NSfOcBMJAkFQ+FMmmd0JcCwt1dHaBCIjhAISTR
Id+VXOGaYEJLq3d5nJ5PZbMQtCEoeUKB+NYfPj21mAd71wswkCsIz2ZP0uhKcWiV
+o0HM0mCFf68DRnzfSys6se6ijgvkQr7JuKJy0szBbERGtDOwovJjGMseY6bAm1Z
l1kysay62AFaaIe8VGTfefrKIpa50CEEOgMtFSuz0nLXayKK2phfMbYuutQQ8xtT
WiKa9uvTYC7TML5EXZ6UvnZZ4krlUJMykYr/+FfnFrJW7FXMUr0RM48o6De/SEw1
RgVnrCYF64ixV4S9QVtVXA6Wt+vGXn5AGnZO+i4+A8OWg2IrBsIcZZzRUb5xLGj1
JGMAxCsPXJw8mqrjmEYq7AFzpmq/TkK95JhTt6/OEoYwqWnEYnrg+K/cLtAYECJ7
WPUrcBExz4xkuux97UpdrDIN+APsvjG/iXzOgCZy51WP3+P7lfruJSyAKQCiLB46
iI1tQJZNFIu/62Cs7eqavgTnHBWaePGDEHK4g2nq8TW/iGwDWRwP8LQ7F+VK7QFQ
xJUCt2CoxnwwuQYAowf2qt7nCM92lCoOo9OUtJ1ySed7tFXobESZQ3eyWJVAsUg8
cMA/T0DyeT64JwTTR6dkuicB0zg9BzgEEaGuBFohWux4ogDdkRL7CmPTCMAuYhFa
EPZfxfc8Ng2HZBpqI42eqapruT+wjYhSKjQR897DuR1R+MjPYCWm1BmqgvyF31Yp
cAlBezEhB5nXvtWm8uq1pP5k195mF3rBgvCcYqzzZl/WhkA6KkMqvcUN7FX4XI/n
ZKoIRh0liFqbq6diegtNQTV1FT2srRC1Ow8hhvbnHm4hzKjqYtzjuIWvH5nvJMAY
s5emCvtkGP1YeGsXlv9FMlnf778wzVssO43C0hvBD33F5i/lzooOGJd7ULyTULxZ
1PDDzlGMILoVijiWyACIRFHfn+KdIfMbA/PMr+/67D0w6a6jgJiTqbjpmXEjPm7O
4g78ABBI67cAwAX4OMsazJh8Vx+pYL/Rqc72JZcGOr1i+YqDfmTdOKlmbIKPjwmz
q4ZSQT6pPknRvKqOzU09+s6HWfSGUomW9lWQyUgZmVVJ73UfSQuRDdj34Egtp+7I
79BjfUg9VyrkKhV4cmG7NsrLx7b3773XVP/xxwPtLvPEDWwvf8Pj/P4bhBRvAmPw
sY4+DBm8KLS1KM9CsLYZGDkApG2fXulKnmi7pHA9akLYnYzFjl8QrHN6A7Hro4NU
0eawD9i2J3Y2YUioBdfpz09+e0VlstaQN/yBJVGgVIGSj265x+aYttXuBQkZOgHm
Jp18vpINZTeoGIYqFzQdFTmevUHTgAdGOQObl/2MlK64ZhoX4s4iyEg2muHxyESh
2LDJqFSwKq/c2NBW38q/9bihOotaTUYNMLjwRH+UKRU6kDdov3hIboL8YMBSdG02
onnmA9wxtSFpBysvADMR/Obrbb/FGEpSzB/3fM55IhqtC8788dFBPKJ3G2vfheIV
5EeXOPiRxyYC5kMFq6sk0MInU3PTJnGPupcJtkq/icYwnglcIavdb0vme2er9y+f
BdQkHRM7y6cn0oUUZfzLO29loLTYJW12viOGM+B031N0K0uu5Yyo6AzmGBjghrSO
UuJu0XVIqw8RJ6KuqxP/hDdS0wGVIvYgQNM2gJwLR007aV56pA2vh7/zNdo4/IGq
ptZJqWpiQtVwLQ89YKrBFlljRhVVaxnZZ5j9XJjiBvKpNKAq2kS1cTx+pGJ6rYcr
NJMikCEoMZuRjrSNyXFMTohhNPIlSMqvDVtHjXfiamu82JtTwzuvq1cyb+NlF6Is
eTBHx9AKJPLaj2q9v5jmPv53cXY8o6da7k23vENmeqN32Uq/lnxPHSL0sv5fCkQj
fRUJ1aOl5ssHNzQIVfTetzOiNMBrVzeL9LDLHjIfzvZCVI8wpYQ3NawLpMy1YKU9
5PtBsnwuOhD18DLt+kKAKi7lj/4W9TCId0I+YwgpbJUgYyL9+v3QrhWEwziojeyC
FK5GABSQ154492zihqW8NvHIE5qiBub5Bxcv6tUML1s8DdD+YAlXZaLO0K2hKqxk
+S7Dv1mVeCe8YhU7oXrZPOcLVsJCdOgQ1Ke2D8S/6OIF2HZaPJwNNXcKKQMTKeaj
`protect END_PROTECTED
