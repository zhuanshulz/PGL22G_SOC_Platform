`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VxFBFGeswrqWZG3ZO4uJ1N7Pcrzw3ypELbp1O5aVXWyt2pkd6DuRj+NOGBLLqyZ0
QTO8ljxjzE0J0E7ZxfcTmIm0o0mwcwbP8nKXkkUwG6G49eZ/CeVShC2g9wep306b
ikP22+eTfTVy1O1mhJCl6wayAs0NzyOQ9HRg6F3wkKRjJ5sR0wLFNu0VNSVGPJtz
ciO5sg2EEc+Oe70xrKc9jW68IV7byqT8MmSyR/yNLYNdLjWrK38Jx6JCam7y7na5
`protect END_PROTECTED
