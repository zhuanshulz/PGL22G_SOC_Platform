`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
acdDvlVoX11o9V9BxYXYxM2EzPQEiHTfZ1x6LrOAChwUD8U60HjW53ZK7+omXE2f
n+xLCRnSEYfiWeMDHp25fcITW3Mi0UlZ4M9Ceh2fyLeMNIIkGoB2r03Xbjc7WRpV
XTcglHMga53sOnnKDxREz5tVIQLneVl52ZT58MgJBZbbPsdwk8aZ/XXllGirxIB1
UFqarwdRbh8tt/DHpcdCbQmYbUnQazF+8Np12Eq9EUa9qAbDS513djOGiAmbNW8k
beGZDQUMf5yYTe/trcdqpTKIACdiwbXenoVsMF2GyhM84ZoW8Ir5t72eoN0zCrMI
Mf0Lx7jr/UtgHLIeCKhjy3p1jxx7s+FMdT7uPrbX+ni3spzNwjvlKB+f5ifqawFC
Md6V9W+IpSM5cn8aERb4EBo+536AfC7p2rUxjEN4mkD65HRO0qZ7yU+0RAv0fMNI
Qz4YIr+aVG7tbsLTSfUk/g==
`protect END_PROTECTED
