`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MoasfcZ7lV9hnK8R/KdN3vsJ00i5s4TGr0f6+sEPS5lBEwl+XvpYYhxDppohYEb7
pG1uK4dPbY4IyCj8U5e1582rFRj5RoosFIPlZO5C42tCfSXnrmP2AvtZIjKtI95X
Ahych45FJ2Q6gR1nCMnq8V60OwBw7xeyGIh5iDjS+OUggkNnrms2oGvIREzRR6pu
YIRCCH4tFVs5egYWR5ZaQ0qiV9Jn/GPX+9tOmMYRy1M1UIyouZsznetFA4iUg2/v
KsUUAh2SmZUkC0iaZCYnILVfxskyhCZFolrxSyiCYzapUQlKkb3s/Wrs85IAIdPs
umGqMCFoEg2vbolW9jqhNA0qIBtYzIFjUysjyKe4gm0TEnmpc/RN9Eg7uFDTyjd9
kqNfGpss0Q9M0nP26LMgHwEgYM/eHp29YUZqfb+cHVziCzTl4DFyNJfgTjTiBFpd
8RGAan6LZBnD54qH03AgZ6c+SuNk2D+4hUhOqUaeyz3RvwFeCTB5YzRxnxkXBQMq
+omocOYYDRXY9Mxfn++pIpaM6msWf3eiR6Z9LX9Dycg1NmDr0lDcFHfeBfqmGSHj
YsElDoP1p69yD2wnU1YV9F8QA+9QvnJRqwYT6u+UbfXtWInC5bagYbeBCkM7FLiZ
UNoX4nsgv2sOWI3qc7FE3fWt0xVR5RrVS6OMXajPNjei22EBC1qMEWLwuk9HANkc
nksRRzKLxVOK//iWnVJAkKCgb1nsQPt08g0pKnHNNr+ySz+LCOTkN9nJiZHeIP4o
CbNkAkvIq0NgSmVu3yOg4tftC4Vksb8qqppedyB1QsAlcs7EVSGKQvCjqw6410bv
Oy3XYh8KGEl2q0+3KdiZ7wXO/+EQ9WuUkPe2XFITPLdGem/HfucY82VZnbJ4UvWV
OC5lA0jDfpC32a3f1IAOVplZ79+dCF8kL1N6swrY21cBArVbl405mJ27XGtN7b7r
FnqvT2YNuI+PI86WTlMXxQ==
`protect END_PROTECTED
