`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FnmGaOMKNvDR6tyPycU9z/8rzwCvCVOSQVbb4XvlJtQXc0c/B7nfCSrNJX7GbG53
V5Y+L91xP8MfR/tU/MHtAMV9NdMU6w3iZA0VXS69Sg7S91PEWgY8jTZC1TnhOYr/
G9SD0LQeW/gwQUFbKvGKQZFInur9zDbavsxDKPhI76zXOdfL4Ucv0zqqF4uSmS7F
/70WyU98A3O7RL+/dz0QhSS32f3ODwABDsK7fwqA+xibuiGrwnX1uULMLN9Kq+Pn
SghR3hYzrsRikcPb0oDfFBDfjPsWJRv2Em5WH/Ug/RTV+Xr3unsGhhPyoubrNZKE
Sherg6pI4H18jTbpOTaPdruojUYkFKtwXTv9ATQWbYPyN7/R/2+pHYE+jIEJ0zFB
EIeyAnWeULAqfkRN0rEkeHpDXPod5lqxHL8sYkApdvHU3jfORaoFy5NmKK0qikBU
9GXiyOYrgQjZTB8yOgXHmjqtSfQq3RDcJmn+7zdwx7Uh/9IBs09dtJRYbved3sDe
X9d8WiSWe4txh/qE+STdn+KvAE3aNeC0nfC/nlHRjaeNcdngNETM9fNMdsDli0Uh
i+NM7YquisMAldNBxfxRXWVyc86E+Ys1eIeC6gjYSbI2WSUDMxUDhsWt8sj0Vyes
EOK4nrN6V6AjhG4BghQcn7d1+j06ZrCyYU2UPfsokFWO9POovWnfvQx57CrOYt6u
jpdXxtZ8iAuNyVTK7hsWlLnQ4W6Ysb0XZ4kab392wSOtMSTMWFnSwV9oqoeQpO5q
ndN7BDmPzdVEi1Du+BHxtHT3REPpBmJPk8yiGO8/7k/CqQtVCqWjihalQjuWRTth
3fzSOqyPjyBk35XjoSWreVjT9A7HWJaGM/NwqpuAfs9oUbl1GwC+QopvBj9aXOH5
P90e4FjRvK6RmZxexEHy+BvNKucY4AeMPURFSpOKdOu7KmiAnVqyfXLD81rD8lG6
O3wTS1jRI1/gZyCEZDLTEx8nDLBThl/n+tdsRkIEHNzriNGPZKB/OE5f88Gyn4O1
dPv0xvgTQp4XLvHL1cOCWsNouOks117AmA+hUKj9U7COjo2gGVqr2iTNniXkqjZE
b/r2ANrrXJXGQTHQWh0ZWgZ6PXSjRceyocHvwCMY6kLwbcqr5ZvvhUWDnbBvDgNB
pNLFeXG51MwJeUEea92VPjMrLOToGIIp/capCXw6w2RiviYSB/ePXbyYla3V/RLI
MpkLWbtoTJ7nCSe9aiHcy/KVwNS3YXTfvsv8C7OsiInkEYVxao3t1OcQLYY3fwH3
0X6/okVE9ugNtvGXcFBK22yOG1Efe98+4xQ5dr5XjFCyiPoqJz5X8YHNxcdHOQAv
GEt9uCCJfKEczotP8nB4OrdQNkvQ0XvDMVEz513QeLPCvkaEfrLGa+CL77lwsn1t
ZpVwmY+ekss3lD9KnsmTgjdjkTfI74mR8iGacbmWew0491FarD/oxjKjrNFjsCNj
5bEpx2UxOZ5jnBSdybzbkPTb9InRl4ZuagoiKjX/Sa1/RlsbphYB+zzz7985cSKK
3f/lplxSsuOtg8oN9Eu22QpcEvndNsKQcc/qnnjBRK1RCzPGC40gerpVsO3Bh86k
BpRe01IpahIj3OjSUcvOHRWtFajHkBhqo9aB/EDzLer+rpMLo/xLfROK5bl37lpr
47zFm+BoiO36PsRUVOUehOFgO1pMyLi4Myw/iQeQtxTBQzJMegkyZrXuU1fsRzvE
JDiuNUj+mJUZnLeb/MOmcktY1Y9MG60QlqMS1igKpOjjfP4yr2qO5BB/v+qIDlPK
fq8AmJFcjWhTUk/mgSH3fvBlIDEi37mzVxqIqNvdqvC9dQn4H2vpR0+FjlDDay2Q
zlsyPoTbAWeXrGGc81uVvqZztF813D6NEhHnQ5zGXOTglqdYkyVM4lWlAeRKkpxw
gddxq9paTbOrVL4vbZIsVw==
`protect END_PROTECTED
