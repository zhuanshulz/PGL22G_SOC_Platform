`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gK2CiBTaHQWiCaoLDIPJEOrtTFfAHpw59ip85sRASER5hAm3bIEFdDDwMg9xwu4/
se96sYT+kBAgIlCafjPnmvZUK5Y7LXSm4Fi066kqlS9TNFMhPs7gHNqJthz2oX/8
6W7JbHEHiPcBQIOaoGUBai67LuUTzVOuu576MnnwOLjO+zNoqxtJUeUYf/v4FZfO
LDx1NwHb55VpRIp0rLrJpNOLntKu0zplkMBt7czms/4z6d6l6TJ95PRJWn77O+DA
iDVakexjZWgdHPuH55DUn/p432WJxYMDOSteWYCYqU8kLp38wu687BAaAdknih6h
iy+dDRfYR72CtRhPk8kx6hEP7MTNXxZAz8nur9NrbIvOkSOo6t7AGRLNnEi+H11u
oB83x1t9oK6ku4PfUQpdvO567p3/GiO/H3dllqeTqLE4qRHnAn+PeRm1EfgoMqCM
1ae9gnqUt6bcl5oWP5I5K9mcMAmZ72TsOTlNm1bQmm7UVQXMZdOZLmw528vF8OiV
NYNT+Sc5YtMf6PkDV4mdj4BewMk3FCQ+bcExyiPwNei2uU61ISNESbY4XgiDUdZ3
BRzDkLvHoDxod9RlIa98eNdmF2/UChX84+q72WMO06QUTrdKHAPKOfFG9+OBcXnR
p0SsCHHd4gIXE4noODXVK3aBgv8NV0CWg3Ly1JoOaizSqSFDqv3dK1n71sWffYRb
Qgth6/N7GA1iLyukZtFQ5X2lUHsQ+LHTkwi1VEODi6tOxgRl0s+f6VBZic43iYMb
6mNdWYsqi05H/PD12ASpmq6gzwBvBp+lySOfZxZkBL0WYrUsLI9SM5fBau8qow5w
yeA7+MeNoeDrsrrpZFYSNYkN0zFkpQF3m7dn9/ODvgg=
`protect END_PROTECTED
