`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G1/tPE2CTZHLEuESl/EGfhaLP9kPJyVMK4zqG82KqUjltqPtew3mzEhNIGvBtFIM
ip36a67el7OE1nm0L5CNU52ibXLCINaDW+kNSLf8iM850ENJYNVZpyNP0FbBnRuX
UmMlF18zu7FWc5rd0cC64TQK7XZHAJ2emmIx/Bq+r2gkA5h8ItPR4tVB9V9uJRre
fpGgWPWvuHSTBb+Z5viuwouvj7WDhemWyJozqr2+nd8RtduPJIR8GEs+IrrQxTOL
puRILbcI5TnOyzLdSmTr+EfKeAXsbi38FFhYNRm30P/gglza4aVwh4SqaAF4PbH4
gIUEH8TniSJG4HvKALzljQe4A070x2XFuyAqMdjXKZyGxZwnAnz+yrDxrppYPPGA
wWEAEsqVDT9LSiqOJlO+EP6yfpfa3Y1575wYhgbs9zrpFkD2Syl728CXrG8+Uek1
sRvUY9iHefxuf35FXhJPZbSoNUT1UjMr8rBrzEo7vDTZA7qProh11ch2xsXAtBX2
5WC7CPvUVt6TS9gvtLnHiPMWfY43eEZZ70hOa+gMP21bxFgPNgoATUtS4x0Kt60H
l6TkXhGkNxKh7lOBGamJgQ==
`protect END_PROTECTED
