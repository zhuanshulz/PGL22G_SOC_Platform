`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oenY91KC+u5yJHtAg+KUPBefyDfYsEC17yvL5aKtB+kUy2/3JfHJn0vvpmvfNVMe
zvK66dbynrA6aWVwWC7lx+Sqr7VZ+n9P0U/q2GQVFqSWRhin4WmxDrGA7Jw0IXSi
IXcTQUTNv+HFF3/+9RWOZSx5e8h6FI0jfsnRKJyPhZsJUYCNfE7ZWPNhWA9DkJ1v
vAkswFm+moHE0Jq/rztJjTsLGoXJVSyyqPWSzB8t3FKgOEGf53qts9qPlcw6Qeo+
dlBe9eIeXuHNjZFv/Jbt8icYn4VdNLMZSZ/HhXTE9GaJq3UjOxnZWLJyBF/YJz68
PJ93YdyOMp7ZxzRS/VT389LUBQkxlwHnr3NfQ+K7OtxNvdgzwOQsSq4WOW7HSfeo
0JUD/SFswlDcqkL5MBByuIqT8lez60p8VeYK9wK1s/xVnXZZCtpGPKMbJ0Cgw6b2
sF9RmUYSON68BzmGCE9y25kEIdO0VQXyZIv5fd5ptI7SuccM9LhcOiiaPKAD5jQP
LhR9aadGawA4WrMevIjxMMI63gi9HF97k8tZzzFxEN38Wo6UiaUmAunWhEB+I9hr
UkDd2hEwIK9rr0/Xv1IgmDv9bJiDc2kgucCi6+bhLWqpvOYXinUGoBByjXsfif9O
vCTXILYvPIRwjeUhtDLIkxUgnW+F71DpIfILmX4uKHZF8Z97jgbTYRlCFAvPjDCF
jVpblaOg10WoLsw/k4WPcsyjbrSkFuO9xmbExKQispE8KiIbf9X3SVsCSK801joT
5xBlg5enZyAE+jjzjjswx2q9TBFUsZ8WWXKGTqSP0+1Pzof45b7kr6LptA3o1R5T
YZq63sF1owk9cGPdxCow7L1cNbD+fCKxUzzHgVSGbFdjrfVjNffR3w5vCHeq06iz
52aui+InJCYZ49iOn5bNj9tDvVwxk9C6i3SEs4Qu4EjSkKZb+bxbdRaKhRlQd93L
MOn8Vu8VftsjqxauGv1pvRKGAlsXi+Qq5mKUR8pKAw5k/7ft3e4kH9OZfCKlStuF
4bzFtS6LeLWcEzaPRfGZzDtvN2+2N8qBCVJsiijFJWAa5+Jlyr3/XKKxf2FhdiTT
ZFQHrFPRO+SoibTJSLe2NHMQA5bw55E1vXDorw/CbaHBn0MVkxsDlrE3fA/Ubn1N
h4kb8b+McbHWWvV4YZkT3nEcv6aXoOzvzXY/DaihIxRSYJRj9sLzSz3qsAt0D/ju
xvteVESD0hIwB54gTueRBefswap8vxz8e1UQ2qctx1PsFxAZYBvbOMJP6bgyCpYm
Ax9uHRKJ4DTHIlKk4Xu752jluex9oDBW1UzSpFEuTLuWfDqErDkwkWhUg/Pvp+aU
KjfSHAOxrXuaQIM2oDG46kpvR+P2pbutEFnYl9nI1hjcXW+lvtBwiT1qRWGiuRRo
kLxlXYfP8KO1Kpdqei/hQv2ocmk5tKocQlSQ1AOEtZPVlLQzGTecUn9vyd0Z4ADQ
xfZ5nnyIH/a/lTM81xDbC39nUHduMLgCOOAimlrvVv+HIZltJMwl6WIHFh1DWUVt
Z0fWg1qTp24JFQ4iC1ITUKO77z8c9gwy4P/xNy2Uzi8e96OEbm5EHX0md8yp6fr9
MIynDl/JcBrM/7/8yM3CEHK1oGF9SepJQB7Z2qfNYzLdY//lnckTOSuucMXzee2U
pDAXk+5cDx9wy+VGRDrkduaefvGUrXDfo16tm9NyT9f1aCDfYfYxFn9HFcM1IjgW
TQiYxBmEItBGH+CNfN4egtyTsG8wQclDRjXSDSJhk0C7qLi98BRlgYYWK9QErtck
Sy8dKcGBGGcpA2+J0z0gp4vnIhbiamJq0+ECVCORTT2Q9dCDMbLHgZr6DZOfDa18
VVhQHE+43zTULlWf+qYfUIo+ZgDTpZXdzDRkEiTDzyIVp9tWLU/FELt28nJwTKuL
Rl96ad816N8f2oKBhZZ2fdJBhAGQNm+KyXX+6slTKMVUTqWvficvzNAcvbq6wPfC
jPpg9+L8z60Dnu2Ly7GdygqXirxs708G/GajQwkjajgLwaLN6hXP+o8OWDIiUpFj
1nQabA2iM3Ztd44Qh0ZkP+y/JNc92FoOXxu/G+Wt6njqZ9Or/RmbetX03iZlHOtr
nV75F0oEEbAN0l/df5eUnIcmuLOiOA6Vrh5In+VPqYNMpl9Q1GORgYQY/A97ObKV
UzFrykPqH+I1KP8CejhjGCf0Ng+ipi94975ardIbulJ8QOxErc6W/ErkZTlNZMbN
swN85GjdSYPdMOS6LioAj/QpZ7YwWe779JHBcVzasgenI1xfN8K/CVUGlVATqA29
4Q/veAYv447aAe7z0tN4RQ5SD+PsKgpx0xkkhFK5l1x4T9NoaDtafVXZ+DhfDaua
UtG9xXpY3W27GuFYWD6gyUmO5RjxAbXNdpjA45wlnJXlqJsgneVk9R0Ge4EXia6O
X6TyDUpYnYKoxJRmzDRYGLZE6Zp9iuQEE4pSKkL06gExhUFHGfOGgxgxvl+F5Mp1
CNUF1en27+/Zdrahica08SUu/dxdtWNDGDMbbrG0AsK2xofe1CguMVAbJW954GxU
cxlqkMNp5112yk332eayFDVwcpyjYqqaSCXJrXwx3/XafDm0wWAw/Gux5E9kJQKS
nnHkHTMf1wrUxiEUNwTL00iKbOB1Uw6GdEizxEWx22uJIQ82XcZnjJaJjHMdZc6N
JbIOaNNYRgQYchMs+XflHKz0Mbuq/Kknxy5zuw/nZbvDUj623g2tNP9Nmv9eO3ve
VxWvpHYkb19ybrEaE3QynIsUG5CFa0NqSPVlNPMuKNKKzUREWBjpaFlGVJ3awUDx
xBbwHGTOe0wiZOEo2jhKvMf5GaLQNJftfhEP7oNi48EptlV22De5gNDRHIuHKkRt
`protect END_PROTECTED
