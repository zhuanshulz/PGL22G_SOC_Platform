`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUt1TDT+40vXH9phBraHLB6cAupuw2KJ00KHNQNpeq2xHzqKp/WiGBeOUwqrUalZ
GB6DRS81Ni8YIU/0pFF98rzl43BShdZaiEEfRktUTl6bTenus1XdGcvXMniyOoE2
OjQAeQvh/ihGAUp3NP+sz3VxBtd/RcEsCnYi7E3Zb0dXzi5N8SW1eO0OX0elheYY
ijreNdSDQKzbzYzH4kQX9MaMRajutqlPDt3oaL68yrTCS7KCTI/ouVbRuMGHiS9V
+ZqjfkHxMq/tBoHlABJaS1BQKRXXyNrKoSz6b5zKxsP6oodxaGH8oMQHMh4FLi7S
OiV0vhcRVcXE1mJrh3zEbqupSdmS/UFq0qmAh1NCDvRFUGaJW4x2eGg+Li9+UGTi
wVynI2VPuDAG5crnpfDK0a8TvmnxjV7mx2ZG7im18PNZMlAWH6gMCI9TLyVh4vSA
Lb/WunNDohxa14trI9l8ZMdzawKVlLbUVbVQLU0rHmQb4qqrZNqNZD9vnChgeJe6
o8jAp0dCh4HHaQ703gxmy3SyuVBI/AXQ0WBLoOLapbaodiKHEeyd74Es5gTAbYZr
Qi8bgBCBntHKKNJIRFtt1KNWvCZIM1CpKYIs6ZydHrZX0Ivbsr6lWumAeE69QEbt
rISUXoVW4D7eePFdd3ccDXM7D+KN6c7nr+m3aNWigWaI0TDbdoNyMnHdJPjKZfra
xGV33Usm5FLPTSZufZmlkjaRvXpBTe8zvdV3/1jHjMBS7fsmhThraVmzFfNG91UJ
uvIZdpjMs8uhYHEeumfEaf2tATTOw2CSNobw/c6/3Xj6tYgjai3BUn5mUoZ0Fj7C
I5T0LKc35hoGBbB8G58lzM1pWaTCKUocwev/Y1UrJqZYHby0K9OrHgpTIUohGpVn
T3XWEhMOCzFiE9sXrg1/W2XHlzIEQUTmCoWfTGK45D+HJtK/b0ZCT4MHIB3iqA8M
wMOy0G1VBoJsFfmnCB5SO3h9veIz668EoKOKt9P4iAP+KK6POUsjy20kZvxaYGpA
AziCi53LrPi29tjPKzuI9SP3W9G3vIaUydG0ITkBZzzsiMJGmYjWIM8i0jzJ76Z5
w3sfPYy9CS5IFD0VF+KQ2Fr7gquZaIYUODMGOdIYVK6l63wXPZeGxSsPBGSyGyKp
aHwv6DZC5ouJ4ubs32jFfXzt6V79Sy5pYguWbVVIzCJmxCwVSx5hghKrl3X/xVtc
grfC0A3jQEYJf9EhHSOS4Bd+KM4ARtuegfUFDeK13/AYJxdsOpjA2V4fQfOWpg93
2KYr39TqZ3quKLX5+A2Vgi30vTazDwDMEcSBx/d5OoTrzZ4gwHYjKQcYZBWwLYxI
yDJNS/C0qOoJQjcaxRL3a5zdUIZFvISQp7M1W6lOH0+3HyR6V28F0PyhV71Te3JP
TIImLRdiwQt6x3clwoujm5oWbgR6Zy01X0qnYG1zv5hF8XuKCqDkA8qQ5vkPZiT0
BdMXGV7rjmXNE20kiZLEP/mPauIRA7azuFJvHsmm8j65MjR2lCgZaZDYQxp+PnnS
A18ma27PS/R8hLeQh9JtZ+sYLt5p7LJlo34rixiQn4HHh1tEpI4W0KidZGmErAkA
mmneSgcQTK/uD4iRUtbG1cVubQ9ydho99YNidf+ULIU0B/ZU8YM/3KP8kOQIJRF4
x/BhXv4L2WA1Hp5vt7b7UaAq056eLKO+Q8I0tgVeMNcznmyhXyZRb/xw9ewqXVMG
awbgDwpvegZO8EyL+/oH/M3868IIv2v4iU1gbHUUGb3boBxUc6JnUbVeiyF/uwOS
awcqNX4TOzWa22XZaMcGZ5m6PVi/ZSEjRZ8vJLP2fX3BoyH4odykJCeRLJ0m7Sv7
vix5Rzsznuj6b7e7ZThNDoJ+wmb+t7dwCRZ2HA7arWjgSCBcw4CzZj1JsR6EPzWi
TQ/AyUrspvlnHXULMjVuBYzFaw4sof1X46fo2L28YNn62ZGalWHoCQ9HfaWUyvA7
KEltFIX7T/BCXkW7s/zzutMWMmOjzV13kVZgWLdT+q3C/hakryJvwbBFtwLwq+Os
eqy5opanRlCl1hSTFRj8C+6ogXffxCghpqBQ4/hN0Xl+AHPFdOwoz5tKJGJ4o3Pa
3fbEDy/2i2VydkpsiFGHhdB3U1SVxsRxvjm1o2FqgpDZr/RbhHCOUCTo4pgattQq
iTszMzjkiM5YrxTNa5bFa8BAGcH67oGr5nAEj+D3ah8=
`protect END_PROTECTED
