`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWqB1qKBfp1fKTopgy5qcji61VW2S72bTaR1RHCdHn2K+Y/o4u54NLmFU0IZPpch
jKSVOh684gEkdNymzx1/4C7BY0auETnNK4ptdOkg3lB8eSDIe7OFUSgDPdWqejVh
IWXDixg1EqL1IGFp78sSiXnKaH81hgGzK8bnu8YxsiGY9S2SGNgBeSIYmDugfTd3
0XtcbSdYb/6LV2cCFmox6yZkZUY7O+Knt/bTVQKEDNg776MlaLteuXTBDM5sgUHK
/KPloqpXkURyptEYcegCc/XzldzG3keAiSMsqa0SBxWIxLXQ8ACNwAn1NE6W6py8
HuIMz7FTkrANBr8KaH+qL7WB1oUmPV0Vr24nQehZ/T28bJBRvy15YcSUYWKwR6UV
q3aFEPP6jBdtyMeTIomSw/nJfTHBdqS6fm9rnm/XzEfKoDGoEe8zRsWCLGEpTNPg
U5Xkv0jnKbQFJ0VecfX4ZM7MuVy8FLFks5FIkUGSvaS+y/keWJz4b2AZSpzsQp7o
MHY8AfAfCiDqfhL9g7wllt7DLIx2dvHb5EOLbggZrLqZh5vofuRbc2H9x4KOSpQe
AeeCEcvrUrZl5obo8Sr7ZQ6pnH9He/UpzEi03lGmMzLQuB0CIK9M8gtZQ2F2oGgA
zI0kD+zjyYH58bdgQGFcpqJdm4ccoWLkji6EyvzFDVs4SwRr26NtcTRpZzw/uf5W
lekKwVtUOChccBXVKxxkQ4qnH6REkSPgp6/W46ebSHiWSEjZhYb6gP1o2PWv9r+k
MuRJyttWUrcja5BAAXCc7xLkhwUOTxv6Knj8GzaGgD6OREiflSmBOoGk1swHr4R/
Nu6r3dwu77RAG9iN8K1XOmD8JB6QcXs3e0PEqaz78AHzqKNIlNz9cgd4UW9l+Rlg
`protect END_PROTECTED
