`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pt2F8C8yPbxvjc0MSU6K6CxWLRDirC1nBThGwtmyju3kcBMUH/MXBD7BbSqQ2dxu
CVx2bZa5D78ktd2+sCb5Loiu6wI5+jLZQHhAVz5wX114URQu/RzsfxJRrRoKzdS+
2tFG8ijNpHQP+Z21/aBLqhMulbVt6TIxiqoLw5tpCg2xDsKZI1ZFEDfCM+9FBDg/
IEWniWkQ97h4ea6xW7X05yRZYLmHq0AUmuhRZOTS1KgfPOWhxkpnDKaczTzNMB1e
bvT4tm2uOxXjXo9aQAS4FoDKNZKO0hMUnBXPtywi/k/KLTLicVrN/uKK8BleSJj5
G65FL7ZQ1R8JCKooPpNRR5jgkkyrqNbyOW2fPxMP1/MH/W8sv3/mwZyI7BOTacxI
cs2WluhyV45bZnVpKyIShsuLfpCKh5MPBLwA2/kc5QgaUfU+r/vRchfoGo23bG6P
Kv5GBBAVCpKTMFc22TLaiS1kLAL7VKHza0CkgY7igVs2A/Gq17h4DaioEzJMlWhk
YL1aBr1qstklxMxQwTGWJIuDjxFuevGSK56xgTQ6287N+OaOOzUc0sqpcMaGGTSK
LcoWabO5Um9HsNnWjq9u79vTSJkjaRWvYfJNUrG0Kh8vX6pR7S+cqqQM+zQ0K6LD
cFOnEZNfqXZjCbSmioazMa6USMXekWd4HBoAPD1Pp6+e6/1KRFz5AEcNlSkaVwE3
JsJMQkWamZDo5CNVy5qLu4OfZPAmtuObIbIjRKcvt/fxOl/GK/sbDi3IvWprsMH7
Mrhp1lNFxdHaR96Em/+wtvd+KHORXRCTGI+XFpZktPw6uhi0gXi4MilAOfg7cakM
hwsc7gPLj0H2XlHlQxi1poy11nLMPDaLax1b9T86LRJ1MnpdvSHTHvNjd1II8d9p
q5XBSNac/F+8T4E5D6mEr+FVO8owwqk1RhnRY+RaeQnAH7f10VeMarOxRQ9PCgiQ
Eu8dHNq+ShjJ/ec42md84cjjejOYtNtohV3+sRhsiEguc4MuEn1WoXKzQuR6la9P
sfM5t0uXtrIfWd4CkT7Fp6OnCXAR9+f0JgkFVledL3knNA9gJ/O/dJjfRb/zlSms
eZTX+K6cftQBOFCvG8iQtA81eql8kKBhzJCVvbKe++bx3pSHiCnN5ByHyCR8kXLL
dvLjzdGw6m33MEllqcH31mg+g+luLdJUEgoiPMcktJzB1/iNPnfKHrxJhmIX1/3G
HaNJLAxX7ogY9eXwXU3jUFrbVHrWQ8StcyabkIDFT6mF7YgBwTnwnG9OC0aeK1p/
cC1UlSEAuW2DiJ9LoFT/wBEoF9cO7qWm2wCYytrydAuFSsL5matVxIdWTZtRwpJJ
9+eFIAqEYOPTQyQgtR4kd4kqNcEG0GNxv3DbKORkY/B1+9ZKXbWEx97Jykc/uLix
mMdaXuxEdXeuhXbPjm7bai8l3B6CjoqGhdcU4DUKhSO9I63Oe0k+BpcbANB7WCtC
kZyrH6qH5z2nbwfvSCjC7r2iryoNRB+yZH0M2vKbGQTwpdzg+yt1pHoyE57KzkSA
pMN79aK3XiYWaVzvYRo9SFBjdfbld1eyk6sACHIe3DhdrtO+3EM68QC0jynMxDa6
j8vjisK4BkNHoSplUKfyzkc+CMlrq7hJZS7yJwR8jjepg2TUnQCe05f14Pzg/u5K
elSjZ7PxDJEKCbEn1Lajqi2CFS5jro5N7u5DsKvLMU39Wl6N177bMQDJJl8q+Ery
WMUkY13+IQFuzpd94ONU5/xcqVCmLOrQbaVPG16io7llz+AHMTkACf+u8jg8bVJ7
HHPh+ydzVa3AZpEi/k6T/rdy552g3t54DhpHI59jCAF3fSued2gtMoHzpRHrvrWP
7RjYWN2yz0+z+gespBrjDPJKlQNotgA06whfXjL0rRL8O7CYjkxT9ePotUL6fmwI
Bch5LsP4KE7eEZCPiU2iwbT4Jmx6QTO434FlAslAOS88306uc5Yrd1P1Jf51hrU2
XD652yw2dr8qvy4coXhOQNIklOYtPcf3W908MdIJY0nWrk/czPlm92c8bpPLrESF
ElEo8UGgwEX1GL2TJv+7D0cbFzv7W0rAR4q5+8NFhsFbGqi6gWwP/FaBI5b2Yu1+
WkDY63uGSFYAYpmTu5l2fK/CJDWcygtwnN4zadch1Fmijy4XKhpWBBEdyAN++s1b
ZfRYTRMjP4rdLzCKdjAWUsXLX6GIg69agg9gqbSJW/cZGjzoW10TPeBEDkcwwTKn
o4q5OjLf82dg6+phrYpnXVIibliRCVjl+HBM4dPVsq+LoPPcMeGYQIo4YFE98MF+
OG6QIcFuzvJWAAb/+7fxssN8oxjYFPulC9GoPHcQyGDVzmxekjRhRah7n6pEHyEh
VBHRg3W2dT/E+Dxr/ulfZHjX4lAkUfZizyCt8t9BxVnNtKMEMeAalpggs5ZF0zOv
zGZwoc1ZYyUXSLBkaYSAfWJfH6SWcBjBko+THqgvB2GYi04C4tnpms181vg3PuVI
LkJ9TLuw+HVo4tZxSRo91273aIrTJLUcqZmpA22l8TRu/Cp+G++yi7ALjU5duwbJ
tboJ0JiQpoyrAZDcKbvgTFUmYLKLmClFXsLOu0sFotB7Jfn31Mqc6axkt1IyMXTf
w+2S446lTL5k1Jt4AGLnH96xTGh9rhrqTidgwrq95Rf1HToZlv/E+eR821tjX53l
a1PkLnv0fXLsEvJiXfneQoh1Cl8HcEUUCUK8X2yeKNZctqqKm8AA9jljSRw20VOE
Qg3kO5uqHY7AgEh+YmgOuPN0RkF/LPK1LK1jmNvx70DGqtimoGCeEm1KtULv3Vue
lOZKndUEHqp4piM1RGEdzvl6UyJy3NqJ/UP9fyaQeJ0KqgpdLly0tEKqYBQlIlpz
6RrWu4PnryYe/mcDzN8enSnyo5i8l1qyDzfAkV0jmwhIuGa0/OLXIUyc0EEQ0Hin
z8qLK/BheiHdbwmTrLC1x5p9qqkXx2sVISTodDQrQ0khyjVzJJzG6QE4Zf41TpOF
acB24w0Hsj+cRtbptEfw2f6rHqslPWPRcAIDr+mjIWbtR80Bvu+mOGooBBSLWDMR
qevctTwV6Y2qOZK9P8t09optrij6jWkpYDUhR2NHEB+xqJI9QoEZxMnoQa32M7rx
Purlcep1lw+ZayVskYMgAQ3X65jVxDN63452wOTLCXHEBhPGKNrGd9Mf/GdvOiqO
PVmlV+FsLqLC2AWD36/W3HzdYGdy1hm6dOfPty+JCR7wcg7UpGZTprBY4vi4MnPB
zCOyZRDl2yZrdCsicI6dt/qmB4Vm5zVUdxWiE6mpV/egn6xjYeT0hBVb+I6E3/q/
hR7YgVDIiKoyvOOpggkT3V+uht6S8SIEM/gmmykv3Gzc6oiZkPiCTfdppDhOoq9h
/n84Z3M0kWblavO1JCUvA05ltPDSC70dHXVcqHnUUhsKLQAhmAr1x7YBdOdeveiE
Jup5q99PgcOgkau1XqXcjlIrq+N+Rptlmxvq8x2RoQ4W1VLRGRt2Q41SlTIH9FGW
UG4W0DeJNR4sOqhd2old6NzowTU2R4Upr6P7HaNNvTL2Wac7cvltHFBwzNmM5JFV
RVJQ4hZqOSn17zWmEEr7p1LI0kQxfqNmy48+H1YIbnAceFfgDKHqpFyD9jkPUM+0
OSQLACIo9SjZiMXwIFeWNj2VgAdbRKddk8r01f+7GgfXNEjzojEjSQ0N8FJgyCNv
HYZ3kbUKMBNkk1Gf9qRRo3jX+neBbPF7lwCrGrFncjyuLaoEq7tToDO0VZbytCyI
544kurGMG8CH+P67kaxVfIi1IAGgDyZrG+XWKwF9hNIMYiLMXwgUM+HQRoKZJZbc
j1PiQ/ZxaeAJ4BD3Wl/nLkojo4iFnC/LU+j6ossyaPBMoybirK75Ffx/+ZZ7kms2
tGoJiSm/7vj60E1HQnmtXCcAk+m61tn71hK2djv+LuBR1ONf4q1tYIPZ45qOQgsg
+u7EjJMDg+825LdH0PUZnor1QzdT3aYqQpRFL/kceR259rrOhi21yCuN76wtCoal
o7kjzRhNWVoYOauVHJGhdI+epQIv/SPkutegbpb84b5sQ0ahC1N5ts+s7j3I1blj
8dqRbkrNHSsue3DQgUIkR9iBQIw/gUvG80xPibt3zy1f8ErxiPXdWRbe2cC4HNeb
/Fl9LqYUgzkSQPLAChXq9dBkKzJs11BQRVZqLoMMPrutr+CraQ7AskGOj8wAYgzT
kWZg44IPi1Z+okqJnOw7Xzqbu6xO/ocq2ld+sVbSVLTVH2PR5zK210WDBJwv1aJy
T3Ax0CmxdbbhmzHeoQEc5RcepDhFVZpd+R1hPF5zP2Ksz3rWGcNErgV62/ynrjAH
WzWRKdDWgVxgx0DktBBwbS1j0cjQWo1AviK9rlCxT/yaJh/WWUxgBgAdP65N2SK8
TSko+9/zGf2ywuCCIDmvZRt/xt9XbjMtROmrqfZBiJLLCtvLFeV31jHP/agZ2diI
mC/9La5YoTxtE0lKEnG6HM+EKIUrbsizM2rGhLtkQoC4ZJwJIk15g0CMi748JA6L
FhyxRiHCKj47ZbRi+s09n+RNHqgH5+uSC/CalZTtpfinLRsY+6/pOKKCFB4yQyaK
MJ8FX6hqzNh96GNNIkshqTOe04V88oCD1oTHM1MKejgUWaM2/EdflqHhLs/E5zb8
gT18l05fjHVCViGj5ZnQ/tRAauSGSqeFJqGrp6Cswt+AiNyEaXwKwGDD2g4cRpWL
p557tVavT3kOUNHbQtIIiL0xXy968uKNDtdlvm5FnLzMLXilZlLwyCV4etzGL/E3
P3m7K8n+xbkmxfnFFxRrV3JEtlMI4a9t6PUfF7MxnsUnQUeheaU4N4qAe4/IjvNC
lGL7MBiQdMFmm4cJGtYuMG/TWhng8d6y65OBLQD1vjJ2SZIzVCYxFXBv+Y64TgRV
ODTj2dnZWCyk9fnDCOFGks8An38yQiw8lTm5DHP2FZnKoEZR6/VvlLju8qp2qbSI
tdUpIpx6VTO3SKdtr1AnkyhgpGrsKVlkolC8a0PDzbOCPSgZ+95jSb01a0pkwk3p
3KMubteY7ERhhp/cYnqyRdulLyQEFqmVl8RObvCAv/YefKRp5p/5cit1hoArDxuW
NEcTipdYEYNM+84I7PLCNTVRTJbfw19Hghs1yML3hGKHTGy14Dck46mS6Z/QD2JI
cvH0gz4Zhb76ITFq5+BFEj2RemfAZ+ZGiXIH5GkAFCGgyM1q8ZGw+cUjjsFfJHFo
tqoReYwid/A6MquvH7hRCG/zOS5WCHb3LcSaqenyIvqegyYx+0if+EDodeT9c1bD
S6l5bRxW/2WIWGUCVhvOhPEidIBcX9ncA2ee3oLLzA13OIHmRivuaTfGLACIavIu
8yQRZFmE/sAY3bLwzFPeZcQE4N8VZN50iwGU1LsQmqcciK+E/wp9cYJ1VYayLvxz
wXFDs4KF9G6qkReJwbm5vbFxER77Z/7B4+D/lHGlopjvu/ZDp4nqFEIt8jUo6Dja
Dn7zRVIbYaUTgns/Be3D+Zu2qCGxMubhheFm84duNQbju/jb9xIuAk2tTJU/id5X
VCoU78lM5XYeyVJW4egKowCQOzcMa64mZQp2g/Kcvq9pFcvTtHKhBMqmblHLa4nN
d159XvyEgaheLQTUoenudPhC+raAn9sXRQXkBeLqdvW+18Lw3kyRi7kgqdd/dYob
nkwQwPmiZ10n/7FQKZ75HjZjwoeSbUGk2jYRs+Oie5f7m7z+YYe288xkJmQMSTql
1ohtKvYmVVY7MEGFp0AAHoVM2UdOm03bFH12DEj5/jrbOSdSTh65/TLMJgoK+j0f
sTsRrmaXxiwEeYwjwimZNY4gCHtzMkopNTBvnFDS0dkjqTFYbECNjDoG/9Ugf7Od
x0/GSgc+OHeZFcNMIUFA0nSTzP5DEQU6sSo5jTO4OIqPnhNHGj44QzUTgJu0EG8d
MKOVZzFkvVvPIO9HsdQxjiuzvRE4YdtZ0uGka2lxMj5FOceZ6GEuaIfCU+tjturo
I9FhOrEod2M3XNMn2GsiMuD3I6Jo3VSrHhZiFrLsGqKGPzBbltOvgrPbSYTId/77
+E+jzU223Ewxcjiy34SnCwNRlYA9cyHDGKs5kNaQkhJh//oCfn/5ItCLUVE8Caac
pjl6KqLfhq3aMk7KbVObwGN82l+uN/KHmniK5aSP6JSVunsq++oH+ii7JUEj6uE5
8h6t0YZtxAF8qOeS1XNNX9L8g0jMeNcZdgtY8xG2qUpW4GkWiJMeoop1ZVJTFuIM
iK0cOhIGRZHk0iDCG64N2OBuD1hfkLQeP2LTSIFtLiP8aV+kqDeFtKhA8YjfD3sG
Y21KpLNeGCBx4o83ylxvBEnyFx97w6bTE/KR/QJ7FK0U03Ay0EQtcmtz9KZF5jmR
UyJaORWakGwK6ZEE3YjDVNc9luF4wSoIlNd0NrMm1RP4orzGEGiMByvqd2qk5R8p
yYaIFO0cLqSr2KkwNiMWkrMmTKAGtT+AXb3DB0SItcjfbvTkvk+cLbQtxAHqbH5r
O0P6Mo2A1+4gyHkRaBruUOsMz9Wt0+KwmWvf2FwouOU1DkCiSD/jFlXDPRPzTyg/
zWwnfM9wf3wGBS2D/TywnceTQMPjxDTPHIxBwghA3ql/sNF5REJtiB/D/8v0SQKj
ZBs8+TzNB+ncBGrCiBDjvC7LRACGzAF9ks0RzUWXSCzdDIi3/y2oXiowes2reFTP
PFQW/cb/vaeginNFGmsM+H1ZqW5vJ/PXOpqvP8zbMv2RFwvJPH9VMrqJY/fxIv2S
9uyPj1FQNqf3tvdzuEM/kQpu24e1DQfYUD+go0EQ91vGiFpgip3h0zhKLKMDlKVi
mizwB/qYo9ezfjHjLhxV5f6TEwxl0955H7z1AFoyRuwaPoWEQ7Ls0z8GX2jpRqom
863gRuRLTgsOvyZ+UNx0jFanPzhTKUr5pdlxGfeW8Jqeymxo87gs16bbtuLchn84
bSK6DrU8TPpyBXEjYCh7trHYsnIbVvzbmdmX4Oo6rYbO3EJDWvxcJP/ZXOwr/cQH
SKPfRLAGs5uAwLFx5meyzFNucCv5PlhZAPHRF6XU6DfKk8tD97WGT1YJbHJspYMG
C+UoSxBMnPK83zXdXKUha+J3le63IuTof1ATFyTeXdrDB4V+gYYV4p2leY7gQxcB
HqhB4po8NIf1AGWTciXIHZOzUrP9mSrptCx5JIcTV6kNybmEPgfGti3F2/KO5P5A
ZsHp7BlD1XFSVCRW1qszIip9eRcg9Cu2MIyRhrfo0hNjnqHADjBz2prNqdsByA2H
kbYvlvCI3EYSNiKr+97Fvj9KN2CeXsB6FXSIXCHcIawsEXeVZLa9kRKqm8OeZfg/
s7+XRCutsajbdaJT61AnlZH9t3Xi3NWZ63cLD20Xi2WRtWpuKljGaf5obiI7Cpex
r4CxuX7EaEVTZnHZixNuVJH70z64nkMkcoRomMi4OypYFFvfgmH0ZiHBg3xII/Cx
6AuD6NnB1+8zzEL+ilhyurQTnBoNRMtvXo3w08IoLs+lcdnN3MGjJdOmpe4SrZOK
6tEMAP7gqgnT8yrBFqEtcSmdrzgOwjUajbkCUx42YrekNW4C4mZVj+LaiLoiNi/r
zqyxFM2odsVksFQX6EH96J+bXyDNotLKglVHBbBUx6LBOqItIM8TnluTF0Jqg0I1
IE1QKPF/7KG4mRbn6kIBjh97eFRzFCWkj31xY3jsRGHX339SoyZWdFw8+gDQsy+1
jdmABi36c9R72bPicqosGHicKwU/YzakyGiCMNHixjX6SR3ddqvqhu9Mi2RjDXBo
4tMJfO7+DlfWJFubuk/2kK2KSIsqR6C9A4oU78JI+yeYaUZS2BX3eE7VDjMMS9Uc
cZXHkOJr8fBooe/IAoIPyJR3IRfkt3kQtFNEIsQAMjBhlPDE49WSIdM492I1nNZM
fCEc5IAP4EN8cDvACgpBYPZzILzmEJRbmrkfCzPeSaTrnw5AX6Ajha4kR9dDIAJg
xYbd9lHh6k8aeq/xjNBH8HTuxBRB+sBdBERyI5MmGgrssZlTp/JfMRnNHifoqh3m
vB43XyoxqH9Cz7dDdjtVa6Md0nwSsOkEBZ+R+8dmNryRXlacfe3cZIyipyg7OBYl
HjDrcVFsYtTBTPAfL3GYFWoWcbXItvSJ1kC+qZ0ai5P77/qiI7EjQPy8O0FHTX5P
5oNw9rgZRYYyPW2Orc/2pw==
`protect END_PROTECTED
