`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKid7ZTpK2IXGvDrEp1fIdUPB5mfBBBDPS2kMxHH/z7iFFH2lk8MEgGekd3qCjfL
6Nb8eMbA7UjM1kWMdzSLGiXJA8DxxuI4StEC/MFYppDsV45UY7V2KSSCOHOEZhL9
l5RMsUyLW8mzP09TzTupm2WP0WrXS/BQ1UJks6ucp5VjcJjJqt2pitsfEwdGUP+r
Z70gzpBvuGVVYsKQ/McFI1E98ORBJaOUZOL2nF+cvyu+WFRdkbtMkwf1Cxk1LBH+
V+SvjoQGuNthZtlVKVg9XgPVe9wKm+pSPAoIED0/0a485CGeVN/E5MAOOYVdhZqK
J1da5ZjLELlmeDUMzatcOk9rZRQN7n+hhsZR9JKWKQazwKvUgMuzxt7tMsW25XeP
W/M75SYNkZGcTvYOV4xmatMYVOore3Y6G2fK5lPbO0Jv5UAHbI6IxkuUq02rjinx
1XG2mhx364Em0bP2ws+AOL3+hd1/rU36XpVRG0PeX7L0PR9UdH9WDNaMriy+OxVE
n1rX7dZjS7s7B4DoX2CWx5mAuwLY/iBGhyGtm+vptNOBPa3BtXdv2n5w7lZ6Ks+1
xbLj0/kEfLcnWUm3SHW5ecaXjNNO6uTt9j5ztwcMlPei+ObYVvOourBTwD4cLiJO
ra6cZYIjlha9tJUNKA+MtbQ4BmmpFDdz1hVsG1Tll1oo8bUCA1IkFBV3nnQhIuiQ
hTTH4xR2VBvweiUHRqMYhAj6EjTipujUPyEhlPjw6YAdeNyh0JG62H8AJY98fkeW
sJZtKFTun7TnMa+ekBqpehwKnqCOyFF3uONPVruJw3cT7cXphK5Eg1dvYzJAG3BQ
U7AcIupAfF9rCmBREOoY6rb0hKuF/VFSgGwXXYGSP1Ke5kn/rd9ZoRHqKrVBGvB7
XWGhWPx31Pp2kVeYB3kkI0JR/9csXB9XEC6vo91ihrPZnFfA/OFhizvZmgBdmBTr
cW2M0MRlbgjTnqW+ckixR1CwJC4x8x4MchCqrBVYWTj4JhEnVLkB8sD9l7kbqxLB
Semvm3+7enculKvlifplKNsodLQSfhL5IgGJjdOM22ymYPrzjvUNQVXg4IA8Ttto
Oh6p/ZHwpyyvdPX68xtYam+0pPv3s5XuOaTsx47fDeV0PD9AYZErkuQ9+Wh9yq8c
EwJMqOjH3Tdbe2XlmLWRlAuVRjvK2bUAT8GGaNUDq0IB5U4hkUNPv+9PuzRqTXoQ
nNA4k75e8V3vM7aJqU5rRa+3wHyrCKcMLE+5vGb1igryvvRlUjY1lX678F4/jlRC
U+kAM4c293+0IOKffr5Qfx9oF6/nh84zefZg1kwjIOIghIyzliVn7LShJo8VWoSn
IzPRk2Evmu4eKLemXwUO6mbClNjMqXVjFzc3aXE/56mSYW2FPx05yx1WEm9u+SDQ
i4HjZbptNODghyupulxLnTSQHa1+44gNF92RRxsGBAwc3Jxy1500PfscWbyqDlqi
MVUR56xUgQADY+p6GbiNr/rmq4HJ3T5xc7rFqImBXU7alPD6VnwLwqmy6HO0p7wZ
5iGRXr+VpjNFUER7WyBw1S9UiFDvyfC4YzV6Y37Xr5ZqsQhgAqIGNFjFNzxfj8A8
l6CiSd/eH98Ee19YtURTSfabz6+QeEtHNpV4G1Du5j65xIeE9wsM3Fh04j+PfwNV
RT9ZC8pS153VUA5rgTVjxW/Qa3napD6Iu8Tmnslgl+6pT1qJ0qRPCkduuc7+6cKQ
2PfQotmS87C4brMkcZTnNLXWPFqFUSZ00mA4ZXrj0tOanpVjTBP4wC8wPW423vAG
Ppn3wuIyaVWibStK9EeVU0S0obKxSScyyFweZ+JztCHIqK8/594F8mRL+n8SrwU1
7ir7KCFJQ2JH3j7VCSAUqUKarfametCi9vHTyGI20F7ZzLhW3Um8lLLB7qFezt+s
qQQ8LhA2CWJnHHUAwWGo8GwGuauCunZIyPUIkIUxtNH9DwwpuHWHdxoO7BuJ5ne2
VYJj7Gb/bLMMfVAW8ksMRU47xx06TWgUJ4m8LYQyYUMMfGhgp/KLHYcjRCpbXn2e
kyr7y/XyVxUPS2msaP2J/XTTyE+eKEUMOLQKsLO0CTsXpItuGlHJwywidFdfyFEk
d14X95Ni3E89x9li0xX7UdXn3gVO9ukxFEzQjQPZYbQqdFNWHJsgr+frs/MbGz/+
Z7MJxpzbSTaiZ76gECUWzwgnv7+pB2cZKEhkRcL4TUtAEXeKNxdq3n8RsFrIAHIa
iyHAd4A/hP5NU+kSzyKy7OFD+0bZw0UxMwkhhNHUhxTRqdleJgBYhlQy40kmNcEi
RnSEy3lg/nssUXxpFvHKEAqC+FmlPgPqs+oBxi1/xNuZc5gax51uaFj+SFztqqSE
1orGexvyRkfouFDJD+XBvkNI3fJlrL//H9iSNeQxqURasW8zGpUqoikuf1fZkJLM
pNYTmjGJ18UXEEowLdvyU2yFl4ghyQSP2IHnEZHXjpFI+8sv49RYEGHDnAQeJnea
Ix4U0iS7BqIG/Njen3j3BykGbMsPUkJYgPjSWsfNY8S6DsZT0sSgIYv+3VbIcqBl
0NBD3P0DGWikL3NMXmg2gGxo57+CVpsggQB8MBJeQve7Yz0yD3+ho85q2x9oVUxb
ltFjVfHWA7CxgU/sml3ZLiT6eErrJjEDCVWi2vJa9tECFpyjDJepe7Fl3OANmB6r
sa9QXJ0YgF3ESGKE/qZYiklV1dApMAJzh5MVX+CzXCspsuflHd4BNy1It69Jzk4t
M0b6NbidPmT9ZCoGJhG+IL8GYsSF9Zu3/5XS54j37HaCoPpbCsnxh6nL65VxlRYA
vh1Cji8AXEsjUGtPDDor1J5Yc87L6iQmSrByZCretuLgCj9meN6vHsIMYQwSY2mi
IOi3osKoLRPIMUs4140Q9PPJ4P/XENeNe+lmHbkCN5nk5AElPWtCWVwt/IYlyjXx
t8IA0QYGU+hvkmoNumXmwTUZMPpvp3NlFCmGAbGOo+VJsljljo7hvvwkzNjflk8F
NBdiA8+1RpquQVV8X4GNhqdot5qbAh6e0s3KeW3+JoY0CTvXuFLgq7oRBjA77c6i
naLEWPc3neuAugdB5eVVAA==
`protect END_PROTECTED
