`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9jsF4hc7I1yFt7mSOKoAc7qVXxWTPof8Ucszxegm2yPxYMu4EurJfk9y0RE/cj81
WTywacjGRq6qhkYnpj2jZLlCnYDhrtuTO6F1+Cb0MDfkyPPlGQUVIpet5q/pXi77
CandwD1DNsQDtEpbLJYTN+H8YeEUn0r1SpeaT3dox6u5z8C2ZeTkrp4lHBl92YHg
y3h+t1XwqVVEDmXCL7hjA+3Z1aXRCkTCBbcvdtS0YrcmgfIkRXPm2ZrWFIjW46te
lx3Aq8XkjjbbYQiFlNQg9qDp4YWnHpBYwI/JoXr5pgtRUSptQCJWzJesUBqnkzUM
zDBHlg0Ae8mLWCvLrd6/oZJzSmlNgyY6YYVed/riIOtlPYAfBg0PYP/bdWjttQBM
MSgvG1mSAUsYJd0fILrkxnAfeGArVnggmdbTtdbnDu7qkmxB84VWU2Twq0z2SpJE
xJ7DVCPx44Ggv2wp6F+ofPksTFTq1FutHBEt1XSPgxi+N96gH8a+N+kd8ZqZLH+v
t8mPhRkGFHoa2X/OZSh9kc/vEUlm1CTSTtJ3S4iq9UPDgme1aGYXuPpgbvIe7Veu
7Kiob+cnH3uNFsukZS9LJIeUsoTTgpnupI42MJXJaVyTHDKcSx+iT4E5r44QQ420
6IdYAI/0gcw3qyJSK63yc/xXxkc9/b+TzqYKYk3nFEy7PJoYlph5xwL7zPh/+W9l
2sb8J+6+VoGSAkMoYW+Xq0WhTjAM6SWGDfwrecW29p8kMLRwGQ7/8wRoe6edzIOm
FCOWFpQ+ZqWnuSYM9ES/3e3QJRmq7eS0GvyBclJhpEk05SF32XSSubW+l5IMh9+H
INYa9Dp1vOQ++ODHp0I+P41z1tog7VQiM3xQo+Oi1wwZnAcIyaCDApdFUnMHXGCX
VJ9thDXeS7VHXFqjq+3KMYtsam4p7wQ4uJjGs1rAt/POaAguaGe3bYAiu4z95tIQ
dSWcT8vZEPvaYQ/lmCADBR3xuMeAOUCWu0nmIZ0Zjsq4uOT0JjelcuZofVdxalJG
ujX2T7fQpnoVQjRdy3piFjw3Iq+wTVbVLgXXtsl5kDdlgjEkDMy8Xlh3Lu+f4N2v
ByJ9aitNEYL29GFhNSVC3hRXzVsS5atWSibSwUjCsHG1GgTGnvLhL5Ey2hcYNNrv
Jf/4HvnkLtJW9vn2jRse0xq2V4r0VujzDTSGyqC1saF+WaCvK2cqPecNxAwTFwdg
HH2srNUS5lSjeqpMweSbgoB7tj4OBNmbiBKPd4KL83pT72Ko3EhrSI3PEUXeLQ34
8ZL9NehSMj2z8tYj4LGCFMsWbc3ZTFG8s/FRLHT2eC36Q1neim1nc/+0vfZhyjC8
JIbEYtRQxzfKtocmKtlgyTnPfQzQl1E1LpLkvWRbrs00/52omZTuqjHk4ONvmogi
GzHnM7iXM8Fn0igv0oX861obvDliVEMIZb7atucfI2DS52zcsXih5fTBjjGfCTiG
J2vRfBfLGceDZp9ds7RvrbnGqQ763L6/ZwhJLtOlQs/rbagcuG2UCILizQGW5DdD
4CuCL8v8UAjejk3HQB4Mzn29XVEiEDSX64HDBDC4Dbd1CGiLY5R51UdlkAm4ENta
mv6yKCRfATcKIretlz+NdspwjRBC+GOcBLbUjSSD/joQAnzF5Oz7aY0bKt61f2kS
cRpTHmPVK4o8ZvptIMekfY9QgnVdlJsEvW0w5vxvW5sZBph7IxbHa0A1CP+TbBQD
tSZXTV6Qz1dEQ7Gt2SkZKA3waxOr3OjdqrT2OsPtnMuDps0x14x7JTHxXFwDowBR
H5Y0AoTA2WV3ORxmHKREpbZxqxM/paOAomNAN/Pr1f08LFDxRjiFq8yljlCp1lAo
gjOSzlPgMf1azA+jZ9oAvPphrYoYiSJuwqlWKWUxr5EyobL11lAPlC3+C+ZS0uFB
l2zQyDnOyuRol/SeeNvJ3S53yocyS3P36Vg5adpDA77Yh2PqpebEXd7+cKosAMGS
ZU0JuIfLCyFGVROfHnW+Z7tYktt+tXzITJH7qrleJElaR4nmWTvxOvafhJqvSSIJ
eFPPN0bTCD6/PQ0i8bvYyZtarQ4mZxm8KSlebnela1gAutXIj7m25YjdOUUShHHk
5EtjMBQpTr9hMFfWZXev6v95V980aBMY3/rgUQpoY8CLGoK8dn1VQa3TXnddQZ1R
KMWUdWYMySJXjr5rAd8jk3bPTEu7xTug8evray4GalRnLsUIt3lhoNSs+IRsjdME
O7OPCYSBfpkMJKju7jrfGw==
`protect END_PROTECTED
