`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1u5ZjAlPxuXEB0BxZIuT/YNElnZmqtuGiDd2TaLkQvZ2nARu+Mp01+Y0FTxt6ws1
/48lg3LZw5PHjSaLhOJoMOltMnhMvtEHd7ecrAEdJ+VpjfIfhRggdWeQ5rpNf98q
mWql7c9zmNecAd9Blvl7vknAWx7ADe3rX7pgqtOKefYkBPMyqAMTS35n4xDe+u8O
cwu2jhIveHrHfqAtgEKNzDsUJhK/GSNgozQYXn/4gXfcKKFDIH0mLFY/kDsN+w+L
4h2Skvb+XeWu9cdZvdgktFwtW0UbFTcTniFJ4XYgtPsKrznYIIUqJ6Ys807P6YDS
1GaWNFtcvCR+3RjfN2pW5JDNDUeMDTYQTdoo01iAcoCMhwO6bJSNQdhO2b/3hL58
rJkEHEqsDmmFEEoyBdRw5Q3wk9DDKmJqkLCjVIT6E9eW08r8X32otFpqzPoGNbLh
JOsH5wzOfmvsjMdGN4SLb0g7qoKA6XBxf0edMycbR54JJdxj/Ohyq4dg8oT29fFL
ipJGA3soUrQ5M3URzMvxUrgeSdv1iN0crn/+0/XcZAbs6b0d8S6nBUn/cjFJeB3Y
Wo1OrTiK58BL3co9kft1ndIg55NyDVInhNCj7n2Nzp03FpjGqylFYU9FXSWMqejO
2qQe9YR8bRPBibeSRcpEafZO6COL6yDOjw303hFrdVJZzPYK3jPhAFo5FRTUQw23
fZGTSVX5r2py41cFmdmzmh5f74P6MDn0oQ/9x44Ty2GzRLo1w5ghQf7/G6pOP7vJ
oYpM9HbMil7LtjDJLKgJ+cgrbzRnS2QTm+iRLbrnzAv8BKZVl+igCRVtu6RaVs3T
Kak2TqGXMt0Ih3IUcZjNlxwxxfeXyoZykRTSixmgrNQztjM5ec0A71mc61UGkNcC
gWMMmRUXnTLfxY0Hg57qGaciOWSnrJhajnhHwJXaX0F0VA8XVL7SJnnEQlBgdH0q
JVTrJnn4T8z7nnYXSQUU+1fhSfc9VktCgx+ug4bd4adQlPDYpjAQ+5vWQ1tClkdU
BFqsiNoBkqx4RZSngT8L+PWj7GZKC3y5bzvtTX3tiQbFMC4T/NY2x4TBtIxEPpgK
lZXc/e55VGMeip9VTpqwwobGvlhUU0j4Rpli9Jm27Yq3slFc00hyN99VJGKgu6r5
INvjbpKGHNDNKgavB9kW3XDGqQZTjhqjTnooQp7pODaJ06r9To5i3OP6r09KAgZk
1vD4QAUKmLmG3dEruiT4WO0gk+wL8exbLQc1nbSj364uEgnmo3lWsuNJfoYdgBpO
HJbk2JILogisamXd8T18+nrIPhK583yz7XbpmGzFx23ZXdige5XL6AjoloyGTKdF
r5I71RSj9jBlIHKbXMc48zvvi4fsypTadyCGoMkUUtuECbMH1WjErRPjJ02uKkeD
IEuOkDHEQfx7w4SKpUkwfd5kitrUfQElQmiXAroHdsQ43C3IBPDFuHR/U0lvvDyh
uYvzFYQZNZR4rNQluDpCN37LlG0fGyHqsW1OBUXbzIGrI/cXOgp/zACa2lcVjLdT
VUnTO6JCv8ZtzEw3Ddv/ZMqS4YIvICks8NjjaL9WqavlDQWp96WkHbi3UrElmPeE
ZYOpYZbllMZQIlnPnJCmWqgtNRal8XmzlTP5J0hICh9L39XWYmM8ThBFMjdK9uRY
Ip0OZJDxdFqpotXxqwyy/m6gwFdvzdIW9fz6yyOseO0LEcWtjdguL8JMhJ71/zNX
ZqtmTPoMEOIu0pzpHqx0jiMOL/BNztTehfEor+I8rb//Zy9ALhGN5B6wtwRTxsPe
hID6o5LaDBMNDd5TlgHzpOV+XbDfY94DC+HCim6o+KEscBCau4geKbQCsJ+SAxQ/
ArrQfHMEMdgVK+mSXzUkwXzbF5ViA2jD45KiaE2DvO2Jup7bVK3IKWQmZ+QGwgZB
Q6qdMQGZULYRbzV9RCuMSmqZsd2PHGkRGd71uSvpQWleVb/gzVRx5CgOZOvb6UMK
QhG0wmmH7WMe49EW0pEEC9VuuhS5LRggASDiNOtyur09dzg52lgU7v43e9GWo+hT
Ba8fsBhmdu7sxtW5FlTwZ2Yr/mwBVE3JI+qrF/eaHjIwBGWmQkIWt4AdFDB6jNBV
fyfSf41Z0BpSvSJouIC5SXL/QC3P/6ArG/uzNEapTr3hzDqZfuKG/MYvlGBFgKmR
vj9Ji3whONAQDcxWf3WDr2XUHO9HNmJFTAOch9XhWUmDa5MYhgGRHqcLf9uok6a5
4E7liAich+Evmm0FjhomxAuqJroeHWDDW/FT/CfPP4JMljInV0HS+l4yIaShkc2Q
3z0UqC1Sa8lr5VnGbilNVF6sBmME/yre6kqamkSCEre66e6VrZW/mX+ePWx+n+Iv
sQLq+sacs9YgKOMVwJ2UqmFam1WvmEwylKC0lAm6T/LN5pWw9CFlBXv1NMkQG/lE
4jzEuyUGyMfMlB8hpcWtUwai1mugJ8oPXMEyTkBKpmHaBLVptN+EzyT7q//wrU6k
hzCNcXJAPweujM05MLd3PojMzy4OLmFhmJoBw2EBkbIFDdwjXuL7qxAaIu/KgS7D
m2JPB8RzncsS73tbid/En7edQ6O4tNrIx4hrndkhRYbTLW670moOultLY7EERj/s
ZelDGDdRdPYZv81PjmOhiXYQTbzkPrpaxPkhbdrkVSjlP5Z7twxvc90X5iLexqkW
jNOi0/EoOxCEAnz0UzB4hoA3u5/Wn9mU5nIEvuMkTpQn2MVxOUU6WcLEZo5SgwRF
wQljpWWENAJYl5AzHD6bMTfye3Qe/HTvz45oOH8e1FXSFlFOxJMXLipsWrTvQL+c
xGzR/u9XX41mt5i9t2L1F0dS8r9q5qEzMn3igCf7MuJaDutLoDwksqB4AMs8EBYS
dQwcizKLCFNfYf57fKAQywVodOSL0QHKmqNJBV2pUzrkpOJ5lU3VF5FWwj79k3dP
d/BpSedKfg5NjkM98+eiY1sOtwD+Hnaa4mI79/yK8n69mvwB7ad9KXFwfTZQEICV
uZkDf4BLaegRnXut8vLNk972FRjhHFwcZFglvOTYyT2FjLko7afi+1szq8TPj8Qx
/HGDQvMSQvrOF7ioKLp5x9unOboxmXwVAfLHGD+/dNXcocM+elG97xpyO0ZHBurH
zlYBZ2a1F/xtTm4CocUFQy9KutNiSax8dXbDS+DDbC5+TdG0iZh00MxN4kkPscYN
TF9u0jGRltXNirzfGeSCCw4d0hsKmcm2utLHrl5INJWxhpfJ7hveVsVTHYkfvkM2
qZztsJsC/LZeQ/97U276mQZyDstL183uzLCapikpqCknZmgnI58AYLe2Q7t5X6mO
THjKi00bdrdmjUza2EF6aXzVMtSTShrhV97+7sZNAOaP1mPWKiFHbNFjjkmZUXAr
pD7EVVU68GHnTI+zhvTdHwPKFet0ZWD9hznMIIAkZPCByzSz6e7f9hs5jRY/JRa1
Z+IpCtfFqGOR+Rr2a15tPC+WwMYU9mLUnan5tvF6/V8mRyoW2QxVg9fJKrpT8bbM
T85q58/MqsBpfs8+bkUnxNA7XQIm4WyxenGzZoKeKq63F9ssGJJbUTtbLPtPxqmb
QTshesNt92H9Y9GrvhJr6hQzZ77IoODbiAtPI6nLGxqsT+WHH+RfIibpDIEZ24D1
5lbYr95XjE+XS1eZZBFBM6wLhzXq/LCzztWwOFErbm4sXCpVw977LBoBdOo01z89
+wa8uO+yGBrd81+qanNNMOfdymM04/5gun3ij/ZqIJvBg+E/5OyfYVvOnnBxR2mI
/0uoeN33q475UJ546RZiMnLbXPTT/xrijpyYJ+NO7t4SoAI7/Xh/7+uTbHFqNIm/
ZhiDc+1UPkjYyHuH6jFmg1kNB8cPtq8exKBfTBD6fe98GpKVzuzmSCy4mP23Wy21
LivKrUJFYogzWivlbXJoGgFQVc3KpmOw/ZI/iZf/4vU4NeeO7qqVXiFUnA6f7scu
nst4ldj8On2xJYM+jrbykVckCn2Znzz1Nx2KyO2uyod9sdKqkUhwTHNs+DvvLdgh
5luXY845PRY88HpWWqzCNZPfE9ZOImRlbNx1UB26BlMJRxsz2fR9iBqy1aiwPAUp
KXxxQt/PloA+iwsk+6YQtzzcDY4tzqp2Xt2gipf8G1foOHtwEEIck69sObeheLlD
qlGhn77UNJibYClmEIq4DlKnR6lctSngDO+YTOrUOKFnUcvcZSMP4xTr75gnDksu
r+xUG2vuEexFOgbYvmuYk66Ec8ui9uykL9j0Q3VXgp5/DyXXLFWKE/Y0thgssQbS
TP/sgxtMeXgYeUeEb43387POwtnSZkVc+a9mdJIMQAv0VqKDD7b2DWzmo5c6HHgw
oeHR/wHsi4DPA6H/TUOryFlNm2XZ2psl9tbqk6Ij3PSVdWYbScREjvYR8dJ+iL6g
i3xKTIL73uLG7xHWrzm1tMYJGgomZhdYv5aBKUzKEjUzYsMB42LB2zw0/E/rd7Ds
smzDUdYQXSUr5pQCKTGkjstzGDVfIKT5Or/2QpKExNz+IHuZe1yeZugYHnfbp3RZ
hpT+q3gh0acUADr2xGwa5/8AIDcXmLqXOyCQ0UmRsouSaJfkFV/fw+b+HzbmJhAL
n6tx3T/hwpKPS3bDkfaW7bD/NHp0DyJFFHhK/mkabRKL+uakU8qSmn66wx1u0vcW
+Q1B3EpQosWu6HCiLRgMZN1mxWTExIakdhWZGBhF17KTnW4kLO1jAeVmF427CuT/
dUg/sKYlrZrisy5GFNiBMPw6FoDpOvCaZDWjTRtt96yiV9nmYXq0D1dTu46Ch9um
CKfQ715FZAnqzytpMIlGpAMnRdq5LSG4z97jImeLlEiVExmjrXoZ8NjpTwDV+qc9
apfbRlM++Sg9TXrdGj0sq5RsbMqblyBWaAkgaRkcK4tPu6vwIRyUj9vYRMbfrS1H
7uMniZmzVdXVC8fR9QCyJKW3edSVqfcvWE+t0S6juKHdrSsRZRz4KanOUFd5X4nF
jV/2o5uHXYaegwJaowMeMew+Fi8J0YMUXyg6HaPwm9mgJmOVT+QyN8aNbTp1Qfg/
HDHlKM1bxMUiBhbaM8G2N/sYPO7Y55i73fAse85Go6MmL/zWv0FZ11GRaR/AbPUT
2qsfEzD/GhOzNFZ1sIc6FyZ+fdY5f6EtUmW6S/M/1kQHjdW/7gEMGBM2XBgaWEt0
S+g+UcF4M/EgfppplXsckl57cX7PdwoWZCf8Cou+ns3U1KPUUNpiQFAnOU05t6YI
5m5pwJl/TIzaM/0jy6VyFVbCDEmDZewwgvfpa+On89aKD3E/bVJ4xxOzjXw3JEO1
i8Cm0GHUBE0tQUOD3CklziaT3nxAZ6T//dzVVFXA4cfSeNT4nnoXxu6Cxdv8ZEB6
PF02e+0t8wV2sixk5opHyJ6ySwjc/rw16qsDHZSnm+5RB4zlApiRtAib8BuzOe3b
hEG7UA9+cPYkMXVDTKmjxokRdERE2kX9s6gge7TylxBROVZbjJiTMnMjNR5SZeYf
ShUcyVhuta7xttsWtYA4XS58IonkWhm61qXm1WG7TBIovvD3A3RGTDgTQWUiOMqd
tHRRu47VYg/2lC9Lnvuey4gT5QmLnFPi0sMLcsUVpYwNdXT+z8e7rPmTSmH487ym
bUxgxMFH26CaC2lflBr7F1e88Ht4CTQx9GM6aV3XGFJpEPS80kDYn2IjE37kPfRM
xI4RyFZaQFK4OmEaZHlFQRW0OMXnU3aqrhjE4Q9kiK1CWvGbODt7EbhEP89yukkR
`protect END_PROTECTED
