`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bcStORvXwt9f9sbVa5nhSllv3EgEzYcy8ncM6+cCnn1ojKtGnfLSsr7BI/viCBWH
n8p1VPJNqdRc0RRrkQ27lmLcKYP7IOX2D31uunbwnH61tlQ2MnNtlmrQ60nJGhQT
J/w56V8B4Lt6vabpkNxO52euFwvkyeknlN8vui2x+yPr0cryhAN+enur9FiQpV+P
lDCZOlB2ujKVuOP1dIR8gn8Ue8zY8DNyIStQzPlzW5ifvZUJ7Gqw3at4IwJo5oik
SxeKAQo7b9ZLHZR6UMQ75WJ7Ypj/XHMOxemQfpXEwApe68nB2CAyS+fkoJY912oG
idnMN1RSztGgJ8q8UV1Q1ivNLbqgLargxRx7kB9sOc5kHS+5803xwpb96K8KBcKb
TlsHnYIfUdeqfjsP0KUmkegdj0BYtkfinqsYaO1qk3bsgZ5gkPFX+9bHXo3StDhX
MQ50UhOBFxlYvIxgKBV1zkzUyA8YQ9u5aa9t636nGErJbCCZrZ5IL420Y/f7LN46
0SX5X7iY74L2Od/nFPaeXXUcwv8imdSmAZEXluhS38fBDz8r2fa3tlLj0WQK1tAQ
VUkXQQPrGAP3d98KFMKmvwAh8fVen1evt0QL6CbppkZxlOvNbkYsbtKYprOWxPvi
VfCXXtQPclYSfLUjW5ZbF83LoheykESmG7kPMpqij+mviAkvglJa5X7C/w+T/PF3
uAIx32hkbAz37++l5IJCOj6aFtHBWc0lY9PB5ku3g+kvhtcVVQGB5/BgnQ5KcNfI
zx4OKI8MwZlq8ikv9jvBxUJ2xEBdsF22rTvCI+Jq+nbwIAJvp3/T5qFCDTPwmagt
ZTDtmBMgyfPQg/kHOUbp6aQ0GwpB2qw1Ok0I1RZAciAZ1UfivmFLAXH31V1W8xlP
fPdqWbDSsorb+eZLVcmdsII9MUgOV4LVhUigJSuCq023hIV5mQAfDcJkwzBHELNK
6914jVMmZV2WmWuy+tdn2bpdJcvXv2T1gw4Yk8SSwoKtWXFYJ+w/ppXnjeN1/iw1
9xEfVCnnGePNqcbuIfzw8MZeUejxdXWD5xoKF7wY8HSpOg+zIvRgJlyNhkG61xnN
/pgGpiNINnInJrXvMTnJeFBnKV5IG5PSbufiXDLoPnxPVFVZbM8tX9or6QA8yI+N
xhK7WIAO6rzI3L+pyz7ylfyudmA7Ag3sZGvuiA3lLwA3JtXidGzwFdG3B74EY9w+
9T6ZBhAmEUzIQuKXuqLnR+jCqx8grwoct154pk5FEsWOSx6AOcx917jgbzSKp7Q7
QmY5ETukyNOuj1osmhgmPUQyMQlvWkwgni4GoIA273dTjM15fh4UgwFUfLYLLdQa
YsccXoVeiQIH/OPxIlJ88dceZnYGFFQqDugFw47zqIlfOR7F9bQCa4ZdkKBab4F7
eV9+a/C+0XfsHETUWqzI+voDkxiXOSTuYfnvw6m37oKJvvINVDrlGeuMC+bebaF8
t56pyTeujdd3+z+O3cEdM56Hq8Ow4ICqtLh0RstmXzzG8+tITtlKUO1uUkxmqSXz
HY2cKZar8m1M7+V2euAtSxdELJRcj5hcxbXPYLqP+8WzGMJGUjXYAo84yl/wqXkm
6rN6hZnrfMxIQ57RUH6evXagCg8IGjL6AZTe4btmfMyHtgRvewPESINJ+BN4IbY4
zoJANikWZoFaICEOVE/dFt1VU8W7sq1/hjr76SctvY1p2vQ4shwa3QnEdX//FR5o
+h1VHPESzZPWrZyJUwnhK7ItMYURk1elk8qLp1E3b4u0hAsMf/QWjU1wOUophXVA
G+wgiX656zAxZR+NtrLwXX94B6i7AL+oBvgoIWa5P1DBaJCeey0eVFMe5oo9PB/X
5eiJ6miWTVQeNnrgcnZRT/JFHLXfpV3Q6hSUgjdrOBBK7Nt6Sh8+w/GjUAdqzyRO
bA38faPWGUlvJUpKXvnAQCACblS9+gOT+G492MeLF+zotROzwL8rCTnzH7vPgFyL
7b5+aKHSMPh6V+gHZVdlwgjsDHiM9rVjz95nbbH+YAmiCQcIIKH91sRD1Pirl68a
/meUpBlfrzNuvNBGnPx/xeACtri8tBhNDiMFDt07HHMcK8l7wYcGXVcCOcKmoXdJ
4y6GnV+fs5DEjI+n4kGDoGXSJvdlLB8z2JJpSVKafgwdgIIfaRhPpwlQQvZVBWha
Ym+j5W2rSrK+WN8bBXWReBT8STx+QnarMnXUbzLaOdoBszcIxmH6r3/M8iUumfPE
iI1djKmdhA3/0PhEbPN29zs8m8G0D2bLofoU/bYhPUM96tIgZXDJ5VBV4zZ3RR0T
vF41srA2qfwssv9xjn2D9HxuztXeOHuJahbX1u6+V1VB7rvTxKZXWoZaJ8UecWP2
qtgcX1i2ZPc+1jXmpAMyfpy5OXQCNXJveHQlLeZXXDXO1+JA1KK90LwpZyXt2CvM
Jn44zTEzlU5jJ91kSV8EYKb2Bc9V6jQYyHg3KuhK1g1Xc8a2UdklE61mMsnXwf6d
0z3yje49LV3OcUPTqoZLf5xL4TMyAPvyzljCoDQMP0pHgRudkSY8yN+xrO9JD0mT
Su4vjCWqhxreE8uOdM7JdvK2rDO3/U7ajW1FfKdqDsKbj00jVbL3nCGaaDBxSGVX
cfjgb1MQ/pH7zq+g77wUMUvKLHq0Uzd+/vTT/G9T5ufpeRvWF6PaxhfVtnj1V+Aw
vNj7uyRKMgtlGeUqPe70hL9qNKGSaLSO1IRpa1wEaQO6qK+k20qBumc+Vw9PrDft
mMkSedpPf47HjnxP6wSOuidN4di4AL/xGAFiE1zMcqG3Wgyc4T5EgBrkGHrCWwPV
WMDiLk1buziefMyQNStzvuX1s8OaRc9a9rMv57LHH/l99RYxgeq5MdRvspzMrpMT
vL3DIn4Omne4z7l23ZtPWac9/S/Nwth3o3A58Edf070K2/mJ8qzzmXNXOiN3MLep
KN9LsQaZOV7M80u2A7XmFoh7A2iO8ZGu5pwXUbfrIMoDf4x7MK10winwzaVPk+Ss
tP95hgjmVfdAkW9jgNZvHexB4Ze7n1Ixx6rTrLadlSeRylLMZgAENasGpu5DLZM5
n8VXJ9RMNeH8kz7jIKA9f8Db1PtmDU2YOAae2vHACSalX9/ejnqdLl2PT2o+plCd
0B4N6wlwPCe+vS1SQ3omsd6sykVoZbChx68q88DnxwoSIf8d2yRjoTqt/bXRcHka
kBrPuIsBfBJ8EZyiAHdOtkNTcMBcJHZ5mlND5kJUhfBVwoHnz+zD56b34QrA8I/X
`protect END_PROTECTED
