`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7DkN7za6Y2uoK4J4kc/7ZWCr5P6FcV29Nh3JKCME+oHbmOSDGPu2AM3TiaCgeIy/
bpW/dIz6QAdySWk7pMxgzuTh7ICi5IpBIJPaGvNteG3h8jbfTVUIRnEseqXKFx13
u74EKDDh0An9Y+QYKWHsYuWmJJNUSGSiG2AOyXJgBDwkCd92VM7kzZWS7nWBa6GL
nmWxSD33PMsz9WQstt+78j7/o+SR9TQ2MLMxPIe+K5DjdFeq7thF/aEsVKkcb6mG
xVlQPODz5pUksoA0aF1PqJkTUJ7fOLvBJlVIYVJDuiYOdXyTeJE4sJJ/7rHAQDCM
HKs2wvAVRcE/K5T9ck5IbYRS1YNA8uvXLcj/a4NDyVZGrOcimY8elPhR6K+JlgFr
6oLlzHSJdd0X2pmVbA8cAqJe2j+PCRvhGtkPTgCUemHg8Ic3yQ/NnqKkQ2CXFE8p
bIzBxrlj8r4YMRepYFFxrz9tVYWH2868KzDl7ijQyQvZ8/JqY9yynnIv+PZ5szm+
ltVTb09xBoetjHuSzG2zwaXzc+ayaZckBf/z8ut8UHJoQN6CVNCpOldWYP6MrasC
KkB/NSfcudyC8DSprw7n073Y72lpyZZfVAJ76gdOHHObj7izwEX203lIPbyoE5Ld
yOFvIn+3Qa5ZASYNCd7GkQ/fSfmEw9r1iNz7TYXZg2SnDAXg8QMgR3as8N7O7ayH
gp//CMd3ckTkRGdLhPxVp+4vaL2Gfa69yCnJhWaFDwTzDi6RRkZfCZK61YOYEHi1
GwAxw5V1o1ivi7W6uuzeo1/2TwsqrJQRyzKLd/Ufy87s2qfqssPbJVV513ZPSCi4
vIA4caAhK/pCIUokiT1BXOPFaUOhsBqpoLtbdAuCBTA6flllNakaPMFmuXv/eBio
0oe/uVBLGHkSRr19aeXW0FEx9PbxLfPhzB5dbVhJt4ebfqesJU1XHV9hFYve91M8
E11x29PRs+QQ5yt4dC0niO/vHH7Vpqg4XMGFqxAZK2U5ILC5K9PaT1hK7Yrgs1sj
vAlIO6e8oW04PYxL1pFCWN6pfCnK5stvNKXcNjyOamTEt4wElIS4KHuz8syT5n+5
PI01hYUX2OKDK7Syfcg/UxyCHJoN8h5g7aHJfj1EfjZL5INbNIurcye3JMd+23qL
RbPhxiVlq7zaKmffwjapUGPKAOA8+GtPoTTbz8MeZ0PwtAYGEHrmLD4ivLG/PJAE
1Rx/9q/jidPJtuD495dnptYl6DjiDiHh+bGdNkcpT1ux0UZR4VYO1OaWYYuqxqZT
wsKoPP7CJQi6IOVYyDZ+g9Ys4aWBl+F4DV5hfu+iOqtT2G2UJn371FDbG7fEImS2
QEKtB9mcz8G1XH3ByfBXjxCee/TRyBZv0cJLr7iwmFnPntlRTeVOTJX3VzBCSmKw
IC8HIY15MFdjAquVQ95VZO1GXJoJSLz3CdqCsyBZbQntMJgOWyQbgTR73hUrX+ke
NUs8l0NUF/n+M60/RDCC0LhQYEOOMiYRowlh+s8f7Hige/uBKZlSU1nxGT+kNhzK
k9Wo9WN6z//LkUZGafI3z5fuzlhJ5AwCjsv7hXCRLDyg3kDtQshAxGsenlHhLzEU
KsnsjryG1+t63+/wpdaWE/msp3krXqg4QquhdXQMqwReMgwp1ztgpo1l4NcJ3CPG
3F9wnMVSuBkgEWavU+d9Caf7bRssuxkjXeuPrQ1PhCh2QOvx1dJLhB6MYWGc/0f0
CbonVNtOtv7XtfatdsTeZ5Bark2BY7k/oTzjdNrhWnO/n1Gv2Jvl02Ksl5JxvsWQ
B28loShSPJZqSXNfVXdyo+vQP2ZQJCAekHduZQPlPsnS6HVy3sl4PykUPci6rrQq
vnqh631sMaHDXeMwTAt44KxSM/bdCB7QlrqyBmnkSY358vtMxhzV8qfP3+eb1nol
Fz+y64AQafQOcfpM5Yy15A7z5brbBmby+I9m/kfPkNNVCIDc31ZVch/Fm7kBKIhb
7rWCIbANjJH1C3hUdB6zU3dfIrS8/lGA5pUgA5diklo7iSwSGsPdS4pUrLWU71pt
UkLXguj6zGqOjFgN75/DtdfL8a5y4InR8dCNV83MAHUyMrHAHWiCUJrkGFU8hkP2
8dR7z6RQ8RxeARNrYtX0N9NerTBEOV1etEutvxsjhgMU5nPxVo2j/siCGCZtc7bP
eW1iYM+xmpgPA+ctupvuwV+hb/GKE5gaSzmzE7f/P67zVXRQAfM/Zg86ti+Zlm9S
AmDhSTQ0KIiZGKy8kknZ/mrCMBFjolZ4KnOTBTy/RDhIwMOhFlWDolrqD98HD/tA
R3a8IyOSdOtp4Wx1z1yHCPjRQn8hGpF1E1IMqEL7ld8R9rnUgTOA9ek6ppIH9E8n
HDQNbs8Znm5288rg5IiQb3+va0yVq5meibapaovmyaHJtL0vxBqHD29DmzB8VGZf
b1DCyr/+NBm0yFCKpKQejKsEtMu05MUZ4HymiG1JjIvKP/fYShipaOANh+pTSrZK
Wq93AJ2gb3IJVw7EezfAqdSlZYD+kpATPAEqFBupWvu0WRocKysKgcbbp4vFmMB9
qdatZgoNaG2JwFg1xBppSdSrb3l0SkRdTWJ7f+RfAn6TqTwHdvRR2PwWAdTczygk
GCqeC3ShCE4Yhnojfjkiz3hSQYFzBakA2ZIrgqFcsvmDQQqxFGffBX5eVqt1KiUm
MjyIEh+u7fQP9mc3lmFLAJSaRE66mKME9HigAEAr2tSE4TUVJ5rO7VR3yxKMZmTB
U2gdFVfSxgJCDmGsiuCKUw==
`protect END_PROTECTED
