`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clKWRPHG31Enzqv7635KWCeurZK5i0Rd3fEfyXRU60Ewj4Y4gifxIACYGreDZZCT
E977ABJ0yP5w5gKDN5AAc99Ato99JdBcyERy/KU6I3dFPlHN3cuqZYUl7IwkoXj7
rS+x/Wa7uEyI/F/W3joDLDllAqGIR4+z7rdANIsLcY1cXMiK6aUSoD3uDtwPL5RR
L3HDSG0jYju3+AyPf/D5zYe1SP3hchhKAyklS8YUB1xAhzocx23zBSLCxx8ouWie
uVO4TnHopzbtBPvJDQJU8qg8P/IFo4U9TIf6Shr6KHpSAPEHEot8iOdDbgR+B2Xo
itvN9ZZ4RI1xfEYWX2O3vZ4dIa+ZhVsJ3fY2HJ1tbFQcfvdNix6Szd1j+iOBuWMt
jjppN2CGVku2hfKiCqNsSnyF/iJcX5HkY7JUewg/ipRliCak7M/vAd3SKs9mCNZC
zQS1dhi/WKRIi0Rcs5dsc7oNnw4O9c0pnjnWMcr/GKHmDdAPPjiAswNSaQL5jI8X
oPL9rZ82D+r04KsZ1giaSmyC4Dc6uGmUs4nMYZLQrApOVe2YtRsp4lpObrSKOKO5
VfBjqMaHHeI2O6sbbh8XE6CAWmhqWSRkxj76Ejz0RbvF2B7ooKWJp+lI2FxAuC2P
iS/lvLPJOyzXpEYVad6LC+UrR+9F0eB6b5anuxvsGDLwOBB5SixSmzbbeyaFlplU
EucKjbsKjVGx4gLiyALJ8J5/lKpk4S42bXbvyIArlp9D+2Q3Y4DHU+1SbKqRgeSo
SVlRJjMIOvBBpg89SezgfcDqbbqklzfzIH/K5HKBjf0P1nR11umKaQ9k8T3M+RUn
OoDnDA0SMz+myfl49kTcsxaK4y369VPhpFiVesXbHTD17Zf1ASuwEQydbwBxFOU8
cPxZA3DTW9ZTv1d70Pk3xO2izPBMXJg6gxN7aanUiR/FZYNN8SlQQOixcpMESg6Q
E537US3PFWG1R+BvVSJn/kZP+vdHbrHVytuoCHBBER9gqJ/bwoRAg0Av7UFNwQBG
No2KKGbkGHlJu9I5vpV2tAYu6cNb6OASOXKy+ELtCKViSYhpcQ0wFTLz1P8mZOn7
gkElWLlyEngle4i2XIEORmmh5/uPT6yu/AYOgyC5Csfek8NBvgbSS9AKioXjOffR
2EW7r1IF9t4bKm6193IaGmgIE9w0uiuw8vMSRGfHRL2DuxLymvl09mc+1zUaX+IS
oWoSjDyQZBtQ+znIZ6Y5AW78PJhh5B4Ki4U4vpCgbr6DzS3K50QC2B2jSzyEyQSn
H063sS0Pt5ZPd887blK9usAUWZAF+5POg7K0RULZSmix7eiidN/e5b+0Dtn/OPQI
vZ0s9CA5U4HTlzi/gzf5eTNNyP1HtDRAgY6RWUDJoE0bwBlOZj34D4Sta8huBEjZ
2cb2zauVvRQ80otkS4i+JrnAUP93SfXs7qpXjiRQKeMkT49ZDbfRHWiKCHycovg/
nqDJ3S28VrXMg+QtYCijeCXDhhqrCNDrhg38uyp/KJc=
`protect END_PROTECTED
