`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Z8LOQTOvGy4yujYLKKpxJCSm9bWSOwO56k+14Y0VGkZvcakPVphgfBvi3egiU9G
bNWt6KIpDZ/9ENdlEhgXhLgwHXfiyJrUs+jF2f7t+Rx0A6GWoySifeBElm0qV3Il
t3ZBkvEgDKvHp7EPEbTdE/vN5+XS/AyZCHXzYJNxvoCHKfZuVsx9kFVfZuUA3HKh
ecWqR7KSz2mJjsrk/M+5QEVgIBrMiD2qCeoEWxfMkkLKeE2oj6CanhxcZQSTAIw+
xKrEq6iM6wNtYbrlk6KYfOxXul2sc+kr9cOFjtZ6HE69GSSh1R88muEiPDorD875
cR70+ki7otdwd3eQY4OKurDns4OgpCOuGUoCy5gWuAj+GsCTpuXGmDAcWQIXfwkZ
JK1ijwqdS0MlS67YFFWBkSyBJcl5Wf7EQramyY9f6nV7GYPaGU4EZBSrX5WCYQIh
6CkvDkt6HRSj6ydq02FVTFulq1/fLjjE8F+G7iEog+OqyOqyNugfujSfU6oNYJZ8
w3ES2hkbcbVw56J8TY1G/E/4z9odJoBeInWQwRVKd6cZFJqEkcyUNS8Oul25L8io
f80R/wntJDEs6EPdH/tVD33EeMHqywm/1mYW1UBuM5ZJ0P2oMONE+XOwEGLJ+aIw
UWu51FiiJZ5J5rcJgFR1j32Myt5X9MrgDoF65tLJ24tP/NAlxWfPlR1jYs7vut8r
RTf4ADIP+1qSJQui/UbQoC5YCCUw3xfxP4EFjtqbs9k96jtkjg1Y+W21AHzYZ6LH
ZmqOyvPHxs27e/7LBPqJbFz1ZfoekGzdw83irIgFiwLVWkKmSvoRtzbsEWyetdSJ
BKxAwltu58Ba4d4QAPPLrEiYKZ8E1jwNFhSJBYsy+qA9iuYTKDHeHdZYK4Gayr7G
LcmjEds8Eit1e4M1DOw6fg==
`protect END_PROTECTED
