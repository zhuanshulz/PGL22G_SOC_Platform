`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o67z/TZ0+8Yhw1Lk+zpu3+q5DV3YorUq83mtg/a7ZRmfpixufX6j4IJ/TKotZMZy
tg5QhCdfkwJqaBVEjF81HmbjzGNu++de6dOgWGnBwwqNoPUwqIX4h4UxQAe8QPXU
7VsjIIAzaPnnaCO/djJDVLzGMEfvPJGWFoZz20ouHLWfg1Af+y2i5hZDc9srNy1A
HbMVAlOTiFNVpAfqIT5bF6rMchjSShRRN1g00vnzN2OpeWbI/+uog/zEh5jsVJ8E
ykg3JxQ76TFx7gD6SIKTYk1uDajoFIGIKyVF8ACgt8YXmUrHTUZHn3Nd9k4L0DOC
IhYwTVDY34hrmWlbzpZP9NRURMYsxnm6A7SsQsBctVHTgj44ATsQPguMMBvYa3+5
x5vF8pTOfv0r+rABBs5AvVjA6fxrSMlHopFvCi7CXn4ZpY4k5dX/fdWtK5vc2Pn9
fMDeDRZO3488xCsRl/TlxktwcgFNvRN4jg4RbKmysBheOHNTwCLkk3rGCWujJFZf
qvv3J+39xio+e9gTbJrlOE5hnp8vH44I1WMuDDTzI5MGwpBZF1M4ZnrovZawdxDR
4oj1fuMp0ao8NO1Y/ySLHzJwikM9hTxOYvp+Hyazituf6+NZ9VbkiS8/MSDUU9gv
Fd405WIMAvgLI6dmrKm+S9YTsO18uicwquQAIV68lXyB/UV/wE60JgG6TAXZgBfL
U81kiVhl67fbyI4Sm87TGhQ8D0+5w+IbEfoQSv8RW/dIbzXz8LkytSITQ8jj+IU8
vmlAOyu7A/6uewsiuPIZmN14X/ilsHCrzudoZvoexgIiO3JZ17+k/C0kjyD9AeJw
KarW41y3AAuaLjacntmdgJSD0mWWztzBGdYyDYS3iJuxtnPgmeJen2+1TygT/2Vt
XTwG29m3eOqB+wQIKT1anJ7KAo6reLF4M5FwHyIGswTfh5PBjrFZFtmBoS7gNAU5
sJzeg47z29FnU1kEmS0DtQPPg9FNt7gP1cfKK6Io9UQ8Nd1vp7FnzgrO35N1+xKo
3B2pzWNG+4TnUkD0Tulkor6UxDvxwXWiMyjCLIZ6bvstx5QCoiKpksny1anMYAyY
PcrmS3xxn0OR7dG1BvFNRVWNX47XNjHBu9tdrP1fwFOaNxC70e/qZR0osiTAmzON
lpJ7PE3d+IuUM/FSSno/2qHNon/aC95x7z3avgYaKV8KIHaLm7Cf96/9Vdu0squE
CtDOfSbo2k4EWEX7JHpOcnHggE1Q02+s9MuUKeZtep1STFInaSR9k307Z1Aa9ZBX
P0b+5NuUbp/tYRtHDaNooxd4jlh5JH2yVEDsNNrtbR59jExtLcxb0mnGgWLTH2sn
GBQtIiE7FY/XJzPsjagXCoEGJ80b/KpJT/9uQyyNaR39N/SIxiNMxfn5TaXEcEWF
fNuzn/hWbQsCYlC6ZftCb/wA7hRIeg18N2FSJZY/0iEAg+MlkVuVYfFCcXr4UeqS
zjQYj+zyJPEp1yw1vPjzSHRdMC2umBlWq3561pHIFk/bNJin/WDEDepvyjNK2hc9
F8fJ5SGW9i+qGbVZ+uIhjR1dq65/O0gm3DV5Ae2UdGemnqkbB1iJVwLXYb6Jd+Xu
izHxa+WjTBKHBT9Q+flazFOEaeLEHW6VI6TyOSgP+IXrTdPNZCq3tu4Eltx3VM8i
FTLfmTtxfsvb/CX7rQgRd1Kbn/3JsyTOGjKFIjP4LxoueTq58RTCONEqu35Irb1W
LfCm8wXOF/C0hicIBjhOhEnmiauDsXQ4u2RmTpRwXUIWTWK8QeWDVk+Vwv20TG0V
NJC2U+r1UAAt37l3hW4L0xVbQXYV5f8+Lg83ibrO4au6CPE6laLjoo1FTEZboSYM
VwyfwbPVGGEGa9hmZ/Hajr2PrnNkaL2yeiEGrzXvtDfIk68J8gS597IX0N3uMavX
O16cYmK0XkyTxqz+WOguP2ZLXJq4dEmAPnpWu3xqKZp2iQICDJp246GHeWhol8iy
fzFwufTZjOhYyfb2KtpuqWlevaW8Jwm3HodvFlJ7EeZmGcf+wvxJBS/7xnW+eA8T
7dYs2Bl9F2E1yOH+DOi+h59XAqyxtHCYoe4HAWsoFX/z8b9/aeaX2wGJZY/m9Oxv
5XPqWncSRPqbV8x887IOgJJXtG6mgNd1qI65rG4gu3rs0cyhq/j3SzTQi/pPi+uD
CB6I+feFBp1DFLaxqDTXcXC2DgkCqM3+kSXorc180aQBpI2W8jr2S0PmFU34Sqmg
AjGhcHC3CKkxq8ias8mGOieKp9t8akbhRwEvCo9WehOAJHftJZo7ERXBVa3jdK2e
H1Fworf5AM7/ixaLprT7an0lzl6tX/Xgvo+KP53EaU0B1OnW+q7/aHL9ODyX4AwV
pdNRRDfhXQjfYNn+Eq3OAM5oIAcpJLzgqk1hzMJ3vPUPv+RWfUNIiENbPfP68P57
IQTT37lL73rPQnReInScwC3rU8siOdnlqL+8NB5KPvZi+6LwwQ8Kywf3Ao3NmTE3
fsVEtMiw8hrejqTnMuWyHtBYoLTVtzM4+aMwQIIx2XJlouJKilCl2XYZC48z3ft2
+Ie9MLTrMvEeqow1SOFpjvDkNtM1ljy+SxoaEyyNLO2gfs3F3Es220+gcoQI6GlG
maOO/AWcyLQ0NBLb/x7DpMUfh0d1rGe7ZbvqGi7gPDtZGIelFr+BPxRkg2FO5gzO
ZVetOyNGt7HUxNL6JcUryvCPfg1/mk9pMlBl1S4Yric/FAH5P+Q22OlthZEyIcNt
tZY/oh44PI2ObUvM52PHTSM4+wJrVBIqyQyZzDUDZtvbO22DCzlZlT8/YB8Xvadm
eZWAQSM4YcLoSiOdK4yMsF/YItA6O5WhABQOroMeQyKLI9gWpkA7sinHMVCzZV/F
b176ZKkBwe/QlS3TsoC8PmW44g40hMHfGOzPTHx9Np1cTpOGMuk5Z+330W+sLBR6
CcrfdTQtvrJOwsPgA3baBPeE+onZS7uYnrYhZqDXF/0VoV4eaOGe9yDutl/tFJhF
JlIkpEdpGhxWfgkkgcNma+CxaZUV3Fw4xfPDbM6uibJWGnLEqHwwPfSNkJTb2G4y
nz1M74mj5BKnrCNG710pb3bvVxi9TL/F7mW1Au+8msM5lp8sVQU1QnbNQXS50bvf
WrwMHFZo18OvByQ36BlzObF5V/BHvymAseM9vA7KTijXwxDo520AuB07ohA/RzJO
NTd3NtOgL83Mk6m000Cvo8SOoKafJNiwYgFxDHiM/2MGizDc/92hA17rChRjxovx
g0eZEskETZH9JNm7pnRynRn5xwHuw+MMagEAaxliUfRsnnTyhmRdGB5Z2Cn5WlcL
1CAfpjqP0tZHP8TlScHYWR0l0ih39KQk2+y1iPbf5b/dXDIgTIDIrvF6d4+XNWMf
ng2FE+DRprVgtYAJqG4h9UzF4is4d4l1GRaQmZU8mEciF/iAQbmJX7ULS+yhxK66
gEjlaxOebjksyelNYWd0oUj72G5kJLSbUm5x9mhmCoyfx1T1RVxiCntNwXLLh8sb
+scQNmsaffblcexkDKH6MmzXelidbyTPdCNIvPbXefPRqS9m17YwgS08kSOUOwR2
kR0mCpv1RAr3/wB8E5IjNPWaPM1zAHGPrpRMUI0lX4fLiDDLD8bykZt6UOLB1gZS
Yq3nyFvODfDZi0ff77vNagDaILWwOyfxkTbHsPu8xUnGoNuLJEKTvdKAE95Hlcgx
7eTBmyc+0JaYgoQyvsvDphVBC7CJDPep3gid/Li9PMOiAW3xuGss8f6TpWpOeFjD
NSNVCVXfBRKeftvmYrUFBMME3TDHDCSdDcFSnv3hDjFvAUDZwBzqD9aRx7pBoWga
nNU5W59Da/M6kyW4HItrAZSvRnQLXbhSI2f04+IpIYTiP+xEzdY0z9c7vVhhrTwI
7qMbvsOS+gQnJaziW1ZgI7XhGwbXU2CE9zGjuo5on3J1j9609wxQnnZnAZE1BdDb
Vh/22UzlUXS4vNrrcKBF+SZV8MKD2H9jGGHasrewEyKUpnzCSt14Prq09VN80mCI
f5paJHwIlqSKUdliKp6XrpBX+la3fi0uidiZ8gYEUqd6YOSAAxFejWA/oYEdlB/n
GalgpXTcXYZFrusGV2cORCMFITkJwlEmoS6J93dHv20+3AT5Jj15PFj9mef87KJY
AFOZvomEXh7Is5sc7MaXB3xYZS4f/sGTBTCEX/jg6dESbRgryRSjjxnP5pF845UY
a5bcKKooK2+o4D7ltQM0EMcUP3g33oyPtqioCxnQRkoFvhvPY8NeWgU3XT1Swt9q
d72csmboydrQsyAejLi8PVE9S40+aAgnXFzEwjwEbhfIZ10v/LG4CloA5UJK3A0m
s3mYFHqsqt+p6wVBGO7xSbN2KR+3juw29MArCZx4F/+DqqPOHncXmDIuyhNl8lJB
1XPw6pM/xwG5ezXG0BIJF1OkK7rSsJEJ0Uf+a6aRWsWqRrzbQvjJfD4Yr7wD97Bh
Ng8FQnhgxiNomke06t5EeQ==
`protect END_PROTECTED
