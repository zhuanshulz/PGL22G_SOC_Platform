`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6cjxD1OHbYmwTLPu4Yg/4fpEGsjri6BN3VfuWQDx1jk9Ny15gijcE35fDRg/4NA
jZu9x+tg9RuUc/R8z3xQfXFOS/fEoXE/UX878V3NQ8OR/MGXYD/yhEaGJtUc6sFJ
jHhIomOvgu2GORYA+9nD08GYTVdOHT8+jWvfaOqa8pZJjydZIQ2JAg28aDoaxjay
2CkjrHCC6kJT+Kd+V3OyaXtFaf0p6M0E40QpnBjpWhXlQkeQM+Q2oEfHCL3VafTx
U2qh7p5lWA/5lbqQim6eTK5o4SBIANte3ijn1H5sa2fvOkL11JgRr4i0Kd+NJYfc
Re0+qs6QxId4dr+epZVWxX6X4IEzLmq1+V5MkdLMVTd91l/+nZm+q8krbM8GlEXJ
99flQLSsWoU6sgg/N67V6kWL52dqgGvBeS3hUk10ANFrmykAakMvBBChMwqY7Z9E
yQOyowjmf4sOXp5lr7fgsf451O8u60xL66jJULTIC9vFAdFuQP3ZnGCLjZXt/gyO
bF9dvoUbtNvN2xqikx4XHecejmF8UVozV6vU5SYIHM5g3CdlQIstsSf3D4q5Ncve
DHzMk30JD/fPy5YoLRJfq610aPkOy67GwvuJAWGPXlqlr1KVT4jcb5i+FefXEiyU
P41RBG/260y+GUzbz40Pi1zJ/gzCRfTgfBckjwVBRjzv0qoedqH4Q+V1s2kIzsdj
lhueFof2OUxplm+yI+X3zNpH+FN90rDp0XgWNxPqb/UoTd+RRDNjHdc/1H+mQGGx
YpKejLKVZlNDSQLrW5VussKhFLM4dqwPFNBUFc2f1edjXJD++2WWdWK/7A8zKGMk
+Fs0KITPBiK5+HMISBE0gMulPLezo0qsRypMiYW3Rv7Jq9e8K42XxS65+WFmPE8R
4cl15ca5NlC0OAI1UmIPqqltYzfjx2V58N4hYEmKQgXC3OSEnal6h2mHbfVp1zOF
IYx7eGdKBLq/dSWkfyE57MDmDNlyr0vGQL5Y36uNwH8rPy9qT5RP7LM3JY9V6VXe
`protect END_PROTECTED
