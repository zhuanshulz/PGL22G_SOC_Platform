`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k6kwv6N/a+CnE9y56Dt2q4V0rSG1NUy7MIiIy3hQQ2shioWAXwojnhJSXQg87QfB
2Uz1mPTumleaow2AzQS81L17UTQC2bEsRMBLQuvWL3A5A1PqUJmhs6l9i/OOs7cS
sqBZMRityuy9QfpppEc/d4KHWrhHVUd7DpW/qSH7rYTRUkgsK6mk0aXwXSGHajKH
W4/yePRw+oFDmXcZHnIOmVzDug74wHoG1rS78u4mOf58Whvfz2+95w8ccATkzn2B
QdztMJ6Ay0ZfPPW8xvmGNIdCXbhmSpE4UNaC47pPniueFIoxqmz5+7z4PgInooi/
jD3++tcp3Zm36TDnBpEBgdwZZnAg3UFNj/ry4dtXd/r6AfPm88/erm0j5H7CXj2s
XM2E7OIM3LHLP75d9aeq2Rw66vlLeySjWl1t2lx9k1rgpUrXNxShHfQr+8o+8w99
bx0iqW4m+XHzDdTBiZXMagXUlQM7WV+tdXl+K63ttPCNfPmSof+4TgQjzQvvL8FH
hC7rBbYv9GZrQuNn33zoXAvQFJtkdmoJASVQF95xF0ke0e0oUli+bxxlUDTx60Yu
yIBnJJa1LmIdI0es2lyqNHcbynJdHjI1lnEXmQrDdE0FzOii3EDhCOHm1xHiAv18
HepFoct+YoQDxABdjOpfL7wdxrmJ2J+xfDWfR5/3NJvlzDkqpmWpb91Y1xjulWmt
YrahzLUbajJ1oMr8wQpkU4oQuuv1dx7wXDq/fyMjIMu2KUvvO0nYBhqkUTREUGEV
qPuDDoIkI2FGZ1L1gFco9EzPdSDyzce5rUbiUM2r8urxjd90Ae0Sn5eCKU7X9l1r
dYDQY+58CAfbxeo4s0Ws4y9NneStZibgMYxLpYM+/m0i1KqgAeLtR7qfcZ0JqzrN
Up3UxfSgAaDYVRcb6H9pvjTsonDeL7UpxTIlMfp90Mu2ZwJy0IcCZKZ8ID2E5KbV
x7Ldy+iLVVv5f1ul3iQjVnnuvSP2lzy3Ohm0FKSp+AcYAejrutJCbXVhYnASeQai
moZrD77RhNnX4wIN0c3EIS361E0H8xHR9vviMzPYD7sXYcqapaJm2NoqMQ3Np8ep
u3PqH4pqtDr/fDWJ/Kd3roQzda36FQj8Id16eOW/K82qlLimQY0Ki8xK+T6XDN42
X4VOhzGAisGOdikxetA9QBEx0EOenMHS0uDRMQK0ojCtD4q+TCxKa6ikxjvitCv4
30dkyFkxRyg4MWkETpLE+jenPA1hyr4HmBoE24ibeCcomEke2sPoW2uGBVjRD8Z+
eBzZw5KLj5yxvc3ZGZWVYg978EqJYKSgDl7EhSWsk7lHdy5DWGTDIXp+WnneI0aC
7gmBpORnORRzvyhPpO8jJMK8ox024/GkDarVBmVR3lIpmB+f2/N9efHEA9KFrtrD
6QZi9iczc97/aln8aG8wdnKNvZ3I38tf1xwVxM+b2umi/BSkjhm6skp2WkmkSREv
lPVDAYci0FXeyl6t6zD6VfjLNdflj0T1V5AqvpOVTxr4Ku2T9jCIhgOQ44mb5ans
c7ztDSO0W2ynliRbfr5VRWFHw+O257Pqt1vrbHwoZQNt8sZnA1XJEgw/LF0K92ow
lQ0ddqgAkQB8r93vKTv17xRzZG49vP3FOUsB17b6DNetMe6KVkdEHGiw+X2l6jqu
7pkHgxIwlmB0j4JMIzJhKr4UdTytQk8yo8Foszz2hwimuypSDKY/Gn5N9IoyfiTZ
VbFn3NIbt3lpg2pNtuXTuyElcuXHKrmTi0drX8/mMRDntSCLUCyBAFIkk5XUWh+c
o9mdYXUDsY3yL3CNceZvcjJe9nlMjzpV56x91Mp/G3/7bOhrXSIIIWZeNnKAa3Ng
+lS8R6nXnfZs7xaYwMyRSitYS2DJXmtCOtTloziT9/E/PLY/BhVf3BvZcCFyXbjg
WqqFktMcS3kXaYpY0CMe+PAo5QyJjrWLSCZLiRc9Jj4j1OTzdkBj0w8y/kkEai6R
WAqnO68llL+kKkKX+oJqMkB83CwQr9Mb+GmAnluJOtrwJyBMdDvgimpQMiHRL4O7
u73nKhfnW01ojv3BkATEEH42c4Pj55bjl9cHNhclbGm68MWdlhXH28Po5B38jsTE
sZhAZw6wVgJHIavJ1BurpiiAKIyF4+O3xA/1f1FFka37/JiFYyIr7fK3Ykv+Y/v1
Qky/DLRazfBPq9h8BxtWJiKMscms9s3uRcezQ5S3oVburK5jJt/5DwX1xu58ijIs
6zhujpoFEVp8rz+nle5/1Nqy9F5qXJPrHL2+m+u8uLrWQyTOZc+6qlM48A8KKQj5
4wBN8Vma/UIJHZh3MBlpHguFfhZyCj9gniqwmuDBpRHzfVPeGcaQ9lcLWFmIWnmo
OtIByhU1LT/HQKTPbALsRk9FiTgKQfN6yozf7Odmz6XG+ulacdOIKqk7u0C9qLWN
cIYQqEd6BGT/njPJdLeKyCxGG/aAhYpMkhAQi+qiyosMQxWhijJ8zzdIoF++SRHR
e/fQHVpBTgEzTqNjxOUC/ZfHVJOzFpsDfAn8b6qzkUMhd21CdX9VcJha4u2zwYCw
RHTZrbeSRWr6LKa3fOqrYjXBCfJs5wWdhzxqPunwoEYD9Ex6h3VN7V1biWPf4P08
14HBhr8Z/u1R3XHeqRdjS0EhhecVTgvkPR17bCTxQ3rvtburKFGeurJv6UVgNo4/
LO7dOLhMPKuYiKAz0heVVu/otTd4YbqOk+kXrP1+WjkXVjAu3WewqfMknTyf+h3D
nxR1FdqZdSoszLU+rdtB2D3X+Tz3SzMh2wX7vuBX+H7ZDjPXGLaNFSHnixc3geDC
YCMbGBo/nePOJfBu8+fTCVshoDLiaXrE5ln/lR2rKKr7/uEFmvexN8rsTjN4lM1m
PB5cAJP7phUWBirnF+FAxbGwo2+RWdbfnRmffg3ZMHpSBEeLWY36yG2urSZkxKq/
RQESUdNZNQ7gHaIeP4Zp+LS9uD2Abz2I+QCo46JFlRg1MWBsX8J4rvunuZMP955c
Z8pXx/fzPEa4eOXMPLVsY1gUYeJTV/jMf72GNbks2rGWMCgXCihZ0Z60lKURG1Lh
54T/WN3KroGXgsN3BXn+jyeP7sypQE7wac34kJb9E8bWKnmK8xQtcvhJayq2x5yY
XD4pOx+eDreGTD38BodjKCrh/rwlqptF4+wIe3ghbIdRg1GywwXhmDi+444nR/Im
r6SEZsKyXH31CtZF/OKQo9yDZ4m3DayrxIlOtGL2fvEZxsg2smfRmWT2wmmfE2Kq
09WGXI7gjEskjcq4GZEpK1c1J9LhC4xJPd0hiO5ijl5iz4zVzR8H/3qesEymKTJh
9itltj8wJ8YKRXPQvmvln8Ki8P3mLBnQgniXdtLmkseYLTOm4Zv0D/p+TMxBu1SD
4gXl11dW5kR3jzKI9A4L8lpHw8lD0+T1lpUk34/cc3yuZNTE96nUSDlqNvFXxSgg
w81+tFG93sOPAg6Y9oC71IzbWeeK9453fElxmkiMUCysmjNzWVfEigCt+A4i+yRy
Ti/3dfeT20rfh8t21aHCxP1YYLNU93N34K8TpXXD2PfQJHufQ7erCK75gozZlN6Z
WKT5Z+AYrz54WjIPA8bclukBco/u44IJY46eNDqeynherFmBMotm6IRVVd2h8To5
S97rbSoHeh5pPSTSfweM2G5kqGiZ70Y7tYMSemZtvRU/BNTO2QxDx2Kw5FqbBAsE
hgTdHkiIi1kmljrNGqhIDaP9LCrqgyT4BaSR6gsAqXvpV8AZtYvyxc3C3QdmmEBz
jPUYI2BUGSlA+Tpd22HSVmWnsIgXOiOkz1iUEgbIJjtgsa0pAYOrRqYBHP2/uVu7
FWd8bK+1i3+2FB7EDTgWNMjn+49Cf82FzkeeIGKUy+6qRfB7PK/9CsPfLBdVwGYN
uuuEweo7emJvr/JXxgAm8SBGubLCJYOvkfM2xgqFdyrjfZH7+Ya1EsXpQ4r0tMKB
oUJE6Ov6OzlH5ciDHDSKp+yNvDPTeUoenrbUB6Ou7SBOBXcTPFPIOXulyEiE/j74
iJJ3+Cjy7AWTi2otRQTyhQwY4vrGfdfAQpkRqbrwPaVWfSzpN6MUw7G4YUqne1m/
eBMZ60NRNz30griFCAJgtg7RcyZyKJ/P3/zlEtV4Tb3WB+dfkRuST+LvvEoBRTW+
jE2O1jv0ckQIakxvKsaqL8TTJbv/I6CvXMZowKMyh7/dUJAmHIFj63xKi73pA6+L
hBv9lBZZxCZrivcpTi5JYzZehtn+PinVkU5J/u7xUDb4w4pH3+Ddj+kmfBWbSOeK
ZzSdVz20UI6R65PD88wWuwKMHk67g4Js4rfVodofrTQIG6kUjvC9FFWtR9rGRkSC
7tAzynDa1hp8KtjowuVCT9WjQYYsdMN1gB5+cjPgICP5Rib4YKbUGfV48Ov85Xt3
7s5f3R3lViLQiCKVXpqkeBy6iTF4ZKQGE8sUppJa4pEB4msGO/XW8bC18xCaEpit
N3XTIHIRxImFMeYD50Teq2Y37MZeAImCAymlIsrxD60dHloytlGGvPMzVKHLHTif
vDNtGhoJzm7egvxVqWlkWIaikX1xZap5Rlyw8jwkx+0M1ZsnOlYJgaRdAdpvgbGw
/Ftn156YSJyg4e+uOSKfUJ2/Rt3ZZpwzeC8haMKNMh8seyT1rK6cJ3DRGhfUznkQ
VgVS4J7ePWjxhRxJDowZFOMWF9gFKSaBFMqYUt1zq7AB4MWRx6Gc0ugFJHkbJudO
1B0jGtwpPpkU31O52juFPRg+nInEi4QHPYjJKJjyvCO41richM+kjXR+VFLxfQIH
c6HlVDl3HCPvmZpPDqUVB1vim507/a1pYZ3qnDBXIEEph+HTZTT5fdgHaetktnfT
J77aOzMnNOZIkCmI7+5ffjR02/t1N9p98WLSa5QkCTFPZ6/fhP/PSbOer5pLXkXY
ocJqb5AirovC1ME4C01pR5KbV2TgiO23UXDmZstN+G7ZwZiPxDb7UDB+A1qveqHz
2i/g+HE2QYzblpGcnHbBRCuioKXP6Ky2a/4B9dRN9TBeopMMHblsLU9PV8ehDwWa
BegmA4tZgKTnxzqKztZ/KQ==
`protect END_PROTECTED
