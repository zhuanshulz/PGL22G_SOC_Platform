`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/6fhFlAjFu7pseWqw1pK4gF21SXz7sHMUjyR2tcSKNsMXLKuGm8oWUlYS3Fjp++C
vvL08tq3CiGWlLpsFlgxmsbPWHpP55TDvV+RBxOCsKiNnuOhem7sCHAyedXVbXLY
P8on2B+NYExqvjJCl0Q7FC6qEXNsuq8deg/NLLG0EwLlg5nYON59nu7VeHLiy4/r
sW2Geajipi2OcZmDiLuQPFDi4sT1hkuU8UUUv/oxD3bEjRI1iVEwbTLuYmNoauzI
J4HfVvtl++lUS44Qfi5LPuNvzn6OlSQDKNssSXp+LDvZHNSP2JvdM541udg+3XoZ
Xx1VbQjOQuTFueEpGbL8YI5zedC//fuQCOmTomnYt7nrnitJeTr72B8U/Q4EZKNm
fk0gPLFFhjKFUYJtlurkvbsl1jjZfUM2VfoCIlTLwnlcTgbh3/FsKH8JosvYkIO6
P34+gNpWoKZ+XZxMqNZ6F0xvOjqPvuwBfWg4pbEZ2BHq6fXkJGk/E2IOzRHBkW65
yOInEKmaQXgteZKjrmVWvpx49bE/dtwkGln+UqkhjXv5Etxy79IYTSzfU6Azt5YV
istReBQUSlEU/sru9cbBpTH2F7u3p20kipLOP4u3HIWZAhn8BB20hkIfkOHdm+tp
bRP9Scz6lma+df1eT7A9Hlytks+1TlxjHmBIw2ZbPUMTNRPhMmrezDACkY0ijRD0
`protect END_PROTECTED
