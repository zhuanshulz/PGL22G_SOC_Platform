`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kDA/+8qOsjacIEDTkE/sprLF+YW7UP5YT//S+tPFYn0O5W6AlbbdXwZHYdAcnYrb
EfmXlGC9QJSOz56ySWcUgKb4HEQvhqD4UGY74qDR99DCb407nJ5/mjfSiV2aGJaM
MgutVHkM5OaqEdrs8e7647s75qtMZIGIQwd40suOddkOcJCyZjPhVqrvUKyjuUUF
RvCo6poddxbDknL+Sg4SMCzpgDPqSiCUFxY2JjluZq703uMWxk7S25qVWE13Fglj
LRAUmpUsCh50PZSIOyq8eKWrTyxQmr+iRmJde0xqplFYeqKF77puLd8E5g41Mvwi
FnyqBt0EtqluaRqdVukL778EWGBUKg5bLN3vkUQNswg7R2EfVD5FYjG9dYcIVlxb
8vi58tX6b7Xl6z/MEZPq5tznyz/3m6WGz+43tbLmVBIxgliuji+nrkjzs3u6zT4h
loOCGvuxW3O47F6C8D6ZzONLevMJX3zuNi2qT8AxP4FWvC+OKomdzTerBWCft87U
532dpsplGHY6LVdPxabpjuI2kBC7EbWoaqLLYFod+fcqWTd4IDy88QcJv6Bt0WMv
mK5nWILkyxm3AwBL/2HQfDMDgIGsMvQgPFzApBUQ82uVE0ZJBww6+PpYRIzdiotd
F4dknMNaZeg3aInQX/aVa/1rLgQTMknzTDqxszYPd0alj7IltISzPjhrE8HmST4Z
vGgi8OtYp496CD9obcJEmQm6nxVNMjGHoUw22Ey39UNk05UNkUScG4haty1lK/V+
60u0C7cf9E1TevHdbqSV97VMf8m95B49VsQhrQTmLyez+3RrHtEaNqzeoNvh3BtJ
GBb1DAEJ+nTruzjkJVcmALvgAahv96WHug2z7uDR+rL7De/4dLyxOLxWKXle10G7
Jk51BR4PXsKbV+x0QkxMPqLt8K1V5n9SmpXMKkeYL5PCM71kuZm3y6165sHQ+NM8
EYORRvkAHP5FpoSUxYNuZIVJwdgOe6QFcaiMN5K84dpIBYhwa4FSeXs0fWyyFVDl
3t2FzFI0pMhzvUgFk95Yxfd5sTHNj78wDrqGa1i7gYKDxiZKEtFsdyzvCI2ggH4W
r41Itis9g+E9LDTIu3XEqdas0O52+LvV11NM2HWMwkQloUpFNqRXPMxfNljd96uu
NlArm6PlgEdVSTcUwtkv8TFaiUuSbynGJRH7DorGG+qGXAeNmFiSfto0ay3S70sT
4//G4wdxiahqLdux4vz+YO4/KebwZ+O4xznkP0yVAd46P2ur5bsH6eBdMRx+uT54
fUDxrGt+sF6Xqvyx9ZgfKz/TU6dYX2Oiq9I0pWZcFrBqgQhdR2ts814HdMotzHnP
BjZoEpJRsGQHGosDSAHVCRwagXEktf6LPl5IYbmIju0qgqK4sENrJYN0n86l8/ST
cDF519g4iRh5+3zWHgzyUCTb3IpUjyuS/leM6lRUeIhsXJwEfCZXhTdocnpk842g
UCSUq34gs7Xi3VIEWhfHRwFzCxyrqRoOqGiaV5+r4Bkax5U8oaV2Iya/UkMc6PV3
D19GYhWQ6Wvef0MjId40qzmCA6uE0VtdY+xY0Nn42R3OlZcROXa4MGekCwnzRIyO
gJyEyjLatLjzhD+bTqKdvRIInMaNUnifgX7lgGe7LljqUL8Z0gehoItEU+49xqFN
x8hsFZ06vpm8y/gdg5mHVKy3o7aLyj0MnnO2XTN55F2aznpndnMoxcAiTQJwH12v
IvBlDPChHgU8u960QTXToDOoJrM71rEBXLFQ/sSA9rFo4pTwcOPlyO6ovgJ64UnK
uAMFyTMYfI7uGKxm1ImVaCvLjbLsYsjdV/gov4V2WPillg3bBc0nb+TtNDDF+bAv
sstRYlg3PBm3EgzYo5Bp+jEcDpBgrK47ocQH8YcmCYoV4Bvk0ZvVxoryhYwYT/PP
G05Wa5Ahj+HuoUexxL8j+v3YOAeBttH8JnisEVEXqk/xnIvF5pkcGmfOB1w1vm2H
6K5SHn4BQxIiKTdK6Q+06bsAvDrhaaxG6I02BvIKJChZXt1xv0lo9bDW9aGYf1wU
6cC5vbn5RNvyanVw0LcFxcm+DeRQeOu7rSn/hrvN48AgHju1esLbJAyTYy32r0aj
p5Z4UFWx2deIE6oz+WGTtPARkv/DsWoqnxzw9Bx2/yFh+ksOW1bN91H5jN5pXYLD
Pt7W5BmLiupuvjW1c+6//lQpDC/fcrDKtdCY0VVucQoSRs0IxOaGjhnCdZFYoBUN
/+YNSMUhZyTp3a2HDbrV5fW7aJ7Glhlm5KBFp6CsX/2LoA+wLm3frNp95p/4XdoJ
ABah9GIxCnwhXzd4hlRjznuOpmyNQQV9PWXhKsgqI7fS3mIdJ+IW7B6F2pgc/vgR
`protect END_PROTECTED
