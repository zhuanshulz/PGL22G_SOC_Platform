`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HkiJdGCIQNegxiDVsMgKiDhbsnCC8IjfN+1Oc7k4eKItAEJuRuc8hHMzytri9zju
M5cjhm/OMuLnRhgEiFWkhW6/tK15tMfD+HY8QLXNlbTfz1kuq7w7bKkWE3OKLSK6
MWX8/pRWXvZgaSCDcSqdjTfUxtj1jL/sjkWwcIqn+6XldSaid2ui4pmEpnSJxwCW
tZeWuvCWFhQoJvA0Ur9htdSM+UI6wBHZwk0GvVmkTcPnjp899TE7EFomnBdZum+/
oNR7ZkrPwg858r7cwQtPU18LmdMZLAR+wISgI0YNv2dcpV7H3QfCO0V9EyhRqP3Z
isIFXCutEwyOpxXf2sX9YIV0IgnioV8ABQOpPEVBTykMbLKz3xWKqB2tcXDJlXCH
9pOYYVOj5xYAWFaFYXtutGVAgOnIS3hnwxVSPwcYMNKxiILpbRf/jHd+74zBeqw4
6Gy7m5eDkGScxs/NDhxSukbYlrI4U/J95H6eRvrG7GNLrtSQ4BzMDpq4GatqeC79
aGY6WU5ld37UmCGnpy0QX4K7svGMYgjPyUsvlj/NI2yY3jKyjAGExqISatIRE/fc
ncNFPTZAfQdNHK4y42DIm2LlzxwUz1Od8S+V0Gx/G35JnJZe8CO0gg5/tpoSsySQ
RS6+9ti/g3tMJFSZzd6ORafNFnWp0BbPzPzK6CdvP04+orGBCkGIdFI99GMC+//H
krAeRe4J0wZUUOJ+EC1DbRUTxi2o/X8m4cMdKJqohFm5dmtGHQjH9/gQYyl0aKBn
9i/LsHEMQkB/bmPFpJ9VLvekWwa4260wNb3cgmo7A6erBiJ1Y1oBXMIR8KxAaacU
w5WNYVdSO5ms91w08FQHxUUCAHWmR8LEfeB3kFTC0PcHzp6ACUBHMNgq4EbPpID2
PyhH1Y1RGRyZYBnIEMYfTW/tzhaBUjW3uk64lZ6P0ov9xlVr80Gq5a8AOnHnNg1/
IokIGG6aHo7quPtdzcbR1eOJbO5YWjAwYIB/SAkwD/R+Dcc47XcFVQGHDOetqBT5
ltR8XN4yNqkvgMZU0d7z9R6OsmSolSX2qgMjl/pQD8j+5bdAiDrFgZV/xXNBf1C1
WQZkpScKYuzZTX9HqRHzX//XhYGE85oyxsfknLbyxHi68ecxhlds1yYkRyW5oogI
eEsPGYBG8GNuXTFbY+y0DNEu/AmDP2IpetddvV2e+YCTrJ6TSAdHDOaHYKXr6hzj
AtbnUpzjZlkf97hZJo0pJnvzWYTQiJ7vo/WTtSqRLkeXFud0hvTI3B8455r8Li9w
pI07qbL9pYCzO4iY+I+QSB0FVyqOq2i27wOYMigNvF5Yy/+xGHnodN5sCBQlAMFS
BNuBsrjvrKzqNn//AsCSiWBgmULUcvODcGZn8Fgx2aYJ2uPmxx24wZOKi8+vX5LT
bTWwfLcuI5iw67LndCAQl7xs4Nrl/hX4V5SmIaMprK5Ah0/x4/FjxQAajjDk/FrL
7ElsS5Thiz8FFew8OL9YBjVQai7b4LWEXMiiK0p+o5Jq+Od1bquonx38NWmukk9p
PeviwJldEWIQdWg6iVdF3PE2stg3SuKf6CeokCTWV45dBSo4bsfqZIA3gMw/7SsM
EfFKaFMTHxQcuhPpdLwJq/a1niNqX7qBpHcFL3qe41Y=
`protect END_PROTECTED
