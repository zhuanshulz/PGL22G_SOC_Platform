`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mC5UFd7CfHHnweK5QIHP+S0cNi1oRNlt6qW/FVsm38yHeuY46n1cwmFF7aYTcCgq
TKrfdM7/xggLdAXJqUwO1fxW+CtAfl9E1zU8BgPsFIe7tTVLoph8LxMLIS/J6gAH
GU2DyKttVAkMxevwNN210E9gPnoeTeitp0FE9ggq2344Xs/zjV9QrQneD8M35omO
uZElR0SOj7vKcyJx+UGONwfRAnc8PAaV/NslZjjTfqJbMqbsTE4+6CIx6YL5pSN1
A78cYNBuBdr42bHG+g6kkAw6CRC5WRXumZQ7KDidy2/nFyoSW0NDA54KxbmQlyHk
OsnfU80nZkKNa0lC9g8J1oCbm67I1ylwo3GNymNn6YFjp12bKbEdiHzMGZm0ibG0
FiMb2+4onUjELNvr2d2bzduTxkO9/XiKDEBPkuBpqHCK0TVuIpjYohLSXWP58iUC
Wfgi81KvzkHCN6cvQEAZ3mEDvnKNTXTHLkafYobs1obaRzUeDMIxvI4VjleSUN8x
Q1X5yyn8vF3KD9fXmYfDTVjM1OUZZnZUba3xIFhxRyYqMF0GhJXqWB57Ya2Ac+M5
yQUOA/M75aH2vuSyUzOZdjy5HaAsntQaCYCn5Nygy9zYFfjS9E4MVtwpsYJW1r6t
SFfr5aoBSleTvToTPSVFF2GcRrZDX5PYJU6mb+tEBicV9MCOw5HxBwqduieHCfXl
LtZfe0u7c5AHbdm07r5S4+iWahYZ+ieQzgs+M7Dy4hvV5AMJoHFxAUv7Ru9QaYCh
iBRExzBQfL2z4wx7kgc16VGpCvxWer8mzfq2JbkxJTmX5Y8fYggP0/pqkHy+LZL7
7NOKK0V6WmEvLtTbV51ixdK3XXmhU9jY20rRQY+7LUuiOnPNT67KCCRk33q4uBu1
lTMYO0396xyvHempJaMsUKcudNi9HADWTHY7n6GoJtl1M11OU49XjW7w6yhn5v8e
VPnpJSWgIqYCcN+dRRenAmh/7R0+owLG4ZpyozCxgwC1lFZU4mBwHSPrm7Jf2C7L
BPzzfvPduvEFyb2cEg4R1/uEu77qvOrrHrXsVkbJ1vYgRhip+slIFy7NX2BHTwHN
Y8t+SRiDK8BCaXQ+9ydm3+ROePSW0LlLMth1Q60yFZrMAGEKsPLRBU5lPug1X2jQ
rWtLcf9cKmjlmS1QHj2oVLX3aRPnbgwf6re5DnI09fUe5sgjRWtZ9Kyg9NJgTmlT
cEd3Rr4ZCSdjLNYFKK6+ZT5GkABp8JUHpfXxBeC9OvJ/keko0RFtl1o3GzgzC70r
NqrBJN+xkdPYCi0GjR/B+bIorXh8C1O1EliHNcTEWv+HgVklqV1s9Z10cCMVhl0k
RZzoFZ5IkO1CB/qnUPpoSFsvZPAui/p5rvRO1csJD9zhbLQ5ESPfp9BTEjWnNmhS
RlNHn8N+LcC7SpWprg1lHvZwvZyLjZeGEesVLcWOdpQIJUSllXAgCpr1itDVBG6H
9FrsBKyjjRUxJnBDFneEW5qMXWDVABf2/Cwm1DUmpNEd7BB4+pumJcUJC3rG124c
xRsc/i3O3JDRjYC3/h0CNyTfCIJ74H3oax1k0J/kPYGDHCvPOWZbymGcg9IxjXIu
406A7Ip0T3nrbf5rCKpkW8MPPYSiFeqhwUIxBGAXsvsw5tgJelVzXAbyqfaEzF/7
Ol33gWxbCzMm7tWfHxOwr05sbuUU+mqwkfupMso2BjGZpdvTcjNLCQs4foCzwoQo
reHz0yGjL0rl/phmlxgJvfcy6t2HWy622XCIBmXDg9cbWoAJjuhbU07uyvCcQ3Hs
eag3umIOo6KINlZ7T+sSsEBpszaJ7UxW9m2uIFcuxhCfNhVhuuqD11BCAPg3cfmG
sWrig3Gwyi6e/9RgRb2dvvbFNWXEEbNHNhLytBwEIKJ5mVpbPR8N6nepdMA+Vht6
cr4rsi0e4/OjSC3t8v7PChxnYHelT5uKXm94klVHoyukyu+EqCjXQFQMeqFVF3QI
Be7SY72QqjNNyyfY7RR6YgkWEGDTppKLUavq+NIIpS4UEAQCSRStzfFwdAEqU0B3
W1Bablqk3LtX0b+tZEFobOtAZ8dv+xiYJXTSR/HhDtIUI2XGSTWwOvBIgIfzIEtQ
Sl24meetBw/LhYl+N1+u4pXVtqYqhDKDtjjRsL2Ti3nRIhoYZ4FYLu9ekiUb/sK6
tfGO4La1VhNRpzhxWbva0xgcaOMbMO2OIX/l360rIq7un7OLZvqcJVByUo6ou0Y7
83Aj7Rh7MZKfn3P+O1qeDYxR9QETxzhmgtGH7Dmf0BY4MGosFOMB1CCan0Pk0j97
4lKl/IYxaHglbO7K76rbmNxY8+J9bvFJFpiL9GgKuxSWzWKvWqwIJTb42OB3dWHj
CnBDwDvFe3G8R8VjjbI7LDecxuUHPYaX4Cq1Ptx/yQS8cwW1Dka7GXLSrmZDTi5y
rzpjEWxWR/QVS3QAlSt/Fj37wrjg61GWntXatxuznPpjeFPvKFMPGeNdjDXdnnFm
SXhKokwOhE6wzm/kUGqtvOYZXW92iG7Hnk9EBx2tSNG4ROIvuaIORZ7+otv9t1/N
P5dklPMvNb+YQqd4VprrRZyldd2rremsjnWl/oKDBmePN/6kUv/HDluty/rSlfwn
1j5QdxvywA6cypTaM8mv4MCfnlMD9Vo7tEE7rxw3deHdag4jkEbEwSK24NhV19AV
e8zaa3B4q00W//awVQvgXu39Gx6Lo6TqHHjd5BPm5YRhH/1GwxM3JUCmEKJ62ctB
LdDAOeOgJ4jKUq+RoWuOagGJJFuujoChaCZI//0ECJ87vSK+Uomqs55ThJzF/7Sj
PxFCDyRVa87jMuTfahiYB81V6w8V0B4sEs2zNFV8Ya+uKkQts2yqLWLj8CCKeo9R
7V0GuIG+26VtlEBVVXV+YHMRjrNk2U5qApVERoKkEQrx+fdc4z5PCOMDFDTZ4HTN
42MELd826svyvwDZeH0rl37WjO8h3zer+0QqLO+9KS2RLtwi3blcGWQfaqJENn0U
6mnvhUcia8+zz9fOgQEXonsU24dpbVmX2HBZzXIJkqlGP+KG4uWhyumgGtPWi6pT
qiLbUWP52cdsphccZsw9arlEigssqBdjWMojjEgCFZrlvrXh8wSfG3yz8g3BnGTs
SpXiTisJYse8t8beRIPzvc8/ODW2bjiav2KlMZHapPHYdPvr/iWCeWQtQqcAKFyf
gCiAKV6kEbJ9Rwl7ZqT2I2ytezPEmYs0Cb1xGuWkpT89ZyZh4DJe9PMyaN2bCbnr
tepLxeO5FCw6AW/4a27ci/GzNu6DBhtTv3noDVzTTl0LNv3602JDOCASRaGe5osm
Wv+jE8M8JBvTPwsCyUTpjpSF6CEZFfJjtLmigZ/mb0oCPcKPP4L5ye6dfWNEfUpS
CNRbXPypIhsi+LBYnSRxrpV+Jz7CZme9HTvQh0aAp6Jvs3xr36z+sCUFOHstolPG
jqu8DVpw913xxnhXntjbZZgIalFmh0FRZmdaaRhWdiQnWqiOHAFi20voRhOBCGBE
ow0wT+6k31pl4OuxAHl5X7h1YZRhGCmQCcMkuRzMyDeBbAU5SnvgBnlZ1z5YD952
wh1wWPs0cKe5Kc+fv2yTJECsZ3nJlwSBvUHF9yFYJp9eP0Rq41CoDPT2PHnpEHL5
4Yd8SV+y/rpUPVm3VAcPQ53icqWGoqWMfkI04C8b5ez8Op7tKJ7fGa/S8e1XdW/1
yZDvP/h0MIsxICgqOVfySSyJhgS8ixQRu0DkBQzo1nArs5tIdmMAatkcjjWPoIEm
JAXQZ7QcZxj9YtZgvee8a1zIeG+aZqj0D8obAKRnX7f0drEKJVaQXnPHYKLWqDEv
/LFu6j0/HVXGOw1LIeXdRK1r/xhW5Ck/XvzJ/mqaXWl9f5uqn4rXuuC3h1P2G3vn
bipAqD/pW7RVwMcUEplINLJXB9+g3FndhO9SpuGm2jwY025ARfpl8il+Fe/IAezS
32aTqd06CmnDn2XOzr8kefJwZIUGGyMr3aetazRjLnRpkNa30bX24A6rOCYq+qds
J9ghOpBAcSP+kRzLpu6yyg5coD31sItm8rRyTeKnbMK3NKOGxQ93gal7qCpbIxRc
M969ujYXIzdfv0/d6H789GQBkc2fsAjMcEw4HXLFrY7FNhU0SLAev0Ymb+i3rrzL
qXDkfXYYwVGKSAAYduJoP+LXPbAR5C+8vfnpNeHqJtWGGzrERjPfRTNA9XznYLCh
WCNcChtN6En6ZmS58QpGDxd+UFfUHAVGYN0c+gFNrRsiRyPICIzO4NtJRc21ZzOo
m5GB3JHLFX5fQnpuareDgvEPZQMySPknyx5c3lU6mYH2Lui1CrwXzmAVLXuwu1SW
FnIIdSvobtn/hOTHJJ4bRrxybPVOZ5OxrAif6N42rw2x09wBHFyyDHHgws4VUzfa
/TFvQCi0R5poEJhGQvFUFrMkQF63dDVSPaiEmooi93Z4ijcVCj11Q5EY6eFaztqk
ST/24BUMZ3eIMvyg3vDDEvjutYSCJgIYABk1/3k5T6NTklxViUQv6hvsbqfZeP2M
KhpwrFw2AtueRsCXsohnp7CHZ1cqj371qF4NqYicXp6RVA6jjr5hGHwGDwsRo8ts
P4kbcUjNM85fb9BBPekV6jlEOjar9x8fm4do39pAbCWElLHspAqV8MM1wqmwqV5t
EEsmRCoS/8+KqysHeN7c0e9iEDA6IL8SoFQu1ZfvNTcVDzoD5sIoyMBaAbk9THPk
KD4CHr4nPdSTMQ7t0HPnOkSKrWopNQLG7pSkjSqjkfJgvrZ+YZ4/6a6id6hXInkl
reALJz/ZFC8qxuXv8asMJyhXlvPpUw02DNlUjGpmC4ERqBCytJD6+pl2aXdtFNwu
lzjAhns5ZrjbW2JlegaAWKpI08esHHmPKMz2hFwQlu1kYtEve+3z1xJQthIIMmso
zgJUuqZT5bnKqwlFmlWrCbK7skwIfWQP7j8h4U/PkZIdoxUJLlv4KW9A1G2KRBLN
`protect END_PROTECTED
