`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WJUTIbh+VGQqcmEer8ihPfsUcN8Xd2qNaz0Ik5v74R/vnsNVouPO3VhEbVHktt09
Pf5/8o+F6fbCxw3zdVEZ9ZCeakV2/x2XE1sdEeZvZHn2s0RUA8Eng0G8rEHhJIhH
a3V9YRLPBDJgFtQ4dL7sTxgocsbkDig4FkeQTE1unhAONFr4UBRLKX5QSsfQArv/
GK0bvexxa4c5ISMJJx0IGINcqoRM2YI89qnhMOejBv7BBNd+DexMK6poPnPZcvgs
ECs9qK442hegI/ivMUGqf/UbWlZVaorJ3wyC9cp4/2eU6+7/YZPREMQyyZw62izh
7iD6/eMIGXmh9a57JRpYVklb01/xy30hG8Lkn0Nxu1OOva1pABggknD4qJQRRb6E
ija2GuTyPoaQ1ejufqYzakZwtH1zoiNoWhCzsQfpp07h/gEukkv0TAKr3F3FBtKH
P99uuOc5XUD0ca8Y5y+tmkgighQKq8b6Lgjr5fwvOgP+MY7ms/lyl/2Dw6tihLWm
TygR2ZGzOYiSzH/MCYhsjB6aDXzyVxOOBxRiOEY1zrAYiNpEJXghSNhc22/wUGc1
IXk1JVnSCeOy/aMz5hrjzQYfrI3YDY+qg14DWXtD3K6s1n0VvbFNIro7jK7yMTdW
NXZiRuw3133nLgZtu8jkQvNXATtcJI1wM5TwHj7i7PK4EAjZObtGd7dEt5626z3+
hjoqDpW6GByb7s7fXAQGYiqk6+bmVEBB90ihe+wXRT0=
`protect END_PROTECTED
