`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yd5vKeQJhW67W3G9nSgkwM/fnThLXIBriNrWvR7lg8WY1nCcrKUXD58dXKrnyfdT
vTGmosIKaSpyEz7gEgh0+poUZtyKZtvaZZuVXc24AobEg7Ah6W85ZxsaG/yCuTxb
lemZ2vO0fdKCaAGU+qJWHz7V+QjeKkZJJ3wi6G3lOigX7wBInO5kV0IUfEO6upqx
ZlNWhvwQYXMz1AavvAA6UivxAFAviyhzy8pM2Ze12TRAYdRNe+3Ubbf8lxRETcta
i9R3Q0RqOGazWVKTfkxjNbepaQAM6851JKmn6l7LTV/dKQVCKss1p0w4nzz9cCi2
TiGgs/P1w7tmpvXHCr+Z9XR9bts7DIbDO9V7vXcGWH/0eybFJJ+wOG3r5v9sa5nk
zFoZpWkDKr+qcBmO8iUIQIqQef1ZTzUh6f3guOdE78xPizUIIq2hofJXdF+x2/rb
LNeFnKBls/3kX13RdbRs6wXow+LN1ogjajLjiPW2kZZXa1XxpfnqdW5FMjl50GX3
Vz5pWwn3thdBag9zM67VgpD8Zpq+VRi9okyo9dhnOKB1IeRIIc15jP9S9lxF4G+H
DfwEdvs55ywzPukzmCnhJ18vyVLODll4mbeD6FCzjWg=
`protect END_PROTECTED
