`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KiMI7BAelv8EEx4Omv2esl/sqAOJxKvJUOmYFKbZlmtvAqCUCn7bq8VtbEY+b3EM
fMFMwTBiEV/x2NiOlIymVhzGoaa28zaVTcd5+/EkTMPWDK9wFi4rhvkkducM/sjr
LKbw3qtjj9XlwJduunoc4OMgxTgM7dV0+/XQgqeUDZ4vDIZsbZkpWr6UOFiUGJIh
hsnsJ6PadTVh0hdQfmjCWpOhOvX+7KbyAhhIQTLbiGuYSfy70nzDvlUFFU94yxJK
SL+3Vus3sid40Yy8/gtmWwebuEJZID6j6l1REeX+LmCF1VNi87L+d2aFAF0hXj/y
tCqnp53WZ4d3jaRdpWcJsqzTiMq8JUOwT89tyjW0TTmTEO8GKdveNuQYBf2Rp8l9
GGY39hKY6hsIVFwCXf35B4AbHyAkN5eK/wOahHwNJ+efjZKoDSC96EStlIkpHlNX
O+KvYzC1rgkjWqQI2wSfyD/luUkzu8ZdKFH2jjYWmsu+5508E1ggnZts8EkxWhD+
0BZqxort02hDyCpZsg/DiB6aiGEgtBSQ7SX7Hn4x5XIarfRJhW9MKD9NP8PyoBZz
YW5mDwpN7qaM92Y3lTw+78UBbX8bwfsnHS/FcF2jSu6U6T8gUPxGVa/JnCM9Pu+T
fDnpbDtDGJRaeoe6T0hNIUQoATnFQXDQCtlRDHReHt7iU7A2v19wkqPlbFXAGc9x
PNugfDYTacZeyfqQZw+nerRtER0chyloxUwg4tYTTAt2fwus1Y/YqIk1HTNJyKDL
huT2oaI8I/eoa++cpBry622WbB5INl2L8DOiM1e+KYshlWJxVRgo6QOr28ZuDByl
17iZHX7up22sPckIzTwKX+n9v7dNUYP9HykxyKITtclKGaH1AfOjCzZbPVIT6IMt
01zmw47zHUjJhipfe7GhIqJRl51ZG8USekflK1BLv+HlW+ctfHT3QgjFtjdZNIUt
0ONOy2OdhQnoG/HsckKa/kzmJcoSJoAf2InlSmcT/SM+WHjhHLG5MEtzMk3fgL9E
hAt8RhDTACo86RGyn3sb0+vlgwgmcRR+ADLPf4UztybZfEQRhXujAgwqUKbYY24X
damEQ3tPeba20sP4QKI8CIfZYJb+iYGvqcgu9VSHBcDRZAmIM/zvEbJ1AocGKdB6
9gjzJcLWJ9oQOzvDi4PCniXN1tgWZ5XO2bZSjZ0TOy3NxoXVlTwUakEJUyzRCDXo
JlYhhcbV3Q+dDCSIyct/l+sFZc3JNnACsPuMrEg6AHMd4pOjJuGiVdmXwxxwVvAC
0d34L1Ii1pjnZfxNZVvC70oEKjf23PSZ5tVTK4VW1ZMWTY/UCVuvpDK00Re3uBHY
oUs88wD2MY4Jp19aDpkuE5jwBBJ1kqOWZW7ZytUicT+ZgPg0vDbiVMIXASwtKacH
LsST9n3MecHM9ASv6NWJnjmOLiSH50KrTBZDgZB0YoVaKMA2VuGs0zb4tS1rC5kc
KG8lRsSg2rrPc1wcqFtCp8j85CatFwYz14vfFXPPtO2nTXNZoyM4/QvzNGowgKd1
9LX9Oc5Zm8ldaLrbJxv6q98t66xzCk5shmQ1Pzb35wuwFfZ41ojqaGJsizVxXTuA
NcB1jYPXf4olmgEbNAUMFer9cphV0VdAR5Wpp7eHmqJzSUKKa6K6gbtgydzGPtFj
ui+CQ6TuQXmkFDbPj1Zov+D6Osyl2UkZsSU1crKYStKYuTGdi7Bbv0Kl7/kN5NbQ
DuwcqW4Xn+S+5FVz6WzziDCGcyg6HPjhGUxWk1QE4lQs7SozwkFvnHy7KurApaqt
UxXllBeqHx827ZWYqTVPCg==
`protect END_PROTECTED
