`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f3o6+gCB8gFeIBvZs2zbKB11HXh65iEYiQorm4e1p7jhz/dj8jVjOy4seRbYIFQd
CNN8IaNU1ozQLyaAR5dZIqiiHIKtFBNj0fIHpVtqvkMfx86BdqgLaaBqRzwbFXES
yZ4Ca34MYzFSbpyJGJzD12kdONKkQwxTiRUHkXHjLqH70Xx+BTvvK+/QSI45XH3t
hoZUq08E+BefDztT9FSnJztCdRbdcIPj9jDXYuqQtYPzhgVsALlQRHfERoFtvTDz
e5C1SZ7HG57hC7XWD1BFq2KjVG1XyOC8XWvXOK3vJUzMHIcIHdJw2OoEaGTWcOYV
N5yRhMb1HFPhvDEZwKE09TlpkhjM/LBVcdNayV7+KxTzmt55Bc2HIpQF9UlFr2fk
ad85iAcUaxoyZ3nOwnrCnAQjSsdQPRd2lNOZ55Gm6U0RPQrk9HEYN7s4+QYg4Nc4
aydgRqdTwT8HulgF5Vy5YrGEWY70phBK8wqjpvKncU9aKS5u6dle1mDMSrjbSYMO
sr/R4auhCxQ7+k1h3DF+iEYL8mE6BYKIZMX1N3SFVOPQN1K17rvLwnnTdd1woM5K
mSo16eRWWiphl6ScXY3J2xOdRCRJRUrGKRqyn/uOUrf7hrSQ0Qhw81OgjzlPw2p9
DSyHHcr0zKOexfbHxkspRJAjuQYviXa8gKsaQ2j5AYvM8f7Yf0Of44IOFliKuiiC
HJl+Y0YDuq91BXzIMyBAS8tf5FJQgFppXb96+cSvQpGF9yG6qWs6ZmwJmqoWc3V+
udHMuzSwVPutHzOwMZ2nxIQT9RCXtQUKeiD9pZXwHdyX0KGUZDuAjkLk7FdJTpke
J08omQf7ENyxXGx8iKwAeWec1TOLUYRWtOx2vb7djuKLe7jKbZfpKNEWlJHBRYXc
nemKToMQPzrSCsMI1vep6zm4NbJ9uYaNTJOVH2+je+0GwU7BE24YYINdn4dvgVRQ
fDwbJoz273xFYzFG/YJ4k5Ys3mwYQmHeeZPIohB6i3DORVVG6WryNIhkk8pNM2tx
F4TVDEXWe5K2X4fhZV3kglPLAFzOjeoykTvQSVsaBs7EpelWhrhLamC3SUUq1BnS
MLRqQzsBsS14ql6FEZermMakWyrRyRskl1NJmuVMgeI5lSF1hywiHhPYVMxq89UU
e6jxhORqydDIQpbO7h/MQTjCDXmdye3V6e7w7mI16ER0/eqb8pHLCc0zngGcIvgn
4gsqm36Uvm40k0bXNsvTcbxxD/e0iLX7iMFutIDEnmA=
`protect END_PROTECTED
