`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zYk4KlghHb7DUt79bsAgQUtI/0c6WaUihW9oE/xYDn233fQCttsv3qQAri25jBZf
UJN62uNKW4pQdrpKCGQBocqLFJ3CbkAOW4ysjMHbwlY5uZKbG9x0yY0x1jmnReST
pyqcLZufZ3uXVMiJBHQ4o0oFayhMWARvVFsyfFD34AmfTyQY1KjuutEcqnDMlRgY
pZ8HOLJBaRYkMjwIeKfa06Ff4nlZudxUVATlb7dw5LvZ82G/HWUTVmSia/niCno0
fSWW/Em8KO/SjjgZnGquFChQtzeITh2wDP/MXYH6gLSHlrqS48YYBI4rvv66Kbno
tftBEglfFyQ3h8wd21o7a3io6/ZzxXWeNN4DKg3t8cL9IeR0P/vR36+XNFinSLJW
k/jVdg5xNrKFqlHzw4XcppV4lJQbpaRn7jqpnBcduN1jOkry4MzcsdjLROXQvDU0
zVIzuGfuf5hamfbhmoqCaR8Fq5ESmTmo2qC8n19lwKzUeP9eEGFSsk9bXpR6TdRs
Xetc7xkkN4VYSE5NR/BkcEb6hgQmqWiOGQDwN3r2jzX83jDM8PuqWfVptGuE9pdD
2+iLAbtj5senXpeeiO6jmIBvMf3ejKGDlohRt2tvLPY5O0IAzBwFq5qi+XK8kj9i
p1KoyhAemDurCPd9ReYhJpOHmg1lhpamejCp5lfn2KwJRvR4AUBbLkpL8iR4wr4J
c8u890wqckc0h4TZECr6R6I2mxPXgcM18r6P7YBGy8zwFTmvZ0GjjXoiWU13Sj8V
HXKRXSdRBTWdfgTWtqE86aVukTKKH7JsJYn3ud7sOnYF5IYZ8dfOEQPQGb+g8pnC
0jp0xPSFSZ2OHe9hY4Zf1NtHhwSq/eOXkWAQnWUZQBo0gzy+XP7Ja8ctcKWM9eU0
2DOkqQ5kzzCjFF3N8SmFPFxhxGIj+1EawTSaRzHASD5RrznME1wN9oO3Dblovnan
NDouS4aQoUFWcPdMCF1QJym4DBGakycbgJ1L6sguuwetMOyBUUbJxafZiosPq6E5
AvNX4MrRQQtIvSnOlJCTUXB7iQl76d1eZHQ3IuJlbYRUWQzmGXPECtbJobt2Tl73
klKClurgmfhPwuIweivs8+JHcZBCi1mJ5y/qgnCUlb078jSP+2pmklgiHe0FYK9Z
llRv3FF6A5JG6HdOMQzJ4jZSdtNvtcOIhojc2BUe68DIATuSGecBRD1STDn9bHeH
lxwMF+ta2Qaq8pT6UL271lyeZGlkPaZZD8hgKj5sc9+rEsB3lWI7ETnDbdeCNlw8
1437sEo4dciYe90S5RAqfWtWRsf+tCvccBZaDv8ZCj0oMihqvQ8ion9D4K1H257U
TXX9vRDnz8Vyz0z04ciDEaP8Qwm9VzCVFydQJ2dWL+IhdObtPLUfHUOId2JLpb7O
k4cUBpdVdgptJSU3dbVjLQExslbt+23PgQHa8X94c10Hlpj7+b2FtwvLxUm/8TZq
AB2LpmLtI/Fv2XKchyehEn+VmTlX+gXM2zu1MVeF0jz8GHp4/efpG7xXtaFoL9GS
RDpNA1uqG9KRuiN3mZauopHJ03YlSg/IGflO6kPzzTpYHmXaz0xqQVJnJibBi6m4
CqD/MQmI3mRDZfUa5CM9gAHjXCL6Bc+vH/EHZF1uiMDbvD9Cuwp2F2MV2RARjICP
YRgjYECTi1175nLcVrU6QPVgFS5qSmiY+9yiDdXPZEuN3Zt+K185MBIFlbuZg3dY
Lo87iYxz8KP30xoFN/ciR934x9k+W9JnqxN/Yk0gR2WCHaRMscXcyfe4unMKb3Gq
431mkLlhkA+TJX7DCqJZ4A2Kvf+7xYvbf3g0kyAdz89W3nQX5R8DKpSnMX3mXo8u
hKkt4dsTv2xTT0wF617oE3M7eK6q8e+eoxHTaCw4CcJPX1gPmQFmK8a9pJBicluM
r+Kgq4HvelBcPYplZgcDrkcZ5QcQ0EIrTLNXw5INQXeTd6JLA0v43+MY7+jVFa7u
WlKLifZB5nx1obi3wov53sE/feNSVMVOXwr8hYmARVfAfztl/Rg6bc4EamPy3Bqf
+9X7W7tMOn0lH0Nxa22NySEWc9sSpI7OX3wwJQXjeeogLSeZRx5lV+ZjezAwkBXK
kwID7RTKAFDPvmLnOSHx/ZtmZvUwnju+F5PqjPWssB2v1fsHYTe8BbiTXkW0C6gU
x70dQksuIspUnSPIdWJ+xuR3q1Ycfi7TRcZu5nBXcZZj5yiiBbPlm6FAom2AvB+v
xXmoAqjW6UeaiP2DliyvmS26gRYpyi2+P52ppJXnRuYwuqjMi0NTFU+mJ2/vtBYp
l61NiHRUEaXZT+2j6xbmruhhVigjik5TZtYaVG+T5FZxgisoL3eLamZRyTxtjaDM
WLLecIl12VxYxidfTzJI6eJI6t6GQNhgIwkmyHJYf0mAVdxGWpLcAa6/MFFFlRCw
CMNoVrMkMHmTo95MToKEVW5HHmfY8VNRLTJVCJrOw5y/suL3Sitgz5EtRsJwDYhg
2wQrVRuW1zqAXDRs5rBVF+nJbK/pVCm24gtjMJUnhdXFGG5bGHbWrgLQkS+12uq2
/uPzpOrnQFXYphQ/pkfRFPKqrhNmmbSgZsyiJyO8Q9IBDMM2sr4SzRu3+ttCje6k
6SWGTSfmVQcCM2V+pERZZdQZ2qkc1VZOh9k1gk/3pjjbVxcVR3hp76Lm9UCze3E7
bRvV3I0oD5sYXn0vwARt6Phm0U9KrUKg5aRD841i+6ZPnusXqnU3vnNNU9wZbFl3
ZObA/uRzh7mNzFvntjUc32/lmIqAVbr/WzPZOFz9yU5gdoS185+NXtuzZP5EWALU
pxmPAvP0NxwE/BIfK5ofTaEsx3puIyrw7XjSkwjzQPUua/rarNwcsQiB03CLaNSK
ptdtwNPViuNJ97aYdRNZmi0LuJ1StVu9FGuHG2hQrM1500dxhPZsFHBPvZJ+YLr1
JFLZ63Bewtb1V4Ouvr3WQ3BNWWutnIWOqZD4BOAgzRjEUQVI9hLU6oq3kqsZ3CCt
GdmxjJ2UprEwCr307j/hY8O1g2DQ1h6VzvfScvlgChPYHORetSRYaG/DMdooG/ol
t3Yv0ksnLdF8TGVzEzjD/Xu+mRroTAsw7ql+Yn8QnSZI6+bUK/yKMhS3q3zIqzYg
lhAMeD0GBnUkVwcal/51TzZ3n/golD7KViAtobO4HjaEN+JWWtzhOHjUlZMg1Sho
ZxrEuJ09GJST1iggXDkX5w8uGFzjPLJMqgwikXh23AamKu0q1sQh/YHZtRUp2PZW
aAom+hMYLxeBq+OA5x8rD06Gcv18c3ufQf77GvrnQEhTcd+Yrge5jPZ1kid4vzr3
+ShGRCzweEiiNV8kHBiguYgHKXDwmQRRdSS4UXs0x1bcEgU5t5X57CJ2iru3Nsdp
jtEikzZ53nn3JHP84VcX/ru5QSExE+YZ0JezBi0GqlkXgrgnk/FGasQ4JkzkaG1n
cy/4RBxrXc9e/e4ezGNPa6ZzFuvnxxBrnzyq089GhkxA0HvYY0PMSGjkvY5xkVro
8GRgWTMTDvlNw9e8v5jpY2SKhrCeyHPX2GaU93TUVmbAycflk/2O7rso5kX/fFqP
iszyiRtNk3PO+NjJJRd8Fac+Rozw03Ft2ZXvVgtuR8WYqj31OstwgCkELRWPvMLe
NfC7LPpwNkylFrY7NxN0scLw6XSF+bvdALTSTMf3GSZJmLujVO4gKGiH1XvAxYiW
/FmqIuUQx/JFzhL9HlqdegZCem2D41EEZlT2Ivm/2FORr0nt3gA9DcE/CNQJVBVd
TwzM4EVnlyBBiI9bIITsNlwpYtkJHd9wYdue4AoCBQgFPUxmd/4ptV3kleJ6TGll
oAMch8EgEEFFeUYeeb1HcYaxIXRXNF855jaFtLf8pEDFH0iSH6FuE3vXPgcuTzEo
tJUtpglNo324H1oA4JuasZTc/O+q3zQQhh41/G8mOITatd+I9poJd+yAce8iRHrE
s9snki2QIVk++XdGfqeCoHmE+TK8Gnu3xtwmahgrIUxArTZKLg11JwyNssx0a1cY
ktXG5u2TdiPHR+zTl21SoeQG5A4nhxrJRYVenitQ5TmZp9u5K+JjTGABM9orHv3/
GLbYfHpnALOGORdJugUu3zg8+fUbDq24XWwzAMQMIn9+/czKI78RSFHjVcCa9NhJ
IFpgnQrTJkcEhXGfmVPYZwLTdd4CYqYD0AXVi8Q7b5QlOL0EqBIC71HCPMJ8gLNB
6JYuXrtOV9jWCwOzUFY1P1qYudbcvSk2P9k2izsp6wqQb+62gEha0+YTjVVwpg7S
eMJtQQqp9XqTIbZnykJpVJZ321hC5psYAlcr3+k1XODD6iE0F4pEBKdDCXFZDPqh
IMfyWYA8aY2tmhIhZbs+T/M8R1J/q5vCPLUyC4UAKEkQGliotQrpm11oG04pnY+0
koBB6kYM2gIlnrRb1HsiCN0EWg3tzESbYnpHHjAO4/j7czgigVL2Toq6XHlUQOtu
A9yibDb0u0J4axOwQnmsHD2BvFlT5uWfnPG/rmD/IrxMngBbEbLxSE+ubYs/WhyO
vp7oH2VILEF45QjbrRCsH4hgaLYe8K1ocAqyLyCZRqFi6VcLZ2nDNVa2Y2K6tEbU
li/8A+JegT4rc+OAlmviBXRgWQYjgV2Q3pfVSu70ueS14xr8JOSnk7+HexRWn2eJ
5dGjuJpzzjQ996OjiJYAdf8vbrlyE0LK8FpaMEyXxAsqNDu6Xwu6XBdYBRJWFeHW
EFFUYZ/OBn2XHFcdIaQsovpNZweBcyyyeZPzqWDx8nXu7iduycsdDJKEYGSvjsng
E+TwwWEfXVIwyAvopbgUkf3hkSX9bROp/SYVWbqrvAT/c+0wezkU15mGJDWVPd1w
vSrT9E5YUV8eNnNshgzgpXWBrn2k9Hxw8klN+2GW2paxCssM/0zh1BmEjT/oLZQ7
3xaP4NGso6yG7cnmm6EpZEVzkQrKvBGnZRPGUmZYb2O5HVROgjmJN4LVB4FJUrr3
T83lJDYpwrP+/zQIDvJrs5fpFTuqywJOa1Fe1I30RS23r1plwcVZ6dqSJDUh8+Jg
rIVtFgup1VHMl5Opg6Nq4/hFutUYOg4XxUfz7ifNhJjBBqxIDA7ghyZ/YltNh3x5
1Ot7wxWPAlxRLl/js/eghmLpf9FDZfiFg/o73vsQH+Fw3YrwYt1BPIWULRduC0w+
DYJOHLxbyjqy+zdC3Z1nWKMf2JGdNCf6EfV5LB4IVUolz89paCL/uHzw44tIk8FT
A9u4YJJYvC+yrL5+5/xoNHBouRLfP+Ourx3ZTjaGDqSATg9EUzLWpygJgH36wJBV
0vKXO01X0oe00EYlSVHc/8UKr2ep3y/7pc0rS8d5uMcfGUdas+21p37fJlUws8vW
EvhH/mG+EeoUmN8IE0gP2WtU4xQF/PX8mybMJchXnpYBNeI6V2Vzr1TOAJVhICGN
ggeemNsCWFKvRbX6x1Bp1c8KibpHHBR07RatsFkTSzhKabMOPQwoI7Oxcf8upnp/
BnBVRBCRLTlGG/iKqRwtSf3aAr8+8HShun0B8MuQ15CvLkWo/T2qfpu/TZEiB2e0
CmByQfPyBM2keywz5ljQCylUoSTyiyKVs+qTt3FOEy2bSN2g5zKgjKeuM/9IEpQb
dxbTLyqo+IPbb9ddLZkJV1011K4bbFFDAGiSj78std6Yfpj0B5VveBfhVo3FF13h
OCaGDxsOwgYulqbm+CzpH0kOJrKz8m8x1gui6xuPxYfYF4G0Qq/6Bpp1ED2e1uvA
CWQYJykp7gDA8CNdD98ZWYmSfazDUXXKmdORbQ+AlT3ayAPw/fFZRt8hBn9Nj3Up
UMgZLmshvVvzoH3uwFGfEfc0vrmny7gsTepTr8IHXWO0JW2O+pMmefgs1KML7U5z
s7GVnA7g2lzExxb6XUHUzUFrzLQtIFZ2nB1NAxOgsCLAd1wVfifhRFF8u7CxjAAs
YPmog3G9TiWqSpjg2w2KL2rbXxZCFI8X5thtSIZm2fM/0VMMxDKXWbdkXTd30NZL
dHluzZZF0Stjm1Tz+fo4O/wfNCb8e196JQTAxuCXLTDS4AwSVFfpEfns4AnCnP2K
SlDvh/bq3hTAiYPGjl2j3bNttXQMxbJkJ8Cf1XYLo3cUJ4Ms0Z1qMagXy3ZL7qL/
/imZoberQFIVRXN1JLvlYc4357sotzZ5Cr4tjtSYQ2vJeshCVma7XCe1qCH304Rj
HJMz5t5mAW6sk3rdWp8uM5/lpOGh+HCJechQvD63bkIKeEIEUfVfKgIyfnrxoSyl
yPO4kHeDhFTdwDlHIa0bNZJEVNBLo7G+2BOu179jNpPl7433mklMalsDMrkfaWqb
ct8lDcKq41Ijf6tniBGGy/r+7idAvVs/hdDFXAjTGIf+uin/PS5hpfiEiavtmOwW
yIMnt3tGeTuJGtNu2d73m1Kx2AQEHqbBy4+5OQ9Sqxc624sexX4lBcqj4K6ktVUp
P/aYxxmezpPqUTxSZ2CT9uSfj36xerRkScTlozYt84Q5/akVh/IobCFXwhaaOyvZ
ecuh505IVwusyalhCZS8OW2FAkX8WLQYkoduhZwl+xBXnWgUkflycmQRUdHuksnM
Crx9rNRPFNPuGnydH+VlBu5U7SuCCfOKb5uSd3Y3L5ek4Dt4hU+1wRryGfpH50aJ
3GMznlPxxYYcKWiu371rJSKFdrFjNiq/r/qmLadF7dB70phEW7AXh7S70+Q/EocH
xHATEjKPDJwwCc+Hnc3ESDTDlrY8gIM7Qqicc8EZk+qyH6WH/2IOJ+FATc4Jp0wc
OU2iGuO/uZmowGTb9KT2uC6/hy2wg9gVB1kI87CwgfFFhPoC7ZgQw960zrNITllr
p2nsbPkDpBC0r6lu2VGbnyveAXqTXYgIo4QBmaq30NYpRQqsTAq2CuV7rvSARDNl
a35OKBUtglbGiNnRP5JWZ7Y8Me4F4qqphOTuykulS9+i5Ap0rGW8qa28nldvUpPu
zYNAnV9M3m5NRbPbei+5l/0J0/TGV1IcgjoPk3q7rJ56oxUo2C4CVni3FZDgJGYq
y7Pe6emyo0vLAffzYT3zelHE2WZiD46ZIu4TjAPZCWYOa0p282CEjRe1bIVQ9t6w
yAqNfLLVCvHgySZQawaQpcZ/KMiVTYt3iYzAa6cSYI4puK0YOcnjbW+vStFm3OlQ
CQDMO3OSV7ywvaSqprtLpw7Q+ynZKEQ7araxY9aDiXaeEZry6scXaNwTayW/+pC/
/NlTTfM4toRFpT7L615a6zNHjP3GPdd2AJkoXFAqllrf1c9qVC24TquiF6mji9vh
Y3rzrpdAb3aJCL9NImDJZMbHlyLLy3jOI8p4SCqU4u2yWG2iT047cNoR1h1zGabL
1RxIPu+Z4OkvblPyHyBaNKsSZPEkWwyumBl42AAp0Uu/KeG5d7tt8ikNR4Q9KtbS
TDTc2tBFKl7HtsLwrg/Vqbe/iSydEfd1ejIHgZjCy+PXvTU38HHMj2AAjDGH8h1t
We3Lfsv6Oh+VllFrNTTOT0zscsH7vv8tnsJ5O2O5sjWhQpcLPPZIaX1SJai1TrMr
EUzhwqEB9jcH/aPrmNAVnbtK7MZkXlvjuxnc+1jr4kIkoNpUMNV5wteaUGc+dD0X
L313wml+PWtNK4TvYwD5jYp2KuOR6tKDtanNQFxYgO3qKcmubb3u4EP8G3QaA3wQ
K23OsEueIXszy9jJ/R5SwwD7IWrXXggpvy3dBo5h9dm2Pd1HcbFDZ4VBI8VhJh5K
VVlkNdD8Pi6tBkDFx9TzWT7C3qx3caWSeLQERper6Hw0E1PnBLskRCXFLKc1/eTT
j8XpAnfvkxE6t9cspbLGaDojaSXj6CMmFHDF57q4fBJBJZMRhKcEkZBDWyQbApva
V7mTgW5jL57D3TPzNFGPMAc/mpOog7m2CS88oDFVpqddH8dP+Z/WvXZSbon6XMmv
pbUuRQph4YJncI4O831wOhAiPy3G0q752O4hiaToyjY/1uZXAIrT55v6YgYgEdcn
UdCHh7r+I0ehwAwdv9aSNG/IsMfa1EuRjzdOigof8zaCTVP1stsqLMa8wgsAGGaB
lpXOR5IWh8OVjFLMt64nzzFXJybfrsrmGLVeDLYCXossbf9yGYS6RLRmeVYt4itF
P3g+dIgVHoIYNyaCIjfNZQsNzXkTkeZU6gw8RfUesW69UShQ1cfKzth55TA630av
G9o8LVTUfHIslb14b97Pm0NLdDP0HRE14ye0jjc8d+v6TUPgJwLfTOYECKs/u27V
6oHYH0Lv0bUcpZ7u3mKY52mWu9FinRVKxq4syPVOSjFdpJn8tW/TVr7zLtdRv0m4
MXbvK4FvmexXULowLMDXJ8NZRMf5DhkSMSrK8tkuV5F7XAibKlOA8XMHXGoB3RNS
lwxNqnOLBIsUII+M+MRQzV/57Kz7k9+8iuri0apU8rgskYPK1zUezEzonbzznwx1
LabBS16ouTyTgteWHur4Q0gQMcwDrZmWfkD2ZfThjK406WtGLtj/lN1BJeMu4Anu
Vr3ExYPtg0CvCymMY4rEdEaqbw7e2Xoh5OCo8mrab9X2HTLZx5D4XCveQ800j3Lp
XJEP5wdmJC6nHRpz8orn6s4z1mV9rl21jUeUAlDo1et69ZGvbbXGiieI9R4jkAQh
uLJxQmDs0yjxIThywBfxjm8VOIhFXHNnwF4dYcPsc01Hwe2+ie45TXcRMJugkeKU
lABDFwelLeq4IyCD3VKAp6eBS1s+3Wz1jEJO7iMPTeuspdv2aIxiTZWehljK1mU2
dsJFCZ4mwpN+clpIg4t65fqALmEqRUn09hRmlVdvtQrCZcRzPivDd1i4lVrigZFo
39EO9RgEFU4AjmlmyMnkQ0ePNaPIsCYlaAJq/vdaxc7Xg2n6Das7uwDcXISDLocu
a4sy+1lZmA1Kf3wtAbiD/OZUsc8lN5LrxWHeLhUVGR0ZlNWyGIi3gHBmdzdNQFaJ
CJdJL+DjIRFsI0RuPWUjLVPSjSlw//X+HcBuHlnPFj/mAI3pWBMH40T096qgA9QD
HSXkxB1MfPY3Og9zmQgEnMHcKYqsHfKJcgEo+l9obR9JAi3JKdfwClDN3165Trgf
HMWh3PupDz0M7imJPPCnIe95qQxZSjrn8BXX8pcBDJ+QFcyQmfSFst0sxKAkJ73a
dUNXRi51FWnQVrSJSTvVN9aZg9gFcjYIHbM7KDoplu9jTZ78s2xJK0QIIaclGCPe
TSqmW+pzW3SUucrdy8SVMZ/GOcqWGiV4YSVBithaIpvGd+oxDrcsvqdvkIhhyH6l
pxdkZAJsIgh8FMlR7Bun7l+JBYOwPN1qeFBDt/rXZwdwviKICWUNgTiRuP4uZc1G
mSOOh3cWb6oNk0ZqRPNyST6WXOJ/TurrKaCEoYEcEMFX1JL3lxDo3/+bDUqM+YZ/
IhlCR9OC0zYYqjfl5mzAWEaFdHCctzi7lKEKXnB/0W8yy5UcmI8A1sE5fI6mJ8cM
Ld5PZ7yCpqtHEJhaNCAc4Xrm8bnGTcI6QJc9l1mw9Lj1Tl8ukq3DTsqmpUmijfZw
0X3H8MARY2rfY5vAi6zC5Y+0+oQCxjOcdUvaM0n8GKyTTWHu2TJYOgPzOj0OCwWY
ca7dx7opFKxRRK2/0ChOYzKhBUvaDSYXdncpsJfFp36TcltheoTeFLVws1IWTNVI
EfZtV1KL84gfnQsiz0D/zVRdHy59NfIAndyrpTqTnF6VutlGXEZdnxljvlicIYsc
c6nROFC85ZtiL/Lbn+B0AJ/irFO3t1C4EsSdQ6vMjfQjqjdcNqRZIkeu8vOcKgCA
kU2Aco+lZqiLj41sotGneDU9kTD8fpYlo2ihYEep3cIy6fM78MYSM/v6w3WmDEj3
rJS/PN4k3N5DBu5tp6VEH1lLcS5JNZrhS698Lv/mi1s0uCwKytACTxQoEDQ2fQ94
+AVQvcqaYuZ4XQqUVgZUfb4jUQVn+ERCFNzOZGpIjEE1PYWbW+il+xRRExFs+wN6
RXjIl44XU3MgAhwhVkhkYzKAHH2kuE4adYK8FP3z4PZJQQkkAQLfWZ8Uv4vRimLq
0zn34hWEP+qQLISyAKon/3FqXd9sO+cy/2LS6RB/9ruH/U4/05X1YPybQLPn1QiS
9s4I5OtDVMc9hrdmMeP+XW9PN+2p/zZYWz91pToZIj0mOp9FeDcrISwVL1m76bdH
WFFrnG3xb8jROMs3snzJP7ZTIqAEJJOwLD+lsp4tK4he4s3XqMCdVPsADtH0/NOU
ZOmBU4JfudZfLs/zZfp8Vk2B5PXMF7n2Qg+S6EJrkqk1FUQJehX/h7/oGZ6nqrqb
lI2MPQSjgC2LGARtTe0ExDp42IaBjqmDPyXO7xh/prBFel44ukiTi+Zpvl25YLfQ
7geiwW83IC13/ovESaTBU5R7d8xtEAcpBSUMkWWKsKSk3dZ3xC1lagsS5toT+UbO
rtO8tx9At6tcc9stJagk1Y4KHhHJysMVXJEQT3t0gQ6SZrVnLyZgRRPdU6vV7RyX
UfmC2/cijKQSWwrfSTwyXlaqaHFecDvXyShPYo/QnoGuNvtQT8L6U0DF7Av8bghg
fDi8zfx9NeVlxeXPA7c9Jt+JcJL8QoOB/SqBtGKObIKgUgC2iBYDTgh+SKA+ZLLw
wj+2z7pneMHbMPaaH8tvcYZkqtQ2rU0oYsZE1JpMnWKC5b9aPXAiq5ZSHgaD+Run
CqH5fXS/ANB5GHraEMzB8oshZU4HGEPdmDsN+PR+C3I+jemdMBgWokfxF5bdeUor
iIopEZpEaUkBAnBJWN69sV0/mXnY6eAjSi0c+It7HCDKYTsWnDpNrhrRBKJL6YLo
uBR473CTlKpDhbvb2pe+yEQD4lUr4l/ga7Be7cfLVnRUMtwMw2VeFLBpfz5E1Sgg
2pwAlmrmfmpwSpt9czJH4pSaY/z8rYccWdYdUrVZVA/7neXBRaH56wnprgY8JzZb
g6gPmYsEp9ntm4FM+rvAOqI/E/Bzu73DqL4GOCfbxvqFouJ/GnsRVfPLFqzZAV9q
B8U0+0j7JflST54apxd0Z3o8nbjIaSllsIYDIwgVA7B58MfObCVl7eKUT0mdCm+/
a3SEtcbDT/h5+WLi1CSM5XLzdiondLNhPiPvUHdhGd4SPBmdWCAHFiBSLmN464yZ
eypBCIsX0euOeo3U6XkmwUZjkllyu+QLPrIDMYeRoAPiuYJ1IuXtx0OJT1YmL+dx
LZgp9yT1zUrJrxwk2VGu3V/wyrsBBORzJw5UiMlL2/NlftsvFlM2aPls4kSAHY5p
Ck3cKwhcnEDi2l7WHZ4+tIId7MbPPLQCEexCoZ6kT8RadXaUpZYHMqZ/SvT5SneX
q4vEakrbTyMKIxr0IQzOgisJccMklIGICY/4NIsoZVXog+/I4U8sxeyIQrnIYg1q
lSLpWLPYXsfYAi/t6SfMx1l+u43eqF7pPSiIhJPIQxkJ3LrZbx6Q7l00UFQXysWG
Oj6mx7CFtrV0IHWZp7xzWMqOlHBm3OOxjGQxbk3+IPnJLPuTVdG7GyTNH2fyr9mr
yDwk3mb4cCUMUk9n/hFzQ7AXwb7n66GaqdxjFA2wUFcG4VmYuk7aqwdCcXKnbHs1
Kc3Z7EKE9NGfdi8XVmBZLy9xvYqOIwKMkIsbryzJ6/G+CKFvqbS6yiUuMWmIsLIe
8r616Zijzc6QeaMK73tRAaeNAcY5V5LZhFxvC1Pt9c4Uq+Qn844jPQMO/3tvECDa
D5ckOqvlVaGFl1z9UVwKkQ43Jgu5mI5jqfM0W+SYR18=
`protect END_PROTECTED
