`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2Z3CQCdm5/ifIDLExMznxSVSfwoB6Goq3M1ZNw6DhtCN5R5IpRh3R2I6tFEHvkU
B2MGEbScTwSsDlieNv5An70HohtamJcW94Yg/E0JsBmeFs2uJIR0kAoprEqbzRKK
YTbYL1cwNtc/4VNTAV/nsejZmlcpALcwud+ORIb6XwLRm29rkrPXUR5cUltwvcB9
R1JVPw2HWai3p3MPVg6PDay8mTTf1s46dEVdT324V1+3gLbU2k6MWQL55Dg4F7R4
IQEhm7KSOUcFzb6I53/KDsGBn3EFc4NxMvl+Gu8q9Esi2QRsN7/BspUx7HqYABo4
t6SJHDzVXSVmDnEzYt8uD22N2TRaPmIYBJr2Za0t9Z5e8ZMoQhg1jl6dG30AeJwt
HOmUJbZtFcrEUoxmYxWJMf0aixwQ+XcWcYxMaUIgoh30wDVtss66lPvifzrz+f0j
I5E32kG0KiYbgOs/zF2KrH5a7AEZHbdy82xIbEyjx6BR5jJh37PkcK00JRqdcTx5
t0LriTbbJAyjZmpvxH9vfyKU3S+r96o/ZJz/GVQODDiyqr1nREll3+S7gibkNF1h
2nI8wJqyqFK6jQbQ6l8Twn7Ijg33aIkITPRQ/UmPj2Fnr6QGx4iWEtqTuSzkZw37
oYpnzcKqBxNcX8LG/qc2/ACjO4kiuIG8EXnJCIwSItmevdS/rS2sMIvZxTFR5wTq
Yyj+snqMJzY9F5fKnMsI6Ma9ZIWo0bac2Pm0+dieqjypSrbCcUve2LZswWH06cXi
G3dX3p1StHawt9tjUxwLg+xZl/ulkLY4rC8y47jABbBwVv1hg3SdysjMKqeJUJBs
VF3kfxV+5NiQiwSpWOhTTgfTd37jubA7odk4KJIUm56IZlkYp2jCsEiGlnPpOfBx
rGPQkV5+AhnkYMJvNlZ3sw==
`protect END_PROTECTED
