`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Hyghgzxda1JNN82nPiM2F81LT+HaGdqqWf1XKuTZKhAmhPzQnPrBqg9za+jUG4n
suRV4VJ4ZCzrcJ+CONKvQZWOxXYHQI7BCqmVJ1wHrWVfeDKu+6w/7lui1dpmVIpO
gy4cihxTUTfsEU8950vRI9ySL8/TsjmZ1qqSH4XAb5Tav/5cAM8Xthnf50MrZMFF
1Lo7m3IxsEGTgNfpMoOmFJTb8HT47EUZCMOfRXtkH1RXy35MqO539Za9kaygmtM/
jsfbGnq9OOtc9pML0qdEB9qyRYcufIxpA2dM3Kpf0lCsEg9xeFQ7ue1rL2q0nvic
v6I0nEGPhZ6RXAzsUFEfdw==
`protect END_PROTECTED
