`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
taSRbu3ewRVDlehWYpYJ6LpSglmA+2Lbg6RNmaI0Csh1q51fSHtzVJILt+6MgAvh
bSuO3X6TUBUfSr9n39RmbnKC+c/+XsGNACm85F+AzfoCN7q1tnCXih9KDE4/EPEG
jTyps0OtsKlPgXzIT5sDiX75uy/ka8S1wbii0d95CTK6eZhVUwKrD651d15S1c6D
LS+QHDfxEOc9+jPQHN+GPA7MC8+Ok9iJJ9cJ957KABOxhjHa+sPIkKLCcnuzQFsv
F8NLDaFhLNcSezqYYmKsK2YcHneoIP60FGzVDAo/EgnYgM3zFfAXbLRqoiaMOXV7
QICB4Bxl6g7bl95wSigAIwCjkF9jhwTg3uAkqjXE8FvSST8HIIatmlroLx6P4Xis
8F/78pH2TMXecfrw4eslXMOCaTBMXXh9ySkYJp+dUwWoEE4hksmMuvCuABrl9lpL
s6bKy4CWDGOY7gUqfMj7zU+FihJQ+G2cKVVU74BaaUDavb0qhx8BAUQM0iVEWIBn
jjVWqN95U6b4TII3mnFyIlQgFH7jkR0Y4uzUwSje8YTr4PZg33jcPC50KWZ+qhcJ
Bl8ktHo88BfcXLmnqDQ8hsqifFUOH4OXJtvT5YhSD77Fj1j7CW92kgwJGvv69qZH
F/Eu07qL2YXROXrWkwcbdVsVzp0GbVQrFcSu1D2PQeapW9idCxPV/Oce0pE+w64c
JMQK2tFYU0qsz38BAPpNDQICdTEey3eoVkGADZzExNAoE8Ar3NVQxuWWdLQ5Ykky
fNYNaJ1RM2HRwY8CYptwDW7J5nAJGDszFPLaY8aiqn2dupQHAR3seMEuMb22mLYj
S6q9HUyHT+SUzm728pEuwdycK8UuF3K1d2ZjARUZ1ju73Gcp6gFAG5vDE2EIDJpL
w8iFvAbal8vIMMf9hBmKOmzbiN4iCAlFTVkQep1JIe/rmTMMF5TYrxPe8O7NRQt/
PxjpVVUDS7CA0mgj3xKGbFX8lhDLJ9cd+FemsLurtOLhWPnGmza/gpZGlQetVAyL
ibTDWkI82XkNe6eQRHu4m5y6rGZi3LPxzLnSeSGiGjHXMxbLy1xzlnQGD2lVx4ea
C1uxyM+mqOQkmfetgDPuXEDY8GLaCGpGgZYnkxhq0wOej3Doya3d0farC6BnVjXI
mJ8joo+97ldpDMTwGsgJoy6a4A4Les6aQ2vYgsVy8MToQOyjq2HM/DW2JPdGoF/R
y+Zukc9a8GgQt5OEUE0YPp9dMQLb+L6Yeg0qhFEmknIT14l1YLaFDpqhMbVwmHOT
v9DxKpOqicCq9gpcskCfr5d+3qdy4LaH6ES9PHh7ZPPsbkm6FvZatTm9Q13hbtCQ
81728tW1eAqSVX1SyF03D4npYwqM11r40lr/Z2TYPnG25h9k2n1tMDh3aladIVBW
r8E5p3VP56BQ2RClO/1Sfho+8k8Y/M+1doDOYBZrokToCCL8g5VgzRPwGo99+0eB
qUGZqGVUw3EXMRL0cnaelJ1XLvA6zUgbH/GDW5LkIV+CAtDPm14hluh0m74nkE7N
EJ8aF2ab4vLOMUsnnfm9fE3ULMDO1f0NbmseKstc746L4ZeNWwPxZhGw7Pq3kZEW
7Y8R5zeKaSCM1Tvh/y8PhA9iL2VvNfaN+rooOmpnKPWFL+hSZbHxcELEfjpFw94B
SvH2PVlDrk5cgvrqSG9VaSmSXo61u1WL3sgDZfu6W4QgDNqFppo6GMv3DmSoh52a
20LYjB6At615qKlJ0Hs6XHfretuIcrfctrbEUDartlZb1L+m0HrrsYcH3D+JtDd+
6/NkZvdBmtqL3PUlGolGatzUupryjs21h2dXIiI2jjz9dMuDwzSCbCHu14tGNlM7
FE6Tsc017arx9W8FtHmRpzh+/nGCIDYhHroVN7UDnQ5XYu3oX+OzqBsqBJUx/Dt+
TvYCpDBguPrSER7o1iz1698dzz1tAQZ1ll7AYq64ZrVV1t8spPpOew3MO9CXffgs
nUlsdbFSuVmzgSf5FeKFZBjghTlQgHlooWLr+UFSGHf3e3a8wsa1RqlxiAhyN4/s
fE478Xp+Jdrv91nyZyRUNHqdsS2sbZvFUJlT91zqKlKLZ1LgG8HTfHxSKYtF5laH
9TZUHRLwk7rS5crkXQ0rToufJzPMI4JPpqefykVK9BZkdSc+TPFH3r9WxNzRKHCt
eKLK0iy3gQW7J5KyeYDwiv391TpDlfFCOz5enQrV3/A4TNsmHKS5Tiy8d3XiUNC+
nfADkUhEucYsfvfnsAk8vmZ2tz60ZJIfO8RB8FnQ9f9c47ZIbuuFJw/mx1JPUTPv
e1hsHnsBbB3SFegWrd9fXJRSWxaCD0ansO9kSzra68cSrCDk/MptKvYv7nob9Onk
3VYFl633ghlKxnqH0n3k2gWHQRnfqL2RFDbqO2uRmB7dvCDl7gLE+ft9U4sQwNPm
U/4Riak2s7nDef1YmAv9dCB1VBGhXRqkTEt91cHfMs3QXPW0XLGJ94LCufzYdNK0
AvidjFAA6dsJDAVVak1U1Bc7ntzpic4ymI8fTfZHqRtouBUcIQi2nv06dZ1DszyX
Ci1C84WXjDOrcd41YcKkzBb6mBr0Te5iGtz9UgJocC3OuVhKq1mPqknRB7EszXkZ
z498T7+XKap+P/7ikP0SpZq19JrbAb+kaKalskNZ0XE5ThECMPssZgkVL/fS1SDj
qB3tPKZhymeLQ3tlmSZUN1R3JhQ9ONZjJw/pda4ut7lMQmutWQH8nzgHy+0wBv+X
fHn/TyBSUGPxJOdYcFa+j11m0M3rQW71IfLh91ocVlJr7Fu+DmQDQ1nfGy2uymKf
pRz4hgzNpGr6VcUVEJTeNDRKI8XedhD1dSvIeNDBHb67L/d4/ytVS80EHQbRuzMP
K7W7fxUaM+SjVhV7wkvt8y7ve/eqQ43mjLdNPovsdpWGJgS4jxtYfrrZAt/o04i7
2f5A3r9O4di00YE2mp3wfTsAmpPvgYRbTjV/25f4I6jGr5tsXD8IUWeOfy7wz8Vw
2JOFSlmdeJjVF2E/wTjo3LHGDYsYenhaGx0qgjl78C7LV4YUEtMTcTo2U+J9jPAS
9dU4c38OGgmLGNwhbgBB8nYIuT1/CcLGHWOv5tbfsVCWNSWRttewAYfsZynVUtPW
AMOVof5DvrPK2vUfmf2bIPFJQcdLLd5ZX0bxBCDH8xdkeeZZnPifMsdE16Cdsu57
p0jaiTd+SpV/NJkcuZua6wooPU+RxPG1hBUDYQrYOo7gPtEfZKkgXT0uWSDICsbG
t2JzovvoNu1EQaj0kMrSU/NvkSiK6otTSP+YQ2WerrOyeuJCenHYQ51tusweXMB7
Qn82cymaEAmz7xNETOxTZnfArHtDxqy/YLaLXF1EOf0cFx+Mt16Jv6hlGLwp+8At
BOMWfWcsT7DFCssDSKSrjnrOaAoFcVJLeRK1aeLiBAUC6ABy882qRip8JSLwKL8e
QLgH98DNBvzri7wqIVP6Lo6wHbaWsjmHXJFgBIgctOE792yNJLLTILhohF86CjVF
v6g/rFd7JorJUDpO+htYUmDjc0wR4dya7tuKH/RCTyZKaBrgrGTlA87cMNE0DRlB
JbW08+0ONQKBkydQpp2abBaqmni9JCdDu6BurXF+r8qKJhkFyV5jtFGbilZEMDLp
/lPb+VFT/3/wI7YgnpT6qqHK6LSPEBEsZMRJFLJCGBylevaC/WQLdgqlvflusYm/
j+3nzj0zGyd+Tn6zZuHCtoX/Ih/n7w5rDt3OjET04TuaQDKCSCdCLpAnPn++wlhv
EDZyRjef31abvDkLZ+aaSsIzrl5AnhOk3S0yJN2YOVQbpk52Kx5bhzJAK/aBqEME
FtRgaIL9CsFrMWgQaTmq0x+135kaLBXKdjEOn8SASCj21siTSLjW9Nd/QXgcwWm5
aqj8xG619kALysH4zDzKtgdGrB+LaHL4Uo3w8UatfhDYXDWP6dFTSvXToVk5iFFm
+EFVe5TLhYcRS72DmGGuH+SHOA88vGs7Gr7NsOTuTvHcMGYv24/EFgkaU7QYhUp4
3+ktX4tVvb/otIvi6GL1qK8izLwZpP572sb2/lMTRHIl1yjZrK4FuM2B2D7klHbS
BMQfCDenJTM+vTpMEn5BNyyW+Z+Y7s13B425i/rJXP7xV7xY0Yq90itDFT1up+Fy
ktSloULDIZqtnejFURtDZtHo0N9Bv19sgnMHPTZX7xNhSJc39manUJwIeulNju/c
oSNGFEdzhuVvpXGaRcQl5aHSnstUdzeqhgG/KVKcll2+GI/VTjXwmr+PxVOLdhVJ
74RC8tA9jk+TxCgfDKHgf8H1foh0RXMKGQSybVzv/+gfXSGUFYBTOutK9iOjoYZw
Kx9lJLqcnjLD0zrwIhpj/pi2w2vXx1pjWfr/SOOfTMMpjnc4pv2hFQ2kUms6EnOO
niMSDqSwi8HLN0r6vgK/XeAmrJr387mkzj0sAK7YVqJ6QYvAixqBgWpiLsjJW7Sc
nppltL4Toa27V2+Y4VgFw3kCQooqcarRbexel4Fc8CdwHv6AjXJ8QMgBgDOVWhso
tAIBVHYndd/z0iyM0Irunf2GwDpLB+Gl5cSckSgWqHi4VvcX/WZ0wQBOk9sJCNwA
SCY7pnpZh3PdpLlUMNxQJMqCc5HTp6CD3CFHkwLix/LAUFlbfRL4HtTTgUAeKRnx
nhXeI+Nkdc059WMXOBpABbLt3mpVY8FTtXjnEYIZ24eyp9OHcobAThOY4eAsRq0J
8ItvRW/D+5eRqh0x8fTx8K7KCBBZOs5Ms0bQ5ZCgIOE=
`protect END_PROTECTED
