`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KcH7GPV21a9PYqnm08kPSl3Hx04CktcAS5ssPKh0f+PjQJoyAtKVxDQs5Od8Z6aG
0+fe1GbHlBqSjLnGLptYs9ToBZIcVkR5lCRR8LwRxElbQFsAHNHopy+y8FBrHocK
PpHtR70VYDoPUympy3GHqPZeMPM+I6VDkPWrIUw0A3zIJM3QHbfhkFTejAPSCG8c
NQajGcUQYDn2IwMRGlLwNIwLm+EkZ8jiN2CXu7Ue6dxd9CV1+Pwh/VFvMzmGYgXe
h4RaAKdgQ41PB0sA8Zfmznb4ZEcUwTRdRMdffyDDQFMUa4gKqVaD/pEFfSS2dUtr
SMS5eVq0B9sC0B7CLwX7cnFTmmHbAEWwpwTxmmAYHyIgWTE03VfBhmRqbsn68oB5
uRC4ajMTF2fSdPulOQ2WHvlOB6VSnfBMfKgM02OVa6MJL5yJfkvFyYWwZV0+Ue0U
yEVb1v6+HvtkkADx4ra+wKOE8J7KawlqnLFmDMPg8Zw7aEyxawbDNc5alHqE6s4Q
bbxXbjcaCoMPo/jddclWbHWaKY5vj259WY2UKdlaUtcWIs8tXJaTrDMky27mLuWE
qdE9BMF4hDndU/m1kRxzpi0xpo+hEpv0zjYtDVfXoXl+maLYjDf/Fru/Iy68BDy4
evsgdPNs5/3H+SdB49wfFefX0rvvDLGfWEP1VmuClVaxvT45ov0Z9/aiKfBuFUkz
31hGyBgrEhAyVLOCAmDGJ40cMhf0vtCK5rHQTAWvlReKQwxB6ClH9WQBbyNZfW97
Tt1gh0ECN8ROKd86g+byobWxCJxt8vgrE2aMxOTQBYcPUWnlwbo2kBWWsvphlSpT
7x8b/83gWkl3LZivoQTHIXrzVjy0N29VL7EfoGQZS77vfUpw9npICD5NlhC9vsjP
ksPZb+31QrJWfl5vClOrMcXhXIUEm411bezKLmEJXO3vKxLGrv6vnrLc4VaBROXH
G8fp/6AOH+wijk09MjoCpUNMHocioQBWY8lgOhVkw0HOp3M695jPqqwSiV6UEoIn
McjWW/vIl7pIm9UCSHNqzXflZhe4aP6r/+yhkeP0wk6HsBEywW4iK/daN64mIGmP
87i5sN2wKmspaFQWRB65NmnFJpq5JeKefmgmC4hrB9DHNfVualT7SNOwlbQZ7Xe1
7QZRak3ae0fw5DUHQtGMrvRsrbKMcJJ2ZBk46nzgVrLwMXchfzRijNzV/XqiGmPu
RJhVaMC9406wDea4gKAuZpxeIukLZbI7tL5RJPjHrylQsQWV7pxvI4wu/YpZIsjS
EigXpsdHFIynG5dsDEH9buuT1mXM2Nl5gPFZNTqQSBUdCXl+4hIjCO64XjlkFUv8
ne+B/VjRmZwJs+yZIqIyIWr85AERqxPxbus86+z9DgNjetFSAhtBVhKBKS9/t4h4
QTCSZbtSUwi9Vuz33K7K5g/DiRmqn26EEsndcVUiBzCXnaboSJ28DbgZlsrNG85z
ERAEPIrmDH1gXIUWmEz8RiPxGQusoi92kex4x1wRIgD5PXKKzvkff/6IFtZbBdx7
EdXT0QWW1zx2iLeve9pl2adIJGxtJ0Q/90+frZd9wPmL6u9CdkYxLxPjepyIhuzy
sG90cUHCodlX76cr8q1Qp0di+MUr3S6BwKI2YEnBed2u8+d13nTCJdMxzDInCjcR
VGZbZ5ZUbmE1md4zL4ZqZJMY/Msv3bRjuB6FLSRWSsgwFpYmAhWYBlFSFblQD6Wc
1WdggiF3ayloTAj/ec9c9chSyKT0ayl/4Z+8dCZn1wr/FE1flX5jrsghcGHB3oDo
k+7APIhQ6E6QlI+eqCt6ofAwTUyt2NoxD7RSV6ZQWhSoUIzZWm4q6AUNhscAi6Qf
rRBmPlYd8wLD0SKMm++z7RhlwllpDSoz3ELKfVxyLZ6WOzTgNMcpzzpilsvQRmeu
JyDL0fV/473noGW0r5Awky1b6XAFbLq4vmOvYc7slu9ulmwf41XiYT1llqXa5fA5
2i98CKZuRaBkzjjZJZqaMtkwd9IRwTk5kV+Hk8a0Ic9ihCJpnsWmilkDLpDyUCJT
W8yXsLh0AWTk931oPeekcpuFBfkkztnXhbuIbKtZ+FwEH3sj6Fw31JUgq72dkX+6
P5mFHtw3rD/eJVZLUDWAF9Wqo4qIK3khi3lC0AW9virsL6SjnDjEed4PgS8+5gaY
FTK8DuwuIrERCFuooAgzolcb18obnRrp6tbrGtdQCNQ1sojIGaDvg9hX5j1ZeO3D
y7CSyVyr3bV9MpcejOVFJfpwGlwP1SF//e6IUvR9J0xJhomafesOHHqT2F5VTMkp
bD6MGE00RD8qTCNMJDigzYaSfuGBYPphc85v2ehDsrRuNznePerEY8Rm6UMi9Skt
V2nf/640tWbyUfpRdeEkG5aClnAHBw9kZ/lMWtCyMLBZYpwit8yzH2YZRbr+g0eN
bYlk57gwjamkk8NB800++JN8TUh/Kgl9KhwrHgSL6rAqhGkjKBGbnLobUisVxp+m
2CjOQT6gII3tA5HgYE5rtNCp0y2H5jZg+Nlnxdl9nujXwPYosG4NsL/Mte9LjF7v
xmA03qU7J4DjcCLdeCZC0/BEcc0kF+kPArqJBz5bLFWva7YFXY/8NtylQ1uHxHA2
0qBiBiEUGDIlIAgAIo+ICvW1AXxGkQPDl0NYbrymD+GtNscya5plKEa9n4gdmF0X
4NuTg1tIf18ThWk5ZY6YB1GuAYL+F5YPARjNqaDju7NYFSjGqgkJyrWgbD0cWqce
ljRwJj00Lf00NCqfYRdLR90DFIvR5w2IEHvTKfGoEQPS7c/QG6jMjP1uGrXJWfH/
qmPWsiGCBkmgqnmCPWcZXdW25frM6Qz1dBa7H7eAtNuUWhXQ9tL2dhYY+OivpA2s
tSDBGkkm4hd+eKdL6aJIo3OkmMbqSmUhx1RW3P0QIC47gAiXoc7SD1P5mQJ85hSw
8n5FB1v21SeJphv8Fr3xSReG0D1FMwOXeIodFrvGLCrW9l6HNPqCvQOayB4TAotT
qrOFvBFl9FB/xvrAq5u8fWdHYciKQhuke8laOHR1Jk8NHPLTCTKmxB/jUzN262ti
rGKrkfXqgEYbUmFBzBOhZ0JZ/eqqhJTfbLWnca4XFJEDHq4B72xTYd1Z/DdxqneO
m+2eKY3SNrBJGYBZX8K3+LtTdrshrcQibVMRqZ/wasQAHaw5z47YVZsm8UKHmyei
Jwf2ffBcCZYdfapXAK3B5tVZpPNrjFDX6C/C1cKrjt1XT0WjQ339F2D0FxlsTUFZ
Eoet6C3hlrUCegOOVTdsfC5tzXbwXitk+e3C7hW42tOSFheIAgrKyuihxpma5QZX
s02buTbZhbR6NrgmvOUPtuePlZ6ijHI8MVzvLScCwZyNMRQPUBjGl0mp/o8YYKX9
Hs4/EInAopGVtj2f+tzBe0zMQAvPm2vU7z89NDvwVp0peCaJy3SlK9c++cU6ecPg
3ZjJ/xs25RQE4Dr4lsQtFr4NWZvRUbuXESQ+Unv9MRIXw2kceQ3tjJrzEy0tzjBH
HlRizN0Ps2uoeMor/HzpeOGodcKUZcdPqdfz+zrokUFcsEgPhza7vK9wb/yrN1PV
vy4xFzKcwYmh5y6Jc5qutmoX3JYUcsOhW0ellddUmow7ONgyscLWqSpaUxdYJ9w1
N67q/6lufUMrN6WIVweZgiMNBnjtfwq+qxpK9dOAWAKNHrz9YFJz+6Lv4lP8jQrq
x/eZsvLyH58P9tjX44aloKZ0YeDcX3Kz8JLZwrzsnHxi8P8QVoiSSJyl6j2qKOiV
OaGnA4i9EnFV7dB2QxZrS7HYET3PtK3ZbC3Y03EkiMJKyIrzy17T8vBC0Ow1F8CC
SCGItSQG8vuGr+YF5evDoQTCuILG+6hNed8fvadD6zalelx8kTjOQTQu0LOLNzGR
HYNjD6Vo/wNAWyxjzm3b3oFeoClzDq1/+sBhET0Wrt39VgkgEaiGTU4FyAYBUseF
qEXq3dtCiuP6zuvR3grQ9KT/nlxd7i5MVbx8gtKD7Fk1XvxLbuOvau1z1NQrfKrE
XmTq0f6RzaP4OzVa7vv+1g==
`protect END_PROTECTED
