`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3YFvbILM44/rONr0IMdEvsAinl8xRIR4d8xPoO3zo5ROwhnaFhXgZbVjekzwW4Yy
qLdN727ZTEWdVrqueYNJw38xrfBxIBmQ1chky17D6df5zjun+tT5cRdiSYjOnwbF
W6qEzVmzi5ToHrsbzUqw4rm07JkMnoejD56aGcnsJ+Gi7757WfbMhNMWA7U+fM87
BAXQ736yIOXPy76wsw6ovdinzOYxFAQbrQYXi/tJYQbx1gpbg9pDZGzvZvOzhg8e
Sv2qapoyaGfzxNUEUO8qsry9K6JRHbtoOVzIaJKpvdB0snTCNgKzbLPxJ4KmkLaK
YAg0hM2I9pnvo92gzmDM8cI9o27+nWXjD7aucBNPvTgQqnxPs9+mQRw4JVvf2Pok
Xwc96LVz4S3GcuDGn2ypW1I+sOx/1QEvit3v/mIt357BH2Yi/kb9EgAhDG5vs+Yn
EB4ZY5jBmwxgCcUGqRvltva9x1/HFFYbGGMd7X+0YCfAL8Xn/ugS0Inj+TnqyPPF
LqlJ4P5DmyZL+BJ5NWf6HU6mgViUPBjtWyIGtjOzBxVN6oUr+duZObpwHLtx0M3P
ivpe6bCDFCUIB+SJFCk3I3Q098v/I6k+FKlfTFmpmP2ZbS457tCnQdDgK1yCkXRK
4I7hPB+ECNKzznuQ6Ii1iyxbq+BwtirhcmFufv3Sa+L3ESFA5p3A2jOzGAOFg9lR
j1sy7avHsSW7AArfE/bMJVljkX8k2bSzOJ6nKmhvBkGPHu7Ja8NTmLYY2ajdendL
PJDgnh+0QvCBr0c7G8yisCaF+PYmUo5qt8amXpvetD0EybIRhE0+QvsQbAAOk+E0
YUvBlSsJlY/vL40XirSKYVbehfvpVIvMmnlpX5ysd/k3xJsY4bhw4n8RHZ7zL3f+
BhRHVxV0B/lkbOyIDahLF4J9TBD8JroH+oCrv4cESoj+fnSvCPKs9PbMYNGAcksk
uLOblrrE566rp3t6TOvxZuVy7q7OypZnI5kgvu815w9ZJxyLJdRgH3U73Wy14zyP
WjEJoBULL9dXvM186oYA6MACi7waklcdimJSjmJ7ZKj4Ft80UD0Fwe8qc7kzvo6l
QdaBBD/w87U4UGgpkQLnPUmQwu8bN63Dn0ShN4erddwL8dsJM/CIJNYoMJtbca45
inaDb3YAogkpGpG+iL44uQAXQfux+gwvrUkQjXXev6tpN7apOzYbbkRW+mDI0d1l
se2+nSHrC0Sq+vBRmB/JWhbjln2VI6bsClnxZKlsuaHuKRd5OGu1qLYAGYlvpN+5
TTIkyRettmz5H8YqRqY4qUeqeGk9XmJPjCPNs0nAipR5mensn4/fABkVbCot0Z6r
UKJWPmrTvt3v2yY+C2ZvvZ22QLWiTr11PU9kkMuKR/msbwABF6yWx8JY5+cr90+5
aeaNYGzAjPWxzLuiVIaZ35o2ajSMxJs9Mz7sqD2/ELIdASONp/212hNtUgrI6WGg
ozQBmsebUe+yNdUxjKWaZ1ZKx9Yrd0HXjuvN2Hwb2YY+CVgx1/UPC/xjssgKzIPU
Rd+dBXYZnDYz8TG6Z4h6ugeyCV4U7ZhlUQpDjTAgy3bCNIeMqSJebqUh7ATNTZcV
CA6mUXxMguwDo4+IwRunSgca1z/5NxxPS+CNc20SVKuwr6UNARgiPJOcVVgmINc9
YX9bLKmrTzYV7A7vwnnr3Bq2/8sYRjxlQUbNU4v9iixDMoIjfYGBpuSpVABSLHF9
rNa34yvgrWzNjeZpgUp1aPthQIVQYhqKlvJgntglNGkb1si6q0LrP1dDW3cJ7XxS
`protect END_PROTECTED
