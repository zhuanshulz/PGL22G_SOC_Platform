`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3yOZfLWmjrLtlvihO8bIrUQ+Qn5Mc1UssVK9T5SGkjg7x4lKJH4YpY0F/hicoBO3
FC2nVtxgLOcy6Husf3WgT20OAPBoI23GrkBKtJM8CLi00KvfqkLdRiuH0QbvARz+
Q/YZuZ6m+892jjhem+5xCDYbnjt4FBw/hkYEOPy9pb8U5lNpL1tuCwqEPRNv/ymw
F6XWqqF5oJI+ADBZ0KFiYrPvNWa+gatIiE6RV8UOkXtFUkWaa0xgHP7CmCY762bB
3aIfztPBs2OzocDdnJEr6gdyqs7qnEuX9cJc7hQE9LM3Bo/qlw7rb8ng/fMsXmPe
F8AQV1RQBcDHHsJ+5FIRB9Vyipsrz8RQOOa5BoM4A9hTdzxifhEcDufIAe6RTKiz
qgIsSdGBytOPot6W/Uwk8wpHDTjYgGMhCGrYttWSDEuy2pU/5Ls2IT9FFQXT6MoL
ImIJPtWL8N2/zPz9XmGbN0BQznIQwE4oJicjqVlYOGbm3E6aN/JqTofrNfzFG9Ql
bOvs+tm1SkE4gcKys5koW0OQ7gLlUNdnRGFeW44MEY2VnD+PqDTJN/18bPdKJMIa
400+rP0xNP7uqzXJ+gK0iDSwfWNE7+U6s0vALkKA4r+5t1lOPjewMB+iopW9XCC0
DJGaaImSIc6uRPBkZNg34tC2PKXqicCVSnV67D08DUZVRAGR8aIM6uosqNQOpXTO
JRYYZ+2EXNnozTGrEBFleRL/3T43MiZf1jqqU2lCcLhJTgMjEJANQq8m8ngegy6Q
EUTIb6wHRVeDk2uS4EoQZCDcGv2hNqqdS7uulpbpSF16qdO2iKKGW1Lffva7V1Hm
+05FBVe3pp2lJPCsPD/45q3P5GuXgjKO7usAiKIdKuEGQ0hSKh6jjUKLSIIeu8k3
Eagmk3yw4CtzDZSuaLhmct6qd666V/1ABuRljNvC4ny0/dFTLrvRV+N1rbNJR92g
sWduzUAz7aNjGz2xb6X6JetfyJmqr3rdbZXGglDTSDZe9pk0WryfiBGv6RiXjTh5
37f0GWZDAB/o7OFMt6MGKHpVhiX5cCPzIR1icsqWpp6rQ6IwIJsHHtMnWdHHn9UR
zi//yjU7RDCNu6HWXfB4z/4lOta2EPHuDaCbUrl89ZFnAEm3ZX+TVvv4bN4Yhip0
Qn7bu2LAhjRDapvwKp98ZTgl2JBvdDndO0Eo0zhA8UtfoRNpfmQXuWm3VhNsXu3A
2CZMp24Pt7vkBVxntE/yT7vhOzIAQ45NlNXHD0c/5ZRgOztT/tCbJhdw70jCwH7M
eCxWWqb3RjMtIaDXMYV5zveBLJzWfPmHYiHSE3gvTyYCD1Kp19+RoGEZs0nEKxWR
L8oe/R2ApaFNcXmJ6ba+DTu0w7/ADlzw6zgAmbARaTBOOv9EdF4ttc54frhK2W+v
3ylNfofi08GSmE8dzl70p/eoyjkvdI7Lehu96h765VbHwktrEjEV1wKiJ+M5B9Jk
YK18Bz7dJFFmh6GMGMBj6P8kFy6qEbbVVtdVUTz5FImhTBT419vI1mJ8tW8T+g8w
qEs9AmcxxgXq6RrQwdrv+W5gjDtjnAM1L1aa3UTft0jDMEiU2rnbuy+6LbhbtC7e
yl2XvbWx5gcLNWNg3Fmz613AtoZAcWqWy6a2UGRQ8925OGfzXnN1LoZkxDnpcXph
3RUY6lJ4mqbMXl8BySEmGqAWsF8I3k+xx5rUX74ms8b0YrDTswS9YBACsebb3o/Q
A9FBMzRqE5AFAlTmmDJlO7HvFt5jCzBq87jJ0KgxhgZzAUZ+aD7jv2TN1wbsv2Kc
kX/EO/rd12nDADJEgKje8V2EndIx3bogZTf34Bh62CYbxa9h1UMFjw77HnysNbia
0BOETuL0VAk6ocEGbYz8fB3sbXEFfa+45Pml6yZ3yW/rV3pm4gzxVX/H21pfhH77
78Wn17TGy7S3TUcia4V2/H4C9ed63ryIQzNnymVVQXblWwDZ3VI1Zkaxh8/09n5S
MNM/xO35mdsZxZDqu6JMXVL9pJkO1VnBTeazhHEQxWk1pcLA/Fpfvigabe5rfPwY
6FxaDaPP+MpdSzGcfA9k6cjWTkwm05BPl4bFPhNc91Y8eLZKC1gHfe8YPIJkE2q1
p+HGJa4tqaBxwCnmwhcYaRZ5X9WaqDsjFpRAcJv9mSnNoNd3UoQxzGUWt6oxUzLn
/jvNVZegZfr7G19byncGJUVZK1m/BQBXK4xL3yg3hxbfZRRvIMWj9x6zZ7k1oENq
9JyT/5wNc99ZLn4k9e7yEn0CG7qLWFV1dq0SjtDYlaGLUQZNZWtkx+HG9PMNI5Q/
UTC90TAviqerSoOsjlKf15JnpsY4QGsQ0sygwZOJAKx9T1tW8GMgZpIQr/3qcVS8
MurtWs7PU+jQ4S2onz0pNIP6ZfpI2Ko/TymHsq92QYHtrCl9MwX94Isv66IfLMjb
DaAq0wjbiQq5M91QMj3yWaeyik30Xdh7mq6Sq5aqPTXxsQsBTdpTUjtOmoV0jHKx
lBaPksyQ5Ni7187fORiggkslB4JwGQ6myP4P9rBFgGTAjxS3cGTrxZKCzJ+Grn64
YWOz38Zr1mjrA+rfAsxr6gS1mpLGXKsJCkuMf3fKjFl+UpQPFAqD69ptIU5GkcjF
PyfGc+jnUSdOQC9fDo/czoEtVR7P37HtkawbWVC5tI+BRwY6kEyx/zB0rTmbO5EY
qT+jb+JzZzcdxNR9qNMDTYk04XXQJwQSTcN/Vwx/WezPyjqFff/hyXD7Nzr4XQBo
V0v1lAZ1NJRIFTIH12z9qmZ5RlyVstktH3p7DVqXnJ6EpgSbEJgJIM3yeOBgPUuU
MNYT4dDh9YptA0yTuuUJL3oVTRrS071JXE6ZyKdvQuZU5U4xdqyFHXIeNvy13gN5
++BQXUJ9TFkJ6uhLOqcGgvJRygYQF/jMdEZSUxBSC0RZx42llaO6qPmZ+vmwmVQG
rfdtxyKKUkg/8TtHghTQG1uo6agNtAYmce6TUwzZ02T6/UyXUQ0kPnYod92gtYCf
yyrGt1osxNBK4upjzszkDNyqy776Sfq8wl5jjcYLhR7azS6dMs0Ype7IIhn/Ezfu
WijfmY4XW8Ss0iByoImYtzXEA/9lja+0nxTVbWSA6nuqaGzcYQ1qeE9imoWVUKYh
aEfpostvCb7kfVjs7rcqFz4m90VmWGR8OO+pbJg6SQCS98Xg4G4euH/1WhQn/5Q7
Jg5GHTFO3g7FpJFCQP5z4+9JTqQd1zPRWHhTmVq9CpGGQ3BR4pvF7biUCsqxvC33
hfSo1Jg37dXDZjLoH92COL5uHuKzlDsRlo7LxWD++nf+jTrZWQuY6K4MBZmwwapZ
IJWJAM8JmbixKqlyMyfpAOXROCRvnvzj6iyrX6z+JlaLgcXfVsA4gI8ozHnZxyjn
vMs8yKZeBS1bqw31vtZP1bCYd9nFAgVZpWFRXI7omoFp19a6NU6hRCj4YAD9gliX
3H1b2JLYZtiMOU3dqZLOa2hrBjwsin8/XAxWJxQvbDnUUjiWTTaFucctGo2SopyC
5kV74+hHrxS+rrLbzbU8N5FKkqCFUAkhzLY1SPZsPx6H1ZoCfFu7mCCs8UJjxwki
9DmJ8gdul1NmiVCsmcfEAnUDFc2BHdIUFDc8Tp4jxZrKWV7Nd8Ylq38Zx031HjZX
bT41qwtIf+oPcy4Ycf3nbC22hah/kaBN8U/scRozV5cbHij4WytgvTmJHhsz2Mvs
P63vT/4QlTO9EraW9gpBxofnoyoNm7CqFGS3+aXliEA+CFNuJIfFnHAyri26Ss72
6PhNByO+IRiIuRL9yQ7kJP8SFJfB8P5XYshQ39uCrc28D3NwZQnGKXyskflFXa/0
9FYTHMZwgmJHjtmkMqHDdl+K+wZyM8ZK9G2d/MRmMOln8DwgUBxn3nIT4anlOMM0
iw+JifaTS3tAabXHjsRSB+5gUNBWk6pjA5Ms7iGpa/opRPon5k7acsDY7NKpCkYq
HABw1AJtS9J5uG3ZmR9qRkToCU6mW8yG1RxXZpNlNJiisRwfnw0qmdq2maGWvmjL
uAWpuGezMrfEiffFoaHx3pe6PbgeREQ86FkZHsZbAp/5dJraKqaxdmxjGkY3yO4f
qCfZbvlzvWjsjfdZSrQCpEv4PFbNrwi3FMpf8JUPMD3TvtjTSvaE00YRpUAlbUD0
HFFwPc4+m17uOHDX/As/y8cuRZXn+H8Bfdax9jDBvhj+Hkf+bW386XVbQWXk3Ch2
QLWRhJ39t6YqB7CUgznlaoP7ac1NOkkAhWG1DtR0Tp2CaBi4ro2mwvYYedKBSXyQ
vJ9X8e5n1f5nkTW+jH4bsuwZtCsHqozT71eNTknmukH2Rcj/qVaJjAshxDuFaNzk
GgQC4RVup+VjNk5MAG7tdWB4Wj1a0zm4MIkDAqnH7ptZi1GamlRUXwN78RdlzyTQ
IxwEnQThuseFa9y1Urj8c5zZj8youC6mcNlJJbaPaGS5KYnUW0WZoK78/0xp+qgF
8PUWnU0p3j07nWO2G16twrd8ZNjTzWciMNqIld14gNYZAwN8RQ5fiN8WZjFstCGH
ukYln+QGd9tAzeE22iHxadDkl2GEWKsWOuvdwdR10F3rKMVmVGlIk8YQSw4bDq4G
8BVW9npwJmbhsAEtYktiozvhICCsyn9QhrOywpskCJ9bH6/j3N9oYQfZ5XvaEzI9
MxAGFb+TUmxN7jDaaRKMTIrmNQmaS51ZwSMuVCfWR/h5B09OEPEGsIY6YHwUEEmK
mfJ409U3xEv031ylWTdjMII5wFrg+FGmr3rL5I9sgidnw8fLZQfeuKOX4gcI+fm6
+hKiZlgSFZWF42e0NF0Q9Cjc0GC7eLUrJ/qaCoAAtPyXdhr0Nw73FzTBKQ05gT2W
k/hMEUq/HHvOMEL0PkdZOS2waZpP/qLS7VIyCEDh1YMxNsfEvm4PqqpUDkJTyRSo
XOq3G9PMTA7gFUMITCorCnm4XLL4YGh9FS2a03l8nwG2zuFuiDuOZzZZQu7UhNQZ
tmYR6wWEQzGtkHB6hQAXlAs1u8BlNnSMB1kQgSteViMorRhCTm6r/fPmpjMmYS1v
xjJCBc2nZOWs+WdmOqJ5x0Unk5UooXhXyhdD36VNO1mCTDPIkzV1P+PhZYQ3c3T7
WSu0z4/SWvbmO0tzXKEyqHNnHQ8Cvbs7i1Oa54nU+CVfQgvJq2aGKbsRjGLNOJnt
cCAak/QJWRBrlQGbyb5qLUv1DszixIdSqBYu8YYiZ5oX6m0w9EuRUFgQDN5xLY3c
u6jZ16mm4iZE19Kx7oge46PN+dw+6FHVfMERXa0RMYLvX7VIkCFIbYoMKtyqQnKR
ZYJlpGamxh0slWjaoM4uaLk4ooEpg3kQ1DlPww0PiFPqY0gQw6lZWqmP8KKV1Af7
vqE5KfJeaqW3P98P23mhz9bb2j7VxrW7DLN3bUK5HmDh53IPLvKDJFWP2QVjzrR0
t52JeYzjQM5HhOe/cqmPgGA6M7Amskfao9eifpGYPhqCo2CD6bWfTrL6K9Q4iMur
p/RSW7a3OSxZ48zpvFFI35Wfvxw3Lxf4Gfg/SKrVOjo9Ubc/OmtLqryWoGu+toZg
uSi8YPSW25sUxJWoGsRESkK3kZ5wTQKg23BZ6RAX9equ4VOMpteE7qdyD+L+PRQF
laSxgvAt5R8E1c7sLxcnuQq490wrSWExabV0wULEvzDZpGRz3qh3Jb+R9tmsQe9G
0r4O+rtHOC0zNZYpL/QqtKmqEpFJQyzsBSqEbKX6Hs6OMTc7aNkKALi/OHeJWIGw
QzEF7dW7tAv8bpC4TfFGlpQXyVLZWnmfWnnQ5TQYqOIlJA+2V4h+A8yAeFr/+uOx
f2Fa3QJILmsRU3CoqutzL4r5uQhiZLBN0ZCZRmsJ8YmZwILzqwcyBK2etyrDWjXJ
JNlxJ2WClyLXCHl2Si8p2zN1vmWvStfeP8SJJA5mLDBxJmPQ4VXheTg4kMsYMtjc
meGMmRLpfNNEHv2Hmu+FEnkM2nYCZXXBrI8MWjI1MSE3hXfM6zybRXluCniOpKP1
CY6veahbzrW/Hev+L41TsiGutgOWevTxVjm22j+x60iRvKX5J4iCiactKZU3EgPL
PXqKzjvgIqLS9E2LT7HsiJRaYy4773mW5Vadx5y6YmA1V64KxNuDJBuJG4O8PeGp
dkGROYscZ4At9LY3Fee4d/efdzTuj4oBZEbkx4SNITK1fbebF6HZBjtNCtpwcOos
IcKjHMYbdjdli//VMytCuul51R1fKPKIlNmz1dtvEqs=
`protect END_PROTECTED
