`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tI/R0XdX7E5lQuFnj0FuCwHT7V/FKtktraOADtJpvX4S/sRtw5wnrqL4QeOnahN1
ACyZMBx/1mezCkR+Dwin2w7F5vGnR8fTXnKMdWMxQOAHhs2P14+vM7Vlkrof5ltU
HybOVkmCGqKmHEuwp+95XiltQhGMMJOSmQv8/HmEkvpgiOOpaVNIsPDq8LLj7+04
beSPCCKIqW4mZdtE4JN2xhGhckL23sa44527RRegBM1jySDqrSlAEwOTV5j0EstT
jWksDT1ivyyLWESY+k/66vAOnnDGZFqnSyOZ7A42ABC6x3d0VtgDyZqGnk9EcTlE
8toH6uQqSJN54YbTPPozMjtGS/64Sa2/hTsGh6sy21AHshy06tXC0ft2ayaFaQhf
sJfpTH5H6ypkHR0vIieuqJkV8mZ3CHR8POMgFl8wbbPAzNL1h0EiEm4f/RtJqv+T
iVt0gEDmZJWp0aotmc/O4/YH3DJbJSRmxyp4rdMojnkB8u1jo/Jsd80lLAlkg16v
Y8SdV6X/bIYvvd383PuQFjSCqZPaWv40euZzCTJOFZOBRldRAu7HyDhb9A6hiwMP
72B30hjZiBZIcuoYN5uzXUQbtJFeYtVdDWL0esvpaYpU8pRarl8mVRivFWmlnVPH
yPvQxzdI3kSND0VxkzGR7NJLtKpx7aDj+eR5lej/41dE/bv/SoceSsmouyYZUtJm
/DxC0h9y015qkaQNxtY/44vEe9+2XhJ/IHoxzOyaaE+rNu66fk8v1zcl2dlarUS5
Ulmz68A7bdLM+VmxIHmUC7gTEcf7/NMqDbEnU4JdrtdYzupeVRrLh7+u1GS5fKaa
GJMHJI/vmixZYC/wM61AEyCV2K005xAnLHipJxqB2ekiGyCc8e2kj0wOkgW+htMk
J7yg9Vo+keRLM4BOzUj2/kmZBVMcHTS46+pukOUHkEgrQEuWKieqnehQBaFBglCr
9GMd1QQz2bDvyE//VyaCkJ2yaPA+Yc9k4hw2pDn4PuqFXcwgPGXlQPo68ddQTNg/
6YUNNoUlvnlc1FVZhzYBMcC3zB24DOXbYxtbzOQEJg/LGwA4BZXBjx1wKfLZA6vN
SU6jJvc9QIRhJ5GdYPp+U0Er0Fm2B+uyXks2eNVk8C7MKeWxpsegn6MK+jk7Mpu0
Y2rB/CKu4WJwq9seyc19a/2qbmvQ+D7mQn5UysrD2V2MtMNxb/XpmWwG3xaBO52j
W9tBCBYItqeomKmuu2nY5PG/sRQbtEjfcHu8NWv0EKOG5uSwKg4BgBYPo4UdzmLZ
e6I5cYy+NHjB7gBlt9MlMRmjwFudApNW8Rp0aLa+LPoNs8ivF7PIrzwJ+B2PfVeL
LiYFQybDyBTZh69pH046gY/45gY+9ST+fQpNxj5N+4m0pennmjz6op5U4unLC97W
Z+kuknoctMfAzQVdOb6tYfm7TjeNfgrBD7MPkwJGbwo/cVLhmNItjfB25Z1mXcDh
8YEVYHIMdTjTma+X2SjI2FvmPjc/T4VvC78PBRSorHx2bBeDUEDcuFNd3tvTrFcb
LQKO5SxMXDMCwR72LWzol8qOdkQBX4ZhFzfSndSPG18f47qrJQb3v6hzVnFUF0Ij
yNw9c3myqusPA9fB47RNcfObj/n/UoBriNPiEWxyTFGNoEvEzzpSxv8DfA7KKMVy
twMMln57qe6OSizm7FO3TJ4KV1g6uehhnvcqUmMEfnl3pN2Xbd8DAOoKZTMYuQgs
kWI+p06r2ieBW0whum9U73LRMykzKxuKl+UuPAsK0PTHoVGcW0P55fPqmj6RAecI
25vT/CWpFKaeOrJaH58RwXBgEYVYrc1ucJIDKRN/7du5sQm2GFMeNmq5E6A9bdYo
kmbfW+p8eQZMxJPznS+Z4NGknRT/L64nplIwL69tv6tPZxzt5LSt3MGVDdSr5j65
N78Nkb1gN8ik6KwfDEcXzOzSkgbhceRKhSc1WGzgQUZe1tZRKCUKXSEVhVNlAFFt
qKKmL3DdfN8IIwiKHCV5d+fbmB16LI04QqeDqg2abVqxWPX17cTfYNhRZBU7L2VX
j0E98giizQ+zVLnR0Jg+eO/yBCvV0cQiDa4t42RBZoYo6s+Z+2sf3huNiEIFW8AU
BXOYTZmlVzV7XWSlinGYZHEmlszOJkp+5LeQ+ViC1O2ET5xkMXo/UJ5B9J44saRt
j7Ocd9sy3O19TOqKwVaJ1NhN+2GVqbUPeyUrN/JaYqqfWp7e8vlgTDLHIo5qc84k
41SUPDHp6oXaoIEdEpe3wZH+uj3WRfttLBdv26BDiLH//ZxNe1fBYA+vghGtAVlj
1Im2Jk4LSCnutb6spE4yJqe7UMk+cgpIJNRkgwvZgoWteo9Db37V7OkDZr7bZ/le
OXemBxvwBFli+4RiRb/gIlq/4IpwWmsZgptfFpEvT5Cl3r1tjKR3Wh4QqViavHab
jzTYnU+Tk8Ptf2AZYzQdqFFVuHE0xcXk+6MFn0Uj2W5XUHjdL7wJ4yamUP09mUWD
ZPkS37mEMTXMAkcqWtJFyUGU6xkbiNUge5CZQIC/HufffV1mWR6DfSlNEfsZb3hL
ozjIV5qOrvF0EQeuXJhVjg==
`protect END_PROTECTED
