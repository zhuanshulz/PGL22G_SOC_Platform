`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WTNIwEPSsrgZmNyaccFvE7fAPo74M7lrdRLDtH1wArKgo1N/e3q12JTM0joQcPsa
Zpsf3uRs/dPh7xcnPhS8HuZzoo+JZu0eixg112cT2EAOqZfXmw3XL4R8rw7e+yks
hr5jELxWNyR/CkOnDXZu7vQin3nE2uHShVK9Y+N8T/k6k5sM/DtX2VyyrwkQVNV5
eK7KMX2Cenp370+ceUaY/0gI7ShGjZSgSfR1ufGXMQqXADe/YmTwbJ4zIfnq0r8x
DeDEwoYO6g2sjkWg1469Fyq21djPf8jJIE8I6Qaj9j5GiekQVuiGNLLbuf0Ef2hP
O/TtuvnllF6G+6FZ2aLdeEjeOLOerAeLcHjv8bdTYY/L41YHGlE+skLhx7N/al7C
CzSjD2RJz80PBf5elWAutitTXG2/MtYph4uvOvuY2RJbR0jOKsqwdzF9bKXVe3aS
g1c07j1T4hJl4M2dSdFdlXHvCAAZNNnLjDDDZ8iRnjDY3CLrocE54a/d58Ux0msx
cMfLgufS/r576WVvngx+/qwLpahx0xC0kIMicC7kj2Lxazq9XEU5AOS8j3zBt1CI
NaGCFMwzXLwz8R9ASD3o4tOhcGH0zfa0aPpyJdPiAitJgAin+UCoDB1NQ8rfk0J0
buKJ0bu+aQKqI6EXTYnyBfzAN+yGvTLE/3/kcKfXcN5ZCsCOEUQC4Wrw21Bgr7dE
IgKHgLS4PalM9V114sypztf+eMsoXWPKl31LX6Rkl4lZuRcOk1H4cTVLDpSyMbfd
tl8e4fnlE/Li7JmexwXL+vpbxqFTndcuD1lHyRgjxW5KB3Ip/wcvm7ZG/V4/HAfI
L4hva6yV5BsA5x441tgov1uUQtCP/7fmBpFct+rOBus=
`protect END_PROTECTED
