`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IOBcK+T8w08FFAODZwze9Z7KZvtzZ0Z3T3u66RyFU13uuzN+A1eHSnYi8w4TAHC1
tOCcQEowW297weXxFq9VxdlrVbtWwcU23TW/WjU4d/5pt4hZq8aSVDoA3GcqcLcj
4coJNzHfL+5FuboV/JpsYloNumN+10FFbeVBIxTOZaIY3xXXjMwVG3aQBYsnuefO
8PoYz9fAija7xopjmsKDulpHtZFbuT67jtrcRBMbnxHsHwn1TPTNbVEhYPTn3B4P
drmMz/XtAdwezEWqxJ7C4LszfM0xLnno4pxNw7g+n9o1U0zq3oj11a0wuMOR88HC
NiEpgEbQz688cgXxwH5gQZa06iOubgLArI/qpUxvV21/EMGgVEkp6TlXjlT6PkVr
Y2dnfnTEPd2Q0RObTlg1IKQctVv0gVZumzWKECe1hrJIU32ydwwklwktT8q7bFVq
727SW780eIT8ODk7OFyNA8bjXbElCJvVsS9JsNRsHMejS3qRlGHr3EUXhjiquG0O
+/1f6NzfQudebL+v7ZnWOgQ/On44V6eeoEEQKoxeh3F8gYjrW0ConZxj5MxZxhvK
tfa76Mxr6gdRt/hSsR5o/kw5wIYkpVhdY/M8C36cQ7gLoNURD0d1b36K5f9HGkLd
Ke9iXOEjj344F+zOHpY9ZN5gJIw8pA9ADfYuoS3rdtaSRFf5c97TbB8cxd0M/s1h
3NhPD+9X9TvxKH+aJ/O9WMbmIdTy6aeZWqYP2qwqYQ8ShrylfcH4KBTlLp3F2vB3
hr37uSoQOtuMJN8juK4M5Blv2wUR7Lwxc+z22ZRXBoc=
`protect END_PROTECTED
