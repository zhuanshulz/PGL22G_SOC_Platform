`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Whc8bEyvdv/dNLYBybbW7d+qPLr1o7xxEWeCvw4br6UnZRllAHU+U2fZ5DOUnbKC
8cnMY21q3omfz9HzE3ng8KV2qKTqiYyMTEd368GpjlPbEC2TXC1+IBmwPX/XEIYv
eEp4Vq5oRJ4PI+6XaNXi/dpaeo/3xtkAaeheDj3Euc9/KI9OFsD0x5s8A50yWW7+
Q+rQevA3TrNRgn6ac+4XF7gODVKqoucCTHK6G6SEz8E82Oumg5zUqLh8UnC9wbDp
9tL6HWDTjf7YVHsXPHq9eiVA86iPtzTIhbVVs+sMIt6huL/fJf9Q2PbCyZtYqxPO
pB86W83oG+VlLHMWRt2wpFUxbPai9TzJxzgKpBRndCqPDHfnU0NF3LQO1uMDWMz5
lN/8qcTspGr+LEdgj9JQy1kFYywnYqMP4d3GaerM4r4aO/cHgXXTf1nGCZw24094
`protect END_PROTECTED
