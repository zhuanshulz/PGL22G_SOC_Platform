`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dQG4fMV5HKZEST4+JTVTEJCZr3FAayOLMiX6OnVvVUMV/QLLqj+qGfa70jhWzNZK
PtHwpHSyzkhdEm3lRuWeVPsp/d23R3VhjcbAqnxYpGNyTFbBdKjaJwO1CGbmgaRB
wcQeCNbACrFd9NmQSy7YYjvAh/Xlq+1MPvDCXlH+PY5wBUhz1ZF3wbXD22SXtx9Q
+UCB1venBS/0NksC7uuUcEltmKVHwKgcZn3QpyXxXmoD9ko4YvnRIDyQq48RelkI
nhxmbRZXJ5caU8266RrfXAKXT+P3MdvHxmjIz13u7OvJuKfyQkCAzEaC+NyOn7Dy
nstnsMFoujafz9f2LjgEBzN6SjR+J6o4Zhb4n3M3er99cOc+uRN1m25vrWA9z/1f
Q9WQUNoO9BH1A92PanFRWMpFZ6P4Nk015h5MuQHOdRdLU6qCIFqzvYUokTzWpQHN
kIBx9xktIxPGf4As5RYilw==
`protect END_PROTECTED
