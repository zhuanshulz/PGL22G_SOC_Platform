`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qew6GnIHw5BoKFHTEsm+jts3Q4uAStQFrFpL8Do3E6psDS/cmRYwypek9ub38490
oX3zaL43QmBW7XQYOYJgO34WkjHqUBaV3xXbA7s+mc8Crx8TWuJryp7fiYJwTdXM
UQ94+bTsXkkmpc9sb2LGn/7JANsiyaFzWTIsEuPxztOpI10JvA3dfcvp7lwflYgz
ZSXwAZTxXSIw1LmFvnOVJuCHun1yrEph5r1a99D8aEYNNzdKqNQQes760UgJy9x0
fEMzBGMU8FGupMQbCgMAL4VC95m4ASsuBDYjvHDGQ74GjDnxbt6F7Sy7Bbvfn7Ea
1nD1OUDU7NDmMK/RJxxP53qsYT2+Q9SPYwY3VYU+5XrwmIHOQd57GWmf6g6YbZ0u
X44nB1nFf+pdG537qYjwUJ+ocbLrJHQLLPl5eSJYQZ0Vlb1FL2T423mVd9zYwBBR
4h3qUj2UURjL+EREet8rVcAgKUnqbzf70hq4etpNkm08zSdLMJbGfthqF8QOQM36
/VbLth6zO5HKnldQRbCVS1aXI9dajucqYRxwgADNPCoQfMzHSYBQ+1dpWR5IZaPV
no8L2+jQdRSQBl+LySJ5heIceQ8vGiRLNOvUzNKdBWjbH2oE8vGFo7c4INoZo/oE
4mjWsn35pIoA74aTn6e+Asi98mLIY9hPWtY5V2eFTd/Q3u8J7gjKV+tmSOiN/agZ
USvuq+72wSqCIIfTiPPk+pIUQyHFbEUqREXuYyOQKCoWH74TUgI6gXcWhQ2jcGQS
kLbow8iNz2dBzqCVuARABX62HZXj9GUEGwn1RWcPhvaI6dL4hHRs53P91V0EaDRr
BxKDszBVVML3FiVlY0N+HlQqnqSTYQyW2gCwSXPh1Yddwba+d/NhG/4weL2QjHGI
eF+RjdtAtYfxjaswAeKlirkG2N1PmKKOJSLzwfOD6H9/N54leO93HZfbRyHKEMr7
WEfWWFHstf3qhc9HiR3030pypbKilWkOOjJvjDDtnGDF4V7lAfiqMB00jh7b/ern
`protect END_PROTECTED
