`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bTY57Wrz+TLU7RvhqBgtrI5L9wNhvdwaAtM722i1/WitSybcTRNYHxZzo6cpMMuw
UGDczq0VrVXjPwBd8EvBN3S3gSGxCYVrQWScBxqlpMCOqoaLlKjzJzCl55olsef9
TZgnLXchRWJccE+Vx25dgNKFc7F1xT25jh4cOCe6aThMMIuWNjOM2c9H/eB0ys8U
+zTNA8ttUplDzCeXHwSF+UJDSBQjgXVqBDJFMHsNowZ+8MNfmmVImON3tSk0I4nq
rd7slH7eEq7kjPmtmKzps5eQekjcDqsnr5p7n11JoLl0rU0CgHxSe/Yky3IOXWqM
dTOlTvXZE6d/REA+Zudr6a2rgaiqGuruMffXB7h9HZ33XpUtBQ9QXuamrj1IZnbm
EUCX0z893CDdNIChOwsJl7qOd0QASQB1ZTCflIOgzGpXFUgzURO+m6UGcSwk7cpD
wM3ULgHYrt3XROO3qTzMXfMTEI1LclKdt8ZV60fsJq//ESdienfEU7Z9AN0XwAaV
VY4nXQwkUnXn7mZVNWqbTjlEdEDmzaYPGofmuEeA3w1OzqCm6aGxjuXZJQwTyQYG
/MzBfLBxy0UkMUcSqnwNGAaviscVtkzD7UCsEm6wEWL/4yzNebxr5FZZqBvNhoOh
SN+E3D5Fc+XR53pCAkkj4bxvP6GIXn8ZNxyTss62I3gvMTRNVytwmyEWDbsJECup
Kd7ImhqO/cc2HBBAVLqmDUDfP2nQXGt7XpQg0QygY/BmOnJJaFCpWXYN2w+RJNJ2
7+dpPL1THAJNf+YCUGC5oeW9jHBAUEf94PNAk8FjBQRAd+Xo5+qtqdIpMO8C/bCw
3DcnnzEYb6VHGVwXn4dC85wkF6Mm5DtWtOorNuPVpXkZJUr7hJuWSsoDy5B6+PHP
`protect END_PROTECTED
