`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QB7hlzwFoeAyX/QwkWW0ngqQef45SWzeUxe/koaquL8W3VlWy6X0X7l9QWlBwIgC
LGe+Cw2kKuCWSCX69JSiICavEqGe2Rcpkmz2Fc8K7Bv/G7kD8zGy132C6Rfp7Zna
vFCOD+FpBpASd4aKRDK/wznfgWvyNVvaZzxnf15J8pEkqQUrjRZYLTBOqP9eqvZN
9w27nrAAwlaXVWIr6B16ijZBRxyOy0fBn1rBvnrV5xSq4WsHbe4yt97KWN6xvH4i
01kzvn0ECYtxtlU1Ihc2TAncS5Nw4BoQxtDnJIlb71DN5SoJSh8L3m6OZM7/dtx0
`protect END_PROTECTED
