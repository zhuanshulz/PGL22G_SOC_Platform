`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGEo+o0a7VFIV19y0BruK31xsYdXcWGpeY6YgwfJ2LyROLutMQVPat6uFZ2uzwpt
WhGKjQOShBfFpOl5SOojjyND4bPdWz3irH3t/sKryLZd/sH0QWSTdIsmCc6rdHB5
VLxDV7g9Xp0pzY6LlPqEEf6QdNUdp4+q7qy5BdXtIZGiiAAUqwiaMA4cAnxitkkt
6I5caaZBPy/SjjTukLYMgP/5wo7dTYTcCGXNV6Am8iqKp8COa6lmPoBRgjkfx35F
M+HoHdvYv/3J62cBSKXKMWcG5keUgEbUifKWvvYkoAzjFYQGU2Lu4MT89joZyVLz
8G4Zb1rVyZMP/+s4asjKiPYwqmBuxb6mrc0u0IsyrMqaxtV3/v+qqmHJdb0FCbEa
DELdmHp8QT+xU88A1CmxNODTNZz/l7ocfKG+JF+UmQpFPF+iktIvgXOqDhtpzd53
BO9IhxahXPYMVFIaKsavMylUQLqCcVbCyOTe12EJJ410b9zdPisKSM7x27+Qpjg1
V9qixQqD4RDu52EGDX6kuMNr8Lbwgefcb+0xw2TOBRDhRjrsSk1kmQ0Hytq7fhjz
h8sew0lVuznC9AiASNsyAZ8cm4dD1HaoXY4zai+zW7FkYgSTDyNz5gNMrQoRi7/7
k85HrRXlH4GfUQcCVI1CZrQzJycMptv+RWSfd8uIr04SCNTY+oAtDnQhQtmPMguD
OzZYXJ7Ako3DsxXphxtkk6P49hj2Z7dEnIXe4aX+GnU2teCCz6YT0cGWMuA2YoGl
NyRbuvsCcVI1ieEfcVX7Ddbbt5fLUbBQBB/24HHmQnk=
`protect END_PROTECTED
