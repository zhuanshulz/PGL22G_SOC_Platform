`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QcPKFzW+8pt+xFDbjN/Qwzngvbn2tCNuYQ4iyU0zdFX22cPd3y/34S1xmFx8eAp
aMsdDkr3eociNq8ehjCfB5mqRBtr6aRQhUeUJAD+gFGzxsrRRe3NlMVcgd45f/ar
FQcansAxZ98eAVgk9OV1a3hbf6mUBk9eys2EJWmva8VwxgKO4469LcQPni6cozKU
BEk7Lm3jxAB9oBeLrngmW4VAMfkpZd69bqzfishjUeWQ8uSBgIQHBmLjOuJtwfMW
wInNRw8qgksxyOgslXutfMqjIsnCuo6ngibDS/V9lUoO0Y83KPfNEPl4aN6jkOdb
/A8YX4133/59lwL0V4LRT2vM1TNf7LusR13r9XzfxUGeyf1p9WNOp1Xs4EAdK2L8
AusCp2PdrsO00FTtQK+Bj0W7zzmyVmJUabA16GR6moZH1aDy694htmCA4KtlNgo/
tvo3Ci8Oddge3UYv1bR8bWMOqS9x/7Eyh2MJtxwLNnvNsk7NOqFz50cEWURRTexj
4SejytxTYsTRGS81Tr2QcefTVg8yrBhgnCMKEPN7AAWs9u7/Ey5qZqpjnL32Fxe+
Rbas2UZgUnSQjiE8TiFlWLrjiY7uUy4WuFNaX4181TdrRrHVZ/X/070UXjdc+wo7
mAqoh8krI8qgKuDAiOwqxq4fWlAea95g0aEGkZhVttjjRRSPa3SkyEBjAZ3ubgpY
7wu9vhhZVWT5j7JlypNlrRQ+muzqnmH6D10IcC8Yiagks1habqf0cKr7p+Q3WH+G
fENN2CqA3lfm14OwefKuVu78BH0J325korEkyxhcZsGp3tFTyLiICXD405sEeyKG
rv8jc9ostUrwJ9cY9EHDHKaEH0SNUZ0sFWzJMX9w4c6sUB4UQKfOpgC3Ph7K07Gg
+wxOMdVPxDBan4F2reXm3BscxuCYsdnR/zlK+DxPPhI3znAzVePolUD0RSnDyZMD
GKMP+UyDtf3SAkf04eZhvMOsnSQcHuz7j1USiVPaxyxwU9kG5xJVMNzdMdLAsR5J
3Rc02wWGs1+x4v3WEDCIMFNa773Bx6T3Uabyd+x3qyhIvNioslgwub9m1IQsRkLL
jhznfAH3lBjOGRvHSY6A0V7hue0473ssyKw8EbS9J8layethCyHxA0YZZM8ESDIi
JziD1WtAhd7CWg8xgX2tLrDdCUIwy3V0IpUlQSRfeCJgX9fWQLt4LCc0ZUBeWwd/
pebBJo3CLMliUGLSQQxyw6/RBTuykxX0ZfvComPkLqwpWhMdPervNPTper2dSofm
KSCtmdhJf94lzu4PsDuLnxrqt4Pc493OsT5A9hm1HXY9W37UeYc9vBAc167KrKv1
GrriEjHb8r7xXXWQfTTIXAKxRovQ0oMZ6IrAFlRrjy/iChJZrWSb9qbCnEeEX9kO
xNDHyeG755EY7/KI0T9mbu/Fc8YzSpAaNOYQ/RDf9bUYrQnEW1OBO+aM0qHBFhOO
I9mFJBnsYnGfhcwcF24ghFLkzBhRkoz2rFPwSF88wWPxPX9/UB46tAgVDKvD9Y+Z
UE1onNPaQwSiCeJbWhB0qU3bLZcrdoQ57PP4jn/Ko5mNCQktfI60PMxsCZF42ME7
TcAFkZ2/IUDotBXUzhmfXUGKUcERRKwQ7ggsy+353ICWQA+XcPX6C0e2TDDVjSlg
WW7xr2w6bpq5wp36c2lRcsCvkC3kHxs1t3EYtmnF3A08RAFnzS6uzqiEKgA2bewR
l0avS0AYaHmVz2Aolhi7D3+VCHlTV7cP1TTuGAwybgqgce/oxwaoEwC2T0tAy+iX
EkUDN7sQ8Dq1/YtC4gb5K0hygl3EGn22L4NKtLp/FCPSjwUrC1K9jCpP7q0pegL6
aDW75oIu4EVFdqcipr73BpqbK8hlUUgSzdjccgNGLzNZy2J0If/kk4UrpRTvvGZ9
fdu5TcYwPrMBMzts8x/M77TIs7UWEeCD6rwpBqJDbP1a4JEsZdpd3vbaC1Crrzyt
bWADzVGd7CS3bxixuWSvSHlTI7jlODmkD8lZ4spATqvUyPWAUJBSfkZPDLSy9/wq
FA0kgEpakrpZNePdUnG1/s54u0ySmoZK9U1mV2AsgIo+EZQhIyA/0XubD7RFJ5vv
X1UZokqmXaagjy5HVxorsi9SMkDQTx7+vuVAPsST0N2PbIujs9UlfBsBf91enLV6
xOpSkdfBCoh66isYz7ZLBNPoTW47s4iiqgCmqyR+vrfpYn1d4rHw+ZCx197O7Oym
8khp7p93fbIZmGFcuEAsardFortRjfE05HZhmcENJ9QqyRrvg07A8QIIBH6JTH+7
Tt4BsAHBwRi19hdq5IxS0M/X3NKjM9gYrqwy6JvdgkXwUcSk53Py2Cjwh7WDeCh/
PAu2twbBG73nTU8zoH8/cFEJ84mCTUakmKFZ3ye4KDT36i/tEFD6CZAOuT4sJcXn
rTtyW3onqYNSmpmeQInr+h90mfr/eh+R1NxDKUTkbeVDK2HQTImKFT0SpmWAdzUu
hYiDuJR5AU2ho+ekQQwS3Y7LRKBm811cjl+HC7wt+WyeWls84vFn/qIQPKHbqPtQ
8Pxr617NiZXTLHYgU2Wv4k8EyEGhvIbwZQrBUwR9DcfTEq+S7hqpEVB+USZlp2dC
akBHtPHyx5KP0O3iP7jrdMA+I0Q60a6PSpZ3q/c84abrZ53kmD7IOgO5ZEueU6Mn
VRyeGwydyu9FkUw1Zo3SjUeNKwtjeKDH6az8cneKNiwDW7blFz+aSOLKGQF6saBA
2ayUyAGd1o0Ccsf3oD6SMN8LqATHvMI9/s2Ne/X3IoanFNHJfSJ+zKDPmu/3w/wR
Tvkc4J8I8rKE24o8zZuCIqCC+6Zt/+QIRXIn0twURIxSEmpusLOLMG6qSsBHbIkU
hy8T1QbsrKdSbRNxhsk5HiJkKY6RHdwXA2E0cbg/DevuiEslF5eE7NdZ99O4Kk3J
X449WWf8Aah6poTmoQXOY0jAPRQT+no8BGJsw/zfv5TNzy9LRrra2sCXaTVXvmsN
0jOz9MJF2JFTydU0JG5o3RJ7LsXVQxh52AC46CBFHsqTCVHFjR8VcS0+qUK1g11T
VTvroPfH1GPCkKC7cIcapqTCFCJZ1d/CtOLOqBycdRXWsLNadxAMWv2LJgFkZ6h9
4j0quUB1id4ZjWqkiYI4BM8nyRg051M5ZxqP9NFlX5JMnWk/T0/g8ApXgo9DitlU
TzkKGVYI6X8gEWqQ2VjuuJ7Yg/dekku8vfioQkOmXQMSUDw5hdKluTfnxioCbWOA
2TquPFYfO2g5byfbVa5VqLaAn/HhiPq4zt29G+QY4XEl4gmx5LOH5VAnXyIHSz7y
woduxrlL/tggFeHxzT6gz35MGvgw4LcKIkoLxhaP9mHmliMmE1LBzjwTax3So8Pg
S4oUZ+xphUe/6/x9H2UTab66tnPWr/BWoEY2ny+yRo1PqN49Co6Ftc2fE0jcLEpy
FUnSU8sgzGs8MCEaZVy0myGSEmUjDJrQSe4ADOQbhW9nCNEGXWIPsBdCEj1/1p1h
NcwWjTVg+PrFvwW1YAzR6FOvNeoELwkxZ5AOc8S4j3O6kqSZkaZ3G/Rgv1zeNIUv
nR19FDWpMbcQXAsEWUFyy1vbNjd62ZoLyWcSGr/7wC3dB7URa6ffJUwGi2HBt7iZ
fOR17Bwj3NPl1Itxlp1ln3tcOOYaCUlvd7Xy+J1PW0IT/Grc/edC4y/haAolP7Go
Hbp9eONA0vu66jMVfL5TRRiX3rwChVFD/ciVd3EKrt9RZkeFvudMVqA0dgkeg3x8
op1mV3WyWVWitWbf+/2b38NYleJ4mQ5fUg1+hjNRx5CujM2xD0uwIYpprzMDAY2r
REi5ZhEtQ3cHHhsfbiOJUerOIIvQ3R/UQtwjUmAnCFSGZGg6KkZFjQLmczfS4kCz
6yZA4uCgLTfsZE9s/DeMSTb1JVgPLX+FVPtogE/9t6MQUbkOZhnIWq1EYiU/e/A8
J1mwQ+ukm2T84sGxpkvaImYhKXPrOwnNoZts03IiXHhx4FdDsQ7ugqwo/o2KiyM2
GmrOgkEdnwCcYlbnaWVzV67CLxduP101If0MuMAhZj9UrCK5joepuQa4HV96lzx2
Chp5wHbxXH9CD7sfTU1o5pIaN/EhwQI5Q+R9GHm9FEXr4e0txVmfpQd0fO/QRAFD
UuJ2CekbUTsMEMhFpxk0aMbHPjSyr0ZwtT90Sra5B6v/KxoSTNZ+h2+86X3ILMPP
9KuFAK0yuBRbggs0gfaj9hlcvnIAuUcpL12kzQkBCh+WxjME2zpVCzV+wwgNlvdb
e3KvViW1a+GGuoS3MljdYSB/f2rLobisrMO6VT/xXVFj44fw+8c6sf1oLg5eyQfq
xy9xsEv54d4g3PMnXzmI8am6j9cbvbHpQ7FmYKvjt9hrdaNznbxbXCt0XZogeu9S
/OmUBE1W2SrZHCfragrYYM1Epv/tQQXvbenznZWlKVbv0Cle/4P2W4KCMGDmVFgv
IixhYBNS7Ymn3gV7waKdbe9/8P1284Anw4dCDiZAovlKuOwRDOdrEpVNTXp2IP3E
gZoHvXtlSFBbiiAM8TwJh27xomfw2WUl2NZ6hbHkdA+SDabeqxshrqar1QmQ4FNv
0Vz60sU+oyuThRYto1bPCxwvuI930LI2gI6LYwU83KbU0ca0anmlDiuwBTBpZdG9
exTkMHuZNCMYAZqcR/gSO57P6Igrm0cBV0sZ29YOolApJXEOKFgS8iflvRYYaM5J
9uLKAvLWkiwr0DVg/tLAUr0sMmzbwDBu2w26//8tp5zAatTD/Y75W6cuJIxiglBF
jnNmBgFfXMpiVBrG/09xiVLJ1S4ep1qZvIYpLWM6TqSJ0n/McFHdsl0s7DyaghX+
9+nf+P4ThArSdNKKlIxTutcucRhXNnYp8M7QkhQWn/KX6VWKUmDTYd7o95FzDGgQ
KDKisY3jMX4OjM8Xxv5WvxGgKIgHi8oNUzQTHC+x4otFiLBLkpGxnop1AsbjGLjQ
FwiXcrUOeAkbfzP43EO64KycmHWRh6TiXXq0LP+LF4V/BKPOwSa+bGWh3Wo02BYV
N2+MT0Lk2RPHZ58+38olEaVaNIYPfXZaORHFqHW5p2SR421ZeC+hG5SUqSplGa7I
5wotLgkhLp0ra9Ro+XoDIkBgGXj8fjRNy4WDWr5RV+o2t3OJDLkrKr3p+XzaBrxR
YyMT9U1RBzhKvfqySpEb2t8phfW6nnnV/iaV+/QzQ2+d44DCh2w1XjL/ylKERgZn
eo/V2ssbjQl0+62bxzfkPBIbUO/GLgybaxYdh4TVgOqSvcIXqt0lzR9DBOfwy2wK
T9TvsKNw8coweCA8qxkvGYjJbj9LQV4MnM39GK94R+dl6TD01hijd8viGkACOa4F
cxrouNq48B/B3haYidz/9hO0jVfEeGuOrdynEUmCl3cQSGPau3Yaz4qdzThKNvgB
qx3cIur8OBmTVfwEr6yUlOfHU3/mAkkk3hmSgKOr0aRzDSEva9CGAoMnhTo3eXVm
JQLC959XR98mN5JRYE98nr2OHs236HY6wj4rWefm/7ryYpRmq6RRpZOZxA6KUUPt
NJEEar6Lc9dPKNNRJWJnNpBVmW0KQl62F/98DWbcyN4y4d/aHzkhmoI0EA8KfiW+
a7kSZsRZPP6y2OpQB6SSfU4BFHlo/rtr7ycoVWl7IqLuVsgxHiSAw6gmNSr66rJ3
be7qiVIulcumv7gnYCta58/m1Q8BOSUnRpOITaWHf3Jnlvqm35+RELLO2P1Bh1BA
9Qq9uKj1DTifWDGMlwfFS9FuAEvsDkzsl3Rel0XQqo3qslyQwdFJwVNrxMA9Qcb0
WErRT/blrtdvQO8KPmGc5G7ktxpXsdXW4bJWTeE7IPgptb+YopZcbTIcihZbvrDy
0JiyM/lbp41DnaNayh1PqRDZkXklElH6JVPAZeEZcySpC912Gx2CIj6nH4POGhOH
uwL2O4XKHiLnHAvrAfgQ+e7S2pLmXzpbbEQieO5JJ3ZZbZhkIJh4MCQCwfUo+h9F
CZ0c1ob742JImrcP07RH89mAM6vY/O/s8Qpfya/cQqSP88u2Ml09BBMxbLFnESgb
/x53kSps3RjkNY52GzToG5GOm2gsXrUaZTNBolPqSFE2gIcCDYslVGopiZogWV65
nFuUP7dSKKVsp6N2TuDRYKCGuUUrHkZm8pdV77VIPl8yySznvefJl6wx7RM8ELKY
skIYBAstA6W+OpT1XrC4j4tsvXoJp6qIAmmefy1ikfyn/K4IJz318VXsJ/hBzlrW
Wg/STTuLlccPHkPZy8z2cOnCw5CPDDlb4ubwRqclCcctFMWwkVE7k2NI3h91xhVp
t27SDOdMhPL0hoIZolzvJI0fHtzr9NJHtaA3LL99qPYIalBR96v/KblRev8VZrhM
DANOVqgcvyiLFV0018MfytmrQ6xYLvn306UE1jHRwOpZlDRTcbd+dU+YVVVi0QSp
aK6RdoFUiFstbFiTtGpXLSKf1sxKvHbW9JAIg/rW5aMzEcyXlZkyE6+eBAjQV3Rj
0gNn19mrK2kdPizvmvn6cBKYcAlKwMpLLO9yqvnzDGXOGuFm50zv3pHmxFGM8RB4
XWLZQy0zjvIA2FxUuXFnEPL4llGQ0tgDZRSumKAhkwOAL+cH2lDnp6ItaeSDYRfM
iVFi9sM5hR7nlZlYpSxPQt81xIxIuXIiIzRxosmL2MAT3xuBMr07OwkXZAdxG+mP
Vp0jdCKz7NeA/ZRsyJzWDP/mIPK+gzcbiedBOQj/pPuReymKJPsiqqvFeUuM59v2
9K+QGgQuKoTXYhPMl+dg2NiV1L8r6OLR6IxjP9lzwnwLsK/6nwy6Hzy8KT3IkVsG
/8kieO2x18JZ3dKHTZDq36jBVssy/0mjCRF3qpqNR9/CbqTdlSTEiEAG/PjhgYdL
HxTDYXyuRixoVYU/bW4tBGD2XYBhY7jwG3WSBUuYyAaje+3CJShVoq4pDUl0JpzJ
CxW8ExEDzHFr7KB8akwJ7GLyNjxQmssixdIjP2OgbP1D5N2/8XzkL1XxZGJ6+S0e
Z9Zl+IcrenGoY29iheAlwhr37HlVT5iOf2dzWaoKespOtLHzGUa3w7qaAROleuCm
SSYnPTMHNnDX3fNYe6INwsYwfoVx3qyyOMrTA179D0Hr6YiH+dUvCgrS/pEPpXzg
R5iNnm87W/cEHQqz+ZqMi2iKrrysE1BI5q7DAGtr/OmCqklBl3+wnR4FrWbvcnos
XgVfemvJciWR1Mp4nxOHjsKzXXYyjLkFZjiKAuhtGUDJ9SXaS1JOMHxOkmFph6Qv
ItYQ/CuAQCiy6wliwK7JenOW5MnkEoN3dBbZhuW2XZKHxcD8pe0WT0Bzw7uW4LDo
pt1AZHJZBdX2SywMvCEj3toao5VmnK4KOi6yoCS9e176YyL6YkhaGKfstl0wN7y8
fDfOmMVyoY3iMw1ae64OJHj1cAudeKV71fXpFZxZi9Yp5SaExMklXNpcCDlu4Fq/
bMPiTq44cHP90ILwYAheZEmKoArOkkxLf9W8dufF/7FN63TZTgAjlfhFUkLx8t30
Ol47OP0idYIpbWNRRplvou3PdzmJPBjVBlf2WMv1oLVi9iTv5kC8Iham1xboB9/T
0uwd4zAmpDpF+WsPIONZ1aiJiY5Yzja9JcaXyGZDE3TyNJgw5hHN+cw9xztYNmvM
+1DmrsyJkpvbwuWN/TF2mekFSgxzdiSJv3PJs16ef+bsnwAd7J2XoJEEC8X1VQu5
4otbciQaWnwiO/OqfqdtowNhnYdCjs3bxzYegPjbGZvQ1v9as+OXEO9btNgtQCjd
7VCiXIH4t9Zf8jNL6GDkLleNMWqo+9dN5zkolCLCvZ+GWyXol+rVcKMLogC7psex
iLCUPQZFjJusx97OZpz7w8WMuZkxoRNSPDJH5sSbBouxJNkCDq8e2gYG8Xml4rnE
eXApc99aOmS4dZYY7O6VNikT91uUdH/g+mDZTlJpKM8AKdJfDJDAdERQ2cLQ9Ujx
E83ySNZD2QL2dKoKuGTD3Au4Im5tKoj02YYXrq2/KbyMm1uCqr3ZHpFBoKTbz58k
ZYCR+XE/zmfrLAy5JTYKBfsIj4andsgu5BL6LCTyB5Ai5zQt1Rt2pOyVn4y7vHMh
OvPDZC60/f1bSGcnco3SuUrFieuCJJdOqoChP0e4t8u9cigSfuUE0jCrkW143lBM
uCm5ZL+JLHJ8KqIoIrfRKOwooHoR8KftpJZvbbk2ePTrN7pmMIzha8m8lgh/ay8J
CcCvdiEjtP3oJ0zaZ6RKMrzzNfcX93MVKgBsU0Dk0z7BMG+MDC7RO0tCxsalS9RR
lFac4EljWIlfcJ+5Pg2WDYZGgF6RICp13iqL2fzEN6g8N/Zd4U0Xr0WiFRGt5hRY
gUBl1csMZDiWc9E7nRNuSmlnZFrDEHbun/YAWAGFA0U/c1YulCucSULhz2a1vgY3
uZCyTHt1KudPr/hqSLm7EjCKtX9dqKJ6o7LbJOzWx08RRWq7WEXIXGjDDMMiTM4c
qCppbu6l1t9Ll+58sfk4cXceN77329OluvmpPAdaUK9UxLLifKsJYnng/JNjm/K1
vgZRbHEWCLCgLd0fcRaVWeDTTU+9RgZbZTBW6HADO1IJMyzIf3UGwnw23nQ5ChK3
S9/KO5WX8gXO54b3zWq0U4L7yaMhXQ0Veg4bw7coBInXYbktUBtectFAlpZrFsgq
0JfSNP57/4oYBdQ2UgErhs20SJiePlF7jDbJE2wdx0VfCO24P1ftDxivSX+2HZsj
t3wKfNWJcdF8qGQSiyN+EgAO1/vi0ut/jmMzc6YcqbAAR0WnDhtHER5/zPmB0Tvl
fWduGy+BDMZtXgQS6RJ/I4/BFFvmEFP56rs2geuqj/eeDxVf9H7TaUkeGXLjCfDO
GhKVFo5rPJSpSUxK+RNIY0VK156jTXRxOcoEqkXew/r8ncvuD6/D+61GL3iIozMQ
evDsDfKru4ZPsSnJ1Wd2Z+LZYRKsbHxg76fF43p9+KgDBKegTh9ztjxCZBoFZhXM
Vb3kv67255aibXmo9Bk09g==
`protect END_PROTECTED
