`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5lzbAREiy7o5nFeZoIFF7zoikkufuESZ4e1tYYNVJuucJ20qnvvvVlqHC7EhzMnL
8V9w/e9nT4zyVs4LLaWxHMkVGb4pppRr9PqndK+kV61PT2zDZ13B9CwC8pqsaEvD
ycHtqfp6AY63/j0naPlQvcdhTlMdm+1qHJl6ca2lGDeSV6ggJpaGGbxW0rS7pCSa
oilUx2C6LXE87uNJLdQCzX3yNeFzglrIlcoABI00XnQxd5//88XEUMo3lBsrR9St
Y+HyuTsFMgHT9rq2NHcR9oTUlZsudcCOoFkwqITRhQIH8p15P1KD/4TMq6c6Lb75
DBcJZSgt7jxt5jAg+t/bAuf29Gvw45E+uvSdjR+EAZcIYVr+Fzy6xq18zW8xqeA8
LL/FKhRZI/HVXEcE3/PTnol2N1bIafL4dyd8VQCMfMFAuWQxnr9E7MBpBBwa3Agp
+TDriBNKKqIxKS+fAbHPxeeKsFQILi+JF4IhgbahnW+/21Yg8H1V/dN3+YM+goNJ
GxiTUp0aV/zoJS+1grYznmbqfapitumj6odpe50ec6HRipxwRFBm5YGDqhlODfm4
dX3ghH9ptTE5xOLnq2RKYiCbhmnvysVo8MhFLi4WPfqvHbmlmJP7JmtHcXoExMqp
oJf7I/+M3e0v1FfMM30EirvYnJ8L/fsMXx7C7mAQKcB9f4mUFP6OnimDB1Arni+P
a0TUlmc72XS/IhDB190gfr5ZR5szqnDoJN49/8/5bDybCAYE1LqBdqPfeu+eGZkv
ZGsFwCgkN2eOW65Y4pciovjP/IVNDsB7VGJKfsp5iT8NWRH13RoycgZ5tX+CX6q+
czLSdrZfpi9KGMCUkKvwMixoCw9yHpVSKgbKsRdMnCS6SIoBo1F5Tx0YBza2eQeo
mTSBgReOSaLS0sYWrgr96xtOwSKkqr6FaKAi6mykcepiqkTsJQ00blwND5VPh1Km
hnNAO49FSW/UZxM0cqZEzpon10G7rAAQyu7khx7u8IFpTT7PVYIbOZbB4Pye68aA
JHxTYqiTFJzw2FUp7G/NywckvjpnAns2oC6tJ0aTy4tau0XflZr05r3xZKQFmqa7
oZ/G8MOHJjY79JveL6afyEyd/i7xJUo0+m4xEuKkYGdLJTAoquCTsWdgsNLY14M9
c8sg09DgTUbX3irCyEZXxLBR9q7pFGk8z0w7/HjhcGLlUMv+q9U26SvjXONEMEHu
eqYbvfqxXHzZ31LiSKw4OihY566M9JczoaIme3sHzG2HoQC+9JofjXTiHpJdz1VI
RQpYNjG2cjmvHNOWQOx+TVgCjPjZ4lYowI7lHwKhDdFGAl88Q+NtuxeY2oK4iq8h
bJeVaaQWumNr8YV9GSxaYJsIKT8391xlTYdRtyO8s8oS63S42z+qr+VF5jUMKqeX
CgmDTQ061Ei/C7fMW0VD8ewxJY8nqD+Up7UbKA2nRHB5sYDPTb9mCOSlAjqhdBDw
0Z8roabIPFTRAj1hNk63WeqSWdfynI1WefapAA48XD40Wzgxbi1x1ylSMi49WHuX
bW//Sexh8mVzmkd5xYpNCek9xgobpc2AioM8ekF4z9ajVPGlobvT07yifPf7RPZM
VWEbIlIwXxg/OD4Z938k1ivVYyKsUdrziciFKZKN9yQv45Egyjh6Qj6sv0D7PUxf
YZBHAexzdYzT2aMUmU+RNdIN476HdXZEqS/djFmPCZnDDtYLSgAWzt5N7tmpl1s7
adYLsYqxuyXm2ptFBQUXMZw1Lz+UEQzBaq+WZ32EThQHiNT2ZUC7am7rTrDKkrvR
991RE1Sm/zWA0e2k2xCxR4vpfMWg6HZYQuggoGWvW/4S4a8pX2L6yWZL+SPnPOVa
bBDAb5XXicYb+5RKrFygCFRSJuHLpdfpFxAfnYYSHDB+ADGwXMkNb9C9JPfyMI8d
IDWxYWcxmo48Uj7R7BFvVB7pinuMw9WUdjLLhMQfjj9MlBVrtTNNM1sXWnhzNz0F
COP3bIYMeCCI30ffzcJ1hxih9qB+t3K+MoKP06zmBQbxW94zKhSG5yxLlHNnt4Rt
ZlDM1jPtj4piRTtPDVazhFC6NwdJDBGDsCQVruJ2R3zPhq1Z/UAZJZX/cnBAGBwh
JF+bXCh8RXQ4QiQN+jXJmNKnnVVyubtqKD6lXgCLFlxK3f6r5I7RfliE4yyPTITi
PkzLzCM3W+GpKCZ6ROU5KrtSJGMkmetpe7b/Z1LceivYX8bmXtnzkqvmAh0TsRtk
KFiWNHqdhvFJWNYXtHQG8YKw7t1/kfFhj7GfejwwveCR9/LJ4pxpnI7rSxCP4Q7z
xw06EO0tJ8G5Al+5fGxEkXJdaEnGX1+TQiUkBecI55m/tKR5t1m18nL/G1N28msa
9gmAUPgQkC/xptzbCYD3MLgqRYaMFPBl1+j8Rq3BxKYMTkuaQIsMvbkPzwj5VQ/c
DWe6fU+ErbNtvdgCVTMicEcrYwyOh2tHGRgx2dl5pW260gWFq9miJswhFqm/ZftE
sMbNvVGs7K2Stnr5nWRtCEnL+Ltw/jUhJOqAtD4LON+/rUs7BShIeDluQLw1C7Cy
rhpH2yLSpUBpzgdunf3LAaU0fC8WGLkoypnUWB3NaqvonyYtyNjSpLrV7aBaqssu
/GJw7bekcxE8ejIbkBmdHhR7qP1a+xdzNCRPkDE8Em4oLpSEBuF0KvC0P225Rn+4
zELk+4MnYwitOg7/gim7Yq2OhHVvd70A61tUzdtiRnwVjsTa+BhoEih/JWNqfS/j
9C61vsiU0QVXhGeyl9Kkg8gw9zmQ94nHwZrUreU0TKe1pbHfLuVSFLx9hJNQozrw
2jaoYLfFRlaPNKBu3alVtMChHJjW8wRb0IIAwtMqHgWHXK0JdEVPkJppGui1ot4k
XlBCWF1veAmos7Cd7KHTkLMwnMfn7Il00t5xNW9+paclwRLw5ZU2QyWXa3Ha8Gjy
Wd7N7JMvsSBFl0N8DfLk4ohA6FfBFVW047nvuqbmR8GCmh1kPPnd+UQokivLNdl5
atQlNYtmqoQRCmAq3gkGELmf8fEHIGFzVH2WR7Gz8PnnccXwxILLgn9WbwAYfp04
nZFN4nYpRfyjmggmrZnA8O5pSrgfyJ7CEg7rZCmrEfcziwzZyWepJ+MWBb/zQJ/x
0BpY4EZzYIHm1E3/PMu7vhr1O5Cw3wXx03Kt1ChZBlSe8+TH5/Dnn68Z/yH58QWM
HUZr5aayOhR4klvLgbGcC5EXkSTpDWJ7vG0/sfR9+CEOhyRnx3nSOZgzgHeOx/Qs
X0SBW148/BiItRbYTeoAA4DY/agBOLx7UYN752HQVChFimgz1iGGk2oK7P9qNFf/
nsZ0Nba8tnRiMd0HqHECefCxKgJANoO2td018IUlkc7jyvejIRo+x+yIrHP/IWoL
Cx2aFMDFO1m3pHt10CpqsgxFdux/3ISWHdKixaJaG68RRz2nRxmmyZnqjuQV3aBZ
OZi3AkUZyGDL3VjeK9hrWywOk8KWVJEQzxk3pJhmbLwddsoVNAIC2TTSGh1lrKUk
1UyqA1vbEqwFUOv8kil5Y5aSE3+WxUOOYAl2bEx28KXkn0NzwQKlrgZR0rodO5cU
9l2oJTjgZRs586Y9l/Gjo2CLPKtJ6mT+fIOCfxgpqvRJlBi9q3RT+lXVjtgsF0tZ
XYzFK7avMmShiEGLW+jPjve53PgZ60om3ulI3CMt5GNKhhe/8hQ9YBbw1lXO1ngQ
/wjTZroEeyza9ptu9bQeW82HhdI/KaYUtUJxEXhCGJKSSYgQBFyrBrmopbT9WD4d
fRjv8meV1kAqZYiZm7Xa9v2FaWMJRdcTsojoZNoHQmW7v9g4Pi7NKRxRd6Vl3YZl
r1vXm9a4F+hC4qUO7rza1Nk96/Hv6QFwQztQyY4NpGunbn2UAxAOaeveXw9yTsbU
9a2FWtiezk56KpcoE/bO/dEuiChY1JYzns/tQ9mn+TZr+SeWo5f38gBJ8OYCJt7m
uPLOptX5Wn0sDJCrctsM5gtHuADICoFnbRwvgtkqMBW+DDK9FejFBEUzoENJICb6
eMe3lqDdjEEtxt+Q9weJEjbJuwI/wWXhPGyiqSfwdDDAtO09fh7KSrLd/aNqMX6j
scSnNZbdb0F/eAh+9Rve+qetqw0P2qEmA4lgczWKd1cxhQfmDvtzL2Z2EJSN5xpA
jRwaVsMj6xu6NMLvLqHevEMl3zjhltbtQEQJwK1kzTz+rboN5iJQyyc8dx+MqqRC
cfkQcwM0TqB7YyCDpKbiae/t61o6bFuSwgV+zUmz940TqEIPRkJvBXYVHfYft/Nn
mgd2xN4MciaNh3/5EduSPN11qFm0Vk57G64evGCfKC9szq4NvnNQ2Yl0YddjR9vW
FuyiB93vy9LFNudbAC2Lu31ekkKH0fJRJ5aXwz9ZLYKpT5sBG1n/XB5vRArw2d/4
FdDPHQm6nJW4q6WpzekoyOYqF5GD29UcoVyy5G9pfQRP1hhjfFTHG76DX255Qalw
N3miawcmmGM3rItD/hZN3/sSdaLRM5V+uaHjn2kWM95L3ySWakqAfL4lJwrDaslD
1IH1dpCYKuRFbQqTJx8DhDo9K2GKmr/3irFv6cOX+f4m/e5wIJQWKhcWPk9qwl62
LH6utbdvLhipB4au2LpVF4lYPqkj9vQA1jFqbRawad/gq/P8gUVmPs4jWttdmRDi
MCtNMFIwz+anjT+/TqV9ftXHyJrxSUWJPdUGgoZ/LRt1wzWe6jYcEplxFEFUmjj7
Rqs9lvZD8tpsBVUcODiSTQlcpnYn8ehQrabS2N5w8bN2+PBelWzROL+l1ce7RdJg
5Np1aDR7TiL34wvkC31OOncP15Ifaqblb6V8haElQaQcnYVyWhgBINEKTcvs3N7r
+kpDIErxYBfPbat6n/B3eVpXnLAbLWlZTwWzthRzZSL15hCGPlMT1Fs+E8kC153j
NRJVt0xC5uYnEwSCTUmexUhhU1K9s2JICCEiz6O1ujCtF14nRyZ8b3Zj+5kClvH9
pwuHVu2uZfeA8CSz9GjaEuzDYOZ1bZDkUaESvz8gJiU04wFmuhPoOWDebQOgP64z
8rztGmZ2Rp/srvcHB7UCb8uhcS3XSMHiYnNs7KMDeC+X+X+kFYXyfbv4Ix1WIYYw
zGWKreVhy0M+Y9w/mO/hESSoAfwh/s7rwc30QA1SFaGln/kmm/658/fXUs9a88ia
G8TB+NxkpMW0rC2lO1A2RQK1diwEOVp/wGFHrSICSm8OgscZY5EjHjIHk8dNA9IS
eoCGhXW0FZLLaBuGBTWuVDhdXXqWsQs+HSgJsXqy9/zNqYvmYeDGmsmJyvk5oept
g38cHjgfMcKKUoxAYTUSX/DlUIS3+VYViM9/84bXWdeAtNenLRSh4kT8kD41OmeP
OJEN1TlrZ86GgMYwliGpIC8ukWXPwHw+H57PN/lLXz/uyXw2oIgyeE3UqBtB2AEN
dQ42UsvXWKRpiwBOa8zYPvv6qcjRx14RdC2ebMfL7zgIny9wAfMUQZyyVthIRQVM
yOBjM7QSe8XGONrRuDWtEjF4CeV4afGUO+dl0TXkb/W0XeLM4//WNmd2s14y5U6n
dVxiZmp5FKf78cxrEgm1EMGykh8A9n0JV+l+G9wSCIphOsYP4n8HXVxnl7Ou3SM/
+KFFrEgEqkyXVZsMD++VtZsbc6qAgzWEuSBg9A+J/NThPobOrSjLPPKof8wWx4OX
w+yPc5lC2ar3ywZzkXrbAxcEkOER2qKrZm/rqIGY4Trppu7gst5nytEEqofLDbMY
IqOzmq6PTh9aotnegug7WK76MblJnycT4NrPfKPU5Jostj1DmzTqd1J6f/DEyRAs
g35MbTBccsOjmhHCXe9fqWGEaU1U/NiKn3uUPRjOw2B3SRzByd6QK5HtJ04v/zEf
SZPVcQfbWX+1ouD7LbcEj8iFbOXX3Myl1wv+qsKAKBW8ooah8P/WZyt0+PJSirAV
DB+1lWJOcRbyhY35OeB8NykulC89o3gbxIr8MAHpznWmYtV3tkUiANJmwQGDACMb
dZw4nlj9sZcj3nicw2X74Fqhkv77S++vAT+bCraKFkQrEgAKwSLKCWBwdM4BUBBU
WLsHw/GaKdA56fW41DfB7G+20LqKFRBrLk8ugKyALK8/Va1a0C+VHYnxKVuD4hAw
+Kyt72RF2slObNxyqLxp13dArGEdxNSv1+o93ToUN3ngTg7HbQ1nfw0YCyzkiao8
7Q5GVNe20AxVdK/SCuqiDhv9Wpd5YnEHs80y8mmkDV58vzIIjuSrWbUw9u1mdcBY
zF+MDZVxWQs/j25HEskVzEoqIw2ZlBJ239/IT3PP0o/E9voDA5vjIFE/mvfsyjPf
chg3NA+R05jc+8+4ojkkGFWW1omLx1ZxfClImwODYB34TGlXWGFq6oOzlHP/OPI4
4uebIwLcwJ//1I+MCY4fpxRRUkZFrqPYRylBX1CTKfRG+BtpIXKT+oo+Ak5eTMKk
shItMim7xL3uCU9i1KypAwTOJmVpYkmTadgCGbzfKD7d6qNA9LULJlSf6BbN0uFy
2TrQEbeB2vo7m3FjUXyj7LmhFTwcRwmtHD1ncCI5/4qOnNCgpaGHkoS+pYUuIIcQ
hidrUTIT8ZKjninKFyg/IPuyOeXmVLTZ0zPxysgTgycf2FsSoNI2ejIRb+CTvB21
mHMGYycAoeCjn7KfiLzIVkDaFk5GqpaEYDYVgS+nb/pksaQOa0IgS3Hx0YBDo7Vk
VC3vxECZgLywjuMEMpBPBeCQD4ZxTqxer1Zc0h7HWOR8jPBDWeyaadjkFm8CD51A
p4MIg6l8PEiRSgfq0Vnz+cIOq9kOwmhitSHAMSGTZSiwAg0rsNYbSbv/UZWjKP4O
d8Npv37/oaMw0eFYDnNY8Wer5B0cqyrlTYQxilnZxFm6fhRXitkdHrHa3PR+eyV0
M+a+sdamTWBt5KgEqSznZE6oGt3ImzTGhHxrlCUOlCQyXXDK40k8U9XfKyv1uxF2
mJM3ohC6flYpS9cDcnLhqfQTp2lU87Yd5cri+SaD8GgPhhYXHC1LfoVfG4Df8dHg
MDQ1R9AEOyLfQuCWdslFZQXsKKEmUZv2HUw1yx/Pvv8pwRtkOHgBL6yOERwZqGwi
TcYYkjWrmsBt0aWECFRZGdxbulYi35X3gYuYZN0R9NxQLczh1iNYvLleMock3bEl
cofhDuAaGjblrmYmVmaMfvbnFIDPq4fZhUSO49ajrkDCylQLFQB4V9ICNqzBIAHK
sKFoOhdgX0drEM2ejtYsrje1j+rHm2od7rfGX1iMb+iinQ+pXH6M/s99vL3bxE06
vV8otP2H8AW8KtE/RrIpkAjp4q06M5TH4rCGByJrXtVHqMa6LbeqqCOA7utAt0dP
`protect END_PROTECTED
