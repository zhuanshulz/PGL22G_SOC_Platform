library verilog;
use verilog.vl_types.all;
entity GTP_ZERO is
    port(
        Z               : out    vl_logic
    );
end GTP_ZERO;
