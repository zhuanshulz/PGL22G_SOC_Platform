`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kMmKBBOYfcgWCAuL3lhOLgqpc2FOV5p+/SqrEV5aPvl3peK1kVC/N3JaHJay3dK
m1aKmsfOmRljL/QGWC/iBWNESuUmfleAsm15p72hzrxW5n/Wo0SU4IGt/Idok79f
GsQkUbXNwCaDdPmHfrTRWcIHlz9ZghOWSucjhJ7fvGtGzCQoI6CV5UsaFsSLEyrf
MsZdKjlvwqDi9DzcXZRHiU+I3LTUMRNUp8x2fV+N8ukCIPII2hyDkW0OEyEiMVZg
v7dvQfSgovWnjk0DcexKUDsjJTg3zfiouHRiRaWG39XbtWi9DDo9PHXMwkn0YwbL
CgZKbEqOZFNHGTCn7PCRcgdRzU0pxM5kgaqCj3aLQXxXtkSA0GwmcD5LEmfuMJQq
Txo0fe33FvaWYMTELueG2fArkfe3Gh0klnT+4P19BbmN32hJJqHFxtIZc62VeP57
DZngTEVboypcS77/AFh+G6VnNSLQdjbNu568jYWAWcjQkXy+mkaWhVhR6PozEMlJ
r/jXONfYj7R8/zO6+8xO9w==
`protect END_PROTECTED
