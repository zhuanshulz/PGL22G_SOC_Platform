`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ygMM4qG/mtbDJt2xjqBGlotQORlt6klnlf8BU7Ha0ViXkucsAhU1lrIWw552ZSGK
4N9VuXBucI0UYGC19U/nqgq1E93pVG1C+J6R/WNcpBd05q9dU2+wDXLDjDAvuYdL
x8LIIyjj001z8cOQg1Dlpvtu9iNoiiaXS3FNXuPSMrJQ0R0pZGQy7ESWRvFP1HDV
KuI0aEnPhsxrraARWqKOHi7hC/oObUc6frkqpl51XglyPOBTKnRMntHFijjr98/S
cWcazaUNSL+kHr36jpy5L8KhJIjcqc4yvGfLw24RrJKs2bubTBdKArZUoRkq/KZS
R+DWs5E6h9j9hpm5OH8klVWdFpxVRJIjWyKLR7E8H+06McE+4zz+DHUDxCeIz5if
Wal9qJ+MBEQbYbxolyoi70gY6ku7Wc87Y62IIRqAH29SwjSuJPokdW1AIQhrE8EI
WTjc9suiNUEqq+zhNppFtjvDMShX4X/TUbpcWzKsZyux/8UqX7FJ27QuBeJkejsO
npGPk6Gc8YOhwpZhQ2bj7GH1rIItZtvH6lKNOrDnFI95ss3O4p2acUxPtvxrGo+s
3xGQM+osOUsV4ZEOA7iI8OaNb4MgvkEijwSPgXJ788KNvBQpAfvyFh5Uz5Mq9qbH
wiMQ/wsWrAhN+Guq5gnQ7GWn/Pvdr6ezc74Ohn15r1jG/y4nBsismccnZOI+/qww
lDG3NfDvpCxYQ8B58aT5Nt3uHNKkI7zMuv5XqkL3J3W9kjuNe3pKFhw4HVoJZvZQ
kO++CLozYtfK4rBPolbTxE8TxXP/aBP2KTiIuVDmIioF/M5b9zYkNTawsB2dwNH6
/pbhjnw1ObpyT7/hAOrTO5P9sESUdG1r5j9zYJSw8id9ts3e4V8mG6+p9zMQ1nbk
mtOJA/oXjd7Es9RVDV/gpuDT6ocIxd2a0em5xqm+Q3G3wwM6R3Jcz5VjOhC7qAbO
pOzPxfvvxs5H2THPEWYshRN+1Nyjcdc/HjFw2MxhyXKG21T7yEhbgYLyz8+z11I+
O4CEy1eDaigtmucaNRz2FlmGQUavFARfTGLbqZyKyRfyAb8lUjVdyftj/NgiTZZ8
pMaVyxGs37BBw9L9Enqqq0NuhsDn6vfiO/SYONRD3lI7JGzbvu/p+NfORVH9DXjj
fLVa1uKniGIApYFOcI4Eo69UYlwwKKXX+y9gteY0dUdrM6shdPof2N0MjtNjEzgp
WFUnS8UGr5cLCoXfspLwKuOjHkpx8qeZeYLtVSbCjei9WybZ8fl158Luz1vlfa10
QqznrxdyOjMVaD0Hz2eTfLcMDMnhzijMELR5Uvixweke5nAeyE57ohOpctyGtOax
25bg2s3JH8L/V0QlcoyAXm9QLPPE9npGjvyM5u/ZKhe/hRUe7Mdj6SkuVvnVD9DM
nLdqxeP+zekZ89FLfSk0t1+b+bw4NU1Oz8pIMAA20UXXAqMfsQeTbM4t/gO5jfSq
C/i8e5mYsCavqMz0G2FwUaB85o4xrWqirdz4T/2g2gGPFV6xIMR32VIE+w/XEFFX
zQLPYG7Qc9SeJ3QLcV0mSKAkw9OOOppRMQgiYgJiR073OcyXH44UfytUz5aMODmB
dtPY6BT62AZwObBjDR1xoricMmSK72nBzp/MB+WBM9gdUgQ6MGr2RAUbMua4xfhR
/0fNFyYONUnUK+e8QwCO1N2dVUFBu8cFGCHzuJSnthDAZYRzBgbi0PoSA2LjVXLV
OAYEJPLen4clClDzPpR+J34dqHMSc11lBCNae4GLEO6rvmXYk6M3aNigg5eGLTIq
LeiZfsThVMhtgeNojkTJVshuF5DkfUBhtbZNlZ5lHhLHhUFs3SR3U1s3Qi2f1IK2
EFXOB95Ma/SdMppRF/20poRtIUFso0kK/lIq53t3+vTf0+nFskXDT0UacdfnAbx0
IQXwGbbi+ReJxWraZ3X/OVS/JJaHqDWRUudoMuwgSqmsGapN75HedueHKubRnbX5
XwvNAkAUoiUfv5zblLb6siaCYY1iifpO1ceymQQXj0YpOU3yHBAxKGcxgAqEj1gY
vrODZC7pvVQiwFzxHGKhHAHOaaBXsoNUZV0WzFZGjEFDw8OLeM7Um5JfwfPbtjrZ
z7KTfbPTbMlhJf9DQb59UGJbPvtIVg1pG58JNH9jtu18Z+Pwrs50CoaSzP5iv1Ks
2Zkid8z8HepnYQUSxjXrTCSGpDjuFmUjB2snZKRUlQeQOjsSI34OG2fUJjV3fl3f
5Md4MiFe+FyO1FHSOuKHeGdsO6/e39V+zJpaLgGyimoKQQy2xnYlYcBQqLOTfmwX
1TLfOlPVAgNV3xthSea4tkmGcGrm4SWjvl7XdzlL6jqjtRwbQcsgWyxB38OAzFTM
Svt5prcw0LvPogPnJFzRWrLzfchZ6srge8RNbvX2DQFU1n2QiWHgB5qc5OheSozi
UhISE5NK08yNlJBF8MhcZQXnW5iE93KAKCfrxx3YcvFrnfDEiQpSnbe8bgNUWOYZ
oYcvK4Ws2vUQMAI4mrMk9TRz3WqKJ+urMpvtoOFYxT1zlLkqNSWe2B9uoO6SqJYK
n+qeISZD4TsYz0nIq0Qoy3fxhqWlke4m56X+okd1zlve36T9kYLllozeE/y8Fnki
TDQ/29BU1J3rLUCNcWRUIEmxwTeLaqtLY7cWaNrykj0cAGr73HGpyeSLXnhZ14Jo
aUh1gKbqTJrYYV1ViV1o4+/UOr3WZs8iXeJK34k+n/0=
`protect END_PROTECTED
