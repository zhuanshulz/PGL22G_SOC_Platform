`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ud7rwtSh4xMP7D08cp4/KGqCe04Flq72f4tkM890YHj5w2dlmwE5Os/H9X6Yrkr7
HI+UPGuQhBzmZRwUybwpobNIYhC1maf+DMhsSYcY5KmcpQkZH6lH0QI1nn8oa2eQ
CLr7TTW8TKoE8aGz0LwsRO3sgaD8UL2EJt9uFVXQPJpYT5rqQcSco9zF70b8TtFt
vMb4xO8DLOue3Eio1g79ig/fsp2AvOk9gW1lzAqxh3vGzFZI8Be/tKNvRCSNU2Dk
0UIWpy0NmwLyW8rPk3BQDvwpc25bMA4K5w/Yg40vc/4DvUatE7JoUcW3Haq4Bnfp
LCmnYSTAI/649W2TnPwU45lJytV0bhQnIK/J1JUsq05baLVy9NVpNlMnCbgzUcOR
afCVPhuCPZJtBYSqp8TCqkW1jarSZx82bHWAuqFh3EBVYrwSAEa1JDMYtxPsb1rQ
nR/loun6Wl0B8lWZlS1IVZ7e5j0DDiZ940CaOIGfdj9onGBLSbQe5dTlbR98xjbo
1p87evz8TsbPq0p8knZawbki6EiSHfSWt0h+nh0sduCDi4JZFukPx9hFkYTphUQ7
9bbbooTQ5M2BXiT1VLCcA6RPrWcyOlcdh6qWLsNnMUsJlgz1u+gU4G3EOCx6zHzx
aH2NEYJO8mhnyVUs90RgrxquJAUdO91MVNU/rpGCvbOo5CQq5XS0lUhs/RUw/58q
2eNL22Nr0lS346RhhjemK6Q4Cyb9DA3x2OSepl6ErvBd+vDpPgQLudmgE4YOyh5N
`protect END_PROTECTED
