`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IR3Qpajbi/fBg5btqs4wcD6l/RNIR9oXQls12kfzcgykDGK7j5/FxUZBq6f6iWlU
TFXjq5YwaoIS+3zOa3e4FlFR9xQxG2hbj3nIr/ENGp5SY2rq81rSrDTIIUFVvaSZ
rFqh5tYsgTQLXdRWmh+HHQmZWONkI78Ep6P4QQkGzbMKpVJg5DM8L9mW8aORnhPC
0vVsxCu1N/29uJdl1VkT1dv7x9o5oIhfpuwiKq5I1ukyTSjzKbndJpH7AtI61r7R
SIytQNRrAAXnp8ps8zF9DwuQAysKIICpQXsYjbf1bJr/mssvX4/MrL8Ur/eyDuTy
EdGtIn5hMY5cF2L5AKgf6eZU5jROb7qPrskjm2QsnK8aRJ0MYPJs/DbDrX9m+DZz
htaytt7sy8A0mEgPpug6loVy30Rkb9CgpFDTluH9WMrNRX5dok7+ffmjWaWX883k
qMoIcaaqmz2bU/1wkMQpLAwBUiJsI0Vjzv2FJv+4CGRKVcr46aFNLG/mxpzGfo/0
aECtVGAIXScfKROJSxhd93qE1ob78inIdDmbYD8No03NFeqLaEsMU1QAGPTOkov3
xgxdJh0DrVplg9TOz/Hvj55K7FXRMIcDeg0bCUvLzucvDwUZ9VLcdnsOMeaspgft
RPixRswHq3b9gKdeFEnIEvbJkxT8N0enlU57x626+EbTxP95dvksnMT9g/22owHo
gNDR5lkm0lkaIQxbVszuPrAsmV6r0jxeWfaAqoLKl8gx7qjdHXqRioIu5dyzb7bh
tZzQQctXxWClWPei3jzLSasCFWB6l1hqLSM1FiLmOc0ei6p+50+vWwDeNyveS9wy
j3wX1RQcuFFFhI24t64iFrAcEmqr83kMWFzlFAxt+KJCgNd0/L1VQ7ghIUlcFEjC
z5QnsvwXwgWEhTY3JwXSxEVF97wh0youNOQEH7C2NqM7ZMurzTIY5V1iawuroSmd
RoExfbv4gNuxfraSjJBHGw==
`protect END_PROTECTED
