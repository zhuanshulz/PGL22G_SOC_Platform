`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hxVU/Uc2Ncn/Q4GkWuSYNv3HYJSag2mUXVOLj9GHVE4K8lFem+FPBBG5fv06tFJq
LhieKFiKWDIgzR/lUD3lFPZpR0FXpdssdtIeCg+eUkH5MDiNYAS5I/CO6w6CDhMb
R4lm6rrGVZMBqLFn2m1O5TLOva/bnTD0ZNd5eNaLFDVVpOxRfvG7IIuHJysg3r60
CTlVpUAyYtiBtZvSI4xgySXVYQiJaGJWV5hGRO/Pm4+rGQJIQ6OYYSNr1qrEWlU3
BgVvo+52o7+vgc2on42866MUcHmdsYjrqPi5vvx8riVNlSJnRAHVV49pwxdwITqo
8dWabuxmif0UGvu8xeiM4Ht0bmANVAyvBpN3dWQqP8bZGCsY7cGLGcjvz/T6f4dK
HhmcgCDChG1EgIKvQCi/70bVMGDWdMEZG5Fl38oI5aWdIakPkD+mlwFqvIwtLFvR
w6uMtF6p6AO2fBkgd6kLyvuvmWrFTP7N0i4DD1NmAI2C5IAm+qOfCGz5hvDdU5mQ
v/IWWv6YXWSFEebSu9y46nLxb5ZE24nQ8uA9dqTWqHNxoLw8/G7OOWcrOWKtnX78
xe2O4vN/AZ3bwOyBZ1NCo4z6FjigoVlxvDn3LvZs/q3KFYUvtuWXpJduDCFsJnTg
HBCqqkyFppb2ShcE6jF1NKr2R8JscLkD6KPSRh9iEOQfDGTgpGxw91XfCWOa2eKU
yXWduFZAa6UWuzlMp/H5Gziw8kVjmr0ow5gjGH4DajLejkrpasGVbzC6fR3Dz5Xw
2pmj83JjxnV/JZcajXA+3mD8ag0TtDEyqfBmK126lnTOl1x+eMHiVOhG2+7Jt/lz
4rVDfObq3x6X/hoAaczCvkvB6f9j8lgULweclr2dDLW1l/LOLpXctaMslXIv5zaI
7nnundkwC49o0LWoWXmiSE6jsspdk02dIH6N/y5RpsrwS53T1efrbp1Eydy+E9Fx
eKrNDq20DKGwM64lfgQF1u/OY7h9dRyqF9bAx6LGdMmDzVVAL/Qk3oZzOWWjqa9B
1YSQq9NF46fc0qY7ZXicpTHQGlAO/1PmkDQtCg6OIfxjPidHYT2hGosH8xwdyLov
qtJravSJpowfsE7M3alZoKfI7CwdhWvc5y8Yn68qrRGDB5bU+JNMbhh5ve3/88Wf
yqgTs9S5NerPufioA/QNh8Tej5u/JMsK/C1WHTc+KVJyLH7OiZNfCoy4J3DAKMyI
dCCbOELIU0wq8N9wvxG0U7dbqFRMG36mTB4+gL8PdVN2VTyycMWa8DccocAIpoPi
bBP+QgY/Kn6m/taiFbMssZr6SyB28k9Jw1JYrbl96D6w6HLpyqQkGz2lVuZaBD3q
xrGO+7iyp4HEvt6n9GUHLZbAyvXXs6zlidrH6ZzKY3htMameH6taen9LWvsc45of
E0PyMgtC7Ei7PC0JWMV5X7Y90tLXuTNlnmpeAVI/QYLcsmP+ieFv2Aq2XOVPl1CD
H0yeeM+VK3sjh6nBK6Qd/toF4xE2gdGCEFmjaPs/5OxKwwq+FQMkIsYYoqF7sLIy
esqCDc3KBoNXA0kmc0zHcPGU2N/Vfo08qMpYTcZPOSffsVJiPt7eBmZyNt3J6DVc
Mi0SOcpOvYY+ssd1M/J7MFtOKe6sAwbrboTs/4GDfNuMDwHyQCMb4ZGzXWJqOlJZ
K25B6kHxrKpwQzCBZPjbqa//MeyrBXXtATWCpJKlU/Bs6BIKWgvUOkV0r/CUlqe5
I4npb4B99jx7sBLgzguBHIvXdVNo6CpXNkQc0CurdrbnXZ67E/PuI0YOmCQ+C06U
oMofn/0YVRP59fDisGPLr591kGIFBeZheinT8DLZUzfkNkhIKLT41xMzhpKM51Tj
SNLVheP6jIQpLydxG9f8pKUfno+FxFCRCi6U9+CUkvA8aYlbhaTcEDvsk+VzKCSj
HseDfpb693oceh9TxVoVFnPEp8hk3i4Hx3/h9ig8vvaOawO6BwyHEANlUxyZ/po7
1t9hPzhshWJ8MMZK1dBl5cSRbtVyye9tlXqdFr2hhc7TWr9CuCofoKbRlTDKoDup
al0CiqYwCuVtsUEATN5OtM8aiuFKKTM4gsr7OjacTEKEUS2dbOZM7s2Vhp0yVdKk
VwIHWH76n/zqTFpKt8m+7aCbYhWREshftNikIAWUZn9QDPlDyTJ8jBguw0clGPW2
sQ9hfozICm3Tps3YO8hxPnVCp05I6TpbIebeViSlPyvsfsZakwhZd14ebDKq7HVh
52aiYw9l6SnTU7hx9tQhSMQuxxVMCC2iE29jQNIjgYy3ZM2YYAqYrp4W4A7GZXWH
REKSZgCjD5kARx3JG9AY1EWD8D+Ku62Hzo2HSuY6UynLx9uimkGZM/b+jBXFxLS6
ZmsrDYj2UehcoeuSZLlF0EceG5PGD+VdL18ZKiqUPhlU8OkJqKM6uphLuT969Y0u
BwQ7JdhGGtRjtQ/fOx2kknClUBwoJ96Ui6csXV9JWQt9sh+LxL/TZdIluXVFhwb6
mCsSfBQtESrlAsxW16gRWvTmWvXNxHkU2IylxS+CQMpONzS7jVXMcygTPwtUbM+3
l9AA27BxPkqSa2hjyp9TcNYwZq2/KpBv/xCA9JRdF2evXOt8WHVqf9qhRjxd8Sh2
ungEhOGzHMewuoSpT4vpzTs7jAa+2WGyAsJOy5i66ToW3WbSzzzvQslLpjLHvat5
CEvASN8S2drRdhgWEMAmCmkMnjoXX0N33wlsP7vv491FVfR4IWBR5rjZU4HoJLg7
sj87o0qwTI+QFLX+5k6CT2KPUKANVoeeS0IEgxPfmBtnmjxofOrD0BsBTvq1mktr
GELDwklEzgbTHZ7eiSd9aHhgQaqluoX+61nhmklnAW0gY1DWAPIjYpme+//m3Pk1
PnryLlC5XgsaLq8QbiTgiaAGaFy8Ak439J2LFvAEToWBoCTEJdICF/W6eB8MkcjH
j/wHG7ShcQUUe9i1pIrW4zW/Wg8lxDX7cJlCfKMr8DSh0t9xvUg21hANnKqocksA
pg3uHPHHu6dwZVN2goXq1OrXd1yRGOA2kDXaDmInexkOr3fVplJlD8QZNs85MnMa
FXESH3STUQnWfkI7AYSD0CT7wyC4faMl6S7VaEpgq320+qZKbI3FHFJATIkgBmCu
ugHVo92TpyIfmY+0LApEHXYIfdL3Kv2/OdO0fY8UOIUH+xT96nRsgFxbgT+FBdWa
QuIorMlM1Xk6eGRMQSJteEqDDXZqc279/dmGoSsmiivL00+IdDoOAJuV3G9TmSqv
N+ZeRKtdE4ZZfyNZkNnRvQaDwrbQLXWvf6L42562LR6qisdCIaCEpkGe0S9P803l
WJorvZ5FdZXpcDTR9pdZRm0Lgzo+2V2MdQJCiI4V1UYX4VAipqeGhEzgi8ivQUu9
j6bdZ6yReFxWa/qzP69FV4j73xhr9xLXEmYzxoXfpYxbVhBvr5VEdC2yihLXaZl3
DNCasgJK1bNN9tyfIfv5Dn0HXGkt660ybaYv7UYB58HSyTQqsZuhxcMY2Ajk/Xxs
ZNv1wtgE0hswEABeVvR01EH0ZERNbvMhjC4PSJ8KMwVqTTTHLYLn/5xhX4eSyUhv
LyokclxEaaPBjuckodLoObkTlrcUwob0iE7Q8SntiGC9EB7IJ7DTRxd+8KI3HDW6
tuzBxmim/82CdfTA0gofXnKCRDL34oNQLPNNyrH0UQzKne9CVYaCYJW3aOMM5YO6
Dl6BbKmX4+M8JLgoD2GpaxPrb4xjLA1rvwlvZ5PY7U/knsh2Dtdrd5hh9m05YdRe
4RDMn7Qfl3SsAYTrHDy4CAPPwPMfaodI4nYWgAS6aO0eGIIBhZOYV6v47zscqG3u
TX5ai3hf+rGUB0Au+5Jqv1/kDQJDIolR6Z/a04wi5mKyLsfY8ESvlDQ8gvasYM6U
ChaL1JoMDjP6sFZ1Z2JsD10gs7YOe+Rx6Q5Ja0Y5x7VLNEzEt9s8cemYtKh64XKX
BzVfhKsoK8PTdiKZ4Cy7mWY1IhRVe4JggM3NziIflFwDzg7KhxEHJLtQE5vp3UZu
APy4e7rnC92kqUlsC1x7kwgncL6dWCnkL7xKi2fCjPAMrGK5Tm5dYo32/6rtpTd1
K1j2LQJbCn6AUwUf95VdOTJpU+Gfj3F/BKG0+ySpu8Z3Qg6mGH9HUBr/FuT2W3Sd
q1Q9Q+svrWJw2AiRdZUVi06QEKGmYQQrHQlaVS0NozTXyrBG568RYwLrGol6FHxH
8mkw2eluXEyi/NnaO1pujTTECo45UrEUZB3IDN+VLdFVBbW7FzH4qviGFMMREdwP
qk5HZm0ak8aoL5DNyYOfl+lcBPHL8iXE/J35NNvTgabuXC02UbgWvoI7Sj4TGwed
POXbVlDqy5q4h+G64cQkbJ/SS4Gl0ABgKokTAx2EFlFgCjz3ZhXlcIf+R2q2Loi2
fk1MuOdcHcneWnUf3rlnvvuAs6JGkbme3dO9XdfcFWMCnlkqkUhrkFbyaB7mQZGk
8Lrxr0cNyXFI4+Xz7xYsw9cNPb+01+NodYLEuzQ1cn/qdBGRYQTfy7/SG+xhIaeq
5DzaDBj8VmdTZl1xxfYtxlj+qegLWZ5T0OulE9JQ0uCieYcUNj4Ib7VVj7aH5FZv
F5AWb2v/gK/CdYr3M4m2Np0SPZm6mSAzmSCUgf5K3y0irII5k9GL6r7EILT6oSIv
DzQ46RFK22dstwuUaiJ0ZyCbcFdx4RaU+x4urTjt5PIflha+f7jbHiVPUV/W3mGM
JwMolmfQt9WwhrEeUuGcWND7/R/xrgAmUmpA/+yli15vsEuvQs6iW8RUs5SqWD8k
JAnr6H9t1dq+7WHbZ0A4pBdLITt9DPSAxO21emQ51ZeQDGpD0o/RO8DSiv35hZIk
dJY7zLucBVTYNW6E446Qe9zSDU1GDMFRlS5KFbXcWmXWglQO92fwjr4H/4/rlsti
cDKovgeEmnoOETp7moK9gZwbuSDbvcxg+NsJkZTup9glz41Qns5wfaJ5l4OcV722
zcHDCQRFBrVRCMGDmhqJxdSgP7SC7KebV/d1SY1bBUf+RWSlhJjPL4Rew2om4Dng
oiF7RF6A0BFw1m7vj/hpVEOCddpGkZigDoKeYg7OhrRRNRfyM3JHeETrT4NX7P77
0f28Hysl8GGA0ClMGCscYI6WFBB/+dJcuvAbp521cmhLo1/PLMKMMe7qqS3zplQi
A12ZgzQrdAEDgt20i9lfEP7kxQU69AJ0A17/MHgBQ7bDt6zAXQOYO2PJS8rb2bAI
RK2gVgIwlP8iE2TEOTTr0P55k7tBRsYnUHaFL2OGGZch0AF0ch1GQSWeGtiMoRpI
3wvK96eTSIOvTsXho9HrhbUff2tyGbXdnx7tYzxiD7sJLWmzSNaQHdgMkhH72+eG
gro/nNY3wJNe3OYfdIL98xtE60pP/RcZK8JhQbu7YV01k3lKNQRof7vFVWYDd5je
7XlgMvZrCN7g80ldO0lh4n7NDtrkEbv3VXVXLJp3ydpupGJnGnmrwwz5A3MB6UYl
OyPQi/u6WczHghkGmTV+OdaRUBDmRGcXclTb2sQgdGplRTi/xyYvJEGo59MoHX6r
niYEhS4Kvo8u4s9TZzcvtJg0BIgq/N9a+OYfkz0UvhZAWnrMO03FTd2881hoe+5L
prG+1SnC8+fAggokYf9WFJI0ntfxiV5af3LoGb6Fn1NncBvdSa6LwUsrgq2dA3Lf
UIYylU3tj+MlO9wIExlTPcSbvUrTLkep3lN1BZJzMK+Ok085vllhPNY2EiZUtGqP
6jtLajWGJ/4H93RKHNOIjw/awE/T1xV64c4LOG2Xs+yiYrvMbMnmGVMf4Frq6NP2
6sVsr9Wz9rIVOprH9MQeBQfw5XEKtr4xCg9sVEDbsP0sTail/4fFFVxk9HFuXn/V
lN3a7JrCvYMPDHPu+TVMjG/oEmSvWnsnjrXSZezT/X+wlIDP2UtNHE7Qvls8xE9C
lOr5z+EFRCay3h0ATyi4jijmp/wWXdxHdEb+KXLz3/ML/5PTnwXrw1irzoOTRJCJ
wPN3UbDYSfJ1AOLxj5RN6S7udhFXobzUlmRKKMZ9Y3XnwjpP6zCRNSFjN9MFuKX3
/cI3xOG8uVkMDC6zhbOgyB0IEEOCmnFKVZOUFtJVSoyXm1N3viXLGARo0ZHwTsPm
KvmhqlXWQ1PaUBNruRoJyicmVrbTI/m6BWdRUnAc5bpPx5FcbrOLdOfjBuXfEJ30
pf0uhYZQ/e5SRCB+XtCFrtd9MlQ6n2poXEANUadQtroVngZf4LvmswDpUsBZdyJu
MclHykU4LL24fAj1/4x+ZipJ/mjkCKxPtoeEbDsJLUQgpu7It4Zw5FVdt/Qb9JAO
TohpYaQQ8zo4ReEFHDNwUFlg22J2fEGRFPPQPFdMFNOm/42+Yuh+fhOxcHqC0I5z
q6j7KvmfXMWqv8f7e8HKHOXMIIYSMcgxqB12pYs9SmRj414iafoNzpjcRvsVbRkY
L+IaFvcFxJbsj/vOU9FD3gDYBs7lxBHvMgwnvNx/OcLLNanvebVB9GqgxFttZApH
n+r8b3e4y1GUVPCU5O+fAIuShIIb1KPz05JJ9NLezJuHedlYeF/gy5w8UFA6MOTp
lAQqPdi4Q0+vmTVTssEzx4ST3v6N0VB3pOz9So8vSlZH9n7g39TzPdKipkUS476W
DuOwsWSMTcBAWMfVchLAKF/Cvv7haO49dSr1XEFS1p8kXHHPBqQO2c0/VzoceiAZ
8+zw/4AnKoBDq0YfxF5WQ1e0OULbakpXJ5BgVX9PMmIbcvKsUX/OXEDKL0vGJZhu
KOsM3yXwtEsG6B+RmhPmXJhV1EOeKphefhrlzWdo+YTBtiLwvusme+/StUDfRBPE
hCd6CqH2XKMwr7YMDsmwmYN4AiXDb2j5T+3EPX7JI5shoppf3s3L4+vogN0oYLyC
bylkmcg6AWn0RwIm4onJ0PnKgaHpORuk5ST/KqCd25NS3SRjt+qu+1Ikc72Lr0Up
kOqBViGAqJWZUf+tifFjyOPFY72ixer2cM+dsZb+oRXbGqLOBdY/CqQ4ovHtalM0
N/rP3hL6jGB0K7IivVTKbRbz2eykCAZ8yvZu5agz+zB8qXYKa9PWa6sh1+ta9h7e
Tsyp1djEQr3NZAmANI4cyjEyM4j2qvLCHc35Z5bmBxcm9L4WgO6vQMm23xVxpCmb
w6+6x7b5lwxR3DwCXueCsWTr+s+NaqWu86hFMrhOVFEphnQIEulrDUmd411AxslO
AwCYFP51RMhJZIu0yMTfa5SDsIw4b2dd1IxH4tUb0ii83axgm2Lqjtpmy74fvUNa
nAQP+tNY7jd3d8n4iv6NzPzpP2MDIlOvQ/tfY/fOaf77SJH5JYoJzDy0IXyNJXJR
Mc5QWge6no4kWZryBchSVA77rzqXmYbRRBM8oAQ1iAthPgRHGKB2rdzSll4ppYHQ
efxnbPkC3W4UvWfOlbd5ooNzS72wdYYyYK/q7OQ8xuYLk+X5faX2wjoIv9VJY8Hu
l7r2alHkMp1u+WPFXUGJJPGrdJBuoVzMlA+yMIWDDMHa8QMqn+9zVYQU1FjVvIBM
i6xCeybyCQh+4WCQfTaEGA+lE39S04YPIt6pM85WPAWr5ns/nR2n1t7CHfuj5P3C
VcvgSBGPWQXb9wmfFmqK7J0rrNIFAKzPvrTfOhTmxV5OCrd1NJV0TqjtMcmWJHP/
XG+9zas8H31N5+50MEA+kl+qLcW6vuHTKmFB2KZsbLf8tCq60fM4blzwxkMvtUja
z6kTjKaQVD43o7614BoZX5x+xy4km+FbbmrH4ipDxFLJe6Lxrm2UiUq7uNC+NXrz
R83pEbNtLJq/ewugwXh6y396/LsuehnVieYNdsmbQmQ6Opq5qp2XLF3tvtKqQ1PP
FpxDJ9lyt8q8/caITs5xTvkoOKcYwF02IltUc3vlaDj5bvN9+n72Jh9GttA8Ksl/
Xvdc0wEoa3PZF3py+At9OzYhbrzY34MzgprokQW5WoIinaQ2jBEdVE/niHtGNYuq
75CTY5N5EkddNak0JpnGheHbZnkkFRincTBib9czqCDz6dsiHotjFLW0BM2yxAt1
DKuSCIlKaeTtDwSyCNNz3AIZNh49HyGerf1wbNsXlvyMwhmDSy+oX8D82zQRpyru
DfMqh+XGk3EZuUY1Zvt6Jt5X5STDSiiwZdvUsOkBRvB8UcjOi1SMBRZ8T2DqLNf6
Xhpprd1+cvRjL4gu2BbpPWOBRvagFZZAC//nTk8rNmjp05nIAGH0p57dw6lz7/Fz
K9SVEGsl2/G11n0TofrErxc9UtJVBr5IDRBif5RzaBOTpCPS33X5jNf6nLK2sPXl
hoJ4hCFP7pHyzdnr+h1UcpEHyQkJr7TfM3fJQOmtW2fBm/81e3rLcikej+eTlaCx
KFNmFoOysp2rhQ09/R1eWVxv0H7trTj2WN4y/dB1PwN23BqbkrRj6xGC0eoN5MUY
GT0xq7A5DrPiSNwLUVVTb0F/IdVvjrY7xBcEmVzbP6WTKRAtu1bT/MBMol/8RHre
mQi5bsoTe2Y/wyJ+nkJI4TuXam5Ul2GFSEjfmDtBbL0y40Jkn7bqxF5mEwm9MNi4
nJR2lQ/MKAutA2/BMc+qFpEQMdsImwF3cbclMsCGUJtM8x5/hm50w7xRiO9wUfcS
WVc3+0oTYdGmrcVGN1Gypt16irTIPNFQOx3wkJV8+8g/kQlOIK8EiEoNLU9QGlBH
n+QIQ4A81WAYjw237YJGHeVUEKTFDAQbwm/iPG7guDEZZx1kJiFhJUkkeE9NE0lY
klzfg14UTwZ04jAZoj3OUcgwGplDhbim0+BBYK3iwnJwoEf0QFmk11eckCiPfaT6
KMtD08JU0BMuBkvaoT/ypdZqO255Tmv71r1SpJ0hxX49GpcopsW7b1WIJrhtR5+/
XQ7SfK8SXRFO4w0S2lDvWQ6vj0RKXgyE4Qm7XULZ5xU9xJfRw+DO1D1/kvUyMBjs
2jWt/B1YcbVLeeZvSXurZ9gM0bg5HQKAVjOcAcHaAWzpmoWaTnDJ9IvYltmEuNqB
NOujqKLawVDTQ9b5t0PRNwI6GAseZxIwfZZ9dA6+d1dy/371tAoMq7mRlAk+dzoV
ittXcgofbF5/ubcigEaeb0eV7vxlXoH/DOvskS5SB8y+dXYIcydoqYTSCKIk96vz
6ymP4/vZLM1zBZ08GTLbZvgTMTdcBMatCNsskEIJLyNXD4clvjfbUaKZuO2rDhkq
nG0V71FTPdN5NV59+rOmQjUQMfk2uUH730W2wNiYQ7lF+6YD2bnBjbX1gAtr709w
dDb06EYTRs+Cp4XJgtETgsMjKBf2BuQlRq0esZXWI99nGla65kMlxIP9TXFN4L1h
AAuPusbM7djtr+vVdvhua3P8DJOndR1C4kIEHDSWbUuVrjP4Eeve91U9bhFxMJsi
TUlB/PyU79zPRCY7QZhP2ZPb69gzxY7TtaqKeZBZH4Yt1kZOVVI78QBA38ikl1GF
dzafW0tgQwbSzj4ylz4DDtdg+8ywd9gWjmG/06uotDM/8+q35ikzatVLT2G25iWM
Sf43ECSJWeyfuFZUWCvKeBhcJePaeqPBltaaX19ASaiiFbfNwTIixUWD8H9A0Owt
5doARCCZm8k3qu6YzBMbHB5RuhqbAbG5qJpM3iugEI25KbH9DrcZNRYQSPRXy73Z
QshI0rk5id1hZhbWZr/G7cjoEGiPBRAKfM8LmMf706eYAX+EBt8vWLVEKRL9ehFl
ZRNoqKFh9dR0+oExd9O0H+0GFX/mq8f0I+ogY3ydOHi2X1bbISZurEYBaAJk/Do2
UeO5oaC55LGubBmJK8htayGNsbpH5pP3a1zxy6w1OU5abrMNbxXMGVka5ozLwMhc
3eLgs08flrMYkIk/d72W1pFOuR3zP0/bLKvIMwAHRLcLdEo/tNPGsat4Ct0i5jcB
jAVjM32G5HlIOJZ3uBX7tu4ODOXqaAz7VwB2vUIxm/6nIMQn6j6VCzw/jHRJCeYl
QCoMwAKDtOqTsF2TPRV95w==
`protect END_PROTECTED
