`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJPq4x69B4vx1z7ewmMlEJvxxmCoUwHGwbX/8FTdw8XyNqtJ/tV6N81He8BGnhfZ
tCotgGLe888WyPEdK4F2OUiIW/GsSGgdjhT++Pm0zGtvjQ8ETM7JB/Y1e5+Yhe0z
oxtJPUxtix/noUAk5+6IcizQMp3p1ka4YmVicWBZdX4mjtGHjvENxQHOYtCZYT5g
wfcRRZhyvbNm34HNaeLsYiwnM20sVheffF2xIMZH8fQ46MWLBhIOjsvm7k4gGV0i
En+DUEsXRkCkkPvbnMTC6snShpx1n0LGFO2gz7iTtR3HUf0yZ8eHzLKUCZyAshp3
kHTpyuQq/XQ7YYT7CvMxrm4GlX8bNsGz2XJfER83KQwr24BoYCS05l0UCX7Q0VJw
BIDyAOUL849eekqiy6gbBGH8YSPbAqDd77CS1UshjIIEI3wwvGrGZQb8O8bbXNGc
ywS/CofcJoh49gL4kC2sYImBML1/0Cxt+CM4WhijizeyrW4VsnvhbqOAJ3ezn7h6
QhhGx9dMwIi2RgoS75pSpJJpTrZ5H4oHfGehHiuf6LkL8vkPTvtbEMj0sNUc/B7o
nG6RIsnfHsNkwzutKsMt29Dr4ez7sD+LdvcIJ1inTsY9opGzc9i53zd/sTTbMsh2
SfB9sPVcpTOSwxvssXU6zg==
`protect END_PROTECTED
