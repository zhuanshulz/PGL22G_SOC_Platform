`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcy6gi87VNrXVTYzT/WbXzfzcFkMxfp0U6+r0EKO0VZzz6/WdLS7auHOLkCOqzFU
gN4QPyfHBVNc4JLMTR6EgDLc8yLUhBXNNvZ1av1ui9MbmX982RD/+W4wZC8b65wr
Rtryzee9GLYzxA11P4ZrxHaQ1HiX49khsAYrwqbwgl5g9EsTIbVwQeO6WoOoLTkg
i5OCFY1x/0Ucoi1DHpWNbiBPb6fqvBzsIe5qogiVkJNYbaL7XcfawnMae24LC6/u
VrtGHWVDT8vV5QPSUHyWEHI9n+ee+Ut++LD6apVIObYd5yYGEm5sxmerwb8+dS4S
g8zM58r/r+bP2ZGp7+VB1Ddk39CbOnWevFDvDOrQ3xhNWiBANKat0lKY91pp9LVE
xP1u47cKm8obIL2j528o64cUuLjDHnBzk3ZB3HFc30O6Qj7QGyOmpNQ861kP43dC
QDE1mrfvA5eeyDpNmt9zBYTTf00H4Gcds+WMTkcRvb+JJAYiyKEMVw78PfPQ3Vzk
0RzvYvnxguypfXB/dVZX0eA4TU2VWaL8uPx6fTQxjEc6Q846uBeoolsOGPlU9CFo
/XmXTgMSDqNVQ+IoHHuBlkmcWnLOPlKtO1TDTu2f9HV2te7EtaGNIlXF5oWrGuFL
4T6p3+s9gG9hnPtZIp53yW1kOuadHBmxe5tBmGz+51fFsBBlKj9FYnsZkaTUJ+tt
KEkAQBU9QvXxBIaJdhaEvpPhmiUtd/pRtzXIB5ML1iaiYeX0woj469iSftHmsox+
VAHJVUp2KzM2822IwZE0Mk8cK/8UvbYKO9USPMThAMd5SYtic28DKo0KQh80G6t+
GfWz1A0O6iYbGZhwp8rOXL9QzSHhJTAoR+2nA4dhJg/C1iDDGgfpmrThC/ff61J8
WmVEdA5Nw0/z/AGrWenkxoyKZqSnBRIgi5uCR3zllhpoA4GPVohzUdyZmk4mJoLm
k+b/xr4s54TTwxxRpO0mYpthZBbjPy9Pt+nOlWA4G9WCMvjNMcrY6Wyh4ogDqblf
rGs6qUiqruk/NBap2jZx1bs5HYgAeUx7it10nS4PeaRAW+PXpxnaOmw3vV4gkFYf
TfbAjzWeBz5I7rm/MT1ZFLQVCmOT3LaLRxyiXqXMpHvpRuSnOmL4+DMoO28WDugU
On5wW6wuiZKZ0LMbfUnD6x1pBW5JIppCp9jRfp92Kp+4YoEYAA+ffMaCRiYeR2co
HIqfIZo61+MxSDpS/8Td+nifH0/p8HBjey83muLb0aPnhk8gEviCNoaPKg7bPXCK
jeUCwzakBOcRJF2eMs2xThHFfveYFAc2QSg6dWuDOlDmU/cx2VRiHiFNcXKUyeXb
07tTD3LcswoLEeFxQyDumg==
`protect END_PROTECTED
