`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qTZKdylcSiL9FcwxJpRIdzQLpDnJWO1bn6pCPX4HVSGpGafXrdvrsSYI6iJvPo+A
xodj3uq6+7eBD0OZXbAweRa5Xy51DSSrFKCgz5N3gwbDZXiZKLT85CVdWHzZLLPg
wd0NCyyAx6a6RsQtFpqZb8gsZHEJWVTZq4Ar8FpD+5vvN1j/SE140++y8t2UfjsS
Y+6aHtjEZ/bphv7NVaicxBBQ1CouCpvr/6k5ydgCdjjlO0B9SUadfwKRnQ7OmzhK
y6WPnx5gB/7LPStrKnpb71o76iosv2ybUaLzYvNlbVJdXMTkBxSbmZGmf/rlkVoX
alKKHvNjKXjnk6fH/6WyCbgPRB52VuSYN6La0Wxqb/golW7jfo8h9koqW/Gs8soL
r6kAcr0h85/drFwMe6tAGpFoszIf1Rge7+UrnISIEomYn4EZI+gqFktJv25zTUc4
VkQZXb93mV7mCqAyda6QsGVwbS347LoW41lnj1kMjV9MiWTfk7ZY+SfhTP09TrVE
7jZyUvNYItqag5/WG3g+aW/gtETf+XDeZaaBb2oaXUgmlFKIDPw7x1/ekKZDWW+C
ucXvRjdirnd/or7scc2DokmZ1VFMvq5EBHXuAKTy39nkJFyQvryqJ2IArM5NzT/I
cgmAWzt1rKgyyUcxbT/ekeHJlxt1X0QknR+VxTQWTQPCc2kUpvK7KEHyOZRLY/8L
4E//TawW6QIv8eNKnoDvNAcMg+PHEfzQ2W3C3bYKPou7rmL3j661gtef1FoFYe38
p22RnV8IFoLjp0PybNhj7k3Nm6Nk4u/MVUJZxNXdkHoX7s2Ui1UkLXClJDYQm3BX
KZYi2gN6DoAyYQKXChUJ+hifibw949Gh6VKHhydNXQ0bCYp50lN27reh+BD7/0tu
hk/q0FHtLsMj4v4PD43fi0DeDq9+ecKM55WtscZ7lU+P2Ik/lKc3OrAxYDk0WMn1
ZLUoMQzSmkt1bKnRvsAJjO0GkBquAAUyI04hUp38S26BPUiCDdKdf++wvKZx5FiV
XOOCUR1kSduL6E0aTK+4q+O31qZUpl8Kh+OmSjjcQhuShQBuQVifeE6yuejBF5Z0
QuEs0owF+fEmZf+3TV1UO2da/Nv8OeHQIhZXHCF0UU9ZI0lkTywpJguPd9YJVGlA
`protect END_PROTECTED
