`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0BrLZ1oMH7/5BpLNUN9m24F0UBYGm0evIns7YIfTiIDG5AT2gCjsSinEb2Gklkix
oJXLbQtwY5oRFd9WiEHNN3SrBDouRZLuhOWrIjaEv5ZjzH3wZMjo5QXvPMC3CuqP
czTNEFtXtdG+mI4OS2mkSKietveYoX0mvHZ3EqnJve9xDvZYVnk3kM6XLw1EH2hs
HCbQ1h4ES4C8wAY9uEFyR3i4pW2yLx/ygT1m1+b97KTDhjmJaRwOGbw+d0kovRJ2
hZOMnllpethvaRnokSsO/4xE5HKuwKCKDlytbqQHfZC9QMO8jScKSPJGgOKzYjx6
kfMisMSIhcSGJnwBGDzXe+RHkxgAbWYiz2YS/uwx0BttHj8d4ORYJ5BTwtUVM8Fx
ClgaNC5fhb+uy/VrviocA9HW6cDZwVq6ZKP0pmCUlLhUSWBsCKE3cwyjQauaBzi+
zCbWyU+UGyVepGDuJH/jsJ8A0XZCvK4M9vFjpayK/5w5rqHA+vTy2nBv5aLCbYxc
CgQU67XibWvNGKTTOZFB8AvkAlVMEPADOlogvd91C4Fggko0wyn9g/ZZtKITeeKp
ssvHcCDtXJNT5on/B9F6M3usBtxOYtbJfrokRg2w4X288t+SLiC5KGmjsnK140dP
9XynT1GAvJE1ukmtAMFAi8JXthZvpM/EE7MPr7+FijOKn3H9YnKtpni6eXO1UWLe
5kqvl3LWxxs6HySQO4Q3sSsBmPQD7LPtqF49zEItxZ8Xj1GKnHkHHdBI7yZouQW0
isJW8e26MWrWXZhOzmLd87/CXKhWTUlMiD+bB2NvyGWLHUa7eO94xPiy5STjkRZA
XkSxs3Xxl+mysFflqMPo3UNXwT95u/Y4cIz2NhsWeR2ARVHHnLoZkhSr4L3jn69X
6SAb+LPSC7zf9i35Y/o/OJa/jRbQ3fkR3A6IsN0TgOg=
`protect END_PROTECTED
