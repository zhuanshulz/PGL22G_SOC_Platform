`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1lHTDvf8K+aUZg2QhY6WxYw+QAVzlnczNpGz5JUhBKDUuhIlNCY1mB1TdLuWGrH
weGQiZvkIivfB7bnf+Au+E/LL3YKai18e5XO6Dvp3VnftoWbGED9V9iaRONzKCN5
LevRwSDJefwJRJB//q8xL1Yljquk8OuQLXIgb8wi275T1HU4k34TjMEWm4n565rr
s0aWHl3BAEPkaWZn+cMph0vVsGvwi93LfYkswtovXpySt9qZpMaJPFLS4DA0TANo
URx90yszpARZmq1KBeqKrh5gPwtovsKPHXlfd2dqfrFyaWC3fpGQTmpd8TZjKS3N
J8nWMDNpeTrq9BaRHaH222CL2xTBRRHn7El2JRmn9zHhi1iNyAq1fYVtJXbH3NnF
lRppn2p2g0PJ6RY1cfSefOxRjbcVNNizQTyJ5eKfMDF1I4vzWebPVcyKVbmJASVf
ZkTKGf63t1ucws/MDqkBG+6WDRiL8B0g1d268X6Yzsepfa3JNFWilk0fZdybcXmr
rse+9WW97dz69283ClCwBynsMDeQUpb9JKVnJnVcI+Slh6na62FzSZFhgsrHlDVZ
p3GKBCAHCS2kZpQSRUsyql4APx18Rd8IQb16Qa4zUXgSO52uuHGV7KHIazL4xa6g
f7SBZv/kwFCHBdrJMiCz1l2j/Rmg90/SSLQHrNSqC7ACWoPDURDb1gwfcXrwIpKR
HAp7M6TqpEJ5xgv3SSBWoVtqHUhKMleDsH6GiI3bIseiLBay92Kg7GgMCEex9sj6
1KjBnqBlWoQgf9R4GP4MBfiQfTIj/0LhA1dTJL2jfrQd4nQzOkRexhSphs0dMw3c
r4dYrz+Dqs6rZo0/WZTdLJubNv/hrnihVGIJu3RuJr+IU8z4+GU135nysdrA0XHI
SmR3mmxzi70i84TmaXK3JZrQ8RMG85e0KZ+ghWhg+n9i9+wgu8zbCBHQxTzO8dPY
hooqsZBKHTq4p8Jj/TZ/ryzamvmmXKsL2oQz5wvq//2mSNTZMmagP3ILFV6uxIZH
zbK1zUajEYFQjsWsy4sF08R6nIBVUXJbBce28zwYDa/JYcPV4JDlnLn3FAaBKyXi
Ww5VmhYoROUC3gGlm4x91JQ9e+KXqqZ+dDA+gcCjjLzFXasRSfq+H6ejMzDSh0UG
/GRvlJa1QytQjxID9Roi08z4OuTJ2gqaPyjEGylvv57U7ipynnxpktEvYkhB30tU
NwvCVIC7ja7cQdXPGxRBW4qVN2W2Cbbn7JyO2RLeAtPcoIO8wJUOrVXcuJNe94ZT
RaQBsJLpMjir1t1cZAiw9awJlYcR0Lnwp1X1PA5I+UGmMvK4FWPWnx4WH1fTzH+x
r8uqM+5nwnKSvhM5NGwUBKAb0Sgce1EHAO+T9IPknHfXxUY0FgT6y1eM+gYUwo0J
CGdenywhan9/qlLUDdOWNFFgQPTBLUPws4aXRidqepQV258RPZjXlih1D4It5PnZ
L1/oTVYNuNCHN/dp0V8RktX4+72YAJUAGNcVjsZqJq8N1oW5WjA1S9I25vQIyT5n
v32DSYbIsBpU7ilNPRsE3iwBDqpwpuQKIV7nwE22Ophe2wJZEXxBoTqPWAafg09n
hbWH1btcIsOuoXbVaP6xG4+PNX4iZ2Ky/pcmRJvaIj1BcY3naC88lRmudN/SOBN9
DbABZNaqvvJg29tELTXZlqsHqg7K00oajB5+gG6uHeZTNuj97rVfXQXQBpF1AJFZ
wRrmbo1IYy70XtkFApYcLyez0+XqfKLbZsUxMgyjbPm5tR/hu14fuI8AU2rr616u
xGXPQWyahku27WPamVCZ52rziL7TeMJHZ0PVmTyON98L1AGBgwWKgLDEJw6mNxyO
7oMR/czHZp1N6al++phO3bjiLyQ9JJHaih8WSdQQf8f/VALdchcGKZHN00jIs2Kc
6cUR9kDKmGgqUphDvHFUEcVTpSm6I5q6fHxG2Y3mnQBLeZtJW8AsY4ZXHsHCLV74
H03J6IcRZau95P1tILhTWWNwcMDTUhu9bdmYscbS/k5zq5hax37DgAo5yebfB6Yx
vQVNCEnynUFZ0tz/pT1aj316Zl1z4MzTnFX8K1IL8ujzCIEC/iJgYehxiM0OcILh
VZDcURN8IbQEujOjzd85seojSC7t7G1DWWvVgEaxugqk9Yuuo9932PEY260sNzy7
YGS70Kbp35ugpZ0BeDyQNYAIL/gbtzkx0ez8azg4BhGjYaf0QD2LtoSp27r/QU86
DwS+owkENzuN/uxHuAk39E5Ooqthp2LzJX9lkHhTA8uJbbFzd09f2CMwzoYnlkXD
a522kOyqWIbWci6qOS1v4tYf0IZtBGeSK7QW9H9gskEIu+JL//b+F3JYsxTWbbOW
jC6n57fuiM0DyxNEgF85kSmgYXrxkiqhv6JwUCrmDlZRbgP/m+mRPYhE0rCXdHit
4Ihiqg++wTka0czHCOtyAZ4N3DKg6H6bGOzymTtfgDqGXQ+l4gvvBy2cl23a8+V6
TYwSwgDPJhJE1vB+H3xva/vXhSZeehRGmFQtn0zmfRj4Ubmx7vdQ2JrfWwKTJod+
5pNhQjn4ck9OtbKmV+3G7wMvY0cK/eFiMvSHNd/gf+qNhjwtqaKk58KufH0b/q9J
ew85b+l9EK3iRkeIMyJ44fp0Vo3dawHKn3t7K31CRTpTRoAkfu+Kv9xJwYr/0dPu
0sPe8LQfqhnZnij4IXHM36eo9w1njQ4ZfBaChHFHpvcyHREmI9jEVME+F3b1DAlC
/WEbZ+6mRRUXvg3o5gihgk2p6gTnwxfgx43YFDUBav5dirq2s0I9LktjCoQFx1Ru
i/KtOXQy53rN/O5KgHMiooJqV0IbVX7eFZunqQ47t2gTeJ+kdpeGA5v83+Ru36y1
fXzvaqDTf2MuEH2s7MvI3ZHHICZNeUjd4hqnrKEOIxdyxEgS0/AjfZzcDF3//gif
QBBfoK66j54u4IQQ7APPSx5d5ao476swBP+KVWmz0/n8yNjC60blqTyzo8z7T4Iq
4key5i1XACHnbmJE+HF1WblMDJTrwh2LbFMmc9PELt0PB73ks3sNvVhqUxbgUoj3
orSxic+22nMzRo8Cjq2aCnTKAWjmcrO4xX935ZJGdQGSL9NFmHay+BdwEzMUvFMM
tU4BiIuQJoaUrNwHxuGosKejGjYVW0tezPMdo9v8FAAUSv6TAFWeGvE6mWUA1jH/
gm9tCTDYnWPNSSfPoh3Y0mLKPLykKpymjFGAAroJOWwTSRgQ+MEycRtCPPrBawaM
IFJjHk4SgWLSYaNEOQW390PQpPLHcRMenv/+yVo+0XDEFQudCngWUFJsvKBVoQHb
6iZ+RyqhvvBJSbEt4UknWM7uXta5dxWyw+xrBE+QeaU=
`protect END_PROTECTED
