`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h967qBRCZwzPI4eUo85O5zxug+gOVyiPBPlPCkedBfGez0eIQ8hGvbq7cEACztQH
jgP4fDgVhOLNu2iURxz/8iVjJMWoZvFOIpipEb47RimpL6sYIpGLBQEP7M2iEvd4
pC4JW4ooI3L7YLk8ClJ+mU7owQ2u76rx4P1yXa75uLn0/e4uAGawfhZYnKJ6twnE
d65MHo2ImifkQMhSq9nDdCK5rcjRp037OZApUNVH6ea7LmFA1V3Eq5atTAv5WYgY
EXhv9eBvJrdPQIXCI5iNEr7GQpPWFSOyfDLSc+u+8ABIKM1eUEkMqyA+eG/kDg0E
uXVx+DszuRhpvuGn5qjGesVxBPekOES+fF9A5Z2aMSyblp0lFZP1HOtE5lHlrBqp
zu/wDUYhFtnKC8J7i/XTqz0E5H1NQspEzgFY2TTvO0I=
`protect END_PROTECTED
