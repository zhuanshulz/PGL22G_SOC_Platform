`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CCP0zqHnaoM9qmk/lgIgon+hd/0oC7TB56VUp/avyF0sKxOvVwmZkAb3AB1f4eX
rXhU5I1VlLndhOiq1wjfcpJCedjVxIUxx6NzF0gm7ELc09Dp/dKXldBXI9K1h2bm
0VKe01E9X3HAQpse4tbyxHhNZXfVXMytJTzUqUFtAfiYnNaHB/g0wHAmVi9J8FDW
9A0i+L2RcWWIrXXPvmioc2vcxr4RWFjBtaj4EOn972TkSNISCDEFfEid65WHSami
Nhf/4qOxfMPvl6AAr6KbDVMXkYZyHwJYzgTGtrmdyrhImGHWxyzGmE/Ga0Cd/LR2
+Y7spv2h9DSkR1vVhWwhF2p30bNEJ8WJXostY6lf04JH6UZoIBvhRtzWx4X3ZkO/
itrRv7V6JQUi9QLA6XcrZR99XT9wh6leUU+Psnyn9/pIemfe+T3SQ1EJRmu4zjfz
R/42C2rFzbiE/ipMl3XmBzYZXxm23HtqQPUbsLnL0THFaEI4kgsH/RgUoTjRBrIK
Mc+p4NsNtj60LboAeHYX9g==
`protect END_PROTECTED
