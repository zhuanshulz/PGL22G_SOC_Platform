`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/kATf4Jkz4Zm1mQDWYl+j9GBA3wJIkhntFsbXzyjQ7mj0YqK5mqbphz+BE0JITw
kyBwsTuMzutsM5o3Xm3zdl2qDmWkFwtmGlWO8nlhhBSQALs51FF0uotM5sPiku63
HgUP4XWER/Lziajr9fdAStGvGm7VQcAPctWzabX20XKnpX1RYgUM/hCgz3Y5Gwb0
SdWnWfgqsM+D7X9Wr5Hp0cQ5xCCAXslW+qlXuO2+00Xl5JKI6zvvOf618dUHjXoG
usVnfEx08quA3BoZvioD2TnN2zKxXWiKJX51OkkJk6ZEjYllhCQoIi6b++54zB0Y
xjOXft+M6w1r2EvPaGk9NePwv8l+ai02z+jIbu5odApdJZU8xNnu0qWsRYdg5AYU
JJm/6kmz7UGCjwcva3gs26lBLXRBJyGu/UK33rwnaMfmk2C4YlDpk8FrawfkuTJc
HTQOdsGArYFJPd4JjnCA8bsVeJLwWhwpmYKEy2tkW0s2NHXxRq1nPxrE2F0Zyuj9
lX3NPfmIOlgIdks3za83slrvw/yK/6JyhxfsNnbU2t4ErTl7kqzhNz2sRBnf1cM9
qSw0ZWB6wHDdE/kVocGAfg==
`protect END_PROTECTED
