`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pFJTQpX9taPxbyZK0UKPzKKOL2plxWZqi2NKjn7ee3tkZ/ZMY1TYilemqLXxSH9x
C71pnkc1L1vbUQP/MMW6TQPv9AG/1NQSV3raQpcVnai0eVlnXmk/HKbQI7J6VieG
BpkX09YyHsfxbpmDN/a9nh/sHmI0r5Mcs87T91efPYBTY0S4B1O4XWVvpFQ2iWBJ
yfBfxmKNFQ4RKJr8dzeUy+2z5xRGowcmofnSZheS37LiB+j8b/9DQdcHF6+lXF8C
u2g9acnk98kjQQEcOZzRupUePgId0B8xjSUBzHicSTGlRNuylVK9j91WcHZ3oVec
wcJBJtep284ivZvQIpIvizRA+qCYV2fx4X3QHkNpFuHY9VjMH3u+0U6CnySyQd3t
dQkIfO5K8DEhTra05PNMHBUoUhdPBYeV7C9zhAlWzFfOyzfzeMfC8FjsazcwT1vs
T0M18hqdD/eURj1ncaLywkIGty6X20thHYUMAttZ6Lc+RDJh2wBiqQD/H6VCO64V
xGqOSVewk1/ZunHjMXcya53WKjQ52zHZQFy+jwAfWht4sTKRChyJavUfPjYOVZGJ
+DafYnHRuRLvRJ4rDPjsBLwhxSQ3nYDMBijJILoBqitfg5HTRL3TKVoXEsM2BTRe
pN2R0RJM4lsexgVIONAzaw==
`protect END_PROTECTED
