`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XX+50a9bwSkpjuu06y0GkTf26jFCVWmu04NtWQgI8tm46Fr9say4suTiZ5ZS3lQ/
bfetMJfzEiQqEEKXWPTmdU7ODMe90gYbzAb6mt4WP8+HvO+NxD77hq/cf8oJOlHT
Gamn2wx+9dpImkt20CiY3PxuL5DXnkOv6Ml0rb8qecicON3V9lRYIuPuEI2gqika
F6owjW9OpiGBhagJ0s4npIlmyeMldarWQn3AnZD7EaXlDQ2iS8x7oXRjN57EgOnI
slclE7glfFkZjxBgJbLhGseLskW/Pmvx0RCdJX8GjvEDy4qi/WJw22MaJ+OOCsE1
4uRIQM4f3eq0rJlXOpzoC6MMqUPC3O0chN/ndrIjuy5tg7xOTm7YuTopJOQ8VfgG
8/cQctn8ESnNA5UbGZPU7A0nCOY7tvq57KR3rgKep/p0dBYWqbae9b+j4IiitaPv
MZpPMKOOHFEGywH8KQuGKjjPzwQQQ3m3Sb3Ih2rAJe1EUWstYqdhn/803NHeeRb9
+8Jz2hgupw8u4L+uAF7RiMJMDGZGjKgGQBXCkgs9/bvP9Hvb0Jo6DlzDMqh54A3G
1n+pY4gWL1Gs/a2zFd4w4Q9b/2B/48LARAWNRyvNPJimvhp9NUDFL+xttitK74xt
xS2YUz62C713vNrR3DoI1+NKOTsDC/lDOpGLNfzvWkLwXnA7tVbzo7fdI6azJrUa
xuEudNFZUS4EYZvsqqZZrKHirmIkYglquirkFvS2uKyduvfb+ERy3s3cWpH2xVye
x8Kp6UZur2P6or6lp2EchVe9nvf3ZhBNZA0jFDJDzR5tODHbXsNW8HLth+q9fZ/p
n8ZiRVXtCUfUD+aJ8GTSOkb/XkFlPYqCiCcFy4ZfQYXoKfPMxLYlqvSYCkpWHX3n
AiXREi1JC8OWiNMSrVL0Go5HlF8WH3Qan4qfTCwBeo3GmUinJCvFKRs7Zj8rjhJQ
Yspl1M6ijr4oDUPH5pujCVpRigYnEtOoDd1NWPGwtfjXMk9WwP78a3+MRVwn5Yrf
udcXXaKry+wOeYJaNteWxUjQjji8HNk0ZloGtwplwLafjHmC8Gt7fIFVc5W/sPe6
x6Vqmdzq+epJlBXbnI9YvEUnWrl1gkwt6G2nbkVDKlaZ53JgaiTdhhxHapGC7DXa
N/jf/w19mdNe0BlpjGudBLCfq5kCXllvIN594OHCGwKWAfWqd9avFWh7pBKle6SG
tDBI1b+HCOaDnu7tYNHvDnwY+99eybeuUEmZzA8lo+LOmD5/RHXZhFNF+PrjOtKE
qO510cyMZNmqRQOpw74FgaRNu/u5haKKALsw8IhPzcuUZk4vvUjATjyRnxJA0ln+
u+sK6sN370q3htC4O75RfIeGZF85z/YgX0+JeXa/DRjbwpJ/AiH926zuylQhEc5f
lDWYmh5laCE6xwHwhEKaUzOS9whbTMt9WrRYMxYaOdzIGrIQ0TcqAkuGcjZZC1GR
1waVQkYbo9WNmpS9+PgWDxEPzkRY4GXN83+HtAnTUQdmzPHxdGPXGfxtxSI0m6CU
QzKjZY8OL/I9kIvgEdCEnmEVFhXkrD2RxTnTbeFE5DF3MAiiMuxVVM7okKfox2Ah
/J/0u1JkvvzO408kT0mw5oQx9CwDcJ2malr+PHzhrCZQ1OrpzNOJD+LD6OE9JEVH
lTufCCODq7u1fzf0MWteMtQt124TkFFJSsXESkvDg5kxirSm2tk+bvXiSyqzJ3Kc
FjbU8AUjeLGX1Tt2HRTrYdG7/rUBM2sdZ2E3ZsNcewzDmVA+X99bdo3WnGP2rdNr
qH2iyb1hhKJchtdVU6PRych7LDpm8aEIuSOh0LUydgSOY01Wk5OFrFJyH/1gDSlk
`protect END_PROTECTED
