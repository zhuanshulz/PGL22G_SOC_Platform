`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T1/XyvoPR/mQg+Z+XcXBybqWMpRiYYmaxXxZBL2Z1GWkeNOmKAmxzdxBv7pLDYJD
z61uQNglpss+tTRYGLQ6IS+W+s7krDPzaF43qQ67t7hYb/2qJnpaohSBnpiPy9fx
V/GSd9JtkQZqu0qb8E6qIaUSXZKF6c9PSFmF9IV3Ze7Y+i9zs4tFa2U2MEJ+Mv3t
ePWOAy8tlAPgTS9Yt5u9j2aAsXG5miRPDRaLVdiQul/haE3QbPy8EJOJpL4IbCrB
Cm9qzIhiXkjtn49uo9yWpXWYf7tIrX6Qryhy4SiIUglIRuRiYTwHNNAChXd+m3Y0
uJNxQ1ze2Yx0T4qBjyMKj6c3UzOi8GBln28kqBDUf7Ui9CExityD5GIChdUNEHCG
i7dWXZ3Fac25vYfTnnZUPi3sV7+Or78q32PQSJkOY3iXWtIAkutyyAvOntL+V7kX
/ArNU2ORgz+srrJkU+5oIvx8llEqI9zQXPXpt1gtfoHBj37dTC3lMqGGJS+A3qca
KgTMVgchRb41DCWyJzFziFIDcPrT3hSlEZv/BXLc8vBa7JpeeNFWbSKSp9cQZU5Q
zbCuzb1FW8vFpqtSSGDRvuyCig2C483jVUYOIfmoJ3sLW5gHErb1eB7NqAFLEG/N
fOocouL+yTdGUWneZRbCb/3Yls+RcBUwY9b+u03hb8dZ2mz6xG5EVi/q4TNDas2s
Mdj9G0H5K3hqZO/TNR3vp8X9oAoWmiomUS/inHZyjPozEr84AWBeifVM0J/PHUBJ
EQqrK7sN38tPojVPrm39Rg==
`protect END_PROTECTED
