`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Nvbmp34mwZqwytMEC6pRYKeb+GEq0xsTv0joCwtVGpVVRN5GyCvUZ1lUH4/odsR
K2UnS+FkXsOgW/CWT3k3UvBAkNvy2D76JGboOg7rS/G3t3ZgARJ9c+SJJd7n34kN
/aBl+mZJLUDMFKpLO9b9nQXpUj/24oBpNcSURmGZFpESTa/Uc+8/HIjx+Bz6ZmfD
KcUCzbEnFTa03V+yGLBRaChIbhm9qBbCQr4Z/7HFBoxKzjh/FPws4xe1mMaRTU0p
nJbzJ/dbhpK4r3ilKzC5JrVLgexvSKX8k/nGEgeg5uX4RcoE9dzZEbBwTra+F249
cQ4jGurJdXTU/gljNXpVb5AEBS+rudnqc+R845rYU41zC1u8OkHYltYpdqv9e3YO
ZLR5SosDb+mOeZPx40UBAr21DSF5UGnXURLaCHCwdr8Tv7s4dMs8Phxlg72QV7qH
jU8BL+MEB6rMrWMm4MLSy+RClL6WGWTTFPseTrSgOZPM4nZHOBzIAPrMOZ7mzdWj
ZLLFr1kkijyYEDq5sWysDprz9ECtblfrBV+PKBbTj/RZjvdzFxDbMaJqrwdV894T
kzTKF6ajO+TXK1rXxL6CrQ==
`protect END_PROTECTED
