`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvfV+QjIvc1c4iZLytrmuPfgsYUh1MIWfSjJ594cYRuDItE/V6jU2VAxFnmwnjJx
l3o2232xKHQn7Fu+xLRQK/aKn4NtHlRq5HkZS2VGYboD/bP9qllxXNsIRA4m4ybP
BwDNDUwy62jzACLdsLhV5spPFoEWt0rhkbEAggSq686q9j2V5pOQkPTunAIir2db
1brQPV+9kR3nPdtFd7Ukph8KnGPzw4AnDO5jqmLY7blh20vh5vya/zon09o5I0/E
V/f3XaSCRNkbrXU+3SlxZr8kEU4nBd6oJvmD9+qEqJjUaROrAJQfuhunJq24DGSG
utbgewDmqIsBHRb8UfoWaJIV/DpFmZDUZZq2SRIpeYXLdtjGs4JGfPYdLsy8bea/
epZlgqWsVCnJofT5bAXS/SnV4oGkVs7v191OA3D/Fg6Jt80dbKulQDZfxpQu5aeO
CqOM102oeYJOcXvoaQZ1TSAMjrwPf8qXSfLG8/4/IyDXN/M6pswleUSf0mQk9thx
eJJI9SeAB4Ddvbrewg0xVWiR3/pVK+f/g8jrDsPQaTiutvUZzf4zmIfa2wzGCcdU
IrnqyS/Kv9KoHGJi0TeuvYKd2TTIdNFL9tgADmTvOuJgAjltPlynF1cj9IjHm20X
3gHmHOtOkd4D+C+FPKk67g==
`protect END_PROTECTED
