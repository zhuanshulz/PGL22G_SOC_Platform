`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmHM3UvaRYOG9vTsgFU43w+ev5GSj2JWvqx9AOGRHnuUoJihxcZBmXhrGiUXkOd1
+vxqo3Re4UzLxeIjFTEfziC+biPpUQFWAtVK6MzgsTVVbhut+Pgz6zNcSRRx6Yo1
HPDMB7UvDe9LYXlHzc05GYwIZw9BbQuPp5ePmAdMFWuwgyvMtWLMd6oei34XmTTH
kIaf5nKW/j7KouwPxoSzpEPiRp69slnq/6AZ5LsESlsNlGUNudQnYkeizWcKMdtW
FXu3L76RcV0el4FB1jdRsA8dFs2R11k9AYiNVHrxH6dpI+agUpkb6L2IJMT2XXGH
jkyym/AiIPn9f1Ax1DTlJ5RdSLDOGOefwt9aMFGlG21bIg8gxCHia+r0hWAvkQnP
U7P44Tpn88an32kKHtk8DEdOHMDh9v58Njl6u5MhuMmhKJy2dtDEIhzO6QwsEbQk
o5GIP83tA5Qg11EKZ16UfcttoZxbTT1yWtBnioswGDe/xZJOeWLzpbEfv6tuj6ky
zea1fBo4d8NOfyhGDI59so0WsW4oJ2SeRkpFVz3/2spEWyZ0QH8NR5Tnra40yaab
n+BE5hjsTtLPnTafH83ecmJKZdudjleIKMr25LmsPVhI+36uVGMDQcdfIGKKqZoe
5wVyM/IQLYjo6P3CkDUXdiVEjBFaANSde8K7EXgtlPi6VyzUXB4WSjCZYDN6h8v1
BQ4fHDzsvZP9OTX9h8cXgtqIEwFeH2vsmecIZg+DDTBC5vOOa1rij5qjmvacQs8t
do/gXrslsDyqIkhwJVRubVmx34eSmRiHIAWJXlHRHVXTt12VKxNSwn81++FV9jBH
CFQdSnbV8dXhKAWYtghJrAkX3R/iWLEe85aTdhk79BX0oDCnXN3KPzZ1Cnp/vUMu
z/ZPbFs+eUGXWpoO9IGUsg==
`protect END_PROTECTED
