`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zekTpDc0Oi4ZApkahqQWpF5p70HSFn3ZJeQa1u4Oy3U6fWhLtvjbK5WjyjtFTd3I
mV4xSHTbGxTHelZ0km9KxNf39RKx4EAt7jAS5it0zY+9XG5Khw0rYO5w3MCNAN6E
+grJlfjveGCa/f70pOGgd1+8tkuSa6a6EDboAkW/aOnARDGsUX0AH9nee1VE9rPU
4XVIzV5XXFeZYgL3wNRUN3yt+tcwCfusVOH50dD4LqmWBIsmsvYzf6XM4Ov/IJO6
3I9VKXpLX65HvgFUifWh2v8drPTUtpe1Xy43hRQlTnsOCUb4c80WO2ufdMQyte7l
Arbq+ACfsSyGgXnJpf/cIC8poUHcaiouGBy1pulSQepW/t8Uxy/g06WQldKxBniB
G5/p2eFrRqusFaQvlRXRBW8bWqAgqjQE6SM+Eanubu4QWC71z2NekN0LKWVCmwe6
o3Och0dZYmJQlNcPrnrM5wPTZ4wzp2139+Ib+WCLmighd3owhB5ZrMozYIJRS7qa
w2XvbUJhRuHqaPLuZolikO0XkM9+bUF7oap85vtaTKWZUJ2m0T1Is4O5Bu5DJ4BA
4cezIRdlxMEdH6Yxi6c8RNrT13aUOrpJcN5O1a+17SePKmN3+9v+6Lv2uc1YZbdu
yxVtjGlAkgZC5e2n3z4FkZdMIki5oDrH65gfuWdrunU7w37zQek8vpsavfZ1XDGB
fY1PBHRcsjX/nMGaVTYdhChX8e3PDgz8hSVY6m9Krt/B/QxXm8xqk59AGU+KOZwi
FAdbG8ErPCMt0jkBLgwFHr72KTuD65jwPd884sSvtBV2/IOg234snrKK/sUcK3H+
CFRfgnfUz11P7comODdMXKfes/I8cahJaw3R9i9KtvEDj9uSCejmtjQ60cVzPDT+
E799ZGEYHqucDLkgpOvx80HIk25/Hpi3U8o8O17rzbdTrzL684Exb2EnwgTGGPwj
gx4RQ2u1ge8EcZcfzw3XEss99eY1ft0kQHAV66CvRKQ=
`protect END_PROTECTED
