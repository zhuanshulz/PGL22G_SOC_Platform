`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
npRY/GT5+croFaDzVeipwoD6S3hrVRvdqIbdHA4do2gEJYAwQgRtwrM+HdxW59wP
8Aq+kSh7QJc6hX/oQV3qNITIpkCrwUMC/eLKrMyLeQkOGfJARTo6Kxou8qiCEcLS
4IPRvmOxr2lClkesIg+EnywQ0JXmXm+cKTyZjY0tQ8gBJwhy/u1TY9gi+BaCVubi
BO1CTUVOBoHkWT1gzQD4BNMYGFwp0GyF/mSjIJgXRU7C5KqRSASbILs4Mr+opFGK
l/6e8/HDKVOtkNv/cKY+jaTCM7a/PCMxUpSIm/EiO76ajM2jR98KM1LTSx7zMOn/
yMRKhT73I+6VYUmh1OskRv0cbEnTnW/K8pqhvlLgbpaPZ1p9wHeQSDZ0Z67vfL8H
2+c5jmSfL+0q0p9MVIzqDg==
`protect END_PROTECTED
