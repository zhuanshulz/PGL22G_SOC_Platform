`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5uz6JTcL0MIz+ZyvY6IeVqIJ1Fr12m+w3febjtGiRlFAhrBNOrCnEFuyLkF7YFt
FUAnbOuKx23S5YO5aaFdX6fSBve+IrAqNbwAP8kkalwl26QG2Ug5crMLvF6HgVpT
1IS9gYFi87PPPO4dvt8EhLb2KXaGm5kTC1oOgyTFUnfaEAa/ve0z7hddXcJWB50T
DZatFcIwDAY8N6EawMkm7O0MdTmc9h5YNPXLfetxKi8N27sH9Vl9MeAdg+Jtk+Or
KXqofWnk6cBtsNQgIeFsag7/vt0iagX3mQZyrHNjEGGiE1N8cc6QxZrvkp8taMcR
441o9jAp/Vk1kv8XJ0k5tjFnxRkXnqQ39x9yGkoFZY2Ci3vVrMjbZtV2BCLhYTb+
jAhv5ULT/tBo1tv6SSKtuhYh4WzYfe2b9NGNKNqj00pvlhvme6HJJ3B5QZ/dueBs
mXgRRffoidQXh1Dcxbr8irwW2Jw+HuOhYRg3Pl5y4h8fiP5WmXmYpTrLD0lxW6mr
hhzIF406f2/TbANWJsMyLXEtXy5Mj6naz0DV83Ws+bHG/dDDXMb5Jfbqd8kkczwp
I9U+Hd7mpuEthArqLJCZ69zVONXgimmiBEkWC3W+ItTMY1Ep7EIQtfbgM4Iq7GLF
CXOcR+ktXq1vIHkzvSQA3giE66pCdgp6I3YGDE/pwDxOo28dtdgbbB8MhMjRHiaR
m3U6Ed814FDLuNjLUK+O/sddIE2ddo0gcYdd7P4yVX1ENsT4LCOA4oIZ/x7oXGSj
CJR2r3FIx6rGfYt5oi9Mbcdg1h88mcyHpeqBpbbGqFrM1/Zt6YwB+6w58Bc/ZSbM
PSP+2AXe9A+u4jPm81cYJbpRYRdMrgh69RhWvDsr8glaXOOWoZSnUw9qxmd022Vc
/ub1n8lOiJyuFe+8KSEAP089CY9qIncgBVk3e3US3DFEj6vh9an5/OiFKRqBRnY7
TMi54gE23KMSsgjWLXJPLYWWzv5Ucwg82SBPlo0QLTTBQ+xcxMhZyvhJa5dC/lfG
3ts9LYZaaYZ7R3SUsWSugVheFAtBCcTOi57t/e86kIzq41tjDNbB9Dqmw0RVYxRx
fs28GxSC1/bgI60ouuElBw28rm7LHOBY2M5KmCAxz+uO9bMuIWfSKFL7q3Tgu2PM
3ogRU3X3C1LwnxuyQSbeJ+zemQ+XZC+A+IVrXL1bbRH6DiuCYpyPc8VKzt+zbL47
ciuiT5qtXtJkco1EKkfk3TAH+KQi+y23aAmEjcw2xLG7pibqRe/7JH4rxpZVazWL
2F6fFaV/seiXqJqWyURXJq9aHgIk7FJ+KeMDHTYTnbY422/uynzVFk9E0goxN/+4
vaqtgM397AKpDT0p5HOcubfhhdqge3oZL5OIG6FMlwraVLEysLgV/VvZLwe/5Cq6
oEG9mhJBdBoGJvgUCxM7sQPtT+UiRfNatZFtYmBETPr2ELP0kWCSU/4EJ6q+SNnH
uz6Rq0pe4DJPoiZvL5a9/69s+BNZlgkWrHPMeTW0HSg2hZcfIRmTT+OoEkNVAzdL
Tji8kUa2GwyvoBRad7gXtcXZQ8Eo7dhyLpbtKfY5rwaCPQ0R7ZEzO6Msk08yrmkW
NKgT5FSzzoiZ6cjrOrSsqbNlXnAvQmVkG60fJghbvH/mHa352a7iJj92db6/DNJF
atL/AO9FN1EVH+UkMeAsgoftlbovWphoghJrpIcbAEg9y7drcd1OntXJNC2M7KYT
zGRhxeyHdP1UVaLRrMne30XT4uv08MsfmfJMdUic0wSPZ+bSvvMvhnXKZlg7hcAZ
pK/qXnTpNquIjgbJ5ryygONbU8bhUUNEWqD5z5jRQCHab6491+8obeBCQwAvOMID
ReR7rekplFPee/JKw1Hnj6a2StjLLQ+9ohBCbYGdQJG/AEOMZHBpUavPP1aJs3Hr
WjZ0m/2VFVxjnpiUPl95QZ++Qy+tjo62ZtMVLhNf4OPDDK52Ircsvdb7eDAdVvuJ
mkdItae4hs0Z50GhEPyTcnxwy6w3M56MpcdO2sO6FrNNp9JqLk6t6GYq36Y0obRk
bqWK6TOLneCI6LNXuwUSGy+1QCcUpIAwuZ9pGqiFuh3dhQDSI1z6S8+ulIoYI1V/
EcyiYlC+3paKepENU9d1d5rmGX97hHx0xIwJ33buuDgTccVlQatH89RenB5Z6OBv
202/mupmSWPi/Kw34Vodn3XnQlm5M11Z73tjSeW35b+1ogzNJsQQNc8zcusnOrQv
r1+zkLxEiHmBBkOeTkS9ANBGA33dEGOUSBO/6s0N3A3jRDUz1OsJ9Wun1achEkPs
7qMpcOsaXvqiIhMPF2Eg+4RCI5UmjrWPSCN3I/lrWVOQgaVAPEkGDtKTo767j8S8
YLBoeJG3xTIb5a5GVYp/uSNLYHkRjpT5L3JWaKG7CCPnDb6D5w94gh4zO1Y1XPK/
B+VnkUkHyp2PLlYbmu2InTbQRbERTUdE5Fo4SrQmWkTAdqki4JrytPXwZV2G2QQ1
c5wRoMoToUTptHwe+ZcObJcX8ax0TGSk2GmrsunTUc3ZQp1Ew5qij/fnqnxRk4oH
DG+nKM/vYnJngx4kPRae+sSWt4Kj9pr06L6dT77B/hCdMP6OEnAZlc3DclYbqBSe
Ll61T+l6Rb9fM94k/lPWcHGwMHFRATVvHVUtJTsKrWlsCNv1bv9MPeqgbzKT5mix
budUrwExc3HsE0bLXjhG4uBYhIDmwloY/42VO4rFxZeWNFH8bkbGvliIPBEN7nay
ptXNry3J9dRLiduub/P1AiF9Pr0Ncf9eRN8av5r+H1XbIwUhWsLxJEud3wH6rDmn
cp8gDYXRHlTuVoaEnqGvyOCcpsgNClnY+rrp0mJBzSFiP13skuErXex0bMqWyo3M
VeciA2PJeRUDOD5Lyyx0gEdLIMhcKhJG5AO9bo2uC1gnyKesNj1K6K3T5te2oIQS
sgkubh70OAeBRJoOeJDaGgjv8JOsKoyerjWe7smi2yvUOP0tDDRwXcM//9h1eJRq
KFXipdtVzpnFnWovRsMjq5WJIukIfIjYum6qvsByfjXZPPK9nCsJqbFP2zFBjWSe
3Tp1Ur0wjDhaUJi6rHRV2PUwc9lT4cAacIDxy8ehtBmANOdHx6nLqCYUVMAkzvCX
dte59JG+prwzNGZwzUJ8T0Psc86U5Crjz4Q6A++v6dYt2+yafv1HkBo+TA+xcRSB
WJeoAbcHxUZvbQ04D9lCq3145W9SZaEyJN2uxHID6WPeiAETj1lPjKgRt7sx0ML8
lolLqXfmqmPHahpmuOC1JVrtqiAM/G+0iWlxbohuot1aqp7loh9LKhS3NO2F7D90
sIcZg4Qf/wli/iwxwv6R8pxeM3DhY7jc3LrEtR+tVrITlvwJbqjY/NGMvsWcRBhf
0K6mYgBEbx7DOxXZb5Na5wkddOhTop5y/PSeE0keWcVkfF0n6CoQb8e5AgsNMVEq
TZF17hyKfzAaTmf5s7GJkQ17DWzLZuDad0uTINfrP/56OMGy1D+sAQqu58GXyBYD
6zLuyUexsx33XROnpGpJ+Cml1fJDzAXmn0A8ySPhbYy/SfgpLIKukRQj2Yj6/8Nd
+DT4j5xO3PquWqMCm47Z26H6T7LTCgOL+Dy7GDAdwepMeCxWzLMj3XlGP33r2x5H
JGZvknri9uusx9cNJ9bFUGtX/B8c1vlDj1eSyWRaOs3fw4MBxx98XsN7rpo+m/P7
eSi/OMkOezyLZm4DB3ooHJ8UAXdCEb87+hOY+cwXNIYC6rJvnsa8Igaf526r1mx7
/fVJDkXgI5x1Ly8SytIKRrAw5ILkf72XL0ETpgNoy2j+qe8JdB/e69NaLdjBpYJr
uxNCfv40UzG9VgslBNUgbz5KoGyb7tndqAM6xNzrviqmdj/flg3vDS+KntyrbL8Y
HAs3pwq8phiDEVW3n87vqIF6sTUt2H/eQbXxTfi7U2FCuXT/qyKGRFwpz8PZqtFS
INhbUsCvx6Tfu35zAaM34jfUqEFu5PP68v7gZQPyytuP1xp1h47UEqIDksK5mr8/
8TLaoy1NGVXKNumUXBcMtGeGoxKzN3Uj9cil4R//odeYA+0FiSdYfP4xvBCVQJ+F
5a40SVGnnf7E6SF533Mo0wLHijGmVHlIp3NtOwNEotvRRUUsnAXb53jwLihVuGN+
Z8Ej5AfQIKwI51dgCyQB5KHGZPggSM/hbxfAB3sA8Y1msyHtokoutwXmSqcePVIi
okuR780mPfLq0fWwhfmdLXM9rbq7BW2nfGc+fDOx+GmjV717EeRtOOk/WsdZUG6L
Hql5NS6Xrn61RqMx0wM3WV5InUYVQlCTsJioDlLu34HewqgraG2XxS2rMeXwTEqA
zshqmVKnLaLUDPwTV++ZSaqYE3AMkAPdlZawldzrqpXkpNzt34R+HsCVSrCvctjx
14hT27X5ZhlH/XNCC+icD7cC3/lBiw4dkkWeaT5OLm12Gjq7KkuFzldLdqKARQu/
mTjvGacuSgszK/PcolcqrcB45PRTJdGgPYqTsIPBnpqEbEfyqsQ5Jol38Yhq9cne
sUnJWCm77WtZEjAwqVYTHWwyrcjJuzkxHOuW8lRqm8XLe2anFSdRZztUJKsGuJGB
3HaTuY/mZbQJvG/xF3DR7XRAYgNmIQVk+S1E3irxtFurSOZVo7gS9FrPSYoSCRym
XoZ64iNZPMhdsEbxvFv/d1fz1Y2kCSfFddCABpuD4g5SXWp7bDmHwoPgUy51YJb6
soEshj3cEv2nx2axOKp4O8mvgjrP9jGokQvHyEueP01KdAW8b8LrmgzWo4kZe+L6
AiJwDMqYwB0DwE9cKjx7vTsLmPU1YRW474hOnjyYxIVizYaBjP/YgN8VjvNSHqx5
nkQMejMR6fLQdY7LHzbuP1VMFeBLMuEzvx+0pPTP591nQNko08kOP046UwWtVitQ
4ES7uPsnLtXHyJ6XhQqK2peFweuWq800wG9X/8/q4mhmZ/esags6RAssjWTHPRZo
QxiKP1gvZLE/nSTt9lBXRYP2XKZ+BbYbsubpead1z5gSnq63U01cXsobm1uz+dKZ
9xBRFdTQnAUvMbHztKkm/rGe23UGBIGt5Qx3VnkkGjYBLrK5MTbspsUJZ8SPLxCC
KMQiZ3cl7W4PR2NTCUCZYF+rToAzpfTU10Wcysyg5s2z2JhT6g4AXWoBlBY5vl7G
tUmqrXxbYLXP+RxY+cbK1OkRMs6uGMW3qZgjcxg5pEpLR1tnZX0mAtT78MrKxIJs
CiXDhh9SqWQQzq+V+JiBiTiUScevLYQ0WKyWpeWeI/rYcjfvNNxSE2u2pJskHz3k
TX3vsyoVvwrJDnVm93xs8HCeNBUuBIpW87tnVh+Crja0XP0jFBYsss7Y1kE2TsV9
y6N1LmhHKLpiq5TKiK7d7Bxa1yYo74bt6Y2FUQ27wLvOANKNovMl1qpf1oENPe70
f4Wj4yagvrQ0lfwbU3yEIrwuXetnZZ14juN6zJ2sKmnvAu2x2VySGAj+/k67C4g/
2SeR0DmJoh+vbUbnFY+rfmdQXVuBResno7jy7IouhcMVfnhvp2W0VTyKTJX6KZO7
tGs577SjBjQfx1BMhJQJqlVdsO7v4gbeaHumQvzpF/Gg+gOTXrRZ3z0SjBiXR4Ev
9em1ZlaNuwszFPfsKiAOYqAm2ih3nlWk9SlEYJohdK64UJrtaV9qPz8ShTuA/XT7
5iuHwSlWrjBmbTNq2d4inO+3fk1k382SQREzBuWf3kk7YXznN1ZFJQUdRwUFJ5Df
/e4Dj2plNQcjb+jJ7cVVDmHJbYpLdeWkgGz4YZ50zPQtCX5c/LFHxQ0yxXG9Plfw
xdLPwVIzV+S3c0V6zTgUnqJbFUL1bNRlBB4ZTUlmIp/XHHpyFW1MRxkynPSkjmFY
dW+OOM4YEr0ESVKuaQQuXIOpu0mkFOmYyXmj3gD8WZeIz0ry6Ywyw6RTqb0MELFH
V6rehjiyU67IpvMkj8Ctt7czZOEO0NKQQuKL8/wPocABxoNmei6b7AdafLqK+PMz
obI4ycnDOtU5m9dO0HLHrCJP2tY3zvminGFWJBlyAVbuz3U5tfj0vAQH0cIkvvof
rOSGev26RlCYB+cZRbjz6/1IrIeHElSRW3LpzOMpi9DLxNjf3Z18lbxvgUude0wM
g0zNpJvcgbFJsTobT+DYUi+cOgw1QgkLpZRLNEi5/alIBUaMYWVEW6wDZggGBLWC
MZDOUhKxE8J6yY78/BhR9oITEIahopOQlQPgRwiwkq6PgJpEhcGJ5RZQoONsKFJ6
xDsrcbgCJ616oPrI3jiAANHeJHJOFGMorKxidNMiqaDQhWBqD1+UPk0Bvs3IBtsq
yLEf/VkxHY5DLAO/nPMx+vi60oqGFZhbiCLNyBRYvjSxlrzA4u3FQnuUAdJ2/U4W
/BYWJ45HRnsCSw1a8iOffixsa8v6OfBtWWICwl2oZaPiFa/mj9bekBvmuA58bKPG
BZJWhJfVf7Kcytyx4EY+R6LLd7n+WNKWCoPLWpt93jJx71ZEMpEpVCEG4bzP8r87
U3O9QHqvfBYJwFR47Lyz2MGqeN4XYVA7smq7qeGly7FoJz1EyYBpSbQuHz8olUVG
KxYIhYHiUHAtqUYenig9cfrO74uoW/hk4kq5QH+6yCKkmL9TWpJ6fI1PT55ZP8sf
IPHDwRyizqhN9r7JzthkYv1d5/ZypU03hvOVLtjlO8hgcSTcOZS1XHQ/xaZmOw5f
RfOW8+xyD3S0tpOQa/5MPkgFyF8paXWmBE/PgBttIDHJsgRY9iAXiKDoPR9PAuJ5
WM7X9wAOH5LE0H6ZvW0GsLl4dWCfHFDlegdvqj7F1F76gqyqaeXG/iKF7ZYZR9J/
Tgr5J9NM3timcgbHiryba+PQkmbhr087D3gHc4tN2xBdItv9Fl7OpyO/cfAAI4PX
R0h6Hi4HDCMMEuvQw6G0OGjXzfhg0tWAM/ERKgnZxHVphmPiaNf44+NbPgO9bWAa
lJZPg7i4UQuuvZcMVrxkjR2Pj6dWfi2UpDvqEPH3uDshZ8cdFdqHD55V6EPyh40t
nhFUbPXmcCZtw70ADzY3S/obrb0iOpm2ypGpHJUVMkjCez/Fy2VwixUr3H4ekBfv
eg6KnxD7GOjJc4cWAeH08sOmcDEgoDoexd1GwfCJi2HoI73stwycOXgJ1PtVJKPk
Jyz9wb8iof56xQxOjL/GYoYLEWXks60mBUe7fYNzuT0PQmWGFltQU9CWx86qiGjx
yjA6PyDGgBZG3w4zqr438csm4nrEBv7J+ZfqQiWbrLVJ9yn9pTUc4VuynSJnZdvT
UYfSX2Q61gnbi2BlHPvrODQO9BoESPXz1zupAGJRvEmx58cUmx5e6JwBwH+ZdkFB
+JHdK4ncROgC36M3ypV3LFl37vtGYTZO9LEz5mLNXYPY0IV56FSK0mMkuLYxNjDL
gawXLiOoOOYVAaNWocn5NGIFQvXJ5GTfaYEjrIcWJHdf0f2uAuxEFFeosVaPqsFj
2/Z9kzFfUEj8Z2I87+8FovOrOftTVoQepXZn3fbGs/Hk/wJ4exAZXDVG19OzvMRG
s8oRJ6yOdc0WSFp01AfxeREakdtl6WuBJ+KFSXGfgQ9LUuBjjapsoUEn3ESBMzI6
O4yjf3KlrEwH0ZefDTvWnQbtrxVLgkqumcuMkNGwYaOH3jJAUsIOOBIePoU9TQuc
hX0FCDgZcAnIFk3ZTAylE/ZVzdPTBDvGYnZI/QQfuW4TyRVWPRpOEjN00BKJSqVR
kf7vzzRHiYGKSY1Chb/pdpZwx46aiR2j1LdZ98eibrIFEOiKECA9YzBoTrsxN1Q5
0lteM5D9nRysoexZAudRQ/AIeLDZBvGFUR1pLUmz0XprHMCxdXzaXObhuwVxMPcG
2Dos00+J9j4NyCloeFTrUocDF5b5vvCUqL1kYCe98GnfLLNtGA9PNK2hb+Qouo0X
GFBpjpyafD+OM/PmM6RKB2k+1mBhKfhRCKhlB5d2XAf5gHda1axsXeh55Aha5tIf
tf+u87IcAn63AyVEJXOUau00oIk6Kz/vD+3wc/ixP8W4gZMJ1OviK2FEC9LLEqdK
qWMNVs43HMEXipoFwXdRscgWBQkNww2WqU8zzpK7n0eArtepelfnZfEalUkMyl37
UZqe7c5rghI20VXcV+e6s7zijB35QFoFTBuVPwtPBoB0buu16b3zX33Nahi+JMmJ
0HKuNO1iDvYE70NBwDi6cXl5DOFAVahBSegz1e/0s37ezZYodDxIvZDRdzxb7dJT
xpJdQ6AZWBWLF2Uf5UllSGq22mWSgmF8IQurgQAPI1Jjdw/FKhRAvkqCswt2Csis
RJ1bv9U+XnOvkguBqLq0nGb3ISk0ZV0J33fPKTUHRbQW3+8woQ482g6IYt8FkcCw
QHmh1CuA0hCrNjrvsyLPuyASgKdDr2+fO72RKtiIoINTVpI8SsVSOybv9Y7Cefr9
S8I/gdqGCpF2VEWYVLdqcDwT4c+PD898FZqsMwRR0enraOxt3wXNZFBjw6REvpYK
cv+Z90CFry2JkpdrzT1lKgCJnVc4NgzxWqMVZl3NQ8zOb+9NyxfSpZi+GOHxXMzx
SkGi+lDEKpRrnIQNeQj1QUv4kX6t3U4ogGjM2GyKe4tQiXeRUTyIDW5+B2Ooc/k0
hEE+GrjoHx8eJh00qzi6EHvTQ1XD2LRDacaqqfW4Sh9NTvSFum6TF7k78DtE3UnM
Y4s09QT7PJHZq2piz4jgwz8Co6sUiiN8L4xi6J0lirFqO9N63nP/m+gG7qazt83k
Bqd5vK5DzBu/ruHVJwCKkol4g0Olwf8kM05qWiMKvigpGiNH7Rq1tCGME4nVNVzT
R3T+qxlmP6Iklb4hJFr/7j3O2H61jdE4wfvaZbI6okeTQ0rCoX2yxqf4750iXHTd
IcvB75st0or4Yn6zkX/y6FBhpBJhbpa0H/AZ+bEuZXRpimVryGXce94DQ+SZ6aqW
FB6/ZCUmXClDnUxWEOCl0dmHcbXw3Ioq3fuSBuwoaWYmqr3qDwXQguJqltciYqYp
4PpfkOgBRaV/AMEVn4a8zNxyPjE1pd84ugzt1o7MmYrUxfvGQkJOYCO/OHwOd6Qz
gMeCwKEWKqwnRmDWb9IBGBU+otsllrs2PFgiw4pmoX/4GiXH7z3tvPXnbt6qv5rC
pVEyWNzmgO1ah+ZBz2wE6aRtEF59G7gzWEsOe+a10jd2u96tIaH1eRUEQg57HKAb
IvxoBtPy6kGrWM189PPCYqrKXHRtt1JCS/RuAncW77RdrKwMJk+u+zIcN1G84XU+
92AWb2mrKVqLPCX54knrBfglhGEI3ql8lwp18z5RM84CCZtewZ66y5rU8u96Koxj
HHf3v6QldnU2nIacvR5Nv4epac03B+tC28btFGvh+zEZ58WdBuBSlyTqXyL88MQZ
Gw8P+TZxgbS5lrk7Y//u05oYCrd2FDyGzpQd5gvWsNrh2Xg3Zv8w8JQFFzGS707L
tFmf4PmlB6vSk1q82/hfpya6jqo93SwV0rKc8eUvnnbY2jbe3/hM4MCWd5nVYKpg
tU6jq/QVC2cBWvTDepJMbOBhkfiDh7vSSQtcTboHx2+BNJUuPfmBCyEEeljNSTED
fKPkL5zC3cbkRcrzMK3F0IgdleCSA+SaLq1g6QG97G6QYMyh8yu8baiR2b+gX7//
VeVE7fAYSjC7RZpF8VIxYwCZ0X5O0aqI7q6jE0Zw9rk/FS4McAPeuojfZukEiqaw
jMUV5ivhuyaNJY2HpOdM7vBy4194PnWKF4XNpprylZ07JPqvtEdC+Pb1kASJsXGw
/LSeLLKv519IJra2ZVKCfnLP2WD0NhwHvhMdplrRHPu6lTp4BOjCQfMr4bNav283
t2IecCzqc+HTWorajZu8zHCAP6vlgNt5t1ga3mmmIAxrzXnpPEsAQbeGu3yHnckp
GBTgkVhUxzxgzc0flb5xQP4MIKYMrOqo54JcFtX2EOVuAN7NGrcHct6WVNpwLNYp
0lVtoRdjDyQS68RLM0VCgw==
`protect END_PROTECTED
