`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zogpnxm+xqPhhOe5OmtUPdmF27cx6yqw4dEeMr307Mt5MRwlNPgloaLPyxyrYi5n
BDOLC6+p5KXMljchWUaSqPiytzbIM4GBXjgNsOTovwxsvvKAuUtwgAKmQ02P01cz
HnGSaJJTqA8XJCGtBoTw6AnC8wpzNstumFmAwbm6dzjDi4ZWofsr5/4PgULAvB6K
Py1Bi3krFxX4VH/J2Jugsie3kBUsRARcn5geV5vhVVgnZfEKfPvGantzlR6xZMIS
IR5s/INBeiY6GOLTwzog046XoUM90cVjUL8b9LWWt2mOggEsAYhDSJUrgCest/Nr
Tl0Esccq0yQv4k5nTD6ljQyl0Jg3uJnsmZwC4+XGO7fDnYSRJdoLH+yh3v/iau1u
zTB3YBlYsFEn2T9/XjtBPbt8AUndZ1PBTOmsl2t0zlr/KbEJjmlcyZu5tcITna1B
uzVhIFhWmMITpTbrxIfleqIo/KfkoY+ZRmD4OzqBjYP3d0wfGrIX+q/orExtuAqZ
80T75dAK04fg7IPAST8CkJUkntfF0oSnB7conE943tv8+OQ/OA5n8Ql4HiiJdOqN
iC9f0wDWLh7LwX24Yg40i5JGI6aGUMef6LUi57Nx3mUZSvz2qzydOZiYNQF9b5uB
5i8m7LKNddpccULaaRKioypa/MMjOPvw7BAqK0i/zPEapa8hAMBYkKhMo5NAwJrL
MvFYYXmc8ZqeCHQts39QYS9w6uB+RreuiUChMdWU8xP/Kh7ElucqtzsYErz6z95V
92L0XS92flEopUDzVDdgFuBWNHFmulaggmXBG+pTfLY9Fwig/00siRBuHeJLdV1L
zAF0FNwtgmoCERRn+Unv87DfFv0SBCPMpEGvTz92zgtSVzXCbmJ2nWRDenp3fghE
Cq2G9uU8w2hCfuwuRRoXjtHFehEaHVvtTxwAdfQ7cF2+3Pjtz7sqi2iGrUZ5Oyf1
QvODJTHaYFdUTU2LSxOGPqtalolvOEJ+XMGcHiSLe9N8e2pAeiybAmtAcCB3LJGt
ILnPjPTx6IOhRaGmE7U1gTv+mC2nJaXa1tqPN0IHnlJCSj4g8Ds0HvfymoJJO40d
v0b5B9FiawOrGmigAtPFLQDkEMoSGKpyKy2PZqaNtPloyv6T/CpLS99vXSXzDN8P
YGee1BsFNoc0A+uo2BHpOrEVYjn7VHiNjkVXfs6o3LZpA8zshM/p9n8LuSHtrk+w
sS191xRMHrFMlUe6nRIbZUndtSyczxabTfArAcXzBG5kytQwLPyNYtO3ehUff+Dg
+1IJPF6dktH2Vi8o7asOiuQ4lIdYGob1gkEKUXSlGvmm7jASmkXANu1b6m5az3CF
vQjFyJtXdoG5ZOJzlBo1jvYizNK2/27OLm7f36QUgp68XsIfj3Hge+JmxwawkEGx
N9+MH7m3WiNTXevwqN9eShxu7NKVlAs6Z4eXvP9ayrox3UDu4CX9Hw5IOm21nLGU
V64OFd1xwKSWIsHQo/31RxVI0pIzm/Wn3RUUonzursJjWpXz/mJ/kMiRG2FJ8VeL
10q5Usdzi9fVAWw/LdLkXKlsyS5j14qn/PvpownPzoTKa90quLfNlbgFIwzK3j8f
Jw9blgwOVnpA0ctM0qQBWGsMCKi9JASpzSpzVEa712c=
`protect END_PROTECTED
