`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vCne3YFxsK+20l338xkYTZJyUh/F8b0ZXZszq5ZfmaV/grF6cx9P4BgXmaZMhxC8
2fdqrs8lcCBHNvjCy2juAvFQhEG1uC8tJXTdqEm5sLnSO4iEwXVj/O92AD5e1Nbz
dmBUT6U2qauuQgVHlV2rEUwbo0Q+Jlt8eXF01zb3hs1stigdbrYkW3k8QCvUZBH4
a4BeZwxFleeOWRZDubeGPl4pxyCaa0Tnipav8ZbGjL4MeZ/y5+az5VbgtFQJioFV
7bcLuk+6FdRS73bdQ3LJO+HfbHmlQleday3Susi3WfAEcB2xvsc26Z3Hm7fwAYuC
kyb6efI3a2tmtTqpjX1oYI+XVtZBgwmb+lyvRMWCadRcm4ygA8x41g0WiOQt9SBE
PxMSz3HgVaPW9whFUMWek0u0ZAASjJu0w/Tq+5NrSJotAHsAweE2doYsZOEnH1nw
HKDjtgV1Em2x896/OQpNkEbZRK/+cipuRQquS1IwN41xYEO07yIpoEwCxkBKW6KX
bsTki0H7gfgk/uunnrpUdg+OVcPtLC81oo0AddnIuK4/fWIduTx2IroZ0UzSpGIa
gcQoZnbtwbRBwxnUdpxhDWd9WRk/y/60Tnt1aLPmvXV4lsutE8FXMNkhEc9RpHBq
YzDgKu+/88/XRVFawaTyvH5sYhEr6/lIM4icUL+850PVEjxd7mxQFI3XB9AGdzhX
`protect END_PROTECTED
