`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiqrxuTo7EjGUL95IusJgmZJ3YxQDhLX4s7//U6ei/vgaXkDS9PhtSvWMh8DxL7t
XuXBd3fwaCefRIBAj4PFIyZXUoNOGDUSeM/MjBdZsEwf3dQgDR+f6H5acJ7L28zH
LSBW8JTP+S+prnOnXTrD894+XCSTVScsL0rnwGHvoIuGCWc3zM759/zzvfHpdP1V
KCULzM44JGPXAeQWuojAsKTeIiNW7k3l0CBTeYHRDm9jqwP/ZES2e/ytjtz2OUz4
H6IyvGixhAAVfYtL3VQDf3DRrpYOA8dmwIJ8tXggcEoVpLG1c/mgm9juesU+LTk9
qYLwKVzmHb+Qf8cWncpq7bc6qZ9Cs6WGYOs4plGhmS/z8hlJHFSvh39CSdUSs3Al
qKeqCT236ZRYzG8pUwUl+OYatg0XpCqBfFG1rbd/T1VmXe7WeATiv/nnSGT5WX4F
SNvdyZnK8VtBB0ZNK0tKNpGqDi9Uq9VEnE+Uk1zV9mT0SZ5sc8g8SML0xxzU3SiA
g2XsIS5ha9Lc7ZhyX25BhQ==
`protect END_PROTECTED
