`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/tZpJ7Jfw5naS7zhxnm3LuH9a88+NjSnWreTL6+XpdAM3edqZPmWBm5RHppnEIm
wFI+kT/cJlJ/+/Spnek06vvCdoKdrLq9lnZEp4hwuKL0fmeuNoTI555a7bSNM/zC
ab7Plkvp5D7sycdp7T9+VkXbmc8PNkiUQ068X4mEee6Y5dT/qw2B7+FxkPLj7UID
ytV7XG8haMs9j8GQbRSBgE0SLH0nMGsBlca5A2Lr9svq4ZvYSQ2/ctdii0ckiz3d
7yE3Qab+gYWhxukk18n6wFTOt3eXD3U6mqqCBw1jCQ1B4aTYDJu+zBe8B4GD5cKO
IPJybK0zy+fMQKALJD+uWkggFPbZEXu5FV+TWjvALMNVo2g8PxXfSMmz4s0200Nc
tFcnLznfltk+sbXFUrWcpEr1UMPxGeLnsBkHY6kWUCBj66oR0PvCEjmSpDnyVT9J
2xNPWRgXWNsFuj8SXQnv0NGVo9uZ/MBCLTdEXVFUl+F2bMYDMR9NTES1MK1sBLWK
a+OUD/aaAtOgC2fAN9GeeIH2MkIX5Npkf1plZWWOGoB2icB/1dLZYNAVshSB9U5+
w4dfDIXIkZXyeMfE2SAkB3KphMuQK2w3wqCvekuIXl3kKoZFm5WNLCZpIv9dF2ZI
hBTlAUCwWoJ9utPsQV35pGFImQpn5skHl9qzEcI2GgQ7N8ew7lYgTCUGvbi1nE0w
PNAETk7EbaviRL3vq/O9ygIyjj125jKX9bfqVw3S8Qeg5a3zw2WbbfE8MpqCq3Ej
F8xQdMj/ufi+cYkvJfav0p28wkuTjlO0pUOhGx31PRgS+V7HJVynNX2fQ3mq272z
DNxjOVDx2ItZFtqpbG8cKJR0QkY/pR7IjN33nGR8fEy+hUnYeIYoiR/OlsYmNmD6
b7TmS7ejSEJcqbn6m/lmIk9A3OwqdEYOL6MGJZONzjFutZithbq1k/Wtmqr8UG+7
TpawNMJgBSQUdH5Pbk0F4VK5tk0/7UUrUtvNiiKQ0C5168z7bhoes3Pk5un9jzR0
D/QrhMBf2UQODwPaiKdLzA==
`protect END_PROTECTED
