`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rutuKDNTds7mXY5EoqI8ithLZ2aG5IV75uHqEbdLT5ao6cExtWhrKYkU3DXWYiBC
glC9degVnRDt7CPikwbx9KqD96HPuIpGOZGJcKWvKwiqJ9pmR//KkYKucVxpaOzh
t5Tf+biKI6TaVEYIvOG1mkaIK+aAMyZKV6GLNoo3ZePq0ccvB69pFm2gsMywi0IT
usWLhuKSuMRvyNbh4BImgI39GNlpIPduAXAx3RbLRgERSGRAnvR7HosgjaNW80H0
NOdzvkFljFrv64V8ZCULgQ==
`protect END_PROTECTED
