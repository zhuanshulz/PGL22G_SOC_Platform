`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYKDWA1VRtqH7ZmwAiO2GyFSwej+zKzgV7hU2NAh/zkABTeisfg5oN4237ZQ/Y25
jP0IiGbJ2ZhsL8LiINNCHJHbBIjSg79dEMTXaHt8A5C9UnHrYdp8AXbabO61/0Z1
CQJFyiyZ6V+LtNZ10u/y8zQq1m3DXbU/m9KCXCmrOULoUD/85nCEAj/1+H899Up9
R1UqG/CviGVp7BR6zgfNT1JlK2xfEIs1a4mQgYypC07k0AF2DhsmMsdwvHvG7TAz
tyrbd/bTrv0gVrOmEMnNprY107sMSMXIb5vxpItTrcDydL4sWCQs5/oDX2Cv0HXH
4QngdjOzwKx0ESU1ZltQj1MjFkv93iqd2KJajtlLFAtdHcY/OOcoBDyTHuu3qXMm
qmJDJNF0fb8zGzJqoK6djRYVVypf+dFslFj/FTz5SH+/2orHHk3APMa/BOjFF5MK
PjhArPKD8I8Pd3kVNu/f7Yq9qhbVJQgkLZ7MHfa+j1ZwdkTwjMWkHpH7UDboIo8Y
wvpG31JrnoBXoKmHABfah20rmf8yof6IlnJFHCPUtW8FpE+CRjFoR4ZG+t2lCKMB
hZnkBXFzHurd+LXdai5f5NzsH5sLC2fgS5d14rB9k3Cmf+OBOSpGEiooUQ/dhSH8
jOpMuslT9yeGF5adgd53B8XhJlq4LdXLdUaK9Bk1+5i8VLB2+k4OMi2Gj9cU/ike
zS25kZ7VQwbyz2sWej2/Tabo4YPiNzd30xzwiObUn3GDvtGxQaSgp1FUagMZeNBh
H7fo9wT/gO1/x7yQZL6PoiMycqJeRJeOJ8FCOILZS3HYV3k7bAY1gLZnFr0FR1cc
Bc58SvsX4V3YylZxt8QIA/P+25AhqsFrKtQlvk4eIzfBs+7fGwO6QJfEJXYScYH6
WXax6kHocAiVboXrlk2N3t6RYF4MdQOllYQCWcHjxxg=
`protect END_PROTECTED
