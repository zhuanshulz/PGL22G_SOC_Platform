`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sC0sSsphjITZsK+cIffGwtdZaXNPzQC6jtSa40Eny/0N9oVjY1Ueyt4gTn5/CDfb
Ye42QKBcJUG7zqKNovHw2AM+5UqtDX2vZ56n5vqVPIsj+GhgyuO5klD5sLeqgdPN
W0cFf4pcHj85H0xXaeFT/PpYQVgqyL44ukJSjDLgF6DkiNUhSbznJH5ppCHlhGBK
dkdyn/yHtcYKdOPwUWXkbrgsuwbThHigPUl4cdLmbQJALF6o2d+8PT4fs3VeElwO
MYLBwpRwPo3RYqwDH0NeTi4utblBZr2P4TaQuPpP97Wm6Wen+lrMEyr0+Jrn0KXb
C8phJJrlAUHpfc/JMeAcm+Jj39D4jCvcF1dy6Oc/GtJ5odhb/Kk8hyGRlFlNbcw6
9COa0Btn5osaGNHeWiK9DWe6MA+NBRTneSKqt4wingVGuqPSXj0tfuY8LJbeDzOn
V5E1f6ixCMc5rWYAlhe8pzT6S4b5C4NeQfEaZOmWNyq+5jpVvdBofGULbkQGriix
RzLrxtsJHtwWA2yQnLLk40npGufuwHX8BcNRWNf7FghucYKiSf+Z9G4qk8yAUUHY
5vPEgg8WbA0jppQMelJfzstXXtBjrkaWwXYsGEZui50L/6Hwp2UOA1rxKNY48oeh
NofFaEc/uulqN19l/JccynYdBp8KCHKkl/SK75/iqbyDYk/G8Zj4tTZCljuy7+3x
FqtBc1E2vMvNVoKW5/XTJTIBDZTobTYjTngTqv1akPXrv2DzTgDpRonvknxboi6m
NJQOAtU3fFZRlD20YWNkEhj2W0g55weEqAu/fv6xzNYS0uBaY0WoFULC9IG/x5/P
4tqrenORH5DoRPXesvTQbTN1fMkqk5Z3mbzyjkZjzk2oJe9rMzjDj2YphtJkhKgQ
T0+xenRy+09UmC5KENh8BPF9JkC+Yu1F4NpIAveEwZJPdCxyURAOWeIg3GH4XiWR
7cEi5nuhLx7VMg46ZpBPtA==
`protect END_PROTECTED
