`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+zX7YLtcvO5+Jiwd/530Dcvd2v88XGsVKW6llZqBEcwonViImsW3R3i7cCYqcu2
EP4mms/ABvl6e1JWkghrTaza0NqN6jJxzAlCTzEMln71/RKnoO1Z7lNk4f7dZzJT
7/LAbF6nmWnuabDFd+JkG1+KqXDjLPYtb4Mwx2s1jhppfLeZoldU+xuI6eNXpFZO
TnkNV5Srpry95BFZLJ37rMWejO/YRyEWDVt9xaBe0JYWMXSuKn8rzEIJuwV6T513
JSztD3MW6rs9HK3b+HcdbBCbvKGUzDyCnY6EavN0oTy0pYlOSu3WHDMegcv41fE7
1WU8txLRDfU5H7V9JFV8IQlQnCbET0Zx8HTXjmaEcO7roHrVBgT9iUog9Nqqi6Tx
fINNWmsRojr+K8rQf6X8ACTArBo+LZ/YJ0XywDJPh/sMwyUNT/T7WQ2YSiB8f0V6
M2vwwvP1+QH6oIMzTlweIIpqEG9mTwGwtxMH7rDnnnEZn6U0EZ5Oe7aB/iLk5fse
t60CcVIahksQ1GH7MD/Ex8acN2mP5DuNissqpheSgTqxSIE7PNEaJL1rHW66SSHS
jI8RJkGgMiv+c4DfVk/gdA8MRPfThHIPOoYOuweAbVK6f9GJnCfM3EoS+1ayoGCB
DuConxKaPvYJQUJXo3iXHao3729hDwaKLlllM5UjVCrBNaqBrDZS+7B1Mqj7U8IW
agMFAZJ84JkzB/qugT5AvX3piILWE2mHaagIsUjJDA68JPgC4JcZ9Mbe69hZbp8W
z4tu6quQq1hJRNqFwn6vP3oLsoxpFKB80DZ0vDlPyx2sXMX33o24N23tPKfTXCCw
ccmrBmmrlulb/hmn7Zbi3sooS58RQv+0Y5cMiY2lY6f0B/BNgO4uA5uQwZrlLq+F
jVtVZTV8zDmvSS9Ntowa+NCf2akwLldge7ZKk/NNtjEwMXDEBoRbkSMNyLxTAkeB
Hoz5FhTrdxZyYgfL390IsLwBiWMDMG+ObZU7/TsJ+m+kof38HQhg9jyZly2n7wbS
5b7GDfVcG7PGKeetLUvpcVgdNIjk8aBVpufUNziTbbOjMEWd5FdA87+LyQBZVHqP
t5Y8x8bN/GzeVnvlZ3yfqh34i9SRAd94bBUr1if2lcu7RYBi3LeJE2EKCZWWhkeI
1LhlPfuIevdJtnx/YRAQxA26U5TgLy1tcXTEEFK+XyX4ZkM/dfwES69LRlOKqjQz
Er2j0XP2uQuS2euMQ6lut1ze2/De6IweBXH+VLaSaRKPRWSKfjLqFs4eoJkm7SxL
wd/Z9Ag05mQV7yWoA6Tr1mVtIDxJhjMi16nyIckHYxM=
`protect END_PROTECTED
