`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4vYFSaK+0hUiFBTWqr0OGOgH7MJpOEQKTDSsxrbQAKhv49P5YK/o+WVMhhu/m9W
v8/e2AkgNrkl8oY3r/j7Ndvwu/F3/K7IrhcUMYwm4jroDoEBlTXTDhpPgVQrPHkl
boybGJGdOkzOFqYLXDFIe5g6B8GySo6zrGWdjcJCEgTbw6hpIk9V8pBnVhATj9BW
8UiTesVvvTG/97h34D0XW7T2/zGTZmVmRz4xiY+FoDznLi1u8u9reVJYNoeyizt5
/E1lNLT7GJtwRvArbBP6vkrCHXl2r1m3rtVUR1dX+lO5b4xQJBg/z+eqg5FD5T77
++/LCZoCh8p/RUnip4qIxxxMB6nVBwH5wcGD8qNbmKn34H2MpRdGWijqCCUVGj/2
M74ZMBJNuGNEJz3RM+yXOzUl22cnzykOvn5V7cK0fI7uaXUv0dSik42s9BIJXWZq
5lP2Vc+FJNoq66RcRiD7heOcyEQiqFSrJBbsgIaNr4782jdYNsRfeg+CpDbNfCRM
CR1xWWtWK/wzKy2j5QIMq6Z9Q2YdXuwsuV89LLX5z19dr8DDfkBwQwcS5GAqX9rm
h48fxOxD9zJvvlH8n6FsxMM9tKrmwmfAGoq37iH/C7EnBygynifuZ0Z5JtKLjJE5
0DUBNkKfk/MJk74QDNq5qJA91nTzLSkKhb6+dh8Je894D+dq8SlavfXiPA3N3OZe
FbPHqHA5vFCeKQ85LDcHbcGI88oGX6BivqFhiaJYw3aq0Yp/hPgBfN0OSNAxuG+8
sf2LAQiSUGMa3NmnPTwfIvXtSr/7wLAgVSQpX/6YJEBgkhqc23uIejyC1Gs+9Yz4
GkSArJNGNp2/MODzSv8QGNiNj+GDAaVh6Ag14b4166JVOkNM2vpVyO0yp6s21p8c
uYJuDX2uc+poKgYB43OrcahZkypBKwvm35814CCIvOAZS64OYPh4im70nTO9tiZh
kQUJAqnkB3G7s7bMRQ0ixzA1SGcZ99hz8UBkglUStHXkB33GY13AR7afffYVrFJr
k0DXi0tfnohS9bzJ7ZiGtoMhUqqKas6UeOGb/2aY97RTeQiuMtFsHo51uO85J54+
TeCUZ5qzW73vVicKHvyxAJEa3KBOiWBcvDznUgQQ9fwb6UiCvuNTbupD15MeGIsc
7AXUv4N4iubBtWx3INy+alhMBH8wdXOs63uECmwEkE6xYLoMyv52DNk6yZAdJ5Go
11YWAKnhOn9JgVx+9cbwPHS7eehzo9O9476crQy06WE4o+F2e1GuQIcxlPCT/u5g
ejALFIM7hg7wZxaJQeDnLBqx9WlW0stTr3KfqkQayUkeST/fvdOjxB93uaER7TGe
BL8DUMIHJGIBK2tgBgwR8mFa8fSuqDYtgLax6+JOdyzT44vYxryDhjtwn0h7C5v1
3gTDa6vZWRzqSF70nCPVqS5xlxCHsQHaJP8oZ2j7L6dS+hWy+cNEYRYhhQCnH0C7
tKnBTqmnLPNXbamKjQoPwHWDLzBqT+1yxdaSsyuUQWEkPm4446e2TWwGcngbMjHf
Xd34PzTQB7PqbBn+TJutSh4vA3GFpYyRwztpvLQy2SfTtIROsYkfws6XBITJURwI
e61BdnQAu/VwSx2p9LRsWUJBeFYE49DfCFvBqOG5DoCuXvH4SYau5flbASa8PCbK
53MQwdYWDl8VP8cvnCgguEeiiRkwg8zIMiNchj4P4EGQOodxShRiRyxa+1lVCr9e
7LCS1uKXjRbsHAjb6mCLAAqsdHT0r8QHHEOVkrw3bxXu5QIaNdjoULU65JtXl+cu
YIrKpgl8GRR5bMsAUm8ZewK1nsPybiB8mwtyXUecKkgPH+NVpEgZXWNJ5432e/fW
ArtuVuaVRXurKEaSfNe9JcZgK8jPwkHG3A+rLh32FtZUzoVkpFoObUMwhActfilg
zY2nhBdQttLElFj/TKEDUmctELSlLI6xW2Zjstw3fpPgkBhGe/Ge7uskKzJ5I0l0
oEgreVkAJ845bfwqrsjr90zUhcpU1ZKuT+8hk2iUxpWxmA/S82yQaQdqA4TZHGyv
tmUCedeOTouWaa+XBpHLLCzyLW5QyevU732s2QT+h9Ht3gbeW/Am7dQ/qG1a/I29
14cLGovNuWMA7Vjul5j7/WlusEBn6eeyrLd8VULbvM2UcFfUXQ7xB3lSlzBs7kSn
sMmALzmmfOfa0Pnr8vZzaXStyLF76R/JjqmtxtRB9cNK/hVgzTynVhXLTph6rKIB
pXe/7XaYAmxrKvLMXFTfmrLikUZbgaAzD7eyY8p4mTqn2Rr+ZkPaLKKhhnBtfLZa
rlh26y2PJBpOBk+m6O3oXVqAhFJrJVjTgIZhlvUucWBjp0zIYTvhWvkH3n7OIoka
X6tEGXv0yKWI9MRa2jtz4UJ5p99KU3OeQzuxo9Ukbglo0ntwFPuroGiiatD5abD3
ymXab8FvHfcXb/d+8JmaXp24Skx5c1mG1M9/JXeH6rySmu9vpvIlYQlufZKTJrQz
rRxncS05k6yb3S/lln+FCaMiTRrxkfmAavLPoAKqmsYNYBNBEpGdd/wjK5+aG6VE
tkj1TRE4f1FRS65KdAx0bXyIuJe6KOf/LAINcEKUYU4=
`protect END_PROTECTED
