`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
naUapDQ2Pc5dIMpRDDHa6be3F+3nTGwauJmoxb8Un09amC20aarAnaHGuGoOrFuq
qC4EysDEa+/CrXeX3pUWFbYQ5/ABvupmgKtt71hCs6pdp6UnGqaj/qRLLMCqUs+w
5n62qnexsef1jqHJF/t3JTFl6SY+HesTydFscv8TXlA/xkSIA/m0+YdGInuJ9rmU
/kvddo6EGcUPYJeDG+8jIzT27G1C/ptoUx5dNzlrZk7TMSbJ0+E+V0kdP9oU7b1n
o5ySRst6Mwc18X8mpvb45sB6FJYaFtbAajTXIA5nJ7cOXBL31UGqwIWcjzrvFpyS
UrSWeY3FhuqqHz4B1Ri4NOu8vR4kgc8TVzm1EC3Ay9T+lJgxqfVdrgDmA0gEl5E0
`protect END_PROTECTED
