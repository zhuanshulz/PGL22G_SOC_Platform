`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OyMJ2sVr98+eTz+Qgnx7lTGj2ei3xp0ZMIbMEaoQSh9QVhG622gJyxBCk5Fo6N3z
M7Nrq4hiGl0qn3UWd29gGqkaHv0HqXdLEJjtNCcFPkmlYcCp5DVn1aLMbCnbQdKk
qCB72nIKjRiWree7eoJpxKFaR1jLtQ1LJcBQg42Eb/kvww+rNZa2qpETEsbt59m5
19bGTmiar7iZV1NgpHehFSsCblvb4rHif1B2n7feZ63qWVaaHr40hMfKbwm3YHRg
b8FWrK3LPUdgJ6lWVdCzMr7wtPaoQfj2py4CLpJ4jLKRIRapIXwTla9pCyZ2hOQz
hpJCuJQ+OLaO8gixvnyEweVPLuqlqE17BR6P9zQwpuiivfPF+w+bSdmGKsyIzS0D
gdeDqjoo/129doFVcvBKityAgizZZInqKFFLJ1XymfNqwc9GEVu5Pu2UAJG+ZtQv
W0TTQJVUailUlMwnFtJL0UlDwKjTw1InvtB4c7RhIuyBwt4sf2An/ltMRbWBFvHm
Wl1bNF/auSVmxq7GkqKe0L8UQGlyTxZvNHhTvlsrArQOthgMV6AJ3597v0GjzrYA
AXomsurVgCWigDfy90YNa9ooZKlBv0vdJXB61edo1SWQf28rzzbQb/mtJeKG+GqD
R00LBW5EFLQ2Qojm7oHUfrE/gDt7OoABgOj/UCZydF9TFtzb2xXHoFvl3EdKHTSa
GruShRAmd0BfFwPUH3cOqogv4TBQW0ICsW6HfNYpUf1rYGHMFIfz5aZ0MNSqB1sj
MV0ipVBypef4LeOmaDmgEPFzhMRaHuRCINmapwSHbSgBIDFmj9q0wz4wWoklJ+bX
T6BJuHULopGfmEqzDNNOWmdd6/nhj0LQ0v/a+0pj6367miwD4ldcHv8mW/X+bYD4
8gldnMaFNRNe5cMtoC4+g96awZufgSuuBr4ogFzZ6Lukr2hb1+P2QSpkbEqJUXad
IIMD0DszZecZQPIiIOmEGCehXK05RKGUhpaRFgHOkJxH1N0nTL9KDuw49PfLe99n
8aT0qvjxRMigIRHwMXxdOjghZzK0nEERAlZWT+Xe7tJiEuC0U3NbEqua7Uwrnoe8
acumOY41SGnhyX0ijHkaoT9aCFm1m6wR+f4LRcXXK+MaEnKv7fojgfO7Sch48Tku
GPJGf6F6HkUewFNNGCugvcxEhde+I4qOlXP5BMfei5tp2L1ToTf5i1T9X3A8zFiw
aAqGSUSbUoL9R93lzfn/0278xg0sYzrGUio+M8AAYbfXrw/tpzxKak0ahz7IGK3R
PsJGZ6bQIVlg+bhCIBtAO08//WQYwkNEuxTtg8u6T0zmbnZBN03XW0LkkdAUowkp
wwz3rqZrivGWzKvVKo22PWYi/DegnEXpuv2yeOeGHacbLcPA8KHlbECb/lkvJTLm
5HpVmjVFK/FPi1US+oHvDzi0D7lJDWP2tOEXpd7UApAVXfE5UyI7Z1oFlWxSWgZP
resi1s7spRIoB2vzqMd+z3MVjIToJM1+H1By6ZhQZLIFeR2oCJT2grQEMfBXNNtq
NfuOOdbk0yhOrCM2Mto9HPF4XJKjcugH4/Ob2fPStIzkMcSszwkFfM38GKxP6LDI
BecldQExu3IElquETEryZoQ38RSlRX4h3Lt8wFG1rZcjOM/CgtXr+7iGJ6eScIsr
uojDVYcglEOSszcP9Byf3axXLEOW+/TJdZgeZmBaQwjT90id0rPQgaQmTKah80Py
0F8xMnVAFQPAdQrCuGIrTJqtF6OhqW7P1N2ASTXL7THD085FdTf55pF7VXYI+uQn
4XIgoCxwHwAmm5gW9Z5bnXkidjvcB/kyruQS7JelMt+KT1V/bVDVnauqyVNWQvRT
dOBG3wMg7dWJQkLUvjpKnZgB5Hclz86mo/eb9bRc8ONA8GZd8RXTzNeGHwlIrUSV
KboodVJXI8a/lERsDL5m29SBlxxv+NDYxv93Fzq3RwJUtivH5CU5OsJVVljmdcc/
fj6+fIpDeBD2qVACK5h0SDIsK0iBIcoPinGRC6PpH0TSSOlmN8GQRtDi+WaXuvcx
YZATEIViqp+Zz43WRD313S28dEU4UURiQG2eEP3JnL6ogbqwx/yWLCLeae5hEcRi
JwwQ3/4ecXleowOlCzCfbUvtdnSK+C6SzJN4h469e/Fu5PSRjRhhQUWD/mOoSBLv
TxvmcRr1Zg7ZTqKNW/w7yGJZFooeZEmvwWh2edTNq8vEjCx3y9PEKYYb1xlJNeuM
lBQSVmuqiYBz6ZTmLJO6qcbNqHM0Gb3IcrupGUlv7B8Ix74fEU9K24igGhMhALbk
Lio9DcllStZaBwvQP/c5iBuFVcTNW8YJ8DjP5sTAswG24fZVxmkvMkgkyvrV5wTw
u8Qa9LYwQd4k4qFvITNMIaUXPcca7Dtjjpoemw9ZWux0pP+vSO1GSgA5hLR3fPZu
uclQBxFK647koFCLSti5NRhAPo7UZENEWJ8eMhrD7pA5JTAI82zWANRvpL9J53Le
U5uNciQAJ1fsTFk5sLMyCymqSv7D4b0lWxZhlc+pyMbCf1RlXG1YZcGXa88bRciL
YiysfN0sTyu1PSA7F00363K1vfiqlnmRasd4e96JnHp99R7NPHFLSDj/kUedkg0w
jrFRwhbZr7MheWtXY054tCHaTilFbuYwzop6vujQAGi/8xDNkZ3fJN71FMo19Nh8
ZNm3C+dWoZGnsE/brKKShOz4Qy+IrKbjmPP8jZn+YeyKoJEtI5T0frUHPQieBAfW
RHRhqDGKwIjPg6W5BWQHFduvqGRb7HXBAFNevYgd/pDJCZU6Gf8bxi302zO5mPP/
8Qxhu7oVLRYn1FPcB2O575yjoeUC+GSLz+2kDWN10penQr9ofWDJt3oR8qhu0z0D
R4NlVTzU4dQ3cXn05dPs9+egeGtwNdDXYMlR/byA6f/Md8QeFv8UvAKkJz1iUmdk
ZEdOemqlm3W0y2AVnXj4iQ==
`protect END_PROTECTED
