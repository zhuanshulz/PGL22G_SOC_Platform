`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVPvXRIdgLW14FvtGLYwJm5l/FxYPO1A438Bz7Cd5cNcKZDZwUvTQp2D6D5sX3yE
XnZ+KbBdzHbpH+EVNWsR/yohsC/gKHcCE7LVUttVHd+LMt4whw6AYKk2bb6Zk4h4
L1S9iNXuR77TH19x7TA98c0XBjQub0KS3jx5yPAYRA+M1+/ziQh5jr0eZmjso5aE
KYhjfLrF6U+c8PX8KyW4sneEmgIOBou783IETSCoXtDJmps0jPWZ8WfNGIKjwRUo
h/l9ErLK9LjLLwXXIEqRuEOSS8CzngWboEUi/vuq07Q1519Cp1Cq9c3IByM+pHvv
l3uJBwgkTPtFC1AvMiHlbmDq22gyYbrPxYeJrbZ+Ls09c1P+KsdhdXPCuNxRE1CY
32RQsRj+HnIDcCf0v1na+WhdrYugmISFUKaatK0kvIpskGbMjPyKUaOJ1EE95iSI
v6vAgcNFvmN986fX4aoTxTk2BnZn96OUULCb/y6A8eoxWkn57eVD+oM87EeQzMGb
1hU2jWsYysdjEmKTDRwNIwMQUU9wxpAbfNoWzBVbmtodfZrkr6V09wnvYWtlBBQM
oT4PTCgmxtwXXsVJ0ImLdO4AR1oB2mlPEO6zvYN7Yu2al9EVFgKIsY1QcPidOrl1
PaFWa8A1YqkaPvmPpoHywj94D+D5V28zqcKplRkJ0JA5HFWscVUpeW0UGP/dHfJf
6oD4emTBjmdnTEQlzisTPTweEDvllNmUiJg/Ay51mXeq0/79Mixi54fylpdNb7aP
qNwuS8BUrqgl8h4OyS1ipw8l3+LtWBBIEkK0Cvyd55LxD67zhFrbIVMNfebPOPMu
3ULj4anAlNnd1JtupFsZsYXT2ulxBaytrkuI5w7V1OUTB4+vFrBWUOUYCl4uyMF6
4ZcKZYLbmNXa2hlKNhr7wAvJUGaPZsvNCj0eCMu0Cgm1MtP2kj5CB/GPH2AG+uJ5
zsSv+4e2IJphT+USmwp+pMfxuG6yWiXOHGXhrlLcFW0rrrgf6X/+BEbi+pVD/e/Q
S0T9VAwEtYzgfd/GQZNeh3WDEtPiBNR/wRiN7ZqRwwz5IfLRdMYkEciQVPF5c0vw
oeg4rSDjZUO7mqpn5OgykTuGOw0EpVolFSMrseu1f9NGbQ9JwrJoBfqfEvDxqavt
yUH7O+Y+i1cRW8GHVBRqxSK7X84giedzYRL8FeeYze7pJt/2aPivWrIvrP/HdQHn
/iE8eB/A/bbXOYQooBT1N5Zvm1HOlIugkNdFcDDN9ElreT0mPlk3+f458GW/1+sz
uGU/Yajlk3M8AZrtpgnLM0Ncy8p5CDz4C+skAzsSK8P9c32mp47IibnU3kED9Eln
YSo7nFVmkz7duc2OTI5coyAc9Zsv6la0JPdJGLOG1UYSZNnmt/5WCEHazYvaKG/t
0zwzgRC00O2JMl3Db1E7ySqpnW7YgBM8BVLEolYZswk=
`protect END_PROTECTED
