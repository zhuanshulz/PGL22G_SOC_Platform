`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MC5SSGm8P/jtt+HwE4Sze8kg25Ul7JYv/O1wk8OXksXJZyopahB2JWUyU4ztqDXY
yKV2llUlYg5od+vlFJQSiKQN8J+/V6vcpA0JDiQ6+KIrdGa2P1Zfkvd/3VbIN312
St5UJLl5mnoGBgAvyaHBiNBh3ggGq5Vneszy3t720z6kFR7uUxrdPHD1HFCjxbV4
F8MiLtL3NSrwK+NGp73XLdXlj/Hahc45cRN4Chhz68mTYslJFKqOuGZP4657EuAH
GqWOvtOQYd8c+Y498O1EB71XzLgrUiweYomtg9iHeh5hoty1qg3iT7NdOOdj3JN0
vYLcbO+Yy3653Zh3O3unZlWwmlNJNlZZ/3ZpxM+oL+wDgN0rejTC1wPig6yZyMWR
Y0C6M5ldskPtzo56ilrAAZalXJLGKhLvSF8jZhJP2ONsxivalSCDzNzi8T/oseOo
C5HaQqRRlUiL7LLnJLY2mC+zLEyD5YbctkMmwhI6eDUCEz3AfZcvXMfD0SXmHVi6
wd3G2/ZflT4de3rEyfOT1sxcg6t0rHM/F/5NMSofft6DSSjJXc0pMfUw/t6fwBB0
xvCnXoqEWF9r4dGtO9UyjTHoJlJHeF0Wbl5zb/pTdwejYzaFKhmqDw2ZgsQYlGwO
`protect END_PROTECTED
