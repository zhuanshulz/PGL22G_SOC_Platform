`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hm06ewten6oea9oNNuo2F78ZxC/n6RkZpgXOmr3SBxWd7sQrVdBRxsdO4M+nN/On
GC/ib6P93tbwUsQB9kikS0OezaH+4JatR1id2ubnqHxeOHjz/jj6aipDSePN9s3F
jfEtS0Jqo+3jxxnQrpj3zbet43Q5ObJn8S+41gbNbhoXBvhVxGbB4FZdD8CAPW4Z
XFDqA9d+qqXftEc2WDlN/O2qMkk8xRhk1qf/a/OcU0+mouAt8QsUJ/xyGtvbeO+k
QMtuBIDLvJzuSpdC999aNPRX1erikQSyfGRFvEVtwxwo9IeGzV94YBEgug0rZu+I
YMJiHDo4e0og9ChS/FQ+GFQJy/pojy+HcjQKr1X5wVPg6muyYGAfhvrMbys6ikT3
UwoXW9y4nkC0BUAL0OLioLtDx5vBDd091F4pqIhDt1R5deZvBmeM+FiAS9zt+d8T
iOQaKOqzpbhCshWq7lG243VP112OuhUcbODom4308fWDvsx3q/8+uvwU+BjT5rDv
0dtNcMpPm+6r5DbqmKkuBnzO3jFG7IGyKabNSkPP2/lEucCUda1J17QeHCjPHNDH
y2CSiXy4Pc3sVQcdcDqpfWBVgpEWaeNp7k3vFeCTzBGg/XpFR6xvEckJUVSpaH9W
VBqAGeh00wtT0HTEd/tbHcPHySZjaQnnIUjkJ+st4H16zO1/M7y/j9EnnYNfXs/0
2MJkjHNh1huU0dGasgwtOvphQ6g1976rAorsqC+FGIWGoM6WgWsX2S1bwg8gWH1D
l9uqKFqcJipWgSVjD85F2LbxDc1sQgU9NqExyXlf4z66gLxAmcoIJ0PYIJxlnKEG
Qgg3TjXCy6DzAo+eD20yc5wqRi6sh/h9xY/2144yD5MrVxtDPXc/8/VYhmnJ8M7j
KRx0kNsY3h7YB9hOElYhR5h2P0d55CRMGjxPn9b/QvZOz7gA6tLPORdPtcEpa7kU
Wtu0fdui892J6CcFT4Mjjvdz8ABWUey3MfLgDhsIjWgCT1ssGkrfLumonsbnh0YE
y5suc4I4VPZiSYDOwNtv6Oa/3fuT1uajTR7gS3jwZA3hUfWhy+BEjPZawcS2xp7k
mb1ry0RcBJxe3KISrtuw0liJW9/R2b/07G+kzO0BN/UfP3pBqnYpbvXKvcoWVKcc
ASSilV5Q1LsgDgtrvgFlatM7ZwkTh0JR2PXUlNBz6jXO7wSvZ0t8gxgttQTPZ6gq
h5hpW0hMBmHC58UknjF5LgdTMfH3XV5ilPPsKoKEZlhhG03GhlJRgdxRo/qjj2Ku
MJdjRMKXO+3zw4C39Vb4SpF3+HI8rQNRQ5AwCq9M4q7dc6F9+tCN2EDYgc8d+LFi
x81zKP/z4XO6yGAxX7+rZQLeHmB8hpAYqYPqj5kA9kqvZBFqTh8/TkDqOs5LTsF/
6UJihP2xcG3pLsjjkWhN+Erj9EeBPfWFABT56z6uVnMOSu5uZ+64WBx36/XsbTqn
KqzsLl5APMHUvCK5MTBQexQCIc0BDsdnrkxfsidAx1R3iSY2QyE42t6w535gsdgp
OouF9KsUIOc6t0r1JAIhYpankVTx+oYmaWQd/poqhaHZo3CIa9YCuOKFcRyKADVn
X9Kz0B9y3jYxywYbAcIjFbe3nSvufU8loRHH6lEVEg5xLIE+5Fz/i+FBaPDZwsrk
71g3uqBDD7azGIU4jRYcx7kgWFkb0v8nX419fwcdT8VmTBzEIga0KK/hdwlW6Q3u
EOoA/IBE6wrHS4/WkR9xhvIjF+jr5ZnjZ2360OhQt8NUc4semCuzdikbHk/I7uvJ
91X48tdEVEYs4TAx9m+VDPu7Ems7AtYmzL9aT2yOwbP/1LNkWhrMnnrZK752Nlx3
KkQ4FYU+sRNsyNBzN1zSLkQ749VD11yClAPbiAXGWmMIrKphyrx0/P3cMfqLtDip
TZE1sy6Ncs7yGIvk5g5rRbYgaoywXM6ZUgooukmPNuMUoBVuJzBWUp8vM4ZLFkpH
ziOhKS4ZbdW9/q68+z+SVllgD8q7YgMo5uC2Q/ZWlSj2S5XcNraBv6FW8JNr7VKW
T1RQwqtGm+tLNvNa6ZLUruSiTk5NIoFYGmT3KWLxw7KCDCBhnuTeybMmmf0VWepW
kMcX81lL1665IJU45u+BNGVSu41ms44jJGNx0tV2Od3hTbDq1cxA756M3QyI/1Bj
K6fnh1qpq/xm9wkL/xmaG/jJ6zCR7wbVYIyZgLxvhwh/FiPFH7yc4rI2f6LZ6RZW
0CxfclhFKuqPQacCZSWCL8/ZxPCFv0d7wT9zJmuRLnozsbUVF10MpmCYvZA7m4lY
7DbJVRvG6u0OIp4iILDssOBy/sjDD1M+BbGe+rgUS+SenHR4wX9H0eRQeatYdyMm
x8S+2teCOYeG6mmCUy1EUcZsGoU3f6WpqTu+g0khKmD22Fg2e3zw1ggS8ktv7l7j
TZrYPy33tTLX4qlwsT82qt75v9ImNbG7fDgjwhndcUoo2hSCGed/sy60/MHrsFxT
8eCQo4txlH3WD7iiVMvFo0Nyk3odAC2RqxxkyiouE2wJKfy+dJpZfVx4KMq2RSIy
RWftbY6Qg4ANW7pyXic2EjOxTJppZRBQOCHX21yn+rkW3QMlxhrOROw5kLLnNu1r
UjbFTrG0USg4pMzMBtieJj1t/c291ut9/1r/RwkXfUThHpJ3egQ7/iDTsCbOOccg
2BKna5pz1581XqFI9D8p4SOLOgKRrud44269d4cMjcPgsJ7JjFjVZRGjAPuh1Q6j
UAwGM/gfhcWvEw0O71KArwNckG32kpKxJCTPw+l7kTY3zQjf9CBd7QpLHc6n37yj
t4KJr0LWYTugfzvGuY0kzMRA09zwcTLlMZxzNSUEgsGQsbAu6oV3L0EJH5FSHxSB
3pHJRzyOo2cmiFw1zRQzxkFTO6qKwG/KrKsCo7uMGKbdz9jNOzss9frbCdItB3Rw
/Gsszfl/OdAxEHS46GpmrUtlD4diWz5A59yJcIrb/00ko2rPOaHzq/igNMlruXdf
Z1DmWnycG9DfYR5AK/agk1h0+yUbZu5qYgMFF+kahSz+xRUsPsqVzQbOBbSODLeH
hEt3/zbVZqgFQCF7NFP/B4AESrKsCQm0tketuZJ2LbWf1By0N09ZQAPEaeV9Db3l
cqc2QMskwTe60sXRsaQJfYJAl9LnDnv/mCHrPVKn6GGE01iydg2F9ELkymJiVEZI
TOw5F9UrHuT31bNAN+rKjYPINhRZN8e9a3MIMsImOLfKXOVjoS829reh38OeDVOb
33EgefcUapukHnueen87q/uLA3hSrCeYsjigFxVTiVIX/7tqdC7KloNV+EByx+N2
wVRHefamGWsj+yKGhYdAHw5TX0fT9D0t+oyESBGPK4w1Bwj7lskIyRJ4ZovCnMUu
I1HpglLev5zpjBTXDidmujdpRK2B3bs6u/TLqcV0tyPw/bRqtoP/e0jW0EH5OSJ+
zx/o0SwZoZufl2Q9e/DMC2MBStt3znMmWmEBxMmPXxP3CK18tTw94gxAqDuuLii3
NoidK7+XuRO6CJ1cqhOq6mNnlrZtl0Y4gAZdiWFnv/JZEcRaDPro4T+ITpjigCpF
uXRTvoUCAHqh0NfIjzhmaqWntzQu9KdNNn0iGLrkrRhgnfPd02xAeS4WsgjuC0Uq
BaAnJkTu0R6lyDqLX/AHu6ztivbHcSE+zYS4jH8ioSbEPkwyUZUUrpZOICqkf/fc
uQkPh6W9wt8XW9eqmcuh//Jug0zCcEihzXb6aSRVn0SfNbLFur9tum59nifepuBq
8z7T/jcdK0SIIt9EGrAWNZdoOId6ib7ujpRBl0Sfj6OJLvm5ZNDukBW8SAdU07MF
IPM4JGe1vdJsAfBWHrYalMcrXBYe5hX66jSjLa1NjxxISDUgOge8NZFYBePJEr4c
8lq/Q623evLbQ7j1WzBzIM47S4PRfYq9RKd+lh49hxFbJ7/5ow8WdfZvhrxEvmki
dcQg2jtEKuJHbygCRdXGTZL3Jg7btnEuhm0dr1DUyBpwgXAhD/CB6INP/MwCrHAE
D3fAckqjhoxTbOPkWW9AYNfDbG4zkL0aNrijlHAzMip0rM2+ExUgMteaMcvzwUol
A5AjXW5wXH8LYvDxBjB2x6TLOi+upv4H3mDds9ROsfAbgBovJZ/0dYFymCYtE78V
FOivPvsPAmR7dPpJpddVVZOe/lekvT3nj7Ayh/KxjOCNYII2MoUfa2PBKQGjLvWe
ohRqaQ6Nj9ifGudx5JB/vMqQQ0KqBSUcjdust97Ft5Q5e55ONMNii9qDXqhsTZcX
DvIb33BcE+M1WzgzHdC6MBiFGtl6xga2zYTbrGWvo6xVbr1rzoRvpy3yeO3ACUiP
FpGinOEePCDpstkP0H+4ozkb7leOvAu+V76Fwly6uAdqusLEyng4EaKMTzmwNhhR
znlhhgc7sir5GddSjR66nZJoJMISDBOOL4Q6TKRtq2RaEcF7IzV8avhPfZzXR2ab
owKGxj3tG69QaO0ty9UyJIcFbhd4sTwGkMn/TJCVIg/3QnlqvnZhmB3bFUAWxUZa
Q8xFw7fSXyqdYNN5//2Sg/E/aC/HLX2D0BSnd9Vdq9OFh69sd4jsVuhd7F1NYhDF
4k0SbYWwJbW1SEv11Nod8NEnjiMhYMrHn4fZGDQi0OYjIFoUthICq2Rwclg4OfTB
HhO5OF7gna3K/kGkbYJ9UNYoh06Bw6WhfRDjGpwn1A+buXdaNwKNaNkizE+94Uuo
Dg4nE7gn8HuLxSa0SfZrxQdHOWgdZUI+ABUeh9BpKnmjkngydm3WyOEygKcBwbgV
2xlxY+yyDV86GVf7rCfNRr5V49uHneoL6GWefUZ+RqVFUb0KU8FGdV07sxhTD3s9
IZ9vLgvGjHdRk15Wg2GhrrtvBte6SibJ/jKZJSlmcxfehaMpur5vYKQZe5GkrnKl
zC7RyYz6bVxKemPCLzL+ldQfg+NXftsotgNfoP40EHAKVNXlT/Tl5PuBLQ/wTxHK
Fe58cbJYs8IlqmZHJtz2pfuMIT1vHqgLkz4+2or/RhdKdR0xor0eEDuuNogSAIXB
ufi8NdpKKQ6xo31/WdM+Pc07cie/vjJLZ7NcOXflOsSniW4qkCZpAGW4uSsNw7NN
8Tlg5CMABXAxOPMgZ+/qKVbqo7O9lEcnJHbPFRjR4iXndKc6dgr7G6+g6Zan2S0C
LSEYrRE1fScuV1ED9OqnBb5q1F6TikzPKuShAvlG0Ggi5FZgEf1mB2Fxr1P8toK1
0Eo90JGRcXVMHJEHAMNkHsyngcNwSxwixMwwWAMUWb6GMTB2mEFsvRo85f8u14oj
RoXWWfN2rkZZ1i0QV6fsMLB1iPzU3zfH4PEAV4spqhImZ5jW9N3smK8DtviHyJ9/
6OVCtFLrl/ThC4fvAc1OBLtGcxuDCrMn0ZgUFH2ceZbib+Yj1NrgD+HvywvSG6is
SCbc/ey+ORWoNrd4g1zTNx5xKsMlW2sMVnmggCQiN1A/Gyl7RQi/J1Mxgtsz70CP
n/cABQ1sWgVFDqtlru6BM6T41LUvRtFD9pQCnib2CmI2eHYSzCRNkZkJPEjCQWzs
CvnSionIvKGA4ZibnmSFpxFJZWFaIDSL+vUj63SO+7sVkf6ot+YXqN2kT6J6wsiY
4qG0TZmhFpmnLLHksWSanuuOEC2qKc2xR0/5RQRLJnfK8RjWHrtkxSYrbzyatTo/
k+blHj8fWSQ0+mlVU55ZlHUAHUJxEAbWd4s/+o8jj44pbIgdP2WxeVu1iF/0/kVM
lWZ9F9Yf8jDnHlc4VF35+h+VrwCuuV4ARtaTayB21EDZAzG2TjoCKcwmF1fd973C
6aiLe6MBFC6UWR8n6bjhdUAkwoAiy7mWmtJ2d6PyL4au/mJsN4hGX8cEJ/sNy+YM
LLmGYbzlVe8gPgIO/4J9zGa9aQp98vQPcV45tWHctHVxfO3rSGdb7usCFL81mmkq
93G8MEXk8EWR/aIBoQ8jhN0Ina5ivsMcRPMbeYZjHyckq0GXfgIra5NZ6ado4GLE
apI9u7DscOREG/qmCX+wUFhsbeXhkKKdoUyuf8QkcXUcLrhIV+Bhn+Q2XLjeaqnx
Aep8rrqgyJ9oTlm8+WjT4t6HY24P4vUJLGKNDn+tWlgAr5rDENBn9S2qXW7+RqDe
VQgp9MPJdRLKA9I8bHg4Q6962E+74IFmbopVNWKxQLA+SiF5mAVcACzxDtI/H+0R
XVGpcyQKpKHGlcvJCnRzWdM9XnXpZp844xcvQMDhL+C/XJt+erkKQgukSRL6rwKv
TODwjvl21Z6p9IYLM+eJkw==
`protect END_PROTECTED
