`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
65hYn8138CyeAewgUBCT1VCqGXmvVAErIeiuE2wdH0GtbkZ3S98JO5zthEMArxkz
syxizlAXbidHcOp8C+TzubuFoWGf+qxlEO6R1SfzuaURLr5c4+VMsWdrNqcW54jy
sHTqTeJ6fn7pTIj+a0CWxqQ+3vKGVAnY1m+pOpIPOL0VKFDvz7FQD88d9rsIdWdR
38PM5wpvs2NN/dJYeqRNpS7FjRMPp+LKnwEWzvetttm7tewHHSBelVBo/cWJWtI5
xBi6ZUx79pL1ac2O6liWQ4xAT8fM/G11yE4Ha4KXtYAgTIpMuZLiWA2AmM1k6vfh
1FlYhGIJzP0zl+SCCjuLPEiTIkDoMflbEnUmOymJJBPC6SO8cIUWTgsPqU0BOKTR
mnVn/neW0uaxJMXO5FAlIZ4G9nBuVUETdYlpWidgb6UvIhhQPXFG8Vcbk+eS1+i/
wmXuCFNSjVGYqtrin3CPuO8Asc1vtl9xrZalh/fG5EDj83SWMKyn0b2hg2lR+1tI
dRfs3fDgy9GrzPM/qt+OmQ==
`protect END_PROTECTED
