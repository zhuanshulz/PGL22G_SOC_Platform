`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G6xpF3YtQafgamIe7qhTgohyxFs/sQ2mKRjFsK1PW19K/ZE36mOxC1kzpPHNHTAR
eOkpTLGqXL7pUoP8lEWM1uhlJgkCRtby0kqE3qvL5lFo8M24JGdCzu01ZcGxZ/7x
1aEXZjsSXLrAs8bj4REXjEAMvs9Tbu5OJ2xYcP7Tv+N4CoDWubssbHBEYvt0aDS6
CKgpPS2eqxVgFVQBTLgXlz6iYi8rtjsSZTQPf4eMEEHJLktImRpyMjP9f7KIi/Et
x+aGP6lGdBnmgfMaC6xLC+vKi/qSE4xfuijVkDhk6IEzZQnCj678hZva+uO8pBGX
jKhf10DfGcavamMOgI+WOpIl4DsP/NLxiM9S4ItlXEZxI+Bb9AT2kfDF2Yapm7dk
VRJ3HIFvUahQey9rJxmE+WCCM5HB0woBxTvNauxzpdz9QHNvSM9zNwP2r31oDxqC
S6vFTr3x7llHrwhJlOopQqfSbXfNmsICpxm4kykRzeT8iiMsAci3eq5pVWs7z+WP
VoiFesJ/9U5f0cbjcNRjDLIK2yaqHDs0km4xs8kGXaR547DFa1mNMwan+xqZHn6Z
Ky7bymeIdss5zyucM7GynAw2fGMTSPZMBfVKCmdcViWukl89DZuIaCzorakNxult
s8LAsNv9TQpIuQhoO8uLG6QzTxOR1Scc+BreJ7SI6OWjynorBOag44Bgg+FlvUXx
cOh6A2fft1R6GjxUFPrJDppTJDfcz8cWMmm965qUNfzGfX83p1b9yQFKHnhQMypG
`protect END_PROTECTED
