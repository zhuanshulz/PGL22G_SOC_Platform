`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pr3evovOg12YYGyVGB2FU6BWvGrfO0Gp4ZdlQmD3NRuxA/bfUnSFRgTuhF0YoKnp
cBs5FxFNxPhj97SCc4zanOWC5/DhROFSVVRchaOHjl4ttlnZwK65Wr0tp6X3PPIe
bDGDYZEiXlAzoPOBJn7Mua2c2moeYyUpGljeWihUI7mCht5M7bQUBNXkSQeO7xvW
RuEZoGp41Zu/Ug2FYRp6PWE2rioi+n64+H6RpgbQKvWYOuI+hp/vVMfEVQCDYu+X
saVIVMXA3meMpLvYlI9uz+vqc5zDEBAtIsLnT7m3ZEYcnL3pYD1QhAd07WoJeQHU
++OWWQW3xKSnGFUAr0nV+zqYxvZsk7zgsccR3KRHh9pRLMxmuHJ2OooAJcnn+mWX
A0XamnuAaJYmy69EVwGNuDes/nPnQjPBwN13iyksNwCq771Z7Z8Y+gg+MPT9DbRR
yDBy3RorGcg9x6haBn4mrUGHOr0Dp1H5EtW+3ZQgVxdSYbtOkU8fs7Rffiv5eZ5O
wkFnsW5lZJgeDa3H+b3cx1SBbrYE1G0BRgQWoHCFp6JV01ud7/BdtSixI6VMp+O7
G7rtu4+6SNaLs1DlI6OV1JjfO9sl1UYM+5WywiiUSEWv3ND0Xc+CSy8CVlfrIzsg
0xmojH2qpDzZHpJkqlPHtVH7jqcilYEEaP47iH51xhvl4MHuKKpX6qDnsbrxec5z
8nBELr7ClhxMlEee/ivTd/XI53kBf/qFBekjO1SfNuICPV2qgTUhLkMt1vGHcpKC
xZ/tpq+esCLd7V4UAWmUV0HQ9+tHq4h3n3tO82DioH9m6misecFvQAc0WC/XVjBj
ANNjkSOChgW8sj6fFN8R4WazmX9HosP4QYzq2x+jPk4SGTd5mjKnotgpum8w2yO1
Q5vkBKO5KEiIRDH8JkcrTy3wDjd4CvpULQcTZxFpuJU=
`protect END_PROTECTED
