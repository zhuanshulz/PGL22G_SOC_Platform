library verilog;
use verilog.vl_types.all;
entity V_OSERDES_E2 is
    generic(
        GRS_EN          : string  := "TRUE";
        OSERDES_MODE    : string  := "SDR4TO1";
        TSERDES_EN      : string  := "FALSE";
        UPD0_SHIFT_EN   : string  := "FALSE";
        UPD1_SHIFT_EN   : string  := "FALSE";
        INIT_SET        : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        GRS_TYPE_DQ     : string  := "RESET";
        LRS_TYPE_DQ0    : string  := "ASYNC_RESET";
        LRS_TYPE_DQ1    : string  := "ASYNC_RESET";
        LRS_TYPE_DQ2    : string  := "ASYNC_RESET";
        LRS_TYPE_DQ3    : string  := "ASYNC_RESET";
        GRS_TYPE_TQ     : string  := "RESET";
        LRS_TYPE_TQ0    : string  := "ASYNC_RESET";
        LRS_TYPE_TQ1    : string  := "ASYNC_RESET";
        LRS_TYPE_TQ2    : string  := "ASYNC_RESET";
        LRS_TYPE_TQ3    : string  := "ASYNC_RESET";
        TRI_EN          : string  := "FALSE";
        TBYTE_EN        : string  := "FALSE";
        MIPI_EN         : string  := "FALSE";
        OCASCADE_EN     : string  := "FALSE"
    );
    port(
        RST             : in     vl_logic;
        OCE             : in     vl_logic;
        TCE             : in     vl_logic;
        OCLKDIV         : in     vl_logic;
        SERCLK          : in     vl_logic;
        OCLK            : in     vl_logic;
        MIPI_CTRL       : in     vl_logic;
        UPD0_SHIFT      : in     vl_logic;
        UPD1_SHIFT      : in     vl_logic;
        OSHIFTIN0       : in     vl_logic;
        OSHIFTIN1       : in     vl_logic;
        DI              : in     vl_logic_vector(7 downto 0);
        TI              : in     vl_logic_vector(1 downto 0);
        TBYTE_IN        : in     vl_logic;
        OSHIFTOUT0      : out    vl_logic;
        OSHIFTOUT1      : out    vl_logic;
        TQ              : out    vl_logic;
        DO              : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of OSERDES_MODE : constant is 1;
    attribute mti_svvh_generic_type of TSERDES_EN : constant is 1;
    attribute mti_svvh_generic_type of UPD0_SHIFT_EN : constant is 1;
    attribute mti_svvh_generic_type of UPD1_SHIFT_EN : constant is 1;
    attribute mti_svvh_generic_type of INIT_SET : constant is 2;
    attribute mti_svvh_generic_type of GRS_TYPE_DQ : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_DQ0 : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_DQ1 : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_DQ2 : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_DQ3 : constant is 1;
    attribute mti_svvh_generic_type of GRS_TYPE_TQ : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_TQ0 : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_TQ1 : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_TQ2 : constant is 1;
    attribute mti_svvh_generic_type of LRS_TYPE_TQ3 : constant is 1;
    attribute mti_svvh_generic_type of TRI_EN : constant is 1;
    attribute mti_svvh_generic_type of TBYTE_EN : constant is 1;
    attribute mti_svvh_generic_type of MIPI_EN : constant is 1;
    attribute mti_svvh_generic_type of OCASCADE_EN : constant is 1;
end V_OSERDES_E2;
