`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
juL8QAUU+1hfAex+MY56i4L/5TFyoH+HYHV6syGKD6Lo9lsxvp+v22Hgdh7R+/Zh
gXufaM6DFRnrzZUrWFvtaLhHkS9NJAl2tKy0xHEbyPlzGgklDrpogDt7+IxagWGA
ZAExAd+xvAuliJWemWYzZvYSPRllVUeCJl32o0xcODESWCKBN+bzto3b9yhxNoUf
nT2C4fAiNSsYRo1WnTE6CY7VKe4FDp7FnPs6Hiw6gBWDUgBCZ7i4QQ3jeoWes1US
TJZmF8ZxVE9Iqlc1InqVK9Pt/ltAbeq6zYVg7x1kKc92cFp4dKE1MymYslC2R6wD
b5H2VAswpm3ZpSIDA0YzIyY7v9YXSrmCRufcaa76Mvk4xDVidfwx0bZ8wx6LrIy7
woRigmWYfWhhfnknXNHW34Qpzm92f5mNltxRLYsCZPGKFaWN+nZiKhbx8GoWZfa8
PiKTCFVVnb0efXBKD6OiU6Mf6H6xOe1p1n4SqLng4MrhgG6x6Xh6MENM4FSs9KD4
2N+PiGM2/bkLZSSJHu4ywvRGvHxC2WgzmsAYp7PLNb7WWESYWHlsBTR1HVmSE6rg
dHfVbmgKJVmXFSETFeEq17cLQjQRBgjrSq6GScT+KhXLPRDajIeEnPSqXb6m5zJg
3AfRTdEtvDKe84iqIMMC0rkjWI9pdz4cLpzer+MjA99AQl8IIMBku2Xy+ZGLtqEK
OHkPPhc2QI9j6D1VtWr+XdN+jd+t7iXIXzjHl4SsI++XRAzyBSAZ3Zh2pnd6Reos
fS7uoRslSGNaDO2TbLd5JrT9AB/PXWTdLwUEAIj+mzlrCceo/vgLmrVSxgobkp7K
CBru5esEtljUNNluo9SttrRfi/1pnYCAr6G+zyCcREh6lM5rjarjudEM4hO81Kdt
uTxZAsSkWNIH2v2IDVKPp6f7ipMeNTUZkMErO/SRtBHNNujZkZaoAdzgt0TVbSec
F4goYEIdrtKGJaWGul2hnaYQCTVRr+znRqQNgmnuK4zmAHmvsKQtBK14BiKNOum9
NpQRlxaAYwHS4Wp69Mmb5npvMacg76nGMjprIraCI0jmcoPu0htt2+5RTg9o2L0i
O+XpTTSnzM+ojfuto8rYaj6k49JGIoprm3OdO0DqHtyX1HmC8MWz0HfyPOJ1oT+k
2Ru/4ANsmYFRXmNxdv8z5ldq2wfsTGIVC4yHBw03nQHuWOgGlUXTOD0BNNFkq3Q2
7+WBvVsax+YyGX5dH0z0piWlVXF4+89YGggvG/dcCvh55ttwRMHbeCp6yfAXsYPj
iJ7EHJvOIoyuCLkcM0m8SWCdwtpVr0vUU5e/5hVdzzdDB+N8RU0tdsTBq6yn/YhV
3yY1oCkAHEjoxxwFyNvTIipvoCnyjq4COgiBjQEC08+IohzKRjXnBJ+yVljcrUeI
FW3ccZGh1sPKZ8IS/2ycirstwr0FNCZ7O6vQh9amNrgZT3Z5B4SqslmmqWVoJhqm
LzQ4y6Onw5jDFob+hGY4Ox69FAfhGcfqmC/TcCVXxrFb+TcITCIsMcCdEPRXKPGZ
8vsMxCRHngou5BUnoFzRliO5SevpdvNuYwkPgodXkwaZLRpU9/vsTnLjZ12/3+rx
WBwp67EFSfbHyLF8iKnQKfyDo5GMabwXCW8V4Bu1oe9oFXa2c7eTJDZcKjrkDTZR
LNY9DY67gBdYxLKhxNz9SyaQNFQyyTsG2M6h10BBrT58jYzJvs7YLDovbwK1QIge
5tjHZjfoeciR4Ox+36d4FQAq91A9Vp494J93GhTlX6sIc9AgirzMKrdTDCbtWd+a
PDg+ooE6D2GZ4/STlWoR1r/fJl9ErHVgUgQxaWU0Sz/UyzZvei515UAzlPJlniUe
egDly8oqTyXWdAKKu3H53t4IwFQnU9AMn1ckLhrBbQNctnNQ6R1BMHLGvjEi9NWP
ZEBgQ5exeqiZO7DaYgpxVeqse9FRdl0kikAx4F3bKtvWV3pnRGDADU6hJZtzuf/D
va8q0KY8BQF8qs/xX6Mggq2YLqt2rkUfGpiMmk524kszu/13t2TOVoJYRGfUvqWw
x8ZJ9jzgTLVLqjTKmw5BZSV9y0907VZshN3ApeLZzJXvOfbMskf+65jsvtuiwS8P
fAAaDmKNOxaqaen2tf3IDJUyCH4ewiG7b9Ma4LSJMKQl1EDFpxykh69gd6BifqBZ
zaIOLp+Ptf7uCO4UX2ZQGFNBMHYdks+JAXEkdfS4osPFRxylZAnrb48M6bSezxI0
sUgqtAb7MxBZOou/CjpPg08MCwHxgTuPfc6okpA7FO7MMKbmguvlKmJ+XR2rKwaE
tfCSm9f4CUeEzyoUmLWqDhVAsA1suHvlOA+a532wJzLzmNBCEBvy2bD9FzGXFX2D
4Xu1uGthPKNiSW4+zLTv5Lf7Xk2hyRn18dgccqDP9YO72OsUmqX5qtJWI8hNs+F+
7pzaJXkA2tTI8A+Q9whvm+Au9lsPuInr3i1gbxGVNOUOhJtHPK7N256kEuwzxOM0
Npdu6/fAhkpk2CjoxstoKg3s6kPFem0Y/Rng8+pm81VZeCTrXGdUyXrB45v7vUbJ
hRIao8SPtRBZNwuTiCyf6dWqHVBXKQNjzrSt1TsvcDBZHgwC7Dk/1bXSEYaJmXzC
7UNpa/6phA7kWVyvCyHaIcKpdO05JxA9l6Qv4JIB/HERqJ9nxCXDvzW7orrB7ken
0Kb5Fo2cBLSjzwnT6ry411fkptcngop29LFCtONyEyk3hAdsboz0eQx/bme8rfNV
c/o4/LPZ93Pieguq/FLkkNGeDC4d/ggzfM0F55IHb7GAU58JvkQHmYldtt4xcDC9
GWE9rggZ4ipaScFTQ4j2f8PtMZ8buGGaLbR89kWmCpQ1sMfXDpw1kWGfarMwuZax
KwAoFVVzqg3aYSN9nKLYeWLDHbuk+dQypo2xCE6t3t+VdPw7IiP0GwnIWdw8IvVe
kWemG0XoHNf+5MONYvjohYEA/pELgVydbSvHk4O/sIClTFogWsCPsXGflWsgoAez
Bqb5a8qrgQDCESM3sRxbb5PADxIT9uDAcRtYcEsWTdO94dtmo2pzpg0MEVnt7V5k
98r+iKpd7P4NsVFABPIIQl3ZKdVE/V7uzwGl/BfVzNdiJWzW6v4iidi1WwhRE1d/
+RLOigDXDgj+bkY71gF0eI5QkNL4L3RXFtMaEVQPBc1CxX86CZ8dKGQpiyFeuP1H
L/ItQWpeohm8PmY20hkFOiPSN6tV017As6WbBugFpNq6vp5fqFV0M9xXyzy67zEb
LCsnwVXJ4IdZsZmKhY8Wu8sC/RQqGhp8UL0A07RQ7CzNJOeY5IER5+bIgrBBDZrf
1BUpYzgl3GnAQG5swNTRQ3SuVpceCKduKigK5q6X8KbWsbQSV0mwEEls50085Xon
8GU3QncvPRytx/syf9xSHJn7ntvly+1qrxm7Nal2DH2ephUCgc/cfaXrW8toH2i4
y0mvs/CCOMHQBeb+9L/2e2xoQd1CqOgjX+yVN/hpNNgoK17l7fPs4twIL7BFXxtR
QgcbDdTGieyLsRLInS0s3Lash7x6bSnFhwoDiF933tCVsikt1BadanDSNOtllpNU
CNzkjVDog3XwIJ6w3JMyFROhQlur8dldJihGhJLfdcM+uYFh3gxtITS5/CAvD1RP
Xxwm0co4vhstJmrrbIptWginANLrz9p0zvz+NydgmF9UT0oNHAFZfzEHYAxu3mJG
MXgKbbzWOs+eJLVFw4tR8xOxyPOVmCsvmf60jvFGuxDgkMEGuYiMRitT+MBNNyPu
Gy5WKTX/fkyfedIlzPdnYNdY4t5HTLxe8fYiyDq8qH0=
`protect END_PROTECTED
