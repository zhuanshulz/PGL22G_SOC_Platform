`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMykxoKjXx358sqUPm/76B4HA35cQ8VFo2HI5KpccZVmhp1XR0TuPfGbAhQZKHce
kscqNQ/OPq699pnAVrlf6cPnZzfc3y3k9n1baN/DfRlSnTHFCw4LpYyf/U/3GG4H
wuAwADrRzQHRBesMR8XVsrXjlz0Dds5p62fichoXurMu05R8H+4hrTYVmuiJQjzx
MC9+NThgGlVaz/hZx61vQu1VOTYQH2W2GBdrZ3f0MXM53c/T0iROQjgNjqnrLGqL
NAmI0Ipv6hn61Z3zrjzHxSUVmjrAJfhaNQVsrGWRzBVr+ER8LCpyCAaDN+7GggiG
UsEAZrGFyFtGPOtepahq9TapPKpnW0N65qWeQBzPuhLrQ7PcNomGDiM1rq9Pcio8
PW8HpkNzpKy9yjLHOAncWFSsmKy/629RueTlhveiqt33i6oaho6J/6mdhUyGQM8X
fmO9Zg3EdOQODTbrDY94west6Fu2Es4QtM9pJnCLhScwoUPRE0uuyt/YVQuWZoAe
q6eq8NbDfp+zSyOsuGi/dX7fFnGjRoPxuJRCB5cj+AF7nCx6RpRC72Qj+zzanAKA
JG/Abo5kK3HI+QZxJ0fovA==
`protect END_PROTECTED
