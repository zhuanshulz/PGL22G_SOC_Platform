`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdOADc+nISNFsgJodE8FT2oyYvdUdiwxqUmpMnD4GEs/lbHQ4g1JhFlE5WAw5fQ0
l1EWyFX/j+MPvUIpQOK+QFpQcNxeRHNh2XuNKQgAmLyKU2aH23KHTYdR6w+/ecDO
PH5um00CgTQT8f3xjUKWL7yQhdD73Ckq4kiUrlahOO6E22B/VHOZwhMEcBFT4Nmp
IW02onA5ro/w3JjeKERfcYUDa+Er7ccoG+VVD6wLCpUAaVvpmLDfdwGxMaS/xtFY
jYdMXPdcYz8zzjwUdKbEeKC4DZgFOb2WAks6xGUVm7o73JS63TphL2yMlNb4/42D
Z57D/omCZnw1p1ZVxFpamBQluUhfy6kS1Gp52M3cJmRCGMnNDKnz+2dXq3XVDFcg
sTaTa2ZHQYVGqKdt2UP0BhT7GIrrxSuxVDRjUoR+sEC9W7NFhAkiAeMzktUoBNiP
DPM8bDad6DFo0T9EG2LDNN5Dm4QXogCVzt8gc9OTTnHAv1zfkpY9Q1flfyaPmbep
e8y293VjxbkZ+okMbXLtEh/zfBbf5r+N1u24SmOxCp1GRcqoKMQxwJm4XHfLcB7R
bB35KE4iZkM5pnrVt1uoamtuW0zn/XhoUUZHXAJFblrjJQqyaWlM/ri1npA1ZixW
mEMhR2m20f7G35C3jXvpqXYtimrSDDqva7fh4M8bXNwGcVX8L1gDxAqfnuLbktUz
EftwP9lcfFlvAEPqLYYjZ0deOgwjMjwFHZExIgREBU7m8aErhVvww1nEiwMokfGq
Ps21jH0JNtlwPzsj3/JwiK8jD1bLhcAe5x2Woxj0RJv2CvPW0imFOSH7ym8w+Ozs
CAPZoGOK0mXOqesfYb/gYUKwFVhyhsODTOgzp6Lg68OEvMHe7N0kMMYEOmbKscFh
q7v4P9s/WU7NTQRo3TWHVrbnxHSmM74cJkrkmeQNBf+auKtBDGGkAFGx35M6u+Gq
fo2WKtuV6sJZ3cE4MsfXCV4mmYRjtl1LDUKjIhn3d6OaifyO3vc883lXSaXgmeYk
6lVwSq6cs6EPt+/hASMfcjnijacHrva91ad7JXxv92hZxcN/qDDoVsxrMYIXZCQR
zau5KvsgiACqIzyZrgRIY++ZcfUChpQQoQtq+U1eAYR8dZ5G757iE1EtoQgGhrhN
JYt4I+mKFRrtJ8ckmQFyO359d/ebBGlWIbhu6DLQS1KmWX3GSM9lVlMWOqUjX+Ix
tPIlfSTXpCf5uinDqz/CgK1wVc3VzmWZoATtHiDLQ9kSZVLNTDNubn3P/g2tmVcp
7Lkx9DYbSjY1Wocc/kR4F38VAfNupfPaPutSpMmLyQfkPW4Y5+KajuXjENpNQ7ws
qsKm9tC9fl91LvuHoL1v5s7SQymZ1N4N8M5G/6gnnIXpQPtmd3oKhBL+i7epQYX+
c/oFOTi/eSZwUr5HwbNzXoXrUuwGr3ydCc4Byleo4kDniqiiksT3xwU4GiE79KMU
VeiSpTo4FMY/ku9KzwmjOgdQZC5/cnzzl02uNB7OBqNhJ9rsPraJD6DXh10cPbUx
QsEjN6KgRLcofO8qKI4np5klzADGbzjlwKdfiFxVKsHdP2D4fxz6bhjh/0vI6IYT
9kHGMqyPfI5N3haeob6J9Dp5x1rrCJ9TdTH4SZkz3q2RI2ShXeMDqYW5RKZkObgw
2pk/cw1EzhCCDCFBIHhb923dgDC3PpX5MBH+ZTC+9PqL22jhFk+lqs41GmoPAVDQ
tLGXjMIF9FRM6FQbl8a22ROYz4ibWHMG6Gl9aSPh/SxfkriqTIac1qPPItlbzON9
hJ7bGpeNGPLs8XE5LrmPl/Ml7/ckEygPS8wnn+97K1ziECsKEJ48k3A6q4xj8pe7
ojtL6WUQeQN7LV1BrvkxFx6g0406iuVAGD5Ao9D7Xhlv2BuTmRQhVdzWBvn8g7/j
3tjwP/5OiT49i+gBUenxTX02As1Z/2raWLpK2yrWMOTUdBoyXYX9Fq5B2pha0nd0
bj3kgKZ73AzIefU6ZaB8j7fJiRr0JQdYlq1O1KkS0n+dpyyksAHcqTZVAsdbNpea
Pk1+JzN7ezSnUnL1OZS54A==
`protect END_PROTECTED
