`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZEeo0dJ9wFf4eKoAGTYXjQDP8f94zB3llAn3zBk0pkipKpehYsWd920Rm4luYqh
5rQTtbiu9cn/bIksWFmN+2Nho/cXw7APrqGvfigfvJ4O/Nwq8gLgbcadegXbLJef
D4BGyr3OzCsOu31Kz4OwpJ9Pr8v+YuP2CHHCrk8LA4bbTECsBbXnVidXU30TVG72
+2wq+NPpeEvdgw29Bxp5ShOS/djy7L2BIMfn2aHEq9zbiBoVwd5fRzUikeMmDloe
Ltbv/raupKmHGnywulX2wJHrf0aUjCGrdTJkW+tEP7z1pabo1MzMRw1t4MoFbfbG
8+3BDnpiyOcI9FcGLXbsdG5Mld/kaPrITffxvn2HgXoCpPVXgkw6/s77YIE94M2H
TdQ2Y1360YaaGv+0lyVtKLn8vnHpDqX9pbqFRrERuMDm3Qzpwp1jvpN+nb+opllW
mplYz+jueOhJ6Vs89/odIQvVouA22C9fQQT7/Fnz2fSQ6s9ECJi1JgzadQZqKWav
9ucvQZzdI13ro64G7tW0lr1o+GPT6MIT5QslJsr6c4GGU8KEddsBQVZYo3Z9JQ5B
IVFTcQB5JmXrNdsXo6hnZbU7RHiHw9JCAoCuN4uyHmWHGCKRSd1F876pgxt0vHXB
2NO1t6MKugpT1GUAIlEq2LM8uslXvt4/Gg7mIy+X2nKxREcC7mZJb498OlNsGU66
c+0kes4lXR2OdpjZg0n2gzs1CboNymo29Tbh+MRoKHCi9Ct1DpQEZRDVAF+yeqhk
arWyWB6gXazRdviSknxI1LGHBi1AAN057yzERvb5TsCwm0vI+mWdhF8gl0T2WDu6
73HAxbSLHg/wQRkStTZ61DY8NGUEnMgIitFi0ooo/f0UOth0HjENxW/vrZEWF1Wa
10Wntp5Q+Sg3akwDihlm6C2iASSesNW+8xMoC9cSunGQkmTyqwPqdJEbpOp54oNX
7M2d7BarNgu5YRxxRPx8+bQn0WXRznHuROPvu+a5hb121V36snDoUwd9ynQbr0Gl
dPhfwMLkTE2vtqw81Bu6WZC/jFTUkSNz3jyOKSPaF9it95T2efDxYmBjNZaM13tM
sP306BUt4LcCVgTIXTLkRbIv7RtLPrNoMTGT152pm13fME6ZAHtluqTbMpN7K+7r
jFPFXWqOz27vR58FflmiAVISTPvsNqxpqYjmzMsadxSmzpP7X7P9EhLiIePmthip
MKzTEwjgCHLJ1BKm0/NM079mJEYkBORe9n0TskD8TA4=
`protect END_PROTECTED
