`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EeV1cFHI5+DD1abmGdTjcXLYXJJsHl4RUp2EFqIEtdY9RUYhFbL9gFhlObG9IkTD
sw9HSC9iRrL3cXl/wO4nnewFJRELwqyN1OWWTlZIUnFWX0I+Pf5LvT6RtKpukU0V
49Yq/y68RrVqbzv3FZX3aCIrLJSQm2Bqg69mMTm6KKpBk41QJR+BOdxfFW6Lg8fj
27C7g1fPU9VaNjusCgRHL4bXSJvl4W0OXXF8nVPNLqI9Yi/vMpQcJ3Qcn5W1vAJc
BEC8IqrEIQubunhCQg/qBGnmjo8PNlFTSMIjXbS8c/BkBF/BUEERkTkqGuLBQwyO
vpyqv4+WFV2Qu0+2COC61asbvrb/L1JuXPgw0ICe3HL5UlNUNB5wL2QAqUZmLKfn
E4Eu9b8v/mdP4nP5lzTfMrJbsfrnNVsesdN20bzEwqt+fOysivRDOyGZlIHPTK3H
UIC9SgB9NwUzBMJTW4AfJuSdtvaWBlfFf+R0+dqx2pKcazrqt2ICBAmuGCbDuqYM
cw3HRR0xRfQqAM0UxpJaqHjoo0NIuUuVjhHxLOu5JS1f7Tp1dfH5g/qxUA1qGJYa
bSoTs9/qnaUXnwHRdud9eSGVkvz5Te2H6lgZXRDGqoNYXpaIsTK8zEpeDC9wj+qL
9pwoTQeApWvY1Vs3u55iAP9TjL58VltY8be1N2wUmwWPbgkIpNEzj8lGU6b5tUXY
VArCJf9Wve4T6u3RGm0GWvvrZDh0dczzkliHFsY9YgujBMPQhMjG3PL2GtOfPASP
ref397MWcdsxdW04pl1FTTlnO618Jgg6XwLUT9p5jybRKCnEKeDbq0iPkVVg45Tq
Bxg2h4pnqDMI7Z7y8DnfLLsCfVRNzqF+XjKheoRg0idfAe6Uakv0qEcAPPHoxumq
RjgWmF46XCL3N2l/ZGawC02OCVGzVF2NtFMhRCUfiTEAlxamiHg48Hnyk87Q5K8s
MWrG0L7RKce7B4bGNXLLZoJ3mHgptsps/j8J+IqPdR+mHMbNbPElKYGelxfuAvSA
iy2zQo49CR2mNeuuxxtYj2lnQVMgAQsqRW7VnGWFotvGye2Za+zdWE//tSAjJMOo
5bclqiXOy3ZWT/TUh7LtrutFkV2I7odLpCPwZtbum1df8N8ucDSjh/hoWOi9FNj0
BblePe+JdHnSGYmsYTHiMQ==
`protect END_PROTECTED
