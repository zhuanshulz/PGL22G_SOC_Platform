`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iP3FiI6Kpa6bShnS3LfYYDIxsZi+6QRqfa7fTwP+ZZPgZLlYBXOpwSzvCehddZKM
o3ei0XhiKMcYvpjdDOmmYYJJm2nqOCoaJzB+SuJ46xwOuiXWODRkB9TRj8hMNgvm
5dLRAA70yyO7uD5SCV7Y16uWYP9T1h/MuBH1DE4c84QExN4woGB80Ta2FmwLaoeL
0Id3hRIgyBhIa1T31ZP6eqQbzQN3rCQhL/pbL+eLQAJY9LhLWetcJVmZf05wQmO1
r3EARtav7qz58CIBOQWCy2wNaDO5ONK2dPDqfxP78lAbImOTSm3vEe3mgZUxnCOY
ft38oyksyNYWbIIPMqDq31BkcEwlstPVYPWhlE8IbiHfyAeMvUrLVi9fG3ZU+6tH
MQ+UdOHjs2T+sNBe2x3IoRTUUTLNQeJOA0+w6Hn2/G0sVKgaf5FhEdOecCusqj+K
ODk6qatHVIpyaFKEy5tyNiiEo9l1FHf/6vMvfwfiIHyoyl7cKLSWfFedR3uwqawe
0Pcp9JXMSv9Qwr0KiffyqUafjY9FIWbiI2xvLv5KdegLVHUYPDUNbzC5NyRJu1UL
xUNawplOqRXiHn8b5CA3YnoVMDQXEQCd/XncWfp1Oz+AhT/jRMoqG/wdnbcFyVlw
t2C17Wm2Z3R40hglEV6UGV8UeOQKV8b1c9Dfs3H/nV0vbC7Vxnne692ZIXF9g+tq
cHunO+rygzYUTgS0kfD77BetLeojqstZUs4/cdtjK5JkSrCuXsB+JnkE0QeEGfuF
Bc4zC/cPDmYim7rQUSMEN6a6bKUmHE4BvCyWTVsA+kyAqxhGnAy/7NA2r0kihahU
mSkY8LV4k9tm/yXRUzrdvP27uvmJfXhaAvo02CJ9mg3/2ZXfKJ3bQLbmsN7lB+Jv
ls68VwOHGWAMS3lK7twAT+SEwhkIe3F+zRaIhf9IAta9KSy/WbzcxxgicrzAvzPP
e7fgyAkVxgB0Af2gJVLyl2Kxj0ACPYfW80m227v1Huplcz/jPscnE07D6B8JVh80
tLBWq0c8/53G8SqJIABmw63miDFDg0vLmDlhYQJKsFGLo/TMUV5+gn9RyHFd5WME
hqq2wKyNhmdiFw25Ef9YGwPfc3CgITI+fe7k+cg4yQyJ2b23ttcu3EdHT/VhIJlX
JQh4OA/lyRRh5us4bxJfy5LEQukFmg4HeFnbDeW0HSF0N4FkmK8fd8yJLAfORzco
sRlDvG3PM1j46hOp12G21g==
`protect END_PROTECTED
