`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rlf//aVfmS1NufTr/BcG3CKlH5Qn7u8NpixNS1k5ur7l07FSANyy5VFu+5+o4DzT
FzURHEfT08ZKmlcQ9n3tGQ0OSZn635KVB5Nhi/e28dZSCMULbWlzpTWubF1aKEtZ
xuvylngVCeG86vXFuckxWoHa2ttbrtn42f8DBDoxG4gcZEe8ruHBliw910N9fRnF
HxfhzMmoDECQxhveZrD+ggrOv+jujEMFfNsI/w/g+cJY+PP5VXO+GfFAorRCu/Fn
iHWmgoxGXnqLJ34Cnz0DI3cUvjt+fc5mkZDpx1QcKqZmfuwEfF0b6XlWHrzb/Xnn
pS6ri+MNNsy+DRWturJLsBB996Xnwb/BkcKB9zNI2a4EWF05BGZ0yfdl1wHxHG2g
s5GntonYopuzbGBl0ussISJbKC2cOAOECfcZK6fe4A5XdMbrEq43ByoRd7AOEXqg
kJRXe+QlJglK09g2mcjPQlqR45E4p86xoWbGjaUcZJaEdHL62yBIsQ27DZN0XMrQ
OYuoN1WipkEnTPHiiOqlIkae6BBIEhpKzJe3+92qo7Z+ns3BOc8hOB0QAq4WLAsu
HktwIRxebXUM/++5h2e84NP0CzVqXuw80cwiMqYlC+KpQSU+/4asSmx13JEpASN5
vhql5/TdpfUp50Y8/ieW6TwNS2Btt0SegvpKikhrGCdH9QZkyR8cmf8nasEhIcoS
`protect END_PROTECTED
