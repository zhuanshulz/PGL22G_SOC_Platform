`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m5kz6sqdRYD5C07YZ1+A+bTmk3Ich9VWMaluyawLu9SzdWMPuG+DyHGbdDEw9FoO
lsxjdGq65egbjTO2V6mdeh8UzMliDM6IoOqmipltCw8O1/1Ga9jC3xT8jyutE20m
3lr1Jo29/qTnfqEzAt8lDEcRX2XAr1E3/nrIKFdEwmWKpaGeATcIWpCfLfI6oQ3R
NE/jixQGr2QepQWBNkBI2Pt1KRiUcsoUSkEF36YRozLrv0x4dEcAiTTzXBZKQf4r
xbcxxlRoT+3xrktt69kDQrAA15AYSfqJtZUdm+Qc66wF84thhBN+8xKv3Pr24HLY
oru/BH3c06Qpq3ro8hrA8NSysTxUtwFN5E2Vt6pVLOWTrcFP4XxuCu7T/U1Nfdu7
3zbNVq2UPor/S0IEUFssZrqmfK+NqzT7/TDyA5bJ9B948TihptthJM/WFtSO5XEc
jc9TEuWrjRfyktfyyyNVHKI/JazoS+qKv/ceM9JAn4epnU3vq8G25ShYWi+mLK/F
SsZr3raZ+tOy/aFxbkgPSmaFkYtp4IO21PheVPFlMmHu8tHdzCyvenWpusZfq1kc
LCtXbJwlZoRmdJGViM6TxRs1yzxQI9BHmn3eqXJxR/1qLNhqjUpwYzho1X1L0EE4
lKe7o6J8oI3witeCsYxrlQ7tgB0uzLbG/fX9WpHWfPRXUCKtcpoI0NiL98ipVsNL
EbxhIOkWdv0jXD2+rQBc/LDyrtIPzJ7Vs4WjVkk0QturVUovhfJ17wjmWlJeSJcW
B3RXJu2xdqhsBJTayPXQ8SJgSG+x9oYDG8HPi9Nf7hWK77UF8Nx6Jp26hgWNGoGs
AcQNQPlyUvivbMLwCBFHxjfTxKKDZhPaD8O75HGA7rFUpwsYqdt1AcKcYqDOMLwV
QrOBSABm8qcSudqx9GcA5I3ioOk3UHgf+fnyFlkI7sf0DturQwfQukIlbeRc8/3d
+Z+NrkGwwI7AXlXTJRteWcWilmPJUD2oK6/5+jzP72PKdVgv4z+EWYiezPgu2zIV
PQhbm4kBvccFpEImD6NJ0Sck4uWrC9dE46jTYXJzFnYdUn5dZACgOEeW7S9Nft1P
vD2rrV8gNRiCEd96APomhvYGUtIJ52EV9DJmdDk4Y+XMh72Ss0D205bjWqilF9B3
iXDrlzIiZOPMudQ+r7NtUN35JPbo11B6I86eURg8HHN9RrbKGbKL5afSpstdtJTh
t9bZhN3UEQ6o5IxDfd2R/ICQ5gSliSBViBsNMfxLCDPXulJ2XxDGEL5qhyhR/tyX
agCfADgXlPr0eK1McDwds7raaTF7U3iaG5N/NCO3pKwGjb7lelSKcUub5LKbviAG
8Q+ifUs6eRRjuc0crxIj8K4iwSQpDHqM6n51yAi5AwUM6Rs1XZs0g78A8OZ4IquG
ptGVS170g3u4H2HDEmZOxCdA8LbcmfYhwsxPFBjqHTnXHDI76SpUazTaENpQXxgh
vqyaPBEBTfwzeUbXrrdiIYdHVPMtLL/7UIHrF9xQ1hsCVc1VzmSZvqO4UvASQus1
kuLwf/tOE9RuWiQ63EtUaNoXAoeHkRl8Jdv5f+CMs/N9GdfL3PcCbrf2G4XWc05x
JzjcBvCODlIMtkokfjTVsBqPRcqjMuzJJlJAQOPW+Q1na0NsSJBE6+oDmCaJT//s
2hPACs0+FRecWtrf920ShB2mxpE4hhq5E1t3Ci3tHJfZcsPeUUQtthbPEhFGtsQz
/dgzmXUL0g97N/63IfPlzFJFsL7PWwvTDRAomz/TcemPN5kfvnQgT0JCsBMzRqaK
DxnzEcoFwlpoE+ILNabzD+XVjSY3a8CYolttbOZ6yh0nEkqdOs/V1Z5dmuqJN3y3
l/gVXpAG1zM1Ic2vJ80NjdBR6vze7S3EUvIYw0u7lyZ5MLvB4kMyQF2FgyD2OCxJ
tufvq1+P+9VdVd5l1c5fptLAzKFk22wtruHLyvut63FI3VhhSajJX4ap3YkeIsDR
431GOs7YlDwE0XTKKuv1xBfu/wu8HSQvkYS2VwLii/Nz8YA5IfFJcold43vI8F86
MS57p+873V8whG5g+3ue2B243LLjdkCQi8y8pIXQo+1wj3q9SiFZiLr43GRb9c6F
RrWUcvTlEw68MjBKjJSzSGjsRwDLbrvhY8NtrJ6kI6y/dRnDBj9kd2DeQhTkJ8/F
IMCPYyY03F0rkrV0gcSNQa3C9f7wtBZ+DcWQkB+PVL434OXvP06NGn//C1PxSHRX
bLf5IXRcMLHwTsunFVLM43l7AKieHrqoXIEjyUidw+gmVZRfUgk3nxmNE+ykZ5au
5uaoB6Ug0LM0mopBEv2cJo246/Xmw3dpbJJLix1ZiNAfI9aXOWOVaMifsYIJQBP/
NN/uI+jrD0y9pJOYpUOMRtO44mst29Zvoap9do1wBZxz1McG89qSFxDTX5gUgORr
0DBtBRpWWEwEHLFelpFEyRslwCyfA9ahkpM4F/4XJlDZf53rFL3tJy//D7DOqV4I
55ynDGatRIBODBXyxnjzPX4RkSq/5TeSYrsLIxqHjBS0wcPWSE6y+meYpXOOUYFJ
+oWsEZGw7AywEGV4AWjy+Xv6G51aZzhgO8vSwZ5QlwwJjx9wY0h6vhE1njJ/dHar
GsW1051ZsyJLzebZOOa/qnwnJG74SNmTMrDA2CH6o+IldHI9ZI7qlPMHGVJbH6bO
pwQ7EaP0tWY93xWkH3Lt81IKBc4J+6bpnnCOjzbvVbmXbYQfiMAksv3Rd6q4zbmB
fK3QuK74x1j+fonY4XyutO38qn5BFkKcpcXceyHKWnEExMaMLFtEY7z0Jd7ODzzz
dScR22injUZULba6D8DdT4kzPi0fb7Dm9HZHuVQ77yPfuH1LMPN5gC4LQhla4HQ9
a6kEEAvDa13WNwFxk1m+sidduoct74gKANzYhM8C6KMGfuVYrhOCT4pW4j2U+5JH
uchlpDt3Y9Ws6hIQBzid444dvuBKIJfvtyosXEu2QPL+GYwzC9jCy3PlcqzLpo39
UbaQFkDcw4mn2LWN69nwYEYQ77w/oY8sQupWq9l9Ry15ISUmvvYIrPqGA9oXGzqT
3Drp2JXYOujzMmHHQz+4UyjfynxZpxdZZLpQ58p4Jr7AFdNlCJjjso0gU0YCLlg4
itUoMV1K9TP0AmAT0qJX24HBHYWNe3HqoD6jqnBg4Rq1YP8Tw+xYsP29kxg+1wAB
Ju6b2+l2a1DbTk9DqLJMd072AW9TjrWPSbApjoZooU8KNy9r2w/I1mmgdbcwTIcr
XQ6P2LhNPaIBH7uOMvcXiggXLY6mBiAJcG2aUTdfVs3CiuIGuE2+b2BB2NTTscHS
cYO/dUUq25R9OmQsUb2yFhFyIForg4T+NCBHJyWt06bumRTz1jmBj5/R3BV6Cfyf
q7QtK7tRlUoqlrvKwDyNftCtLKGB8uKSUNHQRygcVE/agQPJHfdqpfYtdZAtyUjl
en2bTaw1h8FVcrsN5WZVoTRx6hK9Kh8S6ta6Fjt1MGa6XLoCbMOjxGSWcflOf0MO
ZG9rbUa0kj7BCllUCVynlYWvMfFReH9TPWFT6rWMndNyTEq/8ZcihVwTw+SVg6TP
7mYVfHFr9iJaYCMSmYx2BXbMX2XFvv2uwyX1yDWPJQaruj0Qpc51f3tdbMh3u9R0
+3xF1/5CsddduQcpCpUHjP0wQZiUtZN4JI4C/kY29eYpUVSVYHvIKQDTblSHf2ng
SCriHF8JO9KeRY7bxA7MWVzSsqhahoj/yKBQ/tGa3s/zl0vdbCvcEYFsYUJCq4XC
Od4XrNH4glhkOT70sq8uPFMuMBxPEHtJjhxhggx+77IJQAq5CdncFt+FZ6jeu45E
UnxGVY2PuqVVRVa9va3qZjlAAbR3ZyfahBZw7kaipT8C+CBBoe1Iclzr2ogNi9Fu
ziJ2sblCAOL/Pow7d42rzYXIzdJj4MYg0aANy8aUGJD/0CRZ0sSndLTkvuj8JLd6
3JRNeNht7kWsWYgruHrQdgaweLnP06Cz33ei3sWxQoaT/LRvGZPgTDBoLd1sNURG
LcJmmTAlOJ616JPAYgptWqiKTHEWjnrxYD1pHPx8i21ilBA73B0Ol/uifodFbW+n
dCEN6okoHDWH6rN/xAiqgO3+4i9LQL6ZRAosyns/MVpFQlwsHZIMonSTEAbEvhH5
TwQvPYgtay6p8WMnleMZB/lpK/gJd+6l6SvkHfdb1tzZY3oTx+jdaAHROA5UsTTr
6idLMxTJF6ALASCbsMAD/FvVAFkmG18kK/gp3CCzFTZeNsiJiJ4ZJ7pa3irF0DpZ
niJaC2WrluWv/mB+U52LGiddRmh8H7Mn3e6idfGD8dMQCGlsDuenS2rA6+Z4vbE7
SOykt9n3mv2yzOYVrjvDLmd39z5yZaJtluQF14b6ApkMlcElUn56CmB3kUWrtExt
lphueuB6NwoNcayKC5SDaFQPpfcc7gvbPbzo965jgQqPFxj9nF+PYTGzwQXj5Jpl
B6L3QccQ5eM7W6nX/L6tgQ2lSlZIGNV1cPuQb8l9M5vkC7hLiVuYV7dJqbbKZspv
wLyXtsVJoyX4Gy8UL/pe0Qf9O3toozo29FwB0K3F82MIsuQMy3hg8BHyS9n90sa9
u7c6tQ0IZzr3DF4WiVG6xs4V1QD0DWhGdQrb3NYunInol8v7epHS3IFJyw+hRBEO
9XF/M49yNa3fH8H08aENijpZuzfWwotd7D2P/bFDAM7Ka6BhB45Gfx1ldjGLT/Ap
1iGonc7xOtVrwMDJn4i56790XWX9zlA5s0GtJNS87FmzMjewqZptokRePJ4lQn6b
/2VqAhXPUHLzSh856kI383cjXk93O0wLVZuxsQg8Z7XJ72Nz23aXnrpLa8uOvgMN
kil8zk5dmy+dalevkXUUYybYX6Eq3snPmLmWphU1C09UWFz0sDbgwsIvtnizllb3
89gRsE287PagZiC2wx3rAVznGwc1FQoHBWCP0Xrqwp1+55IvTEQLNiaAQ0VnOEgY
ji8RIhxTiZVKXs0ZQtdqEV6r39GZ7ui0BEMRpg3raLeuhNMTiAJ/5pO0Rr++NVNB
QK2HloJdkpVXMax1xjcCWmBsBi1D5Kbw9A72mCO8HYP4zdL3OTxEthePd14qp5ox
aeJR+V34qByaz//JcRue5CpqkwNqFvWgjVH7Ger3he6STANVMkhvnguXuzbSPng5
+24l7+uQy74n7lbyaL/AEv5LaHYUI/gu/8mqiiz/JIWTuQosy/z4HAuuqjnvlJOj
PLJk+67o43WQr5p9mN4HohrcnzB3GeUF/E6+ZvFSnn0VcXoFSOv2I9aBSIiLlN1z
ADl1Kg78WnGnfybptO8J4FPr7fxR7legeIoVt/2yaFWhVLjJ8vk8oyrG4j1PCoh7
AQ6VDEn5LIkNMluLDa2Cdg7Py3y39g5A1S+Ap+kKIaE=
`protect END_PROTECTED
