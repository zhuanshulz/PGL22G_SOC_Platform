`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jllyvVf1uX0U6vwfHjszzKI3zkRDFL1WYFi3o2PQw2U6mEuuPqK1YADWNtP17muY
4n626Fu8mpxaQUXdX4LamNRt1EwVfzOd0P3+4g/sSo21xnKNcH9ui9axiq2rDpJn
DAtfeMlnp9hV7wg9NP3xdPjL1ARhIRVsNKHmjXaStx84H4j4xJ4kHljOVQ/I7Qaj
HiKF4iMJOHxi3DRkYXiSlvdZVRFe9y1I3PoHbB7cXFNNwdm5jJSWdPCRUgEnHkmp
gR9Be9mEwQJlTC98AQpBAyah8S4sMir8eRx/JfwyZtLIWVmZhaOK7amuvvlKp5RE
XJARBFyDLpNPGkiWqHpBNbd6qdEA943GzpT4ys1eGsY8z8NsX9dRebGyUQM+mHnZ
6buzcfT5mrIH+unBq8wKTIjfylb22n2yJsxn9F1Dd9124g+m9imz/gF8HddQGxqe
EVLXI8q+zSu+sNB81k4RUlrpEkmVe7tRfxM6SmKZP/1GnfMBi5PWR+4kbaZXO3D0
xCYjVgKN1u8TGZT+q9GwbbKCGYH2KffRXbrZSFuIroPwkhHTjTS4z/t0H0acqqNL
pkyX6g7AFOkTUANe1aGV0AF/pcsHaVRoC2XdgWP/qupU8KeX+oRwO914gLmpIig8
+TX3xwldBXXZwZHx3TjE6a5xTpYxcv8JPpXQyCdBLjxalMeUu8DUUs3YjHZny4ok
pRaCIJ6lkd7/SaD2LqeV85aOFHq7JN6eWTPamZS2Uzs0DmbBUByHztxMxo1rUGBt
xV5WDQ/kbhA/ImXE+XZJXxgadDFRWLbVHQHQjwopVBU8VkL/rdv1pRQdEIzglV47
6ysSbEtLUIkgp76gqzrOYduCI3V+SCFXMdIlFXFy5h9D4qkMxpP2HDZRRlMmPjxs
j4cfCa1I5/DulUhV44PPdlerCKv8qVV9qDg7qHfw4BNdP7TPBKkGhjHFKlK/CusU
shwKKlaro8Ffi5e8cGi+18GK1y21dvyTuo3+AeAoUUWIB0YS4k7L6jzhyT+nJNgW
`protect END_PROTECTED
