`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kM3WXKZFdcqJQ6FEykUv6oEJaxYfsZOv7SJ3igqfNrPUkFdvVOM/Yw7qyCmrM0rL
oftIv4snvhhDdHnBQLChYFK4UeLrdncnTy40qAwsNS36uGbed1KqbL958pN0qGm6
Hl8GQlJnavWU0b9onw9PoQVtxImTgPBqj97+z4RAU8awVcnilTUowt1YzuaPSAf2
H3zoUqD1RyTZrqvH+B2MMiiPJajWCWhYOKFAKXE7koHE5ExV/VACnmPnqZ2VLAnQ
b8CWXJ/SBMTMrqQM9/cqtxAt7UeXBeOa+Ub+TMXx+xNXWyVyodwnPutgrlsUYeHZ
pC/J8CzNQaGZnLguJ8TflxOuRYuwPoaHKi2LG6Px8H9B1i1XzoBcSv+4C+pnG4O9
Rflcrbj4WXSheFuJJ8oMGGopJju/qdAAUiQfGcLTODw3+GCdaIMDBuOUlICiIo3b
XhhcYbIlaI8b34H/WPIPO+UYPW97b61spenWKSr6v7nLnv0ZBo0GH9F1eIbNMMH6
WmSI+a3jQguCcLPk9qLxcBBecMab0zMEmeabrWTLCaRZ0TAjJ3shzuom9o4cxvpC
IugyzJwn0HiGe596myI7o5vcpAFAV38cWQXF4rjtJAoW9RNDiheozVpOH7wA+q8C
sMod3gRpiVdLCI+sCF4/sfyxehSVt/GeT3vdiawjZF5CO7nzkEBX/8lbELMIcX8j
0H9/nyYvUOOL9wblQXpuvacJZVCRgU7iNWJkctAzCcm+jxBBlMjZPy+cuncl/XXC
pFsVFPFU/k4b5F7XKvJ40BPxoMPUS/STmRY6Uvtm7kggdYnPbt/vnpmIUSdYhOwb
dPgzbihkvKgAKuwk8SY8OYstXJDpCiSbe43rXyipgSDG7CNYt3eNW9F5/F4J800J
ue5MjL3Xh8XZTYkKEZOUTzbJfM0zl9rQUBCSMqX/vT9NDEYfTnjB/kI0nqvav5Xa
V93Ir8uKXJPGlD5+HdCfkBzp7p2JNZfh79qC6wIwplqUUsvQGSP4Z6X4n7H15Pgv
yhQzlJLCK8gvBD2GNkzAMH1SuJuLxRsHBZpnKNb882LkGP5hW/lGV4gQn7BTPqm6
B8F0w9QcJ6Hw5h8fgZ68Pp6f6h2PT+25m4FQj1sK7WJghHT9pyDEGqyVtK2y8//w
rHjUPmvPTmFvpa6Mz5KMQRHyo2sa/ZDfKzdHAfylZ8UzsMLDO8PPUI8N45w0ouL6
tn001HElq2eenflPvBEOF30ymOC12lwPc4arHAVmPOehjB25vzMQBOoq40v0zCoc
CIk6xAqkoesPuH38quE38aOFiw4YDKgTx4NjpYq93l0FpnZUZ9SrPmfJ/5B2XV0y
qokx7h28v1BI1nE1FSFku8hjA3dLYXuBww37sX1h4MM=
`protect END_PROTECTED
