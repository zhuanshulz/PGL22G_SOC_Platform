`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7AB0JBb/ZVMV4JxGqAY9xuZd1e5LCMPX4ja/r+P/4QJQNOYK6akIy7yxoQkPpJq3
kVtntD8GuPUvwfg4e1W3bEF4Q60PC0bgKOYRqZPlEqHvBbi8EJ8tXhmL7giU1wyG
IpLPFykIVSzos1kv863zVhG0pbRQlJhiB0kst/u/kRj+pNQ+Z95cDLC5ZVD5N/VT
4rXQYA60b/C74vZcFvcV4CiCiWUX4ly4D944lGi984JOwqD3RaxYUjcGYfLUjgov
aLqJZ03rsHlKYTQUqjDd18WxT0+VJLEh6IYVhaUOlHGhLu9PeGU2cyHO636HZ/nl
hYEUQiYGgqkqgq4mCrbnUAhgnLuvpNkVgKPtvtwGDVeKLkcLSF1uXyTCkFs9PcXE
VFmN+HT/MatwOZxIQfOl/8XMZ7PU3nF5f4CWfmst5Em3hotYjU3VGUCuzvM/zlne
9/QW3syErgaVIIQDt7z1NyJdcko7SCCMeQxig6D/53qt8orM6PIWgm0cszzVt/kg
bpINUJYTElG7xRPFclVxaNo/YgnWGufm+U4Wtcbtbzo=
`protect END_PROTECTED
