`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2a5oxmLYY0S7yuQkTJyhcudq85YU/S0qcmPkBsHXn8IkpJAtXlM9iYKYvWiO6492
7swoI+ox6tx7OkEnkA+zJv+RVbjiBqw/fLowpJnpuT+zwbboyN72kMbacTSgL0G6
PKlRCDosysOkwMuXg5MdSHf7qpnU2vcDDpQx7y1Fxg88ZJcl4492sawrd5KQnU85
snUGxuJO6aNRRyZVD47O0+r7zTXKzsr2CDUtOQztfV7xDk33a7PdL6MXu60gmzp8
nLUkmfu9LAD0KWwA6tcKX8no+8w0h68x6rHY7lc6hHmfqasUoB7hek5M2IeAC8J2
bkAsMeM4cmb40ASwWF1zGYgEVJpr1P0Z2fciprhhY0a2JdI9CM6NH2ja632ro2CB
DqSBOxQfOKJSDPHNq6mgO8+9qjuDWH16QZkTaAia240x/vfhwzSCjw0NrQBtRKlK
isPousRHkhZ+Bu005rmhxq3fxWWQosJPTkZx1QeDjBHkKHzk7OQ0D5GZuDbBiubm
VA4gRjU+bYENuO1qlPJOE9m8g23zXD5fkFJdsOYfhEzdwsSeltLTBONklycn/fxc
k8DSVvih3dOH8H51z7s2sp6+isin242dgrFr6zZAoCkqTSwwpv5qey2E2yR9z4gO
vhNBDp26qnlmskmjTeOW270Skq/L3pY3wvWJ+wiMe2oBfhcGwKtwcjLzi1D9n0FV
s9++abpS8xDPfIMJ2i4uwy01gXTlU1FtkBz0vopkgyTLyQ2e/+JLaaD1NFVB0mo4
nfXOkUWMlTGSSbdvdXT06UrXilTZiSS2iiyuLPjAQ+CgzZS5dhxlOHh2/Dj/dmTp
aA9lkBZQraNo6HL6lwyWNTE+Uim4euelsiKbycl93hD8UX3MoxYCenszExH/CD1+
GJv8o3IlK0y6BsoLH4T8jN4g2pVkCYmsdlf/AIQi7Fkxor9e8dGMc4EaCHM0IwZT
jmjS4aqUlvSM2wbluTM/CWcMndEoTJEyf+rAZsEyZHuxnhrkDjvo3x8zAd7Wo7hS
HM5xhwblgMUNgzQFW4ROrQ==
`protect END_PROTECTED
