`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rj7bnxseUiGqBjdm8J4plpLBvFZKRjZyugP8sEZQFXJg9oidO+O58a/uQMTMkJj2
yOeQxGA0VvUYzo3zlfFRcdIbyBIHxFxrU4C0Zv7qcYanOeGe4k8fFWD/pt+v7uqq
HlFjWDan9s0UDtsCmn/rliuhRT+3hGj0g/2xBNRJY+bYbFX03BEXb+ky3Hwd96Ll
eN8meWXKIF+FK0xHIP9orhVj/Up9cvDcHdg7C+mlhZmdskuuhrlnxR6Flv6Dtpla
z92wg44UMpYB8p8F49zvP+VwjN297DxyIAQRcDxWtz5dzjsYuHO/jb7lxsjR5OMk
2KYgjwPg2Y7B2C48agJc5oX7Yd0RazIBpzlJPOfCNaQb14zTFfradHthbSrYUa6X
5/WDBL2Yrks9gO5Bn/Y8ZXVJ4wrUQXxtxMlEWzC27pSWDfW2bDOuIEbprbaj1fA/
RABPvkdxHZhSmh1B/UEims5nT+8LvNXWul+RcXJ1CMbezO/O4fR3+TtFAVd2+JP7
Zid+W75snO32g6rEgigiGe4LW0lZFJ2FdtvrOHNXOKHOKV7jElPrTQJesHufSczm
24tNHDp8SUnLO7UA+r8+kv4R3cWSYM4phSfTN/vgPDKMtd+0Yd22Pjdjs870m1KH
xp0EoBWDbai/6Jj/4FGnYnnkiNpknYc1/ReTtLqVmSNfZUK1PeVTZEr5TiotnAqV
GL10wvbNi/hTtEFiOJkxKEAKg5kYSFBMifJzO6K/v49SqibmyMPzAgd8WYNuXy2s
uF+lY/9pxrW2OmpQUgtRf+gBmwv1EkKk3kCLxW6PZmaxSacqD69HdynxeLehPlQ4
s9MzkBEDsJzTnTL263bpM5i5rPLtv/JQUrpT90HqNT0B+2HBHLAl3ZlpHxHgfMU9
tcPHePX53hOQk89kTEqvOnFPUgk3uPZpmJKXwk9q7RBO4CRhIBReCht19hlFlQCi
NReJKoQI4xFo6utEVCY5btnPSpw5aDHYJPoFylHSMvfn71fAPQ+GbcpUWtCGrIuP
meqkScr5smfT1b7bvrRaDQO1qAEt14wAyjurzP97dSoqgOz3pVKUmNoJz2Aef8WN
+E7dKfIqjG3wSh4R1LGXyq66Sggumy1nBljEEhlAWGzoSVXbtFbseR3HdSI484KP
vyo5d2zP06+zmxNagWfuAylN34XC/vulwn9W3XmGnHINOV7h6xubLlfhWZwX1o97
un3mhYehaO+vED0BkVuayKINT9LHs5vUEBQz30BEbiTSXCffFfPGPQSau+b8cUO9
VeWKftMcZgTA0zUZ8ANmXBsrNGbtp0vgiJW60IYJqRvzMSjMjXWbUKQie3PVC6SC
fru784gyxKdSn+mQceAFJUAFzHU0h2QrbbSFsqBUtg6BHEsiUcsPWD9waCjXqcIz
t8y8cWocA6UpYoCFfeRrKbga1mn4RF5d/mlsgSWISeuoUpX4TDThJa72OCG9pgez
DZ06d3iJ7O5QbIIGl+ZRDi38cMrvzy9e78Lv49pdbyoGG5oQt0THnGm7l+Sgjf5A
2QRsT/Oe/RuJ6sjWs39MvRorBYo22YwD4MrkCYXQfNCLXiuGLK0bnNd7+kk6FgSz
iSBOZlex7wKXYzn44aR3Cjc976aPhpRo5SMypqg9qqO0m6p445Fd6YQ58PIL0i0S
m3rwgwvo/M2dDIlp+f4GI/qo/QxCH+ItgKb5TJw8WLU1tWwxusKUq6TxC5Dl95t7
nlKs95GoOrQ98ySpV4/ass4085bPu4P6xkH2DopSfFxBkiorRNfcKOLsodomZBVd
ssbygV7iJnZ5FlKb/lelUNMrHXWyL9POuP1zTSHWzAja91sjX7bId56TWcQ1MuRm
5qNOiWjTzjkVfCnvYecrZP7dZ5I9Qt3LYpQVCG+Zeo/Cho8AaOkw9eqlDoGVzyFt
BVOauWLOdZsiW8g156d+irsXIRkNjp3A9KidT69xp9zVAm2u8RkmZ8Ceimahluid
FSemR/6T0XFEqhl3DiLrHsZFpQ76hGSQ8qVqf7Y2hInQxKw90cdoPpFBZe+7lD+D
OXW/xgRX4mhxklegf9FuLCNRHOyp8OsCoJY7uDbfImaGde3Dc+puVqDwvmeyFDS8
9jGlTujCL+h/Oww8+X2h4YyqrSnrY+GDtEth8NoQ3EF8M9nNRsKwTYQuP9rpMjG/
5SmaPlu/KJmKM23VNML2v9zoGeXMfszowIOHnvYNZPM+gCGTE36u2CaEgjaXZ3CM
9DZ6v6v+QOzhldqrG/qcWj9hMgDEiglx5HMaDMt1ROI/XYOoCYmeHKSWooJ0eyL3
8vv3fiPVYnO5Uf6xIPvS9WuI9xwcyXiRz6WOxqGyRr/crrkFKcDy/yxUWc5FD3R6
4VCQOJvxUm+k6DTX3ZiGLNyojcx4MrJcdjqwoKSWj/R8PniDgD8QivTpIWN0TN9n
3FF2o3Tq19KWmy1gYdp+rr0BkRv48nwFEcWR164a+Gle5g3gcPmexqlhLZJTUlkU
eAdeCpVJYWujPnCmbOElMUssPtMXIRKk95tQ08e9pMXaKN6ird4KLCVIhOTlbML3
H049YOeeNeKxvU2udEqKTFlnSdN+0GKBPOv10BiwXW/bUNR/I5KI8ItIo2JHf7e8
FuWNYlnRi+ywuTmJd1JEJf6JPNbofjE2TND97VL24p4fKjX8et+Rs1fONQpCcHid
z3uaGj5RYbIKtcwXrFx+msg91o/pgMgu0bJvF2ByIfX+rWQh0VSGtZy4bODKR6ua
fE+TWqB+HofdpYnOrPOuHv9EyTrxUelJE9rO3tKIFQ5BDj9fCR83yWBKA1iwEjBK
CxzPoen1LyLZgF+tXtmRXbQ4+8ye+TcAwTr2g+ZN3q/RnHsrx/EVxqLmvrZ9QPz+
g+4g5moWs85jtyOlMDs1CRRm5RCs+lf6ufdxU7+BYpZvn4AaQ/ylKWuWwSUkNMPh
vgeuB6+WiZukyAa0m3XM7WNZIPJrod3huj8yNgx56LOBMlkQmA2/3h/z03VU5S2f
FLWAp1zWZAqRld9xzMdMLU5o0mA7lq3uMwvum90zY1tg6eONVIBr9RKzybmQDY64
KCxk40t0C4Mjk4HBvdIuAN3Xn1V37tiPVA3F7nYK3znTyuWCKKOJAz+tSa+fNX/n
zzc+T9kwEkLzGzElYCbM+nFL2jfjjZqdSCXsXLznCDXPqwEwVv15asluD3/RBfeB
TjAZcGcWZhxQl7fk3iyQt2zUEKZz3ZfgOYMLUzFJEBYBoppvR5skoT0uR8eCEsSZ
euZsE2AOrlLdI7xNiLet1jb2SMyVWP2iNYPwc3tuNqMsztXX+7tYG4cvGCzLCHLN
yvnYw7+QBTV3hRGg2tj/sAEnhrJbdBGphdNgBqR7NUbiYsaOnjqdUFjY4Bd2FYcG
9LQSoXqJBVol9CLAxaFyzfVAuhnMiO5SKA8xVRXaAlv70TAkjFKunK3wjiEIhQqh
sx+EOPZ2ByYXlN3Gd81vMcWWoYyx9+bldija5xbhk4cybGG7EX0qG52Dh3J5JI9g
d43XoKTMUpdMNyiPeX8paOvcqOBqURzyXa/YC5MkryQcJy/VT1kxj97JcflDP8a5
lp/eG7fmIQyg+PfsXLU+eLB2/otRPvS6cPcHcpLD89dZbmapcuY/4yhVez+T9b1g
atQnpRRjktw74Ps5/jjcQEYd454brzPk1GJz19IH/sJjFDIvt74tkrtOHp5MTQQD
II84m2+0aJngH4/vylsdwol+2+8i/+uJ6gw+1CciXRmo0WhxIPfPYDHfuQSiB5ue
1qLZXZbSidMeNJYV0a/CjmKVAWT4/VfMas0oO1FjA1ctJEemkKe2S6XZijdXrrJ5
LC4nQJFjNGbpoT+F33ri1PLq8PZW7uCUVn1fixxmaVqw1F1X/jrkVFlEf60HI3zb
EWaN5YVvEnTkqp0i1uGMzXNmv7nYieaze1LzUCGoGoXgWxLWEJ2XGlxzJQDdFdzU
QmJpE8DZ5dbGg3ylc33Aw5Aopw5LR1WcNQn6XpXnDfqHXUR2xg5I12ewIpBxYhxh
xNbQqZ0j/6AZGHNtp1AuH4SNy13RJD9xsCimdq7Lh9V5g72UlfrBkSCZQu8h6I0c
duGYv5VIiGGLNnxCtIwGtdHogcwJSo5K7Egvvp6dDvYLcDSvmpFBz8FxW7GR66dD
CiKajgB0fYKSY1j8AfZKu7JSSlxvYjBRLa2MSifmKph6NST/3qlXbQbWZAZXUixH
waFKo6m6Dh/mCOEsGv3HpURcsDjh2EG96jvSbDQIfpKxeTAqCE50f6UX55D4+Myr
xGjrL9L26L0FRGm73J86OUrTOXH74GgT6eieE1jEXnISoClD8enUYN5IjWBpjTOB
NPWUTgT/S342nF/+QO88Sf9Uzf28QL7kanFM6oGipapk3Mt59XYm242pC5oXxixL
0qbyIeyv9AKUjBi4Kg6+jxKZ0KybUkC4nW1bq9c4DDEueU9/ZScX3GTUUPFl/7S9
0bzIRuPnYR4tMjdYXqxfZg2bUnEnpTZfBR/Hj59IjKbnV5ESW5k7fnGZ6IBQs/3G
L8t8VYA3jj0WLZRsOCFcHYzfKmSQ0YVLsk9ADDSSrg+XBmLEi+clzuMUT3CvNS/u
aU3nQX+/H6jnvLFFRwFJ5gsuyB0JMNetN/Q9+aAzB68LDqw+HmGviXqjdMlcwCDD
WAXPco8J+IpCmoEWWVG2jWkl1kEKh8Bp3MzmcJOJGy9dnfk8Q/SwYgGqat+WsJdB
OYi9TcmrXnjGIquL+JFFeGFfGbn2IqKAQxmQ0LaGlg3CG6Z13BKXbsGRRuUFlsGP
JR85gXeo/9IpUQbBUdpVJLgq4yrXJMnndzpDp9MY+OeiZT7NcidDsAx4CL/9FuH8
GacxyPkh/6cjJDRtxd1+3sQkw9sdXDlPjd/z69A5SufvbCZi6DCpdaa8Dlgpcj03
OId7A0OEFdaNy0lriji0TipvvcP83HDUe4s6hsvqFUmzVmpnOveMU3566LE0QO/E
spGhmZEgdFDqT8U7nR4yX7wbRyPUyEamaF+E0R50z4QQYx7S/61mEUl3q3Jf8hbo
1Z1NH/mfUqpyoGX0zimiydWhCsXhnZbKq/chdAj8Qap6sMZ/uVkFXkBRFZDo9KrB
yu2Qu7PTJSbXmotYq59e/A130/ToFjLBBIjuRbrjGtTTJvMFcxfvys96iWokEW9k
2zoDcGH9D1YDD8mz3/04HpyE4KzDRKGfBLjYVHBtRHQhaDVyVXGRN6qQdSmkKzIu
PyLEuKR9dtWZ2IYiy4PuCtc4hQQi7OYUqPtiMDN3RuAI4XtETMM7ltx00tzZfaUW
mgVtHImYY+4v78d0myLRRlfa+29Z30iXSZtoyAnlsD6huR0+q22K2o/YvrY7PsHp
0TDSF7jy4Xoc1WETDnsCit2RPGc02pQP9OC+IUIIwgGAOz2KgKbH1EaJImSdj2xz
ndZw4h9lIHishiM6oT8ghqtVZhyMX3KI2MhVrfvN3W0tiwtaWw+BdfZ0cPx7q7yr
7RpRqoFZf9UlD9yMcHI6FY+XDb3KDWB/lc8JiiSya45pIxdkkEMJehYqKGGFXMCg
61NuU/U5HS6nhPYy2q6dHjOGJbkjYBv+hHOrGXtOCBAXWGopYjiYtN+2WM0lQBr3
y78Pth3n7WY4aJxJvZFrHFuwdYTpzjYA+k/gEAWTmaQmeGayMQSrS/6VxhyKl/Od
KFrcUoUXdUxxZvj4wdQnrdf6HAj3JXTirJbd+lT/LH1+8A/ZEoT3aFUSiDD4Ktvg
qpOaeWYWSy6Flzk2WErSdgCEVPbogt5UTix5oIJEzJ0pt4Y0LBeICujzPlleU71T
vsy9h1diafe/i0N4H6kR8E5LTXVe0Om+WI1ezYb6CkWllg2lLo3GL81yLSa5okan
KQdmvlrF8uY1QZfH5MiX2m/Lvrkx+DGxlPGdlvDMKgI0sdpE2Wb9+lXt9t5ZtiUk
qdOqsFLDgdhjTNZDBDFK2GBwoFzpH/Hd7bnvILPjld3wnQreC/pah0ZX5vxrNUlx
eX2l1S9ni1op9fnJeQzIdkfMicbAQ0DV1nT/qYMSTDkMgndoEHJptiJYPPKreQTJ
YtY/j5P3kyAa7tMG+P+Uj9JzlXXjPAB8NVrWU/jGnKUXqIRdatcS7Gra1382seh2
9asO2Hc5hdcJHjS5Mqs9gSdJ4VgDOcE5Bj723FuCS39nORLfuXXy/urzimUPyO07
iG3OpfFUkSztpgwtEw+c8fDfYTTAJYsCdDhb5KuqOizfq+F/9AKrtpx7ZsvX/wU7
QPV5Cz4YEFyNWGI8WEvWs/c+uIiwJadZOc7Bxslb6D6cWEFm6oDBmeH7SFA7KPrQ
mpO0C/KhWBRBuJt9Ok1K9/FcFlG3zgDTGqD97ysQhgCLI/pGgyrneOSFxD4970hX
odPkBhwa0XZgMafI1in8PJBsvTY+nUWgFr9O7RTgxvTQSFkoJxSnMu2WP2qydlH2
xYjBFz/Ca/7UEL/qJh8zi9Y3/euhW4lm/NgUw+yZsjrhkkD8iWD8KOsNgYoLl/PM
FRanAjHh71DyYPNwxWx3Smup7FD63Y3y9aOQTW4Kl+c0roLhKtXI8a2QSa2YEa6l
AXd+nLnfNGOFLNI15W9eZWIPGm10jq6HePBKWYRzzctXyzE4+d2ghE0EuKlS1MBe
9H2ihQzkN6MWP1pqVl4VWl9pC0I+dMPZfxkOgS1YSl7CUGL3KNB93bTmNhDWkv9b
LiGZCZyRqdJz5PpFJ8nI9Aa6tbI+np+yW3vK2BirintbmWHjESlBOOzhuqlEVioi
vrWV6Km/yjXdUr2hdk9r+SFSanE8tpzyS22E1cUB5JITahzEMTF7R4dOtbA7NoAv
BhSm/K9L2Yr6nA9w7TZg0qfRsCtP6K3/AzcNJO8dIEI2pIV8e41RBJlLdjEfMTdQ
J6OcO9U0Clbc64m9dSJRRRl3Hz6vTleI9s70rD8Zq4sRyhjQvgHm2LxWUF+yv1z6
FOFor9gABLqC2AyVAyQWmtCDRKLSwkb7pQlbmIh6rx314MZk1rMLIv8oxfuMUL7S
HZSSzysv5SD6KSYvcLuc+Q/YMWnr57Qz3CLHrkGHzv8g6uaMPyCg6Ljmu4B7rOJ+
Q4e7phuDzPz0xA2nE5ZXynRKGpLLopfGv/Fm4EzxtPoiqvc5PuJqP0WUwPRaTqKQ
CgdlU9MYDQJ2a30dGaMr0r4N/2wpmMYmeXph7i/bg9g9T4XRvT1TPbh0Y/VYOiqt
gfN5VtXgVcasgBluGhClmI52/OsvWHSxPVgppf5tz2ZAfDBcz/M4FbgnoJisi1CU
j7mDEHgeK0QbPM2lCwMJYntTzZ6M14zwjrw0BaGE3TaIyKD58d3CxTTOWnSwXA2M
GjbOu/OJG5HK55ZZnefGqVlWnhj3LxQkltqe5KMBHKwsPM7pOLcfQbNevnUc8pOE
mZGWpTwxcId08TTF7dgqPJ9h9JwNLnu6vdGX81Ivok+fBsGDSq6Cn5htRlT1kvYZ
zw7JI8Ly8TVErv7lhjbKwqPWWyjnFTBd9phP74WRk1FA4omJONyJzUetlv6MtCxg
l77+l1EkrI5teRJWWTt3NXNyH23WGwbKTcWoPC08GQKqx15jbyCFgXs9GL9fHcIN
M2Ft2CVG/8kBV2SX1PUQPQ==
`protect END_PROTECTED
