`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z+8st1DqCbaAu/k+WJJmcUjODqVVdWIAdLXc9eVQ7xTXe+W9HCIKqihjFUITVXQu
cv3pZslNcw9JLyozxEmjYmmXW4gMpNWufb/E+aY0+Tgbc1vgPZTFkDINV1TlOt3X
mT/ywTxz/v/JdOz3Wkg1mLOwXMSb0yHrkAMo8vlw+48keMrBO3v3G2YvzHn0WSOi
KTwIwfvi7jBdoLEG1Z/2YbY8xOMPwAGWciPTpq4JuXgPmGktEMmO/d6aWTY8x6F1
jNFfao0fQtnTF/X7D7unnr+/p7G/4m34XUcs2IgPMkXzlGT2rtJpyh3SaWkssCFK
m047CyOmepfJHfLXiegAbkTn19kCrB93VbbQLwKiFmzN3xc41CswsML9o84VRJ3g
Ef5VmJcevifGxVdmE3hO2y4BsyWpZK+WSwe9FoE9gKuqxZY96qUmvIPHcsC8eTZ3
8ARNLtziKa7xmWV1VHm64Lcq7chI76t4s2tglRB1JnRuAQm3ynzeQlRR7dUruDfE
mHUGgpIcSME/ewfl9v0cFavYd+iAGMdaYiQGLXgR65tnbk+I00Cu0Hqzd89yGcam
vOZsZ5uDWOavWZBv32gjrc3f6Mgd6dk0MJNB5XiGyLy30DXlVsS9W5Oz6jUv0lQh
OHCCqan44IokOHUNcz0SbAV+MZzmTkH72kx7M2YVo3A3iyP3YqYv0xTnllFOVRJv
o9uHU0QxGsO5gWB6cZPJ0tn9mGEeBxrxnVAa9gCVETI5EKJjtA7m/eoUtlFIuU81
mZ2+NGgsguhwbZVwA32zbJ6pJU5S7yz3FeFLwrpeNYso8jNIL7tfPcbxQhbG2Qoi
X0f3SUisoXjr5k5fVGU+0c/PDzRPL7DT0E1nA424vPV1fmWfeJvuR5/9V4XaZnw8
0HemOBBrlIqylaGirjoIQCsumV3qwfHIUR7emVbinz0=
`protect END_PROTECTED
