`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ULlvRxbOtnyIIKmX+HE6ktGcg64KmfP6YWcttXlpOc/R2UEHmcbCRddjRQRwUf7b
vHZCRY9owJlc2qchAfLjawxER10YvPPdYpaRCfTcb8uNAYaaJq82oXs9sinOX90k
HiE4V0LcZIXMukk6EBseRt0uXdAD8boAAnQN4hHI9S5D5wUEkbxfW+L+RwnJEQ3b
zNhlpXbjx3YxxbgY0tl7JcB3l5s9E3CzaTe+NY5rkkMujdnBxwqLUzTHnddz3kM5
KCSjNFJVZmr2v3jH68MFl2BI0L2BwLTLqfYaQAB+J1XviwETt0EYBKWDUt/gG7r7
SWA1Mx2AngHGh0CKk+YPlFV3VBNHwHSSR7YZfW3SomJE1Sm6WZjm8OH9Af59zHnU
yL5bVgECDP8Aun+2GajpqPDuhOr42eVqMRxRNsa9TUBVv0Z5zEnrKGuj5iQ+y//i
2Mfwo7nCTO2IJeX+7lXyvwPbpaj4S0gsqcUfGREPy0+XHLV1HbpOzvgo5+1OhjLc
XX7G9//NEk6GJ4VIKt9wvYd5u+pftLu/kpTRCuPfezXWg2FNQmyChFP5XGn057QJ
tUqN8488K93M4O1a0lmhAWIhViLkalQr1wzePeuaTwAEgDWue+lES/xlLNBrRb26
KMbEBZUtWdd0+GNGCMBMILjN6FqflQtMFRaShUTnsfyDyr1kyFIG1NNuQ/EjOugF
HBy4Z7XBCJNENaYH8oxiNPCjrikMc7jYnlyQxPP3jv0WxuGJbmQam9ObMXn0E2H2
Zt3kLFXgiyfX6b/Kx0EP5zzIHOJHaBHZwS81NGbjhbC+R32jVrrLYrdGsmaOYRuN
+5OYtCCcbqvqyUHt+47q5N49yyTZLYUCMEYwNOHtROmdZi6yvThcaZFzf72PCJGq
qiwp8GzqBaIQ4EH3Irb6HxbVJ0ZLpggyKYd6k2068UgXAqrhvtru6Qy0n8Ll0xiQ
bHDs9N7Aa7IS7e+yRRKhx5ETP1NOysUSvgnNHYOOwQytHTg27X9o1I1VmLaEJ0ix
pOhMjOXueFotqy7+LlQR/HSrSwKlvx7Nqhoce+bpTUVgoJLTm+zrFybprtUVeXcQ
x15huagrUK+EA7l5VtDUyQxXEtwNMzOoL1MUniua+78c0rDa+DJf94929e8v3UB3
222Ii9DQkBrqtLMAk3bwjs2YsOVRfSqTKdYyp/wqOCil/hXb44uJcEvP9975UDmh
fLIdjzrkwO976+1B+Cev9SZNWq/l8RlUS2uh5RfQayke3bSPm34HkSBJdMdXluAr
gQkdF2qjmSPONIV0yVrK863JBYIUH/h4QYH+pPkR/P5ni0RITUjYiG2L7kJy2S5v
hGnpWjmmW79Fxd7pZKZB2N2ltbrN+yg6ssmu/Zeo3B6J0Ht66ci5xbvHKg3zcCcu
x3aJ8YifLVzosA/4XbE/m3PxasznTVUpTQ8ziDCXB4zJSaa4wnMXmpaTq1Ot+MLf
GWiI0JxWoJL1iA1UgzarhKtTkm96dVJ5jlPiCwvvg+5ECrlXc7FObO2tTWvM96OS
ovz4dC7hdeIFUzT/BcfqoIdMxADg74WpkH6pY52fs9POK/IPMCMIXIFJaNRKF75R
kFpAxbP2EDuPl+G3uZG6+tW+Ex+Pq6DdqJDZ/+V20viq4ae9lP/afNXqq7cGcBGw
nqKozoU4fidFvYbhWSLS3zH2Lt9kQMJbn9YFrS4E4BRE4psZhkVNZyqF6qcXsksf
AWJm7zxN3WOB2OF3nWqnxo14YzNfGz6OTsadEyOCiwFOqzdKg0Z/cM2fCVsI+qN9
4uBkLO/t2N0CvxRN4/soY52pHlyTm9UHiGQixgaBfzBFKx5+rHFuqBHTRu3XnzkF
zXf3M/3FNTdm/9JtqHt1bVVrM7gT8V930NndnN20I3bGJ7CD/g3lxdeD2SRyq6Nd
UZTGpeXqt5s6ZeYWF4jlGTlZqjmpMDJuTs5Fx6h5flkH/hCSj/HsdCTUxLGRElaG
x0lpKn1hqXkpPiDQojO3pdyzGcx0r99fHrh+UteOrYu6WZr78LUYyNtYAuqlNlzJ
emspLRsdV/VPxSt9NZl2FFSzQ+432paD4sWbe2J/oMJqicoLzTm9OTvatqUYhrD1
QWc1sb42SJHTZTzjNHppCbvGpNkrrWM756GoZk6zB0Uzc5i9KptbEimur5IL5M1R
xxZEulh/0/yzX9y9ILGpwpA6sfwr6K8nS5YdXw05hHxYs/JivCNkG+LxfSHcymYC
ezqKCcA8jGncw6LTVD4GwB5QhfMFMaKM8EtCMNuq8LQFeSIUOteVr14pfET1UJ03
CHAdnywKkyICOoYK2hX3xB05JX1/mGwhM8Xg7gCSMmFID4hvmRVH/EK8lIGtqutB
CV131xtbdmKoSC0+sd92to5Drj/BYfI/6J8S9CO9qWoivGV9rNOksjozWgr8aNJF
BAWq22RDHWc+lITlChcYxOXB1YN3vsywU5naTZauTKL9nOYvdVdFGkZ+LizvFH/J
n2KTwzt2f0sGty+JdfDDWpeAJmxrb5OJuRZy3swtjTpz8srn/Flth2lt3V+123IR
7StScHTZWDjDYGQzwaz/9PBnALCrP7AUmCV6QNVp7bDqnNkyzUHry+mX8JBQG1R6
qJI4vNx4uD2dAzur2Klg1V7PdEK7uYp2221sB9mcTUfvXX4Q7MTG0ixVsMRSn41D
xa4bolJ0P2cvYRgtdMIaO/P/WaBPghewLyWeORVtpxRTI2xB1tHra8/uz3BDWzUz
kMH1B4krFponUHPfyXtWGDA1hl+0s+pBgTh/6dEc49ecbT28pTqHcYoT1DG/HWHU
HeXwvk1RZyh0pjqvyOLrKjFRoClX+PdQAzb+lMxpy0FBu8Qx4h0VeBS4liT49ADs
tvJdw6McxO2xQsXvnhvRSiYNA84kP4JoD5vyvF0WbQsBX8kLegBUTmKisYU+GelR
o3Ys1fMFPsQ+hzz71pjDWoJDzHydXngLJbEZ78MyPd+j4Wsoxv+UlobKgECUcoPs
UT4UOG019hhcJNnGsrUQ/MYt6naXvGOGQCUWsGXSuwsAnb+mt/EVkZ+HV5167noO
C+WOs6AMa/A93v8r6aqaFZMy/c7Km3JHbxjJlghpJ8uTIf5Tit7tjzh+oAVVtaKI
hON6ZS+5aoODqr68qQtgaALJgfWmIcd0hAV6vkqVeLtAEXJ6ODLmwSAXbAsBKIDG
`protect END_PROTECTED
