`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dEzPmd+DEuT6YuyO6HIE6kntXiPh1sahbgE9My+CELYunIbD55o40LuBpDY5Emyx
t7T2GkT/YrrH+3rdcBtA2z4FbDA9o4LcUbvy+mxV3MlBW2OMK9VuZW9kVtpUN1PW
PumfFr+vX6MjOVqp6jELuWaYtoeyX8VX/0VxUlYjSQepZ5p3pRelsZ8bYZAKchyn
oDSrThWbsbiMNZr3ENJqYEndxzfRKai1nzGd6UjTO4tNVTojRXm64D7NpHTFOSl6
Q2ZU+y992AROPgaTykk4OSGB9kr7wY4BmpDgaIztnkEibRXwGfIQKBeRQXChxX+K
xS7inEsQGzWPjObmAnXOimALNraahKnQOGM9PEqx6yDh0vJKhcbCmKq15IxCIeRI
iTq+5Jam7yipW8tCdIfWh4DSWLQQHgkRdTOqbJtKg7j9fIBMPE6naRjIzdIjNh6G
XhfxWoWZY+CkyWG2cBX8YtWqMUZCltdPi9a0pdcRTzn+m4ekuJjsPgOUR6VmKAmf
stbeaD+2bf1VRm+jbGlQadLnRUbFZwDNmr2T+ZcjGuC8ZgB6Ei1Elf3jwvPsbSS6
AOKSSEMVRs/mqznj5ywcFq+A2DnWk+cV0bVNn9M2huhLN3+cLqgaau0cgrAWaqo8
e/XIqx+EWr8Y8UMnD0Gg3kxsgD67BIcIzn3grR0UsBSeYkXIXdAuluNfjrPQ93KS
jFO7BVi1mHSw5YRjDG7f1CDNRq8JgcdjKTIQQYdwTwR4GDX61CPPa7YhqDAQkY05
Mw2DlL+Ym9A5Y4BbZe60SkoixMPFJVCg4VCn49+0pO0MbWAP3RnNLEbivGZ4XI6S
0XvO7FV7B06HaY85ivXz/69eJjhQk+us/7uBxfiK1vfof++xj11gVUtrodCMxtG+
aazFhkAKIrQOvegi546wbee5RCA6kpdH5Q1L7syy9f3olPWFAOXC8t9B6sVK9hPV
SG0wpcbPuRJhJqewzgStNRlm+5klSHsf5hY0DRGDDSBYyCcODuLufz1M/84r9Sbs
H/xPk5X9oINsuu+nfx2nqeJmlsAm1VjMGEKq/cfq5/1iBz/LnmGDkYe9ubRFHmzu
MN2EAp4tU64t8WSUEyBBM9dMVxjRvbwNQlDgP770P1MJRlE7fNKdCxMt8ufeyA3E
wwRt+fnfpFNoLPcD7ap7uc6TWzOAdjf5hv/L0vQiDzqaOqGPDWICDimoHnqowKnf
E/Q8zT2ut405WuV5avj0cD/nRGCRhQ4Dxufw+QZbWN1o6fiWuUCXf/kp9emE+022
eNcrhpxKoLVQJtZpLlc+TM9FLfdwCMEjrHt2EDSH8CfMDusRdSKYomg70hc/ncNl
jDZRcHQKZmzdyskRuwlJOShzlcH/5whCBIWhe0SSllOBTW/Y+PpeYYxvAnvXSX1g
2hFya8d5ABMlIa+cVnxZPQNklbATIG26c2EAupNo8bUBt2ENjGr1IcUbOyg73yP3
fw5Cl6tyN3tM9M5LuR/cmsvQxZmYy1D0T+i0NfE9amebo/7f/D3ACTMzcELEfCT3
43Y9GqdTtTO8EpiDcARMLDW80dGSDUX62ZIaJK+P6Mhb6hb1f+fOw9+Ztl61kOw/
yR7d3OrCYpMYfOhrGntgrp+3x5Eogh7/ck+K0MyANeyVStDjI90LLsT5FHtnOQv0
L5i8HRpo1N2gHdsgoZJGur6iXa/PoX/nxOLTofJkJVU33JGsVu9y3hsLh7rDKtD3
6mToE2mIIF8oEAQYqqZ3Go+h4oPTBZeWrJCbyMgBzepizWeKmOlAEKhAtYi99d25
N82kDgsSh5UQD7oLSxTqb7DNqYZPAAHQ8kxl/2Q91GOc0ldlpNvhwHXY/C0iDCsk
7Uw9mlDRvHXR4AKT2e3PE9K/VBiLamuO6/S+EbM5mp0v3NpdPK2OUzmo875jIgQ8
r9bgLaZfEk9fM1/E3iiU4h2bELXJMloVszmQnLVBITADML6fBqQVJciSB0760oH8
`protect END_PROTECTED
