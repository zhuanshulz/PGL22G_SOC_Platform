`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWij9GUgM+hECy+8R/Tsyxv5G3Bqvw0lr4+EvvXeM9m4RlZBaC/egMJ+FK8fPsQw
MWln5QaIelb0VCIf/BJAlS4AXUuPL7JHtBUhe5wGqvAjMHB26+hOjNTrY19Z7atu
qqm0d/aaaIYdZUJobkOBIxUGc/flAZegVD7mWHfLqy5AxZtfSDlpiynE7EsLyBhG
cWUr2N0yBQO7B+uPew8e3h0E6TjIGcMCKeuPdjTQRTEWbxmFaWkpjEGcuqY2laCE
iSb4ftCTZByfYO3nVZfKXPKVf+wUYVuqT+UEas1YU5O00axQuEN0pKj5VoOfR5/t
W767ef35yLZ/R885xh4QPw==
`protect END_PROTECTED
