`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XiqlgLT64SKk7o/jiJXPhBejbJZBDgPXd8882FQi1vxxfdGsmHFboHbCnaH5pviB
8rWs9eZUS8DufAbW0DdtwOd7qr6skTR28j79Jf5SKs6ye6Q0Wrn60BVwALgkfgL9
N0vQITNKhVCPvahxcV+nqo0SzJSQjB6ZFL5NYPegPB0lXUSn+oohE0PPs5XHR8Ae
eAkCXN1LcG06ZNHBp7zy4Nuj5QYmsuph7XOL2vPTCO8WeKfDfkOdY8PEKJusUosr
zvGB0uBuLSOocTe7IaaqFvGW+Hvrv6muo/r69yYZ5cGigL8B0Pc/peLF+eOzWCdN
6JU869dSVnaG8gjN9UDzvdzrX2DO1+gKYrLuZsT70wjTlWJgJa1kZOQWV/iH1iAo
FQh45ldfGNoh4QVGmJp+roSYpaFjfKNMjPxT/tkoe8//BDEMwMl4TPP364Efg2tx
`protect END_PROTECTED
