`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2F2OOcZxRGXJwEWjsXaRHr2+DlsdIVCEXwHigZ/0wLmqOGy/EN+xzYG4GoiqBIS
xXFJO8t/sOQdgj7mZK3BxiDzhG+6rNu7rnu/kbs42UfP/XWn7h3rIdXB3DpYUfjH
BlpzzoIflQ/7WwYS7tfPgScxnP3WD6LxNNydGeqBi0Szs1UWvbqpQXu+03KALYzC
nC0vEpJXwfZrQY6UT9C64UoqSGrYOjsMcps+3DLgOfaIRwhbbAlKn3ziD2xe3y4E
893uioWVG+wORCZ2Uq7DfzYm93eHdyjE5avnL2YerUIQT0tZplhUqb0sHFMEyMtK
qp5Ej/CHPGp6Z0lez/Va4BscD8yCfR8tDU4O8Vtnu74tltg3anrp6F35SIi8sZRA
U+fQQGmQiG62SNdrrKeSyMjxzeIn6YtYgTa8ztkI3pQ33xhKHya3iBQKOrm7rpHw
H56qECeZQsbpVJ/LBxXCk0p1nFxP7ffUCba5P1vXrXg1dtRvTemMFClwtDXW/rhl
LrPSr1L2p/hAzU52r0cRhTujq8LzjxXs77oonVGs0SyI2+iIhbQ/EbKabDKh47b7
PB2QOtNZVJ5TFqwwT666Yg==
`protect END_PROTECTED
