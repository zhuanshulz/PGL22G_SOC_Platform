`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMugzaoAnRn6L1W7l5Lt6bZtxyzRM3Swe5i1+EVOpUNX8Vj+RwUoDr7TUHkb6MLc
vCOgIoZ58uvIczg4/0HnCEnyZP9VDqs7bcf9v1RrQrinS3ku59cX6MTqXUnbAVon
p1iqe1Pfc+tfQ93yHZO6KLpHwCgyuxCDPW69t9ZQjI5DA+OsJCjlc6Fgr7gO6UQi
5QDP5tgxQ3sRz/6J5FAE3K6BVhzkW8sm2O4vukdLK+kJYsWY6FyAwLdsYUwHGJqq
aj90URZ164IEZjXx8tKoFzZ/2yxbk0K1TyUuj8Tcv4ysK10Iug01zSoqpp5mxJ4J
oEhE5S/ZsEda1ubYCgf3nhCa0yxLJKLqeKNs+dW6QNAHlGeU3eMJ/OVLSZrAMVf0
XOqMIlJZqxd8cDjhxOzN/g==
`protect END_PROTECTED
