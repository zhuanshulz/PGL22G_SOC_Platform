`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
avC5JA0o47Q7dCJuunvGA+7CF/yfbiF6gQdssGjfriOXVRm/1bjebsgU0nHcJPuE
NJvhpRTritsZ+XiuCzjWNKZwuy65CSj9Pmz7CR2zJ1/FFq/wL9PPUQUWo18rjR/v
yCSsN1nFJ1GfE838TZhN2VllVoliTdF6JgnfSyGDVSXmew8HNAn068bvjjz2Ujd8
KoAJM4XeOpjL6fReywiPVojTnVvn0f1GmqKGTObEukgX3zJSY3kp8JQv3sYXCLJ3
9mQN6Z7DIdmMv/cwEDdyOw==
`protect END_PROTECTED
