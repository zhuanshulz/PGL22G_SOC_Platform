`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dXrhQ5Tu1cUtFWzs5ZpW9BM46KLYiFdT9N4n3bH9wFowRoM+nC8ASz+Ku79B3A7s
f8+hx3dmNcHKsllZ4Hatjb1q13BbEyIXb10REAR9Vac7XatCyZADeGz+aw9LdEMa
TamfYBxlT9XtqYqJPREBSD+AKyISlQA67DG8b7KT6SZuXpmozrpOZN1aN59q4yv1
+emn2i4yWFkiBN9ByxVnHPd8kOYFPnqQll9ho6V6wSctYCjR30UedS7wu2PUIkzN
+nYFQXz897hJgvdTyfvYFYVlpdFNLYituowzgopDvwACq3iWKxB3Xrqnlz+9ZlY3
7lfggq/EXRDOSdFzgW9I/RcA+u1NNU3iGxjvkLXQeRDmd/Jrf3P7jUQDLJjgb+mR
Z1u3PhiWlnqUXqB7xjH9cBHL4kibVK5QAyx39RGbc3zsppeAxuZyRIMT+Om1Lh3C
J1iXWGKCUrnsgjQSBjdNarqzpU9cy8DWx5I8uhumhY9CfZO/q0bf2MoG0eLio0zI
k0YcF/A9cMYX/6wjD9Pj3nEPGd2m4R/f3oFB5fSErHC5Y6A0DDJizRoZ0ewpS4NG
AGAbwgtI0u98OhzFCpPy65hYGP0bXygHm8aS6UVd0++s7Gfykdvc2OkwsqtvSn8g
pDHAzewuK6qbPd/1VgcO1NLAXyUT4RI1X0rx6SrkF5uSnVxxeHjTD5xSA1XfB0f4
edQ7OydUuV9cy90a56XgxRRdnSjMmidw0/LHwT7eMlK3kPoYd0KoGN0x22WcLmOw
zUJiQjluzqeySlznqS4sQKv6nE6tC0ltHiuPf9WvIfrIFyS7AUV9yj9/4DsBKueA
37kGBtNaAsl3PTLVyHyIZNvjejVQi8F511OZUPukrCTU2pZUbv3gsjUbsarGfS8x
pNV1z2XFFYAdrPW2KPBDtLUzjIZCoTwMpPpXk1xaP54/HPE0kMwJsD0gIlmlR7o2
O8hjLtl4Of2Kp+0pS6Zf7QHWtMo+/L96e0yPas3JxIXHtsF8PIqmTOQOq2aynI86
Btp3JGSGfaK8uBQX5U2ngLQivKbskxosPou6NUhOc5sGDLZX7d3sCDcb/OnhVbTp
j5dr0hiv6goxpSbE4sBvrAJIHhR8gddX/NyHk5CANhVlcpshFJ1ivMu4nmFXdY5K
JbhudvNZFUF1oY4pkgWpWfNYdfL+Wmcm72u+gS2bkeqFWEMhUU+8Pt9Mpox+fk+T
sycgJHiQD04FoQtF3x4nSDcOMFJlzZs6g/mCyLm9bXvC17izrYWqV9aQOJ48gRQ0
DPd6q+y+qGEC4vSWrPMLtJ1sdlezk6gP+wVevCnWhbY094h60xISP0l6PtXViC3L
GWPCOp+KBuhSShKdYtab3xqxaZ/Hg5jX9MsNj50KjKcybU54a7oJ6COKuf0itw9w
IDlPY54jolca57CS7YwY8/60BXJmQo/m07HKQ+nYYzsOQK8CO2XEDy0nHHkVT3Pw
YiwQCspUhbU8jyT0T6anJAbgIqMWOWv/HPC5NWm8EqbisKvUNAdh5SLq2ahdSEei
eUm3OiSfr6ZRpH2U+tPXxnDptTcUr5IKKpvvmROalDAJE9ImEco5zqr/6LbEArJy
Eob5dHBKwGTHjmmgBSUSzMmyFlEh/FPaghhvBC29sVKRp6XM/TSdxB5fZ5rPVMQY
EEeuC5SlRb3HmCyoTmh8YSQsk1GT1tXOg/puZQTD1ThIwDdOPdy0DUQbJsSS/n6+
actBTPQ9ie1kTbiS1Zh8a7/SQebHQsIoU5rgrVeDFZn/dTox06XauPwYFbYFSwUM
ll0mNMXHJ7yP4vD4w8h0TsI/lDqfPUWy1K6sX+/AaO5PGbpMMnkIqerVleYmwotR
DJyFOki9/iKc74JATvuktoYap5t1cO5pyPP9NPl1f8deMwIObNXVhCEMt7P4clQX
ROaZISVUGxJ37e2jYvMeicelh09gbMx4SDkk+0RmPPgjQBU6z9/71I3Jo0XVfPec
D3eLP4LXoMw4hYq71X3aLBhkXiBD9JOlg/D5DnfmGYUD18w4fxzQ16OvXSHrOqwo
vJMY2lDo1P0W83bbE5NE38dGg+6eaRB4HuQdjqfWDykXl1BU/JUokbK3QM4CC8Sg
zAkdNZgbeAuiERYwClo6JDiiVc0D3X2dLP/i9hk+zgVxA+PbI12E+1W71P74OxDW
/uZnlGU97xFrbQWWI+qHCcltZLyYdRKzZ60vdw33vGtHjpRDXdvHqNY4IyKU4Ssh
pXJItMk3Vl/yYmxZzqbm0Uk7SSWLLYorCnU4pyQ32Idl1ATcpsNdnMslG0+viVr9
6KuP8SkZkNPIvBX0OJ1JN06+5vLhoDmvSbIvH9kXBH2wCmSWmPoIdm/qogvNWUAX
hX18cjG95f0KDA/i7gDzJkF6rpW72jRSV531c2HD3WB3EkGx+pEpFbmbNlWRqUXt
QE6Bh3Ewxw2XM7AISD96dD3ZvLBHZQn2ZDLj7GZeoiQzdx2d5jXrplCQ5x8O+nMt
GsQT/oqi+rIPN8dc67gArFVyCAYQZlxt44wI3oyMm4KSC0HYCrLSonpvG/dcifRS
yV8Qtom/Oivlqt67NZkWDlBVaN4C9Ez3WjHM03vLGOrPt6EGUm1K4huEPaA0uQBu
K1RTb0lhWI3iQVhpY1ltbq0J5fq11/IiELeqdknqhkaVOVypgzMTH51U+pto2GR/
lv5N1vkfQa95KPcfPSOnqUsvQC+o/2MFqzsnwm18jhcYHpVLSFSocotO6h8P2StA
xJVFEsQJp3zuIqbyWKfdmcHChCmDDytt4BTTAfX8QRMCCD6flGt4pIYU1Qes3MSU
esiCukKE9SurTr2QwxW45JHgA1T7CznSvD0FIF8oZ+xXX7U04zqiRxfNLCXQIAwx
LKIJI6A83X4Em5sAbbxmj6Dwb7lE74cSN1s+9x6ZhjkjzocF6uItG12Gd6vAMZdq
Quq6uVSzfUBnlE9m5omMs9moTRAlLwQIWpupZxWs8nd+IuuczdVwzGA/hjmNLisO
qhN+4LZreNXMHt0WzRXFojzh3fPhcy89Bsbs3iQesmuq0Sjk0eaSYGgCwfvgtiou
Ppd/uzlrUTYaw0ibMdDR8Z7PdvH72nPwFX238clmslJ/rtC5v2ntcjZvy5TJN9bI
TH4eJEU878J0NCOJr/0Pl9fEHIaeYZnhXcxgbaicbnWfZghtgewtTtSmhmvcl1/l
z+tQfK3dAczaR3g8vuuk0iYpQ3hL8q0xyt9pC3kgV8rBSoNpj5OCfmSbA90G6IqS
hvyblXAoUzCeXWWXxHy0gkqysde6qRiqIGS5ceiTqsEaxlTrDAqpqScBoA7NbFpD
btRczoHEWhwVdVoFvb5x/3dJSLerbdVfK5U5Z6a108jj25O3UVqtk+jL4IvRgUHO
5pAhIYUusMhTcblfHIF22XN5/uTi3Qv/pLGIUz1Zf+0Sz65XXnFKWL9E4o/V3EK6
oRlN6pOZhFLfC5hJ1U/qEwnyGYzwkg2noE82Gc4KhNYXNckNXnljy9/nFLQoxWE3
DPslm/O0aggjxI28AJriN2GH9TsLJvYVmtTwYiAkx835jgwF8ClCa1PU1zB2/PFv
tbRAT3t22UvFsrqLfjLBkr1IE8Vd5w2SpNUDQyYQzdOzG20VgP3ihPgP40rjGPDK
uQhMEf24pNye+iGrWWQWXhT2rYNa2pyC03vr3UX8/rCO99sCnyoAxpvnt0hVI7VP
/f5fJpuU67ZCMfPmUiy62Nm/LQbf86FJnH0lqbo+xDoTtVOy5LmQ25sYjCCYUZxE
tZwJSSGLu3D8eA/7EApCVesjyDgw7hWp7FGG4jVsZcgyc/mq/4q3MqYH1meP6ON6
cONlc7oVBkm+GKS/PvwKWGn++Jq50Qh1zRbvcFYhbtXBUFIIuE3T3RW8dIDCMSGB
e9b87jb2fnYRcNYpOBGQF+7ZptrnWlUSH2TeczU5w+9v1sCEGwoD4QrammBpfE5w
Cna6w4oVB/LXhYtzbrON0k4UYBFpGtuhicNKFnckME1S4r7deGnxV/OWXtp8+U+7
CIy87sGxaKLaJdb2CEw/JlGZRdyLA4fPjmF5QXzEChwi7RoiHzTx03t1TcDG1AkG
eGzJm3VXMO5NxU8pRc5DL/dkkKKwKUJrto3427k0D0z1yUZ5SctnEILgK06DfMvx
jm0UmxIC7iztdGtueVGsrDLKRUdXOppu0wEP0UBpVfAObVX1NqI4vehtyb1dmBPK
c+axmdBidnxlJci+jYIm3fesEP6ACr8o8F9gjgCc/6CDk+u5W6tH43eoaR9XnYUi
2KQCT4LzQieaJETdU6qnSjh9pIOqek/Of8NCoDAcCukkn38LzzgzvlXln2zxTNQv
Ol5d91u2SQG/IbpAiN6Ceb3g/cVwfjnNRYGnZKSEHdO+5sMjnXfQG3LWVkWbbydA
EI9kV4KCSnbTVRYYKLP6aXdLVHWt35/WnGyziSAe0DAcCV3yptKa7JwxScV1P1ko
LpDPusHf6OF4rGSq+TtBlIAB+FoDZljyCKSAWQ/7Dh9M0e3LLvsDFo/lrCASpF8I
N7uZNd7bmbX6gqqqm8L4D2itxHoGLhtVeh7ugDe9UGJghJC5xhQsV0VuMPYMhNJ0
5XkUKnUR9i5HDhmSBONFB2r9cj25LgWxxCjfRD8BdDMfp66/X/2+kTmWBhHAWVz0
JSh7eIadIS5wSIo/QfkCy5QqMkE0WGKY121zopkXhpcW+qBRC5Zu73MHgCQ3nPtz
buzjTdj7yWYh6X2KKERBCSdI+S8ZSdZHTjk+bRgVaQmT7ePAyBrMg8vrYGNe7e7x
dQ+f1omwv13uO0IyN5mSEK2Gy4e+wQWrLZzLZYG4UC6DOTZWqaxoiXj9qc8J+gy0
dctDV3cWztnlE2Aqgjdm9cAjLxJkk6fO6X9xiuofG2iyPWjolmmK7gtT3f2EXJFf
hQ6fzWuOxvpJfb9jKyIzkSCXjf11vcjieyQ20eJF+30o7HVJ5ELo4KJUhk8q+Wi6
G76ix/SMhWW8jm0PoOlUonKx6KIX1WusWKhtwxT9833S5csTXfNCQBiMqgGwP3MJ
SinxuEJ6zYUp1btlmVY1DYSyRvsXdly2CymRNMunQdbZ+Fvxw/YF8BnxcEizxQC9
viSIqF6nJeRjqZE/xkZMFqGemkv/RG3Sz+eSBJ3niNkERr7Gw28TU2aTfHHtbfiy
dv9DofbSRFDs1APa9zAu6EGOsKFH7Sf+dLOumYNsqLoKb8em9Xi50waSWHtf29Pz
hbzSjdV5FY8A7qqiuiSdVUG2OBlDvz1uxXct+aFwlYPJ1nL515SyHF2P+QRtY2XE
eZnC46clOOJBulTVDWHskgxiKg+QbVT/EKBLqSeRTWgsQooXlXING/ROwS0vpXI4
FyUW/7ZLtjbzx+RblreXCz6HP3UyADRTaS8lxmFRyFRM7ZShr5U7kazvloiZRXtC
ImAxjtDmhQ6TUfOqeykw3auFWG8Rh+FD1MlbVKxE7CMJpCvKRLjQaUzHsqWzEkyG
BYe/fVai5MlYNCQ94CELcWfd34n2AH9vi45/FBVYGYY8LBF9tt02VfNGKcwS75zf
E7dzmkEyIg8DNJ+TbtBisa+Op8b3jcXL8aFvOAhJQzh3o3Yo5FA2/D0/GmdgldN0
nKBeBQi5No4OAHvQyUhFYcQ1DmrM6Ajp1VPCrXN54EcCDBYc/DYMKXOn6xHxKhig
Myx5FiWhXelIYjBS7PvbdPu5WLooK9EkOeb9GcDqgMms4sucWBnNkDyvk6ZxynOi
Im+H24oeO+WTwNPpmNtmgjr5ir6GnC9esi/MmV0S2oxVUOCDMuwZ15IJ13iZxTx4
wvPIa21NzSScW1odNDFJ1kUzo1Pi6Q8VsSoovw9jiLna5llYHERv3u6vunOFCuww
AVOoHscnGjURqzuDRReAlkHpRbkVZlABxurASf0J+D1iUXrjE6CvUoRl8Ej2q0yg
DSlPUiyiKtPjINXO6F/yuxJzelNZNuzIrWpHO48HJ+GWr7mWlyvjTcVKnHTiLn4L
WIh0CL/G4R61n1ZjoQ3wbKIdhDxFlS0jyLguHpSbMfzWfdA3H8QwECW6zi/uzF3P
/Voi2xqXcDZrg3HYCYCt0QszFR7m3FL6dUh3SP1tWsCp8VOwJFz7SIgDXRI2Q9tE
Up5UGm7roFqF/QoNR0EwBF6+SMY5iJ8/AzekB8T5usCA/xcvSuI4eicVlEqeu+x1
ZLawkl8oeZOYbGFA2g5V50Y3Y/EBfdzoq91JGC9EXJMhbkO8ZGEELFUoMXlGGEa0
+b4HvCxRqFhZ6T+nEuwsdBZCbPTbXz8eM57BJBCqBMQls0H/AJrUH7hNWuOkdpoq
qRCjqZ1Eka2vXohyrjCimlAHGme3A0FzzanSaxJJ8PyaU1HMRsCF3v4UIhi2VvbA
cd/PCgvtB+kXV/z47JJTUjh8UzBA3JbYASPvFZphy0W3+7aFWjnIPrka+pTr83QM
fKmTmSvY+YYSEm34XM3q9qPSbf1zXVlnbZCh/fnaaPkcGrP3ANsO78RTAnTAl0Ys
4R6gdH3Sr4lG6OfbUE8+UAoYoPQ6LNYS2GixhP9nbDQr558YDsU8XhVlhvEiIz2F
dmUBw0fzWM2zAFQmWvpjbqRq8PJy0FRffnn17Ee7cs4SJvgk5/hxr1DOVx/cIZxd
TCIqDBQfRymNd89ENAKrLMUOyNaX93tawfTn8ZqJ3un6fX6tPmwbPFNwV6lDHC9w
rEZ4IjxWie1AcLZfp8kZ+I0Sz/UUBjjjJt8g/M10rqA7OPdjTY74valpMt9trXol
fT/1xnHYcdHPrDivmHlD9DNR1kOjPDi949MNcj4wOiRDPjz06O5gENJF7Duwl5e3
dazonmMsh31upEVGgU/9moro7H/us6HoCHQ4oAw88NX/ObMq+ECNSy03ybW5erVb
yhmHe4CuBmYT4UjNQJ75wwTrPayxciJCrsvcz9mQX0vz1iao0P+aIz1+MVy3g23k
abIKBBJ/YsWbHziwJwsVVrq8AGYvV3fBfq0O0dOL6aqhBzWSbN4TcFjGrMDqpS0X
FFoy6yp8hu8YQmw6FEuczr2WGJ6E+kpLaVNRP0UXynBtsvBn+ofnXxYndoWNx/3F
62mCTFcVYumYJQb9RYZCstXr+XHkiXWteGFx8FzkwfUA0lFMwH0+8fWiSHgzhq/y
zVavzvU+VwDmEQdsieoVO1Qt/RHAc5HwYcsC9QS7up7gYrlHiUJmYApQmqP8i5U4
gD3Zv9/DbkTMJ5flJ9QICE7SiRPeXwhrKhyWGZFRC4xWuCjkieblqu+PG/Tv+QRP
v5icp/LyfrkWutpIfOIDFYc8OtMecSkbr4F+feEIViPHoj1u+0tFTQYOZz9PMnpJ
6IVE0sKHkS0OuSTL+8BlZ5AiLFS3YRGlUqu7VqPalrqcox38VdmePGX/uP+MsFcz
ZYMFjQdpNHkgrBBAzr9kz+Ko6nSAfHVCWlWbVT0g9CgX7VDioUYWHlBkmSP6sUT1
Pn/xjHf4DrE4isujuZKIRM9AbFAzU8pt+iJ72tQ4mWFL2HcmoZ09KF9z3IsxglqM
bfLn0zyi/sXDvasi8VfarqYsnk6uo1FWBh6DvZ7VRFJT+A4VNBZ9NHsD8LleeqDs
ASbywwQxLuMFo/48Me3PRe/88RqkZCpPU0g0YVWX/7mZ5hgcLMAyrBq62i5mi7ZJ
uGtv3i1facJtIocuRFrRaBp42Eexr3/IXBQDTnHl1UTsXHQtm5DRwADzHWK90syi
149WaiM+DfqUvHuG1Rnrt9iyw1tNb+0Ld0zfMcFL6mb3s4Y2NGwdBCtiiLdijjIF
rS+lGv3NFN8B2VR/hA9ePX8wRSvmbmkk4VXRb3C9RwnuvCunJE1mhhNGhNaICeEA
Rcq5Q4UCbpSYRJA3Jv+hc8fy4WfoEYDL3rRnLKoC04T6tiOyVfa4Id8OWXuE4deo
dZkG7rlsZhc00SsjOriKtMSEDdhUUnNHVeaOiUqfW7kGRea5NGTV/7wQDukFimSt
bKtw7XKDB2n48+vr3Iv647enP1FjmYq7kdYcH9y0q2LjaDYDxPnfs3AJTgHOKx93
VzBle2Hk83NGpTEb581yC/74MDOHaqg0YxeB/gs04WJBs0M4g00vuwrMJvqOcAq8
Erl+U/jnPTbeC/AYmUJwcUvjgB1nOW9KqkMj6p3DS2dusQv9nVfx0pDS64WOAFUZ
6qxE+ADaXkuV/wxtSBUkF4uBWjEcWInM/D51hx99YF2/dyDd+nFaRMZbOA31VFF9
IeZx3t8U8ju029PgKdVLDUL1y+ATrsdYr47LIIN9EqDqPh1pFzt5nkrd5GmEEsqA
U0LE1GeDihG00onyI0T81j97WiP9I9FK0dDGrBwsPp72HeY/U8iZc5D44eXcbjN/
1TOz+u55he94439elWjCUA1nQb3+OgtU1zMSHCdCGoDU2p8vMzVAD49ySsCM7e6z
aEfhMYmwONChvubxgbv0F+R8nbrpq++4Ln/pQFArjfnd3c1BGghFIoxs+1NLTHHz
IHVSU5EqAIUg9eGFYEGtoK3Lu0vqmXLJUuoog3Lqu2rvhjDpJRQuxydKC5Ur5oDl
57IjZIq7neYdkK/MZknDWnwZiYTT8xreMOAxEFzr3ZiEDxJtR/w67cbD4riSGWpm
lR7tmRTp4pYAd2HqVSKLoARwrqUtN5zX+WtpCDSHENn+nBmA6d+tbVQvBNe28bMc
Nw7gkFvDdQOa0XlekaX8OfCYVmYFd325XAhEn2xabUs7X/ViFY0nx6x7mgCE4QVe
kDQukZVsX8mhID4NK9CxS67LjviICItPvTTnOiUk5qkKNVCbWlDaPQyiyYksuO+i
5u3FiySV+Nc5lS3eLnlovHwbMFVp0kS3EEGLrBlFHLJC6bQzOr4yKigmS5Pgz9VT
Q9jUiFmeiI52KCBnsz5Wcbf4fVZiuDCL5vpjc40o4TXHsocaKF9vT2rl7jNaI76r
E0+OQdlCUydkSJpkTgLn35Jb3P6cI6E/rvXmAdR8ZaLFw34Mu07SBhOyBYpFSBZZ
vwWhd84xboBoVLDxV7Ua/OBj8ZBQXME2AaRdAuP5dxayS8vw2tZ/IrtgdYgzy1so
M5XVGku6OC1iAXrj9MSNEhkDH+UFvZK3mVN6WUf6BPFVmlAewZNXRObP7MHqLfWt
uXgV3Y6A7c3LHzXoJKCXH54GVN0VmASB8zNQZ74UhtNo54BkYi663J3GYm+7ON3Y
IWczwr16jiJtZQSRex16nSpcS2JHiN1MG0glEhBN5VYonBy0FQgD44uh6r/3+Zth
Hm4HcKQ6T+TtVV5aQDXb8/5ExtH8jbJ+ETesiQ7PDqnyDY8hSBclAOkeGnolCIrt
O6hgGEyjn89UbiF1MgQ5PGPGMhr1gYzJQYqj3+ZIWAJUT+74YdnqwyS4iRxqH2Ft
HqAqNrnQVOlcODnEGlJuYT2iMlDiyF5sUHMHpTHRlmZMd5vvF4yTGtBqKCBQWoDE
gqGlhCnnJEU3m/+4MfDN+PvQ/KRcU3mUCctmFNC2Ar5Bcc06nLc1UhdwNJIYWHqf
rjQBf8Y8OQHb0n/oL9bvZbKBDgqtwibFwNE9WXaHo9g6ea6vcLgKbchIua0UGQxz
8gVQZYzfg1CO+qxQReUfNGMWkxz2rve0Q94JVma1MXUkH+rCgDmMzCx6OCw878Ah
D6yNcRljSWTBx3Vd2Uxby14ECHLD4WIbogkZ49w7CoQTBM+7PQC2Y8mdA0384l4y
smo8CCntJFqf1VWhbqf8hmT61y4cTv1sTbVRZ4ROVGc31EQA0guirBuO1LfV6t9d
1G67O0TF3pV2lJlZLq4jzezLX0SBxlN4OvkGPLqIVHzfwtGSeEBYc5kps/zRB/KQ
SzD3lBHlLqr+Lx0D7givenoaY+4RuCntBELPVt9XyDWy+uabvzA4L5UN2qjZaT5E
urwJrvZ/ArKH6SFTbdo6Zu0vbsAslN4qnIG/YXN/LCUxM7Zt0cp1Frclajys9AFQ
FAh/RVEHprhpuExRtf6Hnvdkm8iHcY1mBRBGwpyFyCD8J6yfGQyn+F1ipT1kpe9P
ROjC3mKuufiHWrQPwaIdkmO+jYstV6UKWwBN0KpurMbGp9AbHhXyuHlGl3Hivu5K
r9R0zEHt1gYdLPsDOEXvjegkmztWkkKRjZZTpdqtRD1I8Yes3gORfjo4q4ce79I5
Fr8gd4Ckem18ZKNFGQf6O46WtIZq4A/pZpDPZgA2Pm/eVwa9+eRBuTqGkBoMk4l9
sDK1rOdlw/TQCGfO/bmW9oXf0WyrdOrL878itQwtKXpjigjmjwyupOKVZTSzRCNn
F80y8RwJQ3KLH5P/Js0jeGdlmSoejdFAQ7y3Kw1iBm6nEv6+dD/2jHJssNLNUm9u
Vxi0cZnD8BbiW9QwCnHCuGZiCNvJ8aXahbErRK+4im2WmBQHpsXTYEQ/9naA6FV5
B/POOqUX0BA4oogDtww178ZrGQC1BbihZBVHJj+kn2Lu/N9cRq7kV0/acEWybBH7
KLBSbq+sFFFahVA0b0hyb5sVmkxemJxl2zWuRJDYs0WjLvVee2ei1ILcBOOuK6n5
pvYC6KKk1sihnhexlNL6tvqY2zHoaAONaj9Ifga9JFf8dA3UY5qnkfGCfDInrAVN
i0DlgRY68YTb4H80uHaE1xZmFg8SrDENpnDxfR9KT2KUKoBemU67ISTu9NbtvpD+
ig6zpdeT8gBZdtVm8gTyXV2moteZskvUmLYMKHw87VFQXvgbpNpZRUzSaqqb0T85
Ni0+J6BPVkNmRfcVuI0U8mF/Ud+Debl2YcjJlIIXDc7D2PjViql1Eeu5rYiK+SKw
E/dJeU0lp4oOwHq03U2oN1xQTYskEm5XZpqBVMUlOAt5BlJu98OMKC7vXVOfX3z/
L0XjeejBmpce/YUZo7APkaY0NM2QGFXyD198fTDX31G4ZF8JVIl2vHWnhMpyINuy
9S73ykqDTR6YgFiV/8IPU0R1mS2BhHvFSeeJ0bJfSjhYz6dN3J4s/GvPOzLX46oL
ixTyiOKlR4UQ2elbw/hQNtU6uuyvRMRsneu+ed7zKYPXlo2XQVzUoql6RGFkNHPP
H7epVM3x3xt+hCJnx2hs9WE8Kw5gNsYJXipaA0zCF37OP+YDxgH+2EG3Z4jz20Ph
RktbeY+D4FkQHT4eSGBIhwV7zdKA6PJDARQGnKmsQdXqDbUzA2aebji2Avfw/eYs
J9pIcM5Hmv+Du7FoFvZkFuz1+Zr/ln053inToUPH0C3ZO1BJryPyp2O7Xtwa02M/
pupLpOZStBflz04FskCq/I3KJSFjJ5ji4KlHrEr9V3CZEsSCvL8cNBq8H8J0bKtL
flPOpYJAJtL9CRGWpYJhMXITQJbKfQXCtPwkWw3TXxSisl7rWLG4caxeDgsQwZ7E
SjkPd37IHGifbnbA//dvaZxSU+Puy9rtblTQtZ1ZFXNbRGX8+M7zdPQigzGJnS1o
faDefm7nP8Y53gg1i/Pq3oFom6XnUzZjegm000fVI85qwyzFeGzAcF3IH00d/x8E
LcgL/k89++xVQcYVWEVsKrBMG1ADYkuT6lk4pAvauS/+63KKCYXkfupYm/KV/rCS
MI7snNZTWQFfrgzH3JSfWBCIvU4TesbDzgna8zfloRKTRoDK5vnjzy9qpoxvI8/8
XUl1ST/p58XjrrTpkZmjNYPH8DZjrLZdkhtf8Ou+J/4RjhLBkPpG88ScnWN46UFP
jzlcFFTusmS5ZXNBz4rGVGcA9olA/N93KmO6lVDCwYSyoJ9oG9LzvxB/iZmNqBnZ
HS+akBnnTBkouWG0pRkDNxVLL9rHQ5ud00zCUcF8fHJbg+IkE/WI2ui1m4bOBo+V
rma8wuFxe50ClebmMDpS2qFnwgcxaUD3o5/HnMZUNyPtU3CyPfvcvuss45D3p2yw
pKl/g0dTpCSH189g7NQwimy50K0XRLVXYawZ/X5DqNjreIWLsa9bFkTSgPGbQwQZ
/B4GieFaHUxmLlHRKvWLyMHzS2kQCiWYZ4tlLXEmWgNrJqGxZhjUgDs/M+qosEaf
DgPPZAH3A8wfax+rdN0YEGRiqfCAG7NmHpeECQ5uMUuyg4i1R/0I5eWuqFrdWmCy
ZxQDrxJiRI1riv17U2Lhsr/F35of8PJVX5vrMmh5blom5G3XLbZGIiWudqUJDyTf
lCu/GDlcyanDKiv2a1cVPcgVBMuW1V94CgnjEGQJqxQH+T/dQLHQLHIEI+t071va
SgnO1ldvvy1qSgAveAK5ps+Ce+F/mb/r8BUE+uQB0NTFbCWAPE9ARiguVTJSJ+Hw
irDQwF1DaXQah/U11ky1uFtQWsGo1X9JqiASZGpLy7RhijTzgNZSwbrK2o4phU7b
mCOIB68fTVoSiUH5N8tHnj0VI8I/eGOODwK/21zidZ1oKZQzQp/Nhq7NafdoP8bN
JH0jUwhefsHUSUS+IfLainIb/hxUYLQpg62UCjGxLBiPrDwWA1+7wcREIinfYn/r
+q/Yhqlb2vQgvSqaBQgPdcW6f+DBavoIYfUUeM3rgwpoKpWCo5QfsFrol7iYweI6
SGEMa3D9SI85ieR1IknVhCyUV1d+90/7BY1f+Lwp17ugF9PQXRDO5RV7xUXnwTLf
oZnWD5spVpQIkpua+lWiO7ltGAV09GxF0HBUb/RcPRPijwTPL9Iy9ljyari01r2D
wwdoX/7T/OF7refqtZ0SOVAcVnDJb4wzrTgiV2gDomq+rJcWEe4sfqIOM3fyWtEm
GPx05N0TSLSaEMN9ir75zhpvwdpo4CBoIHve7M0MDWyl6rhKScUpFK9jqyVtpdS+
4a9bItKhWr/lbykU3JYFxHDu5r6aK95Xs2FeVkVrVLVCjn1mhFyAnI3PdFoi6fOG
w2wJv0uPEtKJVAvJsJF2I0G+fPNV2O4CxVGOmIyBrTbZEoiy6OflSulnxTdxCSpM
QRzxwSzktthwdm+AH12tlYxYmGCTBPVKsMhYS+LFZwg+sShZAErsSQxtgozXDoUl
mXMr7wTVRNuJOvxEvQfMKgqw9/LcGmouZjJaukU5d5R4W6YEnGscHWOzkvwOALNN
HJJEDksQrZXOEFz76dJACO4+iPgAlTWIFqIcZk9MeC0Bx41XaIlJLg3SWqHGHGL3
wofIpwRLKbuYtyKEESjJuDsJHNYfcMC1zSgZJXAIAhBMQD2nQxTRjzPNlFBlfsSJ
B0K+Ql0IT6XofnhJO9U0OA6WunGchfuaFsD2QkTUU+yzA7B03LXc9MO/MvbUqbQC
j+udAKEl2DOKbEu7DUiicf5sz5hqT3+ggPC2LNSVMUf/kfSRq4PSDoKsLwXvcXkA
wbKNjWhd8fSLm5GjJJsKQsWH1y/yEnWKZeZu3Lml99KE6A3LdeV1+yLHltDE+Q++
P0bzrzbSdnyaXKLdRZ1Unnxnt7sT8VVmHWrA+pC6i/r03VorvEYN5knMmykA0vqH
5JSHdcQSsOM5zxEg9DSGpdQoFS0moubPx01Cb+Sxa6JXjxr62Ls6nV+MdHVSCKmC
C7Q8oY/Le1XU6lUho33r/+VFDd8Vnxu3VtPCg9SGx7gbQQiPojv4q2AVOeu1gffo
m16eZPFLQzAR6BdsxW5ZIZz2sf5XAlN4lO7lktxynJsBUEH6sO4zfJS5dn7KrkSw
vesJ2g0cLcKNDefTU6w+EOA8nHbPpqtybdxTqQX/+ytSwu7QrePzqD1dD51p26ig
v9m6Wily8ptGCwAXReEYJK37C5DJ4teKaXh6HhDmN3BfrdbnazGyH0ANd8D6toZw
+xA9SQbF4aeXLXssMaAmYLdSJN9eURrXe8YsyMS33oy5fNX60aaNtnxzZcWUbnwl
rcDIDmBJ61Oi6Q/xg84a9AUeOy54Ned5VUF97Or5ar7MAuRAhm4DXKlchf7Q+d+O
mX4HuhV/hXv39+DpBTsMdjgvfe/LvB4rRO9yGcCAGF3WC7VM/cYkFhdWhwVLwv8F
Zao30hU3lKKOLQd6FXONyybzWMzoUKuiFTfXge+hH5ynXMIqxi4SElvowx9saMjZ
Cbsb+mEbxN0mLkAGUrYn2AF6h130Bl2CAeBKewsnNZWDVDF6FowwMqLsZRwKwNW6
wSRpJ1M3t33m8oYSjiDk65lMxRBXvhyLJJpYWIn2R6VmmCBZR7qs+jUEcSmoN++x
o02n0jypLlUG5PGrxV0hhKXnQYwtVPT6bNWFQK3Qu+kD9qpNXSLewM5NIo3no+Q7
KNHkSKGCKQti4VHY6ONWzeC0kdbbeLu06ohn9w4Yoi2z8e3mAsvMiG2gTWS8ZknA
bj9btYub/wpGKNLHtd6yYs4erqREaJtaFst6FpsUOAORi1tPzahJ6aRkvz31jb+H
OZNI0LFtrAmq9cVNL+B6Qfpr6inQ9F8n0dti8UK6atGuIzGqZvPOpIScU//7HzeD
Vmk93NR3ES0EFyxFLuXLGkvpe6Do2h4e4khv4ln+xO9IivKC+Xb4zCiukjz30F+U
eON0lKoeaa4ZIIvdSco8x730skOo/V8XPLNuw30yvWobIseQaR2WfjqYTJ5rUDlf
HUt97T5vCNbUW78Kmf1edHwAJQ8IpupF0qQJGZO1IJsebcsUf2+bgFt6UnSezJ0E
hGREVeFX80iuVHX+HH8fF+KfupSxPpwmYtlY6N2+HCqLx3gUC60KJDfYajdZiXIT
+DktVW+hFfdnTg19gMRaDjgScXsYILFf3qiXnpRHHjGwXANE0d5yli/bgtS/SVSc
24EPwFa9RUQXhneBkbJC3MUFUQVFMm9N6/XXUA4lqgzMolHRasbNzOnimxPpJeQ6
Lw3Z8YAy5tlCeU6mbbXnzdBa8AH5LuYVuEYR+xTdnHgy7vbwpoa1zQ0Lk2zZIin1
d1PKvPNWbFf71FuO/CstMCLgG3gtX9zi5Urn2MSbHFfrH5UFoPMzJz5h79U8wwcj
9UyTXtFlN7YpAhIkItU1PQ5peTO4qLKRUNTKrbnye59/AqDUFqKupl2tiC40Vu7s
Ty4zviljgSOb4q/KQSSTg8UOwYhE7onfxiQbr/OmuCrFCHOpnoR7n/3HIGTM4z5g
QJePvg1OyTrmBpZytDMvamUhjVb9eYqi6xKPJoIE5JZ0ffs0li/n2mlN+7Lg656k
XGs2pPF5xgoAG9Q0HxSDtzoB0nkqcPfB0vr3FjE5Dbq/c5jxpenRLYRv6i/3aN2C
RqQLZwzBjw5cxMJIQKxDesU9IIthj4asXrJxV1k+7sEbI095t69xwomhDEL3Ej7L
1pOSYKVpBAMssqp1d2nuvQWF9OiNQ8EL2TWAbeG86FrGPqDKU/xdE4HRusK+l7HE
dQ6OjKUNlDIFLkbgyPOlueHyr/5xzwTMmlfRKHHi+e9N3Cp2r3R/S/w2qV9grKX9
emxT/BQWwULF8FcbhZbAUJlsB+Vg6Hzmtsm3qiCwFfQziDnY0zlFEQmBQRICRlqD
9DBLb+R/exXeQzq13xC9RVtZNC4b89illfl2C6yMQP5ntV5zN+2HKKQ/wTdvmlvY
OqED6v/MqQ1fShuEat/WUUmjK8P/IHPI361oJQ0i7jtwl1RTaA8GvbZ6/x9+7vMx
0BZ++N7Ok9nZQFzPkKzSXr7fJ+GnomiHkUeqcNgfz5a8I+bHWS/Mg9YMzyWwmGN/
WoH31evAAJy3PvAMPuVu8dqBrdYfQiRLZ71I/fsew4M+ArT4tqmVlR7E58Ov45YA
p//24aOS4qCWschP5obOl8T29tUpCTW+nfGGDyRn5fTrrWMXVLWTuPJlpc/n65vW
CDWwRH2uR+tDv9Jo0uhiXXWiDEnBxtjl/U8jfP6nqsxnowuDNUsSK0cO5uMkvSWd
RiAPQPz3pNXNn8N7Ee0WMnkUdtTgIbd+puBu9DeJhnNOjnsGIbF9ZBaexH47CNAc
rvYCC6UzWltxofNkswPBu26m6XycC6qmZ4Kx30UWLhaq79ajCy90cVbR6WkiUal4
UqEYZGqnXC787FHlDGQhxQaefIIODT0GO1B628tMWgyyiywdmQ8OHgCOp8YpBVpf
FAlsKc+bYJWKDmyIx1BiSMWoFCsy9ocsM0HDWbyUer8QzBJ1BkLzfMaRLwD8yY10
UMkrtAnprnNfJ36p9lUl/SiMavTVGDe1fymf5/uCMgQJ4ZR+b0PYeEuLb62vMBek
gtURJ70z0cDZiuxnuxwUnXU86GwwgbB46osJdmtFqFgkaegFVZNxIw2AsmnW/1P+
yM6t8OQJoq4skCmVP9bpwsxnRjjfRw5Er/QXMAOoRcid6jFtJsMfro/kiqbXYtmA
xjOCJYMXJ0Qz6sAxGKiF5TiVNw36KzXXxRmD7F3khOwp6YBRZY3jJaq+NvO1RRMv
8K8WcIWfNG9tJyXFyzGqEj/Mk8bPufRZjQUlHG7+Q1k7MN3htVdvyouwakU1RCiN
ajyCebWG0Z6Z/bea2/Zxr2/Xjg8zgj5IpobWm3JhRsKS3kgBpmMNW8FJjXcf/ChN
iXvn1tsSVqUqOJPj2fyPBOwu5KRm93Tki4s5sPbrIVKtrzY2SUQnuVVjzyI30DUM
SM0q3h+3y+RMU/+Tu4hzcoRexMgYcL8rt19Pda1bIlH6mkgxLjEtOJ3d/qqI3y38
Q+Wx0GG599/gsLui1EW2KzUF4hO7bCk6Ujg9zetZNNVjamwxtLbUMsu9czKPpQSQ
LCTIuNUdfxeEDklBadnFpYidzPnQMdTXw+AJ1cFoeqnkDvdecDF+XPP7SANkGhB7
IdTTcUVMGvCuTqaDyyU/bAm06agRjQniZKce8t1il1p9nm8l8RYjw7XZC/z+GQ68
VoW1B6Ejx1lV+3dMniaqD197zsX8WRuTUiVmvJZWHrff0EON5IXljufqA3Wk15kv
3Cw1xCQNTT8QnaPaTiEW4e8YPdTWKtsuZ7kPHh1FtutDYNNfXneRa5fLXdp9+o9g
P2o+//6p4iLUDdPlbVO88bIJebjYTQKZtfc8vPwuo7id07UYke6VYZhZVDmI1/k7
nxA1ZJzOnQ92ATMjRWrGDY+gwCT2i9iPeWzASlIzdRQEFm9d8Mh5HDgw6cVgl0QJ
w7/7Y30I9pZIWd/gnrZcNIUF+SOOVo7vvWmZT4wDpAT/4jZmAk/YJgkFJVsBQwh+
IAVDxrm5PL9utvTGKm5nPvZIqtFi5JD9UFTxqNT7bstdHCYQokdBHCQED4c/ghsm
7WAAOIex2Kxzr18wcSbq6fsxroHzWk9JuA2FOTMkNmB2NZ1CdMzl0AKz2GBCM7NX
kws1zz26q+SJMshvCjUXQOzy2QrhQYA3hlxcgExrVaZEnZxBq/Qk9hDwQJkjVJ3J
hoBbMgTMj5A61W0APOr5Se8iYvQiA6ks1fXBRoHaDqpZffyPSgPFwWzFZm2zDGCB
0huFjRgee3IJzSI4Q48HhJ9WwdSYQt0GetWMvazeHj/YAeLuU820F9MvvucSSHYe
Gla+uAvdtit6dPcoQPjNkaQVc9KuB4wEMKZsVtedD5yw7/duXCne8IAYpoxON9SY
W3ZYW9RxG/sPrWy0jKYrwso4WLfsUcyVvOWPCI4JVbMI/c4YTzlLp63KrvK5g07+
oNDnxjDXzEJ9vkJ+WGF0pVaWIwiv6F2GEiWMvuVu6UPtl9ohEOz9d/gyaAlMOL7/
XF6WKLqCpQUcClVpfmpxBYjmflqc8kjkgHrgOlAiOzdYXm6vB+m0kf9q31nFeFoP
xw1yL8FUZAqB6VURQNg6MCpRi81eN4M8psciUWYNsHO2/XAYtfB3DdLfGieN6ZVm
7iSlo2BqQnN8q68nFYXIkKGDXNSJIIumQFM9DSczt+hNdMF4cj7jeV4esADl3mL8
Rc9a2Wj4WOL4xfVAWjFxVqCakES9zSuGjKN/HSYWU7TMpDxy8CI76HOQyURwG2pr
S2ptsqXUa+93plFN5SlsX3QGI1HkpJ28zdu3aC8Ml0iXwzqkdoZ5Fr1dvP+iPYPs
hOPkMamP/Moay+4kvbqlXYjhKQQ2zqAVg6qVWt43qz1plkpzEyjoASABE7yuMWT1
btiq0Ga4ywW8TRGsXm60Uw==
`protect END_PROTECTED
