`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Atg+HljrcRm4NNPwTOx/a19eMryWlUsOK6TiUyAndPtFBug+U+XoZGk3Dp1t/Xb
KF+h2R5Uyk4cQ2WlFAOPkgx3+ZwK3b2Lsgoh968lX9z09VK30XBWiEqTvaCIVQZ+
nqlqK5Ia52oGDmiSdGhKwMiZK8UiTQSjayjGiLeJN8Tder7L8qlZJc5ka7woAyRQ
utuGHeJd75VPv3R82RP1w+g/x93jAfKb8XAhez0tTaM/rC2XkNrXRdYxI7nnU5R2
/mEnWNwMp9cIM+1+EEWLs39/CG0G/KhsmnQQMV7ePmHtz7EMJKoFT6IKM3TakQb2
GvSJmaqZ8RBrXKST7QfPRW4Qs9MgBY5c90L3ePqbI4/kwWKO6zNVYd9/we90L1qi
aiFFx92c9c5V7cT/vRZ9eg==
`protect END_PROTECTED
