`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLbe9s90uIv9c6RDNyK1uIX+PI0CvU3TYH/Khi+vTqYJCMuaJVraHy7H4YWjrky7
t3bdOw8eVVvydDrHPlOwTN3yhSnAVQrKu4PppTNAFjoVVWiTHKQsGNO5+xGvFUvs
CMtrsp4BhAwh6YtHdlWXXQkKYVZmA10LBYuQlbUX9/ZW9sTepNbUuhKf1EHn7gZ9
s3U1mSgpmzTLUxOOhjWqWkRZdsNN878dsMBWIodFpdYglyxc+F2fncHStaWLz17n
ezSXaLNEoucjqYJDRQ3GJLYnWB1npeEEV4e+4ZVv/YKwB7GkYSI9e1/4uWUzF8lr
+E3ig2JG05mZwNHRqe3Ni+9zjW027d7je03VhgwBMBGqPUe13Dcm65l9g723g6sb
B0GPMMeiWBydZPSIOxaCZKb0f71OaRBB1dLj9wx1EVz6l2S620dJUN503qSXgaaW
k3d52bLs90wvVa2tLY1WcBEYs1JPcMfT3OVIG9B4HFFRhlV0SllXuz5jV9mExBiy
5ZSsF9AIY6VgFvOdDNyw+EtAncHgALIW0zmogUF6kYBa/YQdoR0EKYTayN40QW6Z
8US4EybB+ylA0RnGAV6giw==
`protect END_PROTECTED
