`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QL74ghthb+SGsjFVu/RLiwNDFWHtA4R2Z7KtWVqNos2BlAd6wKwpxsURaUxRyAfU
kIJHUKt2J4qpcQjYtKLFGOFd2GPbkcBzSRA+gq2MnGQPCsXWaACFhV1evvpCNI1f
r5BCROF5JGUpNWDWmba2w56UBNZXrk0qtNKcPqgAmqSHHBdld9y6dedqV+iVhbw4
6aB8T5IUoqfaA3P+9k8nD2wqs/WlevFhDiwzaeRdiXVHupCG1BWg4GIatbfgWTqe
EySc59xB1dxWk4JYsyMn5hYUj6W39gxekVkn8ToUG1abirtNw7P4Xbv/VdNHSZwV
8NeS/y+L1GL4rusZB8l/z7Y3NGMVHlP0CBsltpI1jNdpoU9syEXjh4Z3hocX1ouf
eevdwtQzMbgjVhlC3FnyhLHAFLoC2gb3Zv2KMR93wucrNd5YJy1MYuMNGIEe+C4B
ISqGv1aB5apXcXXNtYcYi/VJyU7N7dFhZUs9PB/9ujkqNhPRAv9H/ZMIIcMOwalE
byU5nTk4xx2ldLuUuRDOghNyXakX7waoD2IpSuCkDVWRiaWTb1JCL8K7FfsKRm6k
ym8ayCVoZ0mmRNcT+IpRpsHX16hU8jAM2eigLD9lMC4kU6SImbWLMgF96sDjrE+F
YulhoccR2FxemwfTFG3UgX1bBVgNUTCX8j9VkvXqHI7gkdqOOcENUX+EWy10drZZ
m+53ABYbNPZFStnIBEFNIzADEMykPHznh21AS1YNqph6UMuUJMTIkwK9RaCa4ChU
COCedtZGOMJNeGrPhgqVvtHpw9hhDktZzdd9cclab0/dhC9L9PzOd3UsS9FJrWQo
Msu9p0jaDdme1V26JQgb383B2qbzDBEgaY2o34o69juaTFgVutGjIycasjYhyUKF
UeIowzu25pbwFmxKzlRO40RHfKW165r5hMVbyEuZUFC/Hv5AptoOBRqKj944/RFF
I+1vr+bPfd/E8tDpzg3UaS2l+Bu/bKTHlGyqZEmkQrua/ENbZ3qAGtMTm3qxIpNW
puPS8RW+la6ZZKrpW/FRu94idvDx+j9UFzB2K6Ebz3hERQrZA7YPn8LMPz579HSX
/V7r7ijk5I1qrlp0B3iinD5Z4eWzHoGoTWa9hMOLATy9FzCQpWGmdkGcmlS2v/rb
wDdpqg838O7yp13THHfRivIKkJ+KgIZDeHukaypACfzESVwULO6BGt8WgOtwoEeK
1AuJ0LTWpj66j0VcwkZKkLa370JouG/qjd5zuDEqp8+tsrLYh/Eer7dGaRlkid9b
N3vGwfCBTI+fu8fXXAnLyLzOnapapSXsoJozX8H4x7+two6b08z+XIVfxPp/kJ0o
19dkip62Im2ySRt4gOFsH5PHBulPoGAHsYayD1rTEh7HD+5CDn9Ghox6V2yrxF0S
DIU9hBckpQm8bD+1Uh0ooX0wc76vnD1+zlT/C+MXoaGRM9gxPdgHrQOMdnahF4xU
/BVzrn041ALp8YT7rq389E0FCZRDwr0pSvbwEgAsXdX0yj7F9/ugUlTamBikn+sZ
06mESu79KKf7Q2wzi8X2oTBH7wftPTyNE/gcOkduAo6Nje+2NFJu0pSzbALAG+45
/p56lwJt9Lbl+fgxhcwi2+zhurzKLrNThztAU2yhh1kAnp2Tlj1Jj4NUUDuaKTqu
VKTtS2DRlKh4jChhQbm0bM3VUWd8Mm1KyLULNTCLAo+U3R+kE+65qxgbTR902cTz
a6NXJnZjj2+oWJOPFSbg5z3nezgip1U2HtZvYw/kOobaQ+5ezf+NhOj2Zj9pXCKW
Ym0HOGK13B4vl10xnT1h0AJ/6vQtz249YHbzBVxv1RRVWQEnCeAz2sGdGFPLpxFR
ONwkBECTH/HMJnpBAi/R6SGPVuoZGJsmwcglrK8qTwQf2CqF4yMkBRburoYjY8/o
Q3A7oOPmclZnYrhlqFKji9awwYgHrJkkF8Hs5x0jVLXkrwy72d7gqUisD3HNF2cM
pGZqWXTO4hTxxcQmQm+/pIYSA2evbyEtDsNorLSMKWdFUJl4g5sSE5QVMp8KCZAJ
5qBP2NImwqzBgiSmIs7Bh2OfQv2Ts6E/KyO4y6tDwZCeWnCBsZxnvHLXb3QprjtL
0lNgmUAi85tZcLWFGPVkYk9TE2u9f1GsgmPMesF0OBF/tddnPe7IBMDlkn2pzoqm
Y9bPkm8vwMO2Ur6AnLK1E1aCv7KOx/CiB9e01rroi4SEuNqMsUtH8MRxKAFZaE/Z
4ynfbXqgJU2FecPPuwTpJGgr30Iq8WfiV+MRxpI4jE/qWsyLcFTvwovJGF96y3Dg
1jzx9dH8bM5euYGC2nkeFJ/boG6CJ4Hb1Hl6evDJmF7853v88oAA54704X1Pbspj
xBxVYQ9m6L/9Ooq+MvYYTIV+Y5+JCYxHzwbEkNORPs8AwzQGUESIDXKinKQJvSSY
dv1kM0Tj5F6Tf9bn+87aTiELAikxRYzrDRjEYoZxzFdPhZl3gJ0ohVXSdOMYM6VM
URrIEqXoIfBSpaethfha75TlxvGgXbNS5EqHq2Zq7A2ztsGh8aW2ZcDwbKD+9LsA
CJVeiPE1jOu4VK3o9xNO07V3VhhcscIEjZpzCD+xHCAY20P18ynOVMbXgjrDeVBW
s3Geu+5tKv7ktpGeOS+8WHBtDU0GnIdrPS/9jZ31TAL6ua1JxLxlgmankJW48d15
jWJlBkbew8K7YCffUD80KBGrf2EEf9GCv7bahWeMQtr5YL6NUygEydpwG9O/FIHt
ks0A7VuixupyNvTI1EqndN5LfJuMVQp3i91kpb4FlzrCWChMqu2pkxpvipK7pkKk
z2cKckaDHHf+RT3NABaYKDDR8jxXkro07KzCQK3KZdlVTyAisO3OBGkZAf975UrA
y2tkNBixnJDZFxyHjYUI7Zd1Md6/H0ijhAGvbEcNUuyvk7MWLPh/5vP3YSCFee68
JMhHd3ed4OJ7zMPPDFsvJozdINNieko73EIzNbc6Tp5NWhpOJbrO+4vUrvu5XTwe
+rVAgFMaU4XADTqME4qoh58VEC6EDicPwo0acmsIYzCt3oamNqQpOMNGThyc/tzo
bMzPAmrjfTOpCl3O3LWO5oD4iONGqnlJgTXk7oBQeejkT1HJbtLvIbnoIQgy6TD9
ejPWpjV6kBp1VrwRUdZ4G0cne1SynZfHbRxRt2ZCxR88alBEQW3/kk0ivXL8yxxE
XL79Fm6OAjvwlPcvlftfn1FW5YQcbzyOTwfAVzATn95R4CxBgxKTW8zhd4s10ZkZ
ixvWmBicDmJ2qZ7CjPiu8ENu+xHYuK7KKR/7NTekgyaRTfcbqpVMfITFkWPnIntj
6FPAnm/PpZFgLg2l9gK/7bgjX8IRe09MI5ORMKGqBfA=
`protect END_PROTECTED
