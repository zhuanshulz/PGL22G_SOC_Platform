`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJRmLassU2z8I86WnFpcvtfRozW6BKPzPt4rw/8mLxTAyCM7RVauyxsvpKIRm/S0
M8uLXBZEhM3IROWOi1cpv0tOlg4/V1qXyg5nlI2hMOOzM7QXsMszvpiAOMUwfg0A
SRNKGidI6TmrwY+cubBe7xEt/T8vQrfI9bJ/sKGxWgDU41KFjjR6yoZMA6XJjoh4
iwfJcDV4Dnt/qDW4h+2R4PXRi7mYms2y7m6HiLV8O3frSVuGMvWMlGIv8WFs8PBG
88fNaOP616f57vlRkVVbKAihO9gq7gMW+l3nIG6G4UUD+8UytRiKHgWphGyPIb3G
9R6JjmPjZManVuU6EKS5EUWyPjy9HCDbxU1k53CAXrTYg6MepTG/FHidREf1Zdn3
Oosvg3VJ+ojcULLO3s2FqZYvdW4YJU0UxiEprhDKa86QPf4e/GelDRjsdwKOGplW
iJxlIFZUqVpD0iE0CL8O9D0ozmsZ+JHvW7KPpY1F6Ik2sSXCZq1sg2EYc/aPu0g6
AAHNd+hrhSyUyHT3Cvt2vFGUUgua5jGIJfqnhEJJ/T4kutF++bN9XGpi0qLgdklt
3MxADyAcXwJC5Yj9Lrc+UcVneXZRPyXenibbVqwDvMtih7MoOKjarwIwrCn/0kGu
czYf4fLdFkX0VNCf3WY4siTSu+qqv8d6wgpf5NCZa/HqHjsb2z598t8TiEXaU9th
WszeEe4zWP1pp/6jZts1fuLsfWjcgsQChijb8rejszwjozaVEoltAXHbpFdkw89+
0t3ZTtlJg57dDbOBFbRHrN7oCgwr04LUjSMDL/IqvNqGuq6lXYz9riYxD+aA4dJg
KmJEthunZtscWHEoFaG/Fd9Js9B0dKolfsp8x+3Jtxlc2XpjUP0cPAL/7H7TILfU
/yfSevg/dKtRKiDjLBsJrYfwF6jPdgJPGUgqiIj6arK3XYWoq6AylEhyFw6ENhGC
qpxtXKik9AjTMZZFE9iNiHnbf0lLVLKdsz9CkoPAJsABIRM7h+Pc9aEeD+HPmw8R
xDIR0YojOdSyLYQaS9OYpvvHlyMkNbuaJ6wXs/66HZdPlQ3Bs4AXLr3ytPUln2MW
OK+h43EbhxJ9F5gTU1OGUpCTbNn74pBLV2uspmlD/heYmqBjXYEHgcKfprN4uK7g
bv6q3n+kjmC9L6zC/U9pd4JAhZ9gDDzh/9Fq+B4PYK+obzZmKCjPGZvEL+NxnXd0
1THRD7Gb7ObEd4EFIAnI5t6M+mUCtW/adykx1edPMQiLLnJAm4bpBBG8Rc8ERoEf
y+BBKUEU+5tGqCDaAdoqVB1EIZUYdU5CU0QcbHqLHfxoaBa068DopwyhgNNQQDmd
`protect END_PROTECTED
