`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uNogR79PbmtEPc8SH9nwExE9JnNw8/qCUb2yAesDjKWiqdcjPH89fwobo251n5Qw
zmOettn6jIXcwW9sEbP15CwJI9UBsvJTGxs9FxATUvuC0Z56ULLHOY5yZTId8IHN
hmjBzxf54H8g2t2RD2AHCnWhgDy86OWRpFMYfM6q+ovD/ONtyte3pG2z/CKLfKNg
OswHY5gTJjEQ51Km38Erhc8UisvhrAxI2ugBlcS+N6Gh4ZHG5StiCK3sLHjw8kf6
MjNOd2ad90uMgMp7pVmB6kJL+oD3KEAOqsQ+MdoTpmvzSaxehFT/b+2rMXpHUTa0
iTKpiqOP2j0xIj+MXhkRI7M9NEaUINLjsTNIateYBg2FxmVjiAUkLRGq4/h6+Pay
Lz5VEdhuGH1unwOpEWUD3AIrHpJIKCn6t5nUHAEI4G7bp8y486i+dGOQSoL/ldiU
UvraKB6kSb8pbjyk3sANZleqRM/nyWZ3Vy1uGudBlQXhd5n1a/F5kFF7z6QW3Ckl
tt2gwXSS1kM+wxRw0Av6hD1rGSItjq/jWDBo+hL0IZ/egVNAMQdR4GgRuc3sfktT
VpkHWgYp6JaYl31wIeUVWFTyRyrfn00ch1feMOZ9PjLYfUaLDI/zaVF11qxJpVvN
KtgN33nATCO0H33xza4fHpNW5fMVsbrMjSIEwZQMd09YI2I+2uMgx5wU6X8DAeUE
ePH8jvetXkgxvnCaU64jKDwOygGljSc7vT17vA6itRRpBLW74PhUx5UUt4ne11M3
MP6i+q7U9tXTRYBFnf/ZgZ6rD5MtI9kK0QFRamYdOXjvLHh5uHj4Me/GM3r/3Hgq
WlBwHaOeo8SBS3Acku3JhPOmHLv/5lQo0/E5wckZ/3Rx4l9b9wej/qVj72kP+LRA
KVyo8yuLXZnHCWAUcsT9woEkalVf+86xeRcp3rAAJXI=
`protect END_PROTECTED
