`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OVJ05dxDl72sa4M4BFzPTSLdXyavqerHkj4dRsqyKgJiodAZpAQkmHn7ye8lOC9X
ewSQJwKoSWeJC461PXJz1j9EihDgHZpQpdDT9woY2ql5ufpEHIVyTXKnY9lsuU5T
bGWHhTP83mtD9s0JMr9+pO2zRKbYjKRqiaBrz4fumkHSIF1OngQEAohuyvrafvXE
V654WSesLJ744TfsYnHsqNZpN9jkSnEFyZVZBBElCXF2ydd9di8J87UKWp9+n0Ua
Zag+yQ/4bTNirj6ea0IQ8ttbaRf27vXcMmDixDljvEI13GAOMfFP1MtzuQ4CDDgp
pvfLjZPvT+CxzhqJ9OGXJ2ZFvNms5seB45l0QhRyxJDE0IAXmjNioBhdh13x8Qg+
dzloRlLthyBs7KRPE3s66cqEoLbeJHTNq7GGb4qYJaf5GiOHFeSvQf5LDuc8aFSF
4Y18za3G/26TPXFNeY5Uq8Q9VntlqFATfQo/X5RoHSuO3ofFY6ncoeEUBll53U0H
OCQsT8SCHUIArNJcKyeHr4jgMNg621HZFqKfkAyf/E8zXS5eqdtaTRB6N/MU33uv
GeRDeWkKRDHBFOe3V+Iutw==
`protect END_PROTECTED
