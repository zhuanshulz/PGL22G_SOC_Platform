`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAHwNd1kyvYSRW8/xSAELgUdDqnm9D7QJ8OJadO4dCfCFK9zppgA9n8cHZTpFnMt
ySne5xtvh2zKuTD6XhDWunf5joXyPi/G+0ZBpkL2CUy/SY60wNqP2epiTRPEeZQj
bG+XBobYQgLVNFe2EwxBhUMsXeErTKuFBY2Ss1nStuq0TAjWd8JfzDyfU97aSpJg
+K5SHKvGXe7yaOEmFrmYEab4Wv24rBTcXJxfdAHhnkHWAnM4kPoJoeHBE4iwro0e
BB7GLmUdycAnQPE9PhYryALZE2dPwmAyesI9mMzcEKfls4XmZlUKdPcI2EcYgMpf
hA1nNIljL6hNY8G2tLdfM0mJSc4lg2/M0GUogcIIJ8oIPqGV732VL258GwENn5+Y
P8V5ojBvvlSu6fKQ52avZdXu9kRzWnkFQujV/I8puEvzZ1v/Eaq+W4Qfnyd1sBRH
f8v+8mvWDrGM+vVvWIXOKpRLwEbWir818fjyEzrXjnsT6pqunlxyr21jO2VoAUXV
jG8JDD/XR21acR12VMbEiZ/Oyc4qvCoTML3y1bQOQv7fF08dqAhIGw1rVKu4B9qq
cr8f9B0eoWP3cMUuNbJSq02135efiyGuGd1/yBWsf5QcpG6NYyCSK845hRIQjLDC
UiGAQSctwJY3TMEo+eUbXw7XNx9LwfHBgaP7UOiI9BCYEH9TsXJDZEgDwRpHElju
g5X5lRW7DvjOTuM7PuLXiuK667cLUxVjJzBTjn3+19qOEg1Br9BZXBGGtF9yMSDC
sLaP3U2cc3YOIi8911r3RQEXZ8WAs9TkJGOuPK47ARGiwu0OXvhZhQoevkQJ33CS
Qi5hAr+c07f+xUtL2fvz1IOOz6oU3RmKr65VVV4DZn5zuFLPGQXrgPa+7rUdeSAg
oE4YhaUdBTByCNPvipRehuMY9Ebg0QB8UiNLbebpeqvDol92WGb5dbG+zEtRkBL1
sPaoT9Hv67E1x3xk1nulGKuDg/EYpOuiLZ3wpJM+Sf3h7t6X45VEawI7qNC5R1LM
g5+Seo8H0oI1HOLjrxeO7pED4fUT/gAv9gXhOgTS88cYdWwvzvbkVFwWDBP2KmKY
D8mKnz1xMpqsEF6Jti8ydGYBbTHa0LpbSClzeyqQLQkkUh007rPP4YIDFICu9zRY
SxBd6CybK9uYdzKDTA4R5/sfcK1wYeI8QwqpzKoQxsDUpZoiSQ8RODIe8rxORzhw
Zd4P5UJDk8YO01mQDCNq/tDQgSbYMKcPW3sCWtk7U7fD2vU3hNRlkyGSZnFBtjc0
84XvRT3PgE4V40IB8DUP8KcHH6kmN7UekghGY5fwQz6Zqk4H9DSXfSc4CSkUYO4g
Uf6kcRlM5wua5J5wdmPFzjZIxSE8bjKL/L7P3R0gKdRGPYeshJlTs6OlD3I8YvxX
xft5usGL/aW8PboIuSgFjMNhd6updNjfGtd4cKKtgJeJgm9gv1sWs7GNhcEvalGZ
g2OXZ00W4DYTRP+zWCM9BCbQTVKOUjgfCt5hM/88sD6ktNTE0j3Nd5fita/diQgG
RGp/Y9Zm7v1S7atxHkJe+ruzuYzHdDOroPYYBi7W6kKTa6OWUSLUIpW+OzUBr9mR
WlYNAv7u7TF6uNYnjbmwaac/pYfPgVyIeJBtH2Oe9ppRWoJ6YFXqfYbeWBnB2mpB
9SL7nxkU3zuiKjeB6gf3n4IRjo+WgbAnnEGfXegw3+Q3NfOfadKlf+tsMzbdEl0B
3G5Us2cq6DHc34vslNC4NR1b/LY1xyH/s0AfPyNduV7v9NeWp+vwrNFZxjS5R9WW
KuFQPMN3zGBxSjXfwOYasu6XWvRDdPSId/eS3Zk/5NGoxGXXOl7POzapnnzDEblF
`protect END_PROTECTED
