`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z6Mvym01BjwCt648nfD2OyDs75cNZVu3jFQdsOcjh3xl/mRzAuypo+bbJgFIiNs9
+Va506z6xoW2H1Qpt/R+p4+yMbj1jTiEqlUubQD406/SnmKjRpDhHIKdElWd2Q4b
2vkuAUYe7qc9hgdMvpB3tBYCxbeBZZb+xSRF3a3o/IUiFz+T7+W+lnVBugnQcYV8
dYOdlHrpMMcV6yvh2YH7jsLYtcL5wWrOqKVSddnLMa2UPGY7gRT6CQ0mTC1qHzC/
WLTUtf3G+nr/KGpsJM3NZE1js0pKYBDla+M2u/DSzL5J/3MvwU5pzRjRRK/Ed9tC
RO29VH7hOoO/hcI4liQlOGM+kmm4uLHoMYj5tSK9cAWAbC5VMzrXJR/XcRlwyddq
UHbiNzDAVPHoBoZV1IA4TeeBvy6Zeyq5vmvvKC8djiDJR2ckcjG+o19ctnpoDhOf
CS6IDiUXM8+OWpuv8AHOLzh8FoYTRVBB5UvGQIe7B3vB2ngc8YXK6fM9t9ZolBqB
+2rgivcPT0TfCs61HcinVXw2iG2gdcza9qyoOkPHYqrUhleF2anuUAa0CYk/+puQ
B7QtAEJOQdyaFDxhFNSWEu77VaJfWweDH/N8BD2tQotBaaaiw9lnnoKrGJ8w3yM/
3ZqPlzWfzckFWJitVTgm9WQmno2VOyx0L97WgB2JnrLgQiqeEAWAo/hKP10M/7yV
B4tvx2etclRnJF8jZaFOJxjLT9OV0CCjcVbwQY+o/T81Tc5W7g/iUp1PjaUso6r/
19pFGBNegAumQtecb5eXfxtGvStL7dGfQ1KriTUNwWyhQEnTOsgfB5fB77a08/l1
/UAIvumzWAY6Jkd5zPwpZFxzaCXY7DKeE7d92Vdd6/AjTNk/oWI0G9Rve1aPHXH1
fafftpgrFByjUtkx0CzW6sV7HTb/kJzVEJHRzGVoAlTuWqmtVu6iFZFr+tIxwv7V
bIz9x7lVBsi/vAAfMyrk4g==
`protect END_PROTECTED
