`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zeTKwaYRJoBxVnu+41m4EzbI8GGfU1RkGOoeb7lcnSqSAtRJfyImkHu0H4FP5SPT
A1+mcP145rH/hfz6+HliW/9pTGStrHy98320rX7oVi3CTTDme41Z7JNBch4MSYjQ
eGPoNflE1fJ0w7XFz6CTuESxmsYtW79hTD4rI71ghLV24uku+j4fxrXUCj4UO0rT
9A8Z9oISv+CdKBjxyoqPYXet5JsbA8UI3EdAhq5GsTDG3NYBDHamYdocYMDrM/cB
7/foMiMqOLIhooJWT6GXBCRQo09SqI19IFfXnQXWRliSuxaIo0DUUNUnQIfWnWff
klJS9t9s583Qzj1p5G/I+tBi8h10Dt2e9e9bsIlNFFl59miksfBphJLBAsYTMguh
Suc2dtbCLe4mv1lof79EP6FRr9MtDOz0h/mBg4qKGqoMFppTRfQ18FZva9LoDopT
vo6o7acqEs+fejZZuQK6i8BdV2UvtgB4frexLI3Rzhu/KtgQQYffr5YnVXDtEVm9
9y9X1LhknOa05MK0BqzGMt9U4xF+svG9VP25Hz3b3MiHYoCLBdJo0IL6OT7wwluO
e7gpDmPulvr19BIXNZWvtw==
`protect END_PROTECTED
