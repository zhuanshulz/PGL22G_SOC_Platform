`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AoHgnILMC5QKbt7brMRFCBqujTwOy0p/hkY8SJf3bL+sC6MMEUmvbTPnDQ/NEUpd
hkFaNdkU4lzTSlxNMfGAnUzdbjEtFjNQocZ+snqPtxeaVKpZIGj2HCPW30HOg/Hf
RQiMnYTo5SbpSB+GxdTse7qVkt94yBvN8PGDiYmYJ75O6Rog1bu/v+QlAy8DKOxD
nJ6aALwTb5MkFFKd1k+7cmb0UHwkBBKA4fGkYy6A/NbjESvAwB5mvpTmUrXwiOpm
hrBwHU+ukHTIgja5FoEE+rA9QRmC3Z52IEeYADjsldJD55aZq1hLTcR5ymkQtS8A
gHUl6YccwOtp4fdYnaPFfbL3iPYcH+3Fc/wecGLhQ3+pvRtA+sm3QTj7rfRMIWi8
Wz8cHKdXePBWzCCDfrgaDpWmTxN7lX+6gYLvRJvay9DD0GpX1DRWTB7jxMPFBBlN
5sGR9ojeCmgwyen/5u19ueSyI4JtRaJ6himy1r1vFEuLXoeAkFcT0DepGuLBSQVb
29U9t2z/vDXll+4N1QSe28JnKhh/eI6RDQypVsQppspdDFKZ5RnMNpUpTbeZBx0s
9J8RUxh10ECR7Dqt0qC0Gsx1NVdRyw4IkAVZf+nS9Ys2t8Mds9unsAgHADi8dsv9
cnK1FyrWTtUkGkWc8+VtfXA+71qoDKhGGaF/EluMrykoAZ61a0l0PvMoaKIHn2xk
JTd3iOOjxjoCoeM8xUyotiyOUdKELYyGWciUBZ96hYwG9XVdYod08FnVu5K/bEnd
rnRHbsSijlLwrDxMzP3lket7ORJcKArxAfxPwF02OcObvcuu3NzZ6QFtkhLidkBC
`protect END_PROTECTED
