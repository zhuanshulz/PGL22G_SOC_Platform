`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85EaIwuaFUgBsJeYmRwexTf2cIZc2UTIBpUkNbJgW+6Wg5a9J8zm8NT1qdl6OkJq
v2bs/S5TcosPFaKGNshWTwhzdnFYXW2il7pSP5z719FRGqXjnGZV1uQQWpBzlVXz
iM54cscu6ZYLMVBOq24kjg==
`protect END_PROTECTED
