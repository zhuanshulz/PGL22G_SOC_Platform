`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOYl1d1aEmss5GF2nN3SM4efIlrKvubQQnI0swXnrP/Cjgt4v8jGU+R5BUsIRabG
Mp3PRa2/STD1wD2ot9bwEHs9K5axPEAsV0yPJOdaeNxIxZ9Tnbczn/Edry+Cl5qc
VfkM7bVVCfb/97c3gSh6L6tHfr+4PhkaJWbIsfDztpiJpItAYNGaKJYZH/KFqKuL
c0cFxC2OwC/hUsW7T6+px/V326wL5xXH0euwitNvLsl70voOX1X2MLD94BgOSA2+
p4vIE+hJsE6CsmGfrFLxDOaqM8gncrspJAevPfiAPOoB+9zLqnoLXkqT3+Eq2bYI
PgxstLv0n6ru56fgv8HAnn7HJpwTE4Yxh7B5E3DLOytGZzknvFjFprdek1NhbYi9
cbFT5VoWNcj5FQq1XSHkbtCS/EPkocnzCzyrDru7SUK5G66r2/VyMvcLNZiyhiwO
m7E89Wx4tlC6jPzLfbvoYmO554QtFsdEpEggVj0MSjl6PbGXAxjyGNEASNh7aCmc
LrjfEGlw6SJsfwTzt7stIhRiMBc+R2IZZNFgklwDxFRzKIO5nCJJknRUiKVOb3CU
y0eOACjZgBhiiO497JFiWM6AHqCrXyZXU4LE1wdGS2f1uyIkVdtRCKJQwOL2fOZz
HrzA24rfZ9to/29Y8DgRfglnxGiJ+PnUTG/csgnWyoP0FIPYSYzaKLAbNdxrEzZe
33bxZ5Bclm7+CpsOYuheAdD1IOHDhSM68UAyPA0V012ZYohQ31s7GrNHvQbS5GWX
vWdu2A57icWeuPcNkPt7JFmN2XGXMXx3p92fo2g4VjAoabQdFeReSOgpUo1METCn
nnr7F1fQafQdRu+i2EEa0Zb4GmfnKHZdo/h6R2GkiEnARFEPliZw294SlWipD/Gz
HykPqucCaeX299teiBRZoIVtOtd70XT27HXr7S16Z5uuxIRczNd8LwQ63mGM6eBZ
+qWa5tOF1LWRgy+7jBcZh7+nRdVd6FVK2WvALNuPb3Hq6oDzqSlvI3OLbmZrarRi
OrBlKutmTdWtZZ+BNCMk93K3o+qYzsrly4mNCKjAOhDx0MmtZwqvk7Hdn8JAHCGa
WVYXsWyGHhnGyxV+8JFZ/VrDwbgkHxorcHqLAMOrmJyx9fT7w6MfL1sAfEx0JkXk
lOMij0riaa4o5rlSRRUeKDaTxBGZFU/1jy3uvhzt6k+XLU6jb2zVjHVKqpR5RODt
gGrdWEfFPpJDCzT+KnlXEVXcOkyBwxiwdkdzOEL3tZiYpQMUfC9QzjnrSBqGhKUt
VU+3l+hoc2J/ZxD4RX1nL1SP7PW48By4KFLganBUA7HCj5G01SLYb4DMBtA0RtWC
1crHanCiVtO+hPh/rfzODMaos6f4sK6nfpfhsCkqykIuuUZqLQLhVIQF8SzIlHGv
1/V34NGCuPTDqsx33Uz0iGLM1uF+vg7uOCHLA+ng8zJvjh56ENiG6kvsu4LQ2hny
xEkfMiHFcSbdymKUKpCigiFVLP1gnPyD/Oiq/lw9RvdXPX8UtCXBvETzQRoxjZz2
dfo9UH0+d2wOz/eCynCw40k699aWjxStYmjLg0UONVDP4Ct7amxBYG2itclao/nB
lzzAjKzoHNPxKnJOjsaD2tcJiMZEdYJviiAtG3g0fgYz+q8YSDnaNLpkpT0yYzDq
oa62eGHphInkol4k8jhAvpQEuRIi3g0K7l0ZmGfFxvL3JedG8GlAphT7J/uo9BTQ
yfAKP5+W12azZxDp+rXsc5rlAw2Td97T9+awq+j47joJP0aqKaQsSb7yKPZAeu2z
WsUtqbcMFLGzT0nR7nMG8FTwa29WlgS7jZJpPi7rGGNvpwSfH3uQQCB+myllHuLK
kOGq7BCjKgxZ4A/rEEp7Wg==
`protect END_PROTECTED
