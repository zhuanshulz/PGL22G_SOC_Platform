`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuUPvd9ORNqTXVWm8TTC5SrPi54QnZbwyBMOJgNQDR/wBLmsfvS3bb/IAPk4SsxU
7S6oRfldpu4xD9gavEl5SvqN9645JZP2LPMIj1ySHaJMabt6RwWjd5/Z5GjWKG9r
lxtmP/vbD+kIKlW8ll79pluvDcGxWzPH2V8p0JDUwzRu9UxgH40rov0xubmxoCcJ
GCy2iV070mc9sjuGqJyABS7TaH0sgFq/RT1MYNoQCnPJOP3Cx8PpXrypFpVKczMB
cii2pw8ply47G60uOJE/VykTrGGUX3JYCRA1Av5chXhlHrHu4nSVY9rvqsdY1EHu
lWB8CD4db5vd+4c8890Fq/0a3Hty5mXJJeHcrknzjJ8Tv4O9jWkN/EK3ElxeNsQN
2aheajHtlnKrfNsXIM8QHo/nPybGzYN3Y8ZdmC2qqBXAKo6W/f1dyNmSvZh/1tWh
Q0e4kTwSXPHarK8IxLPfpA4kbnMXTiCf1+ZvPGb5IHCiUQ6EMRJmNJ7xFLDI/gzX
tEVRLOdYNUtE5Bh9pc0Ok+HUsuLgnQuOIJt8N5SlgQkxM2tm4HjKvcBfActlOBNx
bI4bu48dSKNByu+Cg8drHirRrBYEPDZdXoxaA0FdeRX6wt02Ex41msmQ+MxrvZLJ
cvN/6Zh05aHe+ipwMOHzzeVJIEDPrP99p87JNpLfuxfJtH5/ICB1gZhu7jVdbSEZ
g5MjeaRWgRQGzopA6GWkErancwPGvMVaqnZ2uNP2N4SBoT4gD617V6YsB+TczBCJ
D1gD24W7JZNj6yomhs9zIeKPBQgLPYgbc6ajBpmpD/IPpGiTj+Bm2YWNL9n9qRSN
RAnBXP7X+SJA9oMH8UJcik4YkdoH2rL9ww6V8YRysI5eB7JNn+2XuZ1jKK4MvrW4
BweP1qFfKAjMzs9AqCPv4YaulVqU0HMiT7CjC/vOM7y71mzx2Y9PxxMseppIcrlx
EwOL8J950vI6WBPlhmOoe5NuEZTyv37eMLVUQto0gbUzmEf7FS3JY7GObvjrDJ8P
tosb2lavVFmQXGjRoaN/TzKDm6YOM/pZGw4lD+W8V5MyvUiIh9XtF77bWdVrgx0F
bQ10wWubFrElQZ6tKaI9W0KvjXGQePC8nycrlL6AbIajiNI5zJWCxG7OFybZn/Ip
NMYs4hP/A2W0XsfP3m34HfiLcwvf+yWpir6j/AMPM0wa1Cf7A2KZZtAGdoeBIsTq
o1W1dnx0FmlZRMEX0583CPTw0ca0yXazAEwtle7GM0BSTxsnlSS7wUINSMutVVdD
xHYjQi602j5kk/9iC+N0cvqh31Oo0Qi9jzv+ZQ9v9QnmSGldhhqo5GT8p6Dbrrks
arGjaVV3+esx8j84eS0zBEew0CnXEHAMuPRnfZrrv09b73Sf4ejRCRIDXVa/bI42
NRVU+kuioqe/LIiXGYlA+dYnEsAm67iyFWsJTkRuIyoi7HPhun1hKOnmlGAqKNxx
Bj4pvm4wmLSBjRNf9XbLiPcVjcmLBwPgELrMIhZu2shjGz1CPWNasuss7meZu/Tt
7DIRpDnRtkbevTctf8pVteVdN+izR23gvclxKnIb2fcLOyCQYWj3YZrO1XBUJA42
pgX6w6pXP/x+J/QTpJ8EsaNVMMK+w4bjqpq5z7iunWOwxW8ij13IaSZ07baz1eI8
OCNHoxK5ikbJ5dp5m2TOPfmAbqC+VhfTPdUVMPg1YJ6skFL3SvBSJ8AtOXc9MfGu
xGvbjckNgv+yeoJDIHW+QtxkKBIudJaSj1jtYSbZzbwLqOx6XWB8ES9lbO8d2hZW
YPm7S3RiPxjaEYSlpiNgAnf+34FIEjqFq/rJLD0N4+y3QL4bkdyjLYv6dziscGyX
2ZWk9Jw3Ogbl/NpGQm5TRK9+x+vafiQRRYiJKpi0F8tIE2wpBTu8feJiW/JldviC
ewp0POdE3+ujcv/BJLtxUl86M/pZ0DRMbtbdvV2TYxLEMQB7bl7yHBO1LCLw4eMG
eRjeOtVJo3xLOA7m+GUGEVoOKmYgaiLGCwYJVWfGaCA+fzB/Sv9s1Oy1z7D0ybWU
Ep7nFy6S//Ba0lcYKBvIAmJSY2wwCM+b3YuouTW4tanEqO9WkwX1flnF9oBT53DJ
rO0SpoFC10iHWIqW1DH42ZUiFtoZZHc/1i5CyevEIIEag2V3jLnmvCWZPBwS8J0J
BujQH9iTDdH2SvbynKKv5W2T+DJSPomA9Z4HlbPUhRN+Q3muDiWC+cgiGqI4sIkU
eOiXLNn+k0PxhhJNgBEUBqkBxAIUEKiB58oQhqMXU6ZOw4+/0JJ2b0veYBdDpkis
gp4LJGSPol54Kwbh4WzNwBCw6Su5SEhkQ8jWIyYv5aY6JWyVyghfnt+kB/FLKnnV
7ONOB7Up3tuG+aRjZdEdXswigVsQjQGNKFNfXeVQXBRlIH9+0mtj/SfaRKWmFuB+
DXldo5hiodZOeO2I+N0YTLhcRukDV5Dqaz9r+1VtAnFA3RqcJkf5QdnSC05P/mSG
+Yf9/3/kpmD5WjwmjsNWYxnyaiyfD7zrub0pHZvdF5edszARawWOQF6LSFsktMCw
Fq8tsrmdWSMWFkkO988e4tvaz2go94B1RHBACoyXPNJQZG0huJon68VXlAmz39Ba
xN7HmonkczMUYHEyw6c6LjGD5ifIJEN/K3nznwve1g5LekhjMfsQyIJbw+qXx2Kz
KxC7sB9e/+7aD5S4fEzj7i2a8vyMoOYraB/LisHsgyMhjQhQZjsKtOeoK9C5qkVu
XLxvfiyA2hZasWBwcF7Eip4F/0hvkqcikTQ2l345DrIdB4fCKdn2TbCq4mZx/Cx4
IfEapqTbhymimnfdROonHAiFnCHGA+vq+LnXZsaxIPwb9Uv/B+2kpbaneAJmRf7l
4xUeKPsXif7dT5j0TTlXvewD3eWmYu9Q5QtkZVLwe1tp1pHawq5gU/Ak/fdl36CC
K0uxwTEL3OxqDdvsTWk6kT+WeVogWSo69Nl7bI6G9tsevV+zfLwUVSvFpP40MVVl
EuWzvDT3d1oR6URFRbCynL0/QexeLHB8lZb9XGCF4HbQx9AesZnSl1eAKPjarqBX
62TGNgPeeOhDQp+j9tRqJAz+zsEN21Ia/am+EjoFRQfkB1L+d+PUsOJN2wXBR2Tm
Zcf2ToxhuZJy6GTYauBmtWDrXVnNYCEMWhdgiwFGAIyhi6z5nQsyK4xKnhEJOfIA
glIAnje+gISGkmOYD0eYYSbYR6XpozzxgR61L7uNB1tV2yIl1fslueTcxbsqVmfP
3++BbYZ3MY/Nvxne2HSliUVK1fA+ERFvzuIsJd6cXEr3bjYL/fzWp+WxjFMubcOc
ZrjAKic35scNDaOUwOkg1P+BtKoEuBQi60G4DPjEZMoLNPgYCo7tVzg6kZqMz/EF
KkWwnZuuuPAzMWcBoPBgI/T3Ad5hNQZiL6tGyw5muiVBKDxW0TySs/SU9fF3sWRZ
IHNY+Vlhxn8MO2tKK8I8WC2cgX220kg7M5N01I7vELf0O9yejF1inJ3NUyRSMt3m
Y9rxCy5FJERRFiG2H3UDVq1amDciUTmvkg5AUZVhFOV86spvLRNPJV50xRaX8xlV
oWih8YMidjr8X8VByZKg92IMqLFt2tHXI0Al2Ml2BvD5w3jGn3VgKX9Qxly0CQyH
AZXbQQryUDnNlXy2RTD7PCB/3i4qdbpBO2bIDa7T6OJ4hTRi69Fn+kCTLd7XLEok
ClBkzmHjL7xVwaO1Iy/C2wpElKE/r7BgRBiTidFo8V0WCbO6ck4Uvx9j09tKSP7L
5dUcS76VI/e3UogpZu3JsgYLV3LZSE6XDVAf2NeEev2EWDPruHcpkeNbIJK2o9JB
Ob+rcNpjLZZ9jOLmpe6M5aeBoGlzLcwjrwFMsYblgmocTO/uqZMoKvSmUb4aPYfd
lXQqc1YpYygs86tSyh8hoOm8uhtBpVL4fEQNBWmn70sPbw0o1Q3uJs4FLWAxvc6x
fk1Zt4AtlvX97NQoNaxTNqOpMwkBxU3lDzXqwcnMO/HfQRHrozb0hUROMs4hiAO5
kPRb6ub3ybmB0BXPmYenVv2yNHXd1m9kyV7lEZxuHTibg75b7JwufufxwqSX1Afm
q9myGDYIBfD4tnDGRJ23Ye8ARbvTM0v+gHi2pwPp4U32itsFlcU3u0ylCDRkjIT8
YrbtcyQj9LQyuGub5DkiBhIW8X6fPjdLfyIgkH+Bp9jHVnLfuexJHafdTvX+61DO
uEKlDZ/g3pDPBZlDYTTmvQyuqMnHKVQBuGE9bSszsoxR9UevPoM4de2+N+NV2Zfd
yz4E+n4jN5Blpa+pocLzX4prC9FweSruIpvArtgKF/CymIAk8jiwjEh++YXCDSFm
osyCd6IFB/4gVhdy4oE08P9e3bcT7P08716DVKSDthN/obMBQwN9Bhbz8NjFPWa6
yZKnDFtaq6ttUPJ37hJCssuLWZjXQrqpcVutSo0T1kIksShT+yVeobQ3YJt3J7tz
KHddoUevg2F5Ou2dcELErH1aAps9D8n93UhgB8BTV5mk2Rfjl8rCk8TztPuSRDuk
sv0tb04aZ3YbKCI/rb0/1fNRz/SDR0PsT/wOznyUESPlDc4GP/CsQOT6MGDRMbDv
ow4GK+2e6WlUiwkyFA7A2xW+Sl0WxlWnO040pL3aQ18vJhFH23Nb0RDd2RT3CoHN
ES2sH+sn7Zo/jHWqfKIZyhk18PSWtXz5pNtz7iAKHkptSI/Q2ipAHTKWSLTPENWI
1yZUYd4MNDv3aBG0KJONvQRZmjQr+YFnlEj7FMBU3DaFKIEU+MdiX2oHTk0hlPBb
JALBdYRSQwKFevZ6YzfO84vpv8WByn01u4PvRbcjiRP1mB9bQu5ajeupozesm2fm
Yrit5C6uaBc10xlZTPGWy9zYrDdPxFuQu8PmeG6HrqVqglyHVNpvneAxHx1PhTXW
LldK6/YO2pCU3uPATdJCdUT0t270M3x+hsJykStR7gAyt9+/3G4zWR0DtXBElhF+
lMdBKTOnjU787ND/b8UUdNMoLK4oRpNXPQwQRJFvdntpwaWaOo4SSkCX3dcgtKSt
Ycl6RXOq7DD0F2oL7DWP4IpXyFSOk/qQhIz9ghVTrdUbePfXG9lXwhcOYH8IScGR
2NsJEZkYrg0xGDLfI2ICqku38YKMsK8NVCEOXszhQSXHLLf4CUf01hxNImtR/o8e
JHnpugnOmBJzbHqL4y1kKdk+qB2kHVjctBKhLNK/A/lWzXRPQMF4Xnv9G+s7A29J
NhMlZaC9yuXppNXDGho+/uZstkVw8By25wW3TXMQRR5UJ6ZVbtacDOm2/MAOtstm
NmC9Br6GhJNOS35lv2jDTgnvEopjVRX9lUbFmFEovC0HpUq+ma64bLzof5VJnRWS
SgX5fq0J1/+qJTfJFNdB1FHQWBjt0MYSi4fVSfSCFy8EMA/BNDOqA/2iwWBdTvgL
h12CMa4qY59j/yONsiI5oEN1QaAODuFuJPByfl9kUtKNgCvfkvQJ9oUYb3ynN5qq
kMRQFK3uNP9PrwVDbRIIxWv+dfp6QwGp11JDg7tbOwG2h8UfTxyTXAQlLnG64g8o
UYIjK37sGWBNaciE1aB5nOAPcYGIRthd07LgVT2Nmjx5ZczcCCFxhu0nEBVZ/IBl
J4dpZECUJEaX037eTMldTtvQZK51DjFF06MihyLQO4L+ymvOo2jxD+GvsmZJNXKj
cV2mL9/7EhjmBz2Ket99e4kwrPF0XL3YZS9/5NcirPsZ/n6xyZkhvLKli5bF2WCL
lf9koSiaANPCZxVpgGbTU4AmQzKwnfiqQAXBR2QVFL6Z9VqAeSxBSceCOIY1sx/m
HC4ruZCQjEzKl9Rzz6Drqsk3LYPYYNl6cXEn2ZJ4i6zqbpmJAz1KPAtEKwzFCvfr
+UFSUELU2JTUsrUtNOEyHUMWw7/5j6cDGgoX4Zg/eJK0JJkzIBpQ+yB2AElfzily
qjCS7XnhGSogTe8XXvlV8I2BdwcfjOXNvB3+wr8CX5wFmo/qZXIJ8MHu0w4t20Fp
TwNYIZ0JS4V2RD8mq8wlhB48IRDlxvhnHTKisLfcCViUK+ZJOQfS0R9wmOi2Uflx
RECdKh0KxvE6e2Nk71Je7iaNN4PWWp8jkHvylrD6IGSaxU/HEToDW6y7egpGn/i+
1z3qjUWIaTW7MlNogNvOBQB9zBQQGcEI6P8xMQk17y7FGzEK11JaQhfn44VJ59h7
u56BzzXqALRsYZV6V+QGfGqWUj7JFDLCs3Razyu3Up91uV1nHrmnXWpeFSPLFMLh
aJbA52zourYy5xZraVB2Y1TcyVtvglOiUE6SvrwZ9AqMdSz+XW7NI18A8RqMX78R
dPei+FoKyLOOJ5QMV4uMAsJsPY89xOkRwd/p5s/vdAk5ql/+8Q/2TNjQBi3LBuNg
LIjBXd6AOshUwPEsa3z0vIB3b6JtWxdp0J8AHXBhiZsVv8/jm1cU1p0qC5IkEq6K
Xd3Lklu7kRn3KbknejVVFNTaglUTEYhw9lfID62NaLJqpq8iACDZSxYN09Jl2KR0
zqLnivCILXAxrJT1uezjK7ASLVyMc8PDdb0c3NEZBBrJIT34Dm1aG/FOf0Zbj8sK
9UPoPqKSxiFNQVPMZbYaitDxGtui6M0Uu8ksOOxByjHGPxlD41BUhQgoFkTtlAp2
pSk8HSTw6cc4nvlQiRE2nS31UehiU3qaJcTIU7Un62eglfDWP45LgE7PC1T3wC4q
qOpDc/TB5xQ3/1/xQxd7PAf4fqtbztejZ93gg9ftEgBl+W7U7EH7ZTkYhU2DGMJz
4mq4IMMG8+k1BN+TxsIOY2rgtqUk/Bn4LbxEAur7UDu1HpafZq0hsE/qzW2jHz0W
sl1YWMDP8yMjRmhbQd0vkZADwyP13cih9suCJbWNx9n+MakF4JqxJUomGkUR8s9d
d8iIv1OLwsXt0Jf5x0u3U4LigLM8/VZJqDSv6thIEg/GFgULTxBfhYFtNIh4EBMM
jVrpmNgIkt6t6DoqUsn5aNioFBnc7gsMtnIDQ6uKJYnrux8jwFR8PWfPO75KNFUm
G226vVYolC8DdOJ9zmX4rAt6G7mZyVB9ICa4k8IGRBBqdLOXkNJeTteMygpH2cc2
rDwmQX4GFbyv/PmZ+UH8GLxf+pZCELIm1/sclNZPoDPYMYtN7Cx8QGEzbG4iXTqa
7lRjascup8k0aIYKRhmdhvPnpsbImE4/397qDxhFY6fVKv01Lglu/JE3AX+FwHAG
Smmi8182BcULbZfcI6pyH0CmLVoi3Uio44HiexYsjfWFLLR/2vWtslCfzH5IN93F
inHHMRPYRSNGxgqgATb03tFRROf+DAVJRrOgIGYG8zNVw+1vjffflxxGUeYhYu25
6znPTQoFg/hzC80PTxbytIgSbojZcL2LYg24h4ItCpqhq5uMoYYMTeNbeP75cNF4
l8j8VV8HSoaz+IcmAB80kpE1x7uncskazIfAuO8N71e6Ct0A9FpUDB7DB9Tl8f88
dXBlC+pfPph67cZALjZ55JvMZPylsSJUblE4pezCMngdI/3t8trSXwe65upOMwBq
DkTJqxA60H7M61cc+SQAUHKrTRkL6065jhiaCQQ7XlMGuKp+CP1KDL8k6QLVdlMT
T0xW0q0S3mWD/F7XiCz402Fkcr0efVC3Xhvy1uM2jQ6ci2rBzjRqvX3EUF3wgNbJ
W/bGl0WWw+A3eV9QZhc2huHGVnNM/Sajvj+KQ3HwNMqQ3pqhe7DB4Ep0oNpK0j98
l44HQbWYYIEUrJOxNEnM6T8OILHtYnOGLEunSXMsY1xvI1BzpVuDgVJBxfQDW4fc
tjvZylFmG30Tabwng1pUHYVjUkRFnM0CW5OTDVGEput5AnPjzwGU5m+H4vZZpoEc
Ij6Q/+1WuZtyh/6ux+XgwxZJgIIvRd1i1zM9Bd+AdptaQ7nK8eS+A1/33ThnErh1
/gOyqIPESlHVy83k4lBYM/qUuhzS2rO8mVkqp1bY4MdpTOtvjXZK7w//otx5qHA9
bwiWbhYpFOePoIUQht6Ju8PTg9aaw0oRsNcX+SoiWZ7XcYnlxDYYPhmHUlrwMBaJ
YgrhdFlqJV+zsEW9GX+MhKR/MRNktY48WxXMxSAfuEsGCcH2Ol2WUeNEzgE5K8lc
ztYE1q5bKq6IsbTMNSjz1YbILTtAle/zkUO1SA+62XLlyWaPy3fZMOWmEvvIlW7x
kmDBmpR6aaSK7D9by0wUUh3zl39/lfXdRFgPYqey8xElAK/EGOjhCkoVxi9UqKN6
jXo4op6NVlm+6JFrLX41IWn+4T9SWuB3WfjONSaKwYI76CmALcTxI8IkIFCVHVq2
PnlYh7cprYZYxHs8TGJ3NV8nnss37V9AhbRRTp4xRpNKORnLOJ7aq/bXVwiX8AiR
f5afCgJEnGd+tJsU4pKKUEPsjZ+dElKIFp1XoxmVaBU52qVCBigSUQCdx11xMrUc
hczWfm8K8KmisPM4sEGovZnyS4frYlgdTnQpjyKOyIiE/dHSc69IABNuq9OZmzBB
Ul9eUPwI87gu5hHABsnOsXI2YFpDZ08pUCtOgBp623tMEHVmHmxOo/zH+TCuk6Lt
Ff7f/OyPUoGUT1M60n+9rORnSVjE3EQOAl8Dy3kLFN6KhYWB/47r6DMjy2R6q/0U
poovdI2Z0fvPh3VK4ZDWqTSvywNWgE7EEaFV6/IhWWQyiBwgPeCA8/4aQ6jsJwP+
OcO86on5mhm2Jz7UQye32tjSIut/nsUUqk5iDbyZTw6xLpBu44GrLWisTwYyXtbC
I3JaDwGf26kevIBCxJ+DpJRNrW0MaPfNROuSrtlOs1+ePuRhB+oJRvhI/KAoPewH
BVs/E8UimdeqykArp7mY830R2A0PdT1EgvFDjLRF7IXkjSiAiU9RMGkOftUseaJY
NCCzweQCDTvNhb4oEbEi/2OLFwX/bIzHVAceeee+MwFa5gEQfg7Hh0lK9A4fBRdo
yQCBTcBgIjT2dcj+N+E4oy2D7NBp/lWjC2fsmwwGlCWexo1ufJjQuW4SvEzSRRAO
FVl6rqOAeFoh8FICyp67ife8PHZ9zT8YGFc0lynTZwJReGfwC+qwT998T1klUJXd
oKgZFZcRAoyYpQZTK23KsCHcXaJCL0wrMUAzoF41Gbpa3aHHVc1zkfX9VLrL0DJ6
AKVB3oXC17RcWBm5zMyDBdMuYUI2FJ9BjyXy3GhghZlMFW1T3jby/fmXZQYL3gT3
ixAQIg8G0AIzYYHPmQRmafK6D8J/n3eUDAsESbJY/lM1w+25iLjFL6mkwHvG2Pw8
CLTNKfvIZDYweGudrnKLOlrLe2sfthItPd6BHvGJMUcgTFW6tduwAHRC4OUZwoWl
DL5/s1qydfwpcpq/5Rqa88a7PL09s1ANwtrQiDSjAWjlG3N5umBrXqKkInnefNxi
B6xfsQ78Md7pBatI4zJUotdnm/ixygAv8Flrq/t2IBw9hX5cLFK6gzvCRyKytkAk
zmGyTRtxZlWDcqyRV3b9A4lRyDocx/i7vHetKmkvOfhZBHNPDa8gNl/VGqdA4f2S
IwCwnnEDtKVA4nnIum3GuE24bSONZAY9z5FupESxpkycq63Mp4ozyQYJbB/D2YdR
nhBeN7ge5aoHiwNeonaaEzG5gcQxuRi8PATDE2bzh0vcW4R9pHkiJGCtGjvoSLRr
V5XQDFipD8srcxRzATA9awxNRhnWEQsptW3P29Wse3ZmTtp5hhcCzand4ix/6Zuo
akMjVPnAjKwVB1PGg0XhqAt72LVext/MzjlbxkmVhzkCb9ol7A4ygsAmdXAtIqvu
YR/aBvMkQqvVJFD/G/9BQlG5wfG6X9G0gr4HF4XLQvg=
`protect END_PROTECTED
