`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hFNyqXQBt0hZSPY1ZuzMl7ZcB8cYuGUgVxP7gjPAEpiI9EboMU9c90hrW4tsxjj4
6Mw0VBb3hH274G9SkjahWPLY90G+DIQ+SWDGKKZf3x4NjVD983W1vTT/rSoY9326
BpuqdvF+YClhXUt3vd3Ee5MFPd29WvWs/VsbUxW+Em7lIYHiNFye6iY1EI6rWvaw
6k2nWEnntx5U9qYciTB0PTUgOru9+uF5/G8uHaLPdUTULHPJlfFFm6maK97lp795
g+1HF1YDXZD47g/eB9a3e55/XX5WTUxii4zvQ94WYOuZreEk1sVGjdSa5gk7EaBm
GqyT25YVOWfkQpOyuvvLmyYAPrxxl+hVEOMszyao34hu72HNhKwmEvvh/9dxqd3k
6UdHkkfpFSYwtg+vjjS8TR5h45PBQfl9jicL2kvynBg0MB7jTy5yRVwz8l5w8chI
WcfLP5VF3FGQmoNEqOYhDgDVIiwdSQNdstaofuTrkbu/xZZ9a56FUgnBZf41EcAA
2oJmGV99dyQ7wzOGF/G+ZHFRxM9cPm7E0WJn3GeRLD0n5BW8rhAJAzXy87DWSzAh
PgBepdAd54Y4lu3jyn5nZJbFeOKLaiJS0Ns8GDbhjUj3QmA8hLaxJzyNQ58mWYKj
w+rQamjDVxqtSP66dTD9s0EZcT4q0ziN8PY8HMBz00uyMNFlQHRLrw3oSye9f2V4
3ttriJRjm347UWGF5ClQmA21+J98xwluPBH7R0ldxQpl3Kayr9+jK16x52iqAaR+
vbTlmblsPRw4AqN18EYqWOxq3zgGLpXpqpJfqKMfuu3y2vKsiU9TXs0mVB6HVbC5
nySLrH77UmQooIS/H2i27mcewiqbVCEVlp8m9rbXR4iI808vuaoNcAFQ0nOFag3n
lDsRZuy5Aq81WkbWKJeNVjqa4oB6PDUY9h2DoKVzuuKGlst3Z3dit7H9b+B5/dqi
TPIOm8/dhHwtWf0adxWhGEW1ydpMA9fBpS0uavHjfLnq385xEauEYl9zXmbHDJ3j
ux4xkhu0GfFtJHa8KylDRND1J3SbUHxgsXuclcKlMbSGlaU0RSn3phvyfUa1zpW4
CQ7U/99nm1NsGdCV4L+15sxuDgn73lDrKbLFw9slv2uX8L/mXUaPgMeoGvwRW7fc
TDRJtNL++Sv1geHNSnLwbCSbLth/ajfUHh8JG7/QNL5G/TzuYl/wkKydVf+yZyfg
N7sBGilieLRrayXi2AQsRZSrWXPiKweDuiVIClSD0nUDPC2e0mvoVOevDoGmy+aA
rwtrr5Rf8jtLvM7zLImaiwEgpXmI8gpwbKX86/AtnOsQBk4yI+RzJkMz/OVWCpyg
MqGjEVVS/lTuZsWGCAcC7bwIoOQvmXpZxHnvsMrhFSUZyJWXrEQ5vADShVzdcgy9
52n1dWcLyhuZOt5jO5xukwv9/YbtvewF8KqNogRTs7cwiT/E7amNLCd+iv2A5rhe
8HGr/qHmu8vawxFzbxAS2BOSHeDobPq4VD/T3b68BsWy1sEgW/UaUjDacNVgB9TL
lvGZR8DDtHRE4np/2pAbVxnG7cDqWykyEBd5sNX8qcOpRTRUE3t3ogD4nh5cZ8sq
rKlylUgCaYdeYA/QsP5JtW0ZtOXYzgbT5uoPC86/l2YvpIKtomX3sdYHAJ+Qnnlu
oguzKmYYvlqvuO7st7+iaCsqVwM2So9hrBOHo0Wx0MhOTGk5BKf+E5q+q1NUegpD
8RP2C+IA1Q89jx25yWSfiCEgY6YIUIncftgeGlQ/pW4j4ThyBksqSwnR4KvreE7T
s53iLVu/dQ3PBsABbSOzfQWftGk7nJZBNJSAy+HPBdOqfi2HXaQ+rOVBHDK0MNCA
9P01QtGg12cA6grRgqtoOC7vx5ScqsijZGUpXRlfwiEvPqwRsyOxvrHvsKfJv2BW
cBbEd1Bgh8TumSY8fGJ5iWpNYGjig15jW2AAyLW+qAIzll9z9/mYTapq5d3MpKda
Q7BFBTiFWyqxMHUYG2JQRw3Ac0tp/rThFevoPWs68JiB+wh0zQYmitN2jEaT0Ase
7LlJvwzYutacTKxv3hgvoKkezGaoRv6IMFiFQwtMv5Pxxezy1ft4kDsbscJBm2Oy
xhict8qGMR4Ub1+yWbhDwNV9niXiXezoFEmtI9Wsw22P0fGMTepQszat6nMuyehW
KyqzxkpH+Xo0ah7pqOH10HG1ycQAcZ8uirn+8xdPQaUYjF1EjiOcmlZ0Z/c+Stp/
JRb9yS8IP2zrqY/kU6T86nWek3Kj8V2dPN0qq1yfv9NmQAio9qlf7aRNgjKoU5dX
rGyUTImhwUYcpnAWH8n0SAw8uQh0YyZGujJjdJmIv1kV8DAmnrizcl9Ji7vzMtp9
j+ekYsAhDQmQLsNqcvnukq4BH7ZAIGr+Q81OP5YJp+CXQbW9XgR9NU9tf/fF0sf5
cBodMIZNiSnneo9u1dmcIibgaT8wVAiEe1y4e7PxAzEreUAmDayDMP5TvC74GL9M
vlZOw0qXeMR+WBUUKDHzf8PV/es/sElp5gLZ7WgdKg4QPTb3BtjnRFSQ+Nt8dBH7
0xowFNNtKA9KvZXmK1m3NrgDr11eKF/2MxCOFk7g9iXAd6xzh+1aJpqQTsbUGAg4
`protect END_PROTECTED
