`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LraLQ+DrB4lX9Yf9CiRIbocWHjht1/jPXe27BIAaQ4s1P4OQZrrqveuh70JqI2gi
xF5Ahto+hxU1T0EaoE/7FqHQmYIOp4A5XBUtIeXHG/p4dEDO22TAVhYgsdrxr0JV
M6YDK871QH36cIuinbb8DxqPeP8ii9dTsKrd0NIgGSqPGwmEgvBNgDYR80tuSYG1
XUhbBF3RJcp/C/FXFAKWylFjk69AWQZW+QD887L40uf78ufjZDYUw3+HqR8G61Gw
PqzJ1oKf32QYVbKoM2ftIZ/Sai+Z66ieT/ETuTY3KvlDDHSkChvCppDFSp2frMFT
QYJU5dt3wWC7ZaKES/2TR/eUFthxJFrKx5Esjp90rLVJ5bhfRDO94gU0sZIO8ptN
iO2HpHluoGhrsSEZwzsD2S3Pge+KiT62YuDClkHbkyl01T+7AN0o1Jthky/7kLrw
7a4rbYVymCeF3mEBigOpE6UbAZvFgNqUa4gasu6GCADVLsjihpLszZPnVRas51Db
d72tFNMRsDmg76hcGzSgdguERSNcRtZCHJCe4rCX8qBl6+lWxMvXu7CIEtMYbNK9
noeDw4lfb+9THtaJfJZ++rpj0cSRTk2YCi/QMPVV4PPav41qnKqEWvYP5+iWdfEc
dapUL3GpBED8q+g5/07nh50VDRUfdOKdwT4WrufmiWpDowiSz6kcfxY0z3GgNWK5
bpMm7anWSnhNVu8b5QDOzUD9EvLxkAG+QUPspmjGQh6QrUjI0DCvh8jcwxXu+df2
cT+5j74mkApr0KRPFtHfYQskXNPP64iZG92PAd8Mxg4=
`protect END_PROTECTED
