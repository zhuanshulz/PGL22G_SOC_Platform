`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+bRIkjkp21O6khykSg8YJaiHidy7Lz5Qdco5VmooPaBh41jRjc9On2mabhgqtID
zp3Wm1kroJ8rxfUb04FzZi1nvCRcTZ4j9QPK0Tvm3+kAeShGQhfuB8Ag4HxjKNmu
85HgUNuaUALSRCkE/1UOQjwpnyh5KmBSVCbXjJiTDWKDnrQj0/iCLR5jTecAOPyK
Gw9UwKU8/5EJs2fTnfwUCwUBdx8vdVi5TVLqfKBlqYp1teZwHFFUPxAPM56GVoHo
VXoy6FePAa4hcBnIrwbMw+qIa19AcpCMDuICmdWnxME6pZ6Ys6ea+/1GaXRxWMaX
MVpIibWsZZbaitw3dCfnPY1vQ9KoXJ2khAiGkBYX28gLvP+KV9LxDxdyhJeEUbud
TupmSXfBIKakxi2ndClTC1pwFU3E7FVks6zi3LABn4CGQ6M+EwMyiAkk46DKqN8T
t8ZRwnMhgO0+2MQC5fWD5tLno1nn1ixCn+a7qBzPvAUnOS/zslPYyL0CggVJyHDa
PGweYAMYM1gD41dhgwo+tlzVW2u7jI1WwwXRR1G7x4Zg38cqk8Jlb6hw28Bz+3DV
uAF8PSaP+8OT4Vq7Ar2qY1U43TgnCQAEvZWq7Z7gwM6wp76EcM8RDFlwNZWKLTzF
HFq1u1hBLC7lJNrmoXrLPUZws+sNdwTCeo+yXLzq0CimSyooRA2reb0O2Vc1ynzP
wBMybnUd62TnVW9GPNRMVGY4bW2YHtTSK2P6z07XXzOyQBRIV6Hx4gZ3dq4c6WX8
h3tQLt+DmSLLLAfmAGXEqnAol3wlfLcYteGFqSswmkq+46HRmiaacELdKYjIq4to
q3hCxghVaL53dtFnSmdrKrUthuQJ5I4Zb9c9PFd/xRTAjVvJOiCrWcHuH9IMzuKu
Di4i9XK25fpEW5lDsFiaJ1e44GbyKDdNtUsidmzcjxpBnqbX5iXMQcPXfUaNae8b
wgas2LLW7ZMSsy9VsL7NazIMwRMdrp7Lwab0ifGcnJkHWBgVNq2ENi7LV3BTGgj8
UfL2niYF2BMqj8jIfrJGj1XWN4RjKhcbUSllE6jNUDnqkLqLNr+/8kU3PGBqPjt8
i7zi7gon3h9w4L68eQjGBXA/e67S4lkXWMUtDzQDAl2gbqrXLQt4kx/+PYel064H
TeUy4sa617KbVyR+xcMZDDegr2hKoxSok6UNmqYBYbTh2cW+TztKX7uy9tlv84QQ
7LYXEUWz92w5svIfIg6XXHw3XBGivJTM1oH/RV6FVEsMfggKPOE77R4e6vkUJVGd
r2r6ZvCDM8qot451UGQaSODeP/xJOoSRo1qoVPhC3kMg34YfidzJWQbezvvD6glZ
AaJznESHi2yADhb/QP9b6CyXVCFk1oUtBMgNEu0vP92B+l+zOatMWySwOjZEMCN+
U3swh53aoiAu3LPb3iL1T/zsgDECA5Uu6F06hAK5CfAlp244u1WnA280PlgAh+Ya
0YVD6DgDLhb+yOhgx1md2q77VP+nfoQjYJ9gaHdbGtNaIkAARV8rA98HKzC1szTo
srPk2reKfBwQjWYzoxYoMfLmje0w5/I7biXpafEMnsnt03mATBIeMnphAY4cy/oO
D+7mjanTL/fXR1B/dvIuVGfxf2PVRxGdgZOtCUaiBAQTw47TSZEO4EmpavnF4Z69
Mz2i/42cfmp+w5Lo/X1PCMSdOzwdavumzZO72y7gV24ksEAk78X83Pv/X+5gGT6+
ds8RN9wB1fBmn7kVJdiVg/Y3ggzXfl2Ey0x6XLQ8tr74+FSbh2aT71IeiIXbM6wc
S+Sgn1e9YsWyIJbJUsEvnv7AjyIuVMsp2KH8uJGRwaKwE7hrnEY9kSB2tdvdR4IU
bCp6YLPQnpTHaVjITGmwhXOa1Av6hYjQM8UL8ok7xlxUo6vr3Ow9sTBq5kbQQ7hZ
QB5nn2E2xwhuc+Ib4bbUHLnQDYKvBB4Ib0afFmd7awTQ0AWdIQ7LGZLGVDwXvDZZ
TL7AGfsRpWUZCgcFm1353xtc/YCcPU4Q8xr4RUV/ZPSSNNVcZzBhe6Agqwh76Aky
25QsKqLbfeGXmE0fJKcFE3VpATnOdIxFTjAzQmceD4trxel6gtjyTMUqN0w3vNxb
haIFenY1thBT4rq+r5MzQD9W3SFDU6li/TjQw0V/9ddb1MwbnlHM001k9n20rtBD
xiSspa5TiadVcKUSvhXVm7P6Y2PY0RYl2Zs6WAmK0H7aRXXrQkkXUj9awYQfj5v5
w5/8XCoBuG05HJYkg1qQBanYe1UXBghOLqxCcJDuTIyh0VbXHKjnYK81PaM+wxOY
b/C2jmd3e/8ivb+8j9dVr2oaVzEUDSvFgpWikI7QhaRu1Hq3sZnJFdqcFtWcXkdR
VJG76BbP2IeIvo/tg+m2AWeeLI3YIVspH1xJcJQ1RWkYnu+mU/epf0ChqBMSqgbs
ijWd0SqwjNsW3vMI9qnVmYT0CTtwXjPkCadheed7SKrysbVz01nH3y5772s1gWym
vpynaGF1VYCNfA2UAAE7Vu6B3ROJaxq0v5/7rQSq8WMR+O/qwmCCPmGz2edg9lA1
drAwy8RCDTuj6GYkKhM7ORv0/fbVOD2VNSdLyHpiinPRr+5JBLyPJ0e53QQc90lV
wuv/fDZoS1Niu7aQ3ny0VD2ynOJSPD7V5Ej3RiKJmX8GrFWUpgRbsemkgdgDpyac
+SRMdZ0rq907Ony9zTo9YVlPPd4xNkiNNvkzvy+Q0LqRfRnkUl6TLN2JfFUysrZh
BJYaNO2q/AP3peYMZdj2bp/Nne+c911o7DtbNCcSdADtqAvoqZDzrlXrJEl3DcSq
zw63ASNx8rM1jWfowHdqUjCb3m9PXFZWI9LrooIrLvesmqqJiJqkhoiCxLSbu1G5
V46wAiW7hyKaJ9sWHdRdAyEUT0AONLDhL9aezo5xwLW0IBC36RTllMuPcJ4DDdh7
HSeT7O0z2+KPBNF+aCPi4+/BQjd4PegX0Q/sLOMb+0SVsw8/OobY2gO4DTfL9axx
hm7/QUCRGYnidDv9n9Ox8d3QB5ozG7nkxbvKDiAEasp5WuRfXzkRVGKYoJalkQ9t
G9ptoGeNnixUlfI4pGH/XSQnnP4oxuiAhwmMNpIE8i5tC2GDUCuJiCZbKzew27TQ
YhtkVG4dHBd2BNVBNjuT5YJi2pyLF6T/L1nG7oKYPm6yr2xjCYqocTiydKOlGKHK
2cCI5XjSs4RULKWkdvm3g9AXcqEVrKMtAtcPZzDCYRtxMjKqffyrweeBL+F9jtWn
VPhSPwtWard9H3IgpfQnvMkYF5h8wvr9SmHWN807m6WGX6TytZRPK4jWTwp1YYRk
W3lf3x3Px5ydQLzJxjihtWV2O0T2cVbUq8XRkyUxK7Lh9saeg1PqPlVNlbqp7W5V
lap8kifLk7B+ivPxg6S6XeDFKTOkGKrdiVyYNtRp+X4KdRNghhZR9FcCDrRjK1tM
cM0vzOkK6Nafb82AqIuy8HT6C6jKhtKoRmaXgK+6qHoC44my0r7LhvzalIA3mC6w
1v1+KY1aA8sOms1v8v+J9rQ7BsCFjP3KADdRDfnj5dwHgq36XIwQ5Vz0dTh2WeW1
StpnQ+LiO4PhJS7mCA1R4q0yN2NEisRfAHdpNLtq4s6dMojN8j9EXJED177kvA7B
tt8rFIFxD+xSefc00EDmRMWhUV0pBJf/QQi9HjeCVnj2q+W71NZoc9dzOX8C+ilL
`protect END_PROTECTED
