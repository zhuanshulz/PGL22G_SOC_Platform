`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvhBNZd3W7xHClDSq0mhQm77F6rv0YfNoWahq8g7ov7q2yFXt6+CugYODAb/J6gn
WBLy06fta5/LOm/jV9VzOCzrcTmTn40IDrYkQJylQILv5l7ifT5C/CnJ1Klcj42s
2mt9cBQBbPiwcX7vmYgy6DHpMUHAhUjzaLLmJr4A/tYZvwbITN71o9ZhaHwYr4Ol
uKCMnVtANl+njhgh7tEAlwNVkeB/VTyT8UaOwx8z9Cpz8Ow5R9+xkeVvkMv1fWdF
adtYDbVh/0Mh9rxTZ/EEXP0kaj/gc2PQKkfrJ38YWkmS1B9jKVmqtXCaqXGWXXx9
m/oy5cas7n5B8UiUlJEnIT8F7fk2nJxdf3gVfuzxbhuc48Fe2a1S05sVThS6dRnD
y6Mp3ccwuCKZz3TKWtANW6gswpRG/IPV5CtqJ0ylGjXHccwr7I/SrTMhXMJg0MAM
3zrpFFZM2JNXt9LxPgPHOSxZ3+XTErgiLIb99GodK2sYYKKFN+4+HVJ+FFpiATnK
nnteUe+atDuYC/74U4P32XAzGo69bKJcQAivLytkl0WqdPKQSDOOT8qMCUVC7q3N
ybJKmvnpj2N3tTCJ5QsqFKzi5Whfe0orN2XRjjjqRxhBLy/lTP8NuAFgGnhpQc2+
rXKGSXjdgc/VZyKuztwlmCsv0E/X4i+D9ahIv7KGK1IHE69PTOBOoeHYLVOnpZ3T
`protect END_PROTECTED
