`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9sD2TgGsFMbc0qseC4BwvWvOG78+2MuY5JAgB2703kvPJ1m/Vr41QHEZ7ELclLP3
NngF5vpvVb7i+4UCqm4idPSiQsyJ1poCh9hGg1q5VncI+1LS3GhjAnYHFLCytH/+
UAXsno/1/WKs5xBf1z5cmAvsE9F/oqSjkLh3kdxKH4ShT2C3pF1eYZc9Lsftpmq5
EMh+ORkmfDmLw+ffLbGaKc9PhcW3iNazlb9l9fg3rb5WtmgcNsrrUNihI0hODo5T
k9HqlcrAghRAlhwhCcNTECW2Sw6dddpjzNQ+TsjJD63Wg7O3Ezu55XWThl8emFAw
RIHVXzmwqmg+d1393aI6VURfYAQdLElgEynxBktpLJG0TKqTxDbJWkliY7vUK9iv
JZ6vB8oP16pZsay3UwG0yANo1LTTkB0fY3bl1FlPKuAw0Tv68U9rn/HjoRH+f5ir
+U9rTxeDfUj7nwLDxF1zJW5n8j6ASYzQLm3H2KZ+LujpHl5Z87fw/TvJdje84kr/
MW8Gubm26GkS7bT22dpJMmIDYAXygfW33ulpQF7/qtoXN293m7L85KLZs3/qJ0ty
2pmmXnD924Y/VQIjVVPi9DQsOjZkenK7i/kfJqoRYsTJEN5AYwNpErE1hniT1qLA
3ZhFsxvRDzmxDgihNhUghv43050G6InhPeh6IAQG/c9c65AepHyFaJbqAe7UAlAe
Q+D8IBfQ35x4wyzdMAVwFbPto07U9L2ChSCVhGcZW2cCMVU+2iv0R+1GjIc8IHN4
4YyLQYAGIlCLn9/RdLE3n+RnfO7yYmouTbl+COdsHKJ2zR61bbzXFhWZN5yrCaiB
HEvlWGidlPtNP0iV0oxfZzg/hLj2qqzxXLhmedY5qu9WF0O91u5Y+d53Fkp8k75j
`protect END_PROTECTED
