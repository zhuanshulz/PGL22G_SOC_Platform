`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
khHgwVQeyhNwA/izOpRNaYdS+0jpLJCH1iWS19nUWtqI2EPPYHVXKGPhcJFJDU9K
mR86zL2NQDhj+QJjaitZyGzmSOX2R7QBgoUvIGvufg+wWvMXx3ojg49AQnxoGcyb
OrcdvY8aMLKrb89kimTE5yP1uNRGN0F9x4FVSsqA2uHZRNIwMn0zaaCgl1uwZgcl
w490oI4vAcUKre8jJp10cZ2ZcIzxiNuxI3ZUZMZqIbIFp7Ehp6KNB9y4N1ByxEbC
//KC8opQHW4vXspWtazzDozli+8JmfnJeGQaZ6VFhlAxABS/0VWilNEsJdIXLnxV
XObj5g6KJs+JP81v/61wUV43IKugFUM7bYhQFZacb6smTjakueAyRBXtngQ/MzMw
ZVaADhuq0h7bDtSFwYGNbadEBp2zGo8YhLx+2F8M4x2e7SsXxqP7h5pMONFCrfUN
RTNWXbVoOm2gnKeTRjh7nUtBtnoA+l9rbfoMNOAzQXu1ktipEbJDG5tLoEPUD+i8
HveSSqMzCJRzSirztWqHuQCJfRXFdTz3ZBcVPrfX7ISfjhwFbR0uNdzpPj0WLrPZ
IfDlfqKLyGQLoriyiSrqGnfvGpAAilCef2NJwsUebbvmMafvPs51aDyWgt9tfxen
TPFJXWaDc0GMHrG9z0Lc/DYkkrAcpbvWk1YPl6V9sNhY9gqmYAtFqAs669gy0a6W
PDWnEaK1vHRAvPqTmZD1dZ/BnzmBSg8xco5qyLM2MDG8j721v+OWTIdEWwRnamuk
A+xovCjMbM9X9Uk7ZDkqNYSpNzzyCrJMLgOryV0n9cc=
`protect END_PROTECTED
