`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrIqFIdjXTrjVmpttjUyeKt4z07qrD9uiez/9DsLUaVsegJCWgKAiqTSbL4W19ru
36WBchLNgxrW/BlDvkwSqEqlmS6M7WFEZzfikWQybBD9AiV23hpB2ZsaKH3zpeML
K2bd3fERpfYAn9oQTkeXw9uBa+zNFx1kVPav6aYaR+k78l95vJPvkJW3zWPVHISo
uZy4DjJ4yWtU3Lk98rYKVvudj3Pq92AVmW8xvaJEj5O7WecZFkLm1PIwgYX0iABQ
vPFRs4tsLuiEBDeQ2c9V6oqgranvHo6Pkr94/W+SSTe6WOcBhSR0lfttiT+5Fid3
vPmikzNhYxi91M1WE22LNXJnLLZOnlHhAErqLcpu2iuVixc0f3vcgBWBbrTXia0v
xyKO2enA3T61nV6iWsvePnOYauIQIJxhadVI4kYaN57HwJ796kB4nFkHxWM8KS63
9tcs+oV/cBGVRSuvtF66r3uOSg6L3LDN6lw4l80HacLrrj3/NglvXAynKj1Sa5nQ
yq/ZT4OINkYtMXpHhm0rUknYKCiw1HTNELmAAf7aUg3P7DxvmHna6/cjitLcLxQL
sLTAmBX48Kmaw2w+jOTrYQ==
`protect END_PROTECTED
