`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E97mledRNMW/SBc/SnhA5U06SrdPSi/hljT7+AHs2RgzjxnLwyTkBML8tsHh1tq1
wyv31AZyY1E0gG5Q2tg7d4PzGC50jnBdmepk+BekPRpo0Pi5Z1s+GSaNSiMxGfwn
xroVn2NFxjj/XpADwJa0fdq51RHLi2kEDpakZ3tmp0xVs/7Cm6CnEUjUv7xuOun2
3W/mF6NDgKnHWSrbKczHLRuoeWEQPALi0ig12zsNAukutXsySy6rvoO80+6Id7vV
iFhDd2nAZnzFGmwCDbJlYf0AAxR2e9qoGvwDUdh/CXmcPMbHzSraPhuPSqS1Dnrz
0vLmTt4y+LKM2rQ0+j2EOypQfoiIzzu7h862tivkR7swwcp1yyyPXQfMQbzi8I2G
xdSjeUBYxRO9zadySoNVSxrFKV5Kgup5Nhy5R8GTQiG+XqgNebJov2pTDQZ8wz3G
68R7mTu5J8qpKyl7q6egWVF4cbzGSB1AFCfHE71Dz31FJwBE+zg+aw3R4JTesToT
xTe+G8vGCnHDFIlcdc6P8ScHNt1275nCuz/uJeRTlJj5fMOXPeLS0pkeoImjotPv
z5lc78YiAhk6W38VK6e2JUPOP4YIWAGPgmYGS6jAxLx679xktWphq2rPj4l+rHCp
g0B2N3b9owhaTLsnrtE+72vjHLD1crwTb5mclhwKBV0+Y1UQimUog/JJqqOpq9N9
vMCc0mazcTfGL66E5tjrcinIbMqGkI5JQa0AZEEwPaIBd3rmfwJBtMf1k7CqHKg2
uFGTXUNhmV7vyMdaulxtoya+ZyLxXIO9iSKZwWXiTl8jRO5ws+74yvTTC67oDcyZ
nIhFEK902WlPy/fiKuHw3YhyTa1MPTTj4yvU7mSRoAZ8IyhTMEnNCFuvBAeKjcvj
/tzf4+qzLqGyo4uDQWm7rsaeNS1z9U/EE6+OYVLv+2UN23hsbDiGrDqWXSXv+n6o
zJ8VorgC9uUQezIAuInQPfNxS580eYB3N2G/+/r+c+NWGCD1SHe1A4+0aNr8HyWX
dIW/I0+sGwVxCGP5tFbcff6KAr6+ISqX1qUCSb2hgaXI5Bu/90T1OAdwqXtqCQ6v
HOa3VQXrBUVQAHHlMUWaBfgtbTiRalpNSPkTc4yRaNiGWshgKf9GAtLvel3Wjew+
7j7heyd/6TalGf78TGD8CcT7Zq2FWIAE55W0HZK0beFkqUYJ4z/N7psbPDRKcLbr
L6pY9JsbHnrFCzflWLqSFsB5b3CEmEmh+NFrBUrn3sTFFE6BjQL/nYvc0ZJ65yVx
dOCxCIZJHCdvXuWyh/rifMA3pap8ZQFa6pdrjJsIyWDre7cngZKdHKtGQ40PKdtx
eGenXc8Lf5NYUBfAi+4NcjWbrex7ITlYoa5ty3uAgk6vN/4I82fCghKQ7nH05AuI
ZJ0IYr1HwXkxXgFTRJblyGuCpssusnEYw3nPldG+wTvh1e2xkW99yx83MC0scEk+
48vGFDzi9W+20fHxMQ2beF9NMrluygZH1zEqbdZLo6m8pVCftz8j5MgXeyQl76Y4
XzfHm5zqA2vJw87AK7TnvcTKkEVPdXUXbuIPfJs44ZSPdUGO4bT9nFme6qqj/Il0
pjKxX4C3b+xK+UTDzhMRqTM5axJ+ZtUZqVoYPx4b8rPJvFA9TDiu+ynaocfYgLNZ
Cv9k04KTbjA3ZOoGk+amSw==
`protect END_PROTECTED
