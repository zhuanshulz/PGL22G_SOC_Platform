`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BZpPvDFzVdiy3Xqygwy1po3lUTI7FomkivVxb49A8q1LVbdMjpLbUru6b8ueOGr
DxBJK8tjOaH+9BTCm7lBhAxPm2YWpvbjvlHNsxxkm8BXAewSUvDmXvK1JAV09DIZ
NZxru4JZIYmWdQswetXOtNqw4GUyKW0tCKe9W2c5yRhVKeP61afGGb1Np8gTn8HX
eeP6X7V5eXK4fS6aEDQOKHgTAiIQAImd8fw9FzhgBKXqnlQH9hhQ0pUHUb6nJKEp
aae2H21s69ksnUzVrovSqAROQekEDLI3iXtZ+3g3H7ZVX2juZ+bYgdD3RDauIj43
VJaETkswslyykO3R+jDkuJUD7bwPfpng1WxHdlg2buLrCJDrdyAzi0ajhrSD1bXL
GWzmYBsVeMua/8iZhA7zFA==
`protect END_PROTECTED
