`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1hqKY2zgirKHtt7DL2dn+VEHM2JUZqazi0n2lYoMx2Mc6pItcVFNyM633xw5pgfl
0hCkVUoAaxrKewSkex56imd4q2GSBifK3XtwJ8KG49RAi5QYAcTR09pwXj6sE+xW
Q3Y/CMawavjlc86cK7tkdSs/2QmvdHMFj6BCOGFOW5croHMAPGIjzFRgUYrQXO05
k25GJamJVeicmjbBDC+2S+ZcZTcEo1PTEfHTsDHHmrdKzTCaSkbyDCb03QIlMo7O
aia7wK7AIXGWOy+nNzWLK3Ygs79eWQxycYAMMrFxcjjRGX9gvr6D261gaeG1uMfi
g+ZOUW9/HBBabVh5OtK+tu6NvSchGqPFO/JbnfKrOcU5fHtny8Z1swxJYbOxuQ5O
+VpaIUiAbRkYiLGJvS7hm4hfSsrmIiX5jRy2mNkAeBWvGPh4p43CwVWdRjfILFzk
jiwv6yqq0qre1Xo7M/fzEooZGMRsmYez3x4kXhrm/b4iG9RdzoKbNMlzC8zTXFe1
tuOfwjMCf4QKNLa/BtjDNA==
`protect END_PROTECTED
