`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRRY7U5/Bl+cLg9+dlPJndzRo//uTGmw5NMLvw+xnQojYK0Faw1hmLq+32XB7D7s
kD+EBAZkl2NssMFPdF9n4N/rJOTP43YF16+yxCTTjlw2YtgNUL7ygzi6DlvBtixk
KNz7n+sGkS02PyGqHSVrm40W813edziEMlf632f4m1i2V0CD7g551R19tsvhY2cz
1O9f4tZvFcfJmY++216Lck42/lSEP4bUelPWX6m3FvVnoj+2MDZvLTZuDwhBIePi
DfpkSMQm6vuC39qT/jyMUvPPfLOtgsIW+lYiGPN3Nu+nSt951wz3d/NQG8jOAIyD
LC5tKhXyKDM1wEViMBwPk6VsnK2Tte08V4DbKfsCuE0pLsAqRZodkj0Vld8hnI57
srcMLBR4oRaUjxQcIIdgDQVh+uebhrE1nhjWD1mfntPKZmGneCC24ftXV/xGngvj
`protect END_PROTECTED
