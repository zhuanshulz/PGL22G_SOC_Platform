`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ErSUhBTT54q77lZ5X+vfz+dovK65DmB1+1xkc3CNfYqbnVpyc54vcIUMmudWCJ/
laogOvAEo4ZBiMgb2lzegR1LCo01poxJoF4Dfh/lQkHtE4z9g4S4go0ZtOUEmId7
AgbKdgviFTvrwMZIkq6Qlv95qhGg/CjRkalniXMV6t+ZYr99qkYL/DogEBaEoo3c
vot17ZulXKKXy5aYsHcN4fvMDZVN/P4nMhryRmfOdkBipRKXGQaDN3V5hqFeFfss
SMDlYgkSMoCmkvvfwuG0mNtK9o+75UyBzK/BtLFtASwoPFPjdCZa2n8P8AV2NbeW
r5XPY2aWk3lEpUtm1grjHRdA1ohumYDHHG7hRtyfjKvJKcXZOg9IGFrni4iWkTAN
2iFVQjWLBQlEQc1Tpk08llfnhZwbMH9ZGQrSLpuGHP4n6jCzR/NBEfc6c8ynJjZQ
e82CovNbS73yMnS/xHlLemGY7FbR85+mHjZ0XAHav4SB9fTzyh6arDLmXRizBfOJ
UzYB5bO3JqfK9N92gNZ9Nx0WKy8hjDBF/GIdu1NSQtk=
`protect END_PROTECTED
