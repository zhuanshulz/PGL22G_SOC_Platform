`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rbE3ysFbWPqFbv4zEXFXOzdqDT9QibiB+gja532KQRJSGXZTTqTI+Ui1jQoV9Bms
pPs5KZCPgETYdBs+c9x7umu658c7YA+k71qZVOM8uOE+zYRXQgdwsMvvJ/0vM5Pq
CxlELGvaAGxq1GQxgGCr8DUdhNw6mCQgaW+Qv7S4uvNyjxynbRdpRP1N5aUfvIyB
5+6iqCKqan3jY/aeLbGrisppaxk8pvrx12Z6ZZMNg6vLPcy01BwXv86FCZeyiE/B
j+SmSdqh2Z/77+8OwNyrMLGna20ImK3AzN2us1A7Ie689+jYsq1FcK9bdY+1kfUL
BSHlQLBWRg8r9Ag95Y1wPuEqvnefZCynxq8OvDAcUiI9CNGu/DQFJcyyZ0RlGLc3
IJu8sNvlmVNfnwmQJwcWCoIgIDdpeBgQacOTDczxGDOLoHcbHBZuglnO3vPillsb
pXPconiVWWzkwUjoHFEKZwTxnHFdL2CymNI5dE3+PKH3HnSKaCMwZ0nQZsJH5e0j
Ky9i2ohT9BvWbMJJIbFThx+siQKOGRi5jaITu954HRreYYLTHyJu26Xbf5jXhTVh
REBbk03H34UZwh5GXbR87Mf+Vz/4SyBUTN41Rsjg+VO3gnkYifDOss8Nc+bwPnFG
0ejaQwwWltsZxkW8pvCb721I9p6hRLU0561PyBMqIB8QeMG4vyBkYGEzlsX/yJYf
xm97iuCYSEMSynoZ0FK3FFwCeA07m8xjK01q/uByiLBrSZuZVFayCF/ja1Acj7am
Rf/DDCoGBUbSKsye5ikNXTOlPbaCsm4wwzdEk8HVS94w6sCM2POjv4pcr8Pe2f0g
s5q2caJWKroi/+sP9ctp/0qo6tgPSSUC9kIDY8lR7iwo9BPCA0rAzEzSu3Seg7h7
rm38ShC8KyIFCrcxNVwkiNi9Pf4FVxOdPBzufb+/lOmTfSyOAvWGNqaKaiDPD4jX
Ze5EVD45MWo/5U0MU+I1xBY03cGGvVfCi4CmxSIMG3pUl2S4haoVXzEeqhYDXEsy
J4HlVx27aUqzBG8F8Y7usz0Piz1GClCFcMHT9cB80XAQtT/aeFeT1VgXora2QSrB
MKtACisPeqM9ws0US6HqrX+Q8phtFs9QFC6naZHggNm5vN+seusMwl5h2Qm3d7md
sa678s69kotd899Ye+32hS8wlb/ECMcFdVlDKkW35dvgKsPY15QbAr4mio39Kmi5
z1me9BlACsjHpqEhqDVWC5ZFr7svapkw26Jl1D+IOaJ8yWjQdetGHP1FnhMLig3V
w4X9gBu12PB32kJ0bW2q9c0tUQ2ItSxTb+VqOV+ZE08C9Cip76PqtMzu0Px3HU2s
WdFOBij75Oh2H1q64pKQ3IDy6ubRluZ+P4ZbrPQ0krdY+APiaPK6i8UuQkZrYtsm
zhmMe2lpMbTND1Nm6HAnhWTjqjMBS0ysOpzlKR0VfaPlNJRjIuCuzgjJQWZ1ar0K
jsbk+S+PgdwvZo/CHkzRq34pdt/vGMvhcgJnJMQn7gnMzhLW5X6q+w4fUu4ncdQy
zX8SdnERN0VOvE50aprkK2uXYEP60lrJ7nASObZweCH4Azmde/5stCO7MpaMSekE
nTrMruNze0yhE6Vj6UQhkRivMVrX5nPV3CTtl6M/KcuT0FA45g6K6l2xcMVvlkY4
8JEy7VVafYadKQkBbCsAlkYrZSIkunkchZgnZoF6M6XpangSUcuUcfqMa9tvoGtN
K6TB4DlciD+nLUiQDP5vLpBXzvgi8QcloepMHjZv3xYH/u/tFBsXWtyjDo9sH1/A
EiUsxhP8uYHcGcrPoMNtBktox+JBcKQQs7vBoIFCCn9E0Rs4O7BJ+9+gU8XvY1fU
WfG3VQpjtgOIAT5Q8Fzwd1C/zCmgh/Et/EKioLrHx4LZWgewxS1vUk1YwgtNPHt2
aDpoTbf3PIkBBYEtk7aj+WViI5L7CY5xhglEj7wtyX83VlqTI9keowoIz2QG5E+U
+eKPx16imn7n7CI98eh/vKKg1PGE6+WuAYdrGij7ptmDi+YMoAblRjZD104zMGDA
qHw/qdCe7lOB8+Fo0Hxzne17DJEWWwezg50w94ijHmKkTb2B5+xcHj9pDdOfFaJR
8xz2tiOrG+aagzBP1WNb/AzYgA7m13tiu53mqDp0yLsVLgO9lQYzV6AizZqF/sED
Ezx7j08ased2ldxfJLT9H8HXvGLdmoHaSykDxbi1PlpHIuHTnMcgCaKY0PQKdh+s
ygqro1fMa0adDIWNwA9UZ+u5mHVztBSlD9z92QPpRc9AVkKwqyc6rF8OrjeEh05j
5r1UPirIJlhaLO6dqH0CLUFumaGqioXDwEp0MCc3iu0q3XS8uDn/WHpWeixwEWaq
cp6WyBz3e6+T/K6nOZEy+XRtFlPxDEmUq6psPiumlwm0LwHAMkemL9hvqLuKLkFD
RmiG7lWTvyulTzm+g0KNMXlTH87qz307FEb06/DEI2EGKHS1Hj/qPkLb3oYBeAHc
Ziem/8fLvpT0+Jp7JNaEgfcTeDltl6ZC/xObSoy/2iUbFAr78mLyHj/ebcFORNda
KE5Co78rI0kRvUdXbe8r2G2ts7wlKerGJdbT08SKhX22L7wIjMqD1bRwPCYFNJ8p
HeSNJJzCcJnS/HiKHXLeWZy0bhAmGsUQW6RnVgkzVyNsj0EgdNHRxZZgx5yiasqL
WiLgkiz5GLCXdGSli/QqYNcLHJ5tHa/349iE46D7HmNyGSlU0nl4a2CSXw/6IuHn
DX6falkrvw05//mKCWnbGcpDPx/fK9Aw8GvREhiKgAptbnGF5SLrB08JuXgkoXiU
rAL5E7XF5oobHlN+Gu40OLEeYR45olWvRZ7+zP/QXMUYoiAPwov01OHbYl10PU3i
K6yOqKCajyrcSewzPNrZ61STNleq/a0LWFfsnkN5VUgxBkgD1mN3+1m8D10E6VW1
u0mnAW295oxnf6E822S2WD/VL4v5FDSX9rIcbpnqfk1sL3D/AHXeyq56ChgI9kyi
mptelKrx8HeuxWQOAdtQ0B4uPyLrt58/AG3RhrJgPHZJTFOcKUx8LH4pFP9lhsr3
ia654X4azblFKlKrhDnjee2tkWLT/z8O37Ja8Kto6D87glpvhcvEVGTHWJiJp4Mh
RVT/m4gh+/W3OAnWun3f7fIv/r86YoHhaVU9WwM+DHQJLjnNbAs3Sx32/IeOhkhr
AWC+n99zpYSSX6Gdqx9iMW/v4gCzATxgrP+chlC0Qva4vtJNo04fTmpjWUzsc/B2
M7ujow9srqQCwigpT26a7W8IapPDvnyvSIiQjZGKs59NLfpJgqIm07EuoWMwB81+
ygJI2oLKmp5Eq4xlsAcOyO3TYf8v6GhMOchSKmZzrLb/8KaS617xnJ13B3LQMKVi
P6MHYrPrAI7v/cQGrnbhqGYzoEr98l+nnYaFkC46IJ1ZYD2AgDHfxSgiPMmT4Ntm
O4F8zuI7ByCde8Pd4QZU6zmBTG1Tyyn7TDvre5B2xNqk+kmDFKo0PvQ8quqqqoCN
y42a8dkbUJEIv+EcqqN6QI9ueCQCXcvIdVGzVpCLjD6Pi4NnT0TciipWCA7KX6Q1
0qwgLrHSUufGnws3/f25T//5UuzRefXkFZmiUraSf6u+Y0bli7v5Uq1gn8ZiIP1+
wagGiAZVWk++/uPeIhZp6xUAusF9gnF0iewwwHfRKtOJHSUGWzVMSuGkz0fsWMyo
0tfroV6UkofpaYSMz0i8y08dAEYaH7dDgdtB2sFs/bRD7ZAFneIItmw2h31pSpSy
CjZH6rXPrmXnPhdP1CqDHEzxw1wY5pELjew8n1nh9MrDGEPuxIMr2ywmOVHPJxiK
a7qhBl1uFJ/VjbJw9MU4YGCryryBGuVmkeulTrcw0z59/FA3xNy79ucwLw82l7jl
jftdW1qwws5NEaTMbOdveP3KnQEJ69nTd5Gv29ZQ0pKGmW+A3cqbVI5t44vEmSYn
b2HE7sKY8P1SJrQG6pWg4mPmSlkEFU2DxqdPN1IDhifd3SXdYXT+NbThWZSqvU52
+efyBzpkwQ2QW2c0Asa1hbnkNoc47p8usvCaeuCqfpCruhxiEytKlG+wqSirrvfy
3PR8cH9tD5N9OqcBE5SxENLAyUtZ2bbmOLWEXNChBheiMXT6pO0p2AjL7br8rh9G
IRm6YSQZI85hiDlumb7PgxgJ0xK+pTzn19C+jEiZaGx7StNDEN265O6gu9fSd2hF
fFt7iiyuWjuCnBvhiHOAE12W3VpJe2WsmEk8Lez/uwiMCWc/znslkJJQJeQQXe2V
G4/sCM9FhSbH2WYYyunvmDW6/fbuR5LdCfCgVcrArsp+WMGRzEi1T1TzCsSWbNlZ
MkKEsCxbPHOxsOjKGLuRrv0c5GX6w/6/30txqkvZo2Lu9vczI0FP447Enn9Pv8JY
fmybFU2B4zE+5fZn5bhTqYvRORWndr3Ul2GHqvTAKgZyJw2iNCx+N9ivmohVZgRw
nrVj7o/Zlqc9cgkUnqmXIphxnQW/AF8Sj16um6wvoULiDsc2fdC08jL8jwLgItBq
sGERYahlOsAaBFTU4Mjy2gN7GhqE8zoWSs4rtLUJ+j7Wb3HdKCIAb5M1X9e6TugB
Tgys2+S6IRXGdq9iQyyb2ahAWdyc7MYQnYs1PHcdG99cyN/HOZzw5z6AwTZhUT1i
67Lq7Eqv+1KQCIT9tLhyyr+TWFZsUG8kbGk+RF/vtJLl9kS6XbiZzEKRPzFaykTx
gugHTQ1g4kmQ4bUEU7+A98kbGO7tkY6Tajqv1P/JJnJWd6fG3hR9qTil2wPGuhg3
9sE4GwHLlri7+4i4pwFcbGMAMDblMCrLqehxp2LpvGtWJDT6B/6ujErVTZDli5vp
lXxjx/h6QZWrBUCUHHz8Vdr6vTSdVvVxEcY2lsjCnlkBLlPyyiIwUiwf/SVd7tSU
rgtk8kxZe+3N6Uya1l2inR5bmeK8SXi35knY5KOOBBhC8oAqgvRH2wif5xo/Ki5D
WHoy84n1/gq6lj8IaMdpZNMP+EL9Z94l9rQcpHYrjys3abQ/SOdIQ4fojWv7BfmW
/JFEmahDylPzIwhyKIJlKvipcUES2DiYCeo2pFCDqDxneTZmFU8OPsqp6VAPNC1O
F9/cLORutwEaczCEEYFz3esLQq2oZAil9cQz0U15P9JgJBnM7ToDso8dlpMC3Ali
7hxjYlPise6+jjUL33Cr3rnYWhm7JFkzj/0CKBq2Io0vtygVzjAw6RARVmEhM52d
52kot1iDQIj3KMBhkSOw+8yV2QjNFuCdcDxUGNJdVG37PGzLkwcpR5zAoGA6Yw9x
EfY1UoKv4pxaT9WUE8O2KdNVMIYNYcbe4yhU0jAJsNqa3sgjh8uOVeUh5k4rYm0F
LFgrRXe+ia8i1InX2BkNiP/yti8cP5FwTy61ULOzHgmBh6EN760ILCimsq4RQdaT
HuxL1qh9pBl2H9d3wWO9vZ9q8D9NTi3af3wKQcJ4WuH7c370UPxPkg+a+5dC3ebq
7kMBpnMLJHfDhwz1aoPOaw==
`protect END_PROTECTED
