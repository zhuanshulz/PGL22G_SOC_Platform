`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRhhYNM41mIs6qqK97ATtiIpG6nEXEs089QMlw+aErjiVk/0nPra2eaRnT1LOPNt
XcHEzLcXepY70tZ3nVBSKahDXNHGwZMITC+kqGuXl5px9Rpz/DpeplPQ3nh0Bpma
SuCEJJBqgRRAUghIyr44vi/nrONrXbFBv3+Yo5kdtbPxO2RU3qshfR78vjZcw6NL
4URZFpi+VeLHCoru0oGWlJKxxvY6p1uFBLlv2g268J4s57gPEJVDp7NH3MoVx59Y
8Q6IUKlxhg9jVN4qG316GibEFzxteXMPCZLnUXD8o653qFe1HOZtai7e9QU3m2Pp
+20U7f8se+6PmGcq2LF1Kza2VbBFLZ/b8PhxVq+nGU9bRM4/3qgNWwjmXyPUD4eT
phZ+pJN5u3JdNKtHvqjbkmBlgxlIpxTatJ2HuVR36T6uwY7wy9RNlfW5dCdQBNL9
ScFUmqFetj7Gx9oDR/mar75Y5eRNj4bi+trDx1DpYOnG/nwxFA7ruu4mVrEChglA
CbalkvBzVG/Tmkl5O8MOtlipR1FbT7P4Zz0qdMdVUCWefCIffqNxqYa6yM4xHbAr
HSwELBNJywivA2ZUCilTx54a2qNekUqpBT1Rf0DYyNYa5UKBdZCQcJm4CtPibOpv
wmSjxojLyA1eq3Gjv00Gza6mGiD9sRzvyFNLmYFjNLdrCqz/ufuGc8XOR4BNsOO9
psvWk/16cCpQauN8DLgAZSdPq1burCow8o+hepnk4o522vn/s/a76mE7MZrmJ/Kr
93sdCeVChP19LTbZbR73RxItDDEKkByD0ChJ/xIFJHjfafD5m1sDfflTqz1Dhc9x
dNQ9gD/zEv12VHcQzkjiZ0kojirYq+qXcp/jVTii55mDx+2qC7QSqKLMJiPxRlt4
wpiUduy1g30JuUY5op8mPThsc68tqTIWTEKSUFBlwE/VQunMUksoBp9OFHmK9Efv
yd808LC6inEVzB1BURg+wKqXhfkSyAgTFZuCcqqxfzmgG/G5dZ3L16QvAxmclICH
MXpopLKTQfnfMJB0cJ1utQ2jdC0R6kMLLR58WA169bDUv0HTrHF66ivVJPPzfTB4
lQ5x4CR1uKEgLCj0jTwBUD2ceDQQ5VjostRvAmCGwxtr13ElLS3tMhKsVqSvmzEl
caSs3luKGoUgRvFXRjEh5AsJG7qBELcHQFce4hstEjhh3Ag2eredRHs7UxliUAd1
7k1XJA+VoqAVrKsSsMSJtvJUChZarrXPPdXZQANFl6jqRjZ1GoPyDm1GPCMKDovi
ztsjIzqaL12EOJnm9Rc3/L/xoLD92gLadUMhVGUHu6E=
`protect END_PROTECTED
