`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/vQY4tx5EmPAsHSbqdn+Gm+w9kulpFeaRvuD2yoJ52ngA+U4BtDrPHZfcMh014Ij
J2G/E1r7u6ZTEru0sFJa7bmic2VBM/v6U9D9IUCe+b7B6DvrGWXuqcideGasqmtt
L/bkcsooEKb5bzSYPebjtabrJM4Dvu6F2hxZbkuV7v2j1EjvqAvtEpwbGz7ctiZn
5SIHpF/MZEwxTeKBsbpUrQSI8W3dFsjSZOYCRUwXVl91ExntsereeUHYN+GP5t57
GbnnNkZft/ns+N4+oaQU726gtfapCoGGVYOMHcoSuR9KWkZmHz2rXbeVnG35MkxI
viFm5EATbyByL5N5ggMOYXk7iRmRurUWxj8hnL6oXI+ch4ulKXN6nMRZAQxSl+g5
MUtDwr+XLg+PZW8yNchem7uxbRnbZO+U4Oqnv38eB0UYLFEW16ViVO1eJesoZVOJ
5pQ4P+MquEIz++12vQ5Bq8FWfefCxtwXEoXnWn2aukfqXo8ianGvUXmIGlEg70AP
yXQFwaD9GXugsrciGPtyDdbgVx12fTPlEAvf0gi2qvwV/3UMdtafVJ6SsSutiPGI
6oHMEO2DY4G4cv/WQKMOUTJ+wOqIT4O897bm1dingKh7uh0i/1AiLWfOtSv2+JWP
kr922NyxLopQTUo3OdTpsbYkYuNxIpTBM9sYH5mjaZk9JvzMmyMmtlHiw6uKzDI5
1YgSUQZJttBvHFy5DLnid+iCWKDz27/2pUtcETD+ls/2/hf+PHQ+3xh/3DPHPT7x
4XQ/D6B7usrC7/Wu5OttsDGcUVnTyUW2/XDGNDxkQXZE9DHdg/Hm/0Pk7aSX/M6S
0Jn32q/OY8e2s5B4Hd1JCwjs9PJDwo3oBdooCvJ7Hvy+0XE/nzA366Z54Wrbd6e7
rPV2VZ3hcnLT5H1bjlBb2KlphSdwTBNnzV5qbND6gOWLYtrPSAgaDiEXR4bMtds7
o07G9Q5YOO2Kcb09i7ytUfhnRcPKoB3GuTnB3MB1jzqwRYo+lC7syfc6sFiu9gHj
oLkaUd00nVjl9I5SqHPBBOGptik/j+xWzy7kNZfqcdS2oJBt1/B5iPzwLX7gO/NO
vn5/LNnUwhSh4N6/Rjs7h6esaP/D+LCQGr772P3B8GIs1KxLn7W7JLpKn9jIQew+
o7eyr4QA0dFBrT13ZJL9K+1gcLyZJghu0ofVbNmI5CEGUSx1nTlz8ChaR44eFtQC
yevSO72Xi2Ru4sLGYcfbLzLOlZFnnpA0k04LSY7vdken6Ut5PzNDuhy4cdhvVRBY
oIke8peDv6AwEA2EZjetCVvmxGTyN+n1IFRt4RRLRaz5d+t/8V3EqqZm3RN1nmNk
oNBWOpyaymGSAOzLBc4feQQrbaqRKdZwu0yFOTrMNDntHqqUGgK59APy473sBUGR
0PI5hP8QmqlcUQ/SOeixYzSphiZLksin1+RM+G5bi3ltYQM36eNfcgnX3VU9VP9t
LfSEgSX6cx7atbH4mnHT79O3edaSWvC86kXqv7lZZvCjflTE9/6Z18vHgp5rRLLg
+hjhijnqbqMnPeGBa44FGdi3d0FuIG/dxxURtQMb0eDOdfeVaIjkB8vmVjr8jkUS
r7qnhfxEocXCUtZu9o/T5gNrnQ5obFkNbJ0zc6+gXmbQsBPU8YbibHGV22P59IGs
fnyk9EoUaVcWrrWwB8LD/s/4u0rHIUDVAQx8/fGKATR3bHLm23PIwZwuoENydmZ9
IEbsczBpJsYEJ9NlHNOcCUXbVuNaKZ2D+Z2K1Colo08IyA0qPesjpl8lQDSreDEC
F7yzJnV/8OIPBPVllotIBlBrTK/UUEIOFJM4rU302tgipCFUQr7V2K19MxBbWitB
94n2aG7vg3wSunT4SDoMCV1hMEGfJ2ylbx/DRvs0gghNPt3AjxwkZP0VSbMHAf8Q
Se54e3fwtaxSqk3RVUQnwzQ+2EiExnvC80fLax0kAh7YCfZ5OkUu7Wb9e3o9M3Dq
7hsX4TRYSw6mRIQkz4R00iMNemPLX/X/Qjg+onfJNJQVuZtgIpzWOh3Ze6W9Yg4/
ucVADn+w4Yk7C7M0koRt4GVuYs76bABV4emXqykHsfng2uMzikSqPKGgVAK/KRx8
EAaHn8NbOaZFsx9mRCAki2DI0ZoEhuQZPy+78Z5DA0rHZqrYkGfGbCpNpxP/m9Ku
KFwg8WzFwJ3HNChDQRqF6XpVNR/jNRpRp34Pep6JyFkfLWhv+TDIhtxUZ0Z6DcOy
fXDIL/kONXYsRCuf0jXWUWnIK9FGqH2HzsxTkDcrrkDNBy1olwOebpIMd3EwNFSF
yDa9gYZ5lXpqybFiqE4Ado5BpUU4Q4dLj9zUTk58nZzZbTeYjvEfMKlsEqBEEGkE
x3RSUTW2Q9E9GjZKOfbVMF0piCh67XHN2CoUe9GkOy6/Y7Gok4RRmCmG7ZiNQ/bs
IatHR0sG9NicExxtU+1PMfVjqzjm7JlXzYdeKnV2LV2ZcwiaW8ZrGIsAS+4SSzHS
64QKI14Z00np62ueIPWawLgGsrUjoIjD9T2h/XwPnNX94aDPCfSAns4jUg7XvYho
3Iq3GSfyW+0LgIvk8BhYJriCt9KRfjDQFHedxDCfvLx6v8rHhJUTLzF7gzbwVHG1
jm1CtJfn8K9+3qaJvmBu37ChHaENeiL9xfrDK6VnE/flVGPh+zI6J9e4Ehw7uY31
roSbw71bSvfvKq+SyAkIqu64nWjxkXnM9lgQ87HGhb2DBglqBuDR3QSnMqXib3PR
t81FcsufbuDRlx2ubRIn8V3XHu103lvxB617/+FIpu7BcPbXpgdiAiODSX0zzDQW
kgBJUP9iEyDf4L3CssdRYLuHIygMlZBqEWCCJgIHHmYlqmhp7ZoQq56V7leJqEjg
vo4T/nGttHFnUd0ISTlQzEzjHmNAykcXC8J/PTVnRiTweQMh6RM3ZMGB88pB5MV+
APhmStOFyxAOvT7lNw1RSacsGjEFFf+oTXlCttUX1q5LkzBd/3tV0N/AqVJgc/2P
uIvp/QOpHDlvbZCkm/W81uDlp+gOK1euCkYeZwuWchfWpi3/6VTQg2WD2FNQCCzc
IoMV8pVQ4vUPEyVp4lToucBVJ51DfZn0NGjJQCSR+3zus6WTqFKnPyZq1uju/xNi
56I+J98YTjNosKXdDaQr5Apfb+pzfNyI2ooXDEVB9rseJJyqIF96uOf42zY8b/2N
iY52l7zVzhpLxEgtejwAnMwTJPN9ceYT2F1qixZNI2MeM9UFrY3mO6VJGFSHl5FC
2eHWizlAiqYKdTmsjaSOxRL2leFJz2+ib5Ivqha29j1VypiNslE1RjuRQrVCO/k4
zYnMLev5M+nY7t9fCS+hU67513yXK6mNOL3oZj2Zc65f7St1roWFMKf8bSIx+VDv
xmImbCYwPZtlTdSvYbjJRQK2qANrMQpyPEU8dqfqvWnCw3p04YM2Wbo2hIy8o16I
lrGLZMsfqk+BxlR91ZBxavB5vFWgJ1GobXapfRkTdlxMdSorj2AHd95+fxtr8tNn
r1vqA2lO2Mvz0hI+IqXWPu9L49xbaDdV4bw6Yt4bxd5QHubC5qZZB+hLeNpzHPh0
hB5q+WVgQX/cQUsZFWsf1SWrlO3UWLaFgR/teVOjiUwv1sakwGHOTVe7TuYBXURb
TAElKmfss51kUdjm6PRFPOEwUE39P2vt5/1eLe5rOos+/QFiG/CriHoGwZz8W4EE
26dM94/RUxJoWM5H01KnMTXC6y1kh5mnZrr2lhzN/jt2sAf84qhCPUNHod1TWNTt
bFc36N1QLJtqmxGDF8tuLQ7KiPAEKOY36Rap+XRKmJjvS83OzJXsiD7WlX3jqBJR
NbMI+1MCfz3aJrqUgqpqQFXu37zyLIRUHQ5JyyBqQ8YkYz2eN747fEHtiCNUaRtg
sAL/iwgP0CrbUR2pB+0KXY62VWtfvbCZYKKFR7TsXoItttpyU3ev7lqQnG0pdvux
6FsnkzgxE3EbpxahuiabiMF1OPx9Rw9EFbLFl87fAl2QNslL/OlEmSClx/cxMGsS
HEGBeudmSR7usIAuQIEbJTplEeuUuQIktm9EoW2BtsnPt7iBBANV/lSrGynfQAe/
MU+0Y0IyVi9ZqEEW3Xnhpcdp2aufRJcUUlUoh7/Brh3YtI5AP+E0uXbqM5krobi8
AC93zbHLOMQ+m3McpSL9+zDWsqeq+sGLAKKQXjnujW4wLUMVtLGM+CGaJkY07bP+
CvB7VDiAylXr2DhfNJdcUgYPXpP8/b8jQzOvzELEk8KWGSo24/SKpayDtilMV7LF
7hSrz6uQVT/QUZX5tn/A0oZsywEonTP48cug0y+N7jH60lEwnERJB2H2dZXPra9M
hqvTaHDXqHdPIN0X9xMIQU+ymMENX6Uq0N1ICkCzX+ZyruEy9fcbA36wShnnhdGY
IlVM/bIISlejhu9nEW4Y8tbPmJFbj7KIfgLo1RkhDUQ4M3eAEMaagUZOFab/X9Zl
C/q2WTVIcLqFDuYMBoCyV61hzXEnL/n+nevh6RYBOnqV2FolRjRmYVmiORnQQJeJ
b0kA0cOjgaXg1lgvvgaBqwgc3SKLBKrHK18/37EpFF5kQeFZhx/EqSOv/zujufig
dpmHOEyxjFCgSarQZfuoxMlBb7PX5tsr08K0R1jKoP8Te57sDj5tq454tLlSArJ9
f4I3r4gK3k3yOtYYmtGFsMhwN7oV6z5AYmbDfxunbU6TYGDmw2x886AAfY+m6JE2
eLPPKEjnwY1CfGsBmbQpW3MIvwXJNOk1N5usonmbvK2BVka+zDkY5kZQHx45TWwf
AcBkdZ6iRpZAgeTxCV7UHs0mmTnap19pavZT8xOMzV3R+MycyuGPm41qu4XepmcS
ubaMV7NV2rCzA6K0W2udUnu5wv1FInVHquBbaNXXNTAaZuNqwnhO4MKjnDAihMRC
xua38o9/S2qkeb7qdD3p/tSEtg7zlPI/4/OHoXWrLISHKBmW1aLPGiILYAf+vta3
cmFOFrWqKZNxwcLhys0YaykrT03p5a4cYtOdxKsMS8uoOdKTvKvg1m36BHiwS6f5
+FUbE1Qmg9o34pDwqEhAJI+6KwP+6tWArJmpPRrWPC4f9LOdftff3mSs6aV+obz1
oXC72PIczZKyydFVXNqPQXhJp0JNxJB3N65KdUOqRZI6gRX+LlTzj6Bjtfc/xWLy
C8fXozyBNXm5YVpxeaVt0fw8FaizEQ8gCQXmKXKzf4M4jOGSH6/apmxAMCSrk1u2
NVBaEXK0iLNdn3sPdiBb5uOimSoht1gXduvptV+R+KTt9abv696v/jA0KVJRHdYi
yXWygBe1TKtnScJs83ESkbLiChdTEkb44xOy9lJfAeVambDUJH95zzRT2NmBC+5a
IjFNv3UlfesTSHxYFgI9I8coNIsNyQXxMt9ICW03o6M1MyrEzEbRr/09/Oq5lqon
eDy+hmogiDvhfd9yvQAq648AMWDq0RvTgRnTtlf9MZEHROir5vqnr4l2D6FI6Tfd
XWNGgIAQpHVIf5uTH+sxiaB9WCqBDBq6/ocKY4aixZcCXUdwZzXYJAR90zGKLVAJ
QjN5u3cijF5paNINmBOYKQvL0g5ga4nKMAhBzNUUe2wCjU7bxmUb1nXEboi3Zfnr
Mo6/TTCM3MLNAG6xk80FU7uiz2HpKCaKdMgx4js4w2IHa4Ea9I7zXy8WMLGx8B3c
o4fb4xUGvr+IOyLHUXshZoU3kykOII4fgx8WuKXF1hJi7wif2OvzoyLpuXP2holO
SSfnrnb7bKV68ITJkEiJpQf8l/ZnAS8sKNBdMZGSCzJYUtnjbA4gtAl/Mt+ZoY/W
3hqDMrT1lGLrfEFx6aHPWabsu9k741EHxe7Gu9QOFoSslOrh9E6+jkjjgJKe20VY
kb13QI4fpogGmLpCdzqiQ9kJE8HXONip3uXslS+kyqLfWwNQabFohlvjJ8zPD6Yx
boGZCLvwTIYyjUytgVfKN9hn/3/bNdfVOclZ5Mi1RkQ3gytHqHGuAGwk8iBYeCnS
JV75e4XZsoQOBXs0X5b+8gB4WlOJphz1fIKOBgtxjZImtJEWzUIIbFAU5ntqcly2
AVzWTlmq31Nb4uSwATpBPJ1ej89dVJ5YJ4dEeiL9jt978taZ7mJd2CF5qfUNeRdn
vlxnJ5RtSG1hJCjZLkwBZkTjTBSQJItKUliOgPHuqjp9DTFpk8LRTqxD1ylJY8uy
LNOAkYlxTISM0+XGcKobkccbJPnCe7Ij4jLRB1ReIn9iUYUJ5ae5dexTmNnR2Qtt
LDjmpzpPtDZ0xE1FodC/8bjsR5IDDquVwdZm7MQqjpYmPo1zvmv8gpPkntixYYqV
/mu55BxlWfrrYIHgkGQM5qf9dzGIe8JZQmwCBMm/Qw7156S90Ko+Nk46K4XsPJAE
wGFlk5Xu616G/bk3unE6H/+X6iWfV9ZmMcMqnI4oV8MtAMgfKPz8grfZ5Tar7ZG9
ZWAyTkTgEuV80o+uOIwoGkMPr4YzEBQ3CqXtrLJYgn6WFLHupX/6lnl7iRaje3RI
PLfn14po4pufCt6FOiNrw+QaI5OCZroSaH/4t016w0Z/+EX99p4oh9KNmVRWLqPQ
7y2ancntSqfKheO+00+7lmEQTzL8NJNpVeNLi/kt/VDhvbJ51NwM7i+W9wyfy0xu
jhM09UhKr+AldxXfaMVwoflyripzXNfiPo0T33Tpa4ULbz3UEvV83DTICl6hhkhM
Ryo4ECp+NUJw8zPG7+hmgWK2qtQenWMNskNQwUVf/PMG4b//4crJn/4CAL4yUjsN
oE3fM52/dJ5gFflqAhcqrWgyhwDDbf+ET+LJhMoAFyrR6hVtxoeQ5JdrpznonQ1p
zo69jgut0DVUZPX8kRuq2uSq2CvJptwRafBNY//e7SOqalXwOOvZNZ8yhVuxaEoC
d0BNu7ghgX9RC9YFf4vvLgJA8pZ3kZp23SP6Jk6nKR6q533MFYCD8WgKsWvi9yKD
Vrb3lgLmhs97b08wPIqzpo4EwSoOSP/ut3ds8O3HOfbZ6QBzIGGEkC2rx3dk2hSJ
4O2/GMZMefHIsIlpaurTbOMZOl6XVEE8OHaictCWXW+MFAliDM290RMYWdbg7izZ
C3RvOZ3EHkNgqXRhJz58FVZsbBsrZeLv5siwSdVjEVEguqc7lljYaYsTM7ouMToV
AWoieCO0bM6IVZOhkPZmTuc14n/i9cpzljmlhuDBxe0CspH7DXUSv0c/Z7TWP1rQ
BvrE0DWmvJyB9zvia6/RBaDjQtZ3mx/oIuECrKjaBLX+OjQHBHDDlDrUm+Sx9x3c
Bbv7NMKY+wOXlROcs6QB9PLEIpPbZvxFMkFyGy112Atxr3LGkMLaf77vBZNlpSII
x6c5q0Z7BtP9j7tInXtzggFh/VYP3DJChZ4Lm2J1EW3cjVklKdKGUZCUSILCwrKM
e4nSc4TKyK/fcMXa2DbzA7Slv/PZPkCJrc6OcHVAPs0Z64gwAJybGh3Iwr8f8zed
fllAnvsfbXnHKqHyRCT+mp3Kp3/vsywTSSbXwEk0EOg9jICNM/Vz/Z1SxDPWXbNZ
AnwIq8yNUTOEQlnDCtgImHQmoE7uRgrF3jqrK8NwU+k9CKA9DvkwOq43t4UDlv5t
iJcjOG9B8vyLq7L7rKZiG4qlMj7Zs12DiQkSTVUD24jUpp/93BO0L5eMwzqwcqDQ
rvnsUHTx807Xw1aCh6bfCf8o1XS8+23uPCo91NlrLHxixxQbwTsF+SdTP/4Y5mar
Zw6JHIW6gUiT6quD2VyqQAGm2gtdUUL5lB1Yngs4bnFWOS+gKagLuG+VpYVR5Bxg
Y3IT2Ks3yaC9p9JRbFk56C0ZrGezucZovxH6FXG4fzJeL+xDyVOLxrQvq0Yw115/
6V191sFzLBezQyOvEM3qrxlVl2QUxB9Iln25ErC8LRT1gYJO0EFPWIfAo4+uoDKP
phbtTlU+kYkT7WwN4BhugBxCRbJ1wZTCJnLzc2JxnpsUtS+tl3cD/HmhOljmh4AE
wr+sfppNHjasb0lIS3P3aiITBM/l7oCz7w6bzRKvVxdJW9yRAHEux60leJYQD7/b
SqlaGrRL7n7UPMZL8wu2g3mm5t9cKqR20T3fefjoByAJzcngwB9n2Sp12EQQk6DS
grha9YTJke0NRxU/UZy6RZF+d6WSarmHxc7rYt7ANI+6J361DL3y9zaUQf0xUMNn
K2eZzcgA0G+UwofoVzxQv4oOEmY39RfASR2hw8JsuCahckjytZzwr1BJC6wbAqli
ll22LoaNuhpHlczyBh36hxuGZOVfKaTNk2eS/gLhrWiO9ax5vLkj2VTTAtfBcwP2
d6NCff4MZBXw+RdAvAjPxDXIt3fCcT6dKdF0vYxcVSIzgX+3BEUmMkn0T4qL5ExZ
ZCX01Me2Gf7XoETBd88e7yeM5S/4m3OQM+cz4WFKT1DyaihcIbYfAXd846BXabO3
4+hsiNTpraZ4enQARxcxjEbJ1x1E8+jTMmhlc0LR2vdvoUJDRCp0Lpf4G9Lv9roK
y0ZpvZZ599SgMCf0vPGzgIkg/hBANWsqOadmlqYsNdgymyncAdqWaGeArJGhkysY
ITdcqGmVgbO2z3hrGUWcjSiQsiiWlpGKalrh8TbY+D21NUNCkcV6XIWChZNgP5kW
CsxpKVIF1SDim7UsMsVRJy9Mj1aF4BTHrPwsiSmEPG+cuSn+TjwLBNkbqRVbe//4
aht9xOB9ObzENFDesRss88IWLlHjKBCvLUezezV2YXrl/WMahgXF3IABHIHt/qun
JcM5+B8dOeFGYEzopuEO/BUFBIAvuUDukmYOc8tbbj0qGQJ55d9FxNNCq7DnLDzR
0flxPiuFj+mvo3dBHgwf08NALV9dFUoQEGdSX+VVCMt13XY1E5+mFVU5bUrEXzBy
wx6a/E/UrOrzc1N9aNsUkDNZtlF6lhDxInH3g8sa62tzc0vdN3xCGXsmQ3r6vf7v
3JQZO+mvBtREfxPyEZK4/sHBour9S/6F2M7csPvMPM8UwDwhjLJ/mLj0aF6kR/yY
nS0BflDK9+R1uCBpgVd4j25Y3aKKeuNE8ZAMqSjUW0qWBRZn3pnxj4oziII8Jgsr
sHeHy3tvG7quRN5MZe1H2eFG42dS/3qHF6KI9BBRCYRlnHkHwng0Q1gGuwZYmiKc
i3wMFinlF/PqULRbDmNRyn4uLEXiwifoV2ujQdMiuJVWw/r6qiPzGRhOlHExFfv4
foJFCkMlg7e5NVkO3bY5z2ROuX65xVKlzG/woTK9jyD3mYUo+wsNdkF+NY3GbtXI
BM0v6QbpW9r0GB68xxtiJ1YQUqHGZ7jLtS04pLQZtYkCA5C1ikp/kz2YDMj6tDEA
DJiEGa84g06qZhjncxOf4t8jzdIY3FcMq2r7hIqElprNjn3sxZYssu4+yoif6JCW
h/cpo7/GJJhna3c2TQEAEaLykGb54Y7XsRszHK9QkHW9vUAVvXBIZx0FrJnlZIuU
WrrSJtdfpeZr45F6wcoSDqB6LStjw+jYqJnJ2Fao2DFjUiS2jDlbPB+VNlc7Xtc2
3IvUJKYz/LSDy3CyFoZtt3Wy8DmnOeByyCcXTHsmCM4gcozHYVTjRiBEjvAbgNNu
SkB8/tUoeWFVpgliFwz7Q24vnfDww7cjuScevLo4YZc2kuMM4NyTfX1Z/uj7+bF7
G/fC5BbIajjR4pYEvBFQGRohNmsPF2BOoC4dW8Qa2yStu0aZ4zhiJPERrMEo/X08
9MmnyuSmbwxNAww1dMo3NuX1nzOnzlKesnCCaedTXbabNBafIMMNZHep722rMK0V
2bMatBqP9h4NHVqVOAbLDEidww645GhkB+c2d1X7oR7zWPRssF3pS4eo/whB9l3e
g+9m6RLmaoTbi2edicd/E1N22p2veggY3xytb70iC5o/Bz2Y6ktldPOg+kIFL2q5
CExXDskQ1hEmM5h+owVuF5/8RRloSUlbcl4SmrJU7if5fzLcDS5vXMnJxi2OT6Xj
mOFcnKqQaz701a2UYmCVz5L1q0Nd21s42XcCy25SIMhQWlBniYKUcy9YJEU2mBUT
lzPLcP3T7OvEvVtaXgcAo07lvghe0Wx8MX5xyNW9wpFWiEA+kIQvL//2PvB/ajDG
bN1fV1I8CCU+4n0U2PDOH2xka3lTbEedygQcZE4Gj3zJ00vw9DvLOdWkbdllhuiQ
1hmUGwtClzrDXTeao5xR9XfPy2lCyoedhIVOg9FKJkcU2mAbtUqnBwhIlZoiBhbu
WvpW8SBHHJwRxNHVsD7cOwSkQk4bwsPAZm9H/xdSNTsoeFfqgZU4pVXo8LXy/2vP
`protect END_PROTECTED
