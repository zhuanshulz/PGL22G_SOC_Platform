`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DCy8zYLkiuN6Pgw+Y5dDlzAyIBui05s52F5gmiuh+bMcvVzLYxgXVkW9PiAWKE7B
UGLfbgRJUjkC2PTVItkSLdiLWMV4QUiINy0PMIwVGwakiKatIot2dwwm8dFM8mys
V2Ln+9cTJbI31ol6uZubcIIHB/TfU+6bEScaxWwxjALpIky2J4H/QxXGdMVEgJl+
w/3L71FAD3VtjyGlE/CK799wO76ktF3fWRa7SpQYci431emFVAXK/1zHfSLVLfhW
9L2d3lID/PkBpaNd/pwtd3rKNx77h5Tw0trSFDgxm+ANRaiQIaGoFQyqKz9B/hPE
twWZdR/2OgoWZ6wN4nHcn9Vw4YR/Uh1U1YipxFxdhgh707OUQGW1WXmBAbLrjS71
tBPCveOAU5dfgqoNmNQ2uXaYw9lzPXRwEE3BTZD6v1Z4NlR//Pq45A4naFlvWC2U
F3ztOyRA5K48sLSgRubAyA==
`protect END_PROTECTED
