`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HP377rHcCyzowa6r2tXMYrUuwsjPq8XyheK9sl3OodfdW9WKYJoC8n9ZYIaWC8d
IXpZ316h4f6JRcbIhspTz4WVPLCkBYWACrffZX7E40P8RZEc4EcpOMq0/AUODVgJ
EY2tW9340/HHDqlxMyGu9/SbmLYq8Ue7LjNFXssmq4EPm/fFE4eYpqmzulG7SAcr
+VDH0HfKx7eVhZyiJ5YyBu+FKCrpFFojdPfMnDvjWvQ2dTD8MaDEDphOY46sxaPZ
WQbqejY6Di/7NT+LfGfkD3irg2OVXC6Pk4n9iL51X9aiwo9m+RRkmzRuSwverA25
k3MwCAN/dIdDwfgGshTbwcQ/PHtFZHVw+thUdJmowxbYJELRKozdAOireqOum576
nqsZf0HlehnzSSWb5u6FpO+w1CyBpHr9Sk7L/frd8LF/Y+TilsiF3VRoQVzVztJV
SpHKDoSL9JEFKsgcQkV6oknStCLSHxQZxWQnkph+NrtWrV9ZMP037aiAOlxG/p/t
rao3RUbHfZsecJISm2XXnw==
`protect END_PROTECTED
