`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9rQF7HZYjkgAq0NkW5N3UQZG1j5uGYtFKREi/gI2Bv/QYTutP33R5c6WEy5gQvI
/VaR9CYn6qBD/dOTH1j58WSCFdmXj6w55wvjurFwZ9Fuam85/3vAYhUREZl1aRQ9
NmBDDEA2g5paaLNEJI2DT3U0QuGN5DRgkKsx5E48z9KwCm5xv9vgQlM9Zpq7ZVt6
rU2FNsG2HyeKXmUw/w2JJv1Yeigz4QkwXK8foSDQ9XtG2NEVHm+UeHlIPcf+7k0J
K72lkBsjiq7agmGIBd+O7xxsnXMb33yjYfWHX0+ZML+0QSRmYa5ybdH57TdMzilk
fCvgpOfEIMO0zUQ+hfDulvGYDhZGYiHSpESk2xd7odlH/JI9PIHnMjblXwrNVb/+
QaORnhWc6gvMxVoK8SX+cPUDkVuR9GIX/XR8OqkQYtcqJfTqwdJ6TiPCgh3TZ3Ne
0SUO88WrLKG/MYEd/c8LSZ3ZNz2hmLeSwrM0tjc1qj7RTiJZBHYmo9WWMqMVNooc
Ll9Sjtp6HNyqdR7fkMMO/vxx3IhurJVNa1Lt3aECjx+hJov4giozEPeI7g6IScjH
7ObEvJ87SZkQ5fQA/iRtc9kzLHwKRrUN4bNHL2iHOgx0hYTTNYaixQX0rw40NivM
GJrS7ngxrzzpExFiiXTVQe/gd2bf20YIky7ezVvt1fDpsgzdYecZPEG5Urqhf2+y
`protect END_PROTECTED
