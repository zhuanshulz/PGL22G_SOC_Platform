`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82m+EbVkb4bworoCQJc47P5+bwKUynLDGXzpldIctV2UiwuHRojI1URgLQtGM03k
Q6eYa12DagA2U2gzlPGV3xuqCCfgVkoky7NfHV5+MiYInUhdr3t3fmjHDZBqPuXk
e52oEbShRAE97WDpx7p5kAu+eZbd18hS+kuKOCbe37psZHD1qH/3RXPb1NcH9x2P
KV26t0Ma1q93+DRj5fQLIwAkUXygvHEtpu9EuxMdqS+twZ0C3P0btG3FC9rVrYcl
N4lQPJHbX8ut6mqNrgx1RkDCgYR3iHh3pV4X9JjpIaNBmboAVfVgrpb7kxmtZfZH
YQ5SKCyn3pgU9GtuZ0BQQoDUZ32lHuZGboHEEUf999xsJha8osxjNcYK8xwzA3SS
4jqIkPg9XURyRHGZX8U+WK7QdDEff9xwNAoEryOzmPA3f4tPWKGI0j7693UpKRMv
XVmfdsOUwZe3ygpbxLZCBCDo0JQTGtYLdXEsQMZFejgX7y6kCiEEAt7fj7nyyAbl
m6TG3C3F8eMHVZ95TixPUKJWJuviyJF6gzmVGKQH9W42y9IWpoDEPGTB+O6yBqKh
tqPlWNs4DB6pIn6WMFcb0rnk2/5e7SZFX0l7sz+HS98byYvV3UlakHECQOb94f+R
qJFyezSO0OiORk3A0raD6XZaLdcHCTejb0aHVNkb59QKcqEayc42Q5Jd8Iqqlgjk
P0dTGgGLqslf7NoMMkBNtGNLb1FulqEqRB/mSba4EZRNaGPJNRY1qQFajeSdIkNN
yIRhWnEL4KQobPjrJVlMgLJZkymFZZcKPGBUaXr0iJTao7i9XTFjjxmcNoPi+r2I
DKht2ajrdXRh4a7bxTBCSm06XK53s9jeLAsWzX7nOk1dfYGFivwGlz0l9flP9t69
b5iG2TJms4zxogFxQTM3R2WQvfKkcqDdByEwKwmUHEIXaeETsv0ySSky20eo73wT
grZbWwBiouvX8SdoqrasmYacnA3pqdjzxVIuYqjErjbx2D9yE1AU2J7C0hp8kqga
3cReiCXAyqIA0lI63Y5LIYgqOSaX3BjAHkBcsJDzJBrJ598rfdjL+HKwYKxfOBFP
RqZYpoAmJSWaFFnVacrzMQ==
`protect END_PROTECTED
