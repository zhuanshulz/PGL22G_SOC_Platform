`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tA3flwpKL68laFYOK64XimIM9MBBCgxYcnyNs5v5x2ngr3bQMa2Yfwv9z1wcxuyc
3pOYd9s9V/QLL7VbI1pMqky2YZaxzuVG+qSO8zyD2vb8qo88pSuD3XEgOGq9iIw6
AtKXbcNQM9Qn7F/Vv6RO8Xuw4X9hOuAVuLNL5Bds5Hjkrl0OHWMk0vVY69Izj9s6
X8wV1CfMKbxVC7AGBkMARscRdNeoT5RwcQ1Lhb5rCeE3A8HWYPQwMMSSyayqnYsM
g9Po3yt7J+FXzMRthPQTABUZT5zvilOGn/8O3GaWFUfxI2UZ+cYkzrLUolg7kG0/
i5pZhaOV2aTq3hlZjIc9yBCUAz5RFhIyqTekjwj0a6zYqx13LIs2VDUh7ud2szXs
hHICUaS7qzcTf32lhBDo1G/JepF6RXDIWIU9wKTJo5OlX/ZDrcpvfgVtkOuFJixZ
59CoNr6m8u4YZ3P+j5NpBejOnFts9qH4a4Zm8BhePJyA6Rf2H3ZTKfYo8HxP2VgW
7Xddx0UXKw+FTQg5nvYmTO4epRet9FBx5nVLtBFyqU1b6Ob5mKlce3EfwOnDwKnD
dN/ih8JAtxcU97Vm+92gOGfhH82OwQOPYazQE129GUWofmdw0UxQ3W8lMNVgYphX
pnPnph8rLBMkjXK4u/vIS4VZQOhfWd7inYuhIfuLbeba8o0QaAXEoun5H/PrKAnG
6nvWbYoTzBE0Rfb7LyUWa+/eXto9RugxnGs33jhrjbRumz1k14Uj5PoMOd7QUVcA
z+9rDFEMDYWhJtkNTZsErMjAQeAv8slk0dM7nUrIEzlX8VrqmRyjz4DeOxtCWx3l
XuumgPV+bBRiiyo6BRwCC7LKguaPe+mKg6I82CRn3FOOVFDRphDbm37AIh5QgVtj
ce/JrEyVfZpYqd+7AByDB92wytnDuygtWGhwH73IYvR8EQ2DjG2y3ZQ+BrwBbs6y
cpgG5MiU8APGeRQCvuO6ds1p25Ew/SOzoOn+ephS1XEQxwWlacmQfV2TdDLlb+39
sDKa/2cHzXqnmvjH8H4zDlBCwFw7NzyI9RPoBU/Fyiy7W9a8xBWf3MYrtbm1C0Jy
TXpEfiVmWJ/Xj0ntzFZPnfanqnipgNL/f0VZPjx6zADi8x045p0hXgdEd0Raz06C
kd40zCXCnVOkVvkkKysiXYlNisyer/CI6aCwCXlmOLVBP1DlPbefNsgRZQ5/hNKl
RZ5Nid7bIq1vkzUk/1Ap+wFOm0KyqlrL9WfO6XE2lVNDk0oyHQfHzzZkXSOB3yCR
O75dQbHXw/7ytPGLVJxwxtRWClEWaagjoLmTZv3YBsjqeaTYwNHN6UCf1WpEzcuM
ruzj69E7T89nUl7rgRclEEi61T4Mdqy+1PJjP1PQvPdqMA5hjJIzV73LNkBy55mT
VZmfu8PNAHGsMcI75Sh6sASjCfIpQT0lnINPqciejrSGqTvf7/hssrcqua4VcQPz
Ekdiew3AkVTtoPlbOmEQE8aroXOFzFYkU2IR2x6F1aZ98m6VcQy+At02JCYRLP8X
kSmtEKR1mSMCR7OSYibMwvGydMStd9JO/NR3PRbgZ2qa0q5QDTSaoUIc/KK5oMvm
BqtX76hFZyjkmo8pbpvYXKf0HLxuZpTZj5xvyHPeGDvszO9BoFnA01ADrq5Ts9kd
2rzVa3QQYLmkPeExZvWloFscHP+ccx9kGg2xdZ+hTDg8WWMBP6iSE7EdQ4zVlEl4
ec41oq9W18ydree0WCBRt1jlaOoxoKXWgCF1FP1tvjE6Z1FXMn83Pa6hxEmwlIZp
yXzdojAJJQmhycu+im6mNgi/Wty+4MHGT6Z1+xNKgQFU1PHAvVv+CnbBIdl3tiSZ
8hmTOn3aZOt25Ska81TbOOsWj8jwq/+nFwJ0L+Yt//h/91bX6whgvHUmQq+HUdz2
qQgJ0kVkLvtygK1+HBFdWgJGopH6jDg2Ydi7mp4ry6jv5GSMEa/ftMSsKM18JIVF
ysxfgMoQfsnVftZXQxLFTJwTl0jLH26alhNqHwjUm1bSD/IypcB4rPxRpX1yhBiZ
0fkR4qT143vK7SDgJZb+rAWT6mSn+BH41CmOO3ox23d7vxZPtHucHnY0M2Je1YGi
tEZv/r0y2XwJo4qtF1iNerj9j1LwXC+M4SlZXjKOfP1hCzZaL9olk9uHLCRg+irR
WHow9Bn0HhTeWSG4qjKBWSFU57y0cv2/PXjYhyQNscvaekMtsu7p4A9tKSiZzpdK
LEdAgAUCn90GfAeqxxsU18av8cCt7P48f6sn2TR9P9dWmQdFBje+tXf+NmIrl4vh
EyxZmD1VHHMpufyGe6JXfSQSkkX9bvSclBicHpHrwds7EWJwGKu8rdNa5bR7e9r6
u0S9nk9xDM0H1nDYbX2TsY2SHSZYHZEqiQyrBxBouWoCmcdOo/y8d03JMJJo7aLj
81BHof5OWHTlQfymclZhgQQ2rjU+HXNbTNQ+GP8OaCKS20Nr1GStK0MzmHuF/abj
cPSpxcL1lRkmrYskmIgiMvcP1w05Srbz9gbke6GfNOJRQ/TYwu7Q3+yYigbhj+eb
Uafsj8bC+95NV337a75sp8cNaF+4XUuQfrvFFz1TPOxT8kp9CNtb+YRDKSis1xKV
wSAutb5KD+vZkeXQ/K6tXzsU6eszKyOhx8liPa+7Cfg+SbVPKzgYMwsbHVlL5syM
1CxfGXxNJhF/OybQSdeWLnkO/endw7P/op5N7m2wWEbX1xLjqGRWAUVHgFQJbdsV
DK80HNeJnF9EO8iObNaRkxZzsecxGdMU6dnIt9kjkUiY61hEg9dQeakVc7qH/5NB
0shpbPudNp7Xzje9BHqIYcN27URBGu/wlvNPECMSofGZPiykjLO5vlTM32jhzI/h
Xc/K5GNuQKN8ysmd+GyTRLJbGMgn5fY7SC1j9RfLp+/7voCtPMqDL1x6dABLI33j
xbf2fjQqPLHyElost6E3iio41BJ1by1+eaqjQjy0t7jUdxtR9bpdR0qn1KPLRi9i
4A8E/99fni2kZGWUyLZQCyyleeL6zAPFwIaNoBQLGhP47iJ/c0RREt242emOzDne
L8z3Uex0+Hsq2+BLw1pO1BIEHFOkvm5hrHN6vxtOL65LinzwW81QqFBRHzt/kNBr
tBglmkSG9vbcbIgaK+AEoTX2Df3Ajip+lM3ooZQZ+eg8axEH4GSllGioxWHWVc06
JUxh3robW4zxEzxtef+VZz+EE2ErhaYlSfLynYovDeu0AYi3KOmHNBDSUnTZjgci
zlhiMLOuGaIZixZ7dUhFsM18CU/DBt65eLx5CJWednonrecM/QbYJXwpneWqG3UG
S1d4RSwXMf6sGlLxdc5dEc09g4BOo2Tmq6fxaGasAYwUclOcxjk3JTjJxm0LZhkL
Szy/i+inBVW2p4RyNgtYdfheFfsvGwgiurx2hB5154JL+AIAuG3NpGourpAHJCxA
E4nrR776vmQLmWThuU1vY/1XIhEMhDIFy0bsM3/hKh7uf7Et7j1KHcUpy0lkEBWw
nDztDz4KY8+OxfFa4qdFSr1FPbtLte9FMzHv0TqjZsslwGJLb8tEKTOmkGmK362D
NPiJ1b47BgcpnbaF6XSewLX5tW42YherlVuJM659N4Hou4gyv7AXF8AjS6ZLjszH
tsad6KlPacHOByDnGQkbMg==
`protect END_PROTECTED
