`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/4iD70w1z0T7ZXLoKUmU/4cP9/bXQWHZ70Ppd5S1Sal9zIuIjvSdYQq+zi0+Jj4
qxOX5SY+ifI8BAFzDMG1U5rR7FgEyoffwHwFUN4rhHxiOaPZE+cx1COIFnbWtG9y
zgXCHIpljwNMma1oGYuCjx5M4eb3zlBUiyyGsXjKBdVndY6XLlKoWbW/x8rJ8j8i
M/gUg5Z8YuYhtPBHydPRAfVr/BZDcGXdpSyyLWnHkGez8r9xHayrh9vJEUK8EVpI
D0tCYl4EtVRlbpIGhqNgl3NIgt4FvMrOqNIIveWK10PcYX1xBy621e37H7cFQQtO
jW5X5BXu/2Yv3H/e9QuaE5XJfJVdIg3usGTEdVY/fttwToboMYvs/3ILlHsTmP3e
ekOB0iYZ3aJPXhVoV0BPSHJbGwagpUeCBbStQsOlGMVe5VOOG9El4ObYVY0QxlLj
Bv9GrVsKlzI3kEAPVYVBWF3dScjfdqgbpTD1M2tG/0PeIfODD9pjjwwqF86Kud3x
Sc/AhaKSsoW++IeMv1cj1yjV1aSnTeHDhRmxvFkLYPDGyQDH5yigcyIisWNqbQPQ
r7Sz8dBEhfFPshvUHlGG5Rd1ksmAbprmEDUQFKOA7a31rFtTUiK8/hOlLsEAO+wa
sJi+sphpwev6bTDRCffd812TphBNoc6oAhaO6+j/VhP8AKFo3IZf8+xaWdz3O42/
2tZ9yi4aQVAMZpouE5S09KM615A/MAKbMVqV2aARVYEAqF8slHf37QFWA6UKwap4
4E+cXUSIALob0i6OmfPUQve+Khj4kRVz+wTCs5esjSmhEVfxj9iXPAMeiI/C4Zff
Rn0hIe4mtIPAOtHj3owv4NYriRkiEbry3/4rk1wdrVdjy43T0L1iNC+zXk92L0GW
0bDJCFLyo9heoc7TXT5z21qddN8rXtd8kzG06KKGMInijWc1ECeetj91awpVD8ZJ
dzaOkul87APjEsTSibnh/zK305c9Jrb8eFpSk2ACnTg=
`protect END_PROTECTED
