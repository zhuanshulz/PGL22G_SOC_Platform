`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++AmfORlH7EdxEp3714jPQOLGpjwYI64iOU43GAeX9uFZdu7VQVnNmcfZ4IdR332
MoWlrEkafRmxGTGpTkUIAohSU582FIftwayA/DWnDYo1mReXgbhqJZVCvhX8XXek
QPhpdN5faLRE3S3oSaSRE9bvLwKP3POwywb7HUyKZUC4KqX+M4aG6Ee30IMXeGh8
5K2npRZlmRFLzfd2bokO/VoquZI38oSEZCVi7hPJhrocbFoJ8s1a4uSuvAvlA2cO
gh0wntFRLJcVtfDcADg+Pxsoj7viw+QfJnoBpZ+1EHcOZSn07yfurJoTCraAv11R
zoU4ZfwMjnofaSHSWCGpZMUdoe6I3dZw6Zke6/MlTo9QuMHJ4OyO10x+CYhPSPrD
G49BWDyUWt43XF/atpwISAphwEq8ZKWZ0K5fLIAK6XQUo+gEc8UjoloADhpYAff1
5IK4JwVCacJXYpJOCjwUXtc4hrw4ErxWybNq3w5jd8qrkE8MqIMkgrWahFue/cev
UYaw67aW5OdTRIYECsLOAPOE6l6NkxhPy19jf9BFdgIRbkM631iNdbYTHc3Ey1bE
MSxjKEgK374coev8TCHwou2JFJb08TGOz5Zi0X9u1ofH2CA2ZJMjDt8SyDe0UZKL
DHxuwuCEh/S6Qtny4tc79AMqeynGzIqYClP9lpcJPnQdwGJcn70woSf/P3hddB5X
UA6I0V1QDZiPdc7J/2pQlGKSgECVk+EQJS7dWG1/yRnUvh/ZHxpiHVpfT9u8kRXk
yFNzfT/rgFIbq/R9k2SfVr5BWExEMuQlN9O2aAnH0ZwYym7OLBYCo2RFQVJoH+mI
Bdy0P8R0iSVsTN6PwpOzOC7a2JKQuhbCzjMGUqMRLglUtxTYXFF9TZlBYoz+Ln+R
wiSiQWn/dXeDK9+zl6Iakli09aIAHL0t8tHgGCPVugHN7ZIyyR1664a5hccdpbjp
ezo60xKE2BcH1UkH9OOX7eFIWyGgkjhWRKN/cgWrefcPWaZj6nRljCFgjK9GuPFu
0umJjAmKZD4HiHaaTZq1IlIWlfqXRQRIs6U95o72++TYvedqsLvgInMk1MNCYaQh
iRabIY5IwVC3qEoEcR1CkhOBSdDJT277vIDy0DX1gHr4R23MGIbRCYU+OlWUg+jc
ltRlh2pubIYg1LByvQv7Jg==
`protect END_PROTECTED
