`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSAPhTRRxAVsG3jrrvlkAU9RZWLoSR5BMR/Azywbl/CVQzftczVyRE6whPy8D5FU
GLISmPHzbuJWltReBbrtsjtFkM9HNVS8WonihdXqkEq7CwYmBqbw2a72X3e1vNQ3
f+w1gfDXHXzpiXp5WbR4bWrQRLSL00BI9e+gdzPYmVtsfsvl+SS1xSWfU5+k35DM
O3g+XnAw0Av0WVikD1CXDUmbeaQZ2Ls9tIXnJwm2szk9szvZu6FMO70TlSSYqDAM
2cB9Bd120QqvDMVKBWn+isrRBk3l9xpfszYF2XmMoIOd0DeU76mTUpTxW9OX/+jG
+kZWBXG2nKKncdHkHKch4JfX6KBRAgaRVJGX96+wOcmfrv+nvR8Eim6+l7k+NDYd
0OL5uJuOV6Mtnztx+CkW9Oh6kO4lESje0M+GV93kFIcE3UmWgiLN8A5TMc8gpJEH
`protect END_PROTECTED
