`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmzYwGHI2PmXxs0gvvaJmdq/tjpRYUlnycU6XEauFg4plhzATIjsWYQj+T2esfNi
zq6PHKaqDVSDKt75T19emiG91jYWNl4i5vOe2l+k0UoeiEkgsagdb96Lcry6q3lz
oUFDWoEtyjBO1zRf3Gz49WdyNqXiouLvPhnvDqCV4hIvteShJQVFSx2mDPWK1zy5
+flt+HJH1yQFF/IxP50qbji2+tLBuggH35HCtdgJpxmyUNQjXZdWlxC+SgvN8ztR
CljTsgQKr/HRt96wknJydvPn8qdjk67Bw8bO3vUybJ9XeOPwaGJVddJ/tKDApnmw
oVG6k/HYN6W+gHJ3lAqFeFuBRvnjLOOMrEeVwdZ0tO3dSDQwT4nUmAeamYFV4OJg
VcvKXPPCM+KeQ42Alnev8ukVhAVdUV7JpxlCtpQvP4ZmEdzf0gz2nXcybyhbV4p3
aIWa2AGdOXZIQr+DkK8aljG0AQgytPCKleXgQeqsdgjhsU/zHI3fkCEJ+022V1mQ
oUTNYYGWxTJPRwg6NxX5EFy716ss9+7KnEk/CZ6q4STOZfhMiAVgCBdLF5QtgPm0
h7pVVypSzrXyIhRDWWtAuwodYzHgj60GnTLuwN4RF8LcxQwagEe9uGoB4nORHefm
V6QAGYqmycWfpsk+yeQxNrh0uGSF727NGAwU9XLJUgO9dFwwzuYnr0RfBwmLFutp
Memx8GJpRd/acbs8xskU5x7HiR8TqZlTYHu5RmwtTFpBh7BsX8seyGB4NEfwr3gJ
kwtygOlgXYtn27b1FJsOIbueSVsZaWyeBpnre5KTQcy4uLK1L8ZpRBZ9XeS+N5ZB
xFUYg9YgH7WBOCERrwJH2rj/OsQ9epwmhpQ/iFH38XmTlQx//TPmkNE6wfmnoz/I
gBzZOONA2sjvgIucPstUNA==
`protect END_PROTECTED
