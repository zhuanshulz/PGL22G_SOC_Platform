`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7C0SgDKJ/3wFXePS4OsF+Dsydv4YnK0d8uuJA1tgwuWVowwc0xsbPY3gdRQf4q3q
KlFCtkPe9ZnnuidbzYMt24Q7GtVDs2b49Wlva9UmtuUzJlaxlMirJUFibBgpPbt4
EUcGVdJwnkFB1Ry/0dGoBHkBN6W82W8I6Hhpp43aMC4/cL9oX9lV0iby0YtU769Z
Kik+s61bW3DIHelaj7qsZDpVxyVUd/g52v/QQvbHsDp79ABAAoeIrufGIyA3J0rz
0T+bun1k4maZ6k4saN/MrV9SnDlz5nzudBmaxf2fF9jpqvY72wJxcUutP1jyxOVv
Z1KaOA6wWIE4WNjpubitk+oLkQf5zy3Yg/LAOFCH/oZSfZ5sg6/t2rXapK9OQXTn
Aj+CWY5YPPxyVdeibqExiCOonNXSIUUSFc0Xls4VPoYU+xshWcbtiTsBgARaISwW
59jLtpvArJU4uUs/KhKMowECQamQJ+/q198ome1l1MeRuFUQAvJfSAfAwPZSb1gB
pmZ7A8ASP8p1Wd4zMz1ZWp4+7zSEK8gZq8uPUFQfdSLmgTrHyD/wTscEcBhu2Qnn
m0YxWwG2URyEzYF4OAmQKjDaLs7on9KMSw+on1Bhlg+RvQz3eiNp9Wl18ViX/U//
FxwTcfo7Z++5PD8v8AGfEU+ShuK/3YzXhd1gFY/uH+gEN3qG21St/maNXa+Y1Tdl
098Dr6e5bwae+4+gLleR4GeLSmIbrTSI5b17p9k/NucB4SJYF3m8/xoYKxkj+5hG
DbwjVpHBEw0AZYursHvR7ZAvntXPfNNg3iXnLcWDGMc2sIv4UHFNK7vBohCwppwo
SE6+R++INfd8cggJ9a9f7w==
`protect END_PROTECTED
