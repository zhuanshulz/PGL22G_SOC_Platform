`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4mtTgt38uj5wvsWqd5x5B2kuvIdoDhnJfEp0bOxtUEF6iUidB59O6qHJDK2AH8f8
cnCE0EZNfisyN7IMZbMUyLf5aA3G4uiJpEn9Qi5CRBYXDgrvPviWoyXj9+6r1852
pySv8hEQ3HVAoIRJ2byz+vziNrR1vS+epSD7wg+m/QE678Q7AlmV35vJbSrKAGjm
K7A9NkCSrbqfiZGseAqZt5DbDDWKQCOhzODnuSFZ1RiGHpkg7lq+GJdcaCWP+d5u
wwyIw49vPdvglM4gl5DS9iqjk4iVdLewBSj9LXCNNOgdMxAHEGQx8dkUgUvWN3dW
7+jIb2Z4D5Z1rHhnw5eXbLkyd5J2Mrx/qjgetrdzrc+6dGguPqph2PUAZMuPpsmh
wNRkJVoTPHptXnmWFC+L0JnbMfMkxeVw/4m4XqSInoDGF5Z+AmYOale9nIz2NtdA
wVZSeJoFeOaRrNOGbDfcRMZMcuBtNGROO2qoA1JYZCmLqDOJxQMyhZLhIZIXTILN
al2w5bIQa86cNVpz8v5SKAHC/l088cEFWTjDsVxjd04xpSijJrfGKbpwZ79UGHZN
bKsTZKPm9ai4TntncAZG45Xboo/+8DLQVAvKNcf+PViy81USoshq+2GUM9obIvtg
Rs/XYFlT1iUkyJ86o9Sqn99Z1ELmSJi+KaPB/TGxerminbVIgfhYLuRq5KulefLq
BoM98RdoWrVgPnsob6bgstiLHqCrTn/xxqX+CVqwt9cuFUWHUkY+rEA/RxeU8ZiW
JWu0ZCLLlcP7L4eP8qYIcVEyb9jH0uuy9IKbmlDez86BCNc29YBz3ZyDzZpQwmPk
+Sfp5Ug75jOPK+n4baDo4zFE1PakBpMd3YGE/cRgZXlQjiqmE4lROMLVJ7FS9UF/
4EhiiXyL3Hj0IeDfmS0ow7PbAbBlGr3h2rCSPxTLmWUu8MALRnQsN4dTfqhi7mFs
iAh5Qie7t5qLg27YsY8GFYzBgXIviGeLFbCMOgjK28TKK5iKHM/NkcC0t4PREB8i
x+ycJalitRdIjzv1+1RMiqpAvjU5gZJWvq+3Y9ZFQzoPvN3wBy7a+x7VBI1yd746
TWeTE3EdmEoAcPaWRWfYTisH/58LcNyvWNcm+BW8H8RXNwzNOEt8BKVhJ+RiFsxI
P279LwS5vfsvKeYyLSQ9nlZclzRc5124iR6Zb3TFaykCE1KZoaK3McLR3Ft9eUfF
yztEa0GZbDdWye9QgqgN0iq0wEkZW9n1eLzLUj8wqIitkBQhgFgUnjqIOVK69qdb
hOZp7JVfO6nFYWZ9q4tO4+B3Zkn67w/zbKMWju05xIvH3Y+wDdACGMR/rAwyt5Ix
zH8flXqAfyyGt/Lv5wwmSSwicj29KwjTjDBII3zmiLLOkxyA3q9CtqR/JzqPdRYo
5JLq1Xi4vYBpKquX3O1PDsBzEPYSg2GoFlMVHe7gCRHZP16s4zMrN4uP2Jxgwrrg
p+5mKPGEAgUCdp0GUUcMdfcTp/5xTkVuN7sWvCBrnSneGx8m5TsogLJo+prQN7MG
IZCeTTuIA0+LfyjlS1Si1FMddTnzW2NP+rn+9Uqz4gbHGLTsNPQh/KHbRqtuZpAK
/MKzzlgcL82AN4e+xH6ksSSDy4CK9DutBy/JHpnXlpLa23W9HDkvNYyGeUdtmwC0
`protect END_PROTECTED
