`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f56iQKIOpHwbSc+pqV3r1ZXflKC0EIy4Y7HNOtrb+I5BG1JKUBp5XxiOCbW4Vr9v
hA3fs9JN8N4ihiwHx73bfwECob5ujS5hD7mDVr01hSf1uyxy4vX5QfvD/Dsg4nzO
dbNGr36xrDhy6FeLcbeG+nc0x9mG7WD5mgjEo4PEeeaFdEL1SjlSP97B8tDahVye
QWU+kuPkNWOK/Arx4hFGZFqpK+63XH3Shc+khaNEeugdqbH3ClBjOzCjCPJ5NwiU
zxCPgPv4fSZwLCAupvQVhmXwC6hEI3SxrQ/kypzVPNfoHqegBI1X5UHr8nvwnWZ2
h2VC9B42vRji3DGaerDDeJv3ngg26gSPpyM1iGlUCmszpJY03K2q6cdcNVlXemcY
JxQDbtlg+fITeHuJrrucD4RTD8uo9XCIsx6eemII+cbZ+AdwivXNPOSGYmWTPIMW
kBj7+UrauV7rxMNbauTfQrHA7ID1jZJ8Km80Ovi2TB/gKfSIfuLp4yW8OZ8MEcVj
fCgB+evSUnWSKJIanLieZj5hEYvTNtfzfnpOyzbwyBf7gR/jlgAPBIJu98dgXeZA
mfaFkJ48iwDpL0bceg/6M/iNdg34OOLyp0oyItFpn04n7TfonJ6IgCtHpvhe7MGG
kFTGX4mc4GUcFm92UoLpVq6hKjO+2DavcHAvKQBQH9Etwa9MLzty6LVmX730mqyN
rIYoAtfb+mnVlHQ0JCk/kTMSx/Uiwim8n+v3Dz77o4B2QQBcyWmDXxYGuegZ9WOm
uMpZTz1k4pTHpfN4F+VoEA0cm5+CLPWmJfVoUa5juKwMqIUGvMfJijxad3Nut24J
H7yzz+RRKr4bogyh2u25dK1pXM8jBLqbP3RT2riUp9jBuY3Ek3Pk5nrCKEM/PRzm
vRrSiTYX97XtiOKRn5Qh37gCINGIRWcvl5e7ZPZ82+GUJV/GaOYQOnWLSJ+bI9vh
8mOfaOWX6E8VC+IKRthwr5HgvqKNhI8K7nmNEVIuubBPbsEyNmgmCwWfaNCtDiR8
yB+mzMpyXQlS+fDjK+m+1c/m62O7C7Wo82RKUQhK9nBOUQtgBxrlPpr/g07wFq/i
/E2QJXOzqQoJ2EtwENWYdaOhf+wUzwcQaaVWPBGTxRNFHqnCN1E+F2Zk289lpDou
7hWbkGTxysrG8Fk2eexPUi8DK/5tY3G20BgWmEQmGJxepXaJAwi1fSH3Rvum56an
QKYOvIcTYWkpYQ5sSjhobmbBKo/xoZ6fmKnPHwXWtfhKn+sKJdfdn3lLrzBsSdo4
xr1Mjx3U7clV5N7eo+OjoWFTTwAx/Om6sDqikbDzowDd3+l9WGsHivK14Rmi3Jai
FjW3maqaoxzNAqcou54cO/cID9ixAc6J3+UEMSIzBGySg0+el4XEOKok5TEu5Q8s
BH7OTqv4B6RrleS1HxtEU0Fel8R32z3Ct3vzwUFRK35QXLyV7MVPkOK2bcAFzrlp
C31jmSUWKb0Eq6GrUFIPVqdjhdzSfUYD1EYDugTbWYg=
`protect END_PROTECTED
