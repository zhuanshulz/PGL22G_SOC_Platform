`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
55s4ReHYoaWbQTYzLuu+69wiBoriXW+9N7g+CqHr+ZtuNuKycmaV1aP1x6720Ifr
2liy6T4t3O4gcmzEyEgM7qUs9CwoslddCE0aZshubPLj9gsDzfd+LNMd+WXaZ5QD
3lBTpPzD0IuNRFBTEqhZj2c28uTu0n1dzkJ6Y1pgZBgqEgI89phDNjNwvysnYuw/
EE5NpX66kwNj6/N4eaRrw8pwWj8Om8igpcW+pRRbU9uF3A88UvG0Rk8ZJ5GWMkd2
Y005pzT+xrrLwgvdfw5vemkdgYcRsfslKpEum8SCmoh1cIK8aPNLiBDDykyIJdlV
TzLS7DalOK4EKvBYSillVPIXwK+JFtcuF23VUTOPE1sT/jlQOe54eMLrYeqBODdo
0DOzTKYBnh2qiA7/7Gd2yVSMbqdCCVG6MmAs5xZ6aTMWZQQQ6rrGIUipiz6c7wz+
JQVajXqH1N1BkPBYvNHIdO9fvvgFSD48j6+/jf9QFq99BYVEQ+/hQUzlJrauxB4g
RXzg9ohWCmgFMknFMqx9WySfA3/1fqrBAUNFjtZjes/He+GD0rmEscc++IDxFpgl
zepx4JoHmgM9cd3o9pm0ZJldaOfcdbO5qZOfcMcU7g9TF4xROEG8oObiAuqoWhWO
hmqg7pb1/9wDmh01uxPT2YrAzvKdsXV05GUrVqZG67P/9RUtjTWWiGeyRyuVVQ7r
92uQ5Ll1KUQmyJzHXHIiOP5J92rgwM613w1Q+iso5D6tpG+bfwq/yJgSe8IwfHgX
Fm5irsso/zZ/1Tx1zYCap2CQ3MQTE8hmkcGKT0ZWZNHA2DcYo367x+MS9HMY04k+
BYfY8NJ/3VQPb49jBcZqrLerrdj3uOOVhRMlsPvcrbZhacP+3gvM7xYfKvB+HIo1
Wo6ldc2EorD5JWegmLj/tDD5SLFMuHLHmhF7iRNaq0DK9FLK6INhYI0M92Axheai
3ODtFLoSwaIdSvJ9k/EGZPLvHkL9ORhLp8GiouZR50uH5aES4G5s1jfcByA39nEQ
OGOif1w+YOd76dha0RYVBR3C8J9a1HQQJg6TZ3OHGGQ4YPmT6/I+BImDQdsqDxxN
iFOgzAo2VhBpxWAzJ3oZt96mnGR35ys1z5DFNPH05pK8zw0EmOXC5czyVjbq/NU3
tQO6C3RH8a/cnfqbUJVf1D3FPhOFtoj1UKm0AQyqbilssZTEUmOsrAqLBPiH329i
/coCxZOvAguu62sDQOqXEmPa1HVJfLMVEhlzVuDk5chQKT9QnqV7etGO2Ze17t2W
I6HhHyjOT+DynC/eucP0jRtvcEp6YHfcrpdHdF/TxWLWTwS0+DCf7elXK/119ph5
K36giFVGn0DWo3ofcowwI6OwyGcSMlBfmFufWrPM5nc/vNdJ8in3eAScITux8rDJ
AfO4XdrfYNJNDOI9BewvGaEn8O1OJtYuqc1sERfwD6azLvYRD+d/Vu9mCiYlCLza
+F2dJjlPNkHBemVv39ZOGPL9wr+ZCAaQj18Rfb6gmhbC8xjyUzUH+1fRtt6VdKC6
fpeveY1Cu3s90oTQYCPRs5544aFG3jEPG5CVJUSmL4V5FnNE17zJwwgfsOrY/E4V
Q1VSGwIXBS29S0vbngM0Mg40ch97l8OM6/iB9LrIh7dVExff3eyPFD8WGkaTjUT+
4aDgEN29ecDO4xO6jTDLJIJE3WIONVTKbeIAYc9ozoMf9qZnGuC4/7MkC8fSGrqM
0aS1h60ud/Y1TqwnHk4avcnrxLNtsjhfAs+8wNo/krDlNUPeSYcC/ewUEQt95RkK
fkKFIwVtV/eYu1lMOu4Qk5BN9xa5+9itqY4qnKJlGdDx9R3gRABRa7yHyg/pSU6s
70GRsjpmDHeFj/UCOiGbNxErEQzMRKCkqJD5VsBo3lx+0Gb9INbVGrs4uARceOxX
/0DM2gWvCyNjJf1xeV19jNUZBVRMIwH4XokCGwm/5NAPwO1kqPDR1jFbXhkY4c/n
zyMib5/kwR/xtv788OXwMUlp1alq+pkYrc24HSVKBh/2XcybCxGA6EhGSXcGg4Ub
7HhGaqc+dXg6pfLDR2fXXACJjlxQ0DM84OijdbSN7KpNM/7Tr6DfKiOF2WQkVCoH
ZnFKTHesYfUfMyKNzG1GCmajf4T+DNe9/ABh9BKrP61+zE+6EvjT51P/YR+O5iV2
JSd6uenjJFrf2BKtsaIymEI8S/EB1nVNAstO+MOBT1oomQoXyIvaM1w/sf62AqsA
15QLwyzpYwYSf58Qq0ofU4lQLYj3EK2lI0lIu09slqhUn+CD+Tw5Xyc5TO0ngTn8
X5X5pH3Qg0NI/hqYKRI8Oh2GWsMOxiUFubDhk4qB85Gx54O/6KfuigVf4Fy0zBW7
pZNPueknL2GQpTDzFMxOLEpvLBPeRnyLOerIEOULRRJdUVRPw6ZhV7BKkXrHyHpV
bqi11vg9Cwg/X56pFk4Zs/AjeBWgicNV2repvEiSG2eq5oaLCwjZFX7PDXbFN4/z
LAbdB4pKSiMNI0zFyKsqg07VZvynuk8SeznfbOTkbiFs0f62txm5HRzx71JttNrI
nQYsxPYHcebZWRH99wmNQkjYe/GGSLHcc4VLPOzCYD7gGwV1jIju+8Zs0c30e/Fk
MThnLP0HkZuYtJLEFz3GPshY5NFHgF7/3U63KGMNBxp2Z6/9ElkzWIqI16E0jjQm
o2x8U63nc0dp6heVk08AlRnGX3DgRuChcKW9t25612bp2teqIOAPrzYK4ks9+wn/
ttteWRQx3OaCfTZNPPXJK1PcEw0lTbkEc6d/DvWI4LX1bV1+30ej4HWCqhZ3yNPT
5bBrNtHbb4HQy0dO2t9nagXlYlDjMfi6DrVAjWokqsyhbibs8pDfv4GY3hr5RDQN
23o3aU71P2gi3t6ijKUtx9L6Kd6fcdlEEsnhzhlCPpA0u1qJVYPFpi7a64WWhcMF
5NhuYrb0Q8mK3UULt7GK2RGncXOZTFbSJqy385ktz1wJS5cLJy8M4uyZLOr/sSAi
Fi8UQcJAv1CAzZQIcrZFdzwJSli+kujGfLpPjsBHffqE9fylmMUMNwXkSRjGbN3i
QNKCbYapoxC7H2uPSKSa+uGyOH0A8HZa5//cxuwsC8enkVmbFqAj/dPwGd/sNEt9
w59wYZqmdQVUkP9YK+A+esGx0Vm2Xex/hMyKabLNDE7J69GzYGiczHt1zkt24X4d
+bT7g2ZybQ5x8lS06g/jhEqK/LFEKVIjYfX3P+01Pfx6OK2wfRa+G8yS4vk7BwSR
6sRUtkKJzSXoIgqxMDis2USRx4tDegLGlJhWhCLa3fiI+sw6GxSxxSB2CQH/hbAl
UpGOJLs2l0XpzX6neZWpv3Lehi8ignYL+/AiYLs7+5lF15s+SvsBg6GWWO5Ml0yJ
MltLdlUrokV8qrPBq3cCu6Dg+BdcCk1l6sceaAwLV7+KxxIFASmdidc/RWIwtHd/
SJdpnnO5leYor1eVKg0HsN1SG/V8eE2rMvbbvK6hjc88LbIiaR8bau89syDWWJg/
RNE/IW80J0nDrkaojgSnOsx27cUjgTjshJ+kuKYiJgp8s5WAbLGgu1aZRloJLlXy
fTiyfcS5a5mjMoZIJOHePqryC6rAcPlWU/rjVrh51jOdBtxPEvZPqdciT7/gi9If
sxRjFuRcfANwiS7IEG7ZtD7/ASaCncgNSkiJ9CpW88zqhp/5YBqcCXAG2sjuAHIa
LhUzkWCVfbYpX63HH57Uu59BTbN+7qQTYymMxPx4+yqMv+Sjc5r31W6sFQPcYQPD
P1MQECaX+hdRpWWPL1rfgSRXcFLgLW6p2L1AmwCEYVC3MeUHjz/sW7aAKZYeIPd8
hDme6xgqxfwl0Q4l7IYYDUWbZpIlccle22IEKXNBXoFV5FUozvSgUXFN69D7YWkr
69vG0CmBKRDCy7CJ4VlAPoN/gYpxTA0gIwJtPIC4p8Ua4YZycrvAPE4VsPVRt+7f
hxHWeeqQTSHR7/+NEfhFcNudIJiJRb54E+knvkhvgGqCWCj8rv0ydUwxW0Yb0hFX
yPrdh4hxBF2j0zCtvz841ZIs9CgiKPBroeJZrsF3kvUXXz+44ZSMg4xkP/EsUHiB
j0qPam4PIwAXXF48DJPx58clponkMhS17ajg10X8sOCEF1RmQHU5CrNWfmg7/Fl5
gHaFZokG80YV2Hsdx55Nb24W1uK33qxcU+PVp3rN2+AUwHPbup+i6Y7qQjqmYd6U
ehOiFBdSr/j9n18HaW7eaDfLaJ4Q2uizVUR64AZlfvYCSvT9kXbJRDYb877uF5Md
KfCl6yWV6jqiQmoK32mg1e5yjHmIoNsF4KmnMVJZp73HaHP4hxIYtmznG7tHQopv
SMis+QhWDDwI4BDAUVcoSL63BG//QgGHBjzupM/S/ptJKBUa8BR1xFn0j1ygLBRl
Bb81/kliKONI0zgPsXBh1hf6D2Ve62Kqo2ZMdWS6z6LoHl/9Qtwxuo4Np9ji/WAu
MdxFb1UFZGkeucY4yUvK8yVWwFQzSE3+6KRndigIx6lqQpfO1DaUc7RT21BFLnsa
P/jjmTIIGacBZAyloNTMkxzXF9K49bkNtbhYdtbVgfIeGi4RqiQuYtYjEL/sC1Ek
YnnU7qR0dRMPGJPtuo9hJmjds087O+znVnVFyY6ElJVCx/Qvdtt2DWvz5Q4Jkiw4
bYSLJacppd4iS4ht9FOAvoomgg9U2+1gbcFqZm6E9jKhe7qu5+y64dYf2k496fNi
Sfpz7OZWHE629Q6irS4NhyMXuAqnPDecpO7kdfWypEtvlnZZjoYbJdO/FUGiJOaw
MhQsYUz+VEoeY63AKrIY8iIJVKw1otfvo9wOulJNmALeQBdwTLO4z6JRS6hcJmzN
bosg98K97p56W7zpl+WwFEelyvmfucMefZdQVrv1/MlldorVUYk1Ellai0FOf9OE
PKjDoXsLBfcwgHkRDbj1hr0hjrcCLWgKdntRo7pJDih0t0aLmkDRNlsblTTo/05C
iEbkKoFZpeh14sy+xrZ6vuSeCKU89ylrHKjzxjxXeYpCTpJbVkjgHM1MM7JyWI1d
kvnYj/P8s5KdHtATp2G4sY86tzdzbStQHXICyGDP0lREfxnPl4T/zuB1594J6Gty
KwYmQadeVPcTJ2mrfRI/0eAwP8X4pwC5k5SiwlQ8AsgC4QoVYgn9gyx2GfW7lCfb
3orB73xA1xkVhFqZZKwpd13tKA/NRdjfSpE57tTeATm6srWgStYoEIkGNxkrJWjr
lVsOvC3A2ilGNYV6pTehLS/SFEuoqrtIVXjgxF4WNuPk2Jqzba8WGbcN9NZYyQ0P
Oaqmu7072dHvksaklfEU0+fJKu3YvhwqH8sW8aOUL3Qt0QkRO91FGq4n3SwHam7M
8pTB8D8I1Sctw8CzjfeYi2hRA0QdlKxgFitNXHTfQjsNXPm3DJmt7VUjuX1eIjnu
SzNIgGVI43WjeL5wDeU3yLfWHl1UeZO4z3iWYLsqFQ4oIXmqCAL6pXI5EnfVuv2Q
fexUq1RF/HEwVAkH3Y/QxDvy/8khlW9N2bxHNRqes69Gf1L96YawUrb7zoVL9l04
Vkl5nbRlZrvNX+jlv9G2q3aPW5S9M5NrDz5q7OfBLguS62CjYEb4AzgzRQHzwfEp
FqTK2+s94nQ/OWevg7pSsWEKlbq/qmgDUyz2XgrVABj+SAgwC/jbyTCNUpoVFj7k
TGbR9f688qF2VeFw00cA5MQYrAavsOcj4xHZB/q/rgu85LLfq9BnAx+tIA+xnMzQ
RF08nNtVFTTzxz0yPYDjRSlq5lZ/hxDj87N87zKYRbemwbZj6ERQprUphhpuP/fr
93Xs94e8DFhpBK+mI/oXny0gWXWmI5W7PXXR2mamFub7Ieabi6yrNxGfqdpaWl5U
EbydNOnOfbCfzoqtkejA+aIY1Zx/fQkYJrxJA5lY08lZzBxXUk79Rd0ZVqKwjb8j
vXMr8xRFjR0ZQVJwIXGUqQpP1un2bLi+At/F/Y11SH+C+81Zp8PL57H6JreT5+Jo
oSwHHRd5sn0M5ITwIULR01gder2966nnX4hJdkPg3c2XK4hPAVzcoNnocSv5DRBB
hHOVDpTu5JsW9QL24KkM9mSXKP3y/Y6UAd9lzDsaF0BHlU823mDI7s1z9rYLmTnq
tbbNPBXSRxLugZ3Cc0Q6TE8ifRd72c5IjVY+ZFiCaQDleomtXV5VKGrfnLw5O0A+
FBMa8y64mDugyxGvPGbnWrJGwqg1YLq5VEcCtIeLIdTsaPXAeGjXQAmXWnkujHZ2
gimck520wWawcilxGCF/wW8X1trB2u9b41XIQMg4knNFI+h/hWPhLXMKKfIadwVk
hCkBTUXnoxbWlV/MjZwvvONWTCglI+lSyeVTDKmkt4b0EaiX4h8J+KkOF3B4IiTK
eFYeQlBtj8D5ErkPxkZ3AGZ3opI0cwtHSTkl/sSjMsC3mEgElHTDprr8auX5TRvk
5JEWyWEpSZSi+2C2cEmVeYq8GSA9qi9kLudgT3vU9+JeJBBtnitcL8/tbf39JTSq
lOSAdWDbUmVj3uvp6wIa6BYk6D3O9D/1Red+EY2SAxfCIfdFBLYHPmFkFArD28Eo
7kCcLSCXFbnSWEV6/jXXaOV3qtRR1d83gbAyMrIM6hYn32GC6OCSAHu7LtAvwpwK
E6ZJ2ASeU5q7EdImK4EGyREQ8yPetUuC/BSKlxbbk6bKezPwhKe3tdiTXQD24Kgh
1Gv/rWdgJMan12ejOzcQAjt96uR+u1DhBZPPsDFricG2gW+SzMbbGWFmUqQzC1w+
fIN8ZlZ512tZFnwtGSEe9T5PTGckUfAfEuA12mqAsKmw4jwk8UYTgzx4X3VZiKsi
k0BjSPL3ApDm9DlgcrDG5QgWZwoJpnyIVLOjhTUVqKYMLQz/lwj0j9ztzmrrpl0a
zc7bI4i7UownJvvy/RLKom2DPB449b0F7Qpmcjoxarz61qgv1M4sPmleCUDaXgGo
J4+ue7VjeBCtYFVzRsrOypOFely4y3tYQHv8VvZzZUbGOKlEsElaFm3fF01JyKFh
6ri19ufuTrGld1xWQ8pN8ua+JqAPHNdVoCNz6I929rLv/P5+Md1joGXIQPjsjpsl
utdTlQNZAyjIR2Y3SlF10J3zfV3JDNwF5p3wT4Bo1Xy20QhRwmeX02ZTJoTW4mIu
S6eiaAR3x06ONsNq37hCiIFguK/yryTD+2WmEHt8QVK89nXm9vfPP5fLe2lreWDa
Nxy0aDCEz9vORJrErVSJI1XwRYWbZb3juOPXatCM/h4Dp7eKtAgUU6SlcoomDba5
8as7CCgoUzTXyU33/kHJ1r+pg/TovfZY0bj8zZPYI9KV9PTG7ni20EiyyUL5ppiv
u+8H5gejvQNxKFm9V68wQ93cHJofcp1Wv0vh6nxzBc2DidRK7ZTcjqAclqWQVr0T
BVZIbJd9yQnVmo1q/NBSOgfBxpKpSCfB2YxXvBhkNb7NaLZJI2L7RrS0qwMdQdYt
h7JQ3HALDE9VsjFlCimcOFTD379zOI6OIPFic4CDUTz2MS41z2emYGdov64YekWx
2sk4+DNgWuICyZY+IwiqoU1OH/6Fcz/TjZsiqG3u4RBjwN8KnPM/+rWivYD6M1K1
EBuuw8EckRvnqMDVem85NpISUhTMeimFpk2RlvYL6yKlDmjsIGMQKQLGggiGVurn
NCzi9QYhzDUDjIDOuAjligQeDliDm1gab/zjucFLVgLf40JmOhOVq0dI74DNBW5L
G2XtQWPot/m9n8d+GpzjdtcqIz7W6Sf+hQsWwmC1Di6FapKgHRzqrLpJ+EplMOtI
f5+k+JVAkchfPRx8AnGiVyCbjmUq3tI4KJQ0xNAh6DPnZqkD5BBgPDSjjS6T/1oX
uCzmJ3sztIBRTZWj44Lmk3JoKcnOPqOy9sw6XAls6XAesGFlgWCmvwIzEnJ/GZJj
ZB406mEVaaIn3wr9M+bDQmWoIG4hyq35jJnDR2UF3npRO6Cv8fWP2pEtW66ztVEU
QyRBUZI5oTWOFU0AVOehgke7NWu39/XFJzYgoJJHSJxQ839scAuF/HlEpt2fLt9Z
MeHvISwbLKUzDK3nGITx0qmqHwCvI9c6AgyFZ0oMLve7RiCW3s1KGVOeb0WPM1t6
3uKnQeyMIash52s0IV8sa2+GfR6drDn/4O8gwWM7iS9pQauBSj83pUTM7ok286Lh
JR2QfbTYZgUbk8qzfvPx0+P1oAqY9aR/qEEyK53eyM0Zl2hMgyLSU650UrcfrkNV
X3iB4ImVzzW5HiW258X7VMpejxa6h0o3DKGYNLUzeSxFe5owgXwGtd9RdC77RGwu
uhRNRlAV+xHOocRtRJm3rizOtRvapw7NXnGZEfOF/PZa4BQ6j/S2/Qc0hmaPBzgw
mrhmXXBhIR6z7EeWKZIfghIGI1bhR47mPW8g/7A+kxEHhfTkFtpsJNSijW6pBEvp
aZ9w9ge6cYIpV+KUydOrjFyGStMvwlhuKtDU41yoslDIxVIgj40NSpP2xQdeJ+CH
TYd0vc9KKZ9qkHqrf0I3wp+QTsbLKmnR9Di6zR9JVUjG5rDpv30YM2mEyZ17SvuV
5SgQuklimhG4BLZi15jz3Y19FDKiw8mdzf+0pOluP6JD9DuPcR75F5nbZf/i/VVb
G2ImyC/O1LwnpYRx7YLf7xYSuxEGXedsEgyw2EMle/iZ2B/PRkfbdXqxoLfvl9o2
ILB47tU6JjbrvIiZmP0bHLsYA2pXPQAY211viav3UZhiv2AW21KtPSrXYQcmBz7U
GxROZzydTiR6vmWJZFt/HdD9VgyY8xsUZlY8KdTerxu/99qBUVK3ghF7a1WRi3+e
+aB/VrFLXRl3SnwFzruWJBbm8WKDfwBQpp5xIZZR/sJhC2bO5tRsm593I9lV9DWF
UTLIeeKyN4Gn6OcV5gL7Iz3W6Dv9iZ2Ul1aW1uzVxjkJ57FKnpobDmdkV3lDYohq
FT6sPDWaa3wUeGXa7v2XUbpIlS9Pqp+a3TDLD+rCZZ5K8zhGExBEfCciEICejMqv
h575veebMVywTkoIUvFDknXszJRXoLjQF757cE70XNzOU27L4leMbKhsM5z5z3Fq
otoUhCO0hcZ5PGZbyNaH3tw0Fvp2DrU7T2GFxXZghFzjhikrQprx1hMo+K+mo4Yq
6Xk9GZ8pC4dqcw4L3fJlhbLYRs64wi/zyriIdG6dUrRLNPENySLV1tPVNjNIMXDB
p5N+zXnw/3exQRDONatv+OACGKhV3qmvNVQmoXdrsktwotyPCilNdZ8cZz12Ehmo
tGq6PV7tnp+syEBnyBjVWJWYrKLO253h0qbSI7Xb7P7zSRkROqQcHF2BXKoUmUbn
VdNkWUz+T3VLmlj9VXr+SnzpWnHOyONg/GwBJ3YCLHzgq6iWgZtCLOXc8qS778m6
qcjnuMhmQ61dkx7j9CO57lm6qwTTIgc0LcAab6PaS6MBv9AyvLLDAMjXIsSubjxl
nCbyrib5tw/X5cGVfrS0krP6DGBjBLjalyXm71anQ2Sq01XlA8DSPCv61tC0ghv0
jOBY7RGmEvFtp3lMLN8nJIbPIBROP1mMGKjHio/ejD6tSp7BvLPxSCPBfbvWY8u+
OotZcX693rfTt1g4bIV0WL3d/YyCWd4HT6ARHkkMvzvQQdLPkb2xEsx4DEQElPLV
loj8i5BHpw617k/0aDE6NQEh6Jx7HXevDwPaxl2WkOkPnGc9jISxumB8N+geWDVk
2jOPxlNdFp4l/7iv+MF1YusfFHEgz6+l8WrLSIwvf8kgDHimJKIes4/RFOwSr1aw
IqpGj06mPQBAf8IOTSKyYy6TiA6h/hOWnlEMFQQ8A/YBeH31MUoi3RfQ2lLYQrmp
eEy1kuCoz443mcGwReGtnjLjcsIeHukxYrYqSNLssOrm4PdXRrWqdoLATn8awU8j
Np3RoqpiFdT5QHAQjoCgqECH1EJmp8R94uMHRk6Znit1bZSUuBTuNHwyVegxaF4j
HlJ4pa9IeZpYqFIyp5YdUax9cvFHlcI4GPLaQY8fF+k+FpquMt2Dc89NtBQSugOb
7puMEEuEIZ8Ymmv2wJzeXavpDx+tfaGgrHmiWZkbOhKmeQ/m/m1QzvGvB4P2Qgd1
euP002cRb8gdkCtF4AxZLMnP81cNnVF689HMPMnyY3oJJ381knjCJA1IMHFQLGke
Xnrg108uTXg8qYYTKH+qWKoiGvV3uQv4VTuGp//stXPVGg6CWM+Eg0oBlEKe1OB4
8SeBkWksK/V8XQNG6JaUKOGlVgwPgGstfns5YxzAcaWMUrX8Kz8xu5y1FhcbVlBm
vJxL1WEswpwjIaVhXlHet74/AlH+Y1lJvRaksm+bxzEwWPDQODvNPtw9r9Mj13WR
obp0CdoRoWm/rHfG6Va0kV0TJfTbQ+zn6t4RRB5nueJdUcXP17janWn/DEuzGhgE
GReYV5vJ5HASecUTk6GBjw5MAgCPW2aJ/oJpWVXrOo3IJzCLMsedW24YFhw2NnYp
vA5fn8VhD5873E7pVW4J7oOfCkKfxnI9mkNCs32AGcXLuKVCRV/+uSu9YSg9mk89
/Wr02+AVN4PEDfSn0c8wFFv9QvdOcXWHlrnIXBBnWuRhietfWiqdN2uGuJ4vVXmq
h8/ACe+U0S8Tq/Q1yLoahoFm1dRgYaQ3a7IpZ64jKoZW84Ur8enuCtYCFJWagYIG
hxlMDnlgStu7F6qnucqbmdeNPZ8dMajSCuklTmCtI3HG7TN6X4z5E+9HOAjwANDC
RfKBFcxSvRSSSZa86Hv6kZt64PGkwC1DmAv+57WzfBZUEubKCxY53PrFYPz3l1QX
nRukDvhT1gboaOj+yvIP8IlbLna1S8jx1CKLb7FDqD9QhWKrEktrPyjTCGPd4ZmX
vyMxSC1mwLyNKs8ZUmhzj+jBdZHDpqgFHigDjAd7aVHIO0PWDa1Rnky+T+gzchKd
REkZHF+qR8OBZWiAQZSVoHOXjpNi3BYFT3QJvmvIoCrxqssbbJAAY9UzAiLNApDG
gTo4zt/L+51Od/Nqwp/cHirUYy2LFKUULH5htkAmJguT+4Hpp7dCTYPx8D0AYACL
1xALwVo2O65lWso6JE4plVP9qR6gNsv1iWx/eJO05c58xw1ixZf/sHocKvHXVzsy
sgLtV0/lwTLHLcOcbI1NdvsGZet3TCqZ1daiAAWqYbGwEd5rW0ehTYRkwiIOoG9H
tIUzBFyfB1Joh/2WipSFoEEGrjfRxljk2rTuQFpBDmYSR5ybcV7GeIHiEQHjQMtX
J0kEMMA5jsdYRKuKlJ77DcC29F9vzNUmnJ+lZq1eXu/SJlMYBmpJbaWqXWqEBEBP
W7JQ7m1Vx/F8/mviYBX/OILjAG3O2tpAiX1Eg/ukwm7pWjHTPIXjMhn85qaHKUt/
JiYu8zRchJyk7RWpzq8hqvkEat+d/yBt0LPvELTPzWE0f6NviAPlIWh/T5JfleCk
Ytj3wLwOt9e3OhieGwcj1zvo1FJkfOtosgFu3ffmiD31uhkhzJ+sq0tXKZyODl8R
OeLwLhzusI9Kmy5db8tJdtaRfHInArrl0w6xaMYFtfJ4yyxONzYUN4XCv+zjPAQB
9ATUsWqZGJKZjYyQISUtXS92ju34xRCe9+Z8Mw3r5otRPay2Hu+E7YnVFUvWHhiu
B1AbKxRr90iIbad+/6sj8cjH5ZJLX4pspkISNVq1Rcuxw2IvyctLPjXIV8e4Z/Kc
VkdlFvSgaghrGh3LlyOQ2yLZdJrdUXVZls95v2J4mOYOgYwvzR2/MVa4dd0KM1CN
PQIGyNg5HRu2WMYXtrm8w3xXy/YYL7BDVZHsSeaxZXvqkrr/tazUcgenj29ikRmB
xHyoiM6lqWc15j4uhIrscRQJfNYUPnGqTz9ob/0JjfhzQwJiW5+rTLJfVXkYkheg
F94LLynvv0o7mAjBImqneLA6H8f2NRKwKrIAO6wMAz9k8cscG39Au+8nWPXA2hQh
xk0QQY5i/NOg8/uBxM7rmpeZ5M6rgAIIPF28Zhr0+/krr3S+jFUszzfLV7x20XLG
ncvsrN71hDxOQbdEVBa7oX1hm1y+iLoA2HhJ6qqbk0Vqt3AGCFua8ahaWlwPUdti
X+OKqLCpe50WZo0p0GQljJk1Qoqm87BoZfOocsPEAuz2Tt/RIpyTassDpK1b3ceo
0fra0ai+L1mUP+DeDyD9dBRfggxEzEmS5tkT9hriN8+fNHopoT1qVM2nV+I/NyqG
uHfkBZjcIq65Qinx8jAUwZUfV5K1rSCaa4Jt6nQ/kbXbPU7JKq2YlOe7zpMisgLs
23ttJD1sJ0JKohEpOX206Otk2e9yQXDLn/Y2wKpxZKsNdGjxYLccZXh4Mr+UFKTt
h9lGFg8fffbeGH7fR565dY/mHlyj0unxoSwzicbSx98OaR+URIx4YIL9q2mqrPMR
ucii9oN5r3dhcQLvhP6s+ioL9J2YkUuKXlZV+s5X24EzB4iv8FqBGfSTqz83yIhx
b7GYJIUmgQpnz9VHW7rwDo2355+OsC65MGmtcGioUgEMGE2eGgjdh0q72KLdmSSc
taZF97WfJjnd7HQCv53GjCtcyu6cbOTE62tUtjQYiskSBAO8oLNxzt5MNpxxF+hr
2XB1SC/iagbFA/Quj3QR2yu3ndsAzSdBW6NgJX9f7EFKO9yXpLGBe22+fmA6VFLE
tD4XvLecyLT4IeipT0Y0IrSGry6pcqMA7H0aqWRTinpKiABOdzW7NGMqhGnO+aXN
6fJY81/5PsQIAS6L3UOnLEN8DTdwBId5lCviEvR6M51ByTa+Z1w+XmzhmODB56Jm
IYvbbmIQuPJJ+dBjwzx7Iuh5nnJeeQDaX6BDjW0L7wz1pK1xqpysNkfkwSUkYxhf
xevuGn1DunIhz6GaKp3qrjch+ozejCJL3TiO0dogNyPFFGJwIHcXmD6IuZXQDSqa
COqlOicCIoHtTulNl6SO4eyc0hVuut35RPpmmcC2v7hCmotsqeFsTVlkopweS0GY
bjVuK5PQCLXYwVpxQo7gevK7mT5sX9mBXn/lHrUDWjxZdJjMVIAJdw5XjSpoNkrs
Uf6sfHNyAjD2vM0NnANmn0Qyc+LtnNmSSdFJ6QA7IYwUwbcMk+E7eQEEIYNTfF6g
xSuvJYwUl4gxySmwd3PPPhZPnhSkJkhK+sAdMCDSSZYOWcwnYCknNjKbtlIijpkX
LIWKxHVaSLqr+nuhT15b5sWF2EJRdsY5CMfysEwsreRaVBl7t1W7kWgwEHLoEuM9
uzDoVGxxTMmRgiNBnNC5g9dQeuFyIgMDAHjEewS5GrMHKVBW/lqwEOH6O4+HiFdH
tR6WkgZFDM1Kr3x610iF2qiBmJwd/A+Ntf9Q/ob7KgMznZ9IEHgOFhrgVHlR6eKq
HZjMJacAAfhMsA0YrdY2JJHmp0+DGvEX7ssuz5uZmeQsCjrjEPXU7iZCMQdk4IiI
mGjha2Rx/tf7VidUfBmdoUX5CKSu4Azg7zhnVxvDEdZQOHLyhWyihbuQ245zOz12
MOSpOR4xkBohWpDNSw5C7iODnzrjEqwlRoeAlBLH6H2b4yNdhfrqKHnRwRV9k4VR
hN8TOCn0MhDiEBVdPUhpULhbU1Vul38bSplUj58ycsCwVDbvqt2dOr47iAOIq4MY
rRVMtyzj9ynGmw4WYmJNXofcDaI/Gb8lU7HJ6/pR/MWydgLDd1/oR4PtXjYbCeJU
3ftRynru5+KR8NpyDJH+Ims6Ne14N0KdrKgKJKqQDuGavKjVrmuygYKTHR6doprc
mQtTQ6c8RQOIajAlchOfBaLHDapPX+BKOZZhiAGfO69vc1oe6dhXbj+0ZzPSYa3+
LAfGfqPNG2iBM49ERi2oSSTF6XxoMPoje8v4HeOwcGIyyaZzOJvAY214tIoZIBKt
ZkCcjJITRpW4ZL3I9vszCM0xNH9Xb7MGtjgsn4/sxmMDLFwNCf580VtFGVFFxqfE
XFZFiBndVmCwaONsfFE8WqklDklk54BN3MX5Mq3JmN1Opec7buMxVmjsAyKvi/DA
q9xYxm+7KEx1Xbj9n9spP/kRXv4G4k067hQOQ/xhvJDS9B09G1D5cozTnql82ofs
kwN4VaIjNl/g7v+FbInYrFghU3iI7mQ7cH+/TZJU02GBlZpU22107cdq4iNuJjfx
570kOEVo1e5z0VIqaMsnupQ6zz5eXhK5E7IPsetOvBQF/K1FOCYHjaIhXoBY6Rgi
Rgh8E6c65GwFyFYuRMarQft+uIBxlNFw6tjFZQSH0ql4P+xY3cSd+n/bGMZd11Mk
ajxRC5vU1zUnFPNsTTisDa8HhU4eL44NuKedD/zKE8ls8seer/JKcgr4awwUjRkq
Bupyl9uiict1VD3H6KplprbFuOEbYFtn5rzC+ywOFUzKrvrwtstg4P0A0WBcNY3G
y89dcXuOGp22TETiUluhlaE37ioS6R5oHMeufjRJwL8Lk1V9hYDQB7DqQ4NgVdS9
xJ4qygxwVTaAdtYv5EIQhv5SrRLPm058Dof1XLTJKy7Q1/vtTAPgC8G4L4wl1jB5
OVibdqdZr0QxQTSA7OF7tDGX3hfXnu97kpvv5F9s32nLRu9S1Dyo5BFuZ53CjBzo
zEZMQVyYBeYZFtPVbQgluDWLTIicOfG1MVNC93l+ZSxdKo1eicElQ1bMZ377vJKW
nFkO6fudSpLj+IeTPHcLQ6uQSLTmzEG4BfhTaIc93spw24rkfxBcE10SyiJmlwIM
UtMCW34c1iblbkmwFGGWAVOVZqw4YutWjxo4A4q5Ur+5SZd5h9wi2zgV3/PC/uZH
MllsDTInsXBxPj/zPenlIRqWbkKO8FEDx8UA2f+EHKpVskLa17tJ+cHEn3qxU/A/
Yojzi1C+IZPmRsvzym6wMMOTInif5t8Ohoa5iV+WtyU1OzjPmHfDMXL6EvUu08T5
t2kiVjUUF/UKvNqjv9wk44p2zr/GaESl4FcXZ4pqWYAP7oWO77j8IczSgVThZ0wS
y2xomBtzq3xARfLV52RWAIy6w3bjyxeGFRSgE2ffy6c21jypJF85fMcxfjbYTKV8
+hheIayJHTQLzTk/9MJCnJ6/gy8Rp1YSJ0cvJKVu0z5tkjtwnoCNoyWoNEUxUvRY
z3ih1zvJdH4AhIl8TzD1ZHsyQfHfGGeXyvvnkzIdzuwDshc9PH4tjQiYAwUZBDyj
nx+DamaJxDxU0q8r2Ig7/X0jRj8qv24Q83SkLygkjy9rvzOMl+Cx7SIM331fKeSF
IkXkMh0LzCJ+PD1Ih74LFyMsH6jQ0zHD3Uq2PwSIGtnK4CJHW0efRDkVZdNHTn1t
ejmr9XS2PlOZBIWCpGeA13vzBoY601pQgiW7NuLe+rWzDrsMmNssu0WBS82IZMm/
FqyNuRGtzdCo6O6Zn9ocfObLBXP/pNipT9aLBpGiU+d4laeL6ginMh4PKtK5N9gM
4ZVTNtuP6eUmsjFGZqNrBy2FEg0JevLMA5+4lYoFFOgg4VGcw+75ZDx4IftBtANm
EugJd5cx9KUGbI9UhpQs9q9KOjvmJq5HGoZmjKavArcOLoRctDPRBOZx8JhD7fUp
QdkGC4oMi4dqoe9V+RZI3BaHqq/Wcq9Zezq14gJRW9I46rVjHshsSN16JDprOrlg
H8QCq4qQ/ks6ObVouCx19hCY+5r5Hwc9u7HYAnnniUptc1SuAdftcyawNRjNfnpV
tyNosvACOFzaW3+mSiAczyOS4hErrXtkBXDNVrYl/b8LSumt62MixMbvLsEybeQQ
vBhI1OGaOm3ogDXb8B2pIodgkk+s1iDEb4jT8m84xvxB4SIXa3CHFn2cLy/VIK3G
k8A7FjyZRWk2ZzQCvUh+JEN7EGoaw2weIsDKTbT3ZgJQBjsiGjKHJiKQDVxTspx+
i7pqlucpQouzfOJOZSM9J07ZTtbdkR8SfBtEfbQScUB2+P1cPkc6Ys5HfS81rX9f
A20swVzIVPvknlQB/9RiW11lKB7g4szmFvZktt3auwGnbsM+/sorGw7FDzmVgBNr
vrul/rw07o3s1rpFbnTD94PjKUGUk7wpCxKJH0vr4fokuUBbMDp82WnoOPZipu2i
Zs5xh2TQ+p/Dd6y4yxZ/JfcG9p5yX0H4QgavECN5GUqKxuvQ5Lr2lQNrPJWWesmR
TEaMhl5cdKOWsPUkjEPDIgKvbCGjwZ3Rh4H4qOG5XuJw442druaqa/pMMy9idNUc
n7m3RuUD0d03ZRfe6O4/b10YidFcmWPzJkpGDOCiDb9YzyH8/1Wc1q56qVLRFQAl
tbZlI6Z4OxFoleMRmVCBvPKze3T6CBgnKNjC6A0uKxWXSfcm+NGwiDtCvHfDaS/z
LPP/TNmFrQ7Eem6sF/9pH67gv5RcmxMbuYDuHQR20UBGO4okgEyGoZvnbUL1uQWB
5Iu0uHvVsuxOJTwZw36GChPBZ9zXmmH9YqP87C241HPAsjs7KLgkCEbBKi7rjnRQ
AwGCLBx8WCSVqOoXoL7AIfxRIshW74hrzf16YkP10MKKKfoH0/HQ0WtK67JoTNeQ
bMB+iav0bS+xH9feDOX8P+qHWiqVOtoO4MnrRQVIT3BQncz/euWnFERR26iIepj0
KzdELjqH9UDVSmp9Jlowf6ta4KX62I6eDiEeJ33DeCMeb9jKt0BR+ZkinkOV6CA6
xN2lsfrMYBNWHt4WE77dGEpSIA4hxULwJnEfPYlFnYEJMlWsmFsR16A44G9K7tp6
VXkhUd/neyiMAJJJDWcIDMljyuEBSkMnZ7ptrTlrxiHd+35u4vmc+OGPoQUJgRiy
hP51b/8Tm95Jw+lKNrEdIqpwry4VJ9Sre/MkBnawRqwaDeMFhdLAQxzOl6P8vY+8
mEQ0Oeo4MZk6gnI2lW6Cnq0a/KfwvWqnWH07IiL+0SKyFoURF7CvQgwHpcoyHQEg
QvynmpB4z5l5onQOYpfvg3WPJpkktnWqX8oZSz4dJkUdt/qySbrEKTsC3FySDUbs
uU6mM+0JKUqlH3+e5aUmgoEIO6KqKbrsv1EvEpefWCHBxH+w8vwcpTfEBlPAJe8W
Eg3m6np8gZclTKT1zLah8BDttZufYOHajQi74TOP+ywlhwFG47VT8QcRi+zmIHo6
2x4QCG3cydRq0mheaDucX0RNX1zREvno5sTSIiiloLM6n59/dhyJA/KfZSscqoDb
lfhlaUf75nBBu1Z/hof86k0T98QmGtOHyQvJgw7+XdfUFkuzKtapBhTHk/bVvBpP
9zj07kHYk0yT2EABCkimS9YzeGWukVtH2+ZNRcByEs/Kn19OEkFQ6BIKbJ5hzFGU
A1k7Ft44+PRJP8mZC7bW5s5NfmHyzmSYOahIliq+Tthv8Z97p89yLpmrGCtjvwp2
x4apW8Axbzi2CGIwInhoJXwMa1oD9HhLVV+9msLVNz8Fujb1D2ZN+GaN9xIc48f3
lnWBS1EYrK2+WyH0mIV2pfLmhFXtTpLPJEcWvXDjRnL1c1EB8WJBpXaFp4eJd8TF
O9w57wMuBDe7yvUOvpSC7zkJmtrYqLt/KGb7ndjZZT5HKVXGjf2w8YBLm/HTFoKc
uTHJFavtBJol2RCW0PotC8veko83SK6U9yMZRbkk10L0TbIgDGfOgK7KhA8wEipv
iJPGjobQ8VwfwP299tBRJg9ta+1Lw+Q3Z+FThXJ33vC9+TzpTlLfylnidr8it72R
FFOPh1bmW0jUSpi/M4po6D7eUnHeeT+AO28dfH5lEVKKCTW/lgZeKz76Riqb2Fwj
IlYs2w0erwsSa7WeA/idYHQ9fjnNGgQZJYlNJAEmbFMqG9UjWc57AxwUNUJYJ4w6
x2owzaI0sp/fu+7OElXOtSFl05NfP4+S8FlyUiKyAl21I3kSBnbqQ49wvyuPwYtD
H0IQ23g8I3V/6TAQb3+z9h2YxwlKojtJ/VxMHypMBOHn0yvACAU7+8y2sgRZjKZP
jgn8ve4qGZZ6hRLho68Y20dIjxTAKgarfkbwdkNYGTXUT+1cZMQN0FTHi8CScTU0
+uWet276I4V4ROHAi2aXiRoznIJFccMFa9dGh4w0/FJQ2VPWrO5Ii90td8eUm68e
XB7upFSull9XS0TGosHMCuow4+D3VK1064X7IDb00fdc4mEvSzq5gXgUTJSokLOB
1pfPdljTs6hKNYA1q+Kb49b9IunFmYqmRAIQeW6x0Gpj3zQ7oERlomP7kPwOi9Kj
hI4ZbqbeQvnaiS5tw8+eea6q/2+AxvUN4q50MiCmuZ9W8CdOhQvwaLGQOWd4aYDH
fu4zqbo9yyN+pgxPdkwDoTzyYKN0R07PaSbBAuqu/trA2NPL8q8M0pCaWNQl1Q2f
ymoagX8Pn4oZtog7Qy7jmL/mk1DRBmXQOoa/XwgLQJmsjDc/ZaxJq/ZyTmND1ZOr
dEha0bPfYoUkEuiJyaXcy8OysbJm8xl0tOmc9M6hZVi+yDfvTZPdGGkrbvKJHsAU
UgRMlOqCC9K/ENHT8pBVqdD+pDtc952nFWZqNoOyMMoaZJjSNL7qvSQnCIOpQx+O
H34Z+Ks8EbS2RprNEnKalaEyuDYUB5xNeCTVeGHsv4EEybQbbU5ICdDHVUtusHjD
gjNEOi2Qgx1hQyZOXikBtVRCwtuXSIHh0AeUoLWJzI5iRERyxR49pf60RReTimd9
OLp8h+VUz7VG97FrVyuc3WAe0wFeFXs9/3VDfZ7mzbNGrIHVrzICURVcf1FkeHub
Btewk+clEqARDpxnmQx1dr/wK7LHyLlk2xotZyjgVwFMp6FQc+5VuViBLVjdhE53
c6WhgeUnTLYwIhyKkZ5HBlUj5SaYLmppro1tPa+5Ic20oIMvxl208CE0xXT/WCUQ
T3B0RSPG+3veyclu/2uFhzI5lXqaHFcJqCdaSpMstbjoMLV+jXGIlG32mBPrerXa
84umnMi2PROylELP4FW6C+X333OqM5Op7Dyh9oEiNqA2EEeCGKJkvGZtooFrbk0w
ZzOSq/vDyLp6pIqPqanFlD9QUedwZ5DRd01U1AiRa4HzCpsJBefTcBWIcVgV+TWZ
VEfEEBc0yaR/5v6lAzyeajQ+4Vsp7McCTGZgHeEjAyYuh/r8uHZ/fUY6N1+/yRUz
Roffn9q8mUOShQNZT+BHcaAYr+5t0yphWUXPLPOhe6Ks+ygYXSJktWBP6LqYxsYE
YEh5k3vHPo0o8hK8AkA89cJtvLDxvuKUimYIG+TVSBkuh1QN/snmyeDCLYp45bvg
OU5QtqKqkVuhd/BcT6AC8xOLD05SNxyGQdUmODFu1JUO+rcVy57kQND67eHKeVWm
c5N/ZI1GTiooaq2DJjfqWZa2cflUCwUHftkmir5X/7n+HAvelxmEsnkw7cToCa2Q
893d00osqiJrz8UFcxOeG19lyi2r0owrxyOIUyf6jsj8UOace8bOYpVP4i8Dm5xu
dBvavML3mTVk/EPfN+ADu15eqncr0irjVkDGoLG1m5vhzVpFXfx+Jyx0kz9mhkfc
rr5/Jhhpe07oy/w3vo7HHtwfhS3f+kyiyDOTq6TW0MiYE5gqw2JX1t8yCvg3orUB
7pVI2oj66LnFjFONQih0CFlTReUmZcYOQKATO8s5vsT9iXLCCmYeTC+F0FwRaDAs
mDcAb4Zh1WMF8ANto88tMuVMr/6QRAag/rnrF0A9Q2HRXznHQNgORfPUmObWmLly
cP3jxU2rvB8SuhSXdIOGbQUJVn6PtYwXNQAxYUdDxsenIiW6EfUCjimxBVLBV8/X
R/63IYi76RtFlMaV0GSo3sqLRpexzfQdqQLagsq1Hqma9p6oayo9udeZkD9IT8Oh
F1PobySueuLMmZqRs+yi2fsMLX2dE7EJQI/dJbz0J9yqlWsnZROcjrF8mLk9xRF6
I9TInGMqwzeWonexma8kFGUyJ6tUj6JLwI8N9fvQk37ifybYFGclPbEw+Afhf42h
ll4VPBlHgQIcXC49FZrua85g4DdjghPwiJRwGCLlEHoSbOtGsG7yq90iJ7r+jYB1
eY/Muuu7zX49P5j8Ah88FOOsGUcy1uSh9Ll+86JnaiSUf5JxCaoym2afTIXXTWVJ
R0uCL1ZTlespf3b2QHrzaqMXsxODv+ccLmhwC2+awFmTV3Esx7ylPFrd7LdUVtLT
ZyKE9cRZaUgf+4X7SiGsKBEyT42y8NlAkeRs+S6coVEMX7ZIlTrrBFaUkC17iwZ3
ZAAuLTf7wYuzaUrU2RlsDN1iytrtsjmfmv/7vEnpRYQYuMCR+i+71rlIZQ4h6fHs
4/Ybsnu2rX5gdM00D6z6YKwf6zr5i7IGkdwdqr/tbOm10OVxHHH9LnGAkkOeYvNt
a+SqcS5eRWOoJ1w1VHXBOZxKEKyj2+tCFxmXEzr6Ru0XHd/l7SNL5Yd8/GB+5iXZ
PgHwNMQKJr3ZAMlWeD+93SLRyGkCI21KSwPKORWw9bZbvWOngHq4bG37onEkLSM9
FYU1URq+CpXqBC/hUKygzPItbIKa5NWKYsZmSEV0WVAAqEStgZoS4w/mEq6hg2U6
nyNiNTbv+UtdgxfpM/qIpkC58pJcBsC891tbiAdDRu/2apQueA+1u9jS0+qa2uNT
OnwVyYCkaTAZEhXGT5jUxBYv9+q5jQ7Iua3GgCHQLZfAvN3wSvUQ5V6E3NubeWfE
IDZjxUAl/6oSxiZ9LxglrpqHnS1BEF75iSL4C3Hr2+lpo0iACuMdxdKmSv/QPm7S
oflmbtm6bb4354aTEeGhCI+Ce+ffSZkLya+Yc2bdToX/t30tnkJwFHTKuLb2GaDT
wkSn9tiQoVZL03AMouzLkXj0LSuLcytYShJV16Fdueow9qE5eVpcS2bkTlAAxkeO
aGQUj+KIury9Aeg9sIu8VA1ynjgvSLEH/nI8kaksI4KbLaP1IgF+AsEEXXA2YL/z
ws2/VXGRc3dxNkNEOh8H/jtX7D2m+9JliI/iyza9qK5v3H30xhvZHtepNbV8YQ1l
Tf9oRz5DAMOjCtD0FaYpjIm+mASC6rdB15P5S4fbWoRexOJqprI79qHqXIYV1i4I
l6iDROohA/hTDyoBotLGBTG7W1C3TsJRXSLB2RbyYu33NwDQjggQuU7c4Ny4B5jS
kGk7HkHrWsA0dryw0JbxrlUrYmLqZkZVskj61Nnf3nqryueBIOSQe4NSuAmeWPur
/yG+yAhyKmbc4S+Gq5jVvJ3N/WT7qllaS0AOmg7t30/uAgWkjmMIEPbP2JFJuQq2
owxSHQWlcuGjSk82RSkJrSdJbXb4L5+mZAx/tee+z/OX/eg35ZWbTz3RIMy23PAF
YyOlFjAWJ9iGbt06O6b603sZH3frKnaauJRV3RSJjdC+jFnz0pumJzMn4X2o/L8r
kGu8ULvwMVZIM3x24HmJ9oB9HSv4xg4m7/i4/UG82ekaV2O1uptNpYpZh5HCEPiA
FHE2RhD61kYoSi5H8QTt5HhHecx3JXlBP+57T5OfEakIgNwDsQkqvPAxQrdXXG3v
8qvI1HpboZezQ4u9vgcJ+fmOisnr8Veo3t2yn5pH/qvzsQCuk7nkjxwvsuE1arpo
tXquvMv7emKNrk4NhAYUorgRDXfAWcZVoAkPQTrQTHk7MNQuKAcBIO1NnvMX6GHF
1ZVI78VHlMpI+OHhbiP1U6CJWvzeO2DvAenMJkflLaefzhVyP4gcEFrEbPyEZJ31
Kd61SdweL9bhY/+wtxXckF2Y3RaGmSAbTEGsdv6l2aHcjpg+rG88/cGECIro/XqY
auAbof4HUn91tcMwdAR+CbuqXCyBudosCr2piP4+7pIJ9RqFhI1z0Z1baylwYvrP
Puyt6EBYmaqSlwpSYYKKnExWtjxUq7e9mXz2OeqTbHsum9S0LQ0eekl6ROHpJO2n
B7N1F6zTlYqcx6rYOugVK50y311uc4YTz2DojrMhrAhAmhA2gAP97QNuYq30TODD
7GBCMNVaO+x5dvH9GOCcgfXVDV8WED12MC977/IDvt/SamELyc+g+epIJMGAam/s
DSz/FfQePMrr9L9FL5IQNU3ulF9aYURSsnwIBgxRNhHDy33heLrxcYL9u7xJw54J
KxUSU35MzwgynwWIEYJYvURWtm/jZyXQC5okCDZNWx0VfTo2qalk4b1nP+FaNMLu
OnyfzxHOslMtzV6BZtjpJgLeQ8bKerD2klQHDOF5Gz9As4Age42Sd2jgy2ItJxkM
huuOsD1QbDh4M04IYlErsig0aHszHnsy920dHXBlobz7k5YubL2JUyK1FLYOAU5O
hpnLlo8+fNP27Ye7TNwx5QBUW6Bcf/PX/LKYRTomRvi4WHATVRY+WRAR4R1axldF
IISL50iFeDKSHaQpw6KPekS7J0n54J//QjNsv7e1cR46BkDA1xKHE1Wrt8cF3zOd
B/ShYUjJu/x4ProjdOSk/CB+n7TqpAMS6Um0suo5Dt30b9symf0vZC6g3yeGadw6
oaZ1Nz4jmJ9pjy9OHTDFEsL6I/3Du7x91bLtO164twT2pPBLBI1yMoNpCueMxvSz
Tw8JkB47WtzndSlEu43GRA==
`protect END_PROTECTED
