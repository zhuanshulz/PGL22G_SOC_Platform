`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfrsOU6ApxiiDSOVLSoD9jKzouUx7VUL3ONV4FgRqiYWTMPWJcFCOkIYFodwtGEF
fnSgvi/EiWa1lTV7+1oj/wfgxKw8qMAZNKGtxOHL7FkYBQIMaTblXrbgKjOS/Qg1
RZxHtvSfqCHthypj2tySlhcP9fxvOoWpEtafRk4lUZ7JmkKg4bdcoOoC502EIHco
jDfaxQnOi5Q3l/QRz1rwlPJ43FkgVs5lnvolkIXGDu5VnKapjYxsPpXv4u6IKVu9
7H8GdOoK+Zz+Ll2gQ+xh2RTkbISzVoTDP1qAT/519nDJh2K1wD8QfCqZbHK48lFK
yw4jQSaU+n4JtKOQuwzfnV/B9yQqzQ9Xr83ik/BhD8aQvxW9keTO5KLuAIswMTFM
zrCXQTVo2vh0eVrRtQevTMeTT/nbRa6TtKHoJtsduVyo0DUW+8yZLsb2ZS/TTkVh
Tv1pQEJP41mspZBwB73BfY1nxl+tJ4k+6QFezM/F3atGxKoVoB/DN3mM80paqU8l
QsUBinArQUDGEwStq3nFPGP5Sy4Cz38JYo3w1rKwFiJplA1dUH2IJyjeAqTAqvZB
NId2j86spaiK90k1lT8aAhvsw2cpkWG3kKg088PtS+GWEClr5/ikFIQSNn4TkbjJ
c/8Eagzze94M5q85npzqkKb7b+X98Ek0a+B14Fz3QxLB4XkWcSwTzVHnNdWEBl2d
/ZyxsP1C1kTd8QvmUpNIHWa1IkKRE5S9RApWSaz45v7kS88Kshu++iWjM42BtqTo
Xc6HbW+kwcGjZxU1ZOfehKl5lZf20EOacarY2Qwjk6isRNqlyUtnin/7iVQFHkIc
HboF8zqtTiNhfpQZ3iBG6FC5RGxPULWcLKVmcG9YQpOjQwlm8bU+g5XlwUNmLyuT
XD3zcjahakuLgdsW1eVp7UsVRCLFcJzNgPpKazU7sCNFXlP/E0lIFzVzlG6/EOzW
HQuRjA8okERKc/Gz1Ar9CoigzHBRS9/YFMVnqKNdYnu7xITxfFXTPlBaKQI9gnC1
vmHlHMlVhDvaRG+7/oD2wkJAUPSd8dLG0Kuxl9v3rUwPZRMA6r0ZetfSwo+12aUI
i2+MD4A2x3ujQ9Uux5DNk5hdmRPqMkYu5CHzQCN1kWWTJ5gLzfmImT2YB4dzd/aN
1dyMPZ7KrfXYhx/ufmYA83kh7XQO3HmoRRGTOJxKJ3/xUA5gZ7lMWFyQRaA2/BlJ
peD20Kd1Bxt95TLWrXbM9kK43YJBkgvlx3tIsqRFk5G668IhaJSPhjZa0qoqiqc4
S3AJ8kkSFBDXpYIyVoobjp2SiWWoHQ2MXCwBxXi3Ab0qq7izgzrW1Twp1a4ceBuf
F+HWP+mUuT/Pb/2OH/NTyhoeBMTEl/ipc3hcnhAr5yViU9misfN1X4yh6jnP2ZbW
cQ/nep+6N77IY+rnXjhXQFMbWx+bbIE0SEA93M356TdwlHn8zmdKm3nQIGPAVvL+
o3KgJuWiwuVOSbOiLNk7xcfLhXE/l5w2EAnM2+1J6XEe+uawHbvbaiMV9Idjtoe/
tBiOXMyuAHefHnQN9xp05pYYqI+dZxRqe0QAFZqNacHXhMQS/BglkOoMYC2U5oZO
dHA698wQ+CT3ei5U++r5w6bNdTl9c/1RttFXkLB6y2DGHJz2duu9wY2iuQkV+Q0b
muWhXVXp+9BBND/nhanf4sYAl00VJTe06jyNwi/cqcVMxvMIf/J77vyGvKUm5Uhn
F7s0ywMHT6mR5wof1zr7jNJMLy0O5Qa+adgiyq8UKyCzopI5+h9Sbn5kWy98OBbB
VhttI5kX+b2ayemrCBUSOuSVG4TPSwmEMpEbQW6H3Ofed1qJIKWKZc+eUX3aXOWL
tzymQTB7n9XDwgARSEpjNiIg2rW/kG5N0AB7i5cqugY3KfHU3fdUPigmfODjihdC
W+/8riWxB1q3EfruaLuaeSUjm9c4fXOZrxHNlV6oc52CfLuhjzGiBeYAkfhi/lse
zEJTFPUEx4GBasZw6vZEYU24Pd5C/LxDCo0CU8G15tGKl1AoP5XJYGcN4XZM0Co5
U32Iq9FAJXKmY5PlUrCq6bHMi86JcYKDxtSpBlvGiRWaD4Vz5z0MnGjlL3h+4Ad5
HBaGxjjYqcWfP0902mNhjdp1Gz7Abnn+nZ8bKqN1KPOhfF4jd7v6FFrYQVRqTkh0
jfSz1t/RrV6Sh5uXGUC1uQ7+3pduV0FaIcxvRYAA79dI6CeO3s43z+06CPlbNEB2
bIYxickZ9g0Q9JgnW9RDeRdGbjcrx4cmRXvyYX3jSusWD9EG0GQH+wOPJaz25+/U
cdA5Hd0VllsM8gDIrrDV7m2YicSFjfD7Uc51oD6tKPZE9uEEBRbFKyenswNF9Qe6
c0dDaCP2z+jpZZuAC5/B9lI7yPzzlon6NgMjkz9HBMCQ5EQwCLZwRMfUln0nEwoD
uImTbjEMTJz2X+8p02VcT2HubezBlMI6XXlZZBUfZcmvITrmbwVf0mGrsU4orEEp
dn/0TyvjJB7UBBt4T2MhuPEfr3Jrzt3kU9dBlyHJbeEfgHfbwwOzNj3sthO9ghnK
HloxLFsCTeatizB3E+pj4bO89AYiVEfdnYPX97ywdY6zWDk+o4jufJeZ35MHDaTL
qO8TnWuOoboxkc7LdLa5THCk7F38x7yhQiprOaa6n7pUC6BVnOA1+a+44G7Daq/f
4QHy1HWnKVNrp9y+kVVEt5Qu/5HbgbtBTLXN0X8indPdf3o82mm1dITTybNpYnSR
XnS+hdBfiInf0lkJUN+QZnoSmXuU1p1N2DPg9GGFfnq3r7cz2/Ma8jrmQYVZtPNE
D/ph0JWWLVNmnudpi46bgmzTD3mkFxofByNR5G5n6l28IVMO8AjLFUeluOnfhG41
Txnc2jaxqqTdR8GRy3GQNuI68suBVRrayVBCuY1LH1Ru64na9XZ2pj43R9af7twZ
ZGPVZAaRXzdKtu+zf050HEypJgwYM4PkQmKBkAZ1sh0Hn/01hrgmEHL67SgnZJzN
gs6HHS7HqjrTxJqBbKKMoX0Fub2e8Z97XAEMlJeVZn2aN0LxR/5Vje0kCMRI/nW6
Q2mwL2R36+QFinanI1M16oVHmsj1Oe1FmbPI1mjQnrKsU7W/Ju5Ub0gwANuve36o
GMS3ftEohhM4tYvBiHlHaNYi+NQN9I5BUElCeUiHfTeDtAXTu+hQTTYdXiEUjLCM
OQYDgWc8Lh+Sck7E18m6Wt0o7U5hjnPsNgWy4xJmBeLgbhirkasgFecgtFpu9Dll
2LxeU9+x4oCLpAgeg/vuEBqug6Y78dPnAqa0wlnN6WqdzTofqRzjFvRqPxymRQb5
OlK47B9Vy6BRqO9UFhW852awsvLLheetR/NK/4CXvi49P9MZOcAYIdPgajDopzLc
o2ZyormJTRbEyG7Qc8GxNYBplOpQtvrDiu/WJD50RM3al9VgSJWKcEVEpc4QkXYX
1vEMHcTinbLQsdDiKz4HpYiUonAss19qH4A2fw7Ll+w3dpZ4RUNsxCYBeDihXIaZ
eVHkYtgBPvRNNjQlvGEngbl321DEh6m50eQ+OIDWSqftc/93V0Gu2EDX81XnOdAi
GToegNRHxE109Svo+UxLfLZDZJpzxRpNHUYLEM+5kni5s15I3vLmz2DcOs5JKfhs
NOnHt4nc6tgashyl86rVywuCFWDaKOKuDDICU9eHaGiBoCfmGYHYqyr4OBb7vE0G
1hOb4Kle8cwUBMa/JAqjQE6QhcstRrwj6Axnde9DaMoGtIrl5WgY3YzZLCDMZVbl
4+7p+EYEnoqUHKT35y8AtXuF+/eO7vAt+5NqVH3NW59dQvWkDscp590HCyzkYIlN
vORRhZqNJAmqLyXsApZUSFziXW7xAHIqvWa1+hri0tXby70tJzoYirIexMoFHNI9
/L6M0Ve0E3Lu0lOJEDc6QMXywoxSe/B+f7ljRETvUrtnxKSyglZz7Z8locj2COfQ
+cn26HprmxVFd+LAn+cIiBekEysX67K7fkQzamIsq2i+Uf3/vBrC9AKNhHRH0ukF
o6Jb4Vk/ySXiiWqGmPad1H4VOVrmTt6HDBnVUBB85WF/Bd5kqPmuzHGaGQeT+BlX
CFQ0Z/CRb0cpe5bjWVOjhNCd6TsRVydZOOxpvM+nhZYXLwlBIXrtWss0oxKswNrm
5YqKnHG24Kz3KGCuxhnsCf0pRM4JO+mQ0RFZaBI8LoQpD6TWCl10cBunMimUj/hZ
7On8sLImA4xOZPz1Cuwv5Kz43+nKpvHVVMvnb06PwlKHi8EZ+q+Le/y6McQQgAcI
gA3woakSk87gWXgk6ciOLwVp6uR8Lu77R9ZouNaDgxz8yoTr6ijsWzvX6IyMwjqL
S51c3jnJWDCZKjNrT9CYZ3WB4oFLfsWL8z9EBqzftzkaeargvpA7EV6oNRHf7irU
Kl+kY6Ghtn6hvi/bLpFdoQi/Qhz3UJGaQ/dS1bDa0MyqRDYhExySmLmeFZdnmKSg
SD6XP4Xqx88zSXkF+FGdVCvtY6HuH39PqVzeu4yQKZlYgn5InzEGO4tbPY3SSrPj
xPIBR+4IhtxJvOvyIsW61ZcEYhwbVSJ6MalXFIS/3baj4ThFKoyUtazZDkVHBImu
xiUN/nm35IWTjvbzKTu4g9RREg8oA0+Pjd33JotHp7HG8JX4VsgySirDlOVz4G//
NxKdLgwzqu+aA6s+IJJqifTsNMrS0ySW1SbW9PV17+EGqz9bSl/6mmHkoANWnMsG
gY+z1peVESFdVGdv0QVUDVAIXXXezMisKy8XdfnVIA2Z32c2lQJ/OpH34AdUlHfe
cEo0+KvVuL3PT7rTKQRVQtAuY0GlC1eWWucX+eN1yJV6o3Jf7qC4ddbAUhQ82TX3
OwxdelozZtIthOD2vemfW/aau2m7THFm7Vb6ZpdUdZvQDSS00JUkyoQW0pBNm0lQ
zl9HZhz5cerBCp9jEGE2Trmu1HiY/hICYOPa3pktQMESka2tusuV7T8BwLU3yOiR
657/976HvEu6ZIJMy9vM5o5JI4HOP66SzF/lwzoC3DCnCYpF463E17oSewHSK9Pb
1B0sBzbddryJrRV75KEebDATXdoG5zbKgCsZTwR0DjqSQPwiuH8EPVgBghi76H59
lWO9pnEBTnOAyB9RTq9RfIiP5DRL1QS/VI1YsWyvmjr90XQIF1oLoVaPApj3cz3K
i3ncLTZBwDeUraHSQiAfsohh8xtXaBk18GXqVf9cdYbuNfVvmLvUpEeG2faWTjDH
QDAMk0gHbzioDehznHzDuR97FDjVdisCE7nLpOBuU8feU82qUv4q+RZk7EQINnQ1
UzHmxAljLrs4hzn4bThX+PSQAzicCqUQjqVHPB4Mt5w=
`protect END_PROTECTED
