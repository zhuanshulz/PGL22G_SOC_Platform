`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zdGHr2FPD7vof5aCgawIlItXhr9/pmu//4Z0Q5y4wgXAMm68I430AOo7Iz3D/YW
LZnl7teXGKn0jNTnFJJLguzO6ePe2POlwDz9m1817/zAabfa9uNM/R+Upmq/g5Gj
5liEf3iehl+PkIPTMuB2WgduOObxL94er6rLwTCamWVA+azo5Bxy46yP0EpeyuaR
1enthWeWwEIZgZ+tcH1W1wjCPvrgB/qNbSDgRh3/7UGvPTnOmZQ7hyI+7292HtIE
zrfUsprw7VMpdxuwO3H2bw9xqZiy1DS1GuZWpRT5bVPtCCy9ANTbax0dixXIQAr8
AFDI1JLU8Y1Anag0zMV75gewiguXIg1b7v1r0fp9do+WAuKDwG4SRAA5yORVevp0
KLhqkQy7TVr8Da3geKwS/j7iL4/3XoD0Sx2ayjpXX980BXxjhpSYIW1vQm52B9ZB
/H/NjImiDup8LX6193jMKq3ZkN2YOn3lYqIaKFswE83A7qfcE8tE00j+Dy1F+D5F
xEoUW+3WDDW1ZqUuZ0isC+QhBm4WGFCQpw90R2sVX4Awcr1mm1m7RaJCPWZ1oe9+
050Se0Xg1kiKenuxBoTFZcbtCB6uaVDwjyACZCy+BXQxpg+NxQGnFWtUShTHbe8m
+ZWEsMhVHrOw690i50OSdw/jrAtsqLBKEFBgBeXZv20=
`protect END_PROTECTED
