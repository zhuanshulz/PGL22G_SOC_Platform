`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7jFntcO4LiUy2s+zyPGyLp7SmN/p/RVQtbMCqRryB/LAFM4t0rRIXoGovcJx+bb
XHY/N/5iU6lFPvixapeBs5GPeDU6wKmE3TFnoPu6uCk2xSmwVsnypQd4vMnyNPRC
C9Ai/Nx7TN6w04hdEgsT61Jn6917nMmws7DnwAzL+igJ1nD7xVp0RH++dDMMNWqg
/gWhqRI6zB7mtIbqrzrlLO2+gRmZDNin1aP3L3IGggfkdZmUgtCe4WyGduPadJBb
AZUxNbMu/MZ0JYfNiLq9ZrlGvPBEBvo11S2z1xeOu57jtWK+lo835yCFRTQZXzPd
RRXNDOCoF5r1Wq9+CUlzgsT6IOc3lk1OUYpz5Mbf8TU=
`protect END_PROTECTED
