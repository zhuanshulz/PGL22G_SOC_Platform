`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfm+IEsmk9KQefoedsM/tYLJabY4Tr6tdrhu3ixQcka5t7Ag5pf8oezhQ0kZrXnZ
5pXugtjmnzyxSO0zVdgElZ51yiBTaKFv31AScbXnVmFaHPMbrtyvHVE/QhjdNVBn
qh5fQRhHOGSnEg37EJbst0jTj+CYQMUhCUzWZiPc4UXfe1tElleRMW8DRO1V5YTk
6gXim13B/R175Lc8vlkZYv0x9Zjk0AgTXtKtQ3Ijt0EWGkmF5pagpmy0zh83jy+o
9pdoW7jYqae+zmmmH3R6hObUcLNKhuc4pbgnr/mOYPZw3gPhClOxNDYbakbbc4Ql
nNRV2r9I5t/UdE76jacpqDvf7UPHwppFYxu2d5WD4aiq31z8a+29F3ARKcnnUh7Q
sYWTK0Rruvjuy9TdRz6HNvxoUG6DrgMvSh8gw1TIeDuRqpyxXtvdf5oiz09TtVui
O0xWcPjyiM8/d6mGP5M/MLxqrZB2e+GKmjctltoFvczQ0qmJQdATNqzUWXQgUGYv
1fiMogfp9XpuyT0ODg6v3GBO4fMauFS0JTuNuctIlsCfmOdicxOHcYUtxxN/S68J
rrzZw0SiPzD5ZFcjjv8+tfaklgkJwHPOqBbku1oJRz5Ry+D9/QskbUeyuYdWbBXZ
l1gnUh4leIktdYnUZGqvsECgnoWdRX5mw2OhfpgeljDkIPpcQMoEquVBgs2nLCiE
RQ8VDVVr3WbHI979lz/CJLXQ5Uuo71a+NarRfFMjdVFZt2Ni4tTStqt1AqdDTGzA
fp7PpPu7nzM7GatF9w4aoVwYuylPcujuISqe2X+oOim00a8+f1MHrq1Bt9bTZ5PD
Pun/hbhxJC7d4pkQuDVSZcsESfYKquTKLssfUGkcWWMVQMrsa9qTlspoeK6hdURN
T8Dba09Vus54i1q2yIsqPc34BB4VqguNSpb4MbUYuljgGvYcAfbXZQGPHkdnqo+A
9OhcVY9NzDFJ93v16FFDzyKjnP60U6IQO7JlRvHRWB7uNZZo68RuqF8KAaeMnw4U
i5MK1MeE0LsxCc1PwxPQXzKW8cZOLIBR8tK/BR0cWSED5DKWVUcADypAXxgOVtaS
AY5zjtTO1qcnbmXF2my6Qld/bSShfDh8z7XuFmH4PiCMiz/0Og1HSS1AkgDbmTVY
l6XkOKnLMeEMd4W4s1bJ2DdkPtxK/c2E64iuYUG4FPVhXub61hTk6+aayDCefvLd
jbw7EXyv/ys2W3sTq8Yh4hhcPfQfQT1uDhFhdxZio29GRjJh8dFU2sTk/DxTEed0
h3VL5KMABVSMDDAEJWZxaMBam5zyiZ6gauXwRzhXJcBmdJe0MgSiqA3mPcbPIqi2
l9iSDzk3m+BO3/K6UU9OmnqfAJDHrF20vYFgpaujj/70Xz60mDXbXVMNTREYPfrz
/D7VJ38DachDp040eAM+SPCFJ83y5INUhlx0YM8zkbtm3f7ttZXk/t+8JWbkn0nT
F4sNr8pKS+nuTUWlzs2kakM5VHOyuR26Y0+FmgsL5OobQJfsI+ZsheP7o0NjKTm1
m2LMshG48SZfHPEtu/bKXDCyGubTxgWZWkc0S1khYUUS7Ypg9k1mNkXsFBqQo3/c
mIKUvwyb6P6PvyfqAZOEHahLuI+lcTkOLGzbythNGWU1rSt8e3r0TfeTirTnKyLV
qH0GL4+p2wBxbRqSpNglSMxsnI1ictMgSElCregZo15Hx8FBR/N6eVWYQMRFIVGi
rtyhMPjD5CMamtYx4SsYmDiOcW4ZCE9Mozl5c+8cZ/71p+BZM3qObsOMMXp2RC6J
jTBKNG55oh5CffBP82SdrxSCNORO4jLWsKy3dr6+QQuweGX8xxwESwVrvtA5cvmJ
69cjwi37jcHEvM4+vkhx5N5NNTimwTfubcIvoqzS4Gg8v3u+2HxdhSS5DYrfZAdu
ph8ptZQdchFoPjHT4L2ClTuFzeslIq4JGQ/L1j8jcGS9UU4P+pnV0mg4vdONAOB5
kXlS08+pzGsRDoVod2AXCDkRa4YhrFr7IyoDyZJAKloh4R/kwok7SU4BNKFsuMME
nh+h6oTHX7U7hraE4CYnyNzK/hdINQi9jF24WvmWOKkbjdaqWVkseU1ErnXucnte
lRFJ8AYm27UUNCO73LIeWnfPQUl0lZylIxVgLp6doYJiyxQgRUpsLe4oUklyqnj4
Tf57yeMJAHO4bS2OtnF4YCYL1aqArfZ5l2dGAyIDhHFYrwW/0EPgMf8YbJwjwrK/
+Bx3Fq1dXyXygPuU6JLwr+fflmvW+rbR9RhxfljCXfYX27Uj0cGqMpIu65e4Nqhf
J06pFTX873rAwjkBr4GSH3Z1y7VYb1e5N5ZOCRkV2Xy4RVHNEjjT0rrdxawD4UdO
tOYimis5TFnAHaZGQHMGdnP7+kg11uNgLKdSdUnSVvToybAkZGG3wQE80f6pGgoT
V3sZoA9zI9y4mEmXA7hWfjcEF0WORRU2PJMFpO3Tr+YGYVScpBIQF+tCs9fXBZBh
sy98K641LrbfFzm8ogm4CCb8Wh0jTIcnA10Ts7/YRqeH0MvtTLcaG1e55JFA20vB
f6xCAOyVkBQahIlmLZruCs4Fw2r6p7dl/6s8ZHdSM7f1xg9OGZYlx2P0bg7FdwZx
qyqLpAWHEF+88tgb5VvEvlyYPSC58PP2obacJ1vYw7qtM2Vdc4u4bZe47SaoHfT/
NZToipR1SZIganf3U7kh4Ug7W0l0nPebDBQSUQTilDRuGm/PAzzaXpXSS01GFb7+
91B/onjz2vA5lI073d25oUNRF4OvldMbCXWQuhuBK0K7Ttl1/oybP7BtpPJd5Uk5
NIJ6ej+8dOS5V9PZwN5JaI8/dKiuBLEOjuc3YRWs0fQp+HGAbTZJHZ38y5unN+HL
z4rE4NiP1Es9E2o01F+RZD8KkHInTUpEtBJZO1SzE0qwChZcDFmTbKvy90wxB6/A
Ou+ErTX58k1/7waNF9ZjA2SJJqhgCuCdSCq4C2h18ftF0njsefYgo+tTwIaDofku
KfZbksGlf/1ccRCvtHOqGr4PFzFpgMOUSzRKfMF0dfQ0Ofda0zE3v45meXLxWCVQ
IJWHNf6q4Wjbcs8eEjJAysFGL1siCCcEkujKJdM49tVRVcyC4RWZ0QoLN0MzRjMD
YThHyOClbrnUq/9If1sxAekJd42mYOjvyU8qU26Ubqk9Gc3epxXFbo4oBrQRsWWg
L5REmebAdacT3FaZ0/AVXZV2/5DwPtg17CFV26omCiaq+L+ZzUoqgzd8al6IgfIJ
a7ySKOFUyrVAozNpr/3RzPNI6HP+33x9eH014dc3w7HSP3gosXJDs2lxRuA2yAYm
kgcsPdDz5yQicII7v5C7fFrGarnwa99IXBkt9W2c6NjOBeegC26vz1UP+PfKbR4X
CYDwzh2XpsrBuQjJ3cfhM4sL7rXEB2RYJVbYIP+736ZJzHVHijlW7wYeiQSPhwAi
lJbMsbccVFsWfGUMjGQXaqgYRGtCBfdURNmqZ6DQ3kq+p0qw/41ihqhFyCc3CZm+
ivoCKQcVvvNhpVXpOnpQbg==
`protect END_PROTECTED
