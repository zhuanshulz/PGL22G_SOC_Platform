`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij5N+obPEgEJMLpRSqP/ttaqtoh5Pac696klC2dljmLjeXf/3Db4fd3HRjG1yImM
wc236NVdYGDIhVFwPo0NCUw9n9fum1cFmsnm21HckET2eVS6TejqtQz4TDyEEtoX
BVnOtZRCZi5DSe+q5w5Dn8ynYb4sfwtEkMv4oHplfZCA2kCMsvRYygLhmixELzg6
FZkOw9Tsnq4wJKzNOEmENUT0q2RbYiNGjWB1stCWiPJA9xEsEsSxKfTMJ06/WDbI
y4GP6xij9c6kb7E60QymLsKH6991Xj+XAQTDXEfVUPj8G70eWFudwZmOA+o6B17o
6udaeYGo3PV/7A2Bh2V61c7/tv4i2iDPdndi9TW/cMnpGKxw7JV6nnPK0S9072lu
f8MXEWwrzNiqGTvKEUF0n5L1286iZMEBPpS2CucawJGeQmoq0AmyxCEYWMOgaWFV
zySYTDtMRdU/erLJl1vfNtTz+noCLF+/hCQ1bb2XOapnnjLsEcUWdiEMBcxxuk3V
8uEm7ny7MvVzAwn8yX2IbXIKonLxsud/T1Bac6U47iU3UmCaDELcpZhxoE7a7v8/
9h0Dcutkya2QPw21gDDAf1oFR86ld7Qvxfr6WlDIx+DnQuEcHdLOrPnzZVqudw5s
DoSAA8w+LkthITFSx8G8nfuLGuTvAlPXEatlnTvBkkFhkqLqYEy3YJVU+vkZQZuB
tYmmYtw0xm97p9Yh3wX24/mKzn+qYZeFr4tKzSUEfkEov+7MKqchxdfUA+819A4s
BoO847MkzkP+eeUyEvDwJQ5Asp4rr8ry885yRQ3PULqvwWlAZ4sepa29lncyMjfC
vTE468yIijtqyUAETWiw4j+EtHZvBXa84pQ4L4+d6PfGxUqWobWSVEzkuJEsP+Se
qWQoO8+gjX0w4Oidw8XvsvMsWjnzIoFmhg1bCur1hd9PGbEOGmwFnMjy2jIUM2TI
wAfoL6GNQ4muzNosgeqn7E5KO8WvKVfk3zi/am7N8jq2q9W390kVgX7p1dEJxe0a
oJqNUD0AUv+I4VjKEcMQHPcpr1A+se19hR3ubuSka0Z3JgMPD88ZZZYk87LpkDK4
/BgBlDdNbeNIFs2f85bZz5HgymD85XqWOkHMm7kRmxfNGCq77A7aYl8zLUBl9hvT
DJdifY+jo2aWOaa3WpwD0rjd2/nZUzw4fgzh1mkTN/GBi4lBOyo8JoFrqd7TlShk
CSXiW/SZNrvXTrcwlFcpC6ndKcVlxO6mchnKD6IwiYrjZOTdXnpuACfsin/nO7bk
IVz/j1OQyGGCzqcGMMXAydnlVonaXvb3xfBWGCCIPtrKI5DbK20zaD5CaU+O4prV
1AMnBnAkCUCo1ioZ/p+G4k+Lmm35S5vtiPQAC+CYJ71SuOSE8KjgwRxUl0U9ZJ1I
7V1xJEeY89JnsOIXaOkmEGW5ZzkHym9xxyYiYhVFnPYYJa2FtJu4Bzx8n3MvcRTZ
z3rCI/MgFoQvO4e0WUspKRthMKmDwqtA4Zxz4DbzWNNM/wbkRVhDIsp5a2jrNbRj
XO7i/1n6v8CqeixEV0RJYJKolC0Q4YqhLIBZLzAfMgJn+HP3FgeiZvsiI3ZWgbDr
P7YvbB9L/T3Ze5WdnYKfcIJZ5FQ2XrVyz6pAnge2ldNzkCxqEZFsvQHbRAXjXBkB
R+Q1tVURxklkFoZm7BUoKSbyX/k4WQANKren/4YvFohCpAN5aOQJkio9LFOGWQAp
N2mthiQ3UBtmgl9UaQUDbyw5NFJ5NSDjE85RgF5JSwPQ8fgXXs95+yXzcyB+xK6W
rtcZR0KgMBCsO50hKwiK359op2DV7v2SZXhWUjBexThmV3h9nXRm+riJNKRkzSAV
ryg0SUcqf/KFYPC7+TY2AujQ4E1/nkk8FavaEL8xA51Zg+S4d7walaCUJfWqVHdI
d538fav9wPOi6uo6seS+VLmQziEKFMynwiHT0YZsHD26fEwKTux4UL3SC7P+h8+6
4nEhO62pDFOlH9X1oIcx1O8xnQtC+4NUztSEXarGPeHQLiZblLICDVTe4L/FuNGP
sN06JkHNj6oVa8ex3WfDb6C1nYVM4WY+bb5ox1Fi7SdHcEdJlDPjao/WX21mZonC
ecz4f/WTjCfCAqaG+1865a7g6M/rs1Ktio6npEcaU+anAk5LT5wh9dlXr/rXqgJe
uMBAep9aeYhWCMU1NdH8qQ9ioygLtTPCUTn1fSMbyVBvaf89EJiW5JteWOy0tI1t
V6LCJzFr4FjB8TcmfT0U9GJ4aVhNJyUqfWSGuyT1PbyPBVWoIzbKhZ1VDvL7xn6I
9YhuHi4Q4Cr8y/rLQEdJ/5kL6eV6KEDdhAKKqUv1Kp/pdx8tRotfyxwWZQlsO7Yk
rElCWmoweO+WY8/V4IFlkVpuGGudfE1Mnenso5LE6Z4WL1ICF8/WJM0/slzjuxrg
7qYbrlaQhVG9s5iMaF6RUqk8T/yozYqbj5odbMkxx49XBFOcdKDxMTUTCUxIRPTl
SBsoy5LVuKNPVGBwe6OG2+mYujoYZQqorXO3w04hauZR9OrATpuVda/VEfrkjhoY
mqej5Kepq44leGALqJWuArqjuKfViXY/cvUGbEOtdjNVG8AA53jKK9dohAJu49AH
awbXF2LCtQc3Ep5kroVFmLjXm7+DRh2pwqewKHPCNZCVwhluIA7yAqjY52P7ULTN
TNDErM+YuXjcFjtF92Y57wIX944OtMQUVmyzwkFVBI/IfsiXw8eQi4+YBtCrdNXz
Y4YiKF5pIj43R2whOYdiofwhiwsKdBrqBPUmDUs14MdTmcMYXM5Q9GLx5Ni/MyP4
8xF5wKsqDWQXlazev3bGsz4wIA8SUb5zi62IzRWL8WONPAIYLbp8ttSVL2ROCAEY
IrVT/siHGUdZf9jd586bmMX0xBkn0DodJjc/x91LVoKU0zJB//DImLtMu2cpcsXI
JtKyc4DYvqLZKT3qk4aYy5FhIa0Ogb8Kp4+/fc1P/0oQ40tzFvwK+2cgIXv2RW6t
9CgnsxU3S2ZlHnOUkkgnGOk9ZZNP6vnYCPYSLo6cQoIVVsFn+xkHWEtxsV5TjP6D
b2OLMr1dfhEvGYeI1Oet4dPEFbcAEfjY1H2yVRBgOPOIdyWZB3WDmzjGeCtei0Iv
KK3ZKoVxJl3peIppvrEjUR0rMOunQm9/KwU9n37kFy0QWKMcvnQbN6mfuHS7lpxe
4SwsA2mlFi/4qn1xttIkhcBhtUqVutiQqQxQFDLfpAiM20Zbrp5a1lcymhSEDwd5
6bkKJH4KdYXq9rAO+mrROvuDpLyUQKaM0c46dNX6mXkdaCPFKVT7qmvQTLO8aQZg
++WIMvODmqCQLzblfusgesm7qfCmdtqFzGJUoXpilXGTZ+4EMwW+Ez/NaPcQr2CN
2rpouaF930XGKWWjYOJdkiJChdguolo5uxPdOoBd4yqbjuCRx2rGdu3Ljs3zE9Xs
wIAtt4tQfcKiCuMSr0m6q6VHUD1LFtNit6TGtSTBFKp40UOf4S3sQSRpAqOTez0b
qcnFc8I2UvJfmK0CZZybIFRSyXf3HDwha6PP3Tj59VNg8SYknHx8zhZvejx8MtQS
5enVVmho1G+noZ+J7hKKioFZhetugAHt7SWYNooMqJgtB+jWos0h5RGKyOpvdrJt
JBc1ttr8soqgRTxjnkgf0AaNeeo5iN4/O1GpGSOBikcbY6VNT7uUyaAeBvnxhFgy
EV63Uc3o23o+Ux91yKEGIpE0n9C+KEmC/hfvh09iXGKr1lugpsHNXpVn+JP0Nbkm
GN/7ibzNPNHrRoXlp+jS8/T/uHPAWBKbf0RTzcJVWpSOkO7Xu5FcFlTmRG6ofuau
EZBF2lhS7gXZQVxDZouRA32V+SQuXvLulF8nReeP2lp4CX9V//SeBVTvJlgjN4ty
0rCUF0LRCEEhJ6tnjVLdyuyh82anFXrk9hpalkPZT8edjz6gUp3FQyhjL/VMudk2
L7w6iNy5BJ8+iuctqecmf7nqqU5FM0PCEJLnv9iYIiJc02+gUe2n7fGY/vn6Etay
SWY08yNNGgMzpHBx7AzylO+SrG761SH9B+TrSASYNlZYPzJxiV5njiy7jZv5kpIA
R2bziNCPTstZxGDhiVIMj7Kv2SpGhv5KGDgClxYisxzf9Yraz42CgalU/Zw+kLS9
9aNNdIoWrh20pGt68sJuTIv97GgQNpzWaHYwkfH4LVmeHk2hT5K2mkgH6LuYy/cq
f66KzEDGdaTRDu9h6s8GP2dmnWH5mgqYGCNxAcxPxO5vVAmNoIJfNn27EyJlkE2z
XYX9JpIUZKAFuZKQaPNU2PiyW9JRQKlRungFPQ06UobiPOcuQJ7TbYIs5wsanbyM
tRZAC4xLp7puuTqA5FWqJUrq36SMva5BRnu6LXFGF8I7n0JpPctnyBSW1E36CwkX
3n9wj0fhWerVRCkpdqJxWzPCT21eUGF6M2dGu7MeEusmmkinT7oeSURUbt9vxb0S
fAofvbXxbN6f/IzvGJYHJGQ8Cw9Fmf46rtySWFs8w5sSmqEvCJ5kno8c4J8YvI5/
wTbdBUufqLy1dA5TYB/77UvD79wQeC1z2tw6uO6Gd7lC4elCoLG/bw1wqpPCF9LI
vj9BVpExuhwuoWTQTlHImDa75pgaM7aNED+CLkMP/4yo6WVPqqcZv6fG+oFw5RqJ
7yI25nZluqTqIfk6v+nU16qnVhTiwu82wMTKAxNf3LrtsVAvC8qeNOEVXJmoxZOH
aNbYzPAxZ2HCjbZn/H1PKmgxwhQnW9auXkoXIvBiJjx4xAH+40s6qOw1Su9U1EWl
cfu60du5u6OMGhnBwDHtZvNQsUNvz/ksi+1HxJYlmiytzsG7dnUMtOTp3GcXIiSE
Pd4D7842vUA7AdhhJT4v054ZSMR5D1K5uZtj4yyu72PmCpTA1fOiACAyYLc5eIDa
RZ7pnl6eOAW8RCA7PGInKNsIDp3LT8pUxMMgfMYCT2ivibetItM6xWW47o34/0cM
iUE7O6HjJLdh8egHdVPr8Gn69TepheY9SvmyYiaz83aHs/ch/nJXvYUSKMylg9Xj
RavccdQRJ+JR1N9/cTzT1aVZuqmxUilz7NAuIOc+xzKZg2qGGE9N0Y8Qf2POg0LI
Lw9WBB4A9Goej6R9OV5VCi1/wkamhCfiYspqc58j7in93eYT7yHyZow5Bi6h6rXR
NRH1v0rBXa7OBCVAbjkS6eaGxLe/N9xtfEmTiEl74C9DWJhKK/AGAs3fSf0sDZQg
TK7TEOCmtHzAjaOls4Oo1o9pGW7an/CzWRtoDCfYPv3g/bPqsoG3igEgyPZ9KQzt
f5l5hdV0vD2My9AgnQ2riLfwV/GNC1dYi6a5KN2aB/aeJ2gShO4FiGs6D4kHnCKY
sj5sTGR/I7wpa5P9e7fcBcxLCKLcV6ApaiB4oYjATqLrw9ZlIuP349o5d1MWq4BG
5W31GUfOXRXJRBqdeooy8BIUkIHCAP2qjyvzARdJET0GVv0IRu6EjnVIrww4Cg1m
3+R1HixFFpOssZtoNLDNhW4q+H1C62y6nWEKrP3lzH4o4R/KYLSv7T3a7HwIAGlI
wFNRYTBDEFCaLrUTnKW5g/SF7GBgzytAYxvuRNTwS//SCiHp8xN6KzZI2P6RLxG8
myhgtrWCiuxynkbPi2nkq5Lj+y3XkuBE0Ll/FmgArdvVhDJ2R4NlugGiwezpIHId
o1YccZaPtpfhB12ev+ZSQ6DdhFnXO18ImWN2T5o92ACucCbvdEqY2fBj9qrFKtQs
T0RSYEpoaQ1Fs1Jt1J0/stgrlQVs4N2JTgAidYxdQ38+MJPrr350NKWS0ll+83Z6
p+LVP7dDi07W2cY4Tjwom1ZaSfqf4Fjsn7Jh5F3suIg3hD9kUEQ5Vx5i89nIJ07b
/5KuJlNC1yBOtFTVjZdPE195eDAndQw5Z1/rsM9uqPvLsJmEJriEL4KbqB8j1mDR
NwYWYxN36tLVFopaGaqvTWrBFmT0UNUGqTQ7ZjVkA/hFemDujeTtPdWxS2kcreIi
DmzLO/yTGehbdSX9Vpd9KJ/BtHgW7ShqOrVwXnZ0RL8sOPny2B2BxnBi6IHhrCIZ
Osh0CTXcLbM+t8N2VeQ+x731GRAqRg2QjgXMn8UsHzB7fbUZ80j/nny3VZZKf7FN
SDuOs57KBMjlmafH3e5gmNvzdQNXZvV3WTR2JPajElJGbAbKiElGb+XIXhb03mst
77vnK4stVo9Kv+zFeOGjTm2eNmMxLJnwxF15g3Mz44Fu/sP7FdmKtNMvVggZitP6
TG4Or4IOcxKJxGXi3ElADj0Oo+cI65tulUt0h+sf3gsnnPek7yl7a1Qyj0i/6WGV
l6kn1P6QEA/M0SI1MvQCsWoTQb/StHxx7N4jhCXyZTyklFWrMrW9pdzxlq31LFPL
mA4mP6UU/nNKN5g7VDBKGbPVdpCV0cFvF3hi32SaZRIbWS2K3FdAAmwtkB16VTrT
nybwPdAqJBCGOTWeZ8KlJhqwaISJ0nadh5jDzVUyh9B/COn335OyUJeDcUboBYkJ
u9qc3rnUqgr+hjpbXqVg69MrPSSkI0hNaO4TV+b06BugHKN9Oo/i30Uk3upjML2U
PlEy2A4WzbpTrXOaNmgqCH2RzEIo0b6MCBYbgp0jzV9dVWXBdNRPrcqY838uyRyR
ju2sRmmmqHuZKw8kvENyy51KqKCzGtd49tvJy4bme2m0OrLNtKWMlqLc8MtAV6IB
6W40apUHtVZ2Lp1VHZ/CY6jfC8Iqz8xSZyImALeSOqVDfTnoCx5esBuZnPCOLyC0
z4JmOsKmf+cwlQoToM4iooIEEhfSUy3Ep8EG6/ZHwQuheITjSWoyiRjdL2v1/FTu
vctOe1SsvdOA0uBYgAqegMlhJ9X6fYPIoXVmTXbzl2hY0ey+bP5V8ssbFsKB2lk2
1zzFkmdImulQ4pt5c3MKFmq0qfsoP/csQzmSq2DV2ROXZuziQwFM68TSaoKBZWYY
2lj1OIYePyFia/YcrimjLm4QncdHiHEdNnA9o0VnFQOqiPb+JQLgBkSMxnS/YGPi
ZT7rBi7DEKEyh25SagFp62ryyUfGuhK/NgQzQQTEWJ9JorGmwmn0v0iei+27iIcG
WkzIC2strat70zycg9yJk/3fNIGnKC8Saf3onfAon+ATNLlICxrhyvmbAcBsZu/c
2Xj8KBWPH0DoCoDAu3w0EJV55HfupqPeU9x7C2yYEWUp9m+6EKuuuzaX3ms5oA24
7Jcsof/unR8hrxBEEjtepbgC7FzZpNAotC5+KpDLGUaCoAFFe4AfqQKHWoLbAlY/
reohFwSVAgmHk+TNJHM3NoLhzw1JKGgRC/bTya6syLX0NK4RspUZOhK9UJLV/qUa
HZ7qioM44vh3NMV86bn7EkU7qkiK4UogD2TPdU0kLV8tMI//BBv9skVQVMpUswdR
vv4YNxqSqymwEib6JlwZ16FU9cgHpmisafonpvoa+NJ8mKNDRAe+XqZRtw7k3VIt
4yGHhNO/G3gdMXOXkpyFKIZ1+zJaPnWSUsRfiDOrnPoZMnrxWtEoUPVX0jGATEUf
bosgI8XTXPdtd4omhOFawGsNJnx52GC0Vx8k4xsoNODBiPjBcCymUSSE4XKE3lnQ
BebJrXZJ3rE3SFTFZIE1Sr86HfgSy2zWQnGQ1+rxMhpeiU0317IPll7GTpfd+YoS
6/KSqXDr4D+Pedw8zlTEpsa7bjdySUtHvyYILTsflvy4KHtR51kpy9GayM8RYHQW
4n38PaUjRxPuOj6uoEiYIArfD0ev9yOcOEUU0uJ3eKHYZUNpGIivaJRqOb9F/XFg
3JfimwT9ZcMjiUkzXN0dkzSWYXi2PZYCTcUp9XZ2H2QXh+4C7ENiKbfa/Fkneovp
TG8U5GLHlwYoICA+C+yNuPIPx1GNDdEiFCwbsAlo6tJ4yYvZOvLTbsF6y1mALVem
fOPFig33ahXTqbj4pyQR/PzNvtw7B/QrEOpPo16CEIKTdthSfbhxxDqG87xpnYfK
gI+o08ygBBgKmxLLQtzeYs0YMWd+DLXhJKRnMx/MtRKhpoRHStLfPXAcqvoNvCJS
Emb2J+J33i0/wHurEXgyeLwzCA/VYjw8eyzP3zViXV9vqErgzKn9l6uCw08h3IZy
Wc7tgm/kyM0MsS7YVRfTNWaHnfn4th+0PPQcCm7aHiaXT2kZK18atkrhGPV299m3
SNpCvCADQt76S4P7w/BGdZ2ZMlAF1ZWbthmhp12ehJwz11HMl2jmdTwAzAxc0wLa
fXkHawb8byHCCg1nSzSJ8HcaExxm6UPfMArRdBThAsVLk9QoCBJFHcFiFgIuVjcr
/v1UqtCMqvw29gKiER0MZKlkjw4au2tJsQpVlAODh/dkP/qlPETelN3+T+Jc0WtT
R8mj8JcNwlJ35A6ecmIERHVkV1SL+jxq7SPbvJX4RHxXyqERlxjMRVjv+G0cLib8
NXVLcnrpzfVn+cmMe1Ikho5LF/H9WPi/S+K6teU9Q/tlSVnrx4GzKU2ryBI5x5VI
vIaLmqHdNa/d/IioQAjDk0Xxxal9TmJ60GbVg1if9D+M8wee16UwGEhiqRZQZChk
yjiuDJCW6SbXYDJzac1TMvPfNH8ExLj5DljvH+zL4d0DN9eac1w5ZIrw+tscZoJ+
ZZd7JIcdaTccJTQ8tjkpTZWVH5vQIPBLb56uTQj8/oj9WAWugjKE91uvYgjJ8Qc9
JlzIWJAWhS+0u55o8bn7n4ISWJdHFz/lee1ACOci49+uJe7MlagiZvnsuYoob/AD
hduQ0GhK/+bgpOVqFIgaSxmUvQINRww0AOw1Ofkgn3E2E0r4yvpOkHZpmOKGjcK4
jn1jTpJx8QEaEnQY38izlnQ7MCxtst9RzR2Ar9NmARTkL+PsSojrht5etEDVPy4O
7aS9AvthGSfufHdTuJVaA9QE+r0PaEduyUJPwkmk+jwreE7JVCaOtbAfXBkDTTjL
9jbBM2VZUneuI4TFZ9YvxD+f4CCJSyr3R2qVDfMQBB9P+Qy1KZlUIFm5nalgOOMp
QojcQ2/gmH9cRDxKRx/3V5DghK0OszNhciC8tHOzBj0iIBwU4awjmkHJVwdKyVgo
nRJwsCADGQvh2N/XtnGIvRcR2puWnWU+facvfRGzyv3ncrQJZieUVditFb2ijukN
fdhpzORi5IDYVwFV4sIddR8qYYMyeCtZc1+p15mTfQ8zWGxPi79AIhZYZoYe2ZTI
61OYJl5IWJbHanyzHVd7mbtxkQ6SvkqfjPYpg6eAtDPn9w6J/uAB/ODaRKLf+qq2
i1cg03lGbJakE0qTwL8OAi46yTN78SQ8EUj842Nyn9xvuUFPcZpyNpQhmtMW/A0w
5X7Rl8pwcabC6kKqYqPq2kzm2S4q7k70UzLbHxtkEKCGnHU4Dp8qeyLwki9BlCmZ
HmCOHtcnIKJDWtk22bakHe4o+XEn45DiG44BqI8OHWo0pXwM2F2p0kFBf/tW1RT4
Xez3cwkK+aL1hsO6LLnmvHovF3NbDqyfj2eY9WhP9+mOh/FXSbOHQqZoUTYMYeyf
TtXcTw7m7XNwg0DaJ0f3LZ3n1kc58OIsGyH2N5W9ak4QHdVcN5oJ8y8/2ZNSWRVN
w5TVfhK6iQkMzhdC4b4RmiNCAzA+iB358ci0/FhCFc2w2djnqwLoyZm8uKAwIpHY
MopcTY72LVhxr0+GYWXqeEckD/7Xy2JkhUMBFKOljfxjura9DrhHzjuR4t1Xvgtd
tFdlFF46MnbmK+1GrKhcOyeO8qSRZrvaGoPGdojawaIFDTDvK2lYrSkKFziP+KaZ
+9u97GVuospXA9LgNK0mUZN9u18FVkhLZGUoKFTRhEp8lSWvFZdQESfyw2YmIbBx
kS+KS7jR04xf4C+/SLVwpbPvh+dxSRCLEZogoofUaxDsy1ACzKxGqsySHgoikNQv
H99PyypabHpKPCOyAM9NNkCD62Pu9QWQbCeMrRiRtMKkgVZjdYWwrPTd4iGPnOIq
+0FM+D5zQr/lwOMYwDt7nmFQDGeCNkSvi+s1QMkaAFd9pFaf2yWYKkTaIt8BI1PB
iuUrDqzUg06xhbjdiLOYlL9WaByBK0QzguCYsBF7IzxP+5GOgUVYktvTHOFHw9Zn
LvQdFsfrT+OaUNALv6pXu9A6qKzCnEMSzmcal2zu8w5q1Gp7fkn7r/5YFGJ9fKpo
ZVN7WHTLNXucwbYf21FuPfN1h9nbjkVbLs6SYbhpBmm6V9OhNcigKPTn+VMjDtrg
paU0FoAi1em9zZ9Tdl0pVewEtjUnk/L31E1YaCotoW0+29WSZa58YPqUh+1rchIp
75iTugPIu3+ltnIVSu9d6ugH1DIR2/fSZiu+KjXAww7KM38HsHqFPqAX/JzQEIIn
wio9Hxu4DANpYcsWGBwIeMsV9DFwsOvoqr5YXfJoodpbr7NfGTQr2dqgw56vGyfd
HKyE+LWgpjbsbnJ9S20xzQHulXtoWa6yUnJWypfnYDFPKcnTUwf3kBUk6DaiIeP7
i+erMLtIE0G7K+ViVCmgTlW5aydlG5mDx+3OcfxcM8Pai+Qz4BUsfOCwYipFDEB4
bnQpUhr7ZxLoy6K4mTk0maBxiL0dgzgYmtH4zl2MorsDikmkujKKQDbjn3Nzw3aK
/8E9RLWPlEg5KYjRmAs1ag5iXoWzgVlYRz/XAeBjqUGiNo39zsZekr/ydHCitJ9q
8WaVsUkf/Fl1v+QPxSTVbsspKpbopJu47rKAEB8K55jf1mmx4HwTrN/i9L2/Sshr
c9N9zMSQ1MpTAyTcbPUoN3/srYo0a2GzTGFVrgJwlTU8Fq/2Q2LKAdSYeCsRKsLf
aG9k/yF1mEcORfcqfqHTyAdq60K6Hk+H7PPQkA9WghxNrIn/X1V2xHjxAi/wHUoO
CPYmo4L2OWIIVKETHP02O/hLlkUPoA/ija3m5md3IlkcgIQvNq4rXLDyKI+iI0eG
+J1JwG1yi1Za/z5kmewxGtxwqC7mAsFSalb+9q4Sed9UUwUfkbzT8MPKwP3paBPU
zhcsCB1wJ+rp6NHE+jO+tqj3PahfLd7BxgKf0dGSJR+bY0TIzjJvPmn26UpS+K3j
eRfAq0EjU8vekZbY+vcdugkVKRIUwi1rQkahQIy4Oec28lQdszWXwGz0kf//hJkd
uM5KyqdLe9Regl6jMjzITdyrlR10FdqlllbyIQq+deEFk1XL2jO/9AMNP6rjpNOO
QLo/JkyG26EhlVwpeVCHoxeuIFwqACCtUB2Zj5DdWY/5Vyg7EmWR4KzaeWsHTVOF
hEq4/6G0v3G9EUWynWcE6hfQEAf+aDAED4N4xq3gV/oxMHqur2Y27s7Tmn+nr7g2
TyqGxad/HEWsan0LZt7HGb5j2+1AV6AAHkXUaQtY57E51OTAHo2shZ6KCGhTnX9f
2dmc/1r5IFrkfU2uAQOdwekSwecNt/Bt5Vyw2Kg8v6uWxXIV76r+N5b5SFtW5c8j
EFUk3Ust2ScxIlNOAEuU1KsennJKxTD99Tv30unrlgNAa3YophRS3o9P9ne4gqmB
0BoOPeWvav/HomPv++gVCB+Q26uqcrODVVDy8CcmzV8HRPEp7Ni0v0qUuVfzpAy9
0fbFtfz98UC2/8sOTh6x2hghVPVEsIDOS740fGjfEBkIkuo54dz6G1LL6NW8r8cw
gARTV6CBzFOMu8EZpWFoybYLM3kofNt10Rskp7Sq8tb7zWmhAYH/CfvBYX5vNQjj
ur/ifb9U/dAQEWDjX4BOiwm2CEBce9z5ddcrxWw/Tl0V92wVtkbGYnef18lkxg/6
VqkgeP0e5K/HkL8j2NojkjuWAuXQ2Mn+plUNhxca4GnuyTyguypl8H8dRRwatgRI
TjW4MbPdHnAHBU7MKJ7Gajc4ErO2LDv2V4KtBZdzpivJYbLGIoakn5r3+uaNtSQH
ukaRpflzWJqtJJjPm3477tBnl6TMpzKUmAk+kRMHkcWI8MdYwBhdCbUfbQEKb1yj
hrN4jR0H6HJo3Vmn6JAvUw==
`protect END_PROTECTED
