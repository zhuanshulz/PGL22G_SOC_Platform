`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PbmMO9K/bqWI/lqwHleWbsBTeHh58UloFTzllWIVIGiXqdx1oVWvfB0YHM9JGEWN
06z/BUOFRSIW109FcCVO/r1fwYPxVdN/GbLksALDweq/7ZQvu+8t87A8L5kwhNmB
qVqR1eJUeKQYhKemo/ElWv4mTqzFQJfg/902w2qn+/SJoRIRbdqfz32X6UWLNZlE
wlBqymAVMriZ4U3gx1N3ZdUT+AmwaApCLck8tk1h/EUc8BJTf7T73L/RMIO5cslV
7UG4sq/KYGzQ2ff5i3cyD0ZHzzzZvA3qmclzkyQ6OxP9o+aQBZN8Pu8mJMakbt2U
/++8l6Y7vXVIrP2aJ0I2Yznl8qjzZcUGDYT6RFe/N87y5qa0dOYc273F8kmtRUeD
ijD6Tg13NAgN5ppzuLIXLPPlSDY7sSaHTw5G+kVWk4vRYWAezQp1Wole0RiUSF5m
Pb+eV8KeuSHQr59Evav+OOwb85UZF0A3Bw2XTSeaGjtv+2Q17j902RtRSIXtftW5
i8xeVin32dyZR9eQS89q1Y7PluUETWpYO7raIDyxkGD3JZtX5PJ2aGIr5Lj+Owe8
`protect END_PROTECTED
