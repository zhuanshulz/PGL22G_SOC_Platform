`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLw4LPw4TwSUWvfJo5LYy/2cjmTQ3vq1nBqoVZJQIiGiWIR3J0X8bjVDTEQ1VszZ
OOERpUisDmJGlLZro2qN7/Ic2E/+R9vFOYTJWDzhLz7/yg6R1hPwoH+uIsigiGDJ
MGej/zHK7Qyr/AikMIy9Z0bJX6PwdJAnlRm69y/5MgjEqmZ6mhGinWFPuT+WBNNr
h+rQyScpbePz8fD1uHs6tWlF86x7RBx+excA1IHMGBiCNRTHakygzsVqO8gFnlmS
001cquQyQGs4c1mk9UvC215rgpMlwNGhUn04Q39Fov8FJpOqIDCaLFD3l3/kJ9xD
TQxXmRW5iS6qefyjhM6/zbGK0Bzg36KXFrUhs1ttUj8oXhmK6nOYT8LSacYAaveB
Ze7BTYTiiq9Zcc4m/P89KkymnugYJWbFwZQxy9wTCMcTPVrbdpFm+3Rl0ml5MxNt
n1v3LbrZpaf2ByeuhLv2M6vsutiYB0Hn7ec9uiTNswemi0OaitO1/ofqoqFe8URt
AEinvIQsup5z66BGGhR6zDW8wgRehcaNAULczMkCjrzPTcgdlcqtn7RRgWuN0F6/
4uZzrVPD1qr9D5wackNoPwPJ1Wi9TNxjG3qV8Yu//bjvOOZudV2k+Ony81sGOh+j
Ku2XbNJoeTRfFmetfVQq5TgLGcv3JAfp9+Af9KFWLt8RXx5cDz08g+zFqwphW1+a
+eV3LIdyzBla+xXnf/Cr4TdN23b7Zgk9XRHcBwZjccplVDjPVsoxnOvDZWTIElU4
sUo6ZE0fOODuxoiMhTh9JWo7QW1ifZoDC0uoBvKxXLa5sofk2NEJdSSZ854bLfSx
ROmmRypKDTnV7FJA+vOKbMS0aeSXLiEXy/hZYD/caM8=
`protect END_PROTECTED
