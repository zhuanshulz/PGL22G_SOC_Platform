`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uDIcHzBnWPgWMCp/J55aKn/SMNu3ToMnVzICNXjZuUmVqI6CnqgpRFxpLl+pGc4w
aWXZB6yh6F1T15lfJTm7oD1n9pEu3KUIwHEDZY7lbEAHU2+PJ+ptbCYhAWaOzKw5
a8Csi4a8WZ+gZgl1fYeOe3HKUUIjTWEz7S6u7YCyg+iG4CjpF0Gm7rd0H0bDH0W0
+wXSUM1GWe1eLy30TBU3CmX6PmmGUnsZZRreYbSTjgMK6GCijPoJNwU9f3vbYNBC
MEBKhZ8q4Fnbz3NzTaJ6UuC0Z/AOoI3cfUyt0uBVdL9AgrZXm7Luhh0Nlaa3PziS
3SclNOIRWEqXDwYwzQINckNgSqmLUPgfIcWXsQcxbGVI3pV7IrKT2s4/FiwTQ8D6
Uh0I5SKZE3D5jFPPn5EWwr0OXvIuhMsTZpOT13VuLxCprpFjiZ2TClALT04mXZ6D
AM8GmEJPcH8DsCU3uYga2njQUghAATQ83hSopuLtCtDo3AjEzD/cZKrUQbL25kSI
`protect END_PROTECTED
