`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BuBwwdnrinVC5w23hNu1jcsC1c8AOiv1ROdBVERsyK32+ATAQyjtLC0eTtzvL948
h6pEGfSBIrGGunYM9w/s96KWY/yjtOA4QVApQPYdm4pvmYwIAsPId1yE1OcRU06p
KIKL3x2qVD4kQgUItByBDH8xD0fJF8p8VPKChT7+tTzqGT9p2IDN2AhJ6W/7e/gv
XblOfURF1FFfLd2FhjIWu+8HsLgBeCVrFkpKv9S6aGClurGCE4daOk6ZuogOjI0z
l5joTiqSvBjgrNWK4mR2xA==
`protect END_PROTECTED
