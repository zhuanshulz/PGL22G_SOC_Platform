`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGIAEJnb6nJ/gy/vIIhy9oKVUNX8ufSbiH2soffp9MVFNNH0UpNnt8Y9IJhzXv6i
G6Zf3xhEgiL4bR25T2jH3Iqiu8m8rn6Z9lp8MQXehhnGePUEe6kLi/LickmM8yk3
o8EhLSnlcu/xoUEIaTWN9uq4R/J0TJFXPKyHDjSHB288lGQeMt9EPkU/Yxdv92fL
lfKVdReXo+UBqo9q42YSwtI2biiRG7pErWEflgzlFm7IvScyRzHg4wOs5ywCj5dT
NdocFLqsJwTXPsRb6XHbsm/tvEX6iYtbwDbhUKOVvQDf8Oew5ESOY7om3bGmd6ol
UpVQRGAluoydUgaCNneRVxtZpX+ybveajgcI1xBK3GprvDpvk7UylBVqeqiOvg5X
qzCd8MSp/uxUql0jEn6586+JoX0+AlQeabM8IlfQLj30v6uJBYnAsy4Lz9mq21gU
VetijFs03j0N8YR2WbRN6PXpkGbF2Zs/idY/Ao04FAuXD/Uj1bXurAosc9bmNz4k
1R5PvE50+9xCSv903gD7PitsFvc8F6gouAcEjXR0opHwM7e7Jw0C9wxSSSOsUGhE
aBiPgGTSbaN04IwtdvH8Pw8hcR6CbISWIIwC1Ypnm0c9EOHCDcw9y1go/z1zcGuU
RN/88aqDE+mxIW1MNty+oawPx4OjYgF+DXoKP76y8u/VGStSVlDS3hm6lSD0Y/Fg
4Jq7I4yLD1RqjAKdkU/WSPQ1CWd1AO8hHng6wZTwLRkQ+0nQGFHKAc0kr6SfrmGv
4Wznw2d2HKSbnopHSJ7cqfkedasTlicWJd8sjj1RU8hRnlDViFiZepc/dPK5ewI+
7ZqP8bzYuLGuzikaXN5WqxZfO9lOv1NUWTjaNJPZp12engYilqn4r0nD7Q9HOdcX
LnmB3XqUbl5eotrTOmQPAYB+GGeyF3Lghta30xs5L4x0QSL0xsv7cCNVSN0+jO4q
vWliOA6oWJAJLSn6eX9gTV5iq5odviBwS62IDAGpRb8FnIUg0GMDSYDLWQ4Qqsda
fb9rTvM24/7w+X56iqvrsr859HjgfK140o+Hpjsugp46ImH/V7/J5l7TOop3BJ0h
lJJBwBEqHWUnvvp3MoRayLzp8pSIZMRJYPjxyNLvPIQF6VmQYFYMpnreZHQVMTrJ
HeONdcbv8yzQHllZl3it+d5dCaHqFvqTrAd5DtBrQWudWn9fbkOvT6skrqXbn1RJ
iXcnhegYRI2/WxdOovpP1xo1j613xQyus/4+n+ndfRx6nKyfBVp2nM3BMRbwwJQd
ojnjExxBo2ePYgKQHIDVmLLWrxH+L76oAb8NHcE2dAX1PdJ9Jn6sroPq8FfNY7DT
MoC6XRaC1wSZDzeXN6/LmfVZCP+ibeHzlilazUiEYnEvsYrO4EwZJlTXU0EylX53
+wgbRAUO/5sEbRb7Poj2YjNtfhrsWfG0BAn4YMXq2vd/2Pljc18RLpeYwL6tT6uy
tloDVprprS7PnyHSqfRVlmOEl+7djJIer2pQpXUkCHYkrWbaEuAPibqMr5z/SrPY
Wj4Q/8U4BTzo04nawkCh/nOgyizINHFFXmUu7n5h69PzA2aMJC5Jz2/IN5+JMCKL
LCrhX2gQVVFT7ftSJmEKe7+NR+MTIBMgQKHBi8ZfHMpU5xyPCnpaUATmEiv9LW39
LRb9QwvMKfSlJNOkHyuY+H30IPJ/CIoDL0bf63TSp7n1YpaNCKrm06WAUawoR6f0
erxopAi6JJ36IOnZgdd4o9Wr3GSomOU3ATahQDtY2WA8OIA3VoGBHYy2B4u77KPP
Dq1tB1QolFnxmTBZVOfbLse3OaM0ES9K6JLYDIUB4U9p4eBj04OMijfX2GzwNHfW
hGYAJH4WROxPfbq37IHJMBvlHeg8/c3qxtn3wN6GFd32GpRzz/Dzhkz4tjU0911k
PeoB1BBtxbjXG6Je8onxVUxMX3uSiVEkADSK2BU90nu7AR5JRk8WTxKzB1zDN+TV
8w7Fgupu9RJia/o2t/4j15X8+qCichhQDoaCCarTXZUV6hN38U3UHA3SBndHuNuK
MSnlslMzNi1bVYyfQKyh9yJORpRBz/EdFFwSJOGTxxg7EbzKYJ1/4ydnZTLu6E2X
MFgmTyanHyjh8mUCtcp6SBRpKKwYE4uq+lElQMf2OO4TQf8Ddzd9WbsOu/qSmQH/
1lhaKW8shlLY38C+k7dqq3bS19P5zmNTWuFDl+ZziamFw/yYkJ01xXGlJcREi02o
4CykQCWVLiEe0rA5IgYN/iJzQadkQ/kWsZDDpvuHoVJP7q7GyuFfIDNJ/Yy1se9c
WAo5KsQv1CHf9Hc24Ea/6MjbuHNOdP3RsJlqO5KtG3tsSZ6eKAQWxkeeOAC66VNj
huCrQ4BJvAfCpfOYzeWrF2XNkIYSXYrXw2n7GHuPVWMavqFq7Yb2uMCc1qsRdYFt
mmiyx0Ibsc/x6jiy3Wp21QNE6Rx+CaG/2ccjHfkURe4AyXY1BXtnSlG+zt35iBbR
dOfFhqv8vOFS6/daWYyooaWLXyI0iDtA0O91ob3/6FPRR+yGQH0VrKmI4KLhZ7C/
yepQvNK+oTMZHegu1BAh+pjMrwHtlYSmMNqYisaLkVA8a6PP5V7iBqYhFI/YhYWY
vEyzukmLqZXfj7mnIozH9wNeQOoLo8traUmy9t4TNsz7FJ1z2eVM+bAAVn0WOrec
JB2d/g3J9encT1OXUrHcn6KuOpoiCOjYFD9L8ZexrP2IWW6a7kHN+4yZ2gQcpTaw
G863YJgR0mpDdWiY862zeE7ZFQO91MTpa+idJFqjA7TWDPm7pErfw4EOqVSMBP65
2xkg97bYcWvnamXh0y0maGjd4nKT33Ept0mMR9WHGdzc+d5+r/EgTu0VVJx4Besu
6LB0ygnvP31Dt7F3/eDQg4b0bOh0+tOs6upDCQws8AVCoOGO2lf9zC5FXlWPh9tI
U5DQlbF+FADulFq9rZPORNypAWhYAl7oY2j/S9GUt7f6YbVjqoZTX8BlGLhnqnSI
7aSnHlaCH5EGlLBDWzlBzLWv8v9ZEMjnm7JbdFPIkOmfrtrRFizCIgNXve7iO+w4
F8u+eYmDdYK9V9MQevdOIPcQrZ6k3NCB8mIB9djM0hrFxKS8YENYfea0jaMSp36F
zGssh6WcmYHoiFXbbvpPf9uKCvN+9UR0au2ZbNo05DP95bTk5Nix1kXSn9IwFh7o
pqYLGeAVlVqRbUjv28xO+TOYYBVJIJxFPP6vEGIOQSQ3xqYixiU1Pliv+nVOkv8n
miGyYe5F2V7lwkfRvpXq4k0ArNP27bOFN24E11v1HRgi/i1CPNH1y4R2qQ/lpA9Z
cNR0vuPYLyqeWZI+ob7rSc1zCZFbF8yHGED10+Mf1c+mc+ZnozddrjgC54COe1X5
xg1cWGXwF0Yev5XJ8DSKqdN7j/LJ+VvJmfMZ2yu+8peB17N5zlHtMv5IkCppX3Se
OS/Y7q/lPhW4hOfdGJlP50stUVpUjjy556yoIEVglYVxXFfpNsgEHUNtGGkRtlrO
dFodbsLPYc89o4xwwcm/e9Wdy2QgqOynMtZVE7LXyIgIAH+dBBVGzdFJuXrzEtcf
1+bCpYYUdn9UNJzCHBnsNQbEA28y4XRAtPQ8V3Yc02d2ZlUFl6Lqr9fUIWerCZ2S
L40p3pcyXtqZpUDwKV053T5B23umadi/mqtdpFOJYK9ZSFu4TODJtJngAdqp3sRs
v/R2EX58PGlgdMZZWmsjAbuyP0lUc2b7ZmiTbOAcrejroQFH8w2ODys3TKB+ZedB
cHX9PYDX6GN4u/BusN6XDg3Kjkt79w9mi5VeDLDxi5MGlTBGXh6BI1INrOkh8u7I
aOzaVSGVr0lapXPmBPclHQFQh3loYWAr8wjSjabDZCxwAByiXFpGMs9Wwqhf/C8Y
DnAWu1vyhMO7RPOp525y3/X6BTfbuicO6dysS0itz0mI8BWSMeIp1x6nWLAyC2Dz
H6FQ0lgeZcbxHBLoasYZWlEtFBAwauTMTWia832TOWWNvpzbNVwAbm75+cxQF4bj
EbCLJdQjLNQjXUQAHFPePe6ZVmAUW6IwXoPqAEe8WgNrQ6UP8NT+UBpFgB4FVqyo
rDkx6X4Y9mt80N0BJHPbsGaKPDlRC9oV+81Xd8um66TvKwlfLqeewhL+Pwsl10Yp
xJJQkxb9GP83OqzSL5p1mPOd6CPe4s6ayv1dyx5YV/cJMcf1kbQZR8Hf14+giYWK
ZAZAzJBmaUCGy3HqudxIMFSy71/G62UkltRqlHXDdxbS12s8sdWLv0HU26cx5bEo
fhtYDw0cW15vkD1LquHiNtLgKGNHm2Oc0N1owArWYunc1ZBEVoRec2m9GYWvMw9p
TXoHMH49lp3yfK0SWtV7sJqEYo+b/QbCa23aneA5N/deF/lX2RNIXgWeG4ogje5f
r+6XK8EPj5XpnzLERrYvN9Ld89juGB4DeUI5HkYEgWDd1aKiO59T13Fgd/bCa8wB
wePY33MDg13rdlWS8grSoMSzov+wqnV5GaRmVz7uC5U6LDc0s7rB3mpffKDy68h6
Gov7blCmIv2nztLnO6XBBDdIQ9AFME9xemXJTGvDeCCJkq8Q/tYq2LhG8S42deSH
A2yXU9tgaPEaNlSQdwWmJ/mZdBYlKHWoltHJZepvxEc6NxWevYCM7/EMudOKt1lI
13K/dFA9fjiMSN1znjVH2KLkVbkN/m/vCBKuTJpfL7elEXZhNCOBWwA+rUVpDJ3H
JvtMGB8tgoVWl4xmLJ0VlhpilbHlbjUejD2e8jC4T4cAbybmMfDxFatXAPJxNZwy
Qb3/uTROyfGGnpcW5ETGWtZjun3qw42RjwBRbnSudmbgGLWR5LwKA0Z9QOmFVEDq
z8tsJ/oTg9z0owR0EWCds7CRMo5m08uwIhUV0vWI21Zffrsj0+aZOp2aFQR8cXil
cpnTmE0pN3DvSqY4LlzlGfQ1r/NwS0vGfPLIgILTCxdK5pNXgmQ8d6DAyTq/GpJ8
OU4zrCaMEfjLpDqKvN0XPcGcpjWCR9urzczUyWocKDGUHWqQYZGiZPkC97J1buVy
4OfLs8P8wUMEhh8GRybN62rJC/xi2lr8aq9JQdUyi3FdapC5rFSmuNRmpJN+dZYq
Lr5BEj1v/6ddOXwTA4LEUbT6mnYafUagnu8KsYf9glbP8kEi7xlJM9edtFpvak1I
vYeSLCT/oTCtFG0tRBYyR/38fmJBBFFN/CfG3WKxCmiTmpyVtOxmLDZDnhDqFWUf
6s/OsQz5Zal7YI/DCbK4ZjR3vkVEDW2dKyneDyEh2vnN/XOkuuwYFtAEib50Y7WG
Zj9Z/w9DGN555j9PfD/5D2qcCH9EH0WJgd1qqIRNX2/2uhafKJouNte2v3V0g+/R
Nfkhv/yPLuK8URBq3TQd2OFUsK1YfZJfQJUZsSrML2vHTkXBF3ZgVkLGSmrn+UjE
ks02MhW0wdu1BOORYAbvJmSwsilRWwrlhTRpZ2XN0z3u/njedUINdiUeLmv2WxpS
7WCWpk4d8N2g+hvsqCtBvrkdT5Q5qkH/yx55xs973vv5bYTbMg41T9g2CAF6J1d6
YAs+7ds4THfx+um4cpVc6IAJmABVarXid/ETFppnQ9QG+Qv9V5xabrN4EV2xUhFu
hbKDhFMHpRUNPEps3+CmcgzZuBWkTtXY5ClkzHRurfqq0V6iJG1sF8y7+9bEwyzn
iyD5thCQM6sjO8D0JDSnfAfE+pBtqgEdqS9D80Dh8UuHs855o2KuzMmIuhnelYEI
WGN2Tma5Xg84OKz+HVO/o0ZtRy/Q/jALiQuIpMJeg2UfpiYncHzn8FMQyYxT24Sh
mLxtzSyqCfkza8WfdTqXLFYK50Ocrl8kFqHG2gW0UvoAOdJ0779a/dt00fxFrtZq
b7bGiWWtdeYy4wmQQXF7yV+jUZbcpuHppx1B4PfALzJBllN/J/kxJ3M5KMu6We11
2+wZiBaMhQvFJ6ywu5hDLG5Jd7K411HeAx/QpIVeYL5xPbu/fBr9Y2n4Ann5NPdp
i26YtwqJbZzYlObiihN/yAxtRJSw0GDj4SOdR2gszYZ7WKsdGCXC5iJz3G+TAF3+
dmniB9jTQ4o0ZhXnOKrH4pXhy6bgDH7GpJAs5K1jooE=
`protect END_PROTECTED
