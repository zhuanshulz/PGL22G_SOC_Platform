`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
05UalH5g6SSQD5CgtNhNq8bhC6Zth1wLcjb8W6icpIujc193/SfjX0XtnT6PHzzE
0ltL6gFssZPpx5n9d7aSVrmv245rQ2HBEj03Q7V1TjTJiHlU9za8mlntaAPbDDqZ
7/FifPCT3VImtT2KkkhvmLNqsx8u9wRQuc+o1iGqU+pYnE7qaS/gcf2d0YIhNbtg
cqPwu19TWwk8Ge6jU1GZTt2fNs5o5iedke/CtdbPwTuoJ+/SfYPZWeBA3pbQHj/6
5cGP40KJJYkEDpgfCJKrjRCX6POavy4zrRxiSQ8MFWylJnzENXTMFoz1VngvGwPY
4mhmROQs5Sl3kCW2TIfn7uClkW2GR+XAf3/Bbct8g+boMnQLz/gBYGmcagPcJaOR
UZlsI9FnUhxCcrW97K1YuE5cm78B1vj8JYDjD0pyNrAVxtPiJlK3nYWj2iX2wARR
`protect END_PROTECTED
