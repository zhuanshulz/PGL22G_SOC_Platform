`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FoAja1j6pUyiyb8lHBNdBl/CfirF4NNcvmj0yx+Glz4s9XaiQafCpQcBxzk5mUHN
kfWIxWnJfyjiPRC9uEZg+16Ya91gWKZc+Pu7HVkxfOfdro7BZ1je7loSaQs/ETxt
E5Qy7B0EGbF0joZGN3IzOZZnkYtTSb2FO3i8sbSzYzNl1iRXfrUBvAd2R4GMW9eV
fE+xk/ZCyp35yoJbl+zWxosb8JI/lpiOy+sUp3zroV4nE5XTm04oBuSWBjVgil+g
V25e1KQIt8xjzf/qdCQGYs2qh4Nr3ib3DMlTtakB9gr3vILHy3123jaouK4/EiRz
PeN+JlRpgzLyO40zWTgNDYxmSbd4lU40ZQxRqYY+7oli11VAsPZTEvfDQiQO7yqe
OhbGXUjJ+cixfpfmAX3R8Km/VByLDgkdzlOqTtfwBEHlhb+zdSswJtfrYZLw+tcs
s8V2Pr88VfZ6wqzF23rvnOOWxcL1e4dy9NxkhWd5DNaXtJ71cDAxynLAyc3lYjc0
c00jLfsqdiRXIgqdtnEP0eresG1F9auTgDE7pqZR++mTjf9Xv7z1SfwjpsksrUUS
`protect END_PROTECTED
