`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocfU2e6VIJ4kNTvO8iARpRDlcGpafYdKBTOdLJlVirgCV2G7hCt4UTKLksjeBE07
Ct5ro7b22d8UBM1xIStYIc/D0Dl2FWQ8RwP5rqWPm+xNjNf24fjyzSCb7w3Pxix7
OnmENYVI2nNZULuslWlBV994SW0TgzD2yA6Tl11uLafUUy3GRe6ZmgdIeic8tzCt
1QXv7GhpjuwiO74AU3EWMLgCU9VW9h2/ivsscTw/luUCZObtz9zJSYrlpCB5xWGI
O3LmEoyS+zchG0bP0/4DO5CxiPB98GduKvz3EFKsVoK9Lh8/k+10x+lIEM/92xvD
1Mg9nAnXss0qWcjwsfekr2jTOzm/HvlzY88lbUxzjvK3tnhdXVmIXowpQE5HhoeX
U1BnUc/zgUB4HjNRZtli+ZjdKk0x6HiCoQ8FnZZ+mQY9/dU/NVupkPCN03ZXRuQq
bgdL/qQ5+dlhtjLpmGvLAwkHLbyXNpi0NuJqQkPPfWf+6sFrDCSgf9VFGK61/zuN
UBsh8gubwN7QPsxDeGfxAZ78PBEMppC0SjhQvRWNOTdV5h5PBClwiskHAeqhS1zv
EpkN3HbfAANxCpJ0bXw5t19TNptWbIHzf/SJkFiQDTlPtKqHSZSxMWXuUmeC83f6
Fy3l55ysfct35hMRspyldsLclkI1kfdqEYrk+rWxkUsbNlsk09mPYGJ8dajNdJ4u
F+yWrsGtykRtCfnO10D5gf8ycVPTpLctJScMuTcVSKl4X/r6DpIPq8o/yXVpOII1
wc9cv8EAu77rwuhbcVITTSwJW3XrtMpfxApe7vPF9EFNRH6FODEpD31N4PSTbVy0
jb840GEc25bShV5b32mI6kg2QYDOM+SYpmIes5Qt7AwlF1mHbmziRJFevS3olA+F
O44wdNcX0FuHiYDsn7Pb60x1PwjPb4RTpd+8E48kFunRvly6ktEXqQORc9pPvUsM
DpjF90Yo7WuydB/+jksW+Sh+HvH4S4QF3+oQI9V8k969i6JWOWliKbt3ap4/GIFs
YNEw84ENQQ2spDiJG8JUKEyEBHF5hhT8KPespK1Z+iup7BS+SLkAnU4KtpTQjw7c
b1kRhY7EckiFFCmlqNEGDcVOCPQpn0nj+Yc8O8ztraM4cHUoZ9daxXVv2FJ3XXAj
CUtSlkV4SMydR7lI+wLWiaIjV3FLRrTEXyxEM24/48QQ+w4D7n2bfqnsyiCLfJHC
zvsAv/3q2A12nliJnRBng0IGPcccme742abVBouk/c6l1J3jdMeCLKEIBeK1UN6R
24PWnXmJWL3qUqnIwwpLhxFfFzjWBRdtdCfyMZq1qPl6+nyks5AA0piw3Tk+yJjy
`protect END_PROTECTED
