`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpIsa9CI266s5o1GQntBbLJizYWN+dFpByhCD0nwu7DZF9gnLty1adIIg5lwL+CT
hxLWRF2+seICAZGjY6K5P/VWZ9yDEVEOk1Wclq+fkWh1EVAm64FK3o67i4li4FH0
f/e0ulY4YZQulRtD14KAUyBj3yryUP++xMZ9hoXTpqqxJnNypMlNph5moLx8+Het
CHx8FCW6lUpBo1FOiIIcEEjcp7CMzWPgLDZB7FzIJLXnJ1cAIg2VadX5ZN2GxknL
1JXwuxqULCyO8psdELccC31zST+ku8r2mTycDUQwlYhhA1ZngTs1muADGcVgv/wI
KZNl4xFj/hDxDXwIiip34QtTkXQUiJ+z5TC2sD/RyGeORp6hHNJVIdQskSp1OvUZ
yciclo42zWLxkWXfUhC5awIU91WL7CwvYf5eOoayqWL4tPgaA97UtQZT4/UFmyET
CNYan/WuPIM2e2F80l8wCViks5V0j1kU7be/AksjWBC5oBEdJKLsm8YhG4oWxZBn
wiCx+Ejzf0CHIzbItrngUbvhZ7GK5GYvswEuMS2M2KrNvni2TtWGgGyvE9FPVWIp
lIwEFr8dY0PwtAW9qc4cC1KRrRs0FaMACrI6S03AFioT4COTj/5bwU+PWHulozMw
FOu6yf0a59o/kPSLX+uZkw==
`protect END_PROTECTED
