`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7OGxWRjCpDb4LmdrmIOe0EoBLHiBR+pwVmtidWoAZOZkLhjiTh4UsX56tornyT5
3pkVjEQi6VB6k4xHDf9/QY4h3CO1i+U4wcRvwoXpnioM15BmxjVS2OjgNrfc5zea
1x5h7K4D+75HGetih37j2XDxWPlne3/hwwfkvvLpkfGDeoqT/rlIDDV6awEUgc5F
VV27/JXK8GxAEMnZBuDKfNYI3fVszOSO9Mv8yG74pHWVxJCsy1/62GqAnzntyb8A
hreHWz9g/PyhylUP/1Gy3++oi/dC/DG1lWYe/TIdiLdiUOyr+kP0DLxyjvoMW7mL
kuKlJRR966dB3Dl4uMo22wHKW7D++t2L4HSxvTyn9tVrov7rZ+s/PfWmqPJkySYn
DABgExMTvYGIeex/585YPYWnh9fgJCYXaqmbyeu977Jyz65XdmNggWOKqLN5AhTq
1xflyoSf7yIEGD7ovbLDw2Y6YP1MYoU+i9gvgImk+4lAXgEPFWBxmJsfB987TGHu
K6CDSBckIWquWSsAHRXGCRoaG0WCNQSJxn6reqMkdnbCezy9UoIqVz7I8GD05Pih
`protect END_PROTECTED
