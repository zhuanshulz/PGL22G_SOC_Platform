`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RfVRnKsXh7YK0o1GFE/K0eZsJ8gGEjNRdY1HLOG/rWD2RRo4Opnr066PIONJ3yG5
tVnQahqtjZ1R+2bJLRckZQgMizDcbhQIcxd0KPhbD7qkqNYzdfDMgPFJhT5xj+Nt
9nkvKPR4+8aZbVDhLOEytiv71PjFZWCMqGiqL03YwbSGt1F7s+q+pJL9vywqbJ/2
JzmXXLCDmMqOSS/FqFTPdDV8756P9OWbiAaXtABG1syQNoKNJDlLVfCDDMzyLWTP
Dl4yC4nBWUgqr+O/eBcqo/GWmOS4ONykQmVY5zNpphQ0LXuvTFKJi8V5aBbHjkYb
uCNOL0A3XtKM8WTA78KpLKBy/j+Qnp+9PPhiW/Vhd+JjQdCw+LPmRh4j1ccIo2R1
R/oFJsACb7bHg6OUPw1q6XMPPZJ3nMxuSPSBnpT0aXR/HfXeqNNwDtm4P3b490KO
1sOwEYy12g6NiXsyaxSTi7FpESeyqutAG6/tR93d/wqxz7GNNy8ZJBs/SB8tFhVK
OENvR/p1fzeg728vDTtdLU/y2f7Al7WxADyPZlhXivyMPMcHHsUYsczFY2NTmJN6
lIPmNqrDtoGkvu1dQQdggz8+psGKyMAuTXC9A777TwsRSPWfHpEXJo/YcCO+24Cw
6Byi01sJi4wI3T9Pc6VxMzbtklCq2bOJLTF1byD8RgMiieKVOZ6P3PTfzYeGd8n6
t49+P1ZAwvTdk4vpCfuO3N/o+DVxUBd2Z/SNd/Ba1C2pnm8unxbAA6Sys1BF1oGT
l2sYJj4oA3ycaU2JJHR1HCO3DFQYLSfsizYDSJ62zj81UKx0wg8YqASA6REPRL0w
/l8nwz7BcXyQv2SvZPAtv6joa5IbBFchHStKiH6KX15MmTBstjaLfx6jzS2Y0aPh
L1AfkgN/h3tbt+WnIznfiL1G6EGRKl9MEnyUyLt18uApswgofNgK62UlNtU9B+On
F2kSdajHpOjvQ5nKHNLOXDV7/40dzXAxR1b7uQJvwJowP8KxSWKwhnxkX11husN1
MnyWUk5YN2/ZKdU65bpotIF6NEG95ydE6zQKSQ6O77keNKnDxevtG7515OBwOJnA
ZwwdSPzZ+noEYjrKWTyUP58pRrYubCAKBsObnO/uZxMMo6ye/4heK5yrLxa72eM7
5HvYmrAyLeGPFUXOXYHsxYZ06P1x+QKPn6PftC41tUY=
`protect END_PROTECTED
