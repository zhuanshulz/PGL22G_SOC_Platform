`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mcqrDkphf7W0VsrMFAQm+2DJiPzmew/Wi4fEpmiRzfLWBXkkWl6nU2m2syyDTAwu
SVRt9l1QyqVSPymT8l7t7I6LcE1irFmFewJsKSUj/92Cj0Fyc/Mk6KafnHECtAjS
S9K5R3XfxOZRttsq7d98SvZoK/Pmm7rDbOb9hHoJvEbBFYWFtm2xQmgoFRykCzsw
FClt8XhrsepcDaA2PB4CLVINuOeRn2dL35EXVyy6416d8KYzEjzPE+RHHXoqoDsT
IHjVx+3ZnGU9rRj4lbUURwIl08G8TJxMSQOHsNPIJNVmBLRSy0Mrj7XWR7t9kCEX
kvN2+ZIImavNSRCTo+ZuaU3EtYsP7zfG5Of+jZkXZUwLJMR0lxiMyGS/9sK4/y5L
zmQmaI9/nNjdgvyiKHwzehQHvbKKk7qvfJZkalYTJ2biPwcdzaI8SMfxwhfagWF6
+Qp9JwOk9iWqMPuLmfQCrki8KkN4cT8vjB56cjudeGyd8dAn7AyzuSgrJOPDCBPo
hU43t6rh+blfTdv9PxyV41r3jD2R3IV3/HIh2HPkR7sa89cJvq4Sfov09rkTo/ma
Pcgz3/6bLxO4/sYoektaZgqeP72gWYCalyDFop15PAITsy9LSWH6qRHObQtkER5/
KDlFZoalyo+dMmFZSFA8Ugro1DJsPT1ZiXWJQfC+OkEyGRV4Ld41EE4OVd0lrX61
NabeCwVHrJnoLTmuZxt8Z2ZJvll6v58cMexsb0YZoCeJ9Ke98UVi3xAssok6Ik8m
f3RGldq2f+etfbZaxJu1pE/Z30hQcrYGqHAwawttsyl8PeIB+CdgfHO1HaXdWT6W
eGujZZF+NbcaDAcJYdAOEDqecQRHY+1E+4OqjEBDJsIQdI01jwe1rt+m9XEJ8XQ3
Utjj8ti17xmrsdSIQ6LWjl1mQ/cPH3SiDnwqyoAe42JFDsruyY+XoyCZbvcVc93L
kRUpJPKC3c8X3hXupjSzfWZ4CbJ7b9chCozGodW6BrPPfRwzHNGLJh+9lNzsl3Z9
760E5BegHBOMRGPv4uGgEI7eDpad75FDEdb7RwlGdlIyrvEJc5gY03XdNF7H/Vda
rj8xS9Emkg/HfRG7zBfy0Gkcth8Uzzy0WdpRbYdtCdl16Ma4Mns4X6GY47PYxWLP
oLxvZTYSzhm2S06sF8MBS4kgmbLSZXCuF2m3FANmNRWxjFOWwHfHONscYrFOy83f
c1OhN42YndBztygdha2O4JfJfpbZJ1DWnVZBw+QqC6YSCIVbWgGDE4QyFrsf2YW1
w62emt/4fjGCROPzk5ztoeQfutLFqDlfENaWBTVKpb9czld7yipMu/xxGONfFlrr
wwLzKV3Cdb1YXpDsTbdZQKk4/HWtan9iUMhZOMCy1WzpwSEXr3K21gwKtXV1IMmX
sPdCW/Olctd+7grx18QTdWFFBULSwiecH3lgO8YpKFFXBLahN4ylJiWGyUzIfSXc
0p/yhZzhoqaQfb6J4TiMlOMSdNfbXwdq63BtORiWqEavZoFAjpEHAJFQanJqhUm1
JHvGwa3fCPo/pzGYc2Gb/HCHnSHYpnHJVB1XLZbh3YE64NVyGL+EKGCUUOua5VTt
JNY2k8Vzrj0LqcbU3/AWF//0lAKGSx7nW/uY7dhhsnOL12Cakhul5l1s0JTwpnmD
igwZvubdmM73VSiELVL/zIBMm+OH2FVZgKQzALFD55ZTnlic0o9Y1slLsXVGhBGw
ud7vvGWC8Tbquqq+hmXGZzG0i3o7gkRmvrHeIAy3Q33vMENUHTB3i5V/WAOBs69P
l9LSrLxiRwN4b5jSHnk4miN7TrSDo+1qiSI5Eh9whp94dssF8ONIwz1CixJPK9+f
ptNIwXthFU9ay5FIbGWNqFiNGrLWml/fSJjQgElRZVDmngQLYHpo5WX8qCjha5zU
THRe2DRpRHJNRPyCRryBWjp9cYtR7LU+N960Hiuzic/u37c81WEuUnb5571WsZ6V
Oa1UiouCFG0GgqMJRZm9bUWoJnSXZW1/d0jC/oR5R3XDewl4jLLaT/FNEy4hqBxP
qQkLToX+JrUJ4QWL0a5ibAHjGcEcP3d6k3D7l6GWMHOcLVRoQqsCmniJXTUn1wNi
GYLj31YN6A8gPLexMvD9k52d7vIX5KHmtcRROHokVOLB64JHwNiO8vmeYgGJWjVC
w0mdyBJ4z8pY1nvZDk1GYpGi3aPyusFsE7WxsKWn03BvwCPJqbpN5BxfYZmmgBUy
yYFGwhqmQ1IVcpta9hviDGJmwtquE2ClG4x5fp9/nTONzL4rK6wzziuYX2wRQAaT
yASpLIANIM85oJLS5p1o4YdYIitaEcNpFUocBJGufbyqTkFkJNSxgaay0uEtRVyQ
6K/xA14hdscX+BRHYzzrXg34TQ1AjynrYE6HNdVNduV8AF4rJMOrGQ49fkGfW13y
/he0ia55LvvCfnvL6Fz9eHLIEgDIc6mQSX+Osqche0glDKDCl9/5uAAvdHcIyCIi
/T2cXU1JG1t8Ih98tJD/ggDUyL+sKPISfrzVaddxzNqXa33HhQiVIEL6MFFPzAnq
tk7SYjUs5UxoV1mLyRbwMne3CLe3UKpnztuZidPhKh0NtVZdYqf/QdGgAuXSFWoZ
EjkXSy8BzziWN2KiL8cb95pU09kd+ZooCEP2uL/r6tNRUqPRQ3UbC7mEyjn0ILDT
oCPw+WISCTXlPs/ApElEGcRqYuHxbmih3VQCGtMSAWPOb49ARZDcQ1eFWS2BavfN
V/J/LvqwOrCoba5V6Lx0JnGlpW6T75QOLETlfKdoTuNpiWj1/VVOjvsVgkH3r+wT
TxlRfpzoB17wogP+qJoO1C3XRNBi25iyFpln5WJi0hxV82ZEPbXf/A58y2NjXh7H
AniB0p/Q7Q8zVkUr/SSjpI3Vx4DZF4kNIhPuAUKhqu+zOb1468LfOZjFuOwaAzNs
KDQKT1pKIdY47Mep68ywh62BBJJt/j4i6u4Dy02P7Cvj+jowuZLmxJteCiBc8itH
HinJp3wnRETHnXw5PLvgIQwkkgdNBgrgk96TNtS+ekSpUy6+rfIfTlr/3hDSV80s
yHJUueKaDY7z3gdhlwwRzYGOGUAbULPq7YP8w+TmF2AZ+GpqZHBpyfHc0+cx8biQ
RA1b05up3fOGWdIRQ5ozhrrfHbDLFMPO0osQR60wuzUAMycxeLYHXsYO5+DLJ0aw
lDkPU4Cd8O+o5kRXgtsL+T3+MROGy4eF6HL5O24UFxZdxD9baiYYdBSp+Mh3R70V
QcFSBcGocqUPCk8tJc1b5liKPy9AqEG9aXFOo41zNTnAm4b+WylI3k5gKJBVFSHz
NMYkJ5x514SiOkiiPwrqcvnEguASorSiXGhJvl86aEzIXt0PjzrRFnvrDV8IQcq2
Hm8dgYpGXZCWr5F68dfRfQxMMs8TUv+9Jc1BkIsmZqRJxkIu/qesa7NcViy7jvW6
n9DjzinST1o7OKyKXFcAb0WMwoqxwBgbRtbFfXSlKpNIj7jM6YIAte28myZLWesb
0GXnqJVRP2tuL/e7vPP4JtP+Yd2ehtp8dsBrxeGu/pM+KrZWjvdNpDnZZt9rzshl
12AKVmg2pj/oVCkEuLPB6K8LbhEajZpsK5Y92LozbwJHl5EJQRyI8cuMeHHYbyG9
hixGaJUBvKJyYQgkNyWS7UjYKawveIePx+W+mLwb7LpsPMndXsWI9J7SafevMMmB
RMkRmtOQD7SVkxudHcfgR2OK/ZEVePWL+2tz3nGkC337C7KDyOYXBn0bUGP4QW4F
QaZKHCMl7RR3lM1QSJMyF7SdksBRPtyY+Kjin2/t37F19HwIOTgiHlANNe13fqax
UfvEUfjG16c1t+B7RvT0/VXwHra2Zveh5+CztjxHEFoOB1U2ChwU46a1MgonBg/0
sQRuEjviBNKhfdC782YBGBnGGWNxcU6FO5Lu++mtXfxh44LFgXd75iHRvK3FZqyP
tojtQG099MG4jJgFpiilF48Jyf5Jsx4WK+ifYTX0qUCbV7b6dkgqxpIivoWB+hzQ
Oj1wX2ORzp4AsILcXrKLr/OuW0/mMKYQlLLVwMGcIz5ssBqPTCWY6hEuPQDUKdgC
m0pWkNt3Sjh4V/XJAW41Nij/0xTd5TJwa+Xwt580BAjD/6TTzwGx7SZAJYRtD9dk
kwr9cHdQ2JFtZrbNvxNanlSga4vnVQiuRXVDrDaEAdBB0oRhkoeRT+4Iz+ZVi+ct
6YwzZWixckooyd5sfVem7EolIuXOwaJWGNzBajZf7bpWVRNIcOLUbSO7Z3rIaWiN
FCo1Bo74ES7Bpa8aPGJXZsJ9hO28fpFG3/YJa5WnEr1qy8MguPlD8zPz38T+20Cb
2UucMU0HbAsUFDyBI2O3orSYbjc6S+I1ISzH0TFtqbm1CKL/Z0iJLFjwuqYIuvkF
PGlk8xLUa7IhuVXn8EKt+mtm7kpHFcicnVJ9fHADEgmycnWXf2KYDtdeWdQ1Ifg8
Rqv+iaO+p9XMlbOeDJLWhrCZpxBbxCRdIlfYGo+npD3Zw1G7g7kS11KTEO4J8fo5
H30Go71n25UjjdZUPq9ijKdFBRvnNFikIDBeMXgIkU4=
`protect END_PROTECTED
