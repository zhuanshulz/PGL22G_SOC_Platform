`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WYwigupV+WUK4OA/YjYqu65Iee6t6vQ1sj3NYe2Z/YVRv/iGrM2g58XsFow5GObT
M+GlaL71qY2quGMxHWa+sBEypV8Dgs4IZZlx9tkFkQS7BzVQmmMjjGgduR7k31l2
TUjsQycSNKco4vcfYPyOWbXBzeK2aGxRMGdaevawCgQMdqUK8ZeKW/6GVmAjBeOG
w2eXIRgT1Z9GWDFVJ7HTzBwNn/cjoecd8m1N8v6cdjs60kt+pE+T+yzDvA18xKay
sjNj0kfMy4xhgDqPlX9jjyDR9AlM+9p/dTuP83Uj2DINmDv7RpCRusNhvoCwBzSH
qXDsC/40Z45FIluELBTXoEmNNByR66d1iF6gxNBhQLvhUV1UBgDzneNbVp0Ex0J6
XimfgmzKhVuqapORWopZ/wDn5DdRbPYl5hPmj0cc/VDXg9n4RbIUo98Ezg0OipG8
PZsxmVFcsczikQaldTtSoameGoY2WK3iXlRxA+ii/i2lZbluZ+W18mDjCvtIbjkz
n2VBen3iZNMmJxe2mRqkvD8mVfvOfmHu0SvduPbcRTsGb51gdiy981kOLgGcpqpQ
wRjz+614PSxqlANL02lRElubID5I6q9bKa4DxDDAmk9AC0RUW0G/OWOZ3xOPHlm7
Wn+/Dog9A8tDKKt9C2X9gnKzi/kCJwUlR2vt19RqI85lvpyLF+dVNTeBAQnmXMm6
994QXOx7aVnjzlBeO+LsaBubdgp4h9lFGuaf2Yv0SME9a93GK37BYAUEIGeGaomZ
G4qu5p6jiRQwWwcwp1Lrbp6HENHnco5jM+nWORIXPJW57YnSyyXAnLFh9UZB79OT
QImoY2+UETxsQuKwn554oUU95qX5dsE688o7crGLrFJbX2eRRhKXuPskjWfM9VUq
/k3RmnzzkP8cMzgomzwjgcILoEFdY87fxFLAqj1JRx8otGubg2wqIioFee5WfyDL
+YnG+5b/gJj0dZZXXoOTgd321aMFZAZDKF6RYYCtaiwvHUpo0uayRycDOPL/4dFG
0H8xSbmOLxH8H5oFH0eNmJfVZ7D6CrvCpoD2NCcME7A=
`protect END_PROTECTED
