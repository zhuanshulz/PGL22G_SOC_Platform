`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDAwEHYfL3E62SPqFs1DGdzzWYwWXx2yWs6Fvh9zu7+w+yluf0uivali8s7wfD0p
B+2YBakhD/cKMlwPGvBACq+eEN2Ew2WBkoBCVAs22+uM02nTGED1v/88c/iYmxfB
gd/bfAyVkDbzY6oYorseVS3+gZZGvmk4yyZzGGC2dzCa94onri/3LnrNTLhaQ4Wq
S1QIL3G5FZ+mBqWgGSy6AaDTGV0L8yLAicFhdvI62Lvwm0HjOjPSL2mXM3BTzW05
K0K/yqNiNMvEaD/ZdBQ3TYk+tjV+Gh1GjW9Y7fJiqI/zSmqc7IGwMrhsKsOWEM0g
dCc8L2rSeRGxQy8v9KY8yEPcr0pQ813JDlk0vplITD4galRbx73XvNz4sLS4U3D9
2wg79gAaL5XJh/GSH4ntwGr69m7LQYrCX+woCxlY69m/KPDlZ08MqxkLsSTrCCtI
459qZnn4fa5oMLW2YETRZXLqlQtoHy03X4cKiPpn59RrFxe1Nz7MSng3jCs4S7Gk
4O8v1GBuQm1PdkZD/1tnSCbFSZa/Qm8QX7AET3rOz23DCl8StSWATZVQuWe88O1d
09+23oSXxcj+jdkW8T06Rw7neaIansjTDg/GJKqW5Q3ByIa/WIuLoHihQaDBBAQo
Ue7ammVwtb1k3kADJklPkeG3iegQyQxsOUxwX1ow2T692qgFV02iwc3XS40/whu7
7XfqLAAEbRvr/pnDZyOh8Z13WsuPIjPt9hl+QRMNtOsS1i3yoCm/MjSlYUIyRZ/S
Ki5rShF+wskLkRT3wEO/IVroXTkoL5fv2C1s5QB0vAJYD97Oh+ujf1ps1Z41/UPu
C+5jT6joF5IjCO+Og2Mhi8aAAAY8oTV8x9oXdH3WKxf0zLu/EBfTzJZ2BSd8Z1XK
qNJWs6zh3lrU4jvGjPbjKKMcqBtxwYvyGFtdUFz1IuRtUGeWdba1BoPcmVpf8mWj
BdvufXTun+Gl/H5Q3qz/OlKY+hIajkpVu7N5Khs8XDjh6p4kb1nI97Awp8juukSG
C/nwKQf0rH2iwSdn9rUgdP9t+jN1CQZKC2Z/Xa9ghzHi1NimDefRlPsxVHove2M5
8w5bDQO+2YGUtmYE/PpKxT+mjTUih20BIg1veMAztswqxcSy+723+y+X76Y0TuXF
qGXIf4VpoY34X0NVOUOFa79d1LXRJtV2xIodwbTBZgURQLvTAIdVNmyL92L1pko3
GNdxvM2wLtrMh2x59psm1z6iDM2f2iF6zPU2ZZ8F/qtygq8+f6wdjXoqxh4I9lOb
giatWVssi4dZs/xUUKZLtglN/Ygn+T95+Nh9LINtespCDEKj9yEwqgR20W5ypK3M
prQsYScCntM6vDcRhiIfAYNmAF+q2emvD0mBXOzROMAs+1xS6L4DIq3bdJ1BgWv8
u1Hvh801u9GrTKml9L52yAr7RzsKJVN4fGu+FFV/Q9POrrRTTM/0eYAkMMh/bJRd
I/lE4cnaN6rMEY4MxH2Qtb+hKq6dh1oITQs/Npc8e4xBfnGSZgL3CBKdlgDVCkUX
gtHrhp8uQa2nS7EEiYNgAXyoi8wDtlmT7FG0shG8rCfk8I0UJuhZViLSOLMEVAEq
zA3dIkWyno4uiVBGb+bMzpsQHS9BVh1X5ynvYrzCy4OXd7EBlb9SOW54652zb2ew
JeP0844ETsViQ1exltmVZ5fvqLLjpdlroNGxJSna+VK8EW9ICTAGNoitfPaaTpzs
vllgJ0JIXldcMuM1ZQL5SXlCujET5zexaQHsi+Ub/DfX91ng92VRToJDZCA1r7QV
ah4t23zRxLbX2fvL8r1jvOnMxf0FXT9n8omTR+wnpzkVpVOtxA7yhMTN3+aICfUy
d7U9r7TunImV7yfhkCe2Q9GMA5kuJuuFcfw9tIMEfg8cCxsB28gxboB7/9O1gedb
/uyU2wMjspJtvAnkn5sw0DaOq4CFHuOKHp+MTFUW91PN4TEOXkIJ5p/TWHnedoOY
PJH8PLOlOhCdCoAO15JbeY+OdMSYFOub86ReTH6bWCRdF3S+MvlsXTbQnc9OW72V
39Vk01DN0QLUaecVWAMRWNXECWAHDU/1TD8HFYqflr4xkuIfWEVPlhjodfNLI6Zi
kqNJKLJYhI+sO8ApJySp37tf3aEqkYlpX2Q5JhBMF19PkL45uFPzb9Knqv7KSAL/
ak02HTag96vuDmIRmzU8omomDdo3xQoYgkamBvosRDrj9UW+13A7ZtxZbywISu03
uV0BJJssRJJBnYBjvVI6ISzV8xWUbr5oHNT57mA4CQFS2IGXBuc2ZYS04jSh8THW
qeNByGqa/nM7MRyVLPcsghZ5n5PmN25+5I3EffjATLOe2uii5nw0ntnbG8lO4dsY
jynS3BtePV1hHdqfWL28preuYgdnUnESfNMBJn5pHlyB1oXI0d/05rwGg/xto4Fk
xuM1joCS1YY+t3P3bQI2Q1WqaswlA+QPjD6PWIz98Qz62xI7Iig9YzZFuwex1R4x
2AaPboLnQHqQsE52yYT7drc5O0MC5chiOf4XGD5tISq5TUbLPoQRy9/ik4Ea4faQ
ZONgH7isYv9LlErQxSWYZ69KsQK6acyh1oNvDRvHSwWkwjJ7bjnFctU7erjwIHnp
rN9zS54s17S4JUymj3mXrH+invJ1TzqdQQGbdvW67kpDNBBOVlBvTBkjBJ+p99XG
0eIJUlya2ULgQEmCqXMNVKs5SDHhaKekL7NbpsDzce01uOS5gHKVKaeUKoORgy0S
3hcpatXhADKdcHye5gYB2E1f0kyxdcXxioTMhKNhil0p0QsWV3KTwvBuI/Sbf2FL
R2aIle98aKfJCK6qK9NjGd+D3XT4YUGU+VcsgU2/7nXly3zFu4cy3BXmP+quHWWt
feOJL5fIY5P7HsyPxC+9Y+xyav0wntszkFvh7yBZvRi9oHMCFRuRqXmvB3F6GbEz
LQNIb6kk7uBl1OOfzAzkl9J51SmbIlcKVUzbxgJJHHHhNnMi8VoMuHIWYjyoIMS+
xhNV2nQjikxrZdc0qfVlI2Uk38Um5l4ulfW20uhzTH4k5viUuq59X2NFI00/GEj7
943ZmGQpHb7LUaROelajiroad4xWbkwLdN5PuaLxp2uaO08m7IP3KeCxSYePL/Dv
tv62Ouz6mxmuf8etQlRJ75KXcoHhDc4uUrv3GWgnmJ7B0FvwOqsK4Bh/+CdmavG7
iVegkdIQbFN9FxxgHgdZvSGv2RO06JHgRPo64ZP7LyA2zLNDdkDR2YfqGhw8Yx3A
d22osN5fCDFWAzgT2YQgSQziWsOiLFxivGl1uVFIr0KT9fNvZDSbRvVBKBJYSjaJ
gSTVGWXNUB9Bx+Jw2urHP6JwSK9pPOUid17hkGF4O75dAXNM87Eh4cRJcP9bzsHb
SMvW48eljjhvxpcQ2SAzynJC5Q2Z3aPJDhytvJRejDWdqMm4dk+mCgl1sN0b3maP
29+GLhxXYSkxOf0cIT+MHuonj++Cc8TxcDJQaDZJAEceQLkcjwJA7ukXrHBFFrzG
Rzy0VLYh7nc/o7+5wkQW/jp22N/md/NqUoXQRpq2gRBvs8gGbXwUZG1KNYnOJFLH
dmD7ydUSMXALdysIFlu/uo5ezQmaSH6u4ZfbBnKVU91APCnpJWPwUYWYS+S3ix+/
aRZwOPnmqAtPpDatNIeDZOzINmQXuUShzQ3wTWbJkwahowQzkwT+6XXwaUVZHNc5
OdpDhbIRKbDyb1a8AjbPpw8ifspk/O52e/jDrklsv0uTFkstSMQ/lgZt2argtfy5
T5Wl3twzC3hgEXoBuuHFuakKCG67fsrF/Vn33OUaOfZ9SAMqSX2DHqUnWlKqhp8f
00FOV9MR8uhB9aXGPa/30k1Zk7aDockXuMPU4xpK9NjOXr+N24Fcr9AE7Qel+E+e
iiIk34RDTvqdV4s3gOVFRQEj8MrUw244nC/jpLXZrFTgfZzNL3pdKgnm3E2rTNuX
YOJHPM2TMBVoHykeQhKP4Xs2gBZYJ1R+yOVmDJPfyfaKISjg13oRIcvHvmOgTl0U
23wBPV/+tcNCZNMv5NKebQ8LhtKzZsaq2dW6mOErERl7rosADQ8kUsg7pirJOSIs
N3zeJuL/iWav76PDOyEfiJS/6bB/A2EwBTbmJDFh+5lq2rJuyIAfcwLMzxDLz47l
KRoKzz6KE47SSyZ/B72cpu2e2kLEL4qxILS0GmhN377q5bz18F0MmuIJaARb5z7w
w5kv1H7CQw17Dq2uoahajQv/6G72FM9Va2uR2MhIy76z5LnDT5lr6ssKxLPCy7zE
gJ0Qn2SrF0ldKK0gfwVuEf52IR7Ry20yaNtzTKMM3O3/HVAnkbLOmAyg7wlIDFd7
/g1myqe4SxrZcbanSlQ8snc6ORD1B/tSCbeVRa/U6TuqD+KUboxilrcqfYmZHMZf
q060w+5yN5Mk0XuhARL/DA4YzbAUcq87Km/hN4LPVCvhkXRNtai+detAslzMdj6b
ewy3/cL55eA46RJ/Ghaosjs1uDv1W0nXY2NfPj3ymT0PDfQP8cvn38y0zgQrH9uy
t6DOQVaQ6Zcb4/Fd1qYrPsrahRSU2tGyzgMKXwsXTX6Qk1R1hE9At/n68EZ7oTAP
U9De6QsdsO3U5SM6ylntmd5GGK3AluVeUHp52dfV0ooxbW9aghlKC+eNFxNTxM78
HADIT+3saBpyj6iXILnoRyOxRhoNiDoYmriBjRh9kVasKEeU/AXthcAP5+uI8njA
rObQiAxq23KLWl9aVPsq0sTWiEiIyjrA46rRzzh59SP58lSt1IfG78GOp98qhSo/
fCK1A2HcUPuwZmMwymZ3X5/o+0htVPAnlknKiB8v3Z1M+rCfjntaXiqzTQr0E58q
taeB1iSUCim63zP95oHX3SNb4LJOaychUkoKWAxFralXWCmJAEFToPJXiQZfTttB
3b/sASpvcXSHF+lxMSm5FpNqI/JHOkqXmhO7EQByRwFEjheuX/xfMGy2jKEKqzit
FlCjE4x6vjWUmL+wj05X91c9+oIalN0OnsAiH8IkJz7vISDpg6T4bNe2UAaea1kg
vFobvayQcbFbUH7+3jIz845kYoASLVMzJjH7yYmDsAshFj5z8oXNNVqcN98po1Vr
JWEI9OIKM84CAKSNqDXRXumgE5A3pX4bwU8t+wD2lxg4aTC+tqVJ04ro28YnLjt9
27PCv2CWYP5NXbUpp3ysjNElmWsk4b74WHLfCyTT3W9mh8aGHzjAcNKHNWJrP5CF
c4PxQ1RuVSFq6WWgwfH2hIlhZhfPrkAvXORYhqfotqVBX9F8OtiShz7ObvakgHyD
mviFkiS6UfXBSOiB5U++OYzz8dpZl4TaoqlPGgxaWA3Nh8bm7/j0GapFVd7Y3vLm
cGesHgpHKNG+BU49dmGJcpKRfKO6dYJetAuQY/WmBpSl/xWSOYea16sLvfVM1mxS
cCgYZMxHXuJXgPPx7Ila/faSfV4PNF1w30Zq6eRgsL6a6ydjTe1F7S9KaCjyhE7V
ZR+x+Aizo6R9QWL5jFek3y+ZwzZBCqTTVJ0sd8sZ5MD8x8g0/6hwRm4xuu0QJn1j
LIWiIawkXUfCedPuQocivwzxO7MAOqgwtEL+A2Hyy0lvf+zspkYe5hWrHHThPGJ4
DSj3dsUpPvDq/p/iWvICUn0opC1++AmTvmgmV2sr/xW/oZgV2YQA9sTMyKjAJRUc
bxnM/z32410zKolQIsv5eLgL7ZQEemvtdWXbi+AbgKfOV5Zlpx45ywpbEFRqFvYp
BjqOdPDyMvVLVijP0/zvDPE6m/Yy2/NPkwS/gIMPYZNuePfBdtTDCjfz9DaBDa3D
vgyw0dTva20HU3DPnph0m7J04oxfd2TD70YwLlaNkgt59BZgnBEHFVkLheIntY1o
WqjQmZP5aOpy4XIJZQ8jpEdDw4Z8v0MLTpPJ5kZWqtX+l1xsHxfEX0Mzyq+tSa/o
mjQbNIzzzn0UnI21CxT7hNpfpVIwEbdwLoxsqTgAdGo6KMlunhn1YQBZIF8CMBlU
x1jT4ZGFz/wroRNyEE3SIpeina08DH3JzV4A0RN0z2WTm6I09Et7OID/iEPI8nbU
/gVbPwJEPJv6LvB8OJRobOj09iptZ7PW/zClsQuBWRu0sGkhXM/82lqFqWF9gzd7
KAMdTVj4VV9+RJ/Cx3z0toWheZ/9tmUPkuvF0k+2fSH+hlO3aXaH6Jum+X0sw9Zc
bKJp+GKlO8nrqyEMspAkEHdA/wHypHJphj/T5GfUHw4gHArxIjla9cWvsi/EnKcz
AHkjCkOkkwamBRGBgj3rYNbdxqk3Tec2fcHEzHTRkG5VeJ2sGZLDE74O2lp3gf0/
WSInYaTGPUR+nJflGqvn5zgsSRjFfQ5J3fciITMuvW3mSsBhF6vjiIO/Ep78cn8A
gpCQ6oEGN/GbTDHwLW4fuAxSADno877QIEK1Z17Aj7juqIUoSJrHo0a1rr2z+OGE
4ePatotXeNFc7pQo4EPYe2gLCPU+njuEvSkhEQxavqMmslGojEA5oRQ7hh/aC+be
tp9Tio+aQ5PBeE94mU4vx41HVu9ve0JgiKpxF9VezAaOcZ0eJMShMIRBwNYV267j
5V0IihwWnBZtXQRJno8/3kka8rrL+28QFjbiaNkaeT5XqqBGP8OkdtdIiasmmD74
R2IJuyKLeYaKVr5Rtml8FTqIBMGJPqkfY4C+p/Nvl1/jLgTiyjZf+l2bR8kcq4TT
jn+b2c/todksalyFvoa4qFi498T4dWvuBQQUfmVQqBN6iYyWoqFR6pvOKmbalDin
wr3NNKUyGejzGr/abIxOC71rtHpLGKMHj9yrhk+OgsI7SkrLrTWiUOSOR9WAD1DO
L8bGo4jfc/NRAyloCoG/aSJOn8wRPm6LUBOuf1OSNhxFhNxXGsPaliRSCXF5fci2
8pFujw0bgM1ozh3dzKy+vlnjgzwKKo/0pg2OCgGSVWfHEwINwA7wzAD6vGMx3rgp
wpZHlQCK7gCnh4crhoyvZ1fFigFAkEzBYAce3hO8DwllVsn//YEetKp0WMnyEYhX
7gLoBH2qYKoiDcE1cwG80JdMXYdKZiJaRMAFPYotbqaQtVjMwbKY6pMRa1wN0Cdx
d9eQ4eFiFmYH0UvmVtdSy4uCCrkEXWi0EgWLW969movKi8smsUb3LWYpWw3JjCF2
TeGT6MJOlwExJB5/jZkWWOS53X4Xw0mMcq4XtR96TMiBzI9B45u5e8MvW7PwUW0I
Rws/9NrSRdoyyf21LVJibgwu/wLzcofEV8pJL7tl0HDq/n4S5LmpxAcyLI06bmNy
Hdl3hRPw89iy6MO3ArDY1Iam5hFUujNuX26AlaVygQxt1fJTx5DvF5CGlqCAYRKY
mXNLAO9/44zSvTKss5VF9xnlJ4WGz68DgvWetYBoaWQbfZPXwe4p6BzCuM5q/3V1
R9KuNCRAfDOtBb8/WcIYRwflZSB/Xf5Bw9gnjxO6iorl//8AMN1vl86+sE1/5Ie8
xV6wBNbGSXJ9SpH4a5xXpHBUNj6qwcaWKEJ8CItVnW+ATnOdVXuqSLL7/wAf5//N
7Vsl3pI8ngwFPLTOdVMjJ2lYGE3asFiVx86cXPxh4kas+gPhoBwnZYi1bh6dIRGQ
9SMkuCLvJCa3E1oNu3YD0G17bGlxFqMwERr79SUTJ8xVqUFZG47R/eURUzuUyobL
Asg6Ie0zQyQboyEMAumvkfbevlQ1CsmFFFGO+g6Vukw2aHKPLkj+CCSTL7rF1/xK
rpwFz3S0zrSnQbJSqM/aI/xm/QRNjeFdzrwBG/wnoS0r0M8WW1vWxBDS/sUKQJQK
lO/2dvvvzw76H2/mTTR3/dLLLgpy0HnPzxF6ec0sDhaybwdDfLYEcrIDWi7Qyvek
9U9PMHGJhxjoFq6c3f4ebIwW28+tZflA0M0+F9QUx+X4/2KDnKf2dkhCo6FInrtp
mtw2UdSokL/Mt9n0jNUXxtQPVflXZD3cYlUAhHJxKmI6QdpjWAV8dUFp8xvrLTRZ
yGmQmdS2/nWVJ+pR4Wrc3/jvgqHO1UKgKK0x1HKqgJQ0QyMg0zmUodyZ+PFA1R4c
YzSgee39UKNqk3Z9Kr5JxErOcP258m+hf/+f0r0Gs1gp5kfOKu0RhVuZtNtQZUCT
3ZBYZGpmNrB6uDpxgfXED141y/sJBKYihi/6woWhffwkpdlO5oIf6EeIMLxrYs1s
oufJ/nhXGSOFQ4n6W7q/P+xffwr03GjqCs5lhySw1mApdncAz0FyQfdv54CHERet
XzUa+GJmIJZjEa5t7KqHYqUBP1wECw9SbAqdYaHb/hMJDaaUuWmFqkShe6txzUee
qgnSMmIE7kwHtGFAMhaIQY6LSgRAGtx/fB/nmD6VaoSX+ac8pT41pxVsn3mDx+9t
vq/dBNln7J3wnQd7BkPT6bgsmL4yWdBannGnk2IfYtKlmQG6XaB6tOWftTDGNqlo
wiSw0IYNs3NGeYYuNBuvrqCqKM3CrKWGCs3trop0nn32CqimDN87cP9/HpElxDm5
URHqBG7MYr1j9BL9RyWbJvACBcecNELtSKAppAH4VmzdykPX1IRn3vOkn6ciHbWZ
3ZMawRBhhRk78jVsHhAgmiIcLD7JH0KW1VRvILVxCgF4BRpO6gjweCOZdCGkwXHq
3dz3s0aw765ecajPkPf8J+xCqGVnLHKoIBXGMFRew45lR9wIiTAQSZb01apTPnDI
dURPYQKGLjcBlNwzrE7oo6HYfWtGsGxuxJPS0vhy+ee/B8IBGLcFSy0euCMysD3F
+3BbN9C4HxtW7/FAkrcXi1uUPk8xm6rs9Jfwm1MwKGdRN3H98bWnSnKhzdHGIS7+
YCz3jqQaGkNxYEUdfQjZ8H/GqMlgvYHsynK1zMnb9w9E+TH//Ze4HWyiKKa/EbPL
oryknYPsx3nPjhzI14lJa8KdaNlmVo3bvAXB6QebRFJ4jkE0DlsZIP9uciZUA5ss
dNX3kQb594hhNwy6XGXwMv0NfqyIWq96iJnNcbNY3nKNFxJ1GZ55evfo+DIxqNio
3QYmjPz6XKFNCUL99ko/EX7e6tgbsyp4xqz5x2e3LEGiFaTWcQhVYu2YSuK9FaJj
Z6lvOcS63Kki3Ahe4qAyfb5PLCVOP76yiSnVWjtGzww0t1B8dpnfojFLW33BT7Gn
5ltOqB86RajgCkaSRX1RsOxVctRjNvOa6TLolNke/zkFcVionlQt+L0DrJftvm7x
0Qukt1IDSRfJoTOCHhYE9KusIVE2uTzuDEuxwp7Xpdmrlg/UKBYAxsYvVMVKqWbZ
MKb7a1zmzhEQHnLDiKBukb+UD+AfP8XE/4596uytSldl0eCAbwaojuFhHi7UGlrg
el2dPFxZ5q8ia2e40PzEz73+vGbLKQW8dN+cSM0+7xqpDkcOaTzgV+bS8iCH0wsp
iPaKBjyTSIO5mQ3ybgoS8whmVwLjhuMvcN4noKZsGGMevzLo/z+JA7kMtvFZx/AB
09T1pIWAxJDTX52vl1pGAiP4ULejYRu9kHLdIbUv5XONAjPJrflvMPXPG6ij0PfL
pth3Fc44F+N0dklMt0t4sk6VwA+TSanTMqExIil3x/ilLnZ70o7n8xR8c8UYv2Wl
8svuOCq5Br+o8k1K6eOUS/RlnRXP/0yR+TrEYP0ZjEiUNTfo82Y2G1gqWnwQdqgV
1QLVhMX2xCFR3TdHYB/jub3HBIw2yWFOo0nOEFnemBX4srMijffk4ndI3T77yqLs
q1nG/UVUptYLr9sZFewHG+uEYGwaIxNClIIYt7KH75rhyb/IG13t5zgVdlRKJKyr
JJOTQtS1ks5pYQ33uFaMBegYu3Jky6jtWVb1K5SCuxUncEsygtvO9uw6VIzIi9Uq
OEPTWkogxHsdwWNKwmss0YDyGSGoqNwEaT0j1EGJYZgvf9swBe9WTyMZ1nBzPJj0
85W6/RP88je7lO9/8ok4Dcl1sC81KXLgnvciCxdwr6e4QcsyZvDydbqanKT1WC3E
2S1LrCIGVnaXMf3qUKOW4tJrebMTgr1mrMv8Go3O2Rm1IGbMdL8pDNavfujv9/JN
SQknJKguRUBjxgMlwFUBz3xODHhVD9eWXPNjcrQ1LgbC9GriFGuoU1pHlHuSGWum
0mqbAgdqiW5eQUG+R53ruKI+WkTYmkCO03l6yin+VYrDOCffHb8u/b/s2LBGkf1q
oRrVBl9vEK8JYmmuXTLwErhoOP7dcxz5Iew7Oed3D/XzliITy0acTEmgrTo10gq/
SulMGS72ELyH+Fl/GeBxJ/81D6dGmowOtS+56Ro9Kr+vvmP33/N0x6COEkTCwtJQ
WKC3g1xXNrW8gpsyOJiSxtPXI9NGaVPgXkCU98t0PtuTxRs6ZlWtONxWD8eBopq5
66SUIP8rqhXstOoTsn5cLB2QjB3W11H2agYh81NnELlT9nUdaskOIc2Dop2xd1mG
APrdXeBQMLPYQsKdgf/H3xusUsCZ1p2u7uJ0OMNJip2T7MSjv/pc/hUkGLMKKTyk
Aomv9tkYOR/ng924hpFk+zpfnWf5PaUao0Qun6lGJ6f/o+gG9+U5XzxjKi1WuJiC
DwjkAf9BMUYx7WRhGHb//z9Y9LZEGXrq03GZizOlqdH0nWEkD9h8IHpmHvrzy1nE
T5WuKxsKrB92zJ7+mVUNMlyxFTQyjSeTWanpRT4rjNaNoxVme9W4UeP5eZJWWWjM
KJ0/wlZ1Ptb8t9QAhwSomwu17NeWWSVAi95w6r1TW/5nZwiFDFM5UJfT54si6kZx
iuJALXP3VF3Vbq1w1x4/NWJpkRocS2GQ1GikWXRdXogc0sotFasUMFXOdRlNC+3z
4uxhdHc2+J9ZBrvfZUbexIDtaWZ9+3s7+hwtP3zGjKM29fbKNs6R6HnffniBGrkw
IADXPNlp096Ywp7Sc76EJ4EbYP99ShZJFrW7/qB+N4exlL1PVBcMhOw7V8bT9z4R
MHXWSE/wdR3qG2GmJ02PkUcJr3WXYrGAN6lal2IQHoaAY8QCFEWlDF3gX/vypTQU
QxUc7QeGIrRWRZXqZQ2odgWeMqrcYtb7/EuOyPVcsoLb0d4Wqt40OaZJHth6Wcd/
NIy4L2Ck5Br6EnMDhr7pSCxGcUTFn1ei7AkAtH9ArOq4/iCOTClf0wMN3rL1tRCF
wbA0NiEdhVas9xG9/dX+Y0zQDSck5CHCcaDcXBNAuwA0oBlp8H/dnwREg45ZB2di
ikOJ1X97slZDInNRa+Lfk9ZEEMD0H482kDRszp1DiZuwaw0P5szuSGEIVx21KeEf
SF3cmxMvC3stARu2R5v4hMVb7SWG8b6HLWE5pcgLjQOymP4fToqXqiJMD6+87FzP
2N8AdlhsR6bv5U13xYlkpXvL23BxHtYs4T3aXxhNCWRTMRDSt0Ia/hP1nl+nnH60
SMhGd+G4BEb6p1uq+1rCUHUna8vuunAh6E7l15ViJ5KcvIHWlfOBvC7XlMTMvnrj
VleW+92LzkXbGWQ4zt9z0vOYDE20aUJ6bd0PktCnku7fUTYck2QDQrRy3n8DveEx
65pisOY/quHLLQgN/L1vFgAkE69hc4nK1WMxHPRXhnda839BkpdwvwOZY7Vy0u9Y
lb/i6Mjnyrp++7mp10wdGKx7hYK1+T7NDRhbb+j4dOgkXPfD6hE2Cd9ql59EoYbX
ZNfzhISmZYlOI8iNXI+4iDjiraYXOSBnCK0j4QmU6aKp9mJU1pX4hxSRQXnifpCe
fYJFsMBdloIw9ccjMwb1GwN5lfdS3YF4l/BJ9Wcq6hrduHRZa4g2hAxeQW35fj4l
CHQsrl4I02aaSrh9A7h3M1UpKjq0jknrlM75YBH5lC5RdeUUMAwpHYkwHIuiR1gr
UMoRsvs3i289jQW0PrN2t0giSNs69/3BbvTS2beTj6VRzJA/rZMt5dq3DWm5Mf3L
7X6IfpuQCqWX1dc9Gmn0OL+VYbwMYiohfr/4THspD2FYeoZxGpMcw5qJhMwEAluL
+HqC8j1s2UAN2p1LP0PTbN2Ir2YklMhaTFzgbg/d7AFJKVgLtDD4EMG9SOmKHAiv
/tSZjzAD1TYwSb9i1c6Ka3xr9WSnwG3G6JS6W7qJejnN3uYjn6L5FDyz9Q//3sj0
hy2VcEnAqRtfatrfzq6HQZzNrxHkYY6aIOyZmUTVXYHkbnb/5YBjzjj+V3jfrcFE
7dDkk/jGTG+G7KnRC30vMDX4NHe4uBTr7XDWyX/NP0MUSIFlIUOptoyGHhvU08HR
ELxo6kXS0RjXVw2eufEvMMoHY/fgLUiwMGERb5KOy3jrdLq7OjvyrBPOZRmRR2r8
QGoLaKMjnnypjklNc+T9VsTwlMo6prnihN+csy/xOXsJW9Dqzvn+7JV9SkXSnosr
vVpyG71dSfoceRJZmQtdqQhUxgJQLHecRHjLbV3YUc/bz/1Asa7k4KKfxxCTeOnC
4NQKBz3qnAXBmz7g7dGFALZXTCiIPSe3yP348/3JgLAHVLB7GqhXihuCarD/lRwc
KH456QF8vyrpAA43vcXHVSbbGUvqTmfGUCiJvd7OhiRGK+DbkvORHl8m1nDd6OrH
HKrV6cESmnaW+8UMp2lLg/TOP/Lmkyrw7EiOtOqIb83oSmfk7PEso3bp3Y0r+lXl
JwP1Uk82gLmhlOTvMhhTleV+8NpBWguTbv6NCHxGWXgdo4i/lZkeZ/t+CO7I0Fj+
CoaaSovqhfideXrPCpMtqGCDRKrFPmZxKhZ9eUCOGV/nykif5/a/221khoKcqtck
3VZ/qSWLZLeYSUFGYPCE8QVUO4V0esdFvCKx7AcMiIoOBCYHXd+XDfjBBarCqXtW
FIocWqUZo9b77NrhpizVcpP5nhmaUJMf7CNOgchyF4uCJ3eSH2HvxyELqkGMljWi
nNhkeHgm2cFymIX5PxAkM2VyiYHClS0Si5nTl1YsMX9pC5pXLgaaxlmk/NxM7hMi
Wxg2fADpkUszpTO6PkHJWX+Wfvh72x5ASsHUj8RE2yS3GITgzMqIg8vkPe5hhsfY
cM2poFsGA+Mxog/1xGWpmjCLPCBJVwEaSbpWYqmXd7iyboKb68nOYqLm5fh6Sf/b
OdnC+snPJ6ReGHGMN+JmKMZWMvIt94/OWLs39Ko8bO/qeZTujZviPKcPjM0IHxHA
eV8veY/Sy8kasyttLIZFkBNQARp3cB4WBi5IDiNyNajdAheNOWz+GdQy32Hb1B8w
zOYykiVOoiy4/owG77bvrLFLBsCMC6F5cPtTD6aFQkC9HW8ywzckZc8M0DdDlR+F
M30HI28m0pcxqSRO20U1jj2WlY9RCeYTRje/+jURYwRPkfByNfe6Y78OMOx8n+EK
BKClFhe/6mCE76rBAam17oE3t4WSF4LBJ5HkayX7Nyxv1/D0WEOY4pETmWX9zl5t
uF2jBd02t6bse6cxPDn1hdE9qlvPPo9U5Rap2iOd22mZckzviHakADc7zikKw3eB
VEjyhS+p77urESC2YsPZVmKyNuBRZaed/SanRS/N4tPiz8O/iUwhj8gzaYXLRS+6
MhRNJYUimMWjc8bjLfhPWueA/YQwsUf9urWO9DqdrPBxvzHJeajUenBn2BQx/tLf
VwSkvYbLKIFlC/EH/EKlyTHzTBt1NBOGaiOcE3ll5eUVE3Qn1KhXY8KeNM2TwPRZ
7V8ykDdJLNwKato8ozWu29xu0rU4dMHuarnY7J8FgDjJDZqAbfgyN0u+RvdEtydZ
B1Sy5Wd2D2ERSnrQB6d6ca+RH6qvLqAQNot4rzOqLI22aFTs8t2pEnjIWTOL0DPY
vRmS2ve3ryzbx59ctb2EbUmrnzv47qqcoVZxqPPXLoVJ57/4yDm7Y82I536uAIRs
IturDS29V3gh9GddyS5sAQW7JNaUqcYMo4hOSWA8jO8THx8IvEJGpNPpFH1el0TF
ROHtUSJgWrzTA2vDTfWpai0lLeM1VX0ClqwLWGh/zKV4OUaS1AcGg7i02xPdYtHb
L3n6abQ+HTr0tx7Jk5Uh8bj6yAMF4Zfv4fQkFZVOG/Y799w51MfMHLgAR1t+RAD7
ZzhhYRKYNi76wY8sKAQ/2OjiVF6nMB/s8EWbhM1904FJ4GfUlNZp5ScAmeT7WkD6
TxOAxIf6TMhxLWI+EclT5G4fy4NSoUunHrrIr5fw83AXngZvwvED7rcyEP02/IEt
UjAgo90zUyJvY7gsi/5PGvJJkgZ1uuss9SrRhGKvQT3DqlpIbVwJWuy7I8/ARRgO
Yu1AhM9wpsJYveKeET87rF+dqSmKnx6uf3Mizd6wXWCj0f84Qd5P4Kga7qBBKXHQ
tc180xpIxqps2lSmQ+37xEC2SqnedvhHK8yJz9RS/4GCaw++p1WwB8W72PTYapb2
ts/jc/Hxc+G7DgsW5zQ0vlJvFx5RECBm8IVQb8Rd05FNnUotXGUmtpf7Vt6YHdXn
oCOAlzT0opKBSdmgulWCAs1GoN+2vUiR6WJPN9lQkmP0Z00XRaCNwYFQdLNbX2Ws
jYtt/oLLCgfDWBlVhjfCUFqvG5uz99Ncmmi6yHoEExGEEiUKmYJeboy+YrKpgMQ5
TLoTkV7QVrNY0ekx/h+ORLIPVn2xHQhsT3jyH3CcEQGDO73MZFIPjeWE+vnSwTCQ
FAxJVbFog5cyKcEBkztYjZLYoK/uMdq+rGUWXw4PUadkD1CB2J3fyB6SGsGDx2gv
v5YkLxTiFuGNcTkJkzcK2raQxNTjjTcQytveeKcZrWBhZeyvGNTZYQ0g7HbR2Bd2
9V9/TMpI0uYgzRETCAB/Jhvynkolgy/DtZzjfSrcQCzx0gxooL/pquJDQbX6wviZ
2FUpmRZVL6ZdR8eXas/47jBp+Tn8O4CeLIgeRmE5qxFKVV6XDUBfglXhKPT45Egz
RvKtoxL5YZoBJ3Ljvp62jz9Af5nt+VCSc7zvMFVTO6u44RjvBlHFO1qPbnFzech/
eZLpVQlWMBu/Q76BzBQLXYxoC7xGa9Q0W+SwNbtjWKr7nq3zyiRYcrWEIE9vU0me
Kc7q230WEvo9PjGqTWnuK4I+w3UerebBX0STw27bwURg0K59aBPIMuvRo+PO6sJK
wzvHdmEvwE1zJ5E9pNWIbFK2oRgtUfg9i60O5r0U1noU37dJnjKvRp7UHbi87NCC
corZP0Hg5SFEJhfO8mGZZG+TXLhp5XutQtXbS4JsgEwTmtdpBzwWGsqWenKrHLlX
H18EgCLslnb7tnZfmZFPsIwldChMKLQX7cohBdMl0irBOnL14l+KOGQB8lxjYOAI
DeJZEw3MIzEnzCi20WNTPJWemgc98JeXdRtaS2LmsFZ3fdvxT80pcPB3kBjl2U/2
kvKNQpkOd4W7B/NSjfNZJxyW+LMM04ag5XpIsYapD7xxkePN5ZaD/T91UjiShPmn
HsaGKzO3yC50Zee6VUTU+yUKZpbzXFSTnL4onMqQF9tipiqjcVEWAwMUFmydJNaA
8OuuTO5sXfiSNGgCDlRc9vu/CAkJQdlTLHVCjztoBZ2Btqg2qTIOGbJCGcyuCYvA
f+PD/JnJYL+fWpc91cQ9xFX6WQ2kTOsUDSJSa3+nMVXDEfxoouoCRLSf5tVFrXUC
b4DvLv6v027t4OgdLpzF9xsClawdAtKtw2gHTJxGus6QIMB8rbZQdV7o3NCnPIle
jew0JZZ7lNu1/cOoGVqV+EnkS8OW32HT3cAyqILLh6twc9yVg91iH2GDMxGoMk8I
F+w9F21ehg58q3dObOAP1vlXHg7l5TqGrhu0c7br6K5dNpYsQH+specnkEFGyuGI
H+BFbqI0ZZIBdsaulsdL89ozv+snuRetO6zvevJTvWxv4vyIO/lNI6ODz/f25OyD
T2/5+GNpdNxO19ImWHGnqWSTF1CLj+wM3ASDtZMsuPZkiszyF0Fa7nBf8R534us+
lx/9IxkGdu5HDInPxOfqgvtlvmmd3c+12AmHFkIDEgI3wqS34qMT+tsHokh6Wmva
fbnRm7OYYdgfaDkZGogwuicgO1oAJZ68fbGCBmJmyD2NTepejnh8gsI/+FJpIwP1
XB0NlNfS14ln53ck43PkWjHGGMr4mK0SnodFN9nHEeDP7LYV6hAHgT0Bwn6lPv3f
Yg0QxU7DWWDcIcmHTk2bermg2Toxn4Iv4IPILHADwns7ea7dL9j9YP9eTi5A3ZDP
kO+pmlV+laybIxLoJypTZ09bvZE+xCz2PHw6U5V0jlr5bUxoWCvjuaP3U42dtGpp
K6Sou+I/RwNGKxbbZGgCl3aW76bXYwhp7X6RERWeha/T58XNVHSoXMpVPvSGRWx0
z/ERyQvzWrcX182J9pH+zB8BOLc0OgGoZmBKUc9UCkwBALnUADOyFXB7p4JFnJtL
kJ8cgzvvsZ1c5EXyGr45OLvz9z0xjKIXMnhTj3qSMO57udu+fnZaMMxl6yuctS+b
OWkYqw3vAMAfRkmzzOW97l7yXwdmZ82NRaDBkby80oHO6C/CU9R17EeKedies9vH
2FI6b/UoJ2W2H42iKSYqq6k53R3FcfPxVNg9giwq80rcurPxBAHKDUT1FOKQRGCh
vT1dRvNCdHCq684Atz8aWkoDc+B4eNGYBiL1neyEtTB+kE1qRNmu0c04pzsAUkkX
5qKdhX9nr38LCTDXztJwYYExHXk/uB6xGpu254cETSJD+s94ggXohJ+FfNXYuERe
xuOdpOQXbLbBvsaI6DhOVqRzm2dOqji4zq2MFi6fEv9S1MDdPscl4ONMcDbo2vya
ggocgSOmuxns2ZeOO3tAxTn5ONZyecQpQMhVdhblG1AhZfS2DuyhOMaUapSjBln/
Ch3E3E4LZf8iQTliCE3DYFOC0MNrQiOHy6khxkj7gmPVNfvZlV7LPsk9n/rWwGrJ
QC6Q9vuSMtCtCnHtcUSLcQnPgFRVDWYY4dMX+fKMWKKMWLuHZ4y+bnCJuQQehQ5R
kj8ww5s2e5BBwV6tAy8HceOj7WItp/pR1QceoHyn3k76Yo1oH1wbKBitNPN9CPo9
DtFUddSHPn5+ipWavABGR9pBtGNpNyEAt+Syu6PM6LI83v1EqljbG1TH+rmxjBbI
r5Dn0R2KzL8U4e1twGEhOFIMNdCOcLhP0EeVduiI4u1Q71ClcTGxO/HXix20W2XW
llDEAUi71z+pYwu8WcZ1A7FfJ0Nl/XJMyexqpCh4uN16QLP9EZen32zhz2CLo/gM
yN5F5eO6RzXmRW3+GRznrFADVi9r679KhqRLP0nYah4YKjlVEEWWJj7M/nu5gN0M
KLoDb2vt6cUeSS8pTiB1gUxyvhFYTinVNGYImwbtRjUtIVjcRAiILt7ZjeZlcDe9
gwjb2kIfOPFk3W/4KApSR3YS/jX/Ezddx82ms5mU2DKWig9eqsV745TrHS4NxeFH
XzE2BIJxN/YQKTRdolm0IKlZxKWZsVcqwOqtjk0nkE8K7LNjyZo5Kfh2u3HbUHFC
W8MZ9Y2Z7QO/dQiyNywiFNUAiZov28qa45Xa8wMQgytYN+xF0bDkUVla7V+IMFfw
K69kYow931UktpyHKpEFi1iwdBj1O1FVX5PNV+SX1faUJhkhjCX7Uvox9MKp46HF
k54cWlpawU4B3wNy0qTqtoN2k+1N9XMnLaqDB8GppUIoGzlP/xuD2VhT09y0qISf
LGXv3xqmlMecUEJpLTBVzVwFyHnwgywydhABFUJJUyetuUIUZTD3iSMgMzevft6I
8EkhHmQniVvChPRhFfaAjzvBzEdKPpZxaisiW3rGJX12GGjAmB1yGmcoCrgfLvL8
RFAEz0wIsG7JSVqbur5eXMNFOJLJFP52Ia2K+AAMKhujhJlngEhOi9uRgLSOq8Qp
deTMQgwI7j67h9GqAKfblIs8E+woJfQ4GuFFeFKhYHuJy7VHgyerUYX9pjB0sb+T
bzjEy2T39pgU2lhuTgykenKKSzpkgIMxcMaaZjs9dOeSwVVjlpaA/ZetywWvBVWF
rW6l5kByXJpZ+qLxLy8EijU46yDcPNyOMOrMjxEkzik6cVuXz7oqkbbAv8Y2jPxB
4nwgJUqxUqfqwSGqkMwdD2RFm3Zo7LSi96EDk38peuu4ia23YHFLdk/aiWb237uJ
AWIR6khZxBofcsomQATd+ZfDPTyOe15nT83rgJZ0Lve7KpHvjSeaeO0Kg8bQHHo2
D9fzrd42gw/qpDOdkoRxW5wwcCJt17oHus6CpWn4s5AK6wkJln3sYeTLN9RToX8J
rPKYxtK4gSjMGH2zp27xxRVh7MtFPJ5D4qa53Slqt8DESYZDB/K0m7RW8GGrYDVS
GA9E/h64n0+JyuVeoTJ6MDa+MWw7aHwreZfihWCjwNOOO/YhUEUI89RrTg4vguTZ
3vOAwBbNdtA07IjrZ+ZVg481nLz7ApeeelZ6g1oZHL97KvIgArz/3yfirTH4i7/S
PYQhY7by7meXqrWqP46zdIctJpz53pG3l75WaVc41YX3UjfzxVXNQvzUPDybhjHx
5AYvpd3LNRkvcBO+FZRMNsi4h7+/INe8NepMOAL+kBwfjmdlcdZEbrA3F8+V8wLM
2cAdmYN13BhDoHNoL+w2waEyF1FLX33CFsxmx5NSmrw9Z5RhgUn3Yk8QWijpCbUC
LgrgDWUOUVrL9kIiEVmHiufVPuBrss894NFjHfU5ioHzUp5gv1pMxOhaXyc0spGR
AAd+m4xX9K48hE76dh1tgYwakXbZL0WB7T4eme2vwRmMC9DbwdQqfKWcRv8ltLEF
KshGrwg8l9gjdtRoLUek/Wf5IZs+RhZDdCIfr/VnHve+NAJSVW0lcGt2XqcsdGL2
y5dWh2DTrOJOekfokl/13+xO4y9Dv5j8petCb0Np5lrAQD4kZkXLr0EvIeRgud/p
LaQ8b7V83qts6mqKIs5Sy76W7QpzZTaKTkR7C+sGZzDpo6Aw7/L8QtvGolZPpXfX
hXVqBOrAVPPn3d3X1HonlPGGUohKQGTlIRhjz8DEvFkFs+FMrLZ0O9TWSKEo3TMw
yWsMPGTAgp+7u3WNo1ahCrQ4Ue0f3Qn+kF7WP8y0A8qFmzby1hstP0DvCQSlGXal
FuJ/4fcm5zxjvr4LtWNvxHNgsIdZpXFWhDReWCm027/+R3hmermuQ6U/3+JR5Hxp
1p6jXNHjy6B8V5kscW9fVYcnGzIgRZ1zuNBBvWi4BtM75KsE/d5vvw0iUzisNLqU
lWi4cJEGmFZLirJpZsw2KP3j1kntpPC+g1W35pW3zf8ddo4z1Sg0jJOpIuofqlF/
vaYyXjIxn0V04EpiGWOo3pPeDoaOHQ/E3UXfETDda/D4dgVH+ajpIwD3soubvCU8
EXZqQW82hwKQoGAfo/qnc0b0D4K8FfaMotciOdbNkCc7KamZAd65lG/4KqJZQZTY
VFkMf64ICKBahJR5i20qAkI3rtxoJglS7dT3daExpFymQzteNnkfbXNIp5M6J7Ix
eS70mhPfcY3XyTG+fcczADfw2qqs2eTXFj4uE/yeDm3QQJdkqYCZnmo6a41rkkhT
PgjOK8U5Mi9by7gmQ2lYkcAPN64yn3/fyaKyC8e3mX3u4qhuSPXjGhzjxY5Xa4EG
EvX3wnSsGO4msErcjqEGABNn+gQdK6AwHPG9/vKa6B/BBNIrStaXelIm+w83Sdk/
wfphgJh1WzMhm/LCL+3Ju+4Nyd+xSdIPbKvujQuU/weY4CAw7GlQlP9VSJDNezP8
IajqU8jwFA6OUEWWyZWKr/58O7HlW+NujZkVUr746xP36B3ZyrLS0zexhhQzYY/V
tLOUY5uETvufiJkFDdN8BmqbTL2GZfqOXc4wCHbAzJVvIIcv6H5QAG7Z4mbW6Mp/
5v6OV/Vkz5NQQtFNQOf4bW2zFg7Q5H7mCKADhwjp4LCH7WpbUeuQaLPlEopZ1tgU
gQAXltFLH1wn0DJzfGff8USLePYC39FgcxKIH8hZylB7okLeUhNFz+LqHSOCbd4C
Bf9stBIqvktSlqrcSoWscK7+2NdZDnqliDMGOhRgWsag0fck2O8GqFuCmBavX4bY
cTrtb+gKnvEqX/+6rvnjIb5KFLyOBEgSEaxWtyk8ghaaIKoA49/peBEx8gTxeS+T
qRS0HWMG81SFGVxiwVTJ5DfUaC4E12bbRDcgZ8Cg506+lemSh+AfV8fQ1eR8b64o
YD291QsZkI9X9VV7ajp9cvI+YGpUJK1HZUR4pXDos2+RCqGyCuIEPqVkhUc2wgkC
1XgRSQdzs5mih3uzHN1vnQDjWEpO9wmZ4kek+4kzZjjIO3nK5FGi3pwjGhLBH77t
9ua9o08LBF/+FhVrRKbpJcvWYMQ18TlPCoVA++SXSgo0cFfFEYKz0vfGmmyvjQXI
LiLds2kXGhtRjH0MgukoCmmhMfKnpDUIXwqU6aUSM/g+1VywimKThaYIBLz+89R4
Sj/OCNTsElneYsQG5dgaANM78Qi6XpwOc31lGxkDHPMJt4OWIACZXIQyhlJ6wdvu
D77ZzuwruVtgZLi7Zbq9wCJe5BW7aS2KdVa+Fcd4AN4vWa49WCjvKlztR0iBy1bU
6ip6WtFUmJiLQDZx9CJDKRx4kMgA9Va1k8bZPfmgGnymebmtz0V05vFjWXzxIlH6
rKz2DBcQNQsY9N0EpjpYpKCTH8+KLQYbL1+cBBROK3RNIt5lqQ98UHvaCchAPx1Q
qTHj/6Gi12CmM8qRoIQVpzMmj4+fJUGofswMpRtdSstDtjmZFxy8zQ1rtd0zsVQT
stEGlLH9Zdho15xiczKGddVi/vGC86+mmF8MzGJligqK0jWqgJ2rq2tTaE4CkbD+
eFX/MgbsrcsC07YvrVKvOBzVMMYO+hOiJTOLw24PmP4sLmvRYfVgVdeUjZa91tGs
L9gBiSGQTI/4vTG8j9ITUoBGa45Kgz2GhZavYm7I4tTK0098FJrXYdNC3HkDShdF
13M9+IAX9EqHGVD4fCzgPJsFjm6kbdfCQJjjpqEG4tWyHg1YprATTikv4O+oVvmK
fQ4kxAdq/IAjZYPf5eB/oUL977+69DL9cy1TsM1QgTHFpNyTLBE/LYpECoChZgcA
GpFpaSTsli7vNyYlYAtUJS2MrIPo9zsm0mI+Ces6ELjTJE+vj6aXf25GYFm3kfyS
Iw9kwgwzJL7t9moX3p2EUzwyqZUogY9FEubnKKYFdfhuvhGAhbA8JmfSq7FRkTaU
U/ivKZKlCsXBCPGVhfIBc2uhpiUXX9HcJNtfiTwrTQ6xe98SWv3vCd3vgNAeZ07l
Zb+m/4KY6TZfBEDwe2fcv/K4CQH88qOeP4qiqFtV57WWbkJ0czWpdIdmvnW1X8a9
SgFYwyiR5cudxSxFfoglN1YLrPMaUiEoQ/aO9SQBItrcI9ID0YPWYAve97NXshFg
7uyFTa1ZulX2q5YZ4KcVwX4jKeUOxV4RBMk77qqzaHxG6KiFqpaLsV7kFh0A3DTM
GzEUXpmKp2TWbIVqHV0TnPL4LzICoFLbhEC11g6I4BBc33ab8j0P6DxcSynUU140
P09GZA4vLJrf8UqXhu5P0TW1ourkM5doKOU3VAjm+ku+2s6YPNh6qjm2QSa02hIv
fX1bs1v5hcYQafsEhfB4GzyFyH8TVRHZBLk/H1G8MKRj5Fc2X9pYZ4gmzD0sKNws
Cv542+O8HplNog7JX3rh7vQz533+ghriC/ghjME84XPwDdh8nqwlOZo4WWWfrK1c
VmCpRfHJ6KwSAptaML7TWvkqmbBwzamlxYjfkJqL+hHdaQg9Gctm/S8tR5+BH6bB
TD33aNXwkxaJwALLkjPuASNQ47zkgzD5jF9c2CLOP0LliRYBmc3pdhkEBeZoeeps
RCoo/JjYit4N8hdrJxV5ab8WhRt7JKn0cpe+zwyucjlX0seFVrIpIxRMa5nZxeks
OPf9NKCG3+BDqaAwARg94m336Vst/6rIfSJvZnD6EHq02qsk1S7XoY3yBIpyzqnk
v0p4ODsql+7WzeUVZ0T4Z2c3AOaaF5FaYyz4rDm62W8U+8hKroypFPfKiiObdMfC
JIUEfuAStc8yqrhlralD2UnGToLNkDDK9j4NWMrViCDRCKIHoTXY+6yP/nusS8aK
9bKde7/bvahgPFQWZQRUVvSLXJuw28jYFWeFjKzV0h8Qtzoglpdq4TF+WfOR8R88
HmDzpl8zxYlOT8FTRWX8gFrSKhjhaFqByrJfkLkEHNtCgl32mipO3ssJdH3Ec3nx
amvJhRMDDAXVjXBBmA1JZtbX10P9XBr3jijWNcl9fu1NQ+jigTsc2uPjgDlfdzav
IypEnQnCfy9YVWWwTuJjkXYGAiydj6vjNvYBmG1xEB4FQfEVVJ4sochfUeSy0D2b
qZi+OmOgbv6njyv4iMnPPZRYa6gLk6lsuyaeYtOAmEe+h6CijSgHzaJeCzk6V6Qh
FaBy649yfAuEWQRPfC0E7PgHLNmnZtdpwcA0b9036ICdFoulMVpcYo+YxGAL6sfM
AzfgzpvqfFt29eBsoRCgcdVcSUyTgqOKcxkwXfDxynkI2RAtt9N1Q5OEioFUB/MH
WNxQuZrDEFl0hcP6wjW+3bTCJH9xVx8beAK+NWGk1iYNIvQY/7fC40h1zwf+1Y0S
jkS8g4DuNDrYNLcUgXBVQPSmfaTA+7P7SDCnOmZQy5u4rot7BYbaiO0+qgJmWjCE
WVhuW+0CNFbsjeM5Sw5Gb8rRe7DDQbLjnBrmXYQdSrSrUmQDPMnjGamkoiwxJXOu
+7NgrPZ5cvpLaSzJowD5OQxKnIEzsk8MBb/htHrexQuNbnpbF6m+xEHZz4i4YqPy
QygEOjYZfiO3tXjX7kITfPyWHWJCHQTFur7HGQFdcqhTd3TUtcy2nUnWPa1Ckvwc
QcxgF6d2msWiEFJYVlvZ4ywc06IHGMMDePBM7rujWdClepOIera2nJoM2P4hTKWO
WpuI61OtlqdHxoQfIj0IxqOOrDuhtryNWngpzSEDVpS1NHBNI6703ai3xFk5S8YX
we6MktZ/MvT/J894Jkn7e1tjFpsED4h0PmJqw1NR5+E7+KlNgyXRIOS5I58UQx9S
P8T99RAcu0ErLyKTTlfT7O8Hyl5MmefMXKDp/+zNfBDOxaqwGHxEWVNZ/Q6WIHRC
J7+MbSc6sAaWfpKJtGIguTANu22lV5wlMMjOLGBSGariFtF1jNK2epNKar2hJIFj
qgB8ceX26X9O0ovGd7WZ+93BINwWjOsrNa0ma5N39ebvsQB8Bvr1MjfjA8smocef
Pbxlgd7OCT66whV5dofmVW2ikEgrt1ePbNBFSVyA2nOgA8v1FokDHae3YQY83YXw
plM23AkmTQutEYZHYWC+2xeVcY3DwCV5+ti5iiLY40VG6npA8WMAxI8dcqYv1IZ5
YUBtQKlH0PWVqJTOyWtjFa+yYVEn/PUWp1v3pqELdHe/PwHXxndP9/JxDS5xQzys
/DCXU+FAsJqXCvhwtFIXokGmwvullcGZYWJA5lVqufOX/lWysRmJ4NAFaS+A0iBP
PIHnLrY2vQuwHjOaLuJW6V6jKbqIAm6sUEtJavEjstt0/S2gg6plI6p84u2MyPIP
76U2NOI5B/qDHSEVGhkq3iN3eT5+gQCQwxSb6Q+ZCqPIX/gUEsHNbBwW48Rzowwk
NiYndxRptyzuvImjgT0mg38pFND9YViBoLi5vgoX1O0gjswduMMozwZ1wFG0JmeW
HOPfn/zKoZpVB6q0ykrNxbw1MKVEZSn1jqk0T8VSXvbXhZWJczKVkA9gZmBOy+ig
tTG9A1G9RCHlsPenwLetTq/ZDrLd36Vl3AGsk1ZeaJklKm0Kdj1t++kyU3baORlk
7MnUZbm5pmjvXf4Ge72H/BcbbNaK1aTjyoXqbNKm0weRjf/cZNO8ks+nI1TZThw6
kDvfI1LVwdf3/Rorao+fdUCiD+QrbaKVRYPqANB2OJA1YUsxqivLekeW9V2xRBmP
42tTIZfluKG0bKSYObqQq60KYLKEpOPShDPqkr/xGm0Vcczn7GDwq4PkU1nlPg67
d/4Ps8zIxgv8SKIy7MLQSZO1ft5gBiakhCuOEBGibKWczfWsBt7k5mo6w5KM4Daf
9yxa68VCWFLjB/oaKDCb6XT0pqYgZ7tWo/mpsg+Z2MeYPYq7PFFZaFQ34Hqj46DH
AeJsQdhtET3YLurqQTzGvWJLplhvMSM4YMOW+esiNDFiYrEYWOoxcM3il4j8UqoW
7CMmU53UARbcYPHFSidhp3S2KDzzpfLx1MOt0SKrILLtxWc64sx1g2fovuTKbLVz
WrWT71rffeZflul64ISyfIDPCGbBc12FLlqVsl828QYC3PZRLbgS7YCC4ewnVQto
cZz8aT3dzMxePrLHOIhyEue7kO6FcL2dVKOTEHdK3qWRaSIBT4+cQW2SyD4EIi25
yR6Edv4IYlBwG6pjvcTeONo5qIFW/YhTI23pDrYwp//KdmpDaoPqwLvUnSg7HnEl
Bmbry3fHjUA2ZaREurV5Pj6r4XlAvkxG5RzaSbxZa5auiVW/X7Xz+Q9Y64RhwiJP
/QOk/YD6yB16TrE/qr5I91PTE4P8HHGsWvgcHvOlQycWnWaIUBHsKkcB7RfajKhg
dNwPnjEgiY6GM9mZhrbG0hwnq/cHWF/UVL/wKJ2mjtc3L+ic7PerMjYmfdR+1/1x
E9vVlKTl9u9PFIUhA8XSB2loSU+rRrJCZFpMRrGCtZNPH8KzOYHBapMOCG/J1hxd
dSu389/SKTJV/4RWFshCp3E3x6HfptuMLPBLGXAZ69Li11/NQsWsCKJr/rnRO1XX
SRUWv0fZB+MPk75GntFlkmoWjBcLs1jJpjQlFBKWB+ecA0xskH0yAcjgGV42O3wZ
lvOC2ZAtNLTp9phmbDKdcE+ACG6cAiirmVn/HbLA27AJOZqekQ1cBlj2vsfGDOgT
IWo3j2o2xwIUt15kZQm6ymog+FPDutV94vVPSnHnIvh9vyv03uuWAT0jJMKMjRJF
N5+lVsu5Im8hY2psOE5VpMRypHiqiEBpa5PSN0Crrrvq9eZp9/jxVFRF9PngmIHW
TX+AopmbBJw2jh0K7of195mE/SfLOTbHo13vQWojhJjyE1GGBIRU0ljguqvQawfT
WoE/GSjnvf/o83t8qglmP+9kOVdHVd2bGr4ktfzgpK1gZfhhxgQu1Yj63tqbJAMn
fF3yCvDfTHw6LJwaQMDh9OtSb19/TGNjoKCfIPn02u7fRvgSDzoSD9eHIZMYS1pP
AOD1YsApQ3paBTDTTC6bO+LaUPVuyx2pMkYD5yp1cQM4h7Qgtk1PDhVvFgySPKGX
tElljvvJDUzHcxlTGfDh2mAaPPNlbRShU6w+B0s4RvrC2/nAsVR1vT2GXMehrgQH
6bsAadzP8MJpFSqC70+vxgcIEID3v/FVhYgDUB+r+SQdEqsVPwG5xEmT6tMe/F0d
3f9S7pJFSxUjY33S3T2B1dVUNjMyAA3GMGn3oSup64LMcRQmc3bDBuJ4Q7jUs4XL
p1W04roTLroLyVz839K/5Vf7RE3AjoO/B45YN5exBXgDtDcW2i3FiMfr6XmeSHxV
tOQ+YwsLcrtblz1IhnkA1MaypAV4z97PWDO8rz8JO0eCVghUdADCg+EcAoBaFiJz
gly5ABFkDBp40N8ZbFTp9gyoMaD3S+Aq8MCewupb6Ae7XbhF2GU0L7GjvqJUAZve
1O7isLNgPgnHNWdHU0giZcOx2kxo6gobYlhdXMga3edFiPPlKu5iV57lmbz96YQJ
uYRemJpOXoKnwPZ6DAaVePV6IV4qtAKvN+1CdBDBR3/cxsBciGYPo4Qjv7bFZfLu
95IWbFG0HzNi8MGb2XRpgbnVMm0kWMtqtn0X7NHaz4Ln0C1qkMBLCQ2/uy0a368f
1q6lVbBPufOpMqTDBDIM3vcaZO+uxePM1LjRo9X7zl0nPNCdYIBdg5O8vbhbtr38
/VC7flj/eU2Y0+diIl2vGBbPAyM3KApp9A8MtpZy9yp/UaHB3V9dlWO8v8SruW6P
rUrtGCuDpo5P+/kSQgTl5IwSVXO7a8f4JEMCHR548UXprtXIX8bo1nj1X5ClRipI
m0QXKTendzCUohiWF3xoLS4UZzh9P1eg84E26kYvWhjJcnZnLNblN7LjFcuRQHjm
K1rfK6sGy6dPhSfFPEb4BInTIOfKm+vU4UM5+X9QipkP1UIjnKvFCzJmwN/Lo6cV
pBT67PNcrxTS7d6SfP3tKLJKFxNM8/fC8NqDMOCDK0wwTaZVwdHOLu/lrNMoIAIg
TDSXgDRAtBcQm1hsqSt2K4OZpqaCLxtXUUyoiE2UFLRIChMuWfE3WkOtUuYV/xB6
CPBI/SwVACSXRbHbkygBfblgC3K5r+MSYbxfdlIsNXvdBnEBYnn1DKf2Q8EKW/kr
thZZFAhh54Sp3Rfo7CVIre7GCf9mdReuXi9xxdXcLxjIPj8Pz61NJSInpFIkn0P2
8GA/UcWQ+8vHdwOYhfVNTo5E9CURkfNHIagmbtdd/PhZ45eeeFYJ5LHZhO+JV41p
fZcaczex+vS6LXH6j1Sjy5aDk6AuAS2PqZpJrWA9lrrKnso9BQ0vII/xQCW+432C
F9qVJaQI4am3ir0elzXBE4Xzl5bzxsfpC05eJYLj98wsomW0gKbkQ/6ZriE2J5Mr
D3Rfv0eB+QfnLe4vpaCDLeckSZfx6dGEdWs3XeaTlfqOZhXkHBBKHq1mgYAEIAb3
K9XR7loSMXzFzZp5kfW7HgICGgiT+G+QTzCMuMoU24uq/pnjxbm4WQRxRx6FiSqt
CsADx7cS4n+73bb97NxvP1xOpmtC0OrbU9D984R331tB2OkJIQhPL54yf4KtHKNb
ZmXZ2meVxnpnkuri5Ts4TcwlPpHPbNtc1u080MBA50757o0vRjvgCNcRCBXnKXNQ
kbwC6uao/PSW7tdunwUDyxZ52OJGzkM9F7A/MppEvgcweHR3lm3zCjUW3zDawFQH
d2mw54gUeFwN2HbWjd18MqdOkhWYIurZlBN+JFqXshtk+KhNoWlok9tCSxHllyfv
vD023nSoBmTXPx3hspwRymnNbUFDHuBl4pXY1gaSQLyElABVdJpDpcW9E9sveNjw
WDXdrLMvfwXI2ZsC7GWbv3RyYi3DSJsiY64c92mx+o1i3kj/xqE6o8J1TjyId6wo
MxiVbduk+L6n6xclHi0r+yvS2Ci8IuYTEuz1vuVzZJCcoo2Bm/NwokIXyftvxkfQ
09Dmxh8AkiVWKxnGIoOXI/0uQZ0IrFXmKhipppEs3tb+Lj04wGfpieOJbSNejFY7
cJy3NGGge0he/t9BjDmopnLdWE9PtpPmSk57UqrUYVs43h1iHAnd1TFVWdqnTx5f
EJ+dQ4h7L4MjJkUu4xSXsy8cOuqqvkyveizBq7jC0C1uJrmDKQdt2XcCtYkNW6yT
wiwLKHrprgeWqN/zobQLGrC8a4Nd0Y4uw0tuB3v5tmltFZvTzu6jv/AIGEdn8AmL
QC98ohkN4LlbtqYncWEoPjGkeZieabjowaJyxpnDdYnD/8zm1Qb2qkAuQQjcVW8P
HIZjEOJVC6x7bnxlz1aMRBnjKTdt3ku+htvYtEe7ms1fIvSSMWfWu7buMsSb0Iic
g7oUwPnTQCNp0TMJTEI9hRGmp/c+wwezvVRuVdg9141ltv7HphlBiNV0/ZprFudE
40kgEcgz0Ev8FgtYsFe+NUnD6KIXXP2Q4i4v6EiNnXs3fhDKxVlHgN1azm14gypm
ECDPQAWl7wUjfclgCrL766mKh6eZ2Id1TvsQe9fjjEPEyUmrZ+o5/Lquz883DLES
uyTDHQxHkohcd+ynnjeXTz203zFZhKarJDGg2Q/EM/HN8KTCMJltOl9uc+byuz7r
mz2xS7VWh5QzI9lf+6mKd0dE43NYIRD2Shwhs5c7R3g6WKOaLPsnlh7hQyTMSjRA
kSUUvtIT0YQVHczxYbM2lxe2YWXjp/QOTSTAquuthQkh672pKH5vAqnUhmifbCZ2
6fA08aKhitpVr6pn5jOrwLU8mGHVreA2KvrQdIsCu0MTm+F2x1DiCWjpEMyvaapH
FJbc5iz2401MBBmIBazJiCV/gz/vnsxSinRK8b+pRdYZu5qNVcqAqF8HhFm4BDnX
Y3guZJZDjdEWBLKpYi9taaswl3ceT91Hf5kGKzjqMJMrm0H2Lx3NtklY84fEUkAw
Z5o/IXfMkN+1Lq15uO6tQmIOrrXbaiPm7zHF1rjjqc74j0jlreXFcWYSA5KlhdZI
vznrNES/QSjlczBm8Kzyqg0CZUoOncZV0IrYZ5RuMLURD+uiiDX9Z1etry0sTVKU
XgjJQZ7nnBjrrUwMRxKZJknJHZkbUHbILN/ZIrc45XEiD/FclEFEhKBESq8rFUT9
EDRN12vR3D9/XDBpxlaTYiBRvA/eoayDtE9Iib5Dw6PS5HVqOObXm+pG4GCsIKqe
lXMKHXfdsWqAMLTsGYY5Duu5SbdOhtuwgLcdZripfwYKug+QV9OLi2dCQ0DdLFMH
XcorN2AygSkXyJ6pKfSxdsQgm8u6NgEtyJ19K1PJSBNO4uFRVxfjDjfw95cxp+5y
E5WMmAEDzh2YzJ5a+PkcnEfs5ozoGZnalFxWcFzQR6tkE5jdyftogy8a2SzqGskn
ChXn9mG5qA0bI/k20kH+49ms8IQSCt+OLG6T/Xfo1v9dffe5/0rdPEOCpBoSmnke
97IttRniHVKEtN52OoMZ4fdjnLCgFgnymuAXyLhrJx+lTMJlWjsJV8me6uln3jv+
yHYYQp04l9Ox1uUawy0jbMgm4HywQZ2HQWZ2PDItaRoQ5h7xaKHLCzuoWu0/cyA+
zzkdeynGPYtgpvQuxCsigOI0vEoWAZ6O58Ry+wmbu1etR97EsEibsnFJ4Bg5jJN3
ENf765xFzKL33E/fVFllw4j5nPHPUSxbYflCSchgkcpF7+XSALmonAsS0Js5NW1J
cjg5/X6CYsxnk/77livfvfDFNPkjQTJRkJZoHejovNoynsSt0w3xr5K1CqBd8tok
CyF/GmxjM522SD8veWVlT7jpBCZ0pCKYIquTrbVmCR85gtrmo0ZluYETXTEyZNXh
eIQzWQNSnEzemVZjOkMxYilfRfpYE1p7oxsZl+1LaKnpPyt2jhc/SUUTW0Ee4o40
fkCz/eWu6qK69Cnf9VDHrBZUFNcfzZ1sooHdZo3j6e/jT6ZjXh50KEYPq3RRocLL
s1nVVkWRcYpUIYqcusIKPfr1EpTajDGcCNftLc4n7rW1+f06neE3SM1vVLoL2UgB
2JP63HYX3K/4a/gkz2yRyWXuKivXL7vEcYdImRUv8IA2N/gkB/wFMSle1KRF6VOu
gDaXkdeD25G22NVYIgjjPTdAwwOSKVHLtibzgQmZ27yjhrnPaHm0CyyuH9TX/9Oo
/OPZMZuqqULWe4E4pcw0CKnWeVap9H2QFvZsy2qe+1z4KpRhfBIptieA0+DmEeub
I2PPaf6sdIYnTc1j76M+i+62cM+iDkCIvdyVneK01+jP5Qt3eiXhhVhxNfhaNdUk
5V0A3nMsVRAhdwcaCijF//D96dt1L3Aq7dUpLcvNCQf+OX+NQ2NUSBmqw9tHbQPT
LYqX1kVKiBaDAW/CFsMtN5cAHSV0JEtDe2Jv4GyZy4T2ys+JfwKAmSJSBbpFis+K
jGUuf4olnEO7uzeYPOykEbuuhk2xCR++s0TUy+X6U2bHqUJgdVKK7OCEOQK8HG78
LRde5AmgsUnW/ZGzAnQm/4mEgZl0pZ2yWXW3UbSOPKN+FyblKWlyaKSrWiFiqj6+
jMs+zYT0Sc1BSKTO2e5Vhzz1RdtLKA77sDn8TKZP+EH/J7GWz4sMh6pFOQ7BdBtS
nL153EYHMD42GqjWXXaZJR7zPjPoB6Pv8rgk2W+7FYJPjN3rjNrR9ey4gXrJZASD
F3Edqzm+sO2jLxxGCgmp2Ao9RsTajujU4oniIn6o1vqicXXx4sLlKA1FNsbNNGsy
5qu5GD4t41xUhWXqsqfWxvRP/yzqIkw+qaS7yF6PQWvh2BjnV/P57OLlU8c2wrqy
srdwRjbTiaHroQbj0JWKvrnqRoOJ2mm4RwrmtYl0ffYVpVnWcglYR1qTAj9d3UjQ
PTJiQnoIgzjVEXD8mO84nbNrLvmKKdKT+luHE1TX0TiF8f1xStxZtPaFu/oJ3Wox
jS2Uc3oG26avnbQxMRryh6SUw4t3WSIO+zw/B58pk5WuPfMBYjhEPJx6GMtF48cF
UIZ2KdQJeBf6PUiywJThlyOZjApmy+Vjj5J7TVY2YfP7eH8yMB5wsRnZHJJma7Xp
9YNXlZVfVQ917hJzQATcmkyRVutY8/VtGhIwJxhS7F616NFg8ahwPuXL7n2g+sfV
xz6iIP2e9AXaiHqRlwe2xlDKJFvpdqVCqG76AJV2Ie6/9LX3KdSJvxZJmquswPWZ
Lhq0A/Rn0drC5+O86hQYhC3NFmUVzJ3acPmnNN2llRct3OrNXN9hMuLX7wkx2TcQ
AwLbCX7Qzz2Ff9I95PWXBb/eX93RHSO7IfhTRm4y2OOx1SsRUvT6TSMdKcjuMmvI
Bb0zKClOcYWyN4Co4ZOaQ05pI816syndfhwl95DBCd+bm9bg4OfHsodnmJzytekL
cmIK5f4NRGPAQZ4r5dalhgLLuYg6k5vqr74p87WhTCEHQBBnmrz9lnioBiDxf69e
6gO2+AYQa/wQ96EAtB+9YhoPnXlVrTqaJknct6w6sttuUDzvi6O07l1unifSEGfE
E8ubL4lQFMeu0j3Z9i/kWZIYdGdu6zRrn1vndNDZ+ThOp7/1NmbKU8v/mw2KgElT
Sg5qGqRCH57sDTyft7nAk5frGYwODQw1u6N8cKNVOfae48f+367xIAnmfidneUtT
ZWBeuW5dKiR+dbiNfW6YQYbvY0vbMbSkNNFqVBUtZnyrfpTi5fZFD+6hMKIhC+tr
RD6WkQ5MUw/9WFYly9P2hoQIS3HemjLdic7E7VJy9Tm+Q3eH3ZszJ5mL8nabxzTu
0WFhNTWu2QaYy5sm+LBosu5o2HLw8CL6jhDOX4j2xOLJGbazBhVwCqkWn//YvX1l
/TZM7wpULPPRVFBldYoqXeuJIIywMvqQXEQ0b3B9xXlZVO179x1Nqse8iP6zpySv
EpkU0LaQn5AtkAe/GwQ5LlO5/5iAzXPxVi4mwgcaXdKNgaksisrlgSDEI2tvbSJF
JMzi6dFsOx0kmEGfh5yb/LcrEI1tek/7Cssgj+MDgHE7La9124ae0WgfNpOHXQM+
UM+xSCX1y8uARbx916a7TaXmgMeFPwM1l+Vbyakcy0Kqtjb6o3M5LOdPpFAKgdv+
hst+cIKzTvsjyT0fThUgTSM7KQck4xgH/iL59LK/jbogMxl8yfahEZPbqY8yUcLw
uKyeDkApneI4N8pi9ojXDj2lqv6aKjgMYFRHUAvZ4TPs8G62igCrSSdVxXSCtVBN
4QngIPN79icBYRXCjAK1A+QdawLZeeYcbHIuSLvfX+UWjua9Npm8LzJbHJx1RfdR
K+mVoeh64nRFYqBWIb3xD66YQB0528PFwQSnS/sRgw2FdUge7HSpgZQM0561vMPS
+2at/ICd1PapeqW5D2iZO1ASAczCI5x0Uy9VTxyb01fdUsR9ctdSkYC6JqgZG7Ab
fRAC8T32zCyjbNm8AqSrk5bojEYYDXAWSY7Mg/XfdjoP9KafGV7smxEX355QZSv8
r6ev9b6NPS5m+Qrpa0zaolztfa9DjfEOxj/O4nqSb9v8bfhEpGcxUgN7RpCsWriT
gf2uRpAPh5aQhx7+ngx5VqcBVnQ7POA8iG0zJn1Obvc1UPb7Rk195qqVbqStKTQ1
o1NVtmuu00qb7A8FMeCIWgO1zra2UD5sA5iPsiGNTdzSXXt0zMbaFOFRKmCBLgx9
v3pmT1z0flZkEYfsAurKMGJm38edl5PZxnik77BuOWs4PAkk1wkRLqiw2UlgmV/x
mXjS5tM5MuQmh11Zjb8S5GGvU3kAc/0oL5ngSWtVBAoovPneXtodmpOyEhluzjhv
RbcQfBmdS4ZdItNTB3m3wl+RXvRk04aexzEduoee9tnQpoOYntPMo3BTNkY4mNc2
JLPvKN5w3sY2ZxeZsi/MjU3HlOERfKMYQ+cSHB6aTQct0u2TI+BtBrA4pqGONDFS
q9s4bC5Jq/sD0Cczh2edF7WcoL6fLK4J4hdXrA9gjgWdKTDfEzIl1hZyitmp7ejN
1ukQGifQa1BFXAMuFHSSHj0jxmTtM65XGweapSATqHFne/YKHMUhdd4Ud6DVBldr
w9UXkGdaJSPf2XgfjZmBECdiCs620CcDH+GpZA+y29JCTnCp4LgbnsgeFA1fG3B2
dk7SAOk1odAjmaGGBRLL0+pBSQxC6kjc65NVqgy0ZVbG+Y28XrSwp5NaK51CbsPt
hf6tRlJTrUoD6Dg+toFb4Hqbw0ESkIXnsPd1sq3IjA5z1dzLupQ6A12dnOzaC3mU
kjzVXJFAd4G7lXALFyMg8uoJPp2wtGStFu4i9hcGMbCXo4uc9M+U8JkvU3Ls+4NM
1Nw/y4sNLyySXyzI/4qkwXbRxTyXEUeQx75JjjL0/6wLfTQ8GNmgzzUAFyJcVLP4
Xx6Bx36SCsV+gJweWjQmYa4qb9XihmSs4zI/LsQljmtLD1A1s8Ue60KPoqB5UJEy
dnMxp1KZMj6zppAGKrnfzPYCpGC/ABvDpFStiCylGAhBGD9F7xhcrPobdVGb7RF+
wPVaGQiw7FnAXy0pLPfx3EbGh2x+JzVyaik0vlkstfdMBtJ4tsNCt5mLeid3OydB
4GEefzK6HlSo/Orx1iT0LMOF7zh4FJgym7vLBmE4MA5SFbIxdrhGu6oUZ+gREeuC
xy39oeGpj5hhCb+gb6JDaluXmM2uJ18bUj+D0LVHw/jBPnXnIJaWA6I/diCPKZtj
xrcXVit5zF0GRhuQnrFDpmhWuXhK1oCL2Ex7grTBK1k2yfJb5z7771ODJ0N2ILeL
M07EEnlPSQEo+08Gib3OTVx7xFac9c5IsqHfQchM7F9EY09bDHh+U2lcYmhQeLPu
lASvpbkRUFUp2BqgF4PWduGPL5wJqTOjWG9GbGGHacLaG8rs3j0S73fB8qBpR8cC
HLEvmDz9BZ1+DnXwZPB02drRcyR6kuU71IRndmMGslMicXvhPspLaGwhcnKc12xO
Zbkg0BPgPdvvw/X0o3acwxrsmd365y+VApUmJ6kwe3vVXOq8YWn/exjEkfGroA1K
InefqRwaYtEVC9OjnKXgTwJibHrmeHMtTPfZxq4Yi0funczVEsNk27o2sNGbnajS
kqxqQhgGphc3Vmvcc8HIrDG5PZDgZj1bK5XMqcuyomeSRHrHwgYIhsW05uwzVH2L
FM9T6nx+GHkvida6hE2kLcm1fcz2xuiioPfyAWEbIfIXPwBXtung6XzqYXWnJWLM
N9x7cRkyIOANvGim+XNp24LBjjJv8Wh2a8gWik2xvsL/YxFy79WwvJ/Jig23znnf
i1p8OeWFXTobBa/AqNAeNA4nTEw7S3R4vPbkSUtJw/+gUyM5+NupubedcpcdlS/i
HjP1QX5mQULZWVyBoHLTgDL4wW49K7CkTmkiZsO85EyOYoUj6ypyxvqpaKeNO+33
urcRZP5zLf7IhIQFgJ+NF1bTGsFmP9gT+I9VW3us5d2RFU9Zz7OS6qxUsQ1cElWg
HB8u5jrCqIu2YfK0e1SYi/KrT6o8Aw6h9JP1T87SikiThXmzcT0s5yxh7cXqfTqT
nYvsp499sPIGfNxCOCyk6O8m2c+fAmT6ldaxaeXDbeu+0/jCvBrVnRu8c6lMA2Ro
039h0rlPF8zSvUEmKQUd/PdazInZ4rgoiPPjX9VxxPjMEyEjBxK6mS5+RXwEoKaL
gUZXfi0Vhjrt3Eev+RsyL1VlgWDICG4XsWotPBqrol3Ic1yijPLIT+207rdkV73C
/czdz598a88P8mdljnSF7QbbKrg24B9W5icMcd2p4L7svqJ6nrEJKtnMryMJNS1t
m4llhSQnf6Szvi8cSZix1+taxNOv8/Li+t/tcGFAxZUWUOUUx7Pmhm0OSZcbg3lj
fCPvGn2JJYfbJtvfq+sD+/anG740W6UShWAQjJn2AfxkePrJWSDODLVryiphL6Ew
2Z5ktcVtBZ0tyFoj8TAQr3stDA+z3uvCp6WT/XwlZBjVih+V7SFtk2g+L/7n0Zxt
Ku+ceDb7cMPbi2c0oCPU+H0ua3skM/9daFZ4+NAkE+VuynXLHPYTpVzFc2l/ODHC
enk/QqG2hn9n+vVBhphEKlTf4VWgBeO+r59D+BtA3UosjjXmEU5JhdGlltPLQnpH
Os4/H4d1/Gu84jMTLhlru+MwUZaAs+P61B4LivPzcbjoanv6qL2BOcKGPHf+N++4
RWGi7iN6oqM886fEu0eZMv4lYj8Xsl/pB8Q5pcKdAYo1fRl3hYlVl2rdYoO/15OI
YS7LheGMo71zGgKh15TBXB9am0PqZcmI2DxnqOUqNeL5FuWNxx01rdyEFpY+egyU
s2zDeWb0t5dgg+jUZNxqS99UewoCjFBEdJJm8BzboXV6TOsS3Uhc9RN+HBY88J0C
cwhELEEo5H+iQ/8ebF0GMoMIlH+1bmguBm40zU2X80ZJHn246Kty7C8ds+C8i36U
h6PnuT5reBuyoa+I2BvoB0462HG9J77hTGUNFR/E2URu/vqbF4ye6hYvnkXpySwD
9oOzm1v1vtg9j7klFKugEgrFaCWUb2neZ5L6DqUg6LSclsreu3mdu4a2za+E8KIK
LX51aY+/JGojoyHRxgDdLDJKZfqikzWkTe3M8xx5iFlaCDc2Sa0xNUNwSjLh9U2c
+ovtyQFG13NeYxF2/fT3wTIQP2yjNYhomUBqBpbtybNwiRgizFsdRgBfCsVzFf3G
Relr+7BYuyjeH7VahHJJJ5qTPI2W1kHAtb/ox4ae86E2j2MbB7s+YcTgU+BXrrzF
chQCivoqNbEq5B3rR/li5VqDi6lw3g6skdfIF1/1gBJCvmap4RMnodUuUxWnWsmW
0+sMF2A51ooM40iCY/FeNngwIhzEeYG2vuWOcw9FYRO5rzSLmRswymtCx6PC0ede
hauJMy1zBpNniGgQg6fmSj76MH24YjrXkiQtHIa8dJNixCF4V2ymsYPx9IVkLBy+
iS3ijL2xEi2Qfq3FJrKXsl+skAeRAohr7i34cBwHi0A1eP1dv5Q9ovzcPBTG9K4m
4yUh+VT6mJXBSkMAD3aDYgF+vmPKRBPwUbDDlSeki0z2Z6Wrxhv3ngi1hyWkJ3OS
fvUGlVVXb02zmsd2KIHYvj9ckmxig+OfNI937grpv41VbaphsbgoUF0u1rIg8UYD
vh4aENH2z83ssRsVF69l7758FQVXBALrTvChmQKm4zC3+YOsGQnkiED6rCNNU8Bm
DwFvmuftEqmxneA+VqyXIz+jZKTalf22404owPJxwZC3z56P6ir9HhQ9sozArAf5
6lPu4W3bk3lMHZ6Lqpbp2mFI7Gu81iAYcb+AiB50f7pQrH6Kq0QHdS29Hudik/d1
kI0El1AiZbXBkMsfaOH0XwSeZXKZ6EKWf26g3ojRFcdPjiZ6HuDKNE8XRq5NNm5N
6zsZgUwOIo1/s8DZ7BecrxJm5nWOcD8nzfBIDK7SZU7P6B0s8XK4teK3c/ESoTxw
0VBT+BI6R1RnrzhbK26gxhOaskszLGOzrBK7thDjhE0GX2imu0rSHsjlqGfl2Xvq
85pIf1O6Set82F2LwjTd0y6fvO/PWqNJa95fqdwpVixkTqWDrOx/wMzhHUDrmwqD
sOoftNzGQlwV4Lkj9LiwDfd8mIjQLUbNl7Axt01BdSx2DdE1NI8V6V9AQWqP4KuZ
+DIGRMJiU9CLNrK1Sd4dPKAq9mvevC7cxJcPx9Xtf6zXYg2DVUIFnekhZdaqI305
c+C6kEowWviGWZhICbGUW16eCXgcsu921jGV3b3PDEkcrOqzw9RD2XC8po2ZYVZh
U68x8X2fCwjv4h2hL9mT5D0pcNWW+xRsOxjLEftzvzV1PLiQjrrXWUe5ez8N8g6z
hQ/aGW3dvdRPmjp6RDnXk6O9B9i3M0NkapnwHln9907N+P+W0oRIgDXiK6rCeWLL
+hnnIyQ6RAhLFRwXnK6228sfVXp7hJh1kLcHCwwAvimoNXBkJ0Mh271zmfrphhed
CfqUuIQRhiK+BHgV1GNwv45bhk72yBYhaHMA6+K8c3GT/2b3bfwUTwyn2laNW+Ij
bWTl6p8Cd1b+pxpwRaHOeBXLz6ELIVFSL1JDh7Cq+MWs8yjkh9RNxNk9dIEVbRY/
eJhUYl4u1FnPCIzKvHwoxKmGjcco4Bs4wMQ3+tJU2bHyz1tfzvFk/JADs2fnByPO
uTFdrxspZ7pMNUMHQdP/WdgrTN5sMxw068PimRQE6xNZ07mr5zowfXyLaxec9j9P
+mqLcomVJoOTO2Cf2Ow6xJ1gVBuw0ee8LPDe0SK7cXnEZlfYKiFuPLfNXwbkYPEh
nPi6nUAcCV3Q0xOWojquvibH7VLkiL2rNPMRkMrhmq495aRYjL5nUYUIW56Rlgts
WftJnxATGyJEHe9sNUW9z4reKLmlDI+xlmYcigpWItZnGR9Ct5OZVTAuSnI3As5i
mNdJSSvLbznUlVunwoiAAdRxOqEWnLJGhg4UyzFHvy/xcjWxhT25L2Xag2HQiR8L
ra+R2a70QbxDjmNX3NQni9CsHgFuiSf4qp066hXbktrjXOVvclGQjYOIuYpRjOee
XbUOon47ayAFrilpYlqWqO2FnBqnnTRqwBll5GxZMthAi1IWeQ0KfseTmve7hIoc
3YS7xbbncrobKCAE9EM7RB4SWi5VsZ9Ss1w5bp/FDE52mJKWDFwZV4Ry8EbqybCL
u4MxJDKZbXy0tgE68tY12bGwDb4EFZXQz4X9/k4x0Ksw59iizhn8J88RhGrQCopE
7k34Mq6AqUz/UTVVGYzW7G2oo/FUKKYYtEfBAXl72qX/ol7f3qbkVIOY4bxofsg3
OM4kFThM1hpk5AkN/DlvwLSTdoCSjXas+Qt7WIpygli+IOs2LZcb64Cls6ixVLu+
TbtqjhP6IGCj+VrgIUBsWam3fTQOI+B5bsBPwTkLL3j63Y1VLHNupmY9JJEHH5UQ
wBNbtabU+zxAdJ9RML+W1lOY5SFYSHHncjkKe2JntcllnaSPMyMXgIeiBCGRkLGu
IRagMWqWriT4Z5PGw8nHkIFxLsTrztl20mzuC15E2QN7fSrt209PRb5RyLQfIJqc
TxceTMwdUlHPgKABeUJCxVWQmL+reTmj9DhwsYVDXUutgdLosJm4FsqCnd3kw9IU
d3yShtdF0a+EpNZiUboqB7vID/Wj7V0Z/g7QBYeYUrC6Mt79JrYs8j1u1x4zDOjC
X8D43JHSd8QTDpT3sWo4ck3LI/rjZhVmmjHZq0hA5tSa1r1YEWqwnSx6D+UK78u6
r1PzVHt8tOgYxniEuCwUdOW8eLS7Us2NI1Cqwfvk+Tgrr0gFsLJ7J5WY4JD6gmuH
gttbsvavQke8244V/L0MO+m6fHR0wJOZw+7UDaDPPXf83JL+y9eiE5hgEBET/N7R
HgivgkyFD36yncPWqyhacWHKazyoNp5XXuo8A900a+9GXOoAXmXdRpsEoLmAiEga
UH5B9iKoOSGl2dosdylgvq+tChtkSq1StVRBCaVAax49Bxy9qEe12zPfj8lZaSdE
hCzNda5noOmVbyiovSkKmp1+1si/4J14QYIwXiUzFjxrBs7cF1iCAfL9BkWQQuxd
t/8U/5KFHZG7icwTcwr6Jw5NyCnrpfpY7Yq/o0Z3xDGAhuNYKZPDf0IJ9DVqCfG1
g4Ns4S6DOFY9NP/0gWRWiHC3heku3DV2u05dvcW3cZ1MgRAWyjYd1FYJxgcfsAGF
AuBFj7faox4g50BE7XVO1BdsDs3x4HOtp7RTh7iO2hEl3erCztJ24DHOUA2y0Ph8
/mepWiCuzIjrVjDDucKnc9oSonrsH/wRPjDMRExr/Ffd0HJv+HdIJa59TWWknYyp
VWIJZ8Zk6TReKwrOf5wXkq3kj3NRSre/hJv5aAJwV+G6F1PYX9iXgG+CZDwhM6bN
5DhfwVNOoTBZ5ruZkikIWV7nmGlaL9yL8/SDyQtMmEbMKobfwaoF3yclv242F8+K
rIdq2zPl1vj10aeUJBNMF6Uagpl6gzK8FlmZs60aO/bFFLNhecZEgcN0dN4SqOsQ
ZWchpeZpWo02WEZHDxWlX2sLcL/Mqul7DVt0doB5i0pGTTYZPf9dV+WQMNSn48lu
V+nSfkFuyMyqnPKdZzzKRuh8A7GHz/xlVagdO+s3VQEe/TaC2VrC+YFSSlE0UQ7K
YF9dlrT8bHcHFN/ntMfFZomjieEdMR2SegV0JFJzGTBfy2EuZrZ+ceoQt2e8lTxh
2bzaSWPdK85lD27oA155bPlz8YU4jKkNB8DfC18HzBfwjWe+vUsYFpQmgVgt+7vo
FaKhBSY1rgQsXZaZsyoZZ4AhjqpeNWIji3tOMrm15UcPHltk2E74QrchxOmR9MDx
hGW1LPDEvLqTwXz0HqpU51TVXpPwfOEbU5mv2F7GNVQhA1PLIEHN6A6mS0C0R3Ad
r3iJVuvfVBS4m1Ma83EnIg9y9SRIJoR/EF0d7TBEfOf1vxKGD+FNYv2eQb+/PXFy
/7n5FfhQmolYsov6OmJuPkn2mmHs4zsFTLBk4HDYR6VlheDBv/hH05PUj4IRnLVl
GrrwSp0iGDlR+5nFuAXShsieDZIIc5S7csNQiWKPGppKgmJRLO3Puj6OC6R3egL6
plariMkAmOaI4XcBFoDURamdGUb294YOGBXQR6XbzOGiz00caK1heqd4QFn/0HyJ
B49Uc7U6VwTF23d7FQlTCYFdfE+91z80btqTq4tHGyat+TzkkKzd6q+VzZdCL7Z2
IV8CHMl7iKoeRusRwCl5KoBisu/WxurPRSew6XpLoxrYBYIcZpAjcY0DSGbTFx6M
oCjusDOh0ww9JiznzLawFxh990S2V9D5vgIQx+MBn1alRmtky7TI/VY9nwFW69//
hnP5V8CpOSOTV3hWjQY0OOm8vNjfvVXRwzx4vWHV9VBJK3ARU1L0/GC/QrKcruXP
UUu5L4Rb6fJjBAjLeoX5ixEHD3yjk2gMURNIczQH6oCRDiGopMRLDkSj7LmM/7R3
pZBGk4bvdwcItVnMc7ww9S/8iKyrdFNtQcSP+R5TIk5XTC8lHHMG6pYYNLOjZjyG
vHcW0pjjS2pkLEExskuIjvZft8UTxaEaTZTrslfRg4xVrLvucxuMULcn+YIlby6q
tWskDFxzP5gCarDEj7o7dO6FitZSLlwgsdX9VLkRD0q8H0iTUbuls70pTWHg8jvX
EvoHqDZgUdTaGEpLv2WC1wpZmpAJ+Y5IkpMbZCNF+j7z3B+3W/drmUAo5QhvKNfl
c6Ly76faavinp+H6PeUK7gMowcOL2uRMapwWT4rFk6fHmR2ZqRECMBUsNvHoEOJG
o3IkrPt7FLsVt336e13Bo1sf3KqRXhT9pBlh2dr9xUYcGzkiW6QKCcyS3rg2t74g
lL9NSrHZJtmxQltYpVtMvwdp/QShzFW5SCgrN1mFFboda9UVmGPT+ygQXgbWaHMT
1SNC33jRrQGOuRrwmqzMsZoE2tEUS4sNrQY55u21ufEtUnEqjKB3ReJsBUsWVTUh
idOQfMpxc6qqNNbMLEk4JSwn5Iy8cFTw/YcGrJKVXIRoxLXLpu6w11THRjWCXfYz
Uz+Gy9V0aT73kwJGHOnBTOla9WoHi0BUYMn68CVpQiupWD4MFnytlrlItLV+Fot/
o5EDpsQGxN+vWnCju6El7yzcIwm/aS3ZuBS8pA6Shmfc9iFGIbtK0DQjeR9RrgIk
brWHI82FDbV26aFpFFwfe9KkQ6O6vbjgVLY3D3znmEtxwQv0d76/7N0lUCnOneRI
uWsvBeVCKYWKv6yIgNDcXmFCUNtYjQwRGj6W0OFOWZH+drPkNRcDqKgd01uPo5Eb
yD+SPsIIis8Y+g6IG9LKxPxiOzMASq7HuPun+JkYupgX3vtSDc6zx2IQv51JM2Xm
0zNWyLZ4JGXj3tNiB8x0pCOOkGq1ahDp3JImm0ZTeWdZGMPpm1lOWiR11HBtY3U4
L4lmy/8uY0hyiAe9MXTvDNQXDOfYB1Q/c8iusP4fyOjLR4Ea4WPwUNoG5gdI8W2w
0bqatLJcUPvxLawJ54w+dUBI8aQ5gxUOOSF8cS+n13NiBLZZ4JvE4QpIMpc00ajr
biUyJOnjjjWVCh2s2XT2zggVATF7Icp6aEZzuFqzU3NtRQ9H+eoztWQT96iXkh6b
clQRLZNXbMrJwdsJIXNNXr9bhUnGMpIgny8/KNGHTpIXDGGpEc579CoFdHOywZ5M
K0Dw/HwR091GVbXIW0wGvfxbJIpRzqJLD8uUBlpBxsDSiWxWj6eLnzyvWg4DxZTq
VaJ4ssHvp53kvhWPlhbppOD8kTtloi1LMrEVZjfBNerwzg5TbM6unIVyc5eg6xdh
nUpc0khUAF4wWqAn9Z5qukbdUKVBkAeyHVi/f6lpjDf3XMDGCbmVqgCe4TAseBb+
QB4xMBlu1WhYhIKBqxteefAFonlaNWG4RuypC7HL9l3GyhumbI4caW27eLJXgJMZ
HtovAPvLblMLNeRwBJfEzKFAQKcUuQiaXSz5fL193/7aajvL4ZyBKxe2yEQGS86z
Gyelzo0+FAQpil2vesdBPCqeNXoESz8sAjpLgHGc808UAjRvIXV8GUThVL5czoED
iVdu7vtftORtzIr+BzO98DyRls3o6YwpXeaVxAjz3wWYW8d0u0KbmhGBXowwQw4+
hKC0WbrCTQo3s3rDHempmJFgCsfhwq9uVY27FOR1BF/rec2sKxPtBO4tN9BTtDWE
LwH7H6NlGCuWo45i0+wB9drjByM7Nr8Fu8e6zDEI/2RM4Nq5sTEiM5NSJFOGLP2v
q7HhB3GIeBS4obCS7tJSYIWxO07uqEbNU9a0O55mTMgiU/qYwLgDdlyQxzeLalnC
Q8yaDWJ6ccsp+eYsP3fTaVjmIc6Y9HZevWSjb45IPM8+kH/XiCJVgD7pmpDCOAbO
1Nxu2MtKpPTN14f3ux4WTZQGOeOuppSYqd+slAUdAqG8kHaUV33aRniS4hYf/LuX
0JQdWOO8y4IhMftsNAAGOl0si4E5d6Sv2crzMLdgxnQtxP3m2zfX9HwEMx+pEq9X
ZnUFz7cFwRbtTquqISoUZC5elIGz+wjKVHeougkg81aMr6hM2HjNQrcB41Yf8fqt
uHCMYrZLvgFOMlaC80nlSuU8sAoNklaffUj4y08BwtuuWSBAjG/1WeQjUrfjtzB1
JcAcRApB7Yjch+IGlfLZEzK6Qv0uC7bDINhRz4c7ewr1YPoO4nue1QZFS6JL8BaA
qQAZnCiVKJz/csSf2HqBGWIa3AvnY0LcJXGl/AY2etrX4MiK+KSsjpr0kUZhJLQX
GYGdAhJiKxtz5Jd3vnrY2FlBtI12W5n0yvwEGZOr9ZKiErZ8kMHy001ivtQ/UurC
uF4muRYebjo3jNs6cWGS25rDspYZYJ9phloNxrcWwZrc60Qg1KsddA9UOQFEtTkN
qmLRuU9wUWqNQ3bsJVAH+1RPslMa/J7zzmw3SPqeL8HG4/GU/njZzGdw0u/b/Ret
zDjl5SgdA7rS0njEZuzeJkdtWGACEkN380Z69xwAPnhhySwMNDMPfAcxmlCzn6Yj
0cKQ8JjHUtWyJLlmPFWGcx3APqHdkmqr7q6Rku64q2+d0kDRpLb1UOlGu1N1a0Nf
vkRUCzli/iUgXs5AnkrwE/UZlQRT7mb760dECtlQGbacR8ERxjTBl6vJUTaapzlT
/QygObHPHxpX1o2opPyGjZzhS8KW6rRPjq4z/bweNNyByZUVtYuyXWEY5DAsE3kT
r060s4glLDN9kAZWzX7iVNuJEG9aGBNFXtkNCtq0Qy/jfGWzugoovzJrk23iBqr7
W2CbRi8tRAJmEMuV7//Xm60yj0jxNRKB8lzvg6h8w9lgHsu3L7/tLlMlJSb+Q0Y8
bw16D8hJzT37PHRLUj4nwWFSevNkaeZrCNmWHWbavfU94IHy4D4O4taTwoGa5wKE
4D+cO8poRf6Kx8NxQ7+Ej4HED/MulgnhfWxYEA+4Xwb3BCbfO1aNDR0QkkwyZlJf
nAxoMRthJqbtLu4GW/0/m9FFSNnp7NkCCA/9rt5LR/cS9cCbk988lzwWPM6hu+jR
2B0rJNaWT6l3ke9+r/V0QLGheAAQL9GGXkGQt08GMKgtl/9I1tq5JpJeWM6Uv1sG
1saJ6HjzzQ/c7yx82q3rXFFvo6AzbXt4j9D2nUJsXD3TkHhbxgEVLFFqbetM+mja
x1fogeBnqPjs5VoJVxxKohCc2QLRJcmTAmsewDQkc59TO8zyJ70UdA0lJJ1x9Qa0
xzclwOKIlyAJIdIRWMz808dGs2710zDNkfWCR3ugd0rHZhMFDb+sD6NSO1oCwfc1
Lo0q0pYTg6a20CGINqCeuqqi1KNdM33GrNAM0BHGsZjO/7CARPooY4oQnHpMBnob
zXa0p0ZB104s45d+tiH+AVDHuTP/qPXM8u9Mdh4dHXvAXD6qec8CKj1LJPYeN7Ta
OKt+Cupoxuwi4kbSuhbeP2yJHOq+9XaUem6eT/EESVzRu11VcMrk6EhzJs4bg3dh
xjBLxZaT6iO9aZYM62/mby9mkfMKdodCELlUsoUd7dn0M+jhaO4nY/sROgkWOQXy
jf4Hk4oLDVMrcB4h8b3MXTyggGRSmM0MpuR0mpPJbu9mRyO5JMw8KuP0GQg84CCA
fdCk2hHZ8oyCprIWvFVYGK6KMLndpofQwcd8awE5trJcGaQTDOgCJJaGRNhmmmFw
fLj7+fSp+d/4l3GJU8dhtS1W4rIRyzFk9/4mI73SpmMXHcJt5eizbNwPNppTbIQS
IV6mCLmJVPG7LzheQVwLexnGvf+Q1dwa7c3xZX282RPWEdBVLVOp94GAyITXydgh
qC05r9Zzd8WPOX0cRq3t9yA51l6mGwCH0jUgN9yUv2I/+71+NsU/DjuwLAsumhOA
PsXzL7yML5zliOhEgZTeCT81McIV/j+BarP231cie4uqHqtyGlAwHX/T27lE/1ZK
hCUcnvDC+3qeAKBDdHDwjFZyponV/sWpeINzg2OgZbwhTASBOciPeXtJwej6r0O7
viDmvOCROMOxXZ5KwLqoJrVScHbuxns6BxDnMV/9X1w/+ZPNVruNdjaB7NH/dF6n
kmzcroGx1UvUP1N25EyT8uMBE+SCf3tRN/t3gdDH4d8AxB5ifrsM2awC18k6giVV
upRp5QikYfuotzuGB0VYUXr3zgC9sst7MLCq+XJhn5qSEv8X82gKZB/NUd7nHya4
UwacxbU3uCAnFpGx32ikP6Q6l2JwrL7154aWfA4NYx7SxZ91MBaav+EVbZ3XNN6x
CdDv2MA8FyKAH4IaN1wh49Ptv1NoUjddMgUmMbtwf69FK4LTFp05TCAJ6jDwzf+3
xa1wmVwItSp4jof4wp5lYym4GQiLmYqAImJlAULXUw6M10NxQgOUJ/TMRwMQLTKP
YQJ04LdurjOPN8ynDrR3kuLwVNeKu4kkn6lXRkeMgzi0/rnfgqEcupay32POi7DB
+Juso2+aGuxQxPW5PsezCPNo9y8mTIwzz37G/Kf2NWRce52ul7CxQFW1QL55hs4w
R0fzmj6+CT21/ikZY8LGF8FySkCuBsB8nBuWhQDBsgPrDC8lu4GNXtT/KAN/OTI5
bRWrHbLCvAfGR5VvUuMddXr4AV4Pv1nBHfiTbu01tm0J5uj4KkVWkSjw3pxZweBE
th/S9/xUDnWpdvtz0wTfmID/RPsuOOLSZl88v0zkIaejlmhqhnGnA/1/nB6CXdLj
r+H2IYa4xxWafGni2llQimwz582pGHN8nWd1BM9WAdJ0pKtYDDtspqK9EI207Ny3
8o4lqQjx0WUf1nXewbZ1jt5zr0xqvjWb115lxqsTHmQw8J/ofKoS+jRS8Blx8B/A
z8klBUW2Av3Z96GwZs9W8EGymPKvbJXayjMiG5wT+3J/HJytSDPkWbBFrNlghLRK
YgFb3h/kIVoMepK8+ShvXLI5Wk9Hk2GMMoKYrok/1VMk49twKA62MrDPuB356mr0
W15GhBbbFXXWwqkksi6c73tcGe3JlhFWPAdQpMxeq32/NpNObqtP4NjV4dZf2ufh
deTU8HOjhTsS4qIC4lp9EsXARlnsImhJBV6X2C1Cm4BPxtCCE0U6vohr0jLigisk
JRCM+XHBFWXIbQEiX0u2MO3lxTTJIz93UidP2L82M+sW4SFIGDlYcGErw6YbuZB/
VV1znoGg9X9Mo064NykQbr2aJfeYTkvhH1JeX1JieV47xSbXeGqoKBIxdsBoK6YD
wjuDkY06TOMiKqq2uGbx0jYScij4BQGCOPS0RVh0yzPbp1x2Ih8OPnky0wqD6itW
H0TvjMgN6mysb9PWHMju47qc+zrWgh97MwLCefLzj3aHCeyo/JYBgxtPxM/i4E9M
GNGsf4NwOB15WiqhDRgq/qUFCsznxe+5Qr4wX8ZFYKFFBLw9eHpkRjdwVUlObNxC
UZBheJbOuED7otBgjnsOtubMqCAlsriKBAX9Eqz95mgi5JLiXtvBIM24NY6V7P/H
uV0uFo6ohSwTyIZgKN7G6iPESLBgx7itoOfYDMQrymfmmEDwOdquB3+Uk9Gytzep
rXa0OURDZl+uS+qA/gNKcQnR91QSUh+jlgjnRjOZ9eoVEkSqiNRdpfBc41dr3g2M
fWBiLXqztzDfMJ0idJ8pjK42It250uPL3fZP+SNpDKg3ZB/Htqcl3fH2g6Oalrck
dWLmgEOKUZGbEStWlYx4tAfD8BEdzy7aARqnrHfA9ICNL6oHQWpiEtDviDWKPIHA
pMCJx/cZZSaZT04TARPGtqSdfOaQP68UxK8oRwLJutsIm1yRVqWBGAoIV1Bxlt84
zq324lj28i293WvBYVXQqMPDmZPlood6aLVKyk22RAplKyDO4Z1aWWcZZ7bE2TKq
7aSLIVrOfb7mWZLtWgfN5BL1we3F9Qcdt9GlrmWmL91YnTlnChB0WQBSkbao9aOw
eZEkPsfioYY0WugOEodVNNLTdoKikY5ksGcEKOElu0uipIL33lZI9LPxWf3+CyaI
1xYaIdIpSho1/P2dVglqKBNXw+Vodg/Y2KCr6momHW7fciXD4UZjhSRpHXj15tyP
NBBxIqRpEFhQc2DT2YYhXK7JDG1o9n81FUOBua6x4JKNpxVqCYwidS51W7Qb+SDX
D/BCkWicgOmmSM0PDHcC6gAhq/TFiy44TnZ1JVDTJ51X4yLItmsYP02M/CXn5hxC
aAiUyGy1Uhb0fliFsDi32WrLldLm13H6bX7x3quJ1EuO95zzDiwmH3Y1mbkC5WTF
hHrcu6wLjIax1aYLaCyZLU15Ndh5sydzTHrmL1R5qg4v6P09WaOCRJFGlWNNQZw1
u6oPjmGJYXWDfA1IOoV+Dx5k8vCGhTmiSIhlOQQPl6Ilr4M6pLO5cZiaeIOaxABD
Nexmh1+DxfpPFYZJsTWRpcgxy4I8HgMYmsxd5jr0RLfpgdYst6ahPYzBnFRnQgDV
9AwqmWepd0uS9FrFQ5VyeUt6Ll/89VdiOMqSSWTHgEOqX92MWxKJ0V/W90HrItx/
ao6uo/IANJV0+De1d7DZOD+vTmvYwnQX1t6iBbE7WzHJGIx7L5tc0w/A8qJ5aWS2
RhUJGUKO6v7EouTrPraWFAgRJO7BrOJpj7C7nLYOmijJgEuX87zmeOzFWS+ABrMH
9fnRpHOtnApsaZdgrKI9rt84o3Pb+e4l37T0e+gzt4v7gZhbJZ6R2bRycfNk35tp
coK9vVXrw06POfKJcE9QC/otRHwR39zMUz6uTx6y1CqAO+uHymTjRVpqCnLfx+4q
eJjmkkAYxwmGWFheXGDlHgJ5+Du4P7zqa9ofuJMwnhvm5waj5Cb6Gd505lqaUi0w
Fj2maY4w7juhEfXG5Dijt6Zn8FwWFL6AU8wO9ggkOh/Z/4TTgvAHjgYrsHVIvFBs
3E1HBZcpKt0H7Xsf4DflwT01uAI0UjXDZuyfRqL35KthBjh2To8Dhy9kxdJhNL1J
g6i+W/tHXavX++cIEPbyV6/JewE/TLmSbpZfmWvg55/d+ttftXhEprAUy3NiIFxR
iNJ/iAk62+jED/H7ooIVOwSUR5pKHoOnaqaB5PHIeVQkKWkcg701diLde0TU7m2m
pIYhli7TXOEvhof3UP+f50KfFBBvev84npbTp3LPsn/XABn0mYr16731SjykjTKi
J45qNzOiZ59opZoxYKn9tAEJ1EgPtsoiDKjKi24JEXxh++yYGitkvpAwSiFnSEGT
PS8ewDxPopwNEDUWko76NKZpoHRpnuNbcNG/69JDMUyb3vJoVQoVqlKeJTNZI1Wo
0P0Ek/yz+vkFPnAJbiUttOYLuBZQYcWE0jtsUy5u+xAwy9tZVwlpI38paXEPOQ5X
ev8my3PdUIzMkzvrqOEMznBjwBAjn7bA8HLhGVRjkNpPRU8OQ99t2wKp+2EOXdff
KYMRKvG4QNRJK4Ql+oUoauAQVx3HfQeHlkv8foHux0QH5hAWw2evyjDr2nHgOpfh
l3FzXl55wzcMotI2aH8lDN9KwCeYPo99Cb4usVRSZR+X+06UC2FZ6plIOlVndWBE
ykxuOClEgS9sjXNGorndOSAQ/AT9GAc9X5t/AlJbDUG0yOQsG/P1NVS6ABrEJCUq
SD4P9tcHWxeL9AjIjWQR2onjFAO6+L3KJ6bC65psR69JrE3VQ9G7y+9hdG63J14T
W9Kng/PDtRB8cYjIiqjuG6Di4FHsjXB9oAyKRuHXw3Vaqt7e5oEJ1dF7xHNBvMze
t/AwkCPxrQujfg3Xj1e0X3tIWu0m0uZBFl6oLmohuoI1FObrFBRJn6qI/Q8SIY9J
3xronjP4DNZ1fzCTnTC+MvyQfbK0mXZU7DlbmaelMXQu1i3mjVcWqPvgwWjITGIW
DEM/aOsT3AI1OR1Lq4QWirpFleuW6lpMynqSlofkxvZvV6rE7gyn1SV55WvV8QRD
teEMUb2UB+XIx9R6dKaXfER84oMp4letJxgeNrwkaiDrBB6TpjTXxbhpOi3+OZqs
YmA/XTGSe4aKMK++FHNLrcmwrQAQMNHvCLLgJIc/ltkjCedEaNeCnHn/bI3lt6LU
WU7/ebbYkDgUbx6Jhjui9/6q/ny6FjdCtYIyvKrNV8bhJNsYkjkDPfVUMTxfGVhq
c0UnwqTbBt2PFBntQrjMZjowmzo5xZGDhmUjrmiUdoBDVRrijNkUd0zVctAbl9U4
k6HmC9PYpkcMJHp1NdjATT68S10+gmL43u7uK8Eb4hLEnzX2tQ/HxMifvrztd+D0
el0DmcjtIrcMVylPPW44e4CV9VUQ8N4zuqrbpBmhoF7C0afWdjwxCcv2i1O6wWyV
ZpIZCU2eX/cbRy7m6mx3W9mDKbAwSSR5J6o1DFf3nCP7EvztEyMXWtqitb4cs6oo
mLCPRJHl1JrNjfXkNnGNQ7mK6J5ACKXIBEFmwC9zmsRzLCLdP3nY/6N7hU9t62Cu
To3rrMVpDk5s0XcqhC2Z3pV1dE5upUIIXQdhqJGkPMAnT4bwO5u9WKjo530RmcTt
1FzbdksNzoj3bP96rT6ywB5Xjmim+qZChySHVsvTz53/k7/GrReRt+6zLgOVQ49V
GqaH+f/Z7SL76AwPyvD9Hj5bJ5763zqE59zlbHRgn+qKRmDjZUUZc6Iz2Dqugur7
e2aPcfCNSLNJ04HH9QekhFLdW8/J7G8NriZikSI9wR/bIsYkGUIt4Q4u4TVgTUTH
kl+aA/rN/Da9Zv6P7QCgZmf5SS5NaiNivc9jLlhJsGdo0F1t7gUHr5UGRc0ggFB3
jtoScMTpbamP1wmLU48apbnbamvcN+3zFBx4XeMnlKKRxQJ5CpukNGFTvAhddBay
kfJ4KLmL4QwaAD2t3Zuw7ggfc49YSEXBKIR+tB+Du7dK9P+nz/Ybrbs+a2L11MSV
Y35wqqWV8Np2E+X/0FW+IihVuiHXexXQ0W4nGJgdpk7gymC0uTnMzEvnQHkO5sQd
xxXJdyz2MJWJaBnolfeEGni5HyRWKPFWaVCy8UxzjSu7iHIoQnmi9jFFpziG7UcE
Ilz8PVkSxwzEp0L/aJDq78pOZDahF8n3f/F22X1moLsvgerw1F4Qer+gPrEoT9p8
eb9Fm2IdbvWVc2PaJCawBLk/Gk3WsSFpD8U0UWEoveZHDFUiJ5jkvEOaPcAci6D1
zoflyqk83Lu5QarRImltpy0fFIM0uW3tapmKHbQI0w32f+wFT8zVZmYWRWZUg9FF
kzEJiU8pkjTOXF5QQXdtxUmoLsc7WNKIk3Ke2N1VFs3lNhGPow7xnf/Pr9CUC8Qw
JribneBxYNjCm/fCLiAjI5+AfsqxjZZ0RYyVc1KwYuwNJl5y8Yrt1Sk55qi6kgBf
PJcU8rk2/7vqrQDMegAedo8Rd4pxsuFhRLUkfhmeGqO+tgo8ly0NpBN/pueXq/LG
/79wGYAxCqB06XSJACMLH7BF9MzxbzRD/PRI9m7jsb4K/jusOsB+0Hu2lV+oaCwr
/6Mxm5B05oVwM+vfjuI2Hoi5lPiuIq2oX72FlPLpX1sS4i6gDwNafAq1cmf2bQBV
8Kz0z8fRiTIHch+xZLZRp3lWaFwEz7Id1l6saKpgIuNCOKcVDwfDQjLdAbHiR/YZ
JfWQP0ZfszBQZUoZdew2NhctznEaciPxPSXep+Q3UxjqdYbm60OEfK+8yRWdi0Xq
cVMCbADNiEKO5uCdRQYKxm8zofwwbq01H8bo40Q3EvYE1t6RO592qh3fbt5JOQx+
YTqOIKDNJwwxlJH9Ep9nlbrrdmPYNihPAg0kuc6VsDWMvoGDUm2tWpO3OdSaZeah
r6gw0+IgFm0rGL4tEAOVio+tWaFbPYep+hPt1BYzZPzcFzjs8Z8DTpzqj8AcQ96+
i4dA0H4zSpwSyemvMPwl1iMSflVyDaYzUw71kqaxVrCpjwqSx1iPBS7QDYnn6pmD
6wrotb/Ws4uKkpr6asaRsXBXuwEEoWdw6l8AXGzlcbYvLSlkn8uW/XVLDnFxoC7I
s3nuOJc4R3oUaOlQPPYRPgAjQz6y9W2dZN9INmCUj9DXhwM/cXkM/cuKPa17GaBo
LCr00Kt0dHFlemTP5I6ErbiYr4VTo05I4iHom3ZC8Sh3tAN6m5yeE5GfYHfHZ5Sj
mBEa0rejsvPYNFyndp0pnFXt5PQUZrQP3zRjclsETOk71ggQGkaZmLmqN4Sren24
U8Fx7qK88uMGLpKGBkVcROVkaxXBOzQVLFMrRtBxHlCNSinXDob1ZzXV9dSL8cjH
d6A2i3gU+5Kuxrq4JISre2mj35ZzSnRPha5MND+D1ybGO9D49iF4PdGlPffhfBRA
I++KENu8QcTB/FqAz01+4qx4U1j0QV40yRiEFhxNlSmniQteCQOyAwOnAKNz3IrK
KpHyD6bjlW2rEtJItEj6rAkhW1BezmneZuXA16DS6mnLNR0099+60rohnP69AxDF
qddMdO+/w6i/NKCYD7Sx4mymVn6cn+n2DuaGh5Brpxvw/gh7WDv4E1KSMq7w3DNz
7xdTY09NI+qfGPPp6xLAKB8f6hitqzWSX4pkL70Be080zjQTfQR9i21w/os2zIY1
Jwswt/9zXGA6kKGNw2xtVEetLcthKSL53ZdIEuGA7zVO4HPWtKl8oNsl2q4WLp56
N0FL+IkaSLHnY0VhisoOVHVFxr/Gm+at+TeTi/54lTUvwpwJoaH4F703mi9Nje8V
6b97KujhkXqtxBpgEcQLOfliLRCj1u1aJKjuqtkHrYtq356vewAV4z7SW++r93/k
a0MQQGnMYiMPPc64QLPYlg/lBqBKVFyBChd0t81QF3/hAzwjldbElwByXB2Iy9Mc
m/OTd/ddJhWGL/sJ2Q2HChWtiI33OWCSnTz7AE1GdUq/mVo2VZKW/oQtFRKL8D3S
VU1/mbmM7F7QILG7H2c0xipY2xXUoE0hnwMo4FSFr9TtKElH9dRw1eC4/4nTYyi5
tTVTKBQJdmKBiI0A+My9eOpvdLhCscUK2gd/O9LlKF5ssFgFTI8WPQxcKs1++WLV
5Qr28JtPKCgS6gnWy3AECeDvUTRpxGGoG/4X2LCJFUv/Yshoz9ikyeAdBoL3SvY4
sMzTFGiQzWoiJxwAHa731kE301AA+2jLmy2aupAGMinrHiiZx3JN3AF4LTtL7oXg
s+90zAEUa42+XMmCM8e+LQt0QwGywtQEW/1prSTk35IC9TTAzwYyqLyjqzq7/8F9
ZW+nGQ4MIfIVDcmscmpTPd2TKJ3FkSvuOtZmLJ4yd5kS8QAK8261bFXRmYpyty8L
I2J50nsb1l7fBVpqesBRMSFmHDllaL1COvU3tio75gRFsSxuxcIlNSdERq83Plhq
prBPvb2caPagw/pm37Iauk8PBvgr+GnBCQt1e3E2sPiAmY0GAwMq2sZyghZKmEFZ
q544ZQpj0W1gQB+8/rNgRfgSARmmuGeZr8gkMMeffdNk67oXdQPzsVWGYzO+HiTq
F31e+8Mgf2hol3ENsLehBRbME6v/RV/LS8OS2DuunZGDzMe8XnuIptQEtgepc5rl
E+2mbwh/uuf1n2ehqW/bP4/RCEmOxj8/poGNrIVwRyMDB752rP+izL/OrRuR+Fi5
UEkXWHHQYfkD0HWpAs5YihcM0X7aC32DUARnFUxGZRsXcyCJdn6Il1UMV/pWfk//
kFhqOJyiArqmj+59A12A7/PeXQ7lklbNR089t66q2H4cnbv4R2fIZe8iDTbzXgtG
HZDrLkIEkmxr0ARozPfFOpFEShtP3hh8o8lugLnzrKVQCDLIGO1lK8UCqt9aJkw5
EqJsF73k6B88oXjvMDbePosPGEA7LPX5JArO1KmdWt9uMs5ZxBVNzM0eJ5P817Y4
ePxuc/Z2uArUCUPvHK2YsaIO+lkVDaN6wTTbvctUzvBEU5v1e203IPWTMJdyEojx
Mr7xJMU38PonWltD8yyh0wk4buJtabxONhQ8Hb+ae7TW6bgTbFk8Vi6ofCUlbgos
t7SFl8QUN/enovJI+Lu7c9tiYaKKPPcklqUl8eSIJ9rw8lDoLbAo/RGE0yeP42us
Dy9h/grUPuHaAH5NpAX2Q7mpbFt1Z/2RdGz6L7RL26b4vZLof5+N9G7uOXoUvgl3
yb1kc/POS5UPfa8Qaia4piRYZxjuX1ZrXYAjfLeJDHZtV7y6mNyybPadHBhUwyCU
ZolquPttW99C/M7jlpgRZqptHV4t8HE5ihG+wzNotarbUXQNWdD9Nf1ZC6AjXtlw
MBKSa7lTMs7aTkxZS8YcWvioKeh3tuwrvXAm8UAmnDk8897wr5EhBeaDvL/hVmgh
WYRKEz1iqvfvmXQpEfiQvFjJahw5Hc+RBRwAA5wjGMjT959t1MUV8B+57BASB2Mo
/90rMqXQUCnZ4RMxgQrnEg0FFMwnYPqIt2a9A/U2alQSiJoeNM5w3/t9dWMsMBVJ
N0PXVh6dlVTuQj1FOYm2wkJvvqekYfWRC5iOiH/N59J1POZj2PqIb2+3Y4RqdrVt
aWbBIbFQYW7z9h+aaSl32DviTDK+vw+QclnmSyoiCbTQkIJXnlAHeBvCANc3/CW0
gLncAOdEKQZZBbS02s6BUK7FnTwagP67STb/0j4EpK9IsWgBKXvROnqtRVxKpRyO
c3tcq67T/OErgDLphnkNgNoFKsPpT+NBNOUnNLcAAtWq4EnXwCRnuu6DFCbV3hmt
cJg9h03LLGOcHwiKnLOrVMVvY6Avq5PQEKLwaUfn/rNc1SadoK3uC+xFNu3ygSpG
vODxeFGuJPsAXwZyzEvG/FhwYX8WlF1V98n67h5PgH8Ms284jcX6S3RSMFu0dd7R
Ko2UnNrgmaVf2fFnPYwqy4tNV+QS3NrOyBGWfv9sx6h7KJhp1xg085u7dM3qRzkE
bfzY8o51/Bx1HH5azod6hrsL1Ef9NVjHsnFHuWvWQmuSsphA/ivU1GXQsjELWhrJ
YwuC0zZ1slErAEVppPz/aMlHCPoNtl5shElKl+CXU1Fp4JNqxYBnR+fJ0fyHKyS8
qG82p8wPr+zsBYCExUxW8B8rxPPbPUnnkmDc4hB5wDQDxn2rLFjmUE4Akxuci+NU
zAMltPYWQmYmT3dwpkV4RA0clF9+Sn7IroSjWymUww1tzEcOC4qBprSRcHL0uZhw
0HbEtkFekBZ/9LdAddc/wan/A6jpqrhy8LFv62O+r29DoSTu/ye5X0txI64WsotO
dv1a8YOtsIWOBB9k2zA+8Rgb6zneH8Y2xmue6memjTi4wgiptSK5euz86pgA6it0
ZheEhucWT2JOJWXS08fjV/Hh+tBAKqOQI2DeQjHSpOlApbiLcZNS6gxsSqYZQHRF
Pi5zuYbcz7TB0IUP8KCdcZ9fFiXdEC7RRqYmu8fwkhs64ejQoTP/h3shwm5G3y4A
BqSW1YQQhVR50XV2enSKXh1gyeBX3wr7/UPxfsyTPf5Hoi3czLaD9RSA1KNq3CMK
3Dkyu4BWBa5FeNC249tulnYAcxTI5OdF4sn7/HAJD3sAyXGR7KtIlLMePjdkiO7F
nI2lEVwV7msfTpJhb69Yvp969jruvUL9pO6FzJLQ/Xx4YAq4bScg4M39s+eFaDQo
LNJazhavMcpeEETCfTnRDwoccoKBxBy8IwdL+cG79uQedJKR7q0jbxRKdajnOxex
YGftYu1dMJ/dSDEXJk+T1Ch3YuHFF2zNslZkTE21ybMqwYg/YlS02OsQ9EdMv8Dr
1CTAbqt7v8g8xhhp/4Lr/SaszrmuXMHmMIB6p09C8qXlJF5x+EumfR152zruPq0q
gym9h6rIrYUWP5fSmm37yHVUtKhTcKnq5jjAyYVQhaDYfVGKB0eqCVlv2tduogYI
N3IxbKFOCjbWyLdlNT97a5jGna4sDj592ew2j019f80SHG6kSQksrnOujPsCTBYM
cghBQMbXfxEVKJ64hUrk3RX7a2daiqfVIdpp/z10QZjrASuYK4TwYrPBuoeP/1MB
iwDdqkexHNDcSX0LlS2YdkljaWD2jz0b6oFhEOl9301SkYW2vURkNu5CrR8BdfgU
f/WEkHb9Bcx4d3/uG62BOdiyKatEK5xcB3sEdZICJL5eQke0AFqEfJArKxoKlUwR
KUWPOFUjqnoEb0vRuLwDZ/rI7ZYBh+Viyhav/78lkmvZFI7J7xQPm47ZWt2Qd0Za
m/cy+FVes437fPfFYe40pPGw+JlfcHgAgwishr1x/lr4emidGHZf+aYNdszfym7N
RvAD1hJy1gTVuAldpf6InS/0u0vdwwvYhB68dkiLX4pm/QgoZRx92BdH96aj09mo
T4VynSD/jK1xpJgO5J6tQE/Km+EDWxtlfuX2cWXS706Pg2yzHR1gH4bS4nXslXKe
yHZkVacHNXkbSokpAlwvbjDVDv/FDXP7XLTc4rUGD7QeyZKG3f0k1X9Nyc/0nFjz
4deehx2zQ5H9PrZIpREiVKb10zKHGtyn8cPgKVggDVL53ghgG4iKcYHVDBf0EN+/
XIPbDCIg01wwylLshLTypIwuBY/eLDAOqWUrMsYesaj6j38ONf/0HcLEwQPYn41k
HNYv4SV8bSw/SyFhLKPy1j6sOSpUtQjNq2Sq39BLAcytFMCRbwJ5JPNlunF97rPK
1kP6cCSOYFtTeggHxtooZQn0zz/8TWFZuoeYVlUphJPOLYvRoI6oR63Wb3dmoD8C
MH2lz3zUR5zOliAScKHjzGigQTGrkc4M/Gyo5lVfD+VPKKS8CWNn/UjV0HYR7H3C
QL3jOwrPocwWBsiea1tI0bb0I9ip4g+A2/T/dfRRtsuwXug6+TkGUPetErcVhMI0
WNZ7fQBI5OP0fCjhzGpc4kW2sdqXIgvyXs2jubbBqU23SIVp/okms71uLt5v6ZU+
K8I2MuC5zsnkfbsc9mV5SFDg+LcH7P8NGMH6Ssmtt0bUdiD0SV1HvdHeGVm/NER6
NvfRDqalGRD5x1qKB10sDs+PdijQHNhJMkA+tDswgpZ2vZSHg9xBLRcNZTj/GsFz
Oc0mctoYIdSOl6BINZp6Gfqz4rzrWdKoxQ3UadjbAfIR9aeGvNj2KmqVMhcTkGcO
5AHpDIBz/v+RTU2VuATkgUNEtysmZHmTd4fVdkh5wOXwNFFGA3cWDK5ERiWNTrlK
Ace2kYnZDJlWmUNEPXxf5WIrxRCCgLsWYXzTR9quJ57gkk2h7GvD/gg+PV2FNHh4
HO+RYt/zE8jOMUr0Im/j3Z0O3yan6/tnYlkthumb/bVQumzhlibQ8jp6+44SsRuJ
WXKSqjo5KPnoeuJ65DKcFooNXAgvzO1sRbK3SHHzwiHCrSPzynweTKfA35Nj3kSG
3JO2QdXCeCpGgtxCTF0kX0NKG7pKOL/oF+7DRoChkq3kASlFMxWzmZSbJt7PZo2F
w60ojQlwmP1utJFt22gP/IMFfm4US+576k/ewwoeeaVaq9Rsb1lzEQ5oBHPHhb9Y
RWLXq5tOm8X5M72tyzSrnAF/1qKG+CqvnAUAuS4BWpP3+0b+NPqfOnRXxODWvepD
ujhYOpb0mOWXVwIi8iap4RjEgTP9t4Qi72sPKI6KyPGoojC35K03PfEjeci9rnrG
T2m8dBmE0MVD4xU9LFIs+AX6njzsTrVzyc9CwA2xNxTO3hrePSTBOhVCMHFWjX0I
pf8NBS2fZVEtzSWuwXHtAszX79f2fK07qMqhObcC7swiaMJdKqCD202aulewi6Hc
E/RPxuDTS2TFAQ9gWxHR6AsB1saVS+wj9cI5r1juidT6XCPvatOEYNWBgl06Ptz7
7Y08RA+Of7gRE8ZnCCP1MPnmUK4Wv+sJllMd+yAMvDRCwyGCFNxfH/wD72IbOCbN
hznP+3XixWfZdw6VFUplPQQA97JaN7/HEsnxedKJ/OZknPb2Nnh7fnaxID+i3P3y
1FeO1nAkvpl+l4sRM+gNMlOAy69iypfIKoP+hg7lCpC0bpCt4z6GMyVWeJFlbjcR
a1kf8YEIbVQ+SKKnRR1PEQhn7fzMMv30ZK04IsXjWbCSCVNk6ZP3aVXc9O45Fs2w
cA6BUho6bn+99dQSgwgKtp7KXtaykQT24dZO1V7LDxSlAuFnQFMjG/vunQbsmfrD
dNgLvCj5qb7q4jxVOCTP/ijKbFJJkopxoqRM5n1pRkM4T0wHWUCOmuPiqiCJnHdP
QREYGAPGPdsphopTRgmwRzUcKAYRHZokHaZVPHko/wg+PXK1tGlzVoAhFWT2yB02
DLypVgx0mOO/oHmPXVGOIgCkNCGr7crvXZ87ubBBIcoBeil+hCXep4PfvPEYGMOt
gbyrLm22LnQMXWFBwPIbyj8Juq+eMcA3Gfuh2ryGbYVi9PnThHYH1hF4zSWmVojW
GXN0T5r+Ihz3rzb48qmBItn+r5IK32qsNuKTYem8WlmM3Gcn8nF9ysOXQWlkVbya
m8ar3sJeiWjUlIw8I6kuPN74laR9ulNPasfEyCWXEL7NxD5IIIR3/ZGmtx71cMWK
8borD5yz/54EOMw2cvGYOpsyukQOcyKJZRYaKtiwyDFsk2+s64qAg1rEjiQ1Zjwy
epf5Tkapupra3qf9ecC9q5HFge0V/sCmlVR+t52tixPp3jQHtBJNdfXrbQJ5PbuC
rs/H3rc2t5NN8xczNqzX2KVa4sdavCPJ+GPdbK/L2fz50wYFMvME6tpkl1cqyfX2
LoakuXXUJm0uOAbifWzDj7iFnTEN0ASa1u3gBlmCqA6lpySS2402SGbDAn2RmPDl
cgxyNwp5AA/dQxFuUxUnJehORE1+yDedDV2TPCGbMaPuyB8gkBfjWnfHcqHMd6ik
9LAXtqh13/EBuPogfIkB8dpMdQ9DPUPlbJGtQIUJ7L1JKW/MTiECjNPYdAM3Alj5
GrpV+jd/YnWURN+8OsyJYytDu4ZrLD6X9dbrxD2QkW8+YSBR+rnQYTHQ48y+ISpC
DPcfZOrOLEN1GibYD0RC++OEIEy2M4APIgkmf5z1zIV4hRkqmiQLcjG4ojVoSb1/
IHrX9me5JX9+nAnHmpcpctnwbBQCVFAqLL+36AJCdUO7NvAgLk12BpO7a/i7M2gQ
lWTrJP9uGRC7hBlNaLBDBPTdihm0Rv8CaoqLBIxHljIbxC65Pw4rN1XU3AgpaIG3
2b+60yftIs0jeQnCaGt2O4i3qw2wb3BUkiT6OwasJh2FZWh+eNtkKS2kx4ZVJld9
dbITy4p2ae0IPLrJmXvYAaEP1IgGsjxe7PdX+RF8+0f9N8WjjkKQVTFeLbpJ3e6L
9MSv+pBLmMEBcR9cXZiF+sNMh9gDhaau90e52q7rSIfyPLCXa7or3SOPF84OimRC
vVZnVbpg5Vmu4FPNByAqbSMYNQS9oUXq/Jkldec4OUFbOsXL/E5EXuEy8K36+qAF
z+SLACSkcFEwwySQiAdXUq25G+Cz2G/Vf1AchjESa2vAOU1O3LQuFrPhHx7hW6DN
FqLzbSZJWeSfZK8zXpFTVy59zonaCjPNNofh8JI5Uhsh/UZulwQj7fTipCQv7GAL
bmFu/4F2WCScE5AmgbPJy33p0iqoR2nn1TcMV6jLDRW90pPU7MW5WnQNvGCOuWKT
IyWhPpKEMBQ1ga3lgl0YPH27RYXspmSLvpA81M5zprufho2+728Ta4OeNFj614Kd
MbXfOXHxlwZfEtXpGl2eegga1KrSxjSk5TYxIDOzdT9WsbgxPSX3cKp5bfhDF+vk
2j4lkb5kbrLc8F3v8+YthPYfrtLQ4RlOPVuh1ecUIK4XHRUCel0u1Y5/Dy7VYMry
KrTQ3vmNjRJd5McZsKd6QaKa29v566B6jtw5diqwhvTXOIefSvVaBdStgbLP6t2V
NfrGFko5X+byxRTg0KBX4feQD6ihydMtJNcHhTRJ40RP2HAfRSb+P/pjeSjDreRk
spFRlMBBTJRsUN/o19nmvfnWekMX88ZaXYCQBbNzbx36zb7e8lW2Ierci1/MsNZx
bzdHexJHe45Ncm3x8BVvcCm3VVjudcewTYYqQrmcfMTnjEjSL0nyEvih48i1RkMv
rk0m/LNl68JglmnC0bLSkJTxwm8Oz+k1cH0k9IwsHt9EcGodd9LUvA9txSCvEEfY
FXabHvZ/FKQFg7ocKuJDnPO5qxYWTnNX07wkdXmtTIz9FQhMBw6dOMhghXIZuSpQ
o+htC8nhU0vBKjIoTk/wlt5UhueO/J5xDnNzjVUUdKn7gJZQoBdFMQQaKeTS1Vft
ChmvVVTAyh+SREz4ZUcvhWw4Mu3fp3rpDp8qYLDUS8cg9UblD1AIlR9xt4/pt5jP
X4NILVMcg+KTRO86FbmWig6Eb1X0uq1OjFLs1lYrpPLHhzSfMqcMUloxy7YJT4W7
sJyKCzR83YZp9ebx5eZcQDGFphROHTMaD2pKGW/+Fen97Y66VS2k/vLwyWkJG4Rd
V4+8E5euQgUWrz0+u3WhYz97BmxOiWdjE1MdM8I2wzbXxKLdkFoEpBWy/GufLhaO
ZT9jeogOSvCbRlWCZMTCcBcqkw61JUElp+N3aRNZjwaPT2WXLAHBBD6FBlGbRudd
n5xJYVI9hcW12OoDFSbfLMXdYK9HDNlrTXpaj8tMTOTssbtmtvcOMo2HZjNZ5zEr
E6hwSdIegqiWDXS1ta3iCleIKlSI4n0oaOMM5bzQ0fi1LHuxIlLsofrY0jo6yop8
/1oQynvmx6jiiGD67pCjzTkjXFZfNDsR3JuiAf1IlZ8iKprYQ208KETE/jkj0McB
P1FciYlwWX659ebt9Vzam8NvhZJ1uB+ZrakZvzSok6gC15B0hgrGyd/7c90Om6qN
T5vWPQpY+rp/cKmeI4i5J+of4DytB2P0g4/1doJ8E9XnmnRXeCoplizIi8xTPVS8
Wk3vV64XLUzHZ6OpVRGntEghErrl+5kEGcnX9RWkJbkbXbJysTGLIqJalQjm/Jkn
DSnydmGUQi+ThqrFBfoxQ+YIPpVtl1Qsf+LLkLr8RFvHz3WuJ7Ky2PUg/tF1eUMG
Uz+XI/OAzDaeKT630wFecQPvEJkm+cNhO0dpYuPqxnchOSuIXmfLiDimTiYthtma
mfTNkcMsqrb228f57/cMxCw0dPDA2cOJ6jwjKS4e7uybg6n3KN2k/HnX7aQNgi0H
RyX3PtAT5fSqmOKF5mgZweWYH3RFGvcH4iS6M70yz6mLUC3xjJfy58k6DKbN9l0R
XQO8XQaEZLDA0RRGg9Aq/JHHi2y+GQTnwzr5Agq84tWV6MxA60q1tf9u0D7V/uzU
KK29D9eTZRKkBHgoAoreF5hhNnjzfUYu9rXMpwAiXDfG+nezGkwuhRHqj92EegON
2Jt0Ld48YLVQbcADOQrDKHKAgULVy2DSedmPg2puxXAkfKGpfeFm2Wo5/E2Nf62s
GJMRyi4ZQB4WzA9cjb9A7b+bnNC2zirtyB9F4xfXkrSpZeQ6u1EMGwna9IgEgnDV
mau0T5dyvBauJ/9txuHmOp2xnHJ2QPvY24//Fyi2xd2PKj7nMdlKzeurmfpxGKMc
O2NuRdZ8XwyHs1aKtWvyCZwq99taJy002Kd9VFTQz4BWM2PeFH6lHvy3p0PfyTAv
VLxo8QpD5QsEaIajHxeklTx+mC36Okj13jV69steJEaBJZqSo9zloXe/Z2GwRq7c
KJR7K8Or3EazOqimD+4H2nqk3Oh+mpST6ourC/45ifD9nEPLeKHCrTuz6/dQ/vN4
85UE6bejiJlz/nGI5HgOqbR7rfJT3dJGnn0JceI2P6kDBMlqQM9w9Up1hJno10db
M9pZhPsTg1VH//BFMLWAN3r/E6+0r8XT9Ray7Lc7rs6KjR/ferrUEYqMKzkK14zD
SOdCWuIzdc+/jzgJFOl5NajNXSFy8N/1NBY/lo7tlUaCgWKnPzwiVRWQ5zkTOYGT
899+CM13croh4BAUic9PVYZUUw/OpnHMphPyFkOa3L1PC5RH9NcrOMrttoEBY/4p
aehlz/aoWW1njWSklyG8VGsfgyUy/70A7KB2vwMzsDeIYq4kmNSl7vZhV2qXC1fH
n7IYrn8UFk+a0w1KPQPp8Y0rnynl0jjbrUYZeK09qF4zIF2/OxtblnSw/qDV/nVq
ouDbPmSAYb3MCXN9JdlqE2ZMot7Cc8Sa7wAM2ckBxwxR8Ny1lcyLT/oBoUCCJUDD
i1JAnLr0u7dkqIJwraZSHIyNpAGivuvpZE3EUQTMYqz4ef2My7rGxyGFpa50dHM9
ZYKZtU8ftaAUSWBIdOLFgrhsj0qtOf99pssVzX8eXGnWppZFcvUicaypE8Bp6F/4
NYOuh8nhe6BWaVeIWOe6sy2A9pEvPTBC7f1c22i2nlJtS5Ybi9laceWTbI31Tz04
kJ80QHwkD0V8oTl7WLCkKWQgUBpcRoTVIgdARwQroLQex1Ni7KdIGDpFgrZrpRn9
o0GgooAP3jIe2sIroEJKyIkDthyuEG6jcoVvaYJOWaEecdKUMGnmAx/F/KD88NwT
OySt+CnfDu6WGez4TWWEaq9X7Fbi2Yj1ZNjg50ttl3x7HHiO7PnozgcFeb+1IFPG
lSKlulaJWG8Gkt9xtQvaQpVKDpD4LMDEUmMq3lnJmRKvwd/N0ezmt9FEpTFN32fn
rbGuxyFfN/kNHWqmsTYIu3Y/4gOF9IM/OWd0aN5jGbK6sxXjJEwNw5bD4dHAp1qD
Ayd9X0XY4dsnx6Vx7TJdsm8WetY30q6IJKXM+2M2ui4mOEirllf98PNIY55BX41R
4CTBLeZtW3x5uFRXkdF2oXy2UYOHJQO+AiEPPytQY+Zobs+hb81HSIuyFIZOTlI3
RsCj+oFTcIvLaJnBo2cRikgs4XuArxFMj+4cxlTIlQN3iPLgXX8iUuudT4F5ifEu
1VdfZCTT1YMQhwPPYJaKFbM1vSPm4BjOnDJMxl7kLEjsSAkPq62A/+wdp+u1Sswo
HJRhTB6tyrT0jpUnv92gQuraFhA3762QRZvQOXpspl1EYM+4+gSpbWxy2TLSt96w
0w+H+j4VM+eFBo4wqwkISdpFf62Wfq6jH6Y98aQGBxOGfrufQq5fgaD/zPbx7Ncr
heS4pMj0Rb+jemWXQpG8H0Cx+jDCyFyG0V08U8Qw4hAwQ6Ya1h3PjMUGInrQ4IdL
CRVAHHdSlAPWiEBNR5M2UnP1JIHt9QvDjwi0XtPT0cjsTOIokQ3SJvQt++9YS6fF
xWK1HcmAAhCRVQ5o/EpGCS5PplxcbHVGOXMjtFMpg509pDVtSMrHpkBP110YG65D
Nmnr8qHXxMz70cO+4aTiK/azwCnEf3GrwUHIEBngGSqVsRLt6Qaw01yr4hk8c37p
NYReshgLuIPkriT6BlS+xlnyXrSutk25NECXRAb285nca3KbaOkh9Likbgnxr/NG
iEkREuqvGmap2j/D6UX/dmfFcoQ/U8zP8R1AutYbAMNIcHUAolc9wMFiJfOqW6eM
1j+/U32TE6M0dGKdBrcZN7ZjAVyzwIxkikfvlvMpb5pROme6WIx53ES7flLkMQbz
gjSl7uT8omoOvak3nP5Rw22m7xeks6nAU8j4etQreRyeUpxxtYmlHEGRlVUT4pdC
QWYRKhoHZcn9FathfIasUz+Zvaivtqe78B6HRo2oZHlS28pXw5YivwMhU5WKMWQY
i9+ebIZwLX9/W6O8rUEd0aeHbG79SLTl8OMSjota6EL7Wd4aNRY5RjAU3FOemzxL
85Lo3h/uQyVuFfe17n+J2kXV4zS/UpshuX+mN6LMLrFlROHbDAEG4H6jCG5OYcfx
ATn4Ea3ENrbbVZJqIJ6K5qBNy7pbDC5aepfMp7E/ww2IgP/q1FPRQ76tFbc42XJ+
5DvVA0/rXYA4NBSj0oCgnabDODZCdoya14TxXwPRWIqi50uvms3ZFkFlQJd2tKbP
zksYiwfe2YCdDnaBc0n2C8PkUbQHuy49IV+BWd+CCIHf9SBzSYZzfFZe/HiiWs+w
Ajnb/a7uYNjG5ZvvXgDWsVMvLxzbJnKfKUQGxU0wf671H9f66Oqu9XIrScYjhAhq
RgWFbkHt93iGyx1oG9ogbPpgp5VPoUhTYLiI/uq0q6ygB/vSb1swbU0t7hCX9xGH
//LdhWwP6Mln+WWjKovUqknDkvy8AM2o8iFj6j4d/tdyxbTN8q7U4n0uy88jZi3Y
WlvMFz1ITDSAmGRSCrGkm+sHC3oTxTKZl+Crw4yFDQKTB/P8r4RMS9TkFpZs1lxW
3e2poRf+GxIfvuvpiBzd9kXUVQEzArMP8rW5YgNMJJ8W5NZnJzivD8rpV4IbMVUj
X/YFfM/brhEDdTzgLxV3gXVWB+BYjB9IJsBrIUUOjHMs1HzVXuVKQD+6OCRqq6uU
ElL3z6vV8lgRlfLGIzTdsKHBleAPkVUu3F/xvK1bkc/m5s8qLl6+5cJ8wyQ+eI/j
O9n5V3a+JAVCJdxDqMJnxU/Th8N6zU1v9vcO9UVJlM13/+PadzTRP+yORedRlcJ5
fy53YPAgujuMy0z08xJ9trwrhRz0QUbJqs1szq1/fw43Bp2owJoxrCDYOYLyc/wJ
+jmG6rsj4uPKAtRNE1TvB4rvCBuQhu+LeTGY6hQwjoClS8k3HTAkaRYQcmPWT/y/
RpqZYtm2WdP6j3VNZ+gbrBMZe+pKaVdZwXK/SkE2g94f73iMpGScODGj+HlpsJiC
hOkup04rur32iN4For1YwK3dk5v20BTS0sIO3CxK4H3+FxvhOmltP+HiIJJJACa5
olW+HmgcDDkyHstPN4iZqGCwe37IFUi1xfW0GXVujz7tMG+WdLLKbj9PFHwIqD9O
MntU/PciVz6Ccz2OOAwLSB1DPg1Ly3mPEUzhEZ7nkxQHVE3h3kLXh04wGpQ8tPGc
Y3P6qIgy6XLcIp+Giwa5hwB+25T5OcgjerZ/Hc6p0yvVXLhVDgXcEF1VDggVdg6/
3YL4XUnohgVrmLrSz/6o1v60JLAjEIwFxGl3zOA24poug0UFKALJ9AE+Kd/5fWml
IqwdwF/pju9+LYYw868ba1xsj6BESmvbSSuwaGqxYO1QQkr3gJM7IGrnZPPpJK9S
yl7j/um5XrjjjrB8UEgaQxrhnTgOyHigHNSRQYrBYLWnJ6SwtAqCcdwvxhyhr4e6
+UWLZjdunBscjGIFw/v1xC1UQEXgltewA1KJTMzwvwaNcdW4+jHh4axU70mnp2bu
Bhh4LCpNQ3it3gw5gi+hVFEZBxFRPVgk10sTzKs4Lj1DhQCYKufmgARxNidPYfNk
6vf5hQfS60+SEVNkrsYgKTBt1MoYwuyOtIAKToLykWmDDE9y+H+WHmVizvyBcBdB
C9+HWE5Qh3WEl2GBnI4glHNNld+FV/l6smdGX+RQqL/JO7YCDthaIYDO3aQZOBPZ
izicQj7L1KxCgzDFzb/PzJWoBhi6CxOp3k1P1tNDwP+NEe6CwMXPB3LOoB1ljE1S
nMBJHKI02XqQWRJ5qJilvv1Ux8uzPVILRC0Al+TvQQ3fsvhC6wVuB+9tLsN80iki
Jx85YQfeYtDZ2Hnw42au8GQUb7/NMr1RIyis52zItWNDNhvbzozw+QrnzZFegIBT
zzo/l6j7v0myBIVX8BYU3b5oT1uL21WzdWXx5BLZYSaRjMqrJi/mrz/uKCJIcMc9
HrEb+/j5p2uuVSpvRGXNkdSlsgJCFjNoV436AOtQ/rcMYmtvSR8kXTAqUj7Ct8+x
JMyRuE3GvULYyUa8DlK16Jw91fkrvGlTDVZhaApgEyh63PXFkAvw+PpUxEKFfdW3
6D9paPzDP450f/rpF8DYX5P7oBwBt0jJ/id/iTz5gd/4Xrw95sjzxQ1gMFxJulyW
6r6WVcq4DcY2HLx7zoc0x7vvtqVHKp1GrKeklDDrv6B16FdpYb4J/9IJBctzBV3n
f5kEWyV+sHoAKfdxbDcxxJh8573Sm/PyP2aY5tOT5sKML0fPKDiX1yWwoRKiB0q7
PKjwIger/njNkIqiHNxhqXRNXR1zBS/te7W3QpPeK0sAdi7NqD1RFPkELf1Pluke
c0W6cgo3QDRRb3PALeeGICmCDg5K5o3N/UHUPNVzd8wj9MPZXkQq+OdrxPeE55gi
2Yr1Bd0gsMtDCS8ASE2bN1psPS1uOWvcMiA8d64+Kbw1rFmnP70ErfZ8wtdMw3IG
BQHVuNTgkhn4zSN3vmu4skguWvH75X6WVFZxlkIM9YOolzU4RlKV/OevZQH0os1s
6VMebfOz9w2rdNojoLMWa3nNAg+fiEykRZsJXFrhoelD+1UOo45hnYlbOBWubWfT
vwG09dZEYhMZ6WakZRCTlxdxzc44sIJvvq+b4sbUsRtJP0OPkuLw07E0nOrVTsQ5
OULIAZdzz8tpV8Xp9n7zcFBW2yZTJgsyLGrBrflRcglEqDh1mrUwz6I9yd1wN9mW
gcojZkCdRY0XznckcwITduScYZh6bJKZr5Qgf8Q8NFJSee8oFPmK2onfLmmy19Dk
zndE6XLmSUmxaG5tHtxTN4UOdGnLUYNCw/+IAAuO8SvPkdqPBhQnCdrqqOp7pkZW
ZyQoWoDTiawnmTbTY0gkhlDyJjPmgqGo1sEFC0O98L2IGx1IfBsVPxtiW8enaKKA
P/3cpvvkTzuSa6cZvGII9L8bCwu6Rt3zppwcdwgX6DUowyj7tkyJFekcF5QztGCM
GvggTwW3dQkNhU96UQAZPqQ1+o408YtSA3KSEJx8MdOhw3+OsJ9OtsvGS3yl8Ydr
oNbZDzPH9MWpl00LtThZ2cD6FcchatuR906SPLeG8AB5oaukzVv7CCKz04kC+QxV
Pl5+g2CoscifkM/l85te8pv4baDicGv7IwOcB6B876RV84x2h+tbCevZgZvhPomB
I10S0gknB7ehJf5ha7y808OT+UgztlpSkKHYmvLWRl+GUxrxdrxWKiFbz5gn5H44
KdfWSDlhcO9nPf0qWC2cVtqTB5IREWaH6LURxOHFt48SP79qRxXrjJo4CpKfMCkr
HOgBcmCwDER7aIRt0zucOj0vBlMW3zNbMXTbZzR45jFFlXaum1wuDf2ZTkOQeJlf
SufVVGFGEy6kR+TrBK1C2H05NgmK5Ds6Zi0ZtvXTbNuFc5uzKxWnFhEYnOdqOnJe
ce8tenXRfYZEVk1Zi8DL7/QziJUiIkUGly6q3gTUqQQuy73QERpTmt/PqBHaQO25
eTnei3vBtw2B1H24IQAgz/wE2NPYiOrgV+m3UUlTV0js5n1IrkDLR4oWLuJNlcZc
6gl55otYbMp1bMpgss2kNsDFASzyodsmnPmYveGaT7XmUfY7T9pVuI83tMuDgggV
7H9+goROXZ0DzQPBJSPkc4ni1zjLwXWi9m94TPXfZbsoNWWL7LI2zmvDJsT2qbVw
wbpPhdXPyuVTwHnlDq+kuoaH7qv5CHJsbo4xmHXJDyLBkdZ7pMatogshTT2Cy5U2
DrWK74RjiToANRjMzq6OrKQ1M43Z/RircoG/GXZfwx7d8SQoFgQzTFNPYV5B8SoE
0+hDKMSdstrqZy03R9Ky15moP4UjsA9ZDkEHqcbgibi1mQpEiNd46lZpSUmHXoYt
0vk1zOK6WQ1LHXXKqIe9ch8h4uo7KahWWD4k5vnofgC3t/CUOsxlL/3+rqa61GaC
PZfr8hl5AxGc3wWKXb0/Uk53acxLszOf7srzP3p5IhX1L8E8glN7uF2MulcIJPUP
3TUSo+jsB0ntMKi0dPjznPTIeiwPPr/d7QKCWhBmp6gmxWOqvfxhHZ3+paMaATt9
Mb5iDFiKcNDEhu0yINRd6Yx7PymRJUeoXI3Ko57a/PoYfWGuCochffS5FRyXqq/I
i88qEWKJM87xL4vonid+ALy6caxD8q3ukjEzBbG8ZiFzhLZr0lbordsMAVCZB8vT
0QXY4LusvyLOY6ym3URSAJMo34JbJZO2x73Lmp1SlOKR+MDqP7f9Svx4rmwGPAJe
cRw38aPSRb4RAFT/86F0/nE0YW74Zxiyokq6YMKFpaKbKrkuPmJfTi3Boo2TFFVx
zHO2Z5ajL4P77OaF1vrLKH+3FC4uwvULqNI6pRCYE7EbYe68flPto87P2u662P/I
PxXblDi8wPyVRmds1LlIlh6gPL0W4gryfv5og6yi/k98/+aZ52hH+VEE9Ul4aYOD
mnC0MFu4sRclspJEw4gqe8/XDZGo0yrBm7jaFgQQ5UEuJcrjC+sEaTXiUq/32tcM
HOAymcfYTFJzHSq6aOiF9kNduU01w8s4ORZ1VQbzx3jTBnQadgFrxBWKqs3y6e7S
iS6EvJz9wIALr2fnADvU42grP1ciq8re2zin3enwwq8rmFt18QScj5Iseho2NQEL
5Bi3fP0/oCaV0iZrN3BhfizIszZv+6SmLi5NGacky2LMOMaweFuU4mhKWc0Q+99e
bHIJYuukAlGar0kYTw8EfceeWINBuO5SYL9Lt6y7SfvdvSeSzw/wT0riQpK8TBOy
ZIz325KIA64/ce9RYktgMWYZ1udCl4ECr6W24erSQFk2FOw78rrMwsOwpipA7kVe
k1A9uqh/qKNZcdFBgSKHRH6Us70Ra/rVTLUVSn1nTVEN87kQXx6EQJ2bcKkAt/+y
yfVZui77KwZdkLnTg3xdD3bA3KWwIIiomiDmzINzj7AHYEQgAGRH4ZijuWhTBpDA
GOc9oUvJGEZ6ZQBESFZAV93HuHLWQ9RANz5r/60R4fQqRqGVPSz9bWKmuXHPNx63
5DA8m6cLF8YQJPtvpwjjWSMBGD/JxBzAnFDUJB9QkuHmVMFsus2n5zKROuXyh0KJ
DHYlRNeoqEib2KXHXy4UtV66jfVVMrjTmsXI4ipI53Lvm3NS6ucTCmLoG6g7wAZj
b5niQZYW8NpUG9e0oyBMWcpYDWMblEEfCKQRUs6darVdSzHyBblvMO5JNgsNH+2x
+yGl8dNlUng74O9/QNZHIGbzqHfyDhVeWM+VvIxyJD7dwGL5PC5EtqbdYpQMWp9W
PEIUNi11Hc8yngDLCjqwCeagAI7qh37YsMRSSOeaKQioUS0RMWnVm2xZVY+WkHXC
WS5YisU2VVpqMctL2gYxTuZ1/pbq478CiKlsMoWz3GW43oBhUtF5kYsluz2yyM23
Z55nIDOLo4b183A0sqDMJi4Fr7XrjCWQEKCeZZh/LyJpq4DNE/oyFWy5oUpN0bxx
DisIZ/DlXRvuuJuO1ZaKfT8o5mz2OsvYMpNiD5seJFGwyHttNyExFw5yvvShW7RW
sI7wsKekY9YHCqp13tqyrjEfllyJGyncPu0DEMJZScLhUF4Ii74+4j6s/jQoIJsJ
KQUoIOp435Kn6wzkVHDJISTxvjax7pGTy1BQHihoh0eXgZhPJ6AXXbvNXXzZPzqY
D3wbs1v+FsHd/aoCTO+s5wJXPQbObF1yhNZnU3pHomVes4ilITQs4eXCP6aTg/Q/
4q9PU4KK9imdj+nyIwcOnJwHoOzbbymxzO0HRNPfg0nWOcuDmSv2Od1O1cuHmRru
jhQHVi7AwzgPqSfcjIV54w40bCdzfpgBuqbFzK4oUYAo+j2j9Hk8o4gdtzXJ0kol
HxrQGNIZSI8S2feHRPYcMq8QDM4A8/vSgzhhCO2iECd5fT8zArCo5iZQlhIFIEW1
1On/5/mcgDl2mPQSsJihEYKZM1aCUA4CldWYJ91Lz/2Tq6QdfWtE8aGcG3CshDIZ
ZXTfPDn2Dho8l9Yx8dhQ8CHmT18alvbbKSf4XgoHrE0WKb3wPPOG5rpgWS+GpylJ
WIbFLatIVmphPZDyblvCE9zgUSbwBE+TIatC15+LudXZH3WMDozxqpnf66zuceh+
tth1eRW5E9U+WG/I80d3PM1WfLksmW0mObSxlrQsN2z0f2+ORODkxN5pnVD1qc2V
57X2WcqIoRLTdZS9Y5TQqifwWx7quY3onSLD+6zfNNNGj9VE3Y0xB9tQRX/fgt5e
XVIZbgdYXhk24efz/YmCCDi1ur3IFj5rb2m/pfcoJImZEanaNwmIOePzBdG6CvJG
TjosEjO16iM33S0+S/JLfo3i5aWH6+Q3Y8yF59rfo9+cH7qGXObMKeR4RUYycXb1
4tLScSEEA4kWLmDwWwiznWxpuKZW9usEkwh/ehtJNe4lujQHun5NGy4BIndzGX4y
PTVREdy4w6mhrjAISnNvevY3jnuaLF5fRkshWuSSp1pKt8ONaJqpS84JZ4b46BNR
wSjjsAzCavDqRSF/OnyU9ZSXEjv3KtivS5ot4MeDqTK2plHmHTeYHLrVFxLlfGso
pPOJaXHpOwWS+vfL6jQ3y+sWbtMhDhl6GC9IVZhvUYV4X1aRpGjVVF/x2gfXXQ+p
fwJAF7SB7WeJoU1b6Z8NWevY6lCfouNyWhbY5uii5s/LDQwG7wmTOr3xeVAwqfBd
6w2tQP/azYs41hRTFc9SfN8O+Bih+Cq5tKpk4EsejKb217KbSBCPRTanTm/lpq2Y
axsBCYIjVHGgjXdQs7cyDOr83xavfU1/37QtDmLf3VvHTemw4Vl2YrQvg3QAtA2V
BVp1EA5OQNeqeg58iBBoHUNz7iHHe312hVACHZFRx+X2a5Ep5OFj6KEjz4FvUBE9
MTrlLvuMeYNjsrgk+yWycufyOfuaLCeD8sFORajWz+GBrr4OKfUoAfZXt4kz5LnX
wBZ6RGUF53LTqC2mO/f9mn7BXSIKhjpGUZ3qiX/9HfhN0l9ilfBGCrCOd9REuBRK
xztUH9nIfmvi25vJl3pVmcPdaDgHc4YW/FwUf2jJR2hUDOaZKaMgLmbiLrnVfwkC
La0wZjv5MKULLDOEZO+Voog+5LvjvGpA7enaCDqRalOIi3LraVRJ6qBLpec/zgqu
M59WBsExqaWIwNtz8TjrnPJjJgIbWPjgV/kUlUK9Fem5KduuiVkddi7VfA+NFwV3
mR3ZGl3tTjPnA71beGt+vQ49mezR1QQry0i8jS3+OUgDdpIewNWoWfLdp1VSjdby
TLdpeHjsS0Kb5D4mbCyJOY7MP8v41c/Z8sHu58N4wdx5EoJMKifNHL1ujNDokjDU
iGaSvnXG9bwwWr9yAan9UKmgN0tC+Y4L91TRrKcDdwLZ0tlEqEznTi+Az+dc8880
FGYASuTlekby3I3B2S/yCU9TRKNlQCVQFX5FABR+dygA5WIQBwDeTNXhXSz1Pm/R
Qxjug8F0/HrZbuo/2yijArIsIR71XTVlQnG0ev8gP/Tsxx3bjPqsjuGgb2l5eYz3
YFrLKd4o7Upe7hs52k/G7d5c0UvuXK2ilnSzOzm8d2jJzOPJ2jXOi1XBw3MaNlPQ
M20MRwsHVnsfJ3P65wx207TXyrE/+iNfL16LRvZzyTX03Xz7cDqwxmN80b6qavm8
u/EaD6+9gDRgrlPwNCyTcPupljoRxrismnaFFNXXCmVS/lkiMixSMvmTtQHqo7nm
aQlT6qZ4FDSOFyTgAWkWpsBzBPPjIW1g1A6uE7uaU+NZ44lfWN1vYxmusOxVWthL
sNNngBoZ0yqzYH85bAnNVPsKemL5oXDwy8s4dTgVTfNtUAIO0srsRyqHDfieJ9Co
tjmFoNkgqlFaheJOX8wJp1nri5i5GmgvmbzUM0A/ssN3m0ijkZOl/JH94KwkWGAy
6TYVzB35jAKe7cEO5juQ/jyQG4WSaBhdQybpudek9MousqMrxA6JjXOFYap8SYit
vaN/rvXC+xMLE81k2J19fsvA4a96Q3A/8+0pnVfPqv31ubFPKapekacRL7EkMnWF
RHBw5hXVCUBk+QjV3Aj4yoeW9kGtCKEIbGfHZ3gXdRppbeHhpuHVMtUsM7UPAjqs
bqhknbhOavpiSe0V/GKuObOEQpT9f06I0F6vI4OMTAodmJKYq1jf4XEXcuDBc4WX
W0djArRd9d/vZTYNnt3BjoBx1wnN3vNd1FvRzxAmTpu3wweT6NDIQ5CJ5Un8UnhM
JhtU4mIRDGkeYZ/d0L8T+cGe9QChck83FAX4L4vUkWu4attz0UiySB2Y6MW1uS7M
UcgQFXv84U2PV0GTXCM0I6eSgUc9F5Z4J4pfCjpV0/73TUjgqlBaLBygYey8BhWg
uW/27c4C27GZfSQ/Alb5XZh9lJzpEXLWuNf221dfuk14F5xJeKstr/Tac2HmWU41
zY6u0Mj1xeSKp6RJyCDJ1mZmR59TrmLWpjUMkA7hX1IJMwjyq8AUXwrX+7KyKzc+
DBvYXRYP/N5ols9oQ4Sh7/Pvj6ukZLwq5H8Ap3Bc/HN3cka3bUJjnOGkFyEqATf8
a+hr/AYMG0v8XBx9gSrtCmCs9hWS62SQ1lSGgKZxAWcN+AAgr7ifcwp3va7LW5Dv
f8ZOcThuZyuvzSmj5JjhhJxGOG0pbn2rk7k0Lfu3LD9ziHEwFeNVITXwZSxv+jgO
2L+HdsI0U3zYhWUp3izV2ZXQVs3vhlf7jtYiGsT21gsxaIH5Bu7/0WtMY9SVZgix
7amb9mh8ZHp3YKd2WctE7oU/4l9g3Bqlx8wOqgqf7R28eqFdMXCwyOrt6Y/+uyT6
VyHHeP6hIB0Xap/k57fWgwNxcmBQF9OL2DddOR/jkDSZoNQTSq1C8TR8rsdqicul
5GKvaIHJFSbd+J5hUcJdmw0Wwe/tkrBHGChd/0Uodn9Jk2JBcKzQd6WDR0trG0Kz
KIfilpEIuy96fccmuAJh5SrpvGkQ3uMBWZg1qOxMwO3hcmKpJCSPokFS4N/k9pgO
pVjaRrhWBq0AN1I/+XuOKdWSmXiumJ1IONyluT83wsJXQsZr/8hBrjNAVB85Rsog
AWYxWqqHs2kQIrFV0Bzjx0bIempAF2oVms2VmgyRc0r2REKU6V8/32ru7dQ1fnKk
ksS9eTXZY+CBjf7n0eVlZe0ZIKCC4qXAhs/2FWvqoiAZNRC44aez1opiNsGH/b8f
W/jmZM/6p4PAmjPtSoKYpHbNe8SY9mGrpkrDo2CUvatJJ+XfMp2rhEw/Y3bZv0tb
ISSuGHw9p5FpWvTcSx3i2rmszmClEymNG8iziW1FAJLfdlK4n5zKhB4+vDCrpE3G
r8YLivmAKzzuDPshZluGKLoKMZO6G5DL4sIQMKdZc0GCzVp0TwIhd4snwxys042U
QaHXdG24JiV/QIWIGNP4J5R1/FNBPiN/0l8rrZOJxpvO1vPgf15jkHJiknqt9+DE
HDv0o3BRzh8c3+SDbTjvXv906z76VKXI6D5s+l/Lb6O9XaecU5JGjwboKWNMox+F
bnpxBlHuxInBPtaPpq3yNOGDnMa13qx8InEiH5AqJ++hAHBtgkatZIbDeH7qwI0O
AVk72HO9mxeEhY4HT0T13CZ1pHG6zY8wsswW07fs1kQUTg/j1RQ9BGlA0Ch/cghG
vY0BbeYKvcLO+UPGHq8OjXvWSG2OCMGWYVvbA8FurLFyFmFjhTOeGaSlYRmQGw7S
jwkQv0jkBHqMcqD1SoB4aj32QOYNMvUVKs5eEmDW+tc/LHCqGxoOOtGMgkKoXQ/W
JuGoU7YMud0eBdiVgbVNV+0vITvGdBfc28NSB5aDbqe2CL/uhrO4MIpjxzDZ1rPl
3Jb2lmAOJFI2fA/5p7IrkwdGNRubBc4lVTW6k5mnlkkWLFCqMLHxE0mdCCsgRYuM
9dFCHoAS+Utdv/GOPoRU1hrBn0ZynxF2P56bZFqpzWezIN6/k/YHF87ARsyqKkfd
f7uOPMDYx2U6hpdLlkudKmr1g6gL1SyUpZaNTu0IJ2p7eSJ9LMqsFYOGrx8S0KKB
2cbdHmwFi2CAoXNWCGVfrmZ1PZ7l5LTgenrPJLmYQP0RuckkboZmtSEw+Frj7d0y
bJNdtbKuJMo6HuPqBwaD5VdiC6/Ml7KHOdit+AFul7ZeOYETPmCv07nVXfkK9JUD
qeAjywzOjHz5ZflZ393//+bXSQq4m5PadABhjYOJmU6fn3EIsnBlJ6iYD7GlhN1s
Yh798hUrdEn0+g4qeYh47BEHRh85jiCw3411fdVOHoETNxtMy3POivGrPvHp5ydd
X8BCTO359/wkZxOH4kEmk4owpdvxSDpaHY23njZqdL0kz8NwVR+4A3QqNVZ2rDbu
s0LxY3+uZ0sb9k5ep5pmWwhJmnknJvX7n1eIIjeFtmV+gphIiE6gT7O56I5TnLeB
q6kLZDidg+h0cma6S1StMHYAYZEGJ1MHXVCd/rXJENLm00zMde6QFEImAn627SFN
HRxGsunV194lzDdJDNs7OgSUyruQL6ZO15urZHoHNPtQQcIcmijQ8MAQpN/Jo5j4
t5P1gqusMkMZO1FzlRNR5CgPbRlmM4nhjQjx/I8Wj+mr9XnwIThM+3hvzqnYpjeB
fnH4sQuk/ayCorqsuzdWwVrWbZCNylpcgu+vMhr6iBOJKvVC1AA+OYSsmBUviFeN
wmdtub2I8KY2EQEhNRYcii6GipesOLIid3nWPQZ+VC+39QyyrRq9Mgm2p28wIsgn
qOPBXp8rSjF9B6cQ54U8El05uf0c3Gu8qXgJThSj9X2JucDM+gcW3urX8HFZsDRi
7VBGfhYtH3lTPcsqWfM3G2wTeemFRFSv+zxnjuwVlzqlgt3eDSw0bJ6LXGYAm/vv
vIhaBPIOKMZkyBjmgs87xOd0rlFkOXAknZmwWsei8FJhQcm2wDiVwcP2Ku3NfpSF
Gi92Or+4F/QBBG3IN7+2O38fuho1vP5Do4pQbP5AweDxt/46KQ9t9JcofXcQsaWF
G+SDHOHCsLTX+IaR4MHbnWOwKFnTeTZw+PIMzyzpBkgUZtQ9A+G+GgJTnfFCz3rr
zl7AzLKvmnPTdYUj/s73bxRCZrL0b4TnBijB3Cvnbf017+cUydO7LVfwVGw2WVaG
undOv8KSUuOU++TA/Y+NzJP4R8tgwUiSPsVxYcGnNgk4LB42eLEUP+rof0A7dxog
qGHcX3VANYKSKTPDVc9QkBjO9ZPFiD+ZpyVLQOD9IYh/BXSw8fDCeiMENg5I3Lkp
4Pb67OX1kE9eTjg5F23d7WGyhix69bRBhebX0zJWiYO3cQ4meV+R0suSWHKc5nUg
P0e4pSWqOj45Z6dAIBSd3XXLlRetl04lC42K4p7vZ8ZLKfh893QtpCCl1qAp2ny3
A3XMv/xMLcZxUcPxaJLMxAjUFjoKHSkvinpsvB3yiSs1pnrA0Y78O58E91V9RBRK
49NpEPt/UthGk1BPPiHzOYCeiZcSWQ3e4V+olcfqbkEiZKUSv7KB33PcIENf6nCJ
sH0p7IEeBorF514LDOZiwhYNizWooEfZRd+lUAuwUHRiM55BPBNlO/OQQwR9p8dM
qucv6KUrNeT2W2+3zbremkxLrwOLodXAGErTXsIeRs1B7oJ4Oi2p9dDqGLh0BXY/
oykff8WiWUzuKkEfftDppg85NjDY9OQwUZb216lsvnTRLCfhUtE384/dRWmeScTk
Evm7xYiCqxeWfclTkrslfy1uRX+lrB1O0wGeAv0qiuCoXFezJdlHN40F19s1YIK5
MFPyCancM3V+qA698P3RSsVlZMAczMusIXgPyUePTYT23An2Jj57fWXbbTJoo3lM
Q5Ptwb4UMGrS3z6X2Xfsq/KHfJHivLUxIPPpK2ZK8QHjIifGqdkLkGt2L0LoE4n7
SYlLyK8w34tRvGk3PTXTt9XH/L895BZh26fzuStf2Jb+qau4kuK15EiQvm43lHtE
1PLNN2WgJadLU+AGR+PfTY5DCdlQgYAPTj12Jf/2/finNqsPTpVtlRp/DdXb4tI1
+m4s43epf7pP6LJBqa4kXOpBNGN9VaDLaw9vQVoWYBOveUtjDCqya01LAcfG8/gO
tYSBJ67d2ZnsDuEciBW1vaDdAiJrPMT1DbxJEpkxEgJ/bjNXiswJyxUsOZ8Ge14E
seKmUtudbo+YFpUre4sBx5Oyab/USs35KgvMf4nOEuH9k7WYSesVw4Njpjnk3AMP
fYU5RPvQhAcLc04MiQML1wKWEoYmRFKTPqx7DAEszjvxbSGhvRXaxykCcSUB/cyk
4klsvweoSEaYM/Po/9zIHB09HzMhHtNarmLV4WCjfpd252NJ1/lr1AQmZH7ftnri
Fb2Gn2VhSkZSsEPvLS1GYnawVDmSJ5xDcAu9zT6XvgRXdiovf/BQKUZgp264VRFH
k/Arx26Id5hhh2mXh1jtwBIf1wPJv3EomhiDD+JKGxyH31gfRVGY5Rn09pAKV3v6
7hHlOBR6ZOc/Q+bzkJe7G5WjcU5otihZWM1O+q9ukZIbSBsHOAzu9rpFCFuzZtl3
v4l5wjMsWw/jggChSUXWibZRFTbpEMO8cKxoYghAFQroMhE5onrxsoBM1liNh5VD
P12p5p2p4OPtZaqslwf5LkSynH9BnSFqAfuzLZUjDDsmsDT0FthsvQgtXvBJnXTr
K13HjGIocgTK/8O/rG6bGFxPjUOjLY8y3yeK2NrVMT/bdYMPdJd/4zoT3WL6N/OD
xuA8qwWa+X85lP7rHGL5fCwrFYc9so2yfNVV/vlNQ2AbsvvFRRkkchCVgsqB4bUx
LxkdT6/1HOOu2idbVIg8tge9pkO2eyVbTL2XZj6KF+s2DpnFJXMb57CLM1pdqfzI
QNP6BRQ/zSb69sily/ipEaLLVsoQJYZ1UXQQ5hAIPaGbldkWTFwWw/luXYoAwBHf
XjrnSaBewx7gTn05Nd6VTHKSeWtcRxPsn27pSd7XS7Kc/857FZdzlkIPQGJbz9Z/
0ZGfeaHIvNcsBuZguj6FUU9vDV1nQcXeHlzYehkkE/drqe9wGbnLTrohhjqIaPw4
N5F6xmDo+9QbQ4rcFvthWHRoMIGAeVE75nZtwsPI0LiljNj80O3ryc7WKGstn9dE
PAHdQvN7Dl7N3NMWFXD6jbgk1cRoCZgRpq1LGmoWUBrYgBhqUiaOQzvwb512/jQ/
lGOr95TdfU/NUKydti+4H5HgSPigxEZpwe//0qSjj1p9s8w407tUA/YI7NEQbGn5
wTyBEvYloI8kUFOnlKqVA3dMXbh/wXA2f6KwVF62POkPi5rXCMCkMsrE6jPY9V17
oECEFb5EkTNSHDfdlyW3Qn57PKjoNs2j64eQ8gkmZLsLd7BVvSfJ6X2sU80nL/Kz
uBkJR8pIWYLFYzJcyOLyvswIZMsXGHSds2tV9ZPdGeTUFzHE3G4md0M1x6wZNbd8
8ff5atMUxIlHCu2rMs8FEZzlfw6VgHVmsjWV/OKwVJf9tJdA/c98weU52HSG0VYZ
QFybOsX3zmSOIxz29WsPKFvdHMkdHKWjng4NS+cHX7IPN7DOVr57deMpXFOklfWz
HsKi4FrK3r/5joI4aIp74dFZmavCPXG/fhvqEXAwd/ASLhC/XwyOdmT/OaRXPrQV
nmd4+SSmU9yD8jpDgJcBXVCFqJQPcYRqsZDDmf7u2r8wCSSd8xAqRRSS07/l3PaK
Mbv0Sv4trQslJ/Agf1MMF4AqJOa89jJtn6byoGz+oLYUm8vvh8i/IVd1/vrgIyhk
1vqzUzwpF9fl5Yj//uB9V3shrQPyKNq3ZaeompWcx/GYhwxCdwOZtTa+WtN89Mfw
cd+SeE6TmzJCQg0tU1m+OwZWj4xicaGdLBmg2xf9MvxLGDbM3mHFck4P44T+U2dU
Zvaa8GWk4t3sdn3NjJORnLIw0wjRzypeR6BeK8ZRTZD8LCV739bZW5Qr/6YdjQPa
olVas36CboYSEDzpOSRyxPpOERqUysbY9eh01XftUfs2BFGsSyWlFRk72Fyh2Ve8
DJ7J3RyL6x8tLw//TGBuCQCNydFM9lIoooZZhIAyeHX3q/5GLwDhPCDzFMzf7x7/
MVaCkAsoDTbkkJXe4FiPbjCyTeDZaOuyJZybsqjkE1HMLutSKIRcIPB2Zq93cQ07
xnWSRhPZ122Och+PzjJu/+l5xhz92xyWtndwiYNsv3NRbWqSNmILyK0vEqbpek5T
7N93USyObJdDxcXkJJx1YZ2t6o9DSMsFhSa/95TOFijKD32XUXHVHOJ4KsPPG9bd
MNqT/Vv1GxpotrrQNN4jn2Ke5IXRwZ5YY2CWkHtQw5GxY+zipBqbX64WoPPy0X0r
WI4Aq1BqUMFukh8bANjDtX0Js4/PoM1GpLJu8WF/qV9SAJ6gobz6r75r2lbQUL9P
d4rD1zpIRNPrzCmllXq0mtk1jXGgPnIMgxYWVvU1nzoARgnrqe4ZzmnPMS4DG6LO
/rV7tWf1/olhfk4lagulO0H/fOcgPvycgqVjnY/RWt5E5lxIn8OhpETS8XNaxtHe
74hG1E9AJPaS+fjB3PXLFuPbNChlDXdgiDyDD4A1CMh5BP1cj5b83Xpl4BsG6Yxp
ckfS8b45EZczoeczpjR74+0b6n+PtmAXEMKU+f4sIykQtKZ/3StkTulW2X7HADDW
fGmjKcgyOQRrh+UfD7BvHxiZ3ggdj25Fc9JjjpBw/GcTUYAehh71J/HyJxz1JoYk
bNaSPRqdwL3QSscsJel0ry6804vXWxra31Up6vhyNqRCBqjKZLHHR4djt255TFRR
dYenD1BK/gO+YgbgwRKDEbI8Pf/eoW1T5P/g4Dv0ATHuLCW/HzSePqK7cFNO0mzn
wrS7mukhRFHbje3M0nqDa2tGv1U8mn7DNumhQAMxXnFrwHZoyQYDhrB1ok/VZINE
zF1nfLxQvyKTRHDQtgUKRObLngSn7HBwZy9lfYJNkmurniZTo6TDma4WebPguPsX
EppCQlVBc9h9fBDPHYpaS3+N3cKm1HJfFNBZdWYq0nhLa1y59REP/go+FAbEbmiK
nNGEuKPRNKMJiyN08NwLVfO7pYJLFF1BA/hNFjGrP2ZCzAR6gcSK90cGypfFFKv5
530kV0hxyt1TOoQScfvE6+f963p43TreJdpDcsOYJS1oIi2IEH6Q864C576vnjAB
Z3GDKgNiLkq9kbgOVuA5/1rPwVLXxC5eOZ133pJpklm5kAZ68m+ez0A1FNxCSuLz
TaPvd8HoUFtdEVXYzkxtnJZCEz3dFiTmm+UfDgCExo5vgSA3zWD3YOHq0FufeYCj
8EtJw2wrEHTvGnN90aFO9d4DznALrJfU87upNCrtL73yua2ZpxYwF3pKZoc0Gt8j
WGJ95VHfAHXhkX9QIfARXQfzyG+/QH3+JJrSQfL5obS5xsAKeODsHwGv4GQg6Cag
ek5deVen5N7TCZbv1D2Co9F7JGELaYpI7HxVcFFxxe65JkgeoIw7U9UoLbYzOiBV
gYbAMK5sdmEil0QARudCuMlAFJ+6uffELT+pUs0dlZNYQAfcm/OXu/L/VJJFX9XB
cy0fpoDf3R/+eKdUYR0cJBUmRweHy4oEHU+H3g2gTF+WWN+QQeGESQ04RrVYLF73
hVfCB0Mo9NQlCXQqJMtBWu3OCLtdl21XCesVtmW6HjDMP3rx6YEzHTfwLYY3JKrj
NPAWh1rfaAHMccESMbu6JgZOOdlE1l2u6NfnD/JaybExyb9S+yF9L8VyADf7MyjX
Gyfd/OLi35JQehNGsg1HhzIGtE2qRda5Z5tPtEfNw5WFRiLlLotcOvv5lYFYCEw0
qMJRMW+ZlCQfA+hRCa+omwnrxKuWGCgHSfFsrPMsUvnGroQBOWYrA2pPTcAxdnoE
cj1WWhogEgsXaj8yBobw/Y2/nVXy84w/Vi/Jnlj8X0gHf5j38V0PlBDDv5veNtVU
pJhO6hygBAqdYRH4yljKEP5lUX+CnjHiSR0Vgk85UiV3j/ARt5jPLLtmkplhAe4I
FAccJ5vtnxDrdRcId61RGQzR0ssHfItgOIhQyM10LUjcFtlMeDOWFkUFUiO0MIl+
uYF4Sege4srgjn6yOGSCkcfQSDEnoWwDBal8l/VLOypQj9aiDJ9J0D8nlAxILvYu
NzW5wSjT5GOCfWNmUtOV4PkuOnklCc0XBSNjWdWdBqgTItBpYF+3nWwH4CMPsGfg
NC9RWSAvhKBShA6sxOcTs8CXMj+I5rB8RVCPR15/KyY35LlSHOo0/HnZJT7GNcWy
j2vpyKWEgEqxx8s8wJitiMDJZL2H668vVt7UVgGOSTR3m2MJP1urXmFlP7xYkKzU
IlNvzfUjejPxxfQyqkEDJ6u6uitavZhU5h1AfHbuhmTFFcRlZsB3nXUrXJbKfNai
Hbc2fRRtPyrFkOO79rZDHC4gWmh9hMkIiRTzRC76RQ8CA//BQ+KC/sgUThP++lkf
xM747cuEKepcqa7/3X0ltEuQrbZPX0GxbpAv3SqL7xZYDrRdtmp89opRCuu4nnJ8
nqEQLEu63ZggfO4QzjYodswR+VRRsJpfnpF86XGvfwgJ5ja/U9HmDPmMJxgAiWFo
tCb6mmQdpDTrnFxqXxy0jN258mhsk4oMOyPPhXkS8FwFtjRnhRO/3hahzfdMWk1c
HxMk65hTh2Ki8ZsmNP9+9eJw2Z2Ja8sYWgY0z7j057uZPsPddkGcJ2m2EQS95bu9
q/eOe1v7jjeUX39iF9bmYijIburh6zTkiv8J/8e4/qF0MMPi91jlkyReahCHyFje
tSyN8sopxca5ynBpxLDMJeB119WzQ3kIyVdNLvbTa5WiljKkSwuscXDZJIICV6FS
ZF/d1a+TfFS5a7Ov4wihKgJn5mU0uCGLNUQSC9QWVOsqgs+hal1aDcol0y68kREW
x5vqOPjUwk7maEcFHzZCf+Zl8hjtYPlNqmrcURMZXiKJDZl+6D9eW2TTL7omsq+4
bhfE9HgOeMVLVR1X8FvYDvLlrglnf5J6iRAXHImT0DAx4sn7m/NHUiK+ttqHecTY
ye5IHzhogbxqjfLNeKTWBL82KXwaDH7iDP8pm4GLLyHgUXi+/Bimdo2ThD27Q+Mv
OubASnqGTCmucYuuQ2jO6rEU45gVJxAW1GtVrE6MT+Yc9zfd6i309KrLkyvYLRkI
K+Nw9cMIjWhNE08lfITxE6BG5O9XI9sd2q/kLF/DbZBuW8wogEJXfkphz32oCVUc
TG7MQUmMhmw+/4ZAvsTMR3hsOj1qUpdXx1TBFHc4dnlrj03lIInoMNwOF9DABZ5N
QRU//W7cH4J1ZLQifVPsP3Io+fBgx1qbnaoV3XtWuvdXUstXXEyc7x5x/1rqBUZF
1PluVyrABOkTVhbJGWjSPZX/dKZwqzGAtcPQEPJHu175Nogs1xLwOmggOWFEJ60e
QH4x1d/+WkzzNkMdzCH+9MSoyRVh8DoSxsDy1w2grnqCi1Z6tMEGDJoxQ2gQSbjy
rkA3ODGcCPaLx6LICwWpfkyjWKilKsaBWeeuhNEKXMzdzVo199Z7ri2HpgMl5Z7w
A9ZClNqbHKXwHPM+yKcmXvrmAlrCXg46kCGmriw/WggrfmQ8t6bQwK83jY35HFtk
qMbT9EmiYEAlPk9YZ5r00W6QrN1iIz02EOeh+lzSbMt8xEQI5drECFdtnb/7y7qR
beYbwVRrk9dE7kokzPnfh8avGUo7Otdy3UlVuANsBfAH4wQuSI2wpI/8k9zlc+gj
sGPkYmFNeKIZToFp8PMrDwVTdhwn+WpXROxLt6VRqK1lTwM9DOQ9kMApFXhMcJ9m
wQl3/dTTSIId3K/HyL4Mdr7qBCmTseO5b0lEQDgoq7fJiezfgRtmb/2g8AMdUGfW
DoHseiqd0h5RNQWE0VI7SHtUbY39oAtC+x2GhnRRUnygc3oUvlp/HB10C/y60sd6
uiwXQFxNcwE1sJi/isBCnYjw2tMK2sVicn8fVu2EF66ruQf0l7W1NFyGV705+1B8
epygibzuuEj3BUG9kdYyHAuEeEVCefygB9twii9l96/rUgtY5ndxCyuQ5RBXsBxJ
mWfL/xE4dzkO+l7SFm3KUlpXCeIF5IuUenAQaJ0WpvwZfM74lqa2AfanR6Q51/2r
XnNnpbtjhzQGenlHWpy3Fclc8J4WL176J38xGJPS+W7lPOsgcQVNECkBQPRJGKCA
vDkNYx7EiXmePKY3wm8TSkR9c8HEiAaXn2AVWgqbaS/U9Hg1vSfpihCZrbiCoSUJ
xaqzYrN7VNC6FQ/V37U/xe4rWLg2NB6WGwqrZAsqq4NMx391RIbQCnSDd2kXYgWH
Mvfd66BuWhBHAHxqi3M6D8FbDdeO2N2JwDRaTF8Sg9Ys2ILm7A7DHMx+VH0ioOgi
YwZSLt29S0MFRiPkl5oxVtFdeFaeXcY8zR7wjrj6TU38ddMKKk0FzUqMJlg+Wjk6
MTDdyEvSAUY07iCRADtfdqvzCwYJL/wgN7GUaOxYs3/0aiIbyOnpjbHev5tamrfV
4jcUwfTkfz3waNOasXoQftz3OgvnRpswVJ5Lc/BEB7U6Mgf9n8h3h4lz3Ja0GOwn
1KJGclJ2KswE5gFT3rRIzkl8gAjPWY18Oyy//UhKZi9Eb4garHfVidYtEGrlmOpU
ve7aOxTUPJlEr/TfK3VOrEYlIJW+TJxzXUc0WnbFGhKsftPAIwGrvxuQnApuo3d8
LZTrt89/uNVbROXqydWAKAwBxV7a7uH6txFJVo2jU+oUnnyU965yat1aMpr9PwAV
K77HExDyi+JJ38sw1FES7e2As2KPzRiQp0wz8agv0hfC+8CRnHhkkxh8Q4MRv1Ql
4tTDXnIYKA+lcURtwTly1XGCZJhSgOOckG6BqsTu3kkLXx7UESwaEdEWbhogwrhY
4DMcuAUcGJYo7SxVQ5vqtK38x6K2pkbgZGqVj/PQqmj28WeVDQQ/lIVCv4S8w2k2
q1b0Rsm4/S7SFAvZVB/jT7e/z9U9EXffe+cCN2mbpiyWsH7Vu8ixlfLbcQCseR5N
VXgVKCurfUFzl4Uxlz2hgqQ8o3PS2QCemXoGyZ9IWuPI8yp5DqkB+mvic2dwKFQo
poMeR8azGH6OBK6DX/MPRijFrXS0HliHpSOn5zz8Fhstyu9kINZqpiqqHJdrtT50
LjMtqIc8uBakrqfM5n/F352o2TGVbILlNk/AUn0Gn40xLRVm4DvIiCrmyV+V4ILL
GQf2r262ub/t34JV26H5QJAYoWlVbvG4mGaSGlKXeXHJF8ePPqbktme1j6ffvsaW
h8dhmQnNBPwdfOlzKwN/QKlXTCAkNTuTUcKGkHqyLJtrlPi+qYOLaAwLHvOxowZl
XPmjUBliXyXzazdqNUxF7WKA+EZUMltlbI8GC9qiR+kmXefQwfi7zepyl+bDjFlB
hZUpZBMWNA8qq+3ZKJkxvAKBaUHRsm5COVMyufxdorywruabHGv8B6/d2GttkxGG
hht+OYBf1ihNyySkbgi9pi8Rz5TWsdtiVFa6XjNmujKyEMHUS4+7xZiAK1bCXWRD
whl4oxOKYUJT02pCizD7w37uDjfU34wc1s+QhDmXkx9FM441Ol1h+E0wC+WJBhin
XzlcdIUj6+x3J2BpYCGKNJ9wSJQwqFwNZv5WqINVNIJuNsMHYdgI4lA7L+BhKrL/
x+ngHaSl/tz+46RBKltXXln+iTUsXlef4WCqEmU0pwIGyKQ0Z4uIA7vYZeTuJzNg
ULPtBu011uHl6P7RykoYhGR+tqqnllk9XEiFji+BZwthnBitsSRhE3q+Nm6Z8mWH
wwEg6JYvLeeNoeSPxwd8liEwTKsinCwr651ocnDJhs6fi1aPxbfO+K5C7/7y9EGb
/6Ka8jA9XPScxLwnXThcIjqmW5n6neaGUtxkEbV+RvG3J2G3ixKSiYz0sbaAx4lE
GBA30XAbxbLuVqus4Qdszp9FFY94RfQirE665otDByGRAFBmcVmneXC+CFIHhKK8
BUjGe1x2qQFgHPz3m0Q9988QQf8CR7DJJOp26V4VMr7mTDbCBb60Aj0Nh3vLsUyv
LKRGTbZnYdBvwb6ZUu9T6aHT15YecOgv2KfDNXT99p0loh8wA77O/w35brvuxnLi
MOLKXDvMEDOz+5UmWCum2k2ToLzohsTY4ClTtoBdWpKHznjNcJrWSMjel36ryX07
R5hbtA94ZabQCmkXMfoRUYGZ1u+rsOWPyxGGI4PA76na6dFYs/6vDJj3Ht3OEbKO
+aWo8MXeUUvDBJQDGeVH61VsPyriMBWoC1DQ0jf54TlZ1KYh3CMcMyiAYM8gqlrB
E6zuULZH24XsNv5zGYhoPoBv6ZT3WckCwvb4zCwzSB818E0eX3F+hJ+EFKzIx2LU
8Wz6eAejpO07bimvgB3hsbNVD64VUrTdoNWA1xV1iACu9ITgAZoOc3wBqFydIP3p
SwoaVTNUzDlfsrH9CRsFYyXvTAeRHwD46M9bDvX2ZJfjlSsoeTXFFdWOtLQI9+1M
fjHmreQDEQarRZb/eWSZTD5QaEWWo6pV49pqcUteNg8lI899XI4xOBrJfrszAOWC
N2Q/tL5ix4A6Z1hyegerdaRWvEFDxwpJOrdPn0M9jbTdh2wOaQtHydQ9+AuHzJh6
KwyyhiuVOQODWpvhUHwIJDcIf8jRjbdHxXuWSCHkQstmH8O1kZGTmRvlAQGP2DIP
Umtk9VlHVVtY4oYRGdWqNcO3Uvc+gRqkSnQlRf6Y8CupHHWnK9fNRi/AVpswq7VB
3pWlfoKUvrP5zJI1c9OVs4ce+BjGW0yjGcbxGAa/XhMhCX3/ihz+If38pDasVXh1
0Oj0VwcotLPTRSguououseQhkws7kiwrETPA+bTA3JPrMQYiwm/d114GGPE9QtLm
Y3PYoujM6k6ah2vNdvMX0aQMNgiNhM1w/Oso2DHOe6WYPQdKHhiUVl2bml2rKJ0a
oZYiN1xv078e3hM4xSGRXRmndCF9NXGYVmiFUW2qXaT/gNsjpJ5MQPs8ZgXHmx5e
qx45ZAa7lbBTQwbptJHwXGAPBT8cAWrguPNXwPnAdq2cLgePkCn/qwivzU1VDMFZ
pN+Vonhlus4A2vPrPtd7D/2wnx8QQkn/yiWyXi8fL4chhaheCBRkndGi9VNid4eE
f7XKoTRkyd06vbKEfm2CFhxlx3wlfU/D1pU9J2TqdAtXh9ZrqLUjW8dpjrWXdecN
Z9CCcevpzS6mAUq4AImQpfVW6V5u5FZDGy6Dnpq+tf4Jy77hoyO7a1yebHqtXvLK
NUo5rFyL/R5i+EbEef6pqD2KsqATL/dLchhiZ3ykoW8krVKh12SzTvWLNgVRFpih
pnaq9usZO3p6wQFmGBupHZ5j9aP8UQ/4beVenqbL68Mtt1YCVlUsp5IDgElaEhd9
WK9aAenPhSgZzlMNzCJqfdtNBor9G/lDZ32gXyOAHKiXIKlRpvvRAUjbMHZodAM6
f87/PNbCuY2ytjmhDZqt2+M3YIK5mQytWHfOEVrcvxPBYfV+lsVJUCRWGaMZWDY9
uwOugiZIQJHZOhJNaMGxjQZQR0g2c14+EZwXHo4klv788Rh7d8iy+X3/1X4DNjXt
d+kl2Ajs0BzifKiKTwR8q0SeIQ8GBntF8DhabrfwtKkdrdB3lo56NfS2L3uYaG6+
/jrXPG1LaaobAdf4oupxFWkm8x99MYxC08H1nj1A6rJO4aEJGf4f8ov3UqaGaiWP
qb87bXsZ2gAMgAkxnOadeepWQbRqxBm6XpP8xyH3q7gjATqulJXcmnqIqN5h+uIj
rv8FVWHvdh+wlY0iBkl8UJdPXIb+nNXqg4Vr6G3RvULPqJICExgRNa1l2utELqly
jfqQCuLwVKwi9O/9fhaDe2o1J1e8OuEgjkPMXQW3qSQpMfU25d9Edr+9FFvz6cjk
kjJmEbYvEcJCNYcrreGfk++12NoWAwGsTtaznjCYweG7eaPfGMuMDFk2pPZ4Fwtr
FV/SwtdNn1e60tVl0rwcbqMPJo7pqlLyUIRzHQp/HUT6JnB/kBi3vjvHQvMPKxpW
vj9dCneRjROrOi98M1eE02HOV67skQecXLApC2j4HPbkxVfy5GlPqMc9mUksUgEC
QGD3U3lQPZxEgRXPJYccDnuuR8rc1QsyUaDKrjaVBhD6B6lTLEEFqb7Bruv+NXJN
y63cyUHs8fepK/RlICeQIyN3c9/qJJK1pbeq4Jj6bbiVYOjHAJgNo7thQxLowgxu
+zj3hUccRSZTLbqXiBsP4YGZBDeO+AQUbcP68BmiXr+qljf30h2o6kg5baqKxsoP
zE5IKDYThU0dPmxI4xlWmvPWw123Cy1BDSKw9o6ZbpgndAr6KBCu1hPzsngTXqnm
R/IlqObuYGAK+45qcImt5gNpMF0YO53NVtyTwwkuNwHJlH9G8JLo30X4qepH7Lvc
AtGwyeXkaWCwwL/dsV3uRKEXbKw9MfbBT/elvZaAuRomAQWDpf/B6qsCjAsLQEX9
MLjdluSPzKvNONAodq4n9DeAgl5izwkzFwohzryTrx+q6+wKpZZoD+mxXyTJ6C46
pfWASN7O+d0BZhTZ2rylZ2vFVdBCSRJ5yaFKyZW7Ai0Q5a4I4UJT78sCclToG0kZ
e68sgBRLn5g7846mpp2kMQuttJpCi4EEhZEpd2VZUy+zh3FdSWr19HdtQ1Av2IZz
ouhjmDuf5Ep6aIhJL3i//0DxVObVLaFdsZYfMg28Yzc3wDf04eEBxH2hWU1Vfuon
bPUF3V4MWcAMWfSbgqWP4M5hlYr/GB+0GMOVBk3kp2AkYUD0BFn2HERsvj2Kqgo8
Yq+PUUeM1pNtNxbUWonPKPyy9f5zBPWs3EdyjEo+Du/JlOmjsHzxDzVRvxpRk4xU
mjpjeAnHFJpKm1Ft6wipgXD4uCqGyhbvUaXF96TDdbQiPaosGzzIgq475WCk2IsU
gUNFntljql75h93ePljfOZruI7boNHjoCsQ6O9FykHKOgybGwzv5SLsr2KCYJ38h
BApKKICaDwggSj0wmwDaxIotopGL2zMDIttYq/n4nhDYgwovAcogpheLXGYBgCUw
tD0v6rk2Dk0LgSuiOWhmp+Q8/71U5X5S+xlIJ5h120NejfY/TgYg8xYa1OIrqLbP
EZ5SY5sM43pi/AxZ8plOfMsdsz19CUX5UFrKJDm/CGdGs8EIipkUmqUyqBkB2bX0
FsaKqXoBQlqH7nFa3nsISH/B3tkGMjL4KUovr44wtDP1K/9mmlTW4wcloKckGKj4
K2lm99J1vsjLKX/+aO9QEO7PSTeo6qJXPhbF41UM/uHWzQZp5lyRkx6iqQW0ln3P
nldy9lbf01rpbqt5MUQWyfhL02Oq6kduYxJmAVNC/g0tU/4PhCrLIfsVW1akwxf+
iINtYWa+xFGLlemI9WwLKDvRQiTnK0gB+aM7CU6clSUs28r0WMvu3/KecVw/AGVh
6wXqkSYeXVarrMwJVzaHhGEPROjBvIHhL9WLbcmLJ/xLux6rkKPkc+eFrO5CUUyP
CxoafTX+D/0+7Xy75mLL/8Ph40XrBZ4UA7RK5WyWHxg5AIcyz46NMD18+9lCZT+s
VBKNa21AyIzk8d0SoYiWbpku18taZ2dEJ37HnVNfjv9NZESG2KJriLVTjym1RRBW
2bA8UGF7W25JYp0MLqeZioxQ7e+a7kZv8MhBQPenqUQTErjfhLNyEjg1T9OILpI9
sHVBFIOz05QnuVwBV6GEJxtVylzS5ZR81+DAQPSWjZldRgQAbJ+nvFcvkRwDMYjc
SnwU4caHlETFYiee7uECA85PEYOohEND6BOdU5Ny+nIGzP+ackwv6jsYrysgP0TB
gYxi6V+AytsBML4rLAKV0PrzvaPkrxQyRqmKUH8CrWnEzfVOttCRzTzE6UZeECeY
9YToxT62TLjICFopcsxryonOCw08VlvWxhqS99pCjHaXdXWCKbf/AaUuJZqea1ms
zCS6XLPtIGCQNPuBOVVniwavkYoxPQMx26kkfshUiZ5w8QItXomYGgE/kRrywStH
oNGolCkQNUq+4dZEXHq27sUkV3XgmX5lOA7VBpMrcjFlxrex6AsIlBuxKcBFD8EL
D87FmqxsoOtPeoB3TnqUQVu6OWDgLTL8OMmqQpAo9L0oTJZr/qBFT6t4Qwx+UW3v
K4RNSTzN5RbFAmyXXvqqxBEy95joY5B9PSHxZzX6k7tKL2/3qLPDsn+g3OU+xueo
9qCPgz+OL08zhyQsvDm1S9jRXHdjW5zCw06OVQK3Z34YmccRTUn3G/lyCfA+Xvjh
SZuR9zL7M/P6l7+KbEU5yVKEPlvIgz0p0YCH5H+gTm0vkgL51RhIPXB7qEOwzHcP
Lga02AOeZR5sGw1jOcBOLdx2GOtFD++Sw4NLPo61vS8VVqwlhluAWXUvUVfHIjkl
6+dJclEELik7AV9wGL9q9tfYkfCJP888c6UWCPqyi51y9Eta4JpDE4pKhsP865f7
7zoFrl2m9d4hrjayrRlAYrg2tWQE9SyM4qWQkgcyd7wFGesa78gCiEGzXMStU2IV
yGd5QBdQBFTHavCAlnIoos/c6BMI1bz4ugriOsw86AHRM0wKcI+sfzBgmIsIRSUW
kjF7Y5QnU4cuInlct278veg7dds/K3hmMtBddgiLJCO+/YCZMNllkrSwEfwsbsyb
0reyoHou9QXMcYlrwd2S5xeCsEm5wfqiGyjDI2UJziJk1RVZaplwhYW+3ijFIeQO
ieowlkUg1ZP7zgD0jtQFePGWbMbMr8w4sT1f7SVAI+Q0XSrX5cvmxvL2fSNeSG+G
CmrCvp8djCeYuF3LpvrbEO3+NOE7nlJo7f9Mrgx2eg1xk/xYwnjuhqGXva29DAlQ
Vc0UL0VOrbJhxuS04IYS4/9wKSw75zZUr9H09qoMido1Av/rD7fTRymzhMlIqU90
vH0nQK1RT3eDZ3qhXYExcFfgwtrGIyeEgduW8BQO5KAhgLj8xplSmJPrYt/J9vQF
ZJfQNQh/Eax9Emk8CFKq4QTavhkqKR4lRcRGWFAk/On3MbFEXHgh/qPZzXo24YWF
LTzNkQ8oYoK4J+fAR5rC0o5lo13Zj+KMVQBMw6f7WihRNBthV+YfCeWPSuwSY6Bw
dY6D42YMdCXfE0mSTh9RUzOb1qgb3EJ6ZUBaqDRJW8OGL7ol3xPZ3o6GUabDcpzL
fLeBFck9f6pTpHwG7zhWG+X1yKzpbYKt2pZcsxqIU7dQLZW60LR28ysUKicwclfs
u3VF/KAZVuEZ0hchqJbeR7z/BdpnKC2XCmFr35LZC/ONV+l4p5dTBJ4vePtVt2rk
wq+zwFCaI5BFjRxPgYmYMlu2zTIt3X2BDsHPA6kWVCCgxGyuwAQnHb3Dpei2cdBX
7iGnGlnWRXv7VeNoaGYZxbCf0vWZlum0yDmEcR/icqQzLChfB02VRoK3fUzDkqpA
3CRaVhsAmD0/T0aYqisSCpX6FJtMFB7On31BKWFULGkDFSIKfElQZLZ/32QV/fFb
ob7E9SBpZGy1GKYJhk9vPc7u0Zc+XpxeodGvbUl7aM5OnNn/BTvdEijzsb6pw0KT
l4f67NAQU2CSx/Vlpcmg7/zCWu/+bL7TbAPcccM0MGFGvlQxwKt68Dfwa/yxRl47
KwRGYSwk3bsMaE5FCovTuu2VNAR1LtaTesDkr98zrW7kx5/0dnD3hLob42KkIl2l
2oQ3VLumfUZWIl/8BuhFGbsRaaiM4kVr3cWtZ2WZmwr/wxXMFugpH0Y0XWys75xJ
xc0M4OMUEPd7HRg+W2IOqiuN4b9z2bzBSVhw/TNOeUFrD1oDOohyMWBsbb7tXNki
Bp9WEhlwtmEkveNEvPFNhCez99vLsvy6rlY3p1PJBau+sDQrePwhJe/yW+USWyn2
sKwUj+mCWRgvh1CNt/vMOMs/OVOS11mKryL3mEugl775pd3u8Aa6AZYW4GupRRxd
9T7SzdocXDL4th0mA+IwpLGmrcCW8yY7a81W8LeX+7CZBmxTrT9743RbSyEOylcX
o7RKoYqOomiy4eXitAktQOkUp6HQs6J87GAZEriaMp/J4cYZErRNyHQclnKBUPb1
PrDq4OBNZ/gqd+lKL5rl293s1tMwqyXoPuUwkWDilRrYGVPnixHFShSYmd/M7kly
67iLnMTKorhiqYK57Yf/JGuzKeSSZjc9QTv7/UKRG9TYgYO+KS5mEmZnwLqAeyyQ
cPmF8aRnPRQ7LRv3z7sLCzRp7VOfzidUMfVmqd2yF50lP1wVVBnb2cCZJwwXqG1P
xOGc4bo/T4ZIu5Zb7Yv8DUph0O3KLhFZ/wlAaR7ponM4LX/UshZJ1GbBiu98s2Bz
H2ljkkUmJrduTKQL6oKvHws0WAgZxXLmyQIN7nYUmiBjaw9thdyNwSIOzpfD2Ok4
gcfcKouvZjuG/e8KfvnrNaJjvOi0O9Ys7f3na7iUxQibj1P4/o44wetb4L1dYvaD
sqhZ3L2iem2CuGSFQb2nvTcg04FAoEGcA2BZLL3cKry1OmO1T+j0FDcy22iSdKFb
K691y1c7nPF6u7Ja6G3zM31iCIcr6ag2SQUnffg5pJcfAs9GHEwzDisqMHTWJ8Va
mG/yTMNTdEpcFD7QM7JIhGz6+KEOEEGm0n2EHIlL/M6qm4RqOVQ0k80HQty3IN1W
pKDvyrU+M7hlIFkaBXrDYg4FoNkKYai8zk4wfDPPfC75GPUFyq+oNB244o2NoDtF
RaY7JqCWsagZuWS0xiPyRCbwOB+imIuIuiieiaNNW5bnv7u4IOnwVMiPNpS3T06h
A9w+oRijNq+F9V+5HyU9Jrr07ME5Cd+xZwxWtOKxJHr9qDqjcsVLpHT7OuhsgKm8
GoN50fjKif6f4Xtg94sT3DgGtyTKhW5oEywffiJelSM3im3+OA2S1Zf7GV7GbmhI
HcIMeSjO3CFqsKyQhlrTVFKXIBTWknmwp7AsTvYMwb9T4OkKBbq8HQXC0sQ2hs8P
X14ijI/Pl+niUzPA9D2nBA4D2Id03vryb1NPHIjt/fyIcuey74ScLx5UEDRc7Vo8
L0B+9qt2E0i/onwSwyAnPKPmu9FmXuabaic0jmpJEF36gRLRHx26+ljkOklbVs1D
ln64xofnMzO9tUQNkXz8twT2tZ/oLbrlDt1kIO+yoaVY1LLgawa+S0EzaAh/6h8E
DEYZ2GH+RWrBjfwLI3Pil/ZNibyDzFNXgGR8gXLp6+PKwbuqHSviYjesHq8972lu
M8/MYUeeLzA5QiIdDdyu1iqqnWsMHWwQIGe1HRmA6QipU2bSXsJlxt/yX1RuGJuE
lX/aOxMQhvPkKM9nvmomS2Lh8SFuYmMPXz9kkq0MhG8SIaZlonUI6uHV+m4kcjf2
3uYwlmrfoijTolUTc9+xL0vFDloGJOks9OdRr/R28VvpZ/qdUI4LhFgpF8fT4Nh5
sLZ1n3juZlH4BBLb544iFZuv+BkZm0NzzHklh+JL7tbGD1o7y321DyyZFXYw7gqU
vFe45ROxtaq7s0pR3rRacTrVYVlgLDYMIcFQZe5rJxFSGtb/YQT5XKRqRLsny1rQ
ctssnHWpwPjxZ6pb6j1R7Za7Kx+bbCo4fkdT92MPxEcyPsg49vCF6hOBVAW2AJXx
pOC5AtgftYc4katlW+sKxJqDW82m3QsLaM3G50JKH43O+Z1JS7yy6ss0ndNKMaLo
dV3C2T6iFGGw9APgiWFdzpDg4xoPbcU5wF9SZcC68minVfO6gW8CkJ9ng+vGB4RX
ewy2znXvpb1rUOfP+5aOGVBqJ2nQGSPZ/6oeX+8xf2wWHI1EoJ6kCNlOkmFtlYv/
SPN1VjrNb05D2gWhC355c8A7GmDZcFlObZyFCPxhBtMRJXdlaV47s9YNv0P8dqLA
jKeU/Eicm0c9nJb4enJx51LUuTpTcaT4ZgUHqCjRSEhF9ego66pRk5FAoJ8LCvUP
Q4LkyF8jfXYB9tEu/TOcEOSI2yGLLy3J6olIUZeKtuoZWb0ICRwtvQB+xuJfTEHG
SYHLq6SOlJ8mLuKDdhcMwZCETfoCvPqxMpl5VTAXFWcNB02I7+xU/1EHd6ZnQioN
Al256v35uPGsaKa31ywifQ3tywuOB02e9BB8bpOlw/ZNHwHIWav5eHgTAMmnyLhl
FxF85r8IbW5lVuuD3xu1eBR+xg8rwb447PHidT+4DxAIhkHTwgUJopEAUQRfRyCE
W4Phjjqck8i4XZ0s2/KChi2mAesppLHqUgX8brxeR8jx3eS0QhZ6yoaNXZFY4YqL
mkwZYVvtGwW1SQysBvgVc2AdgrrgEl+stx1BI7ZwPWKCokSlxXgol5CbOsVkhh7q
ofPf+bhiJAnVQjmErzdPjBMaFQu7j2ztAfXLK5nfMO2wFunvXqM2gjf+w+z+MG3w
tIa6bPycSuatlYDUQLFCHBvtsRU5A3EbFo/4X+FWJxcTtz5+InRDnLIWNmcQiMy7
geb8zFUZTG8eaX2Csv1TIqprIoE9YqGU43i1sTXy8rNM0RfJqMP10qUg7NIHCYqQ
7yp6HPdJyuTHgfgcjmhDIYTISCTzH87W58s5yFFJbCbTPuLKVuj7+EU4VuYxoh6E
07bqZPLfmcS1xY+VwrAvC5AeutmRgh7W9uutEBZXCmKrDUswTClqUNl/Xj6SEp2n
YrJFe2um0kTUBJfzQr6su2/ZLmyw6tPgvDY4x5Y2BPOqvjgIbQ71hkdQ5AWYIAN5
j0YUeihqtviIGR++NesrYGKA9Jg+ImEf0BBk9AbD9/O0rDLB+8r7PMrW9LOpPnzc
w0LIYLvFjLrDKK3goo/hzpO5OKuzhPR0d29gHResC9u5OC++6pWdHOwFbThoYpe6
WmrrzekB7Lewzu9wkbyFY0FPtwgrTuvRlINZcDIqXVIfJclzeVHgjd0OZtBbTJLy
xzyCp48sYkwjjjTnyOn7HGv7XLsH6BpZSvShlylSJOgRmPssd7uYbtRBynmbnsx3
GZu4YjabTl1W3kWAu0mOPYcdRPfCJYQ2QHRZGPIupHvwHylPz3WwV306TBXru01+
UQYs/E9+oxIwS2dszb58vrHEsesjl8S9oZQxW3ZAaAtrOEM03uvdTzC380PP05i/
jqCIVTqrJi2akFz5hAYzRI7YmWYc1OmMZeZP90MqrviGARg3pbf8ulG/y35KnWsI
999jV5g5ja8bcSlhekft9DCAvQKZrRS0/L5LI27pWrh+FNdlZ8rwaxYZ+/TLM19d
any0eSyn6J6RyPOATjS3IjCZ2FfuVPb2aarqXtIVHjjC8Td8wB7hzapGx5X8Sbh7
TEcSvBkZWov5F0ocA1pR2cv72H0l13BjhAy22VOSYVQl3O1WipQ2YOvyve18bX2W
wGbND8dzSNVvkLvjjaVP2FPN6VDaxr568Rtir++P+Ul7gThPaG3UARTpP/LGbxWf
8Nt50pBlNooQ59uSuAjNXXrKswa5cdfg6xY65lsuqcFdQnphfQgdotYp2NvWxLq8
reXnS743CLvQXcu8j5msMWxVB1QwQvDRCh12cYcBh9CziqZd9SsPbKgkNqUQzkgH
Pa63M41lRrSEszBKPT+b6PkpAQKTgh12HF4928N+d3oakdFy4SiYYe/lYpydIWOl
ExBMLAL3rNXXfWmOhx7z1CQVdhY8zIbSsRJNzCtKqxZ8GDfQV+rKBI3uuTplHLjo
Uq+l1nYZTzPbzcydRIxjYSD4ZFi1luZrSgRyUUM0K8/qeqSSqwQkVIbeNdBPzEkO
jX1oXCcwFnfdg2K3RVfPkoXzlbyLla9fAVllAoBnOjn9aAUFpjLiRL7IkCY1ynsh
pN7FBSAVQeD6e44bMvd3U7y0Na2LKmpB/+Wt/EMZQME70TzQ6UQB9/LnvcMWNC1H
ETgAFE65XF9wJZz7zWKZTlt5Sw/6/TE3SjRTIfwJd7nU2Hfpd3Syu9v+9kAZdJ/a
6psR3fPUn3ZNDN9aU72fZ0o5ngpmak4KtS+oW6qhfacbanLQE/5RfCqYqXC/Keek
xJ8fInSo8td/1xR7iwtIe7kJtzQMydfxpNEoYbx6Ef23rcB/3+X5gLS1FqILDzxC
jdh0duN/9JKSXrSRUQm1OyEmlweSgdYw02rysTAYzDEOPzMKmRKGB+eQEY9L/0Qq
EAKr2TY4iPONSg6PrbYcZmFQOXSDsd7XhD8UobFOqjU9SeRuhXzjEqgN69yNCWDu
ItDVSK2N1/KYjiwI0dR2kfGKWoMtbCwimySM90N8x4bciIHslouTLGX3g7F5DeeO
Q/WalfDHZ3PTuJuwjLtITsP1eXSrEumyuGJxVcy/4hm4+WEKgwudxyzdwUNfMsG6
VaH8m9HTELF0OvPl9nYQJM5fEUQtwZ6MEaSUmoSmNDRzNeMIyzR1jvLMfsP4N94K
LwEsd44mg6pjewhGgZrnCZCpQJJSohXzLkNWm/PrcNhBqmek0RJz1DL66Jul2I9Z
Dq/IDR2NMkYkGrT81YIQI5NbZWr/pNKLX1nAOVNUsfhXCaEa/Ha3ZI4lc08jJcj7
oZ0XbNpOf3oeUDTIRbs5FJut8w2rD3O25e1Dvc+bX5KMNpKtcWfn89i+fgW9r9Od
1iQiqWcXLxjkkLQSYIE9JCW/AqoqvcDCJGrMt3W9TtU8AR2b5nw56Eh8Nc8U3sm5
Ojs5khCV0gKzZHa/XCKoDkOVBnOUjExs5htZtjd8YlfPDmcROLZgyfvwZj6h1MDS
6zZ7AsJUJr0SGipQDHGA0hplSE+B6zor7zu9nSzDoYHZ5Xa2AHRVbn/AXuRJ+Iup
2W2LmFnR0Cnajt63pDQMxA1tss5TrVdqf9Y7kvxohDlCRQFxlsiOJvrGrvghubU6
sVoLbMoofH34fSb4UgrshpBuaKdsjmyvF8lZhZ0SSERIv46bGnW1JzvWTC/lcR4u
GiGKbvQVOSOjAbbiM53IvufI7M6t9KwqKUZI3ye3UQtVyfcAaTTw7U7SoWPMIkuY
iNcYGzZUVyj+zDIIwbMpEIYH83jMxsnseFrPmspazIck/r8D4bf4eAKuVxsmksH9
1IaRwMI0OPiw/X0lxIeXd8Ty0a7mWPLpFwCXCO89CKtFiN7EVbLgs7214qqSyeW3
RjrncS0LTROZQIk3g0HwzrVuTOuCJX9BQEEhbhxHCQ1pHMGO/mRPtDMwytpvrxqM
Sr6EGS0/xKVZnsDBMrDLFDN1ACmdxtIYPkuLFpcUbON8AAlZ333CAKUxcr/wAaEZ
2+O67EVCra6T9q+gqsObbSsPeXtMv+WFe1MDvUdptjT4XznTqJOR512I+aIiWJEw
q9OxsmxlnZl5Oy30wUYgSPAVDhbliSd+mge72S+B5O3qbLeKGuNV67qbuzzOMdhQ
tOTZ4xFUFMX2Iw+HMMDIZ2qL5IAiENSNaHlCqDZBI+JCCQ5x2Vm9XLQJBXBSZDqW
KYIUAITZ8/9pCgx4ObUjZzK+z72X2uC0SFJURS9grpc7zOXTQoSzvam8TtYS365M
ZFmNjI0cqhcy64IaCxTfS37xvVZIUp0flQxxpA0yuOalJ1HakWphyhpiDi+xHq8C
fjAVCfXl88Wg5mjmVAL62Ezm65hF0n827wPj95uqMzCp4f7KBDNem5CZ6+CShhIc
xcN7LYXMUpRpZ933+YyCEbXvvna2GaglWLfuv9utFYjDaRW9YM/aSPPuAmfDQ0FG
JluRnyszd/5F+VaceZI5gdfgTxs4yBkPZobBPci+bN9/CeV92OgJL6PeDefKRzlz
httlwxWcJ2sQwMKBIN7Ih8boD/t2PR3BQm9TMP988Qv77/v5uS04baezp/Ims08G
VoAhxuDppHa8+WCMSi5364GdJZRyqa07t/g5TJIrYA06ZJaei7nLkn/Ff3LDd7bK
WFsRBHAfvuT6wgpYd8FHgnb0bLZyTRvS7Bj2sg87Gd+hq0bR8FLC7MsDa9uu9Ju2
WD3zFuxNAtms3JyScbvP8i3sajOYNESm8WnwZO1fAoaoxG+WJB/kSCEtBd/KX48v
P4V50UIw/uFZeub0imqb6MtVBxyuca4OJbgt6VqV6yOZbvLSnRIb+NYaIWr8ClLT
ZGVLmSjKSf3+mVXRVwH8KIW5JaQ+GCm6OHjUG82ydE+yh2n9oSkjgG9AL1jzt8r3
TzAAAySuOLds0fbVRk1gxJg4c5EISdjzSBhTHvgSgYIs/Izq/yyOB6rXLeac0h/5
C4zf8/aFGnIxpKHE6qd/M2uqflbhvAIj+cEa3ydBzq2Xa1JAih5kwM7i7AgAIkND
RbLcJGffKeoEXnCGvSvnd4TsHoLrTC0WTl486PnTS5A/2iR6J0QNjxdUYgrspr9q
+vprDj49e/gvdXwrvscqEsW27D0dFRFcKeG072GUA8Fd+o+B1EcpvJShdgtmQwbQ
JIwFKSUODzysVd/vAYr6qRTOWmDS7fMkKgTLvBQuhXTxSvdEHlIuhdfNRTh0wIPQ
sBpZCjZw0zif/H16+qS76bSHTUtfEs3Kw30Mqflt+RV9BbeLWexGCTnNb6uJnPl3
mjiYUWbZfzPyI1TzRSGtuXyykSGMMPrwZNaMlT8L6fD4l4kMFXnaw48YIc3G6T0Q
27OlJoB27LyScQdwlJ0R/KVNIhvVm9DRTJ2qU5W0wft9o+dbrvztzHHELFdMTPkz
LTKVOEA87FpOQcW/DRxT0B63t07OgYX4ypenL6e+kcvbcKHoYyQWQljFItJEdWrN
WBN+0sExyIdR0G08VIiZUtSXxOm6df7aTRSx0q+dXG2VMmDHP5oNo62lcO1RmKIF
UyrrSObN4+Enhhm35et1Qlpo5ocnhhsnS2AXPt20bnFwAX8kP8zuL16UqBPIvlvW
/jc+R6IV1N+9x5z7x5gTf+EzrLw44/p/dsQFaXctnC5GD9rrhtIp9zcqmHtr1zo4
sX6QhtbTChaxvTYuHCFNMfbpPiBmolWQy/ylF2EpS/79Hc8tamtWj7lktEERF8AV
COau7RtrvP+0YcmDktR9B2ohRp9awvKJldPC9VPHAUptbS0xHBFtjPX3inBoVuve
xwKTNblam4bj2Zz7SUe8DOtiOea/k9VnNK7KqVBxfKAeCyknBjImJClmPM5Uox4z
4r2aGKbc+tpHq2i0+aut0IGcqpTJ0vm5yt//6w5hBUSRdd9uHoYjk9DTL7JsjvtW
cGA21qq87lfIP0y6V1cASVhK2fiyBDguB7/2ow8a+sbatEgLJ+RZI0WywDhO/GR1
ETL+ihl+6t93kgfsS4H5GH30E5FJpe+q3414qsDuKiKMRqM68HwPd7OENAbLfJeG
Y7waBwQuNu7GZB57T73ilKkFpv5B5lvFi2STJcOTdpxnLtU9p8lQ52IhVECnVaU8
y2uSQLpserov1nNlo6gSvaZ6z3gpylVBBZa5pOY+KJbchyOMyIYSTCWzwBVIVVnD
wsppzKDO/jcn3VWNYO/57QkLat/qrnE9zHedOoU5Rti0Kv6P4JBeWq4frnePHFIk
/hlNq957Vq6EqEa8QqM9fC53qb/mDd42/q27j4NWyfPaw/+l6zRDDdZeeZBCY6cx
m6JqB+Beitwy0ONP+MbvjgvEZpH5G1fC5SfxTYTKGzXamhnoTlV+APCQXDKzTlDT
4/uZ9yohO9FW4Z0t3Ebmffzs2p3NGzgnd6gAhx2KjbS4PO3XryLffC3bVWXlKt0J
mOoQ+OwzyOBU4PPXD9v0nNvtrXrDpR7jt90pUB1Zt8K1UdawzL81+r2X5PdGlctR
i43V5EMHr8+Q3vdQzQ1tZw21BJQiYbJbDQq58HBgVFsowe+tLVnHGyLAm2CZCsDy
Qhe21XsmHQJ1J2FWHfbckKo2npa8IyL6Uy+cPSIhn1pAK3CU0Ay0lewSh+9mwVdg
X2zhpnzZsssNmV6fD44+IGgww76Uu17VoOCXlReWd3BtDkMHuvTXbNJjICArnvxe
HBJXWNCNVQttVL7GDWiwuMNsk7RAjGN9G6DepRM9hLvrpzVQu55KuA95qrdyq9G/
semzBmCvKlMi5t98kBEQ7X91rlGvbHx69vW/HS5gJvype87KCWr+T7Bh82jHlkhJ
JJg0bSd6qQXwRE3gqQYF6C0liWA7T7PLRu9dVIowpPxuS+mWFeAu3x6IVSPKetBg
7misbk+HAx6xQBDBkg7Md8+/sJO/oIDwr7pqbT/58LLXATH6Gb1Yx+vklfFK+01l
68w4C8712lV4wamIgRaZF/s9vWLGh7iUJEXJ5fHwEsa6HuN97X/zDXU0adeunHSJ
kSalUqZ2gFhF9VxEuSU7BCY80IGvPLSbFqEBzDJiFncvXL2Y53ehFlM2MnQoEtmw
RdIuJzJGv4dqnFfX+RFLncqgmIfMbYsyQejXRQ4FcUVLnftQli7QA2Ek5K3oIjRd
V9tlK/+0BLolQQFFr4D3kf07xytzy3soxwhUvyqKQRRBA/PTRDXm02hzhQ4/4DyW
mHI5+g+tzr7G91ztyOd0/8dLLjZQkja2sl2aUw8p0CQT+Xp0pU4K9Tr/J832AwE2
Mj4LqgnPHl8L4HMw/QO3mJu/S2ldnqYfqW3W0m/KG7+EURs71ks2+XDVDLiX1yyv
p3tVXjpaWYwbfA8/wj51s4Qo2Y6HH4Ms5u9lhMUOmKNOALjjO7wlsKHc7NGOEIw2
zT+0OpP12ZOJUI16c0PdKPq+nrMiVjP13iU/sA3jeecXcHZgFO0WQ3h+NMbDLYsr
iirkGWu6BdEOMYM+q+goGHk4GY1wUQe7stqWGyZgNTPmk8uO1+eX98wWVgVSNq1u
++V6T0YeMi4k39fNOOF3cYhxDlCauO7nUREJi+6ruhvUu5dnGBzUceIPESbKiFOU
WhV4QtTYnS9uegykYjhFiT8sf9SMAvm4B8sZfy4A2hvHGIMXOCQSN3S3woP0WZ3/
WfSufK3fRn4ny/Uts8NSLglHBIb22JL0kiMo+7PfVp/6tzRspKhNw51qmLKa8D/i
+7dvxN9ILdPqMsfoy+EA0ysZ7f7JzIzFhlZQ6V4pyfwkXyytg/1xp3wwlyBBSTPa
MAqVkXJtZoe9pyz88HJoWfXvaf20Q5B+xoKp+qP1WghgWXbCv6+t7Apbjx93ZStj
vo4FQeOTe8Dpcjc8f27q1EVGhw5a8jg4Nr/heOMoVzFEqol1bXK7oNCmEc7WfMDy
FPdkIR6jRZRR1RDdM/t2erzzvoEeQeviyYd1TTG3acaokF/7sYk9YLhSZMJbn51n
5aDp4ls6Nr+JkaHVzmRHFwi+Mb/GGkKzDqSg09Ka9InonLZ8eTMkUr+rhUUuHOvD
0mX0iCe6c2juW6YSPNaORcUo4/Z9Dy4KDuNB+r92FfmLZvI4DQn8dHFUM1g/lLkx
m4kow7Xor2ZKiZRAhSWCdd1uch47x2ZgvmCUI/8EA9o7g/zaEWG6oOsO+iDH9/di
V23I5YGfLMbI4nC1aOKrMgU+UmmMkQo0YbMUWO0kzRE0kMleNA+GtRL7i1mDQH1L
uyOwMmaryDTxfQVNla0LAxJtOP4xOQM8v+MbxH5TSwnIhBKWzWy+hmMYoLT5rD0W
OjLYUOqDsvCni75E13CN8Z8UTrzJqlTXzNVVHyiwBUW556rmOYJAPhYwis3M7Fjd
lwJEwzggCMtFloiaYzz8/YlOZZrESavXW2I0+JBY62nL2nnatcK4ekN774pt2fWG
rwb7W/19sltN/oYraet4ri3OsbzpPp55QFZlb7Kg7nxiGxlslpdamBvilELcuEsP
MpnGw7p5gOMMbmuG6WGXhasdyTWVN8Jn+aJ1Id1Pi3lTV8X0RagMwRDwv9qFKnQo
0Ic0Ic08JtEqI3f1SqZuhSfl4EfhnwahC1/W+gicGph86drWt6uUroNRAr8JZIiy
mLR4wK78XM3qB7pPhOvlguen6QjtTZuGZxJcDfz5HNh1IICKK+AIaO+9H9WWzEV8
D0TD4GS8DuTUdDmW4xF576VHSHAYrS473Ve+n4aBobpBkxRjup8Sy/QYcDprKdqF
Bc+xhT3G3UC1bw+eY3/ox4agdsVS3i4l5WuStb0i7Oh0ReyMUUs6WeyOm9KGSqMA
CA2C7M64QkKDEHHedLsgXOQcOVnuI0CVmzgG82irl+MptauGpASxYTBje5LJ3Kv3
7GUf/Gm5Cn8tEa0mU7Y+1bE74AqYrxb9eky5jtBg4DFFje8dG4kCIc70c877XERE
PnQyuNWNiLr66skzELAbyDH/O/z059fXaK9h4apXbj7lEfINs89kS+lOH6TncCLn
UwNx4Dm5/27Yc2pfbHQD5D/rFFd9rBy98XFivSDV7yL98MZ2o4UW1lLWvU+RpZMk
97nbw05njyorlavOtavlORijncTL23t6M6uT5VbSUMWej2u6cbMbdjrBpuaQOHw9
eLnrjZLEVyhlHFoVxQpm2Tfj5+/eJwTod7699hq96J/o6Q3NM58XxqRYJNCpeSMY
rZwJkGMaFTDNIe4HHasLnx87Pe/svCWlO/UUkQ4cMapfEoxqiOxMmBWCxWgjrRZi
3Oi98rbmNYEBaufPTGaz9jXIo5uyahyUhTuwuicQsy3r3J1pMk/KxRUPMjbZiO4K
bayV0eix797XY0LMy3EMA4UB9euI+YdKtTZTj/ywbicjJQLsrPYY51yvpRNsMWgQ
AcQVOc+chnkM+7UYV89DVZvjMA19Fm/Yj+EGyXNzkS9CbTFs84yuY4SlWeea8a0G
QhXmLNxUvbpvWv0BqWl8+qoAsvJM9D72gipEv8vIRUxB6wODbQdUFRwcfleb7IG8
UJrGK0ba272C3kAJU0hOx17Td0dTUo9Sp0PKgtZYeRl/7rFCcK3JYnvEaTaUcLfA
aP83qKCvMoN5WEyPtQcrFrAKOwY0ji0VLNQhM+a3XPuFRrLQdCywclyeWaUcPhmI
4ZCVivpCo/K5m7nWez94kUYJbJpKXUoRHzqcEZo6d8HjQZcvgrADRpmaRC1xGweY
znT3pjepQVxN6PbqRXCpQx7sE4JZHztqH7bypLb7+TWYAHvhHkCQD2nCYpljfav+
j5rPAX8cJwGDRCoIR0upwgc7ccvTeW9Xy8tBo912X4a2WYbbKNYq4H9sEbhKkH3y
NtbCiUXPUIa83iDZjhfCCjcDMkxTaO2loPwX4iV7nYLyJwlJIYNiZYDzcTgzYxd/
KT+bxRSWjlEyzdt8WGuy0JOrlkgSEgplUnWCsTuRBOQcG/vaYo91xv7OOh/un2ZK
ymbFbjjrTaNXgbeiY0Y5yNlgWlNGxAGzbXJKqoPWnKd8RdttoMFdYB7zEkl9vjyB
E+Nw/P7ehghmlTxiviDAib1SDI+/NNTcO1ZChRknqgU5JMKJLyH+rChWSO5CsvGG
jZW7WyGe5zNAIjZ2a2MDy2eHkxnFMBqr1daqXv35iW5fqW4mgZeYxa/spu33IU/m
xlajiJe0hnh2nY8IumeNN+2JgX1B8d03u6n81eLHvNpG9slzEZz33Ta6XMfz6g4Z
MQPQr8XtiGhOhJhX4CILHuZ5s0M2U2Ji9KgXJBLI4cWEYMwCMaUO9RxYUG2fSidc
28EdKWncXuTINJ6Agz2Typ0wuPrDL97DVwpABd1IZJ9pFlgtK6QmUhBJOo/Ne3tI
Y6gilYoFgD9TbObnIzav2Vi6ENVT2Xvg5qUr+fRoMPpXY9IOueGSjcpDgf4Mk+E5
QnGJvNb8vlL1AoJjKkdRiSvh44Bz6rzYmBZqmIWoZftwwp9e7+47+n/2+G1bkCL0
3ZK4XhtorZaUUS8tKTSR7VN/ntonQhWfsM6XPmpcOo2NHSRZChaVmV3tYFlm5Dsn
HPXOO+qLVUKpgpDRJvW9/e1w7miJVI/Ov7bUXY7V2VpqOGdJ7TdZ70L8K/od5fVp
mZR5h1QYhJfm+USLDkySiqeq7VbBj1LCXxMZ+CMsjzXdlzjv6EPnCY+UpcENhEbX
XMVYKpwVOKq5TwlGMfemhduVulC+OX8g1X1wBUOScjf4WnnWZ1ywlhiqBabbirWv
Uvm+f3XHZGBkZCMwBKe3GnZ3bsbrYS5bS+/bnQvHRTNXzBe1+iMqNKnYu/t1D216
BJHwdBJPrmQrlLzixL1UPcEVYecX1M/E+SIJS1TGcvHVSuw6YpQc4cRewyLUVNVN
SEmpimoxbB/3x+ZDcVcgoRGwYqJVvot3hI8LP3KtHkpV4c7R+XAH53SO1fm5AYGU
stfkEV2lfjEfVFxKFTrxZfAXVb49duMYVrXojS3+aNKpH+XKbzJzmoes9rHzjl2M
RcVsuPCZ9WC/+4IOAXdnPMEYKhSMHfRheVRotOPg+U+7OnXsb9D/RJWzCVVzNbzo
X1ZCVr/EAH76zZ8EffnEjPaTHVke5wEVFRKSJv/TxR2WcU+rg20yH71vNQCxp9Dw
waugo1Q2w25Jj4dXgoo5VWRuONa7aa7/y4vViFon8h5lKEThhvcpt+l7Qo6HmB2B
CoG0OpU15W9TXT+KrJ8Hvr2nqYW1Gj2j5ihphjSCEfOjY72ZgbnuNF69kJPaQngr
cTesVmAJ4GB/II7hPFbXpuS/5dAHgZHpWrKqLwwto4xckScEB2QKsyxK4L5XjOh7
OUsxG5D24mFAgAwwYku6GzNFuOBqZvuGTPtYLdZRF5LY7EJJRFYKH5Osu7sRQWHM
A4IusN2EVn8PFAF1BNyK2OVsApkvOqBCWa7DJQYXaOCuPoeZVrjHogUykd6Vr/ee
gTzXGvOuc8ZFQvK0Kiw3RSgSBfDhI2eF/ZcXV6Zz4FW7LY2CNXwf1SiLrubA7bqU
M1xnxafsD2noPcZLT5GYHdc/PLK6A2yR6ijYuEX16lwxF78farCcFLRaePFGJ19j
yq0He5bECaI8fDyTChhPqI42yRv/R+V5vC8PHUigk4j1QzVt2nALBANrggjDRz9O
LNR+sCD3uoaEZ9VG9pjEJ6K+vvISCp+1VqV0dFXyC/gC0RUDjYXxDY1wnpwloKug
IFvVl+8JKI2qB1ZP23GDWKQohU8IU2jfPvEr2LJkVTXERcnSt7u52FHFz2faF4hK
vgerDmZ6kbcilnVAUU7L0xEWTHyeHvMhj7X5RZWzkLHCCWzz3mZHkDTnGUf8e6bM
fKYzXRUBmxJn6Z9nUIlVkC9F7ynawU7aLluKxQFbyy0a5vlSPdB17e+Y8jbiINJJ
CYz45Db0muCqnMnMW+KD8vDaG5Motb9Vetz4TmoQwou4uXx4xejqf+ZQWD6vk+TA
ZpOZd65EaHFAecWHhJpesZsQvzG5QpmDeuK/tfcSC2+v+jQnMsGjpLZqe86DQmnq
VJXMcrWqxtcphm7yjdfxvYVoOQjKsAk3zXMidNVRBX2LZ4ziFd+TJGnEq6ehVySh
3Ck8VHMZnBBrC6O09vK/vaa8poWYT6Y9k/qj7wpJHo13LuNVyZHW+hhlRhS89WME
+t/kqK//7Xj7DycMWTTfdKq9Tu+CstHdHWyt+OtZzTx9aLiWThhIzVbD/WVj2pJ6
H04CC1+69OH0ijok+O108GPx+fcJ4dWEy/4zEro36OF3pSyNnY6eLHDIl+OBx0cp
A2TF8WSVQRPpWxTI2vv3zisx4VYIA1ql7NkTQvmtY/71f/BZlJ+b0vBiZp7ZG1uP
vVSd/Tj/Rx+mQy8Yj0L2lYe/ZavTQ52qjXUkoeHy91m6vs/YgshcH4mxGGQIkaGj
WnLN6Yl7fbM+PVyZs4kCjQ2H1ARqR7dkb0YxiY7n1UU0HyecUL/BnUZbFljJmVen
YuM2sJ2B0N61Ht22Td+gsHSBPTR9GNZO7RCS7MUcK2e5VKTUrdl6d2aLa0I9r75C
L/I1EtNkJw8V/DZlTH6LGMaIfzP8tR+dCGHajDh6ueXM73MknC4sDfgJtWOr8yEW
U55141zQA4IGuuigvQ1RKF9jrSMghbCW0l6TTbAP4H4hB7CZQz1JNVXSfYQUuhpz
VmitVruFWsmrJD3l9KFWkns1lynSC/KqkK1I/5NyqNfEkjqRgYHIznzAsJXJQ2jl
7wEE6+kNXzpQ2gNkoEZwjsxjj82iOKiyzdbP3UStJ0wxUb8YzOI8A4C92K5w9pR1
VkS69+HzzNS9RSnRNk6wC/fXKnCJ4RMDXoYPUDMg3TTkyg+3KNwsZP5D0SEt8TdD
4P7Y2B+dfwQBWKy84niSuP2GVeCNlHqrg7iWqAPGbxgM6Dasp5n0kt0w/77uSI2l
Zm6ZYQaFAk6jXzEwxssLmh0y1nAXhw6e+gCUSQ9H6xRetQ05DIDo+9prvGx8W4gr
rYM1qrgo2UcXq0CDnVVAbLyc0PaY3ccA6H9mcP/Y9WfkplHHG5+S9da9pjt5xkUr
7j218wuYToXP1FurSaONCXU/VqN2Hdzdzol/t/at/kdMFVizjzA3RSMseM72kWdB
1KyPhqn/+R1YwKDDzj351MGBMTSxT/k8tVAOk/rKJ/YVBP9cnq7eYIzCPbNir18A
fLKU0q0ziYj1zzqCcK5vlOClSQswjCDIHn2OkqvgWm+0RI6FemanEQmqv6kk1fzW
r1H4gGxESRFDQF4/BzdQ85LsMb8jjEIBPIw69RyIOJZbTA2Yao61JDBWeL8qEN22
0rTUSepjLtQ/DESHxKSGj/lvQfT3KsyfEaMEWcBW2ppUvrqYi7hJ5aYrbbqeaTMm
f6w2Ob1sJHQXdVrB0jrGMtaf1pxZ9WNt4gKVCSyDfCTCG7UTOOwb7HF5a1klAhJR
3rtqGlWF6FXJBFyhMPyhiBPJHFjmkBv50uAfAQL7oGmWKCXm/LRR4NMxu1q+SQvR
0UNxHZ8OpH/cBAY0Bpbnzl/kpbBBLdop4jIANaMgWQtpVsgj9Rg0Z9pKxMjPBY2e
ejJrjM8UqrBNzlRWieL2K2mai65E5nFyixpHV8ndXGHZIIhtiaoR3kCp/sLnxceT
ULGm5148WBShAaHbVsC3OKA7VjIVBuWffk4hr7wI1vjnSRPH7Tci9eeOdSgYuKjg
34YAaBwnyb/xgQtR7YgHgB4u0/zjVvsZmjeHQHAC/8tfHuUo3krOqScJsYPN7dQL
9KZsyDtlLxd3AtazS6RbONSYYuKI8PWJcxIT09ZlJZDB5jhL2bXdYJ+NC+9TANjr
2mz5B5kTqPNhj6AmozQLSDa37uHbb+eUJINW8VO7SEXcPppQ/5WWPoMKxYhINeF3
i3IV0tsAEtuBJ8vPc0iiwlOHMESob4sPNk26LqVuIPMumDqO2T7HeM7pnd6Dv9T8
o6PNX8RMoCMgKE3iVvJRm7yz3ZZZGeY9/Uwa+3pq+pLnDKsYoyp40dBmwM4cdRUw
dtoz/y30zH6D4Bhr/BoVll6haUbgCH19KMA3+y/NB82ubaTb/4gAvoqrXoITlErU
j7uIdDOBBdPquvGWB+m0CDDANOmHQ7PRoB5zrd5g/+bdoY/wKijcMuHq2bVdSZ3D
OobaVQcY67R4XbA352XN2kuu899x9OZoOGwJ6WLE5yfLLAQZOa+qBmjRbOjDpGpW
rlvnNvc1CZtJKY38udZsuf+zicY/I47eSf3PomB1FQUQ3EwCUZ5wzAkuOnT0STax
RrKtfiyCOY9BFm0AfOuayVlX4YpzNm4Pg+z+EEILbfVEifd9bJP56Uzx3L9FK/Nh
nlPVKrKNQHuV+UplgCeubrCTUxybqOU/EaYOJTKTAF8pS8PmeGYpAP0CMm68PK6M
tioRMVOXzc3VxxIEDEh2cshkm3c/uEI1G3kKeqSCQyI1BRHKIvHSrjLySHDjP9ww
tennfu9lwGN1JyIuhfXJvurARZqKyUSVas9eu9lCynNKu7Rwpqu14Uw/9aQP2hx0
HdiYS2vHdTNRLQnj0YABoPFl5aIO4t2GlmjOfRXIoXRj413WsaeLgKBwEt0h5lXK
vHDuwVlPm0mdKRD7sVh/LT2kIsNRNq+qARbwfALdRcOTrJEUxZKaU489SEhD3d2l
JBz7ADlEQfy53uzj6qrkri2fgJkfYJ3gB2DIos5fjnBJtOO+jMwPKXqMySd9YNja
cQuAFP3QVvdxEp6KrCgiMZsGAoCfYbpwfIzpwxeNHYlHAIESjcIPHxljlMIIECfH
Ae/yrWtIBQYqInLCi/EtWvcNZaRCDbp3aH0JdXGlYQFw+sdr6PVglZO0YLaf+F1t
YBgO/jy2MhHfyRx91SYqgmtgxBVr475Rz/BMNrsl+4c0T11ZT2UwUHcZRGlvr97F
RgA7LX177p0N4fySq5P+LBGV+jRyG4JBHOVJXMZLPl7LvjLGYV0phyQo8p5fP+u0
xx9piwAvldkR85E75CxvuKrER52ehKJdu+0QJ20BPRCADJsSi6f5dt39Le8reWUZ
gg6pU2zmj3o8lvF31M1haDhKtRt6rX+2Z4z7rwgXRczzX1h7brnbdnr6SzXCYE6C
w83WJB++00hs12BzYOMUL567aSgjqCgAJQnwFph/e+c0q6sY+Xi2HBFOeOhP137l
j1XuRWb7prsr5SCRssSr/8SzFOU6pgb4EFYcOUprn/UIIceaHn9XE6X2nHwAJPN1
Y/muXCaTpRP7P2P93V8139llFWvq7wB2WkRsc83IcOIXuYVuqK/zQ52FdEQ3bvXl
yBVCP9Qwa2w1PfuYGcSjgF1cvPzqzWIm+o3jFGUhyuUK9CeL4Qp/96C62VgRQoYA
5iKPh926f5R3Ou55W2slp1Ch/hBmckobc40k/LUoNq44OVL0qyBO8hXPwxEQwx6d
SzbBq2Uh5l1VDSottkU6Wnel2/v0tr2VzzKD1cgE/WqdnMgOIHAiXitHRfb9m3dx
Amkh4R4d4c2FgDG20TqN+4IuwsC4VVUz4uGEaPTaICuj3moaA/UbUoR25MJcyxkI
oXg31T+PdG+lES8bnGueMmdpb0EzL/sAbqLDb1ZxchgGzC8rkB0US5zk3109aSjG
it8Wr6Ktg0Y0gZ2qGorxMrPXYPxBIPMlh4P2WEZ6bOshw4BvkO72XjdIOkPoNLxD
RCprr6azs3Yq9bYWLwol75DftkvRuXpd/I3ixHU9O1wtrMbErHre/w0CAoB6QBKM
/z3sNVWyApy7SqC8wemuxWZhGPIxSphfrHB1MyPoj9WGLDRVCErkGxiULc44oY3s
6NGNnTi7UUpj7lDlEM3fJqc/Qv9YjAYlrc44k8RGIw66+6ez57ePD2viXjGonf5b
LsTeR5ZlUmiwvJltCDU9lH756d+Y1JU3cOgnuRp9wCA3VXxcWpGW+jRaOmPpSmhv
zsZ8ewUdKpHOeqPphCQLdCCSKs+teBzrL9ATJ9r0cEttOg+ikA3Q5LJOk+NpQ5MS
vjgPMLKLtKyQjZshRwvWrcBLdLjLrOmx7ibE5o5z8LXqhtIvjQp5l/pqwyJKD9AG
tPzwumZQKiSp6H5x9JxHHLdAzhhCV0hGpKVQak5avTthAcPQpNlYq8kdmk5oyjvV
Pl6RXJGO1Wp4Jy7GS4bX0pPDpNo+06ktjaFW2ulCQNQcUUWjRhMlyrQL2E9kaiIS
ouZ4mFM55J3jXObi8vmd04QqhuSpoOYojNCShifNBYruYp3yzOPIeHJVZ5ajNlI/
t7lHTNvBMHzBCYkBnFZCDoarwYV/e1etG2A9lIvIT2R2xHI2O/2QRkfDS3SbEFIp
b5h9/R+AF2oikgzHknX5PW3X+jHlZHh5mqcZ2YkpsgN3tUPJSzJ7RAoJFBHR9yq4
CLMWlXuNAwpjOqy2afMFqVIF5GaL5YciWeJ1mTGEGhr5wj1dweEqFBanCCSuWR7G
0kUiLtE/ODYN0eQVc91b61XsIp9G2ykp8jmdawGSII0QodFkymicjwwo33JxNeku
zVeuKqCou7ecK04gH2qUAaNRQgwxKmpFKMwamDWGrChLxqULdOWI0jTKgKG3+yET
yCqFkrLYJDUVV9d7SfLz/Vrl2OgJbb6VH7R0DCnveZ4EysSApxAuYvErAWgau4Xk
T0NxIi5oolOAvClSWIE8Kgr/MKFVUAa7s9LIa6FZgcYip52Ja8hmRhXrEiYjSkUa
/OcQ2oZRKgMncwfWzsCgpPTX7n9MM1wN/0PNX2OVAcNmdyvZpQM0OhF1gZMfAllW
W1x9we+uUAoX1ZegWDF20pYLwH5jY3M6P+bHh9Q2NRvSyDiYkySH0vimYsrZgtbw
ibog6XTbLzLGVzoiQDBsWOT3J061KZ0yqN9loctDUnf425H0a3qD1XhjPG9fzgYN
MT06pH0zYtR9f7pMSoLmqVCUkZAEvz/VSUQW6s2vK6Krt7BgVHj8x6D9sapfNwRt
f6s808joSjLbWm8bAHgBzZVN8u+/hM2F1lrqYiS1e7ok8r8gvitolRQk9WspyILb
4aE0d9Q0ObZTg0Ti69zefqPwISf8pVbKgeRHKDncyFun/4CCu2CjgW6JBVjhQWJD
Eihv9Ymm9Yxc37rLsQ1g7Ny+H9VoaDppw/hGw8HjXE+D0YlFWIwmX3+7cs7dsMg0
P2GxhF3Je9jg0nsL/Zkqvi4GoXAwf7As6bI9rfvgwtoD9Cta20D+e4Cg9JcCW83H
tYFCvNhETAg2+NXE0e3wh7e1FAUd1DzkJj7xyTZiznUwSDNt3ixFkoCiwnmYoIYY
VilkD9jbbTiRwyBJN1bFlVmN7q30y8ATV6UEVbfQmSbWbBLUc0el24cai4b+qWMd
wCl6GInc2UgwuFr8AjBWx/1gnaS0hZ31oR3BbiR3Pdnv4aKEHV6NgemkPEdOuq/T
zBxl/jfo8+IU7IBctaj3y1RLam1Nlky4aBFihy997gJFJbio876ZHFuf6QN3mrPG
0VN75TcbSN3R2LMQc5Wvn8OW7A+cFWsaCtZSf7VZJ4pbg0GKFyiN+1T2+ZU9qiB+
RtaElXxit9X/6IVdrS03NU3Hj5FK5Uo2//h55L/E1UVS3Og6ncB6Jdpa2JoJWx9X
T7d1yK+cR58h36Qg7rXBHacxdnjvDmAgeOYMwWrO3kEDo/zQI40n31DhrwPG2c7C
fTe7rIx1OD4Zgee9y1HgAs8C+nQ9ci7RexRA9km+er7v7L1mDkyczjhO8/+A//3I
IJ1alU9wYlEyP8XFGCOVgCeEkcIp6KuBmvGf76tvhGHcKmvEXY8E2RcGKPTkawuk
4G1Lu4OjbWOgrDf3aWAb6Z6ra67LK8lWFBHDIzfaspfAbvYViGcbtOxhRXlFHOOt
pkIQ2I5a0fFSSQlVDgzjU+gRql4E0hlZWgRXP+bDQ20rNUEkOwr937gR6zoLzt0c
VmJBWCdagaMsf3wEMrKm45ObMDHQr/R/mp+WFBynir/uZWBfUbnk8ZgWhvyZes8E
Z/xzLne9a48PMsjmYMnfw5zLPmaiFX1B0h/YCU02euncVBBZLFAJsVQoqeV5aE1F
2xRT5KcMj4cPBDJGEXPubo3ey6r7VMCKQ1Qcapcdlfrc3sEr8MiYdwhc763pzE6T
+l9eNPJlVMvChlkNwxhBF5Rr1btkEXSc1pWuM56gWHocDR2VyBUUJEnuXaYvIFde
AXbvWn3HBB0j0nECG00rVipve3MyYVfFmbU0jUq1LK8abfwasQe6TE5lSjSxlEJ9
6ijn4zBq2MXvSOxNKlfEIduP8rwfW7rWsS0oGfgNf9MHGnDSPzm4PKmWNAPLH8v5
m3mK/wXlvwo5ZhkBckkRUrieLRG5BzmTjjMCARVueVxM7gFT7l4RHwogixGpl9Zw
TcPEdYt7gEhR+6hRcwr4mpw7eimBO44FLqOHqUIvhqy9fKpty5ExM9Wb+xudaypz
4Dzr3gq81tzmiXw3IloBy7cORkT5zKPCFkruPY3UQ+gmhYvvZSgv1Xlkgvj0lWz9
9/5yVC42f8JfRXxpQlbYZZRnEEAldEP5HNcOYuWTCbdCNCzCG9uT+dipRJs3ZP/y
Tf3INhbLAIfzADfgWx0e1IBD81stfvWyTYb0CWrShW7+ANkM6dRNV1u3WoI6y0EQ
zNzlMLLIRXJJ725JZ0ZFh2VhD0HOdUKw2oLSFJeBORKmuOCtTEA7kF1hmhSj3COw
Der/8M9oeRg1oMVSTrBGQu1NLIajA2l28Lu/iMl1q/TomOmuDHVeEm1BeUUAYDix
qC50LPJvBClvr1GPxDBMDOwDX+sz/MJeeipff+dG7hrzTX3fIEMxGoe4zsKPK2tF
MOyE6qMBG5o2Ex2c+fy8mMBUaUDH9IWj2QR8H/n8wEV5wKxzLQO1K0YVw8CKsiR/
FKQeeAwKvIylfnOMLwkIt5hx5D3wDehvNsAoRArTVisxtECn/9ETytGDgd/AEzQf
DSt/vq/gd+LvPOmM3KvCq4w+Kjm03Ssn5QJraqSsZ9qhhy+zg0HPiD+M3HbaByxA
PIYB3iUKUhIJE0bYGMrkxw8gASBQaLMjk6HSDVuHeZYBtlXbk2nNvNUeiH1CBrpg
PMTeJlFNWxCeqBn3GFtsveyvYn2pO5+zLj34Duxdvmzr8zQv3QNTeRLIXnAVZ/Kl
aOKa/JrE7fq9ZZIDeaPMO74KbdyGa0mGSNFFpAOA47ByJkU1gTtRyJkASJAaD1FK
zJoRzDosYeCzJZvbAWZIBup2NzaFX8p9S1ADwHRJDHFDzcZ6K6N9RElf9Geb8eRE
lx+u302tNqUKkmZ2ktKYk6bEw5/HvSseiWbEuDMxkVkcVD8U4tMYW82ActgGcfOR
dq03zLzZm3+HSd21cKmY9Fab3+jaoovEaud3QHqXiI+mkIZ4LneOKD4Jmx/1pHmG
sx6qvpmbTzBzuYwucDstprusy8f5WlWGn1mc/qH1VIjfUXBLmr3+QQlu7Vkf0VN1
wCEwxMi+ktIXVVYzzyvW/K4RsW4D4DCQc9XvuvieK7o7RUM878N/8RiOGlOTaScC
n5tz2ValrosHnjFhXZ0vy13wjktgg+OCAAH/fver6feXco5N42flN2hCmlvU0fH8
uismxn0Gbf/k1tJVExcR93l/exhB1jMGGApN+KBVy7C8/XEohcEGsj30Vvf1fr7c
D5mvwCij9m/RcFQORjYuPIScHPrseEL5PNkwDMRudXkQPoZnA1EjnNBUN6UASeCU
/Wk85TpR3IensYWbfxcnjnkAC7NwiwmsBO+ZpahLU+8pg3GHSyRGG+nKMo0jw2lL
C08HZfBjycIjXcHXYIe1HzKx+vRnaA4JmPOHeQy6xeu1V1lHB/4Zow0xbCn3aR2r
YE6lzBSEZMHYW/eqxBG2BEZE4x53IdAlD0fX4LhZ4V6vIQeZB3QjA1q0r0y/FuWe
RMuB1Lpiq6OeUWJYKh3nfZx6jTD0VIcv+moEwxFFEpXJqJSNS/OXpPwSazqBaA3O
ZqcaKInijks4I4XMYNIfX5xRK3gnQUGvJ72Rrzrd7d+c2iUmFbLuuiPWCUHHyX6Z
13zYJj1yKSnzXlxRtAAikdWaKa3BjslDNNuXaoU72buYPMe+VfFh54skg4iZwE1N
xhGBEWmrJHVzPVBWhpY2tRCBT10sSkz08VpXgbp6+ebubQvT9x0pOniG8kUfbppE
EdXIt9Bqm1wnrd0uy9s9eG1F646tbJDfue9v/YOI0m1LypCso5Ody1jRGdwdpqBT
wEOr4TIqX3sx0xqcOAgBK4gMxSVcXybZ3jcxMxktjeHgb2uLZA3P/Mn7d8kBVX8v
wiyadpQoML+capWHFwWetGNh2pXyeRZ/orUt4rpnCHsAIe7zyhnOQAd7Qh/cJpUn
R1B5iGNElCAn/RgsVHQ3utZz2zfDfzIVvtmvaKYCVAukFUbSzv8ok2t1hXfSosza
7KV0hDizZtONpYBa59rjZqAbSQYJjSq5Lh5eRwOSVe/fhI27LhCy8enxUmO4bpjR
xBoDAqBZQwK6OJxQWlJr9EL4NylVMHMrBP/lxQio1oFgjpLcUnusU5Y8yFwfwCS1
LgvHvJCY2grT1LmUmq9ur5WmX4kqPmkz4oXgvX0rtJAxawz9YyO0B8gI8EdWD3Yd
pSWTg3fypSyJeoG8inFenKyuuxLG8ZmPVBmbutTQOHeHJt1qCdht/ATLTKSI2fP3
Lhh3Vt7ch7JY9O9qP/t81pH/AqPPBcLZemfJ7IgJlMS/DRpPHtJKWu2JXh0dleOS
4YY8PjAWJ9vMrnjvWTuyXNEHvDm6YwDJXANsledZsOiRs603vBRQFwK05jQhP0jH
1vl7Mdy7Z/I3HHRtrfzs0/Yi1zXeDiof1wgBlCVkQeudvU0XODxGviBPoeneHr9E
20ZAgPOgeYRXBm0A+Ot1ybdNJBnvrWoEtIR7mTXfx2iCdTlEzGIXXVz+gJg0dxVT
SEquvW0aLu9NoDVg/xy2aK5Iban1zNw6steebdO5EuKNXE3Uwf1I/wPPdDL6sEJ7
zx9PHBDiGKXCS9Yx7Hgz1p4PZsCZ3bOaVdEFUr/+SKC7lU+CIKudf6RFnE71VWBx
dfyhyMFRJHPZG77OdWSDVzW5uVLucf37INu7WQfvFiy4EaDXzOtV5lgFO2ojKv0V
wPQdPOpJJCkYL+TJYjAUJRnJb6eViFBNwMWVJ0ti99xLpzyDYb5r82RdRNd8At9h
LcpCbQkj+eqMkVu3jw1tK1iscnkXeck29Mky2ASD41VeiYIQ6WU/atSLKBnnOlaw
hIoRzIzBqgTWXTO1pSIqSb3/utnMZ5WCxpnMbJU64+nPTzeT4SCoeop+5487tgv8
bHVV1qKEvPMk0IvKaIU+xzhyKVJlo6jMMLSECu/s9YOdnuGpE4LRSWOq10zgk7ii
87LFP0zBtL/7yP8V4O/Fe4wmbVaLCZAqB+jupcdCsz8kT8/LLxO5A8pD0VKnNk+1
ruIYXM5EyVmY5b9OvEWFpmPA1LU3begVrcIIC6gb+VagYkAf0oZw9UtkjxjsWWDf
yYH8qi6aZfGzCXBc8Z4Qzc2tAlJx314sOWfOvKtwCS83boo74NlCk5ajB25o7aBC
x7f+zemxTVkk5iQLJzJX7pKlAI/SI/5B29l8Yh0wErQCssVvaNLf16PYxOstKQcd
BoKWQdexhzyWliLCeHKibu/191vL4AXFJtLf6kwOxFt2AiKiMjiJMpSfBbrNYiWa
vblvgDAE/dOrRYaQarFgPxq3OyQAQefZpyDisy0HndVepDC+T1unU/y/PNikam2b
QIPfYzaAE1QUls08j4X1a2R+Kw9VqKIpT8RdVIKMKhAhbLM6CHo4lJI5Fpm5pLxO
HNaYjYGfhWBMqySfH8t6nP9Pa7a4LrnQzwV8rKsapV6BqE54qVF9g3mZfhFIY/c+
QQK2t6bbtz2MaH0+JZKLqcl6H4WK9epyqRz3+LovGxH9tg4qxSGNNPve3OVJTYny
WKgpv7MOx2PDH2+AiIC9fBoniug4zWmj0k9grsF7CCUV6CsdPlVsxdaTaDvEtkoR
QR/RH4POCBETW44EPupTJATHnqUsz+AGnTGR+8Gbg3rI5ho4/IR+2BuvZ3oanNth
kyHRS4KH4+OEoEMtVRsbhFcECvRpfC4NANmYCArW7u4E/bkzg8G/3L6WK4h9mYol
QoaAlCZk2q/be5bfWUuKA987+eKI+7kSr1GgiUpzsBBSh/l4rDG/rfIMm4Vc/vma
Es/SQcEC6rv5BOjbgTIsSnLDkR0aGz6KyygQi5DMvrRU/A2FCD6dbK30LvD1f7y9
4+7nwSy8KIApveECxpl0LJbiEqtSvzok991KUlf3SItPJ9nn5lMwYe5IJQvhStGM
tGEAtYo52xHeBWa9Zz0yNCruZQob/ghdAkiWf8SRCJEZQLAOojBecx6OZOw8Z/M/
06Ia0RCGlYenJlZ5453eOzAl54hPLr+zmJjbnpciT28T4zZxua3H2FR4lDFWRY6X
QKqR7oFANqQG0fCwR2/r3Ijjt4Fg0izdfm2gn3CLq8Ct92lNJ9KuoJwlm9/m9djl
b9dP6wgRqQYHQ9zIXI11An78OY3QhFTY4DOUYXQ3V1FT9WannhGUpDw876hNAxsp
mGZLJHvx4nEZt59uw7wxdtzfeOmDzWUxpDPRxadXC2ZVnXgnQnhov2prJazHlS0s
BK8ONV55hZEiCv6rZSfGMc8N4vKrKPme2on+iYKLs2ZtgATSr2se/sYNj1MO1jBk
K2QViXoASSqof5DTYIgFghM3vKIURqgUUDsv0HY9jDW2kNlCWcdF7tVAVpe52ypO
Rjev+c67j4PdPO9wfNXg0GrnZa0Gya9j6L3ll3hn3+hZpYcBVuXeyItAR0vxbnbr
2p+Hw/xz0yBW8E+UHLbwuti+qRTWuElBV/X3USDXLzijYOWalnGH3pVb6x64BaF4
3hkb39AWj8GXoTIXJ97LgtYkcTv7r1tXiUs7Npg++0n8HvvtV4Dhu2wM45Tot3KT
IWUaMLPWSWrXLiQ7SpMTKesxTFjdkum81hQVgHLmUjyl3yRyMOyoa1xA0qFTzkHJ
hKgUSQw7xBJE/t9ZoG0AIa7RcJYZ34rwQdVUivIak3Iv9V1BRo7Vyj/0Q6p0/2Ba
4aSMpM/Ju1g4XoEkztgNPARrpS5sNhzNsf5mWJYBVJl46bdD/t86be7Q83wB1cPA
f82TCCJ1nbb4OstwDFu5Wbuhg3MNRhavSSmPefmSVlMJ/lRUvCBnKJ5XEWg/1jWx
Bqj34d06TihHr25b/cEEgyX1SGmBDlEPCFE1Jxd+CMuR4p0Dv2CDb6VN5Fy3R4Jy
Z0mYLZUpOqjE/hPhvfIwgUkLB6PvIdok9eYqKnNIcPus5jUu6x5s8CCRwI0JCaay
wlapajzO3PKnO5XRxe1uvPHj5Cl9g8o3fGcuvTkoL4BUl1MPljl3l2KIgAp0jDZD
BEVR045eyfe7fqeIL+I6IHm9PO5Bdei2dzDDaDkoUVoU4L88kcM38TsSuUao8kfw
6MUnKzlzySzix5KlzbLD2IUJ6cAw9sJFjvlvEjwQTEXjXcYaMfECs0kLoEhPs3be
AGd5S4MPluXwRI4hDv7h6XsEvhWj7WqNot38gtZ2B/U+VxaxCz1gyQLBQLSlOloE
Zd0MSpCN0qDcQMjFTj7aAVzQEUQr69k+efIxrpauVubjzp2E+ElMOFj3+ugjAZ6a
yGed6yEQMZGIWq5BZeQX17eAVrMOYxPyGdh7OBgQUOEGuQZiOTk2HQa7KJnVGAME
r8Bets9G0RjNmUob/vf9c1kQC7YkgNrni6zLTYmiowp9oUi5P8jjsyAaPwJ7n0qF
9uncLTwy9YNhvMsCG/otJ2FWv5+8LhtJnoU+v2aam0rhwjIJLyzq+j0kgYRyW5+X
bto1ZOBNQ8nb0gsXJ3xPJWHVQs/9u3dzbL5yNbBTUEMYEMC+fsZu6nG+v7abRL9+
5jrXK2QqbvfjKGKPWr7vkWb0qX3Ga6J1SRY3usN77ARU4eR/XEjtm2QpZpNacVfe
yZaMOWL6ye5aHsmVBY9PDYRW6i5ccYHruA3v2JRZD+QnA6ZerVIzvc/PPtbzbgyL
16V4M0I+4/aAez8LOzlQAHab9yf6JJcrhC9KqtosQXqeZwFkIF/6rexUwRgoP7CL
vamK9yhfiFQZ7nlB2OQMFGftt0bJI1ZijaGTDMzGpojr4NgqlBiunKT9WGNSl0lt
z7JcdzYx+nqsgPnNr6xwggokeyOykSMRPanYbtZTRDxIzTFStSekpr/2+3bXKqEu
og/2r4MHHLv0kBQ5LuDe25A4CvaLWA9Ar6lonuRoh1SqH81PA1J/cAjyAsc4EBzL
quTeEV9GjU8xtwCQPWlipbyoln1fTfVN479KH4mLVkg3v1TqWV0VmNyWshEpdIHS
qHRFnEZMqYfFesYsfCS0Z47Qmr/dT975MKX01p4/Lv/1nya0NU+H+X9FaB2cNnQ/
oVgfFVYp8e8seF8Wnki5zhI0nKmgNibBPwmLB4g+iQJY+vRTv5tXWAgU+N0DmxBY
se28/wlBZvp5cQWa42aSyw//NeOLznlP7VOXsAEkBgs9AZUhTTI5O8H3E3pleeu/
RWnXCkCM3Z+VSL4CYGxgATy9qGWq9Tmc8eiHgF/H1enZhMtvBIDYxi/botDaeq5V
a16FXrlhAwqzYFk3YSbZTBoQ4O8VYfs9bL9MbVp8JZ2aZCo7QztTPtiFNwJI1VRU
UjQgdZi2Cubs42KQT6u/FhYyYeoGbvbgPkFOU216+s45Xh31A/ysSy+NBKgQ+dlW
rQ/veHpInvJaCDy2Nq0mtbLEkqQyQ0Poz/5S30WERSIrMu4T2eImnZTtx9v5b20s
JL5WBgnW1aFWF0LSVlh5k7Wxu1gL+QFHA/dblkyYry73XCZSd0VolVCU6hDieAfk
H9h7MrHu6EY36DeDoj0vvEvpWXgoyBoojVywii4lCnZWmAsUiaqCcVZPG7Gq5G8/
od/bnd715K0HAjuKexXghK+5IZWC1rM91P9ZeSk9gI+iHMJN9eBAZ1P6nbGV2U81
heo4BD4Nw+Kl6HVPzvyvqqBF8pjjbR/xKCgUGsQTBLHQwYcDmtmizw1X2D1qSUhp
GZ0pqYnWT/brEn1F4wZkrPFEH8BWGmUuKkNfHt/DoC1dfzxDSDBhh+gfDh+hrVNK
F09lKq58UgJVvNcBF+5gXOj3BrX2tMPn0DJtx9MFOHpGz05zEeOCPS8HHAmsyZ5O
7FJW9e+W4usKFFKlFar+B7YlupQHrI0iGttO0KNvsnPL7rnbBDvXD9QiLA1amTUf
2eGWHbjXZe718atMNBZXZfR52VMJaKYAfz3bX8Hj5P202SyFyo455kU5nlnb7oxd
MmWSeWc4uCTe03FgIciOyZ8AZiiEmyzlB9iwkYybCekcXv82S1llCx0jMp/piuby
SJxrm4o1nrHTp7OVicbdXj/4cuMAXipZmBqYaeq1Bt5OvoAk/T2dchQabkNmKl28
lN5Ln5uH7z8z6FCtV3RRWdKoNLqsF98kKQiwaMTIPvh0eSsKRhF+c99P+vGTeHPB
tpoSHq7m/S/QesLYfsFl+Jd6W3Nj0X4PJdTwC06isEJEx+4PG+wYWHCMo9S2+wFm
vgB8Nk04JGG8KoIGpXXv+zjPNHyB6DjV0Wvze9KIup527xMvOAI9sDYIhuO0BFqP
ydLT6e36bJtMqsucuUL9pxTyJLO2s2PQs6n+u5GE0gjNrP3gWOuoP5ndaJbf3HK5
9NKUDDufUG8HNxyneo6vLd/vsiNEh9yzrCX646r1Emt/q3Q2p2q352zI1BIBnp/4
/axqWXrPz5PZnZ0/9AL+dZbPRItjbvTxuKNMzwnv2lU+4+VxKaa2ttf5svGg4YAW
sxTg4qXOi9sZjdn0MGMwbuD9b58s1hMWvFrbVSQvPmyhUVLJbTSPmIaFjp3JW+un
1S3KjxYPZXSLPWB4mjjVWooFdEtIsc9K2zO97t0fXMLVClol9vK42nPaz5TFZ04r
98t0WIF3U9dFfd3Fnt6DR/uh+WMRLG8knKdOR3c41NNAwMp0HhyApP5MCUdYOEKh
yDtJX/d+SThKtHS9d2eoZ79bsJ2WaLe95wg5Lfd93Uld+QqQnR5LgESjfbgLDNLT
etVBcSLUDJwN9PUIDQdA5glaxTYFbGYGSQwSo+3Cphouh9Yyu6PpmXT8PzYPZSra
qBVx1DkF6XShhYDuwQx0OmNsdFlw116iz8O8Kkvnjkg3a/7kNsGSxMDkBK2X0dhw
elcNjgbYV3r52xDxydbgoGEN0NELmy6HsOzffYEob9Q15ZokmJLwuiw8v/Qs2oSV
0ErDTIAlDiSBSwsl+uv1lpLQeI/B6tAf1fmr6+BYPp+Z/2GaFO3ytJv3952vyhsl
2ceRjRJoBa+kNqKcBx1U5rgbsU8Td38ChMqPbcIWwufHsKU/R4PQiKKMWcxIT93X
OqDTzhrYniDWutwLfGdU40/4sXBAL3tPWC8Uon9UIaTDoA1rehE7FrEYf0+lYTs1
VpUBfKj1NjmMJ2Bo8BoGB8yyVy79KNyo76bwplhz59gQ6q724Ujpr2kurlCG1sq2
TaaloKlCQyoSNxGM7r4xsdOg0vMUPUR5l47GAyH8XQRAF9qPCRlRo/YJF8ppCrEy
MQfBo82ft1Qk9zWYuYZ/klrsdRySqcPGhtAVopRE4HUzBgunB5ApnAhV1fXQFvpu
p1m1sRrnX05zjXzk7m1RQ46Z6tZSmndAOtCfR8EAr766n5WWsEZfjUrBdIXn34lm
RxaatpSfQg0cgJnmUwajsOWWg2dZEhNGkc+Vo/Y89fT1xlQt+PW536OYXQCm0Mt2
wikZB5a19Q3yDOkdeqkbP2LL5G3y46i9IpgriTEQ9iJqvA0Xp1TD+Pi/VKXpU5pn
SUm2B5ZM/OsqfC8Mk9XCfouB/p9RzL8c9P8rlm9JwrNTZQswHy0GgGLCgwmbQmhc
JFzVjbs44GhMRuVrPgryYMw9GGguBeG9IeIwvq8bMg9oAHAfgHAoRY+BhF9CceuZ
cpTCPixewnVsUJMIwNfwyf5IpZvwh/cIzT1XIQNwUb4+7Wn2gbBTLgdd2OCQWHK4
QnTiW5uSMEHOkne+HR/fVGRH1Klu5uhUQFYdgRZGiFFtQiYzMKZPdYk+fdkWH0aI
2vSZrI5OdJjPPSmc7I5L/aBZuHn4FoDE82+c8EtanzIVms8a7hqfuk79ZuqZi3Fe
155aR0soAj1jKCTOQA0a+SaepjyQvuhxxYIXdaA71I6v7Lftz6mdhEBwi0Z2cerR
gbcwb4tF25kWUQ2z+J3jbIbdhtdHqj8cBLhkJjHkNsSSlMLS04YowU7KuTIQFKTD
dFbIjhVj++YTVxk5+Dixdy4hDSUtZRPzmu25zUVADsZF05Hn+HgrNB5w1vskWbXD
65VvkZGCryYvlT4W+KE564gfOWnJAURuNsMv74uLTnztRofKWT4SFXZ11kB0Nn7J
pVdmGa4kSgvXn5+UJI7enIS7bPsd6BDjcaPVkxRj2pC86m+44pZgiUw5l1QnN6ci
FJZxkLJPVlJQJzMS33OLfioU7Ox1rg1ucQy2O9Gf449zw3R9chKwXH9afovH+4E7
RZ80B2rsBQSYmsICIlp3WOOptlGDLIw/jmaVv7eOUMUae+YAvDaVjbEzDt4YVkBY
I+XIYzkbG5MJER6A2dv+qEHVbY3X3Ss2cF7itAOABXwQRwt0RRCZG7TL0oORx234
aKMqQ1e9QFnnBXOz5crSutZO7Sr4d7ObJEmSwzInmadRvmsGONpmh9DwvNaPAr2f
R+EyUMmvUsQ+yjT/XHmH2zTK7eExBAlLSnD2LPtHnft24cjrS981lya/HLt1HDhY
7wv3Qcwd1xDvtZ6t4QfDc2D9D4IQyuKFS8Dc+1goU/aE6TXdNN+qzL+r510g8x6E
EaycxiIkoLiPA5P/EFAmZwav/eQnHLg7l1luBWZrcJNABsxgj8BKi8xjEtWWCEN6
7VtnEnjKeraOZmCBFEsMJFKbne23nAMvHEMdPbxVo326q+O5AN9T7TQ8n2qJJeqz
n8y9HhAXP/Q6utCHXVmssGNPwSG37dybqPzvxJ/x2Y7OYB3WmjHgIClv1XvbnSBt
10yLQNdL1gvHxv/IayrOwjytf3szm9S5tWkiOU8bAM5LgEFqzeSeL3JVlCw7ad3k
vUWLuna+HmHDg237/sYn2ShwBhucRl+2fOKrOr8SHfo/3QIx3avAYdVRBR92Hcsq
bG3PcDL8f+WBdE8qiq4XVoN5GYoZM58SWS4oHBHHlSjX+YW2otUnB227mqtry2kq
duSXHSH6Ri061W4CmxOqjEVgvIKj0g5ByIcli/T5+coVZVeixLowJ+z6Zg2z4yYU
j/SVQNykh5YOVycUlpRvScNfw6bNFH3sREHg0IclVwwVNd6b6yb8CMdonh0pMjd+
vaiFTpg9J2nTWBusMBFeDrn9VOE4ZRJR8ssN8hLvPKTOWkGqnHYvPi2XNxWDdjE6
dJRk1y7ykJ+7DrgXySJMNXXhaZckKiXisJfEA1pXBaK0/ZbgTIbqQz0XcfeLb0ik
/Z7DO4d4WvCzC28oQZ1nUnInIJn7GcBoFBPGg7yhhK1K3eVobi+ZMpLBbwtd112G
mzQkSPmlV9FuNw6f9pgR3p4nyuYbtDNKVLNuQTqAs3WUgDtCeeisS3O+XopW38I+
8Ne4AL9+yk+bxU/ZXyOrHIVDkz24Pqh3svmPV0G4QZ1HXB/FwWkWQvhs1mbk0eTy
reMEAf9qKcHivxFufY9jz4LV82+GCjqVGOAE8dLuLu3Shg9h6DauolWUxwTCwuOK
5iE7XU+ra7UHmu6DrSZznVAhMFA5/t3D75lqeFZbNa+Ncgf8RWqk8ziqNqFy8v1D
PWB/g2N9+hppcpFtUBcKbTm99KznDbR5v74XR6rn73Oy8MKDCbXEFX1wIjcDtz51
62qT948TsobZ9KIDc6mV3tOVAiezoo8F2if8OJMJJQnEtcR0xvxa3UY1sgdrkLmq
oKA7S0nsmMdGzTU9ejg9vDhmQXghLkO35V2Vf1ueTHsrrRXBURLL1PeMHshjQpwn
xnz2W7gqN7AfiD5ak7gvRFSo2BuL5JplycuvC40TGc1BSCZLhOAcUQ5EwSdBDSBZ
Q5hteeCiqmanE+iekG4UTYG9T5em6z/xYVP/BBtuFN17I/Mh5HEVQQjt4xMn/4AT
/vpqpxO7dKW6+qePJ+2n81IFzcClA5hSfcbjKVMBDLrRzwWM/b6zvKceCXw3Gdkp
BYIxOhdtV1dxI7WDt7FxWasQB/ZcEX5V0r0bU3xN7StLqxdL7erGnO6rPkgfTYK3
cW6pg/mkfesY9uyO3uuiG/apx+DMPUqaPq4/kCY+bV4wbopKfrK/ZPOOT/uDUeoK
KhdKjBMzpoaLZ9KhFyk2Y4u5nvVJ6prg7cz8Gb5q6/YpB8Uk1Y6ICtVHtt+bOjDU
pOg+N+61v15YBBonHr9eZAA7kcbJ2N0FhUE5pgaUWpPVXBEw7nqdP+KkqJGd5awn
3C2uabOJv9KQ0MD+eq7nrgfoE0EvFtsIUsXYwOuZ/NEj2f94pEW2LevzKS13qkWe
aPZMzye8XLZVEiX+HevdniGcNYu0pmu/03NgOGLz37ZtJh9rNbwsR8HguWtOGx8t
RN5yU+1aODGRSdMKtk3GN979RRuyrCECniY1nydJLLqjdRt2kgdch89bvl1TQYXy
v2JmyJhoRB/4wxkUaUqE51KjjuNOb9xNOZtZqqcmIYSev7BAWGi5AypiO0hXGlLb
ByuR++TsclTA5vbQGerVjgmO/8OaS5Bxp+rP/s9LsFfDiMKaKtGs74yB2XGWgXhP
rxb1zDbgfHU33L1xfcwyJyq9CaL9H4/6JfLkp7hIwK+y3d7d1eZPUS9s5beGXlZj
O3BNDtF/iZuAgvH5Xlx0pTC9v/G5mS0kRpMRk1/4ZilpNBgxQVD2TohKF7RWb7JB
XvU2IYY61dxTQBhwLu2ztg2eQteqVFJPYhSI6X1oGldnHJdlYQKCYBgAbHQ2I0c1
JrowxMoFqTEpCLtNCnEl414PhnBJ8YFIC29C9ZaALn47wH91uPJpaLuP/ZsjWv/o
KKZeXngstISqQNxVnTYDihe2hbo079wt2ls8qFmp2myCtrtnmTKYND/r1/5Owk0B
XwBaL9ka1SuKaNJamELOZQaj2OGd61go95NjnLn+dQHKK/2aDdxlt0K8Rzs10tLx
30UO75nAQcuMFTorTj4g8pHVhC2W8eR+qB9yj4edwC8+czW1AqILcWe7FSRcghLu
Ny4CqC1SG+HwrlIYSy0JF1+0dbS3W/+dke8Xbc+8gSnzLst2H5bgc4gnVMgkA0jH
DDC0jKpQZ7ieEAmz7X/qUPU8wEN/Ryt7dPxw/XTb1WJhiCXnwViEDxcFUmcpCR/N
dc+0MPK5TwNUGN2st15thF6M9qCGdXgXjnz19zXoJJnEDcmimZnAc/nEtYiGvubq
ptRnp1YneuHmIeZrdVYZwRyIj/lpztYDn7D1Vmqqf47YHPZyNLt8PGX+qdqVev+x
UiAshAjtMLgTX1naDxKv5Cs2p8OG66sCQ8pQCjAStSGtDQc+Vzj6mbxnDQ3z7PO4
a3xL0LIxz0uqgTwn4SCYdZ0gqM8UlWlVIIwfXNNIpA9knBU0bCmAwoJjBpaEIRZF
sNudjrt13AVfcnYKF/mdycThewqbEeVjWHTQ1av9h4CSTt/Mzyo7JdRiG1lRin0O
s0H8QDsGKKgH9knBtQ6hxXXtQ5bvw0CGLHqKtLwHFOkm+6HmRPvUQsDWVU2qLgdq
DFS8kKqU/o1cauIlNCf1t7skTh+q8KitWj9fOjaFjXWbY4PDH0/VLtfgIZyWZhIK
vQbdNf7WyhNTqVhpg5/JeZt7zWOMBqn/R022lutIhFRR96FYnsjaw881Lnh6uhDu
Sxn0JtQiD5qxeOEzK3XyGUx8LIIk2rqtdpo6Jdq0b2N3Ks7YEwglUiPPowerOf8D
Wqoa3UzzFWAq20p0HcJ3rJCQvFFqCECT6Phvrk4dueTBIqWmQXZNRGSeBTpURt+4
YAkRqecCEdcVlDYCNanlXg4OaM880KLmOzy2qh3zzhQkp9VdpQVzTL4rp+jwQOiz
06eUBTkJXBsJmOsiw/3JVZ6juN23+6UZU69aaovQUy005rGMnToE3m+vionkuyw8
ua3wi2zLAHNoUvzZZz18dJxzHmCrNJz9e8GG/o4g+RWk5YOWq6vai3wrBtavXBdY
YZPyJarUjAXiM+fUfk92ZDRafIJY41J05HZnLKjxsltNH+YUDMs4IHUXHs4Tcg+M
siY+lCRNoKsNebFrUlLzxpxSnAHLpq9MWXxuwqZZPiG9L1AtpnPdKXA0G+ieFkX0
Ge2dIN4zbvDJPKR+u6Vrtoks05OKsp6WYXrCPMlvW0BEh02oC1//9n+CWYSeWO9G
xpw2yz5Jr5HJL/hVGldH1nWMrtSv94KQXSPL8uRrOqVAY2Ftqj2S0W6fZ17vx4VU
M2rB5PAb4ycA4ByRMIrtnsv8YuFPT635+iszxKu9JQpXwpkR6HJpn6K/XGHyaSn4
L/7pLjAd/FVL9C3vC7uKZWDnV/cSD5B2CIDRAPZYrfWpJ3OZUUMa9Ld5MazXdIx3
zBw8R6kstX8vsi5soKvrCbuaOAXUQglsVXzAW6nQ4POT3KlUF2epGWrPS5l0NbZQ
yO/6rXuRqkzgpeeNr2l68sVk4fJssKW36ugFOLc8rqx9BCSetshDjledHlSuvlHz
rE8p1znRP5+UFGSEZwlkoiGRv87Nr3c/GZPLntZMjkVEPJmk1cKCXMx36Kz8b5Gb
76y+xF1irkJWXqsok3hX2t2P6Wu0C1rrSdknP+0lGtw0TJgMaQCBtSE1mVVFIQiE
+qHfnqnpJ8buLMg0cXA++KP+OploZ8g17/GpmSCOwC2K43QwVM5tnr3zYewjxSt9
B4J6OmZ/tsGYveGMt3TGpX3pFGMRAFZ40eLerr+Ud7fxKG3BnC1mpqRW1//mC4+V
9lo6e2CerYtFvjP84UMVVr+Z5P5YMhu20pHX7fT2SI675AVTy/Dt7/d7T8nS3BJ8
gFrT55HcRPQyOJf7LaJX6mnq3x0gqsxdvvNHjZ4jmdcbWLG3PG45e5O6enQEdGVK
h34jMyLKKihNmiQNs/Tu8E4zBjqrMjYamciU80n+mFH8NH5WhS+LfPRaGqpSN5MR
UiwUIHI+Idm4LnHl/k3hugQSLrWqcTKhigrECKlox3YUyQKpBappfYFy98/7AqbR
HKNCbkbZM3Y8jRvxl47Y/WyiXQorVpWuNppgpTX5GFirDsx1gFyuuAaybDEG/Df1
6ry72U9AbiufrSb06L+adQL2vBrR130uZqSBjB/sz6Efy9+e3fyTMZMZs8p74fIE
BtB5rcDgEV0XSsQz0mASiLpv/nPcZxmjQb23z+q1un/M9+tfdO3t4kk/0JdjBDOl
fz0mrBoFlmj0aUqm2aJw6ipU/xayHFRMMUkBBi0kFBreyb0YKhA8QP2qyNNK9mT/
sazKMUgCH6UbJzvyazeBV2FLePEMSOco1W+DTfpBvjdSRdpq04sxq2sPCypqomjm
XAq3dHvhcn3CcCeWA7av2EfWcU4pHSru0wagKKJKeSELwgCMSLFNsI2YXznCKOIO
lYu+3RMCsDsSaZoB2glb9UJqQIWLd9nkmu19msXhs3YPVVjWsl4oNlz2hpb49ZiS
plV3zuHJZzsiGoKuAzffBOcynj1atbyT4bidEfkyC5Rl55mX3HzNTQj0x3QsKyTJ
6aRw5hgbxAtJSQeOc48NSoywVw/Vzagt+vjHYikY//y/OWDdg6UTtDJHdgl/mct/
LcBspAwK6koEEdozheIIX83ksOsxQcBlZ7bpjTVWnTgBQ/MMF1bkiOs0VRmA1BFx
WBjkHJqs96b7fbQf0LUhBFdvlfr3TezQVlBgdq3SvhfEVQGe67ho4wn4e9bo51L6
r7WyvrwrofuSYBAD5MAZpGwuEeYaRVatHjicb72kua1eN6H0Jo2mk6bgFVJI2Erm
ePECJQ24I9u+FfpEurKuUmn8Mmgm/bLN30ifSSE8CqMGHy/adLo0FfwALbuv9Mhx
rvxosDreVuWEcCYKeb43OAY0AramZF7XqeihJQk6nz67gPugcXtjEwq4/wFE3oVr
kbHkgz6tw8bRMt7yvv5+FA8wtMmEfSdYkTvhLIXWWIwCp2ag+yPzvhiTKVxIY7US
DV8Z+SMc5P66XCCmnBeMLfP2J4pQvm8pQHqiCMDB/3yETX/9MNTSsPCiZO4X48FR
WbrKzBGNCxT6ih11Gy+xWnjTWsqwtN4a0UxOHybUx6E8xIfBCX+FBpnpqZKdmW2l
fq2qZiqTpr5PjbuzcSUhGSo086+ZWnanCGA+Wg3HVyJ4Zt39VpHfkwwBYG151GFl
3xdlrvuvgN9R1uOWrkbb6eRXqRkxRlfGXk0GDNPMYLXwbWEV2gECspjEFjiFjtrZ
E0S6GxOJ5Px3J2FbrLEz83MARqshyBUUBeMbRCNI2ChkSXPVQLV0ZSI6jPntYhvP
WDaDItLfhmBM6kNBWfMRYt9PaZ/bwgHgj0mYgp4NKYbAqzACYAgUd8oJ7srTRJxT
lPgVIczvi//buramBOGw7WRI1jskRezfPLZO0HmQJF2YLKAFrUyB2hJarj8p74lo
Tb4JhZjBtu9Yo3qAruOtbechlZrflgePczBKEPX1/yWxxLMNfkY3l/kOPHIUkrAM
jRed4HkTdiNzzOcQqbFMh6vwIEUBO36RSt36xtCgR3LsUNUk5h6lCkOQJ+ZQBOPK
/6cryb9UZb3EABhzIwad0fDMYEzZskme7BgFyV9kF4qh2QKBUByg8T0UVF/nnqS+
e7BFMIc9VoHRkzpTy/nlTC04Er2esu2UmoidYdeyoyOEOQZtdXbWsPgrNT+gk00n
J01NkW1VtaISUK2kRQh4upO5H49aBBW+owzTfY/6nSqKB5a7pzUCxvzNIaJkTN8q
0fbOg15Uz7a0Y3WbjDmPp1tMsIiD4+5m3WLNLl/UBG66gUvyjwohhFW7TPdLXGao
Q6U235h2z4P1CNktLAfY2ZS+Habydy+pOt+SeouibeENeLrg0BwrbBHVnpT9y/FP
Pa5tWKeM8RCZO2GuTteYHKy+qekSabdskuQYE2m/A0zQ0wdAt4dygyk84bYV0koM
IqEoKb7cy33WyJAK5HLJuWzk1VkhDnLtW+xSzdON5a4/TMrVsKL28gBdNCUkFE00
tSQ7CMSz0GC3RA2kgI9wVpXFYywxrA2X1bk0GY/Q/fH04ybrcEh7fG2B3FGnrPdn
Np+pSeS4vL9hZiYzRlOkLCVLP0E7RmfGCsUn/deyrNVVuBA95mS95fzjNQRanfQp
AjbyJKQsVYOwVUMywjZRdvfBXK5MxnlL+pRZKTia4GFdmD+fxNUOipIkTf/e9ETm
JUH+1UsEJKgLvKWRhaFduAIBEtmKA4reQAzasfzt3gheIUrS4uarLtULBMof15Or
bz6fh/PYuK4Og9PGHaec09Rp5KxThaHLjzdZMBWaJImfXYffduzQppdB0tCceWJ4
I9eDpBh0eWwKU4emKAJrJBeBAzFXkdgS6eCtxA7IcjCyGK2He36vptt0QJY2ogiL
qFP2DzW/RFH4C6OUD2OPX5OyW+Y9HeXpZsFBGOFA430iPnM2IFVuJHqyrFdo5CUq
10OFt2kCaKNrQIL0hhqyAjyOjYqLddhJ2RC/v8NO3Ldq41TYBCScgDAM0xSLqYKb
w1i8Q36ezIT+ij++L5FV92aYMIjW54fCCA1OSN6HQILkBkWPKjgyWiSS6SbNIftp
1un6q4rBMYR8Cbn3qPZDIUA1OgSGs1MaRs74ogRG8nUA6FGdJcwtQbJT64QOBFer
9gXBBKHEj8P+F2GxLB3/YOLLwEeQLQOASEW+ln/D8F7MMMLT3MlilERSl2NFpwnE
nWghFDjKl7sFH28YgtqLwbQwIZyrKyla00DuNjIPGBtnKumICKmqsfJkD7iJ14bY
hHHj02F5AIoPl7mbjfB3k1AYRV7Xko1Z3oMZ97wQWc/TMc9J52bnTcpK3B56WBw4
OrTAQ2AnoYXqQpYKTJJNdT1AvToav7uMWGMX/b2Aqvn6HtdKxf+zJWPjaHRIFx+J
rQnweesKOSNqb3IGuwP0OfJGhmmCxUs9bl93uIYB9SckHhrmazdMfzuZqDCUntLR
mka2t6T6FHRKg8K6ALgaZ/9akd+kqdLOC9CDf1Z7wnRBUmBIJdShgMhHeAh9GWMf
Wy9WAb6lmrJBPhjjjdiCHxENXRuMopHohHGZeJM18b9cn7rUiZ6aeI9/i8vOj64k
wxCvTfvkyuKI4IWuLFKmnvbuzKjEqUpQbcSTfTtlsM18RRiiicmknyqGV9Q97pst
SnXtJ5s3Ykl3Rj5xafjSC85JzSKIIGellbJdC+rgwl4x8+OlA9yRsCXrA+1fekfN
zGitiDrDik/+/+oDaR4MFy4hnq6bt+QwU+uOQrHv4svjiVd2x81YcLfZM7vYyLl2
430B6jGBqcLWmb1gA8fVVynzLfFLdEBvG/8HFWx3awDmMXQ9Z3QQWAfdHnENlC/O
AnQsIV2EcYu6B0wbMo6Xz3umtQmRRIkcUX/VB4SAEYWK2UyqPr3PPlw1r4kwNOEs
ZaQhUCdHeOQD+gt+7vAWNO3DxAUqRYHqrk8O5yAR6Jgs+U93vnp4hCQ64Kjr3GYj
efgW+sSQde+hJav1EXnKG92ubwpkdGtwtaZtU/u9TVpXe/6XNX1rt65F+w5aKql6
jFjmW8Am9qNv6X0Pn6n4LbnhvUHlxnmxpiiKpgfVZDBjSVk9edTzoKgDGJCw5Wye
A8Rkgm7jg6E2MQ2MwjqUUy9C5PnlHLB3ICJAcY/9Twpf5LDYX96VogDYtCevS0s/
LJ3AVVuB/dh9hqhH2qsfqfsVJAuMGE4VqxAwsvjSkohFH4FB38g+w3N7fhGZdkV1
G8MXY2dP5OIT73EE8xzxfw85T94Mbiuh0SXUgGlsEWqUZ/SPKF5uRmzEQ+xWbNGZ
Y2ZDsl/ehw3ZrCyu9gxe3aplhbGu+NUP2zxVnegmGw3ulzg6F+d4frbSfB5mna6k
05DyRBYJGN80he0qlkts+IwNZt7TVwOLm7jbZE5KBwAAw3O9idbN8Vt3BZCwffk1
V3KkSVd+9zzcbrVK1Z2ubpzet+NyBqIi3ZAHWyRWhv9Z2JGhv+eEolSMWmrno6Qs
MGyZP2EWnDorfIM3V+Yn1iWnMnjOk7Ux/IBRphOcNOwFxgSmz0kY1Z+q1fxg/D9/
KtIZjuGKb9aw+fibHXkmtIi5o7u7BH7CYkSCuNgSxj3LAKb7Ct+Hvy5kZ7DFjqQL
TJf8gamWD1C/SqWBE+0gTi4yj3bBxao8Zzpw/AYHXUU1U2nhovnq5syHJwbbyKq1
W2n7t90ttD00XQ1Yh7xY9WcmdT9WM92SuA5CJVy1TFzLpr55+DfUpVHSZOUQtV7o
cH+6hzyuuiyCpnF3xKSIFlUA+PsNjc4be8ay64oHCJgGVQZmAZSdGoyY0P7HrOSz
huCGYcEjdQo0U6vgGb4jkjpIs8lkFdSDFyE08FWGlq5Cuiueg20nh2l2AR3yL4fC
nWr4scckOrJ3/oYXqnRm5bC1fML7255/qDDxQd3ePMXG71MkQomgdElCBVPM3Rsf
9RWS4DFI1WXWAuGzaf8kCqW1j/nSoac1soFtE8gTdo0q9yRTf/UqSVHrlXylBGd4
66v+YtYe1JfThe3ySNE22cOdfdGzo9WEqJ0uFJXWLgGEp6/bAM5ZKKbXvmHbvv87
Y8vBLSNEyESSchkkPlilbiMQFsjO03pQtXGFH+auzpcPyVH8XcyJLOMqhSWztzi8
uGsQW63jxtHaD/9KduNiSiNbOl70e+381yGt++tGxoPuVj5Cfcc8kmybyN0TRd+F
G+ymJbGj2XrLC/FcIRtGMC5CK5Lzi7x6V/UABkD9KMVCMIasd57mFtIUxHZwlhfr
oTFPPeutR9bKyh1dqjBpQCLAVaipCVuX94RMPdyxUOPOmP8oN+jvyBPVL3GmivS/
XjHklqUIfvuPl1IxANF86o/UZheh+wNIqY8VShKLoXL5Oh/2SdY3dPSuLupXuqbB
x9Dr1Lac7EVEttuV7Bx81JJX10ZjYsV482I9CSHo1CcU1u3FNOS2QId9orrf/x6m
xgW8jVO8YHe9/dy7PI0XfIf/hY3HnxbdJyWZjS8r8a1RM2lG4aXyss/5otcBWhiU
jHBxBs6coOls2cPRKWhxn83m80Jd3/AP9fp/y350RSLdgAuZS68EQ3c6fBkeAiBI
T52hWjsqVL5uLOBk1UdCc4OajQvCosWeTrSxUHS/3Hh0ATH1ky0by1CsvyaYEqrv
ul8rryDcSOvlNwTpJo+oZzTiTEmsFaKEDkigpVVzkfQwSQ3PNMgBRAk1olspqoIL
JqjsBounNPjaUP05sMWO+4TqfDq5JjaA0watnywZV0swtZE8oFw8/dZsytgluwBY
ylCfMrAztb2HNsIv+759GZLzOlibGW+JjhuudIU22Bshx3RuW8TccLG+Jwl6gdtZ
pQtYpj+Bp0Hz4F4PoitV3s2vIqX2XXI1tcl0baFBAtVSIh4MjVxlQDvZc/rASrSN
oPcgzVEHXUVDDGQ9bVYVxvBaS/fWk041NiVQftFCwd3iv010WVnzLmU2XrViQx8B
UF7/QsvKfrzYT55Jg6pzFCJ8xEBNTGocIc9rQZ7eFI6DA6qO/7itpKBtSdpigwo6
TOHov9+c7b4UrD0tTb9aRyfkGEnzBH/nZxjfv468pkZvFqXFrw5dFsag0PVAlVX7
bTL8LjeCAhZ3vVYr//ViXK65LUWQ8jtYUD0UcjuH+Dt5tx0Y+OUFPT5SBLZFq36V
mYbjRmhCxMVLfs6DNtcFsa30bayGzbTnMfX2UiJW5K+XZlPFR0sRTem+7e2RuQji
QYuAwIU8xYmmtsqlj4ENKKfxLz8WrugjrA3sdiZhPCcEhPiHBTAyV0OuqsDgZ4Yk
0QrUYKJueyLfvk5rt+M3I0eIH0aerafWv9hL+RYHqsY7mJ6MiQEP1A515LCxcG3H
UFUygiiAK0IfQihCHYnqiRXFfWVsrNuaPV2sovckGeuQM0/KNWOdR1PUpxawu4Mp
44qplOQFADRdcFQ2Cc3dKOsZ9aHbLn9KnKfDFZjAxbST79xGAj/Bd+c2afeXDZWD
P6Aiq8piE1EmmZuWJ0MnQaxOYHBOGozNjpO9oAYu7HgIj/m0t7V7wTIxqvbbr7vk
bDLjHBvG644U6KWHQgYZIxiuyIhx0+yEduKqZ6yWj+iaCYe+5iAckuUEzx7nx9uv
B4PQFdcwxX5FMcxayj/UdrQPkaBSm/ILWOIhoRx/VrrIX6VW9xLjPq1gVgnuj2/k
YA0UChSBDQM0ApWJKfVx/upI4tyGwNM/opbkzSonl4iUraUUuo9wYeznVI2lVlLM
Q71SovAiyvhVljDRl7WAIhNhxBiFtSZbVFBF6cEK6tzpRT1Kwpaofjd6rcCYVvzn
Z2+nGKP64nYOuWDEblAWYiFbQ/QwpO+d8HyWly0i26DCbwvQVqtcKBDI9rbT0wbH
cbX2MlTrtODmiHEfCgFdcTQZW3IhOOwtS9Lh1R8L14ICoq/AcF1MctvBZqmIPXa+
nIwszAdQMA/7597Uep3qx8RdKvsIxgUfbGshtQjAI8RmRC9kPJtLfJzdwMbUCt/p
1h4BxWxKbNvlxgeKo5AUNiNgns4VI/96Od0HSG/kyh6JxfKexb4KGhWKlTDToE1y
wLbMSg2WGHDEkz7aJTK8qfnpyy2XwLDbOPlNhZC3ACxvPHZOogquESTevlos5OXn
5y9E9j4+tJWtj3ObcoG/AJ6nP+glwGuoRlxWrk7UpovC6o6aaERbeWvkIX5C1Ezg
AI5RIsvw8YAhq77tCehZ7+GcdU85Hq6pp4tw0adOL+sJhtx4WlsJWzAT8TBSsF2f
FHACapczMfLwQ/FMbvA2zE39d1xjfx9jMBvqZStUU2HCslDze8RUk7YIpDZRvVZp
o4vS9m8/sXPpfvlgD9CgMyEePXsPmmUxiXNyMyJb2TPLNJKtaVPlGdAagj/i566/
gWSWonfEkTqBC+W2YwEqxcydTtM0RlbrUSn3NaaPrpSlpFmOkJ3vr2mI3+ze381h
vmrr+cCf5krODCnmb0ssX6dGJBWObQghE8idzMESAUJLCvUKRWwF8Q/VgnflShAs
vzokB+OzsdjV3NgBRMAStkScBXy/3jenW/Vuo4FB3//V5pFgTJSKlfYi2TKiEcYn
DIPqlpqUdWk2UUgppybS0ydqJhEF7kLKvrbcWlxFZUmQM3DLPfPmJ0O4SiQ8o5yD
Vvrh5MT+cLifMnbvhOhy4llW4QHUHtkFrtR0wWOZV4f1ipXqp9vSd4fU/+KSu5YK
OyDEEduT5QhElu1Ppf6yRnO8/Bgfd167Q/Jcq7D2CBxu0q2EsU07y5+4+V9gJJDf
ZH0SD8ysGZxrfbw2SlYXeQw0yNwjSlBqTlpfOboZXfMKpKH70uBVWx75qqlpz1OO
JlABplxVjDpmyKdOJOuPGy0fc+EjhDxbCFtEO+tN2jbVxfHexUBTcFXI+icCdvYs
IF30Bz8ZzTKLiLrHiq0dxHHhx3/a8dNIfTR/AKcv6PQNOzTqXI8mMfvMuR/W7+g/
5U+Bl/W0h3quZFCcX45iFp290uGGxlpKwK8YLMyyhH+2nCvqnIGdF0o+itHSZx31
8n5xmbHGdpfL17z0zOdFnps5fHiNTXts+ZnxslVTqi4l3l+bV7RGzabyEVTG9w6e
MKMEXnSfmyYX2ceYJFEKQFVMbCWsBRZu5c1rd00v0e8Be8WBJReDcri1cajONGxi
m/ER745dj7gbPBUs4lOeVcLFjes1ogJAmpvb85Q0CUXWc+DkxlBRIV8YkTvu7/ha
w/SrnE/1zQ8o9HelOfzDCaJjSH3dwCIyJhm/goztivIN3dYQQkI2edr5Tox3s7S0
qxYUxpClk8yenkoEkSDMvp5RCYB3gd3WpgUmPkKdiX2exog/LXHxAl/Bi591aUTh
QJnnb6WD8PcymjJtCMFBEqIZBH5FH+tbwDJhr/+Zt/b4UDNltldiwf3bSHb+6x97
giOUXefuU5wjxV/+lko9dc3IcVA2lvDyfHkvVxOxuj137XyvqBqiAf2nP6AYyHpE
OKfeOfQopHyNbYGsSJkMOJFp97ziEDM/do/9XGkHjhb0TzAv0AJsanGzBm+Wqj5i
+5nzyzhR5c/N4FRYVj2tedaFEochH3a4ltfyNSh4qZlQrbXdlhCMNbjum4syk0Wo
t5Rby0LsJPvfvOCC2Ymfyii95sfhJ/5gGKGTiCyUYTeR3jqGl6k7FFH34YB7dClv
nHdKP9pVZd8e9gdYJ/U1dJTVLUnoO+/BhL2VT1JvxtOcKJZXoW15jbwM1xe0uhUG
uHAHtGZ7sEpDbyfKaxzB5n+kYTuIRNvVtLa7u21U79La7FCfTkBHD11QcZEYxkWE
0a8kZCCk4vbUfxUDqOQUQBw7dN8tClYQsUAc4MI/79uCeLnqi8xiKlOdab7eeIyH
OwjJZMG6yWlL5snjrTG8BmjPV9jbyGfz6SnCp9mpgUXoOuGq+EIn/b0CDiPXD0HH
ASt/ibv8tNLV1Icwcizz/a0JoF2olCHIOyVKwFd29hEzsFY8dYdumNK4uXnvZPsk
ggyh1z0kUq+zQovy3qdFiDWl8nFvB5Q07xOo3nsQVdB3VANJlCF/SngPJ8crmBBB
j0+qUph/FBocs7BSH1paFIND740ubXaWdhcV3bVU895u2bluG8XG5O08uIVqSImE
/35GyxvlOOSREXphNIwG0Pkxsi5EnfiBYvIACtZuhVQsZ1XEtVRWQgDKbe7GV0zF
8rO37sdE8DNVFDQtVyHsuAyS3dPS95vvewjl35QjQCI5k0siGQicFvs8EB4GPizi
wuqvEExmPly2OP9g6G0yaNH5nbh0sU8U1uS+pCssXSDDb5mxkHO/ULC/fs4+u/JE
wxo2OoGiZVkzaBV6YmxnNXXmwCRZFZd6YodGeEgTaDvvIAWYh/ENjvUMrcDSPMhY
2CDuZ1GzW75/IbMvfIiNeEbjN7DtHrFoS+Sce3Jy1p5NdO1FynaQyskEMmTdPwem
H/ugdxEeLZLRFZeJGdMyXCs/243OPA2n7EJ/I43iIVENtgxFK2azj+PmhszgD6KI
dV3MYBK/6g060NfVuiVaEckbJBnZqs0roYXR5iCTmrYd801tir2rUHNKCJkYcqlM
9HiIMS01YC4CWXVGlox3iqYbsElY/MBCH1/RQMzpvAA8wHdhP7QqXpN4YBJOTZzG
He1Awhx4SLfp4Wl4bRYYwiBW4P0yHH5MnpsUboLdJ+UN8Stg799ub9/lHiV8o9fK
w/rQc5FeVKmVuFivM92vVKnejh2wDAW+MgsDW4crD5G7KrEAhaAn1PFxJNxNWTJ7
5bvm3lFbgpWYn7tUn+m88BGYC2g5qEgmYPkXMaB6tj/AjENz5V7/ww0Q/jR8hNTC
DLUyooYqYL3fMc0Tqq+HeJMZydVJlpBkngt6xIcuZLUrfqKtov6RWG4vMoErG7gx
ZMuQcmS8vU6/CX9FqDWGN5m2XXyib3nmiU1QcJ2tTPit0XvklYvN3iiUyEx6bKKe
5X4V/jklmFJoPuKvPVlHo6ID4weNttXJlYUjszaNTL6+HCmG3WAo6mYVbQ584Mhg
mM6SrIRqucABDHJDUAkSKo0GvcUFXsq/lKb42AIrxhot0mPN1QRHkAnkp/wfFjvI
/25h4pNYQQszdPv5oWIrd4vdoyQzYHsafFn1bUOF0811I2M0uBlHm8Tarx/i3ctI
A9VCg/8V7usVGjIsg8u6iGlXv/n/4ox8bYo1WwxlKqI0t85KOxTRs+b0SIJ9PrYE
xAZLo9FKqwPnyLD53teSW0WinUSVWvIyjDUGFNnvqsteFPqXLeZqSGRk7l5gq2Hn
7o1v63K3MizW9i42nzss8yUGr/IOZTpo5SY0eICL+Dinv3fr/+4HOnyBWlMZvpG3
O7+DCh0ji1kgg3RL9+CnpKxTs3GLD11Qh4xVkg3NwFwApt92DanA79p/sOfGdRTy
x/PPObq37mXOxfXRptHcsYkk+2ob6RsENceJ6kSZh95jhKwlua9C3iKUQsCeIoLQ
uNsKPHHlINlx9JjRR6saAKLquWuOUkBiVpbqFYjNg9vQnVDB+yBSd+2tXhF7O5AP
qzeL2j3dEFDHof2qFILqCiPgEWU0AP6YwKxnw6qxXhxj7vZUwIRt8LU2+8toysX8
WUeUU9nm+8v64YLgp8125dHMrjx16iPRo3vPOI787GjM/G+aSlwkrRXp6APBr834
189xfCx1Z06x1Y4OCEviD6gR1yT1K/ACQvjW/YY/x4lh1pck1BkNHDbNyrTBMMUy
UCg1DNserqcwSKuC63urbaDdbbeMwtgYlmQRAhDHPh4QviMBpwexa/0fVSvHwvq1
eQ7w58znaHtEvBxx1E7WVIsIofEruW5QbkIs/LZQ6WoatLTFHOJfjpnWnwv5uPRF
1vEaTkaHDnHSLTcXNuGzXxbXWkqKhPzdKwQQMrYcRzhiLfUwQB1T3yufZHnupdPt
DobzeS7KQ+ImPySHz5YimtLzQzhiE7C7kw+Ylr1+wvaVf7+tGLDVKFQ56/0qfIC3
B4I/lsHaaabWqFN3QY0oGh6NYRkaaPKIjYh1pfZIq8wcj2WYQknuVPwi/VYx+kO3
skEFtp8cVRqOJ1BaTzU6soxvyGsbJFdcGcMg1MJ5fdICjr6FxJkQZo54XC+1RDpQ
zHg8YupYonPBkjBj+OQBEIvKnQsiSV3EH2HKjugjna20x80IvOFEx8XXneZTYxqP
q8Q0+DSno8OZH45vDcyGNwm1AO21QSk0PuB71ZKbkAGDzCijF+yQjYTt72mxyRv4
72O1vukLHTm/JpotG5JsTv4u6Ve0NCZBKtgXDSoDgUhqvGAFMskKLw9nuia8UCDj
rMB3WZzqwQs1qxjnMFULNwQSbkhIRIH3C1HyOLm69ai0edWqu9hRiSyZYQwxfNfD
z39tVL6qviDMwWVtjjJJTBK2YGlodNogoU+cKLxZyPkJUy78QPlmmEcuFlgkkt7O
VSwwfOZi9Tm8ZmP+kZvh8/zTjdlueZfLBJUTn4AmnwmlT1jMc2QsqOqzqV1qH5/B
/EJ/9Pc4A1bLuaLafguVnbzWXssBS2IfiZABNCZEoiZv3dbE9N/vI86l9sE3RIHf
DYgNTdLFE5wo734gK6HD2p1gt5GqCUR9eNm//QzAlP3PyTING7G12i6I3tiuR84M
0wb24ySAadR7gRGWMvRVrlgzsSWyFpsDa53s73m/ivUGAqH5zoTvQmdKiw357Uq4
XOEiyVc9T8kkOM2SyH19o/kuorThcNlHuj5xfpbQ4qfnIIt4KDOz6bpJ+/BYvC5B
9AMIMQGtysnVkSgzNpC19wEgKn63ltUNmtaGRcQUxDdaRgaGNUr9Nl0wI2n74HxY
IwV8Pfita9Klk8lNtcBS92zQiMNQcwood+u6npDlQ1Y4F/qFi0cUvJy6eN0mFxxI
zAM0MgxmmCbwClaIyIG8UQTbuLWWmNorGpAC68kg3i1uzvSHGhRlGZTjz69A/9Gu
rZXmnl0Mj30DvTAUGRbNyDOk4ttWiWjHWwznq9G8g5cHUNeocC2+HQLMszrDptkq
B/JOk2NYJw79nkJCz4StknplcqJJqS5jJ60fiTQewjbaf2G5rtZtF0J2mOzLWOeP
IMZQB+ti7K5KD1ddblRtp432wWKjz1saU8d3dz5VxFfGur8s+BoE3ypuBrOEyjK+
GXAim15d7IhvT0WFGA5xpSiI8igKsTPBCL7VO9ckQ0OWSSnpc+GeK9st9ZOoiUDJ
D/g4u1nzyIVWJULHA5EsVmk3lDsJTv7klyUdD3haQ/aHyGsaJWgcqt/TLl3feKIk
RyYyEEIc9xytGYm3Mvzci/f9rQ3FrP8aMHHyAFcT/7F1iAYX6zYNDmVr8lXblFEi
hBQFB15Lt0WICrvZMj4y+XtwrHSfWQV/WOCyp5zcM5n0a9F4duTj5AORL9KG4sRh
rM28AlIIWWGaGU6ayZ+KbJ051/DtIiy4AISeuILgnrG89R1XGb700h1/VYZZV4XG
/fCC2REVzBkmDsvRYl9NkxJLD6norj7fa0aggLb37IvaZNEQwccyeb3g0M37AOMK
is8SieG1y8HNqUm2xhoVgSDp/qXfbHSvj7unwHaPcMGIGJk9byixFtZSGI52IIfP
w7o9l/LuB4xQnrraHiaAaMlN+pLKJQwwLJ3CQRn+q1l+tHEnZtQEwkftvpZkmPiY
UlCdOoaA6pEW80l4d3V23feTcU05tvjnSU4MyphqrdIJSaJ4HJOiP11O+2J1YONJ
Fovzns+V2EyI5jWjuBvwVA1UakC0sarTyHCwvJ8uuZeVxqEuQSmhxMpu1DK4Be2s
ISQ2ufttu2m34SYvB5lSz+7NMmINZ9+bSvBk42PmvoX5jnC4ddjEKKDP2gHtn9Go
KZAfbliEvCdjNaPKXiUxvB/1ignIUBU1uL+YKTZaJXllKWQZn4qlMJsWauHIaZLI
8NImO2EhPvjxCl63Bm23uvHNNT7RKWubLt9g7ZoQZv7yi/WOrItL4M5q0JS7taed
Ah5Fs/sT55Ve/of7hBqrzldFELzl0Eth/RAoxG6q8wBxxjSqQtXqblPJ290NAKXX
UVPBv1W7KtOcbFlG3DXSyKh0gXFgmu3nFXJEnp2GUq5ObnswCrlshxWI17JE7BAn
yaOt2V69RoFvqiDHDbXUa4ahl63GGZmBw7aMbALmjUziCoDeh7Jsj1Mm7/5NPpOn
GTkOlKoEqdRgq/bqNAXpwl2G4fTUCqiT/U3ssw/r8hk/BFpUUr1XpscsXor7seKJ
Xa6UxOzTOxejq4p2t3d66DwOECurdOPszESwHoAeNoha4M1/CYQuRXctmBSv0IFG
3auw5EFhiJ2BmWYF96oEQXqMYqHWAoDoS9N8qtyJwpUOWHtQPmqtrUnSzYjS3D8/
zEHqeV0sCxKuwJj0z4cmAKgPleX4zp+bgKwQO+r7myoxFrE7HZbfQzhKcW9M9OTB
Q+DSnKgzqYfNpwqnQLiTUYHFRM2blc/OZd6geBzQEQKejSnkxLC5tsFz+u1LOV29
DGgiamgFLE69CPZxCaZgGXsZ5O1yegaajLCyhjZG69ekuhg9D7rbcGa4TFz2E3+i
eSkmjV/3dvNW6byNhdMcHDLJDT6RvUAiwIvDglFANjUoPnBImXJIDnrRSHhSwq4v
viYPA98uQ9FTcDRVPrw+prOrXzJr0RwgvXGD9ViCSJwm079s1LONSSnNJ2OTTDjt
sL9/OHVyl51wiJdIKDmLt0Ve3d+v3ILagV/R4lph16cP3sNqwoPfX1P1LUl7xYCD
+aHLsaYOsWOFlxHIndJEmJwPk59gXGi/MxCNphqlVUm1d7aZFPjaGtAu6jeKqC/S
LsilNjC1FrsaczXWWFLCkPIrHKtQN3BZh3rIhDdVs3fFmG9C0aqyS4mrhUmUuFNa
3fOZCL3+RSxiU+tGoNJ1+s1LUc9445sboXGuSliDdtEao6oh4fGeACUwpu9aCa1J
RVlD/5ghIwoDnI2EHIjDRwJUa3TxcGU8ggWgEzPrgJ4iCVTJNSfuJBROOZcBw9g9
zeVLfU6AaXKVQiysPeKVwpdYA6LKKzJNapp0ruBe71Obt+q9DrMb6/9bL4su+l/3
bZ92KptgiCCs/DsSU+R2Jc5/UykFafLaMrP6Ufcct7m1s+3b1j9O+QnVWgVkx5vr
ddlHEOiqW1y7nvOSc+5S0BU4wob6N5DZqSpw0lHTZzAjZIEzrsFq9X4TAC/u4IQI
4qZ3pBRLTkjSF9LnGT+IfmIBNwkmKV9Nem3tRoaKDrQbabCRLjjdApxnApA8RDgs
ge4WkgZTWREN0gdqSWjYaY6eygp3TqKxAHHrcJmU0GBjhsVNRjjTxZ2gwTdSNqVw
h3Nrdx4gqS/Nj1XAxhY15+oAGBrwXnI5POl0Ph4EARH7Dl9bRBaRssG4ZH86LmWS
MvJSSA2E7kYEolzt5Vs7uDzHn4jUlwUrVwollHD1fjzcWLBJKNajKPyFuMRZ84BK
0vh2iJTRCoDkjJR5coKf+7HMpZbqS+dGevEesTBmivJyDkotbj6P9tintRh+UWDU
EJgeNTGw1suL2IHx3HlaTgAKrlCxCZ0ugrHhuEeFrSl/U7szzw+LAYC7UW0mNHx8
tBW8WWNTJAbNe/zRKUB2p+VhOrPhbGdkwLZ0aEAZfSsoPjlY4Qvd0ksB5PEfEvWa
qOU6hpzWZeXcCWU+5p5qbU4P268xfYWQixKcGuh2l/lzvMlvF6AvSH58+Do0bkP9
7WYxGh3lyCHPs6G5jVVZsy8XvFte2LVvcUOscrudh5fAL0X3NVC4KTYXlqi4wwbG
caJqXXN9EbpeqXxugmcjeyL0j/9gPqZNVeb9MdWg7xpSoGOdYawBMWQkQkQu6BZJ
FXByfzoMwxtsoUPTHz7hmSG/RL33dkuniVJk5rWpvyBLDxKr7/Ph2voMRPfsY+3m
oztDj6OzuzH+18TWFrW7anqxz0BdIcG9rM+4x9BFYTMBzudhycQ0yvBx6mXcmnT+
v+TIIh4SkH36Ye5crHnUEy6kyuuZA0x+QBebv9KY/IpLzUX7fRfkc8HV6BeDUViO
iQvov/b+Jl4OPlNl93T6D/OHtZXx+z52xfOi4xoWLW6vOOxEt2eDnFe3BHDX+N9U
+C/eKHY7fzXc9s3HLvDP1CW6iCkPWHD5pND66Torn981Gkt20/D6GpEJAMpFAG7m
Cg04qbx2jm0P61oZEE8aojhKNVW2iGU4sqfbcG+PJw2IcoD3tjM6e1fD7gLIG8E6
YhWzr9cC2qFiKHbap6aGO8yVBItztjVCf7Z2l81p+a7cu31Ddc+7dOEtdMuAbaI1
5YCtajz+3peujTS/j9M/bu3tnHAxN7dPMyVJvGvFoYDYxgJ+q2ajE1FsJ9yORSY+
Xdy7sXr+V1lLzXX26P3EvOjtEHlrEPqCfDbiabYPb4w3LstWjkZ0tkFSHL10wIxp
cpjTW5PPlPKwi7OS61Bp5wdOjn/WF+eli4NmZCFZclU42XMSxeBsmnyWghhMVdLs
ujxzREd7bQRdLKd2OLL5S0zHgrJ0wweAOiFeoA/LOEI1Ddpyu9j0aT+/bWfcLSwL
zlpcCQA19fa9Ux3jI0boET4x7T+29uiVnJTicJuzIetSRhL3UjL+GgWzAZOGS66O
EsK8O5fSjGqYTeuYMmgAYThTm5EpwdZdL4eH3mrR5ia1TPyuCa1K9pTF+W6nR7Fz
qFtEL4alq7YZo67uLI4PM1wiWULKVDI92/M0QqDUQqTgTk1uRcnHsa1KzoNtuh25
oyyQK6SA2NSlu15dwFVp7XwVIv4nugYOT1t/tSfGUXwbP1H+1EIMN3TOY/dyRB9k
E76lNCALmayIlY9gqPVnZhLDtuB+dRreoTauFnN8Z4Gtp/k7Lj300tBMaEg6sFe5
rucS5tOfTZl7xIaFpFbsR+i0RiFZSDXNL25iNcQi1P9w6w1JdlrN+JWTdPXrBrCR
gt4aTTYVc5U9VLFlXrHM59SevQaCzJJ2nWM+7HfkQe4YwXVlk0QmB0VGBbFRBuCP
ICSym7W7k3G0/wxO48Jg1sVWmupv8p/tEtbuzmbFnWYDvS34AeJMiGO9ui3xAPNh
AfZaAk1tl/+/y+l73O/kjuPMs3GZ3B39hD2FY+0LHSp9ME/gP35+H7WOYnF6RihC
Q+XbH4g9o8eUbsBM/LqOW2NYIjPoq1HVjb0lUO9x2yOoOS3zC0rlnWuvtKtsRjrj
YW3tsfaRmyqduwPzmAy+/Zy4js20uO99RrCodJHnYByLwR1f0Z2b7B59jKfzektT
cpwQ517rZX0OUSDc28PNdLSlwdm2W6FNHeBQG8jLkfzj7XWrTO8/b1wHLC48Tz7m
nFiPN/8P+7kPkDdEfhlzcSoI9AJe0kwLc04L+MUGYWpNNJv6Kk2kK2DSPyBTHpQk
yVe6vFimlQTygqz55q7gtUXlASCVodzuJmxvtasWJDOnRDwq5M/XG0I6rzg/RpPP
i92I7E58RnZAgPpMZA9yd1q1tTjsl71zgDlyxplJp+RzH2FDmGfWuVtTLTTodlAL
09Z8H6F0tVfFvAD0MUR8z/Hw4vJv6eBLecXU9jngm1CN0z/dTevRpHLJ3rmxIP8v
Gon2h7PbZjnlvhEbZrfxGK28pSUSV0AHDAfX60sl25bi3bdmOfSkyThyMc77Ru3g
Hv0nd5uRJAPyFO8RA6bogOZhXZtHqZcEQWi695rLVDKbtEE8EmvaZ+lPZJ/p6zo5
VLguoP0YDv6EaojHFo6D2AEzj1M8Hpp0WK36t0pXrWvQ615RBU3va7+jWX7iWnwJ
vqI8BPggj9GlCeRZAwU2FHKfBaXyVsxuzF0BKWl80LQ3UoqHehwsmluDzvOpYG5n
S2SMTx9z0NmxkGgKmUboo1svHGWZzngKfsau5fV+ix4/JMoEvzkEEHwYSfCD8hqU
rlbHKuVcSXaZhpA2Kgsh/NV0ZgvZwmiSfHtEEm8yCixiR52AvWgq8jXlwwCQJEw8
AymopNBD4kEu4kYpZUFpytSiZSTipVezlI0cY8EFdcs8v0q8Qb5Pboy73pgREuXk
K60yDgHPgfq3kM9OzhoJR7ZzhTb7kKtJkJfGdcnYbWkOP9J1n7ygmtdo0LrDONQV
lpJubonhyzf0uJrmH165V4dnoBBON786Zj3DkE61jmcKaPje2mttjdJ1vgRIwSuf
+jOg2XtmlLA2W73nFh7vsyKPXOTg1aoJlP+GGyNlC2y8fIjHFXWKOCY+BLChcZha
R3li9Qdj6gjwdjo/E/7beF2qtuRDWRkTuXBGFXQ4nYlhfEvyfa1AzdRhq9kz9qdf
tRtJXn15UWF7V8AdWMtt/Pkf7JJ63Dez8WFZWID8cIC2FFJLfwctDLbxh04v83A8
YCM/moO0kA4dBZJLtM0pOo2+UtLaKIKlFrMuPkbt3IdFg6tmdERSiNHThuZPVQzN
vQkE8kejTmMR5u+XWn2cDUfG4qqknXzQzXnh055nqKeGkDwCXydKYhPGL5xiMYYH
HK0tJbxK7Qr+jelG7x3i3IvbvDY9h/iNnu501WnJ/yWNq2iJ6MJI0StgJisibXLW
kRxVjDRuYbl0zJK1YHB7hRWZKwr8xiRqsiUfftTd9f1h//Dr1Vis0OuBuX4H8amW
CZAKPKUaeceENOcE6GdNT0jgtZgXYMCZmS1T/XyvbmAXODaxUAgQT6b7NuPn0dtP
n3+gfE/OnWyHqxjpL4zvUgxoKZbLuUAGQXQTTVmck5ytFzEkwPqRxq25sy5Vz5e0
kSiHKnyv2xD3kQbNzEx7rlItgLkCDbMSVgB3nRqrTauQQxcfZfbF07CIj3oNusP6
yuelFSHlT/aej2ZW3KrjdL8PPKjs4FZHDpV650wvEre2O7Qj/m24Wrdc/16QbQqx
sxaxqpSItCRExU4qw4suDCnOnykm9WXsX7YAskSWtf0myuYmnVI3K4U9tI/zqoHt
NrzfMIBUOfuVcTSjsWQhJ1xwQU+uSUk2fnCgNkrj4tlOJLC7kwEn/eQOuchtXrvv
rrcCIgHc0vkL8oXvfXSOfIWttN+ALVWhjzhO6scxD3SHAvqQnzrhYl4cXlLAzJyI
UH7LIe55xcA7/K634hXPoBSZ5626fFDlhBb3xDS7fQbtf08gMxp06u7JRRJe21HH
VCreP02lWAFu1KCFe75dXRABnrSpOCi7U+D2ZG42tdJCF9SFxnj8icHEhuu8vbxU
UFRRwP3sGYqWoI9pfKepDLRG9OjFp30Xw0ZFd3hgxEHw5Ijt6ehv8eCbOIUZXynJ
hjcL2gxG/gb9APddoikUbMgEHBVM2SKfIbBOcZQC+g5PBS9qFjSiJ9mJwWXkpC1u
zj/CB7e+oFZlXHfLqHNT8R3urs8fECmBSOG9uJ0+7vPI89UnKAXRqvOsCZ7tngms
0sDDASQGYk5FGgIVoovBqxPwFqHJ8PUWMnsGcnAOUfJARILTns6IcdAScvhiN7Eg
vAtG0WYRVmomdrZjooJ5OyJ2o2gSJAVMB3AXXeNG8Gwt+dA7G+NS5tTK4bn7bkrN
6RQVAII91YjgtvbhBf6a+0zXna1R05LjEH3yDGG2JlHS0Bx33bgR8f6DnPzbV+vQ
z4p9dUUfzmNx4B0Xq3w48/lxcIJMDgd0OddlgHu8ABwZTHU3BbtuSFgq9q9GFl9u
eb0Qov2/pOtEsMhgVX7+rJkJwkKF0enS1JagY3jLLgn8M+ZTHtVyLRdWzc1BsSM7
tU2e1StEvE72lisEOzQdeCDHB3YLtBgEwDTmijiDMyPYPwu6ZfwVOGNoO0j4qrLV
loT4nbEu3qp+d4uOt474Zp2RkHniyH5Vb5YNKJw66HrTGExpnWiwHYFrCVdi7g1O
OVI7Cxp0V/xCgM189PwqgHy9Rt9rDFZaHEk9Lebb+h2y/2tHabHRyKvs198sXm0i
i9LcZRdd3k/srW8BNBRxiWKQ1Mjgo2tULUL0ukV4zerrC3ICzyDhB/8V0iRGfk/C
i9LqCDoesUzAqVv2myBCV9P8RBBseekC3rkj5h1S9etGAyO7IgZAw+kSHrHi/fHU
yGYqEVT9FMbHqRwugEzUtqotlyKe7a0Cpoex/oXSS0Lca8XDU/tkjL5/Erw6EZ9V
iVKJ+44F/8NZZj8gq0KoUhOC7VUh9LkNjWzxPU0LXCK8hm3EqzN3QhSw0dGkW6nP
dy5G+fovGzGfD2z6KyctO1Sp1gTN/14rwA8B5EAVtZhmto0WMpDu2FCE/igl38KP
pph0RKs8E+6kBzRUZVAjk+clRQTNNKBxBh/mFo1+w3/l5asa8aOt0h6Xv7f+zcwF
/DZWDWx9vOjtxxzocQ3zhyV4IX7nw3GPjQlxkH7/9ja2yaHTO2VBh8L4pMvgL+0A
ugiIxGFp6nXg/fXUViibr29HeboTS0ezrkq0f4uizfRb6fDQ6Htgsyqly2PVSVEl
9Qoa8DlfGC+OZRdtDZ1nokINmQKcwiAzoi1kstGUpBgkHBTbjFHk7VV0+ra656dI
phnC1sTk724EDdwUZ57FmA0UIFq2jPG0cmRdUgGWcxGwaapdz6CePJm/TNbhcLyW
dwzzBjHfqCUX4qPz3J67MDC8hV1q7AwWQf6bSwB5BUtpHwe9PGj6RrAOOhSev+Gs
7ddk/rxox0tb2mifrlODJIBECYRkyHUHUTsYcRkriXdrdgP5rIHpcDD6lcAGzM5Z
yyhQZiV6kcmkQTeYZoLCjrpSIEw99mluWaf479ACmFHmDHX5StuvsLqiK20ZWZvp
jhaQUEGuDUle5mI9PZijjufkL/dVf2QwWOb9+LIP2TvJvHBBNoEoaQn9yCgrjMIi
pjfzBpFu/qt1eO2q7wiqU9w7yI2tvawso9c8KL7PkW0woe4sX0ffeQ1zlZIIamJG
mAeMGPzPRAw76qXdwtWl2LpP0Bhw/LDUhYyNuHDcrTrOIXKoGZIAg/wCI1p0BzkY
CRfctYCcWknXyR/4DaZ/JMYDpldK3/WyEVz2jpx0LSghO6bGubu9R6HlvxFggVRi
OPhJ4vqRoZndC8tKaGlU3XOfQhajcCDUt8OrVmIKr+CzaoIWHB/biBtYKMWRfTSh
tVqncyCmYuOwQhvQsgjTGHM8g+v541ql9MBeoYZtJPBymVRDh1tv09ozmh4MLqzI
hlAXfqeTPCyER5a+OqNBay9IGthj4BG1Vwz4obK+Sn1CRcRM0SmhATyVWdQ4JK0c
zhqw5gfG/BB9gUGBdpwLJNaCNlnbppqFX48+WQjck2iikOIdNhYz1V7UDErFEZqE
eSMntu/rZk5VN+iXCgqMI/ZMVnSJvoYd2aA4G0Bz6R8x1pO6lfkdhvoi6c1OwHen
33DaOxpN9PORrxRLrbIMgslV/IBjtwy8Kuw7mwnL/PpklUxb+k8vh7Os8Xfnk8Lv
RvKFoPhs3fiW4R3byyxgKGhKRpIfAflR0WSqL01DQOk4NVi/jbX32pTV+91GEDD+
4JnjSMJOwOnK9Q9sl/k+yl7cAUSJl6d7XfSn/jq8b69PtvHE2HJgccuzAfwfhZb8
RsxCie2k9amXffSBNoqDgu8J+ce+aQ8gk8SQGdzbw8WLrLnYequl3SEuvfZE2Xh8
kB9eN+kOUwzO183Vdd1IIOd9hKgfpRXn+hY/YuWJV8ETe+xdwBaZreBV28lWyh12
KMFX8j/UtFSHeCsh1kOffX/ViiueRO97S/3H0+Kuc8sIVydsaoC0ZfEkw9NpmwKA
xfP7VkV5PIOg+1fGr5IM0F200oczbeBs7HPsSFVJZo3t5gBW9FQgUYGNsjBR7Vy1
RRdykXqP18pHpq3pdM/6NzKxRu6qDUAbLlxOFx8b60wvDu2IYZyWrl3QHKqBPrhq
wxOs9HTyD3rfnhc8TuUKuyD3H7VIn5L5mNWm7QDt6i9uUx9PI9CMUaaZZiskKxge
8Ys4vMwnogYv+h+jv0z271Q9STNs4EmfVARrI5j/RuS2PmeSOyz2tphSjhIKhREr
7XgDaT2iXUufQ9QduG3YNL2Fjs0noJI2C0fgoQC+9dVb/I9VarXT0OaP0Ur4uVQJ
r7OkfepOF4T/muBwIMMoN6hkEib2azMoeW8DWI6Qm97B0U7S8isE1vKttT8erzBe
ftgDhcluIHnFe/1mIlwNPwvheKm1a//wKxLFNAujnHklWmKznE5P0G+QPHPvF8RB
fYJA9NWIpO1LrlG7QgL0R4O7ZCMPhpk/PWkakmfNDqStIkcllOPX5lYpgtZGPRut
se0acgVD6EzZb1l5feRRlXd8uTJBvD5Nyaw+hmZrt8ZCFWiXWdP9cXjUmEiEd+8c
1OgsqkJ5/MoatFF6CUhR5wejGH4nazo4C3cFw2klTNTRPl4/Y9m/Xlt7QOkI2Syl
ldfGCcvviiWx/RBwU/C4f3GKuomgqrnoY4r3+mpijs41vNEFnQBjSPKjRofAYBS2
LdnhGHmUZabZtttOI9QECBpp//8L34UcbXtER7FoJbrKeX+/fEYXpJEqpWx6wfOl
xb2EU/xqsciyexwG0iCci/kWN1nSDx8JjsKLzFYmFwCCQOhmuW1uSegxvDt7q61S
1+WGURao/iIsjVnjzvGnmT5dRW+pP2QgUXaJsl2uPyNUi9j8kWILX00fQYdNScST
coQ2X1jOKl5/MDH3QwUDwT2gNo3KOklQulOoUe/uelwj9g8PIdNHJyKv1yHu5br9
omEOjguGDVjCE3FPrL+nnHAB+wXR0c0a+hbpl27KDxQr+9o0wdWJhIkPgk+R1FlR
g0EAev5odulXOKxOA7WXhPLSQ31jhqlT1ajSXCLwT9KGVQYyxLI0C82VVbwa/0Kb
ZtUjOdK7had/EaOd7BkdpO7/GLg3vJ4FqdKvIsjD59la7sg4wkLLFLOUazINo6d2
iPaCOlfa+HIthWuXfgAJFJrEjdzIk+Stmw+nWo5XpvbUeT3B2I42dEs6BD4XrfN4
9QGA9djqXNfHzatGqSX5/lF1ui/xtz4FLT/skSqBcte46aW+dWDRZPmJAdfa6a/h
necxbVEzl8/2s1wxDDRlgi0dqsUyXJ4TC7+oosi4whMLhWCSHXy/TTa6iTUFedNR
eMfa/YCg3rzb8fXVPWbk5HKP/v4GhYiTM5IGPJ2OcULg8nTUIGigYiWKpLiqM0so
eNyCDc1/HPuXc5lyEBlN9fvv/WdoScjcxOrDyWxtlXxSD6gBqLgF0Hulcq/ZEYBI
Ocs4fv6a8LzNJ4e9YjMPRKARnTaHDz5iGwVM4xkmGN4QafkRs93kv2FZjjq+gL+S
z9sttXkh98NK2jLaTGL2dTGYGgCJDbzVqxKBfNuR9/+chGtnDyxXRBQ59GHLYOOU
6MD/rJh2KJdamsBAE+z3D+1FXnpADObd1uzkZbsJwREt0QghL+K5dZXuR7YVm6q7
FD1E89ruGfzvPDFoQ+gAqk1KK1gJdPHxRpn3gXmGEY1BIPhhwyyamMSE7ZQH25C0
vZa8BbdHXBzWGJjK1sfsiPUxWa4InXZfDfpwJ5s8JXEUSo8qQJp9HcGQxR6KWyUo
elFBqeQLhnFvMdmfBIKpXAlgTVSKX50EdssNpLeEfRZZ/3/iTIU6vNcLEvh2bPNY
wClExZj9/e52Wit7fxK9dzcEOHE7hU/fArMhNxt/1j+69QB5/rcZtrK+RpxewPen
4Y8mkZ5Wurwma9UT7EA5JeV85BlQq9CmwaoPmydinChkbCqrmNAdIQSIBWMi41VT
/VI9Z71jIL1J5HbUkNVIKf/qp0eb4OkhjIQ/0IMQKM75rWQm7Q+UWZp83dVrIr8g
jlMuh8HJjrl8bViHbGyD4mTv0DUSWy9zDT00BkOX2rVgW7jBsBvkUirCQpNRSZth
xtr7i4mCMAcvsDyvTdVdq/14UpcnN5R3731VzWnnRlDVD0oj+RywZ4LgVoo+Vrbq
fCJCqUrnWPRnbKCo3406rbAkvCDIkfSEV2UfaCE063xd5iP7yabVCAZPYotYjA1W
U8GmCJ2dsTGv5AHUh2OUNoSJDERzHIy7e+XiAzzr+DOmd35z95bBDVYU3T4uBcot
FuBxx5RZPnrndXK+zCcyUKDqaKkFW1TWVpFXFBbFrxNwSp2yiR05doCbcmmoJoTy
Y1R5TPc7zj+9uKHf0/3rsK7OyI9Df5yfn/2ucUORJA4yJZshii+M42kN6Rwq0/qA
iLIKeDA8IieWGekDbbLTVrx5caJRDQYdT34jC5wj44GzGr32lOebJwiMeQF/pU3P
ImD3+J1dHPi4Yjr05fWFq4Fqa4lrXB9OdQ+lSyqqcBvn/1KsEfdcJBbX3ry/5f6K
XNYCd8sc7c4tIU4jyFSMu7SYeOvTCo14TVn5kjxuc3Jl7rxEU8byY7kLf9Wy0707
4R8MkelkQ78Kmi3YmvVjKQZrZu4YTdKc3bGzUl1MFQJhtm7ZbqUsG5C6muyu0Z+R
aRKm20OsPhxAyFJ2UhhxNQbe84irjKYAUQsLVm+EmBUi7rDF4+6SEyPCahNNiu6D
xLQds6bVkWQ/+pJIZCJQJGIHfHoyhPNKzlwyyLaBjz0CE4tD+ZQzP57vGNw/fIs8
gSHCiCcuB01pW95NyGDjLe3LTXhfJQSahsflb7i/y8vnU/sKLOWKpAVo9Thy4zSw
18AvmdtiOBSUDs57KtRvU8HGvUfmaoMU/0yASciMTINNssD8mlW/MB5CdhdC5o8q
4ARDrj8w3G7J/8RMDmFP58LG/uCD5oRavnW1hpT7Gx10rwYWClzPqNVSX6KkkzoT
iYsp/1V7RmYUHWMkk4SRfpR8yMSrTyrLNb0wG2DPzMP6lfQvzYgipCkEV/ewevc3
AT+5wwrIrOYJrIv1md6GyHOo7J2Y/rye3H7fv3xWYgQ5Oev4vw4mUO/dqE0Yog8w
3S5yn+uKM5APAE/KbKb1Z8413I1GgCN2MVh7UKUCQVegSuUz3JPCR7EKjECfUUQZ
Lj2IOGj2cjT4i3eG6eqIrJA83D+Dqfx3HZcAXINYXvgx8na0vsq78qbfsA8g2CNu
XG+Kb7hzU/M4I4sC1oLxmNgNMYGOq5de65fMt1g6kSDIQvU5N9ybvlnUopZMNOH9
9W0aMVLpiWnjQiQnd2XzgDKaNdmPK9DdAjE+Wu/l17qgZG+UyLIFr/dAWbWym0Ru
Qjbs/GsowSU8kXKyRBdDlNBtMo+pwJg/oFcyOblmLn3dy2T4naX5TUrP2MMh+/uC
4a3uVjYj9Fgnere4+QTbUuuCcghulSBv+YD19c4m/4pR4MA7k5o7nZATb2dZcZv9
zDnvVHi2KymPSn92oApJa0DHq1SMlCOf27e9roCXd3t1dgiXnd3UdjsHcU7Tovfr
+iXEisPxJv/PWfBTP4yzA/MZxBlo3T0+kPvcIELKqXdxXhf2Zc6E8ijzsRdchPjG
xr8uyS1mOzaT4PWVrMMQcVQjCnus4FkmOZR8EpXgteJdwH95Ort2OrczrG6vN2ND
afmTh7VzAq2TjGgYq3SxOyB7yHYtwcin/UHZYiPoJcPdOD6n6GteGsZRxKD4BX1i
/hKw/CKpqohXzKOS/o3xSjs/uDIMyTjHIyGmDgp6exsWGFFjOY9OYypfhFwaLR2m
OGSsQrTGVoBPe2TacVmpSRfMZdGcu1qvoTxGlcs+Z+ccEG6z2FiPNu+fN7Kryn0M
znrZkvziiD9Hq1TRFtkHkmHTjrWMKu5MYvOF1wHUWu7eOb54xZWk+LuXkC7VhNgz
9W88/URXjsffIsB82gP4KXWwWeV04a5Ky9Z1tbWpJAv5J+F+Yh6lyALERueMeOlu
iUvkB93zTVQUFpfkrMaVjDkvV/Hbw7TTiR2zpxnei1AGdgv/RnfREa1OwsQKavuT
DDonRUHyOZlY/22qJLW+tfWtzDFqm1OXYCUWRQBcx/xdHnsueZu6qIOs+RgYRIKw
rnCGTmGPS5/TuwHCJSiA3ZKOqkx+46nTIBMNd2t9VH75Taj8t0cnG9eBhHkuJEnE
DKT8ShA6sf/X0dXotgO19tLfwpNDumwLjnabvsqK+EMFwMtBU0fyLaLDsqDF9D9L
1BLsS4cP/RJnrLpZSO29c5RjsQ/Jk9WB8TMo8JbPxxNWplKKS/LQf2ldpJO9Bug6
j1HtpJdxrhJTZ35Qgv0p0GnKoTFgbSjlNn3GgJ8lp+XglfpUngL0ntgcLe1s9MCl
RQfNfVsIRe9//pAW6faQ19PUlZquQRPRpvX5YxOg2N/Vi2HPT4+fMr0T8K5euFv3
aCOgPLMY7JTTHUVs67uxcSAoLdqFwHgEfxJ4Hg+vrtVgJ/1AtI8nwVKoP5JG1wld
y3f63ptJSGZw+VnrxKjefR0SIdFB+anApMgKXaxZTVMR/2xdaqngCWNYhM+pUdnu
57he+GI7Sq4lOfnuddaZtmbBPRfgB1D7pOEQNh+CX12v5KW9cRPrwZTm7mF67tty
6wo/+CjftgB6Q4WvfJWpClmutQOn+zBFAH+oLTG/mPL1i2djyrjq5BJ6fRhA0Cbp
bl6/Wd1/x2/cOayy1GrevAzbdsHbbpBIt4/xQIFYh0ApagOuK4DsV69I+IaoiDbp
YZdsMt6nQGvz/KIi553mnTsqqVarRqHujNBWz8Tk9+ntIJNpZr2P8gwYOzy66U5L
Orpx8dxix9S+HDlB2rq0S5udyvuCw/1+XPCaSqscxsQUrPhbDwXThWsfMDmfVoMB
sQ82+D37wakkw5Wjz6/+QVQQEcNYhEC3jySHIDP9Rd98I3SWad/fXt4IRtyfJY1F
oRmEBRG69YrHO9pJWnq/4LY6Ut4TzNwSkUcN+M52IGNe1to08E54JnyMJ/bGnpn7
z7ctCteT8GDdBhJ8JetcCcE09z7vuE+fu9GoeIIMKrtqrsvu7ysPyfKCBZwdYECC
JlHiq8vsJDKLeKP+uFZK8Xe7ykJGVI6VdRzsb065RJznfy7yN5rJZ6yijs14int3
+m0kMmXEVzjQBPly8T56dKSjcNWzh/ncngZrkko2x7fbotbW6KCu51bNfeVpJSMC
f3bBupD4LuHxbxRRcNYYuqkat8IgqyEOxBE4DmnbhssBK9KuEmxprOFVOvLnhuir
fUJkteu6NqtJOQAt/ui9UtKAP+hrbhoAU+jsYi+3js4UHdkLO9d5fmA+Dw68onID
W8S28lJ8Up2SEJkbbbwak5pntCqdDL2hEhOQVxrgftGL9DvMU0HrRjyR92U42KIL
8RbWZMzOWRAa0vuIzMp14y/4WynWr/c9LyTsppVZxBMYEm1spzaZuysOyqUXCvA1
v9DWztmO40LR7iff1UB1xLQ6ZSYKpoHsInKmI0H6G8dAFQ+pxsMe75ea5mVnyfrE
ERVZpSB1GSYZ5zfasHIXvbacM30qz62vlJfYbtPVtpSyKCZuCjDkdnhVoIcGzr6Y
PIUhHvDMZmcFhWDsPuw67kmeLTDq0xM2ICpvKhu5cq6ghduIlnCghfM3/gfUQVY6
iGObOZvdLtHakeopsVt+c8ytxCXq4ahvudPxyCVkLhWsPXBjBP0YqRr4AFANSzA6
I99RC3T2y4erB9Y0YvaFt0Bls5awhFWQ2QX8CvWsOA19rmqLVUUXQStYX6VQNLIb
kE9j0uumRIyJRpMaFk9VTkewDq0u2WzX12oL2EQP3GLj6rALf+rEtoypId/cGR6B
6H1ucBBpocnKp88Jj1enx/1AFeSgd+M9beQEUpFsPI//Jc6aXGt5weCk3uSK/48x
49f4Qm4uEc455YUXLUVmF93PaFWTRHXLrCOyRp8W61W58W6Xwd6ozDSAoWDsMCsx
hpe0ejPznbn2ZgJjEfby8sF8Q1JcH4WSXI1cUWYyW075XlWi7HtRMUee9Iwwoj2A
b8MVDQcVs2RiTS7aiqB2HHLj6b/RaAcrsUfAmiXzSc5MdATy+BwxqP1ropaiRA5b
SbFsu+pQcxeN9KdE/blDdTClBSTfKjfMrX8IgRusyxb96kio2qTG7xOLvYkHHY1C
B50tb+kuBynCUWJL7KImY03esQMlSjbYC9Ue1ca0zfQHrPP8RlEAiuSdUuhSbO1i
PUkeY+nfVhq/+b/c3cvdPL76pjGu6FvuFgzuwuf0gkEDTbcJfwQ8JJiMln4l2HT9
E1GI+Jrg/AkejI3Yz8MUa5LyP/USUbBtbLPjNLL52TfnYWsduPyvC5uIe7I5P79P
NEDNw3UFvx6V47wYaTIEmY+Kg88gekoVsW6N6G94f7re9paCx+qWMNnObM74/KAF
aqI2H2/nK2IY/P/btX1MmUM1bfyUJhMsNTFMtELcbG2ghCQcMdsSfC+vfgxkEYeA
rzLyGESyGRCQ4wWxMgMHtQzsEETI+tI28IpRBWj29sX6rDZByuumo9xXJYvarkv/
LfRiB5li+POzVsZ9MdBNaQIThx5ahjPfgGxn5A7d6QQzz8+5H4E3hVtPlb1ZQ34A
tGLjAR32w/dUPGyNrjlmL/yGTzVYIyLSQe+QP87OIIvqn/t+pzEQRd4vPZaHfrxa
/DGRIxEynXOYjFkxocfhmCkh9qaQp+6rWQPJOMUXIqffsTe0xBDrHRgDbrjRYNuQ
1kDx80/s9vsm9/IOMB+etCpObtX7Pu9AxJeBXXTgSTXo42nSoVV94J9/s9X/wOR6
Q6QSU9eP5gyDJZJ2Q7Q2QtLjvKPWTWeqbdH7S8pp1EDdYvU1HUTA3S0w/r4o7I5Y
11lVM7qrq6TVcK8P2VD/25huItztJzC3fGN3P9qBbduN5a0lftw+kBWb0JIGJ/Xy
uhnFnCbhxqhRmTHqDzgfwe29s2SQ1wJYeCjhTxH3tldXyA2hc2g0QILLE3t4fmXx
QyqkK8A+xcLvl8t0EvHDJ9ozs2vq1fx2nW5G2OKbYlPwn89ppAtZkpu/y07JQ0o9
gA0/c90BVzexNaWDKJE2W+arRzA7heLalFHT1++KFdNzAfJhP1szovuOBei9JRB1
+WuXXSA2R48koO3ka9PuUET1uGlgl9vudJjWCMmDHVL+CQ8em3StH4J51u2jIuMo
8CXmP8FoesSZ0X4DekqFIa5hid6PviFWZrZWgDbaS+pU8N7TbFxgcdNPfWflMfq2
J34IabjhJT6j91ZaeL2epo6dAKwGUPMi8TVcP7VRLBB7RlgzCbxZ94cqVK7+9h4P
wROGopvWJD3wdbTfW+DpaY5xqT8WTzOqt0qbFnzHy1Kgiw/FyVI7Zsrewmg/g7rW
uLGGFsGq2HeGVYKnOTWxBfBM51LfwQJmw0l6nBq1oaku/uT52a9dYRdm7oyk4J6T
JtECM2fiJZz3UFg/8kKu1Q/V36fu/WMugoDm9A/3b+LRBZcXrOiFWu6hgHDzX1tm
0kjdxgr9JeV1aIFoJoqn+OoICVMzKsk0OqHdiAR1UGuMGQLdCRstHF9A/EXZJxIg
d1yaQ28lye61x22FgTLsSOrbPEnghk+xjg3eg734kUTN/cFtoe+qWL78robWA5ga
wCRyhlE8lWyUBHCKR9u17oBO/upgtzJ2BDEoxrsDir6nGfq/napDVdt0vVqP6V2B
+B100xus24mRalvueJz52GpsgfNP/nw9XaBP8U+1yMXytXe7TMbiro+lBiQqxAVl
q3PFUg3idnqPE2DE3SoCbaE3962gZLV/6sf1kV6Fcx6y37qLtu22uGnDB5IAxiwY
eRG2M2IFZkQvG8MfneynBVOMgrLV8yhP5lc/5HnYJ7Lgab/qur0RoTR06lyfPoe/
KXh6cVqU/u47aMTxCsLEkIz45EdAgJOJc1SDysTCSIpqPgNDV9xVKcrZ/FD1PwY+
yF6UHYhXKAiwDxtN7+DGMo1Zn+xZLdylsYAK/S/8DCW8fXcL3p9d1sQTse4WjMe+
FJfd3Yo/y82+Ah1RiNXkiWYxrGh/X8Jjsq0X8uAWxbXKDA065Z6aW1mJAuSinr/q
AZHySO4csm5b7iOfPK7TDjkfObolWl1+9QJMsQGJINGgAi+s66h2Who+hSZEhW7L
hkC/nmKQ2nutFgJesZRuDtsqvAOo0qncA19tT2wXQ6PShRdaiwrL99YQBjBfbcUL
ZpFcxRx6pc9t6FrWjGEKhFslVCgen5qvEG2arsr3/10mxd83EUNLDLopw6G+yWKu
jKRnP4P9K0yYAFCZ1mPaHkWWsrEufU9KZ3mIFTYgYXk4M8vijeqwOzH5eo2byit4
1rkJoAn6kvZxdU8tyxRfRfjuEvZBSqhOCOCb7zKxou8HJ+R+U6l+z2qye6v1QuLv
WVnrclSxNfY8JtCGhUL+37dBlbsEznDfScwetJtSo8cqCWGbbyzG4PemrmOZ9yP/
gK7S2IIbViFqRdolWf9Ztxl6jLFN9T25PcUXOMO/xQWN7EY+wjHwwtUckKX+HTBE
nz2uYAx1lKYvYiBEL2CoZu8BGk4dSN19Kk0Hek1m+0cWKnnkMNiFP3DcwqZ4Yeit
+0cq98CUxgcsBTGcRiMJszOTOGH1qrlhJZjwD4u5ndNy1QijMX0EIFfMY8n7+IdX
d8MJPOMDomqy3sVYTfsotNWORN7u3kvGscPV/HFs4Bl4cAzcqmvcq0ey5IxhLPLP
ALhd/tfDf22W2HLKlFqdL+CAiyeSMjDvW4EBb4vCgP04o7uud4oNH6UWIBq3Y5NY
slBQ2V3vA3/R4z61YNcDqovHLEPVN+iRIRbP+IK3oPda0KCuBJ3esL6DqP2sYIut
6MvRDVHG2E/zZb9uRyCmN7MPBsWR3YgGPAMcQu+tK30rUTvlzf7P3wDI2plN+V+T
cuKSKU5/hfqQNE/ot6sRD3/2ezmMZiBlaBkPt0Ls6+CD/Wpa4l/7KB3pz6Iw6lav
XZqqGg54SnxWSSR4Rx0rWwEHP9cg37gcOlwdYbKmhKKOv+/f4W2jQfhtkv3c3QFt
O1NyRxfDc1/k71oq3AhkYhCBmRxjxn/ar7hmuFu10yzXpgdD2yfW/lbqaIT1bs7K
PP993eeQ7iLVIKcjAA8E7sxNSkajDvTU8ERL10ru8B1VbzaG1OOhrmFfTvwMqQyd
t+jvXeaYIhTU8fmtwZljkTBP/YKhpb00/SFSILFgBjz6QwzCMGGMsgf9s4WmHNmh
8JdChTa5gVugqxSr7uQ/pr2PRL6uXWC2Dfe0pv+H6nZrNDXv6z2GTfly0Z0Czlmi
AQ5z8SM0QUj5VvhaEIqlnMcnVQKtFqfgu8WH2ZXFUYkUBceDPbfmhLR5eMQFo8IW
AsNWtGrHGQ4rflGdRiJNsjfG4iH5Oxd3mcQyvI+sOACq82aRLS0ZMPHxSJDQgNCf
MofUg2Xtrz7PYPCOm6vY5LLj/xnS2/IFuMhypuRmF3w+red36teXknG8FOSjnTEQ
9djAHJvYG4LxhOe6GA0P6q6aJU8Ier2qg+h10N/zMFn6yZ8UZUFxHzCl7mH7feLk
tgm4tong3uSxpjbGe6SY9QjvwdAIWcmN46v367pgo2LXUvkTnLGrcUryRC1i5gdP
ZDGxEay2zO7gyL/6t5QnZet2S1x71wFCw8b90c4PC15wc2gS3/JJ4i9TNefUY7cT
snvY9DviyQzEP8Go63uuZ8xng9Avvfma1PdhY5kIKY8lmhR1grjoAOrgoaOkQvvt
VLNScCy4WmJi3erRwjar6EtH6fKSnfXwUkrIWQnqOYyMPTlO63lyWKdWx+StA5Ii
ynQG5pNstGUfYrH46YrLE5tig7D326e693+BOxRjU6rabA/9TPDiIWm2vfLoFi8s
2o5QZuLFvSPHs3C2ytIYk92U4x8wAxU+yyUxAvpm8PlNdZtf64c7VpJ56S+8aDP9
6/pC/azc+SovyAKCflXjWykKkamz85gGKJ2c61rslde3E0eXxbpL/7hd2jFeJdfe
iSsSleSYS5SZ7PYPd1rkfWsvR7fKyJEsUgXw68rs3ZG8YBHMpWym3R1rRgwUGhx/
sYaEMAJx/p7zA2mrVs/0G2C9GqiQlNgY2L1NDfVS/GKLSLWSIcqQUA0hE7pk0zvi
n0THxVuhj15fffbZW+tBqzeNj2iwKw9ZO9v+gKbrGRVZBZpoxq2yhROWvUPJ7XNz
xxTfVMkqK8YfjiFr24UARghb99eyYzi1LN3+NcaKJbU4iA9P55NxRC8dKvWNopC9
0iglIS1/FsFhonjE6dZilNyVlWYgjEF30iNVRL4QxmL7QGO621yQS20Zxgr9Kndd
UIVnDfOEoGBy0l51qpv3W/JcndcBRKbLJ5zWuKRxtb9IFqxM/njynM2akozIB9tj
JRiAnAVs+tPyBb6ZIHBaYKRUvjjVbfpTtUktgNfisihzKXQBMTGZn0WElaTA3/oG
d3Hpjym8E66u1QwSxEpMc/kGH6oWiREkMd34VCwQnfvt3HkTA9claQsVF/7uP1Nz
wt20NXn/ZTHYKRZWL5SKidHlv3RD608iePqj/oTVuhtKMOEv5G5fdkU9HBoRC/rZ
hfsND05G1NLaM7PubcEOdAhUCqKmZP8S9Qr0YzYB9S9GOMv1pG2gHPwH78OFAolQ
O+tTK65gHUYueR7ihRMMh8d42gP6A+nccxkQwYSB9wqyFCKI0Udxgi1vPvxenoC5
z0AyWSO1MAZ17KWoI75oCmVu6TSdNn5dsP7+uALmLWVXfECJux8LhzvCXeKNf4Ol
9oUSkoohNMuPlrZFrt7ED7Y7JjqdArfVP1MJJGfokS5buGGR3oLdt0ljOJk3TTsU
G704f3EllOWpEsbjpugalUxnIWqv8oEivvGuvVpz4e9YyB8nis9wWrkO4bqH3p1D
QgzQkTE+NjxcEchtoI7tRY5Vlui9yOu4vqCOde4jSNUQUJjEN+CUd81bt/7QTxlo
XxGSWeGGM5HKq8W0tnvuolpQSPJKVydmp8txjQC/oPsd2qV+YaiBtELRhc3E+8rs
mD/peQEBU8mooYfUTI3EfQoVyF/jZ0VgjmTEePrM3NryCY5Al6/N1xL8Rhq50SY8
FruxLsXeaxtNj7NRMM+JMoiKz3cxwEn8eCdnzLC39PXF6g/KV846lz0BJc9ULbaT
YDGObCr5Qva6SjIMLA2DL0KLxoSKngv3jLCmzzNw5+btj+zZPplB8WMd92dZIvgh
LzRTaKmgmvtpAd5+NY8FNiUuO01y9zXBZjfcJ3SRbg9Uj1i1XyBBsKH1m9rtvP+p
QXsluRdReyYQzDOeQ0LDc0MYcSRW/K+R8I+EgKylxML/ZwAe1E+Bh2RkJTokRsNv
sqn1Q17d8epydarWfHjKvZWGFj/KtC/na6jdV1rGpXgEF3yRaIj/sKngZDJ0bSF+
9N9qDvhHxoMukDkOKFghLfA8JjpbebOtG7tcEcJf++D5Xpu5ZtTqTqgB0vqwOynF
gi+NA976B1GoEZRipyUwT85XThf8MwhgZ26oJbkUAVkj4rNigZXid3iqMgo13Kcx
latNOE537zl3fq9dJTtHihsNXAIwcg1Zgs+I1z1drjMPVhEYtCiK29dnxOaOZ5Y4
uhDgtTA1BDJXsdNvKOzK9yZdsKjfTSB1DMBFeHkyWXIlbS2+/4UFvOy0H+SonnJz
b0UQkFCnQWtAY8vcVTOje83GXGGyLKrvNYmUbHVsVKDFPgFgOguH3AgE8DCqM7n9
u3lXeoTbGcfNHzt0jYzcQTJs1mOJqH+FFkBvb8nExqHwniUFTyIAeN76CtTaB6Lf
Z+mCX1sM0VtYEIUVTSH3OnsqzyJX8k9L1DJSX/L2fXmESL+CJWdiM6P1UcTaXw4d
yaI7Gd+hWenC5xOvNozbQCAwGz2V7HI1BTx9g5rQNej41nLnZvOY4HDVdhqBbmpF
Ws+A1IheFE1VK5LNdy2L0PZTpK8UAgT2Rz66OrxPJCpB0E1bZ0tLHZTa+IpdFa/0
e0+Iiy/0KVixuM+2TayMQDsRIUY87RNzRNsIJ0GFTK3KsqNZVDUEBF2Hlpx+Nw2Q
jEkoHL5zIuzuQzUfo2CpSPIwaSg/55iIN0a/1QITZ6Ex8S0/0yC+DootAQc2zqk9
CR1jhIRQ7opjZ5VzQvP0UafZ3YYb2qOzgrrDvVgB48J18JrFalu3sTHTOeRA6iap
/d6l2xZVi8LdCQYb8tIjVLxbvgK0ju857t404M4iiaDLLZclUb1ZxWl4h0n1QwVn
mSQaHFekTM1n0LDCQPnUNLjHzcb32Nulx+QL+FDItBJ9BMduDG3NcvIzOz4ZpTY+
+gbz4hCZUgI3yz7CWu1xrvg/39cIDAzJb3kgWwyzNTA2M6Y6xJx6qky/dHqwnWLu
Lcuhj8+gmzUssjbybtAhslDNLcM8YebCUz2YSZL3+buryxPYCtHXlz6XOeQdKoiI
1SGcdV6oRhl1oXO0x2NrgQNNMFbwJ2By31+k0cxrPknIuyngnDmiQgzQwpCEEbFb
xJbtnpqRNc1N1TaHUPu/m3bBTnVyEacSpLiK397ei4Hp1XDuNs3zfBDpYBeyF0IM
iuB3orAGqKcDIh+uzCNwXFW+gWk3cNwMqYsSwf8Zhg1EzcIzMrAsGJr69ayObLhS
+eu9oIUXEn2shspm8927kSwZLPt90msIxEgByr1AO1OTWQRDNmlG/d0B9FYGOC8U
3vcye+NMmkY2aDaRmYkbMt68hT3JC6uQ47P2HbbKXnRGKAM4Y8ZHCKlQvhZoyXcA
fOm9gA1wLpZcHu+n714dLoE4tS1v5hQKVYtwFJXNyOGtJkmeHQghB9hNxUGDwo+V
K/pScuFw+vc3NTwG7o+Ab7lFM+Wx7NgpFUd0wQ5QMbMz45OfZr6CwGgcyyWa1DB9
ar/3EDZui/GldR9PHjPhhb7LoEnsMxAcViuaeD5okRmHB8Vmu26vLFh60z1r7/pf
C3h2PYfx4/3Cl/qMGjYdp3+af2DfEugpLhufHy8fpZ00Dlz+2zYRltn8p5gVDF6h
RwZ0WogcGGjbU3I9GZXcVHBBnB94fc0Se8cmDWEMO2JwjHtnuHJDrJotkBphf+t5
Wjr7dDP5BayJlyG5kiFz1+L9VXaqyhyNKOOMp66JXj/37iVlMLr+yCz2+836NhtC
1nAej7nNq13owsR3I+mxauWcApwp8RTfWwRqNFxnZudGJyPQ03YKKhQ3duHTUzt2
HdjFfqg9VNvZLRlvMX2FSGtxuELt7peC5hyd2iDEnlkK9YFHlzDWxmgY2bQXBHWK
Rvm1x5Q24d+KTQ7HQ5dmK13eaWx6vIl2M1FWqFq4oBjwHZCsaUAhdwgc8iSdMtve
P+evMbqAtN2QYV7YaFMpGRLrO9hlJl3+UhpjK4lPnvuJCedqXayC3Sx8eZnFp2aW
aPa42vbJqnTRTmrXiU+/dgRIDCVLkzVoAv0uog7nuLOn6ZILximuYNeqPdmTZtky
t4l6adDlLmtO15SX6PsGxjbc12ZAjrV8d9Vp3LUWtIFlM4w4SwwiBrRFlC8MGGv3
9BzeESN+GWHh82ouQQ3DzZoQSDQ21R9UGUpr+i3a00E9WeL3ix/WSgxw/Af+o35X
F34VlFfKx+1ThXF3DORJSQFhsHm0XkAS19iSZPhDogep/QTvVKNWU3EyhOs8RPUv
MkCdET87dNHLJmoLiOaHvBRoFbi7VD0GAN1+RB+W3dNZyNz/oa0/ylqyLbMTYYaF
1Ee0PpaPGXtFxf1TxNKuSfGyld/a7s+An3b2dB5joSHgPqZPMDBaxRs40ELoXeu/
j7bQ2JCyf7DbmPh5BG/fchNJgNKAIxmxx2MMWTT9UDYEmpmiw5zAmyVhj7MnAFzo
zissaZ9bySLu/mb3tVNE8FcFNM+5LGZcmcQ45AiqVwgyX33hm9oOIDnlUAbO0v/i
soeAZxrYVnPy5AUTMVR7x1AJVNTMHo23nw7ntpgf9fECyuRnsix0ihozDVvqCh0j
nrsL5GHkuB1hmpCzdkBDhUamx07C6fQYljUjJcJXC/u7ykwJVoavWo94UULYN+T2
KsOd5GgZdGA5PrwtikFF21C+4dne9zNuQr/AJY2LJCYlWPaN2wLDV/7GBh8Ayo6j
0U1S1dtbAFa6wsP+Mzyl8+IbSkvudRRZJzZj0DCvxhgCLkjSJlkHAfa30Z0n7U/Z
G3XmwgTcnN8JhEADEzhEloiFloMiguMfYCLV9o35Za6mdTaPLGgAcfhsAzfQjb66
o9T0yP/mDVGvQ5v267WLgZkLS8WiRYk8+O3eNtjnGVdSfsxYGiC1yTlhCj7B7SYz
YkXwe7A3eysYIwxg1PV9SYbydUyKUiOjnCBzBtPdSRatdukvgyKoN7AiCqQnSd61
TMhZ71zCIL/FcOQr5FQEL3VbFXWyosGYnpTvVETY96HmusgzL+mnnTH0YTCCXGJM
SHu4IzMFOiLrNXeBhHrohDpA2/eyFowB7Td2sNDEyWMEEvUDozEwtrDLpxtu+RGC
eXvsTY5rBXPFTVsmTP/1d4X7JmpoiR1Ji3NEiDW3m/G9hDap3+kDBFT7yt31znYb
82qyPYQz2fOJZbZxdxi500MJEZMl20pGG4E7Tz4JIYKUG58ER7ekGp5zBD6tQemK
8O1AH20nrOLeeUXST/JPFsZwRagIqmEsUrXlEZexQ9XFrPMVEjXv3a/kI1cW/NPE
DhssfkFaG9m3Fgu0VA9hLAPoVs4gb2sDHFOtz1KVFcyZadQejUThZRXcUR694xBh
UTR5tWFESyDCiTKb8x7/ieZ6SfTixZrN4zgccm8CgixTS9qSDGD8kTwlgcWdHhYb
z+1OuRCESPRxVcQPKToAU2+Ki1CVMuwWP5ssA161dNayhMO2ueHTzSDsnOCEfze8
OtstDw1q1bI7xVmaCyazyQ3LJxcFfwAoRTOVqzZqU8pZ6r9e3cSOvnHqStLNJT2W
24Jf0Gfn3MMJAqMHtXlfEuU6rnUdROID5N3phCk5OLS5H3A7v0lc8SXeolBkxe7k
OJWX3dy7wr/mPPhEHEK1g7AiNRx5aVaa2fhpFbjXq/Lq3zVjdL3LKU+FZHjeSDUU
ogdreUeTHjdF5v4Oduyh8iFCblPm/wvJS1IDrMO8acZHRhSvsTH78rMH7keDe3Zr
UOV2BU0vKx9exmFT7dNGb/eR45YqQDiqb6RHm6pbgwIRnmejuVcorFYhG3F9Qw3b
Okqmml96wmjAr9U6XcV3Tsay+JpM8s37TCbMJ0pvGE8PVcbW1mYXYXN52bg20RPD
e6uV1YM7cv+q0438zcY1aHafKi41tl9R7lBQ/AATHebzIi4TAeXgU/NPyh1dv06i
ArSbOkW3f04dvcb1nWM31v3x5kMHpQh96PbBbuSnai6Y6dAnMHfztTeIw6RDAiRh
+CbCOkg2mhtmgmpk+ViX1bv/PfoBBGPdaND+fRreWZjzAw7DC8v5rPgLteMVk1hL
db0XW6GdSnDJF69iuLLNCGFOsADQNaV1bfzIYb+OLBLbcFDPxzKvfDJOS23rhxt/
igQUqSdrceX4A6FboI2j34GhlZy3oDXkYOCYjaJdvQsL84RwTofERaMPqUOLtmzJ
OmysmOrRVYDmSMSk3PBLZtVw/41mpHcQMKSbg2GotEUbwmY/mL/+9+NLvbH3sXxI
5ne1fFdEZAk7so49wL44ZY9X75skC4QnhQB2QysfsC/8oXqi5NW5rZC2xhTiV6z0
mN5uUz9GQzI6c6N9fg6r7Z3jTxciCMcrB7wC5SiLgxfb3DI8HydQjFH+flpWdtRj
WHAKKeWoq3N6rR01YMTdPvjEJOHXIzaXQnq4hCe8cK4ejSaHi5WTBdWeEpFVPdFn
F8M3HaAbpukUm+UkNOhUIZEZiamLV37EhscUSz1uk4T+oN2L7BemH0sN78Jo/Xdf
kBNog2WtNbh6x1+rdIfVwK6ljS4G9D836+HqeUs6poxL73k/GDVieb1nD4B+gwIU
dXo3J2eto9VfMiej9ed731HEO32gw1LB/YGCnsSbSQlvDm3WEkgWvhnHM80HwRZB
oBrY672VuVAXrf5KWglnVxpGdCJSEpyfM/O7ljrarQMKHYjZ7Ed27uRKfPIod6VI
i6j6dJ7lhfj505f4zQehnPHhIse0mIxxQmW7zI8aMCvYuMbvdjt8kZJGF7qeq2Za
h6sEu5zILrjTLL2sgCeixGdvX7GnnodJaM6L3cPjv9KwmXPpE1Q8QLU4Ngz7kkcq
bTsUZTika66Lgp9+bAjaLfc+cyIAjU2FYWdgJbLiR9PfsPpwHj3Mn6NUJf7cBaXu
aidgx5M7KDm/eDApz+C5wn4am36BEboBL5bPs5viDBVXigkcI8+7BnEidploisX1
ptIx0H7hPn1ddYgjPMROW4ZJ1Kq0VtIA8XOWOsGADZYCixe6Knr94ENrPigDBygs
dCHFQAis8VytKml+DuDwDFMsW4z/OUXvEn+3vnpR9ZKxml/0o2tnojbjq6TxxKa4
yWaEIwTlS4qWI7nRr2wAvESARiQbm3bTNFu4J09qPDTiLVtvCuy4+lHA/Jj4mIgP
dyjEFaq7adOP92EoTwb3a4JoqcvUojAZQhXEbAPFnOU3tkEJ+qte0cPQ3keXMXTM
Ua5LxiFb4GYn+sHu2rUxoyBbtOe9HmY4o89zDJ+5TINeNEx6qWopYHLD19bqNojM
o61ZIZxaEMsJqrlHQ9Y5DBSgWeO6IK8aqNMLpS6FNMV/63CgfpBMvGxQ8+iWnCai
LTJzGi4KyT7OxrrxqqtEpPTgTXxWzzWeDjHWyJRU3I2eugTxKmapnShaDd9atUUz
5gilbgEQI+1vmfHdiMUnHC+1H0EomAxS+qAmEBBEbKZZeglBfi80N+P1mIaNpUqb
hX0vsdTz2O55+/jSAKOkUGD95WywqRcSXpu0vKGt5a26/mgiDnX2TeomtGWIVI1T
JGySFyfoWjO1eFRWPSrkfurbhqQWoTFCb8oORkkjt9vahiUVSr+LzhOhpPpnlOYZ
F7X8/8uc7Ik7HS8iiqVutKVn3SF6pLWcLXShoYdFb6PDimG5rjMi7pcbm8r45zHp
1xG3mPIGMNIpWw1Ikip/KWb/DgtCDtVcQsRWipXT/yLXWzspBS1Jy7qkB4A2/f8G
y1qVqrdx6mvJGDLHMmuhsogRrxAcCrCVGxSgYYoQfaOsfWIWJifV3lDuMK5Gn1uD
Fpf6MU0NK9Tt1BMYGZTwJGEx05TlHutH3pJr/TSAMr5zCwFNLRWyTOUhzxL9W1lx
fwIV5J+Irmig3QSb/G/UZhZqV7J3WKaMqBKVhygWKGFlG5dmarKCQEKFU60e4Ukj
Gn+fVLzMKsJK1Ac9uYj1NCujs1xO4t32wSy+g1JIct28EQ0uTtwpCCKX26Ylouht
0qZf7EmCe3f0kDLZf1GWzyEfYLaQFwIyf17B+0B97nltpz6lKWLY6J6eVfGzXfx8
KD9/vtDHkJxuHmj6NBUF3o8EIcHwscy7cQ9Hxq2zo3RZ5B6ShonwI3IIHyRtpNLD
+Yw3Uj6y9Cay90WZIRXzr/lRwzFXabrmkJNaJex9Kp3JfXyT2VRVNIC9zrbEQYHK
mSP5U9PrWlcduytMt1cSYVfkwPJDxDXw/nBAEdFoGlw/Aucfk3YVSawECZpnrNVQ
s5ceNrxF8gun0pKY6tj/PFacoye5rqpvX1mJ8mAL4+/uZS34PmaG0mes4Z+hTEVC
idMZqS6Q0162LnpRJxLJvkFcFTKAITiBhpjpbiFfELakUta0mULHux7JwdJL7Oif
zJfhT+sEaA4MfcX5NWhcimVWesipkrgX3MDuKAK7VbMOjh2qODE4L8hlGQVZX7Sj
s44yFVBJDyMW//MCCdBnvv/h2j7LIHFxznDoZSuK2BslsI0zMU0VhHsyCuoinqQY
X1m+rOdJ+zMue1nQzQghqL5e9F/foz80CaCIoDidGJCSbF2DQ5q6SpnkLiEDyGXw
UJtkfaEJdsksksKo+sX6jsjxuulfgdwPjYFCqOMZc4ZX38xU6vcYMRu7I18+Ztuf
ph7iE7Xx3T15wFUAbyxB0t4h53etbMMaDm/6hX21jq+wx0vnlFlCbt24RY/HxADs
a2RZt9O28kOGJ/eFccOy6CV1aqFEgzMCcAxRxkbrlhvWmFbPrP48L6hTwgCud67h
Sn1dntDjlBCmNt/Pv+YcqpDrDnHQNroEl3XrxuhK54EnJWA2TA/k9VHoIrHo5XHC
mgOVkrjFBgrWWQsWtOdPD/CXpupN8vuYigsR0bEN6xGY6EJNRO3YWPA0QLdCsPsH
sKCohQRWBpAuQbyHdFeIRgPMo0/0rDN4RphCWmYFMu/1Px2DXw3WXQVMcREnJ9d/
1eNSXdRfj3hZq+AV8mwmYWl4cBCvFziyP9iFpb9H1lvXgYHqQIaDodb+q12o0Gkc
EjyQd+WIxAbWXIpoSQLY0Oh/Qj/2Iz/pAnh4NAQVTfGk7z6REkIeX/S2xN/QAcrm
mYtVhXBhzs5bAAGNu2BY52nk5e8gUoYNpBTqAWAoSt7r52j4i1NXvbPv7Qme4Kmx
Jx+KMjYcNcBNEdkonsViJn/uk/1duGpbyrhXdPeWbHK1QvPphRKXO9nXlwbK9bOe
u8xQFNkyNW0ogeMBZPpyVaVBMafmZ/rncNDiJlyLv9VBiSjtSBEVadPkde4qZsq/
hYoxSNpgFKmAmUTj5+b8YqLbIbk6xVkl/kAE+NiJ9i8uNQ91NJwLw7AubpFX6XfK
rRlHpHRIcy1FDsW8BhKN4DkTnl8ggwgnm7wg1c1c0K/wnPcNiJtI8Y3DfaJNcyza
Mtl96YT1wEnR9nKcs1QfwWLVMefC7DuBO9/cMBEsbDB7M+bGeAToLjm7ku7m2LOX
KA7TWE5zjEKOBMI/lAHAE+Gkgg0vE11UKSozz0JDYLxuzQEspwqLIkv1y0YOGEZI
ek042Be4ODrkPrmGRTaYYbOfKW/3BWznMnHlNgGMUHlI5BuOynQU/0MbjdEuN35S
fVTZJS142M1NwSzJFC9ZuC3p8sE/NuBK5ZKf7/NpYiVPEb/gDFq+JId28ih3aJR6
HTuEiNhH+iPWi70au3ZHS/KxU+l0Vv598se49tSyUb0JKIG2syvaj5VCAjyAPVdw
JCH1w4BsiT5+13h1WQ0xlw4DgeGyvd4ZrEi5oSsG6bJAsj2F6rg3002JaGBmmJob
Wg+RsGcE6F7K+JB01nYgtdJMKxaejAFosugnl79uLEzaMasSk6X91026Xb9V4EaN
tb3AFgWlHuwyq2FxYDxJ0SkDI5eGYpeaEwum2khRCes3c9ZQVPBvVdC5bpTPDyKM
oBKnT+2miiphOk8NcaggpluOE1XOg7sjmEEXnALRIQrlZW9mf8BTwOlORPmeix+x
3UvdadtzwKUmp4q3fJxD89pE5xKd+iYfUJR+wNm0ei/0kpvsDhJcyS5O1Ps0FgYJ
53HUpt2ACedjkEmCPa/Vni7C1R0ej1GfG13gPAZ6jVJBWD11W1W37fj/zIIu8Ad5
28DLVx3v71VMVM1ntHLacHQOImFiol32vnxqr3UhA0/omM5B0DRvIJPuXpqpR9c3
qyOaUwpZc2CrNPT63d0cUWdFNDxG7f/zfJzJr7m4a0Tnf77Sn8zAfnzIchOHzZWE
Q12sk1ef8wWGAvSWlnEJOBj6PLurNggW1Y3ft6x/V3bnrENGW9ibhvJ3k2mdfZoe
AN6z6uOKyvX07PjPOXEdtYvN3b0dF7d/OtUtNfH7c5yolVuUdAVVzDpse7EclwgR
oOTkKdv4sBcozCnX31OkSvX6Ih/szNcKJwSLH52bWomBKUwsEHZKyV9JJrwxq7Ms
VB6NRcVbjYuyG3Z97ZO/Z6alG9LOPcgezKg86zKJ2JZu/oeHx9NneCCGboxxY4Es
mYFhYUmFrlHA3feuMJUHj20GkND8XPeYB8J8vMygZsAzpYrekdjBq4EVYO6ZGDJW
Bykm95ObMzUnXOHH8EDnSz4Oo0jfL+Qz0zeyHpmUFqMScPNrz1jQF549hvWBazCu
/NfVw/UZqle7iVPFWxYmdHHBLdzdWo2uHzshPeSchSdXDN7HTjPq+Rx64pOuETXa
opZhxDuWBu33Exj57rb60XlGu9ylmL/Bz8UXibvdvRozr2yy+Hkc1LMN9XEtvbOt
Z0oeVYLwQVwkj3W/aaMTJHt6DPQkMBsld3hwkFN1hMHh2mT7jZB2nl1vacaxv3GC
umCK06A8RnkNt6QodJrxYUrKw70jvzma3Lo7yvCHqLyvles4hOgtDQ7bFz5PGJxp
QXGfZRBo37J33AwUz9oVCK6FgHnZqKOHNbBMQ9wHRSsxSaPYH9vvtrfaVNpirga3
herKVXXnZJoLeMISxM0zZoU2zIrCuCj6KYRlkRjyH7IRqwGeNR/z1/+VD9owKHBc
pHfG11QNR89gS4FhObLNuKSsvS1VSvzJz5cV76y7OSGyVdb/TL28fFSsX8i0tZT2
FbEvv2wiSjbkV8gnelNMWoTTaLj7ya2+qoIIf3744AaomgGdDco48XVRKS0/8Rdt
uBwDg2YoHyk75o//iKTnbNUtI4O6b+b//xGMCBwv0wdJgU4DVGeino9OcJFWqccy
vRyYgPd/FDWMT+GNx8ZU6IgUd16TAiDzlZBw88Gki82TPNydnItQwYwxNp1dQXuk
ouvKXrserWqtUjC7NYBJBYmVVWG3u+/u91ila7Den2RLsD1eh4nMAn9wBSdVvP0C
R2r+oE9hPbIa/psuw/MLq9b+napNzrNZL32s3+08rSJp39MfP7XJ+QTQEap+ibw4
W0R+XgeUdu27xy10bh836xQQ531pFNDaVPVh4uoHy+O5f6ljCsmkkDpq1qoa02uj
a3apYUPFsP2EEjaX3RbkTgbrEcTbccociVkaw5RIxIkqP9+NLR9dj6B0UPTl+F88
nMj9vy3GZwZQwnj+gplZElisfaooQEJxgD+in2mn/9piUVRRh/rzd6jG0xJQV7WW
b3365riA8SxOmU1m7ruvVPw1wm1OKIJq7zA1AqfEZZ90ZPko0meqKdJzW4HvzR6n
jM7P6KDt0TGfKrpArisNv8TGiPOWnTydIB0WLDiV+tl5KC0/s+wVxymKiKeCpu46
J/labt1++kYtifClQVirmluarlH5f/apHukr35BfD1Kn1UXjC8/REEqMq6Cq5Gmr
nWc1SXiy6twHRR3bUieot2w+j8fd2hUY3aiVr4pv0163n46Ykh/tZSBpBBObSzK6
fh6MDT1mgTYX9bkM/2UiETJhmf2a7fSWxhlrPPCbP/4qBpz+3JZW1SMeWBO5rOvN
wc01JFfMEQlQ+/eBDPvZpCndgH56XEsEfFPTjInFWGCGuQXWzb7rt0n+hyh3pN3D
y9LCUnzV7of5fiZFNkjjtap3LVyKUJcag+Ft4PqM3Ugo0qj2E4lsNB00LcvmDoa+
9+g6rXoOle+2UXduWlA/tcdnNM1leWjgq1WpYaNZ3FpaCZ5PRBU5e/Ng47ucqYbr
Qyi9ierA+Rry0fPgFdvjAV0Ocdr7km4IDYknIMrTofaPlF9fqnfwqfYTVeOoK+vt
v/+toNL2raSm7STZwXJZpp5MwYdUxzm3cqdAsXdmOSn48pByOH/2OdxjlkKW+4MV
y2+DLXXbYrEKdSWCngpkOzMfOGQD79H7mOl8cXFCRpt8hB3orCdj9e3MChhQt9hs
ZixJ9lLPegcfseu9KrvqKa4SJp4HdR/iUyc8RoASQxKqKchYTWZf4Hp8S/DdjC/w
/RK4WK2EvXb7ZKXuHkvNGftFh2usctS+/lGrITJoshImffZXof22vBETjyOM4RTm
jFOSH+52zjnZKESonudJiHsAQWDwXEbB7RPoatj4cU3uMPoIdsFBn9Soz/hWZwFr
YDQ/jOWL6zkz1NAvpX4b7PbHfzHG/2PJ4IbFIVuPeMg4iVlcLm2S9yyc1CSy+XMJ
JDi1FIoaY7AyuJ5GyyIu78pNZqjLG8dxCG+lsgkK6BdO82aq0QOpDKlUvc3LWk1B
/JMNhyxUlsNMiQTJQrgFkGS+LZZcij3t0xFjVPRvzixWtCF+wGxtQE3sIG3n1oNQ
1ioKpLSRylp/Wq/7LXWlvIq2AbRUP8pBoz3tJJP/f95GFbRckeA2jdD75RK50MNL
6rAjb0VQ2DGQJCh0dpU/18iwmlUpOcn2HKvK8ytLIZFS57YcEhNx4WjRQJG3as1c
S2iMANOKNZhfxr/cilQLGb8QRMh8ESHvNj/yMrlxlrCrGLDWQupR240apv0sx41t
gyAaJdA2UWqswiisTR+UhKtB4plQVGwRE8GH5MLfJhUx7WOg+6RCzRgQD3MYDurP
DA5vCvFdXMY6nPdpQd4tSKcC1lnPIkWqYS1zkAFs+crR0L5WPir9xNjQ2Dld+js8
G/o7KtGNUVoWZybDVLbk7BTTxzaTufLE+qZctjMtOq3nbJ9REV8lUfPBlvHcYI9t
PJ5n/bXrVw7McNCt7QQpSP1WN8F2AawcB2mHXN8blLPugQSAnaQEMZHV6JnY7MgK
2KLfD6S9kFyOUW3TvYzgbUy/ao+74I0XaqvrCG/E87ZmcZPV1MLdL5oDD7hCqRZp
FmHdVuNefqvftHH/tYCf9eBsgyXEv/K1lzP13ppa/qwbt8zIe9ndOdJmagJc1j4S
5oHjLlZF8Y4nilgQY+zUTP70SHPbAoMyS8yPkXABYD/f7tLZ0fC1PYpToFBPKFXF
OlI7rDwNF+pMRT3+yenPenFZQrMj/SS9Y9bhwhyiFa/w/IBw4qC21lySuG2CiS+q
voHaaoJUtPi6Mo7QAWftiuEluGbonPcWv7EZxaZlUzWjHy7a8Z28/JhKowUeD/CB
SMU+2fNtUhJ8KIdjw4T2RcGzEuX3ZryG9r8u1st+e2gBsT9qiD25xkiy39V0w/Xr
Q4H8XCApDEpKFbKvkAaBJnPR2lsCJKqD0XbR5yFYZ45BE/bovw+7YCavX326szQb
Ei39mgZ6LvM+4B0M+iBMJsJq+I5b0EHfWxsOPUgy7br+VYzOpcOHGiQufq0t33RW
BpZ6SDS5bTxFBOcJLys+UoTpB8KyGu9sVtwz2mPE2/zPumGBmg5tkuqSLGXeEE8+
k52B2OK54KpNIdjUHrtQpXe8/7HXIqpsKbNLL5aO4sELmdRVM2uNir/vfkPBKZ03
+x1a1dnKWrdQ9IblxU06fWZaCZFY9yfdyXl1/PJBWu8Pdehi9xOMx78IDlsMzp2z
7BVMlfn9GfmgD6f/PSJPGghCfk+r5krIHsSUpsVJvdc4d4c8clUgaOBUi/8I8WQq
ol4ix7slhy9Xb/4FvIBlkqhgTCdQc+SlRoIWjQVKf+bTCgqeZLDaTb8845hBXpJK
81QYjaeo7NtT7R3igRGWQJZwB+ZHlddMYS36K9IwY35+ttRUnq4/C2UbWTJok4IB
sBco2ClgdGsNhzhsy8n3yLYRjDSeyhvn3bHZSZn3VAXwxkup6YC58jn0JWESVKDp
tAQcL39T4dOxX69SuXItxtj403P4qPO7HsD4De9hiHSizKjrMUHtYdywAXLavFpI
jOPDHPpkKrCcCUXrNE37mEdxmTcz2zyin4b1YqEj2ygmLuQlER5NLCMo/uMmg61Z
6XT2HydwO3Rp3BTLSFzltxNDjmYcbHs4Z+CuUzH2ncXRqwE+7xoCa39PrBHOn9YX
IYr/54xZsXvh9W4imb0bAsW7ufct9014qLindrIrPr5C6Kuac+/8rE7Vk++LHT3L
gvys+4f3r/ywIahfrsJRD0qRFfHw9ExVj8jdeTQiE5rMLGs/IumjUKVBnz3oA1bH
d+WfHpIoApSD1VOZPPTb5oVCGUEe2qeZn0bkPdGcUiodUQtOtH7yuU6xqpWEPCKH
3idqPakgwFAMXQNpyfRt3n2EUxOwCu0ntCyNjlK+67qe52JUi6aGFh+td7Vp4NZh
VnhCJSsg3HyBvhjCS1ryxwf9SxUJdhdm2A4teP3ElO9CWm7Lq3OJXzbcPhTCcfg3
GxUVuh6MrTQI3vukcZPdvBK2vi50E7I39mF4aRcTB78hl71lsCtlQzETGaYIKAVX
Wp3hJS6HJc7KCsWcMXm1d7/I1xX7ZzWu21gtPwnqZkX9ccoDIw98vCDZES+npeXR
/eQfGm7Kx9lHO8acCDlmOO4STFesKh7k1URX+7rEp0f3U/mUWQDUHWsGjr8/P8yo
G5y+Qn8rucFvNi1lqXFa7ROpf09wCU8IuuuRfmzXwtRRHaG9RKUXuzMMy33OTSf1
AizYSucwAiORXcrbPckDtlapT57qnJDKn/5uPID5/2l6YZkrhBet53BvVVmKPbJ/
bxll1+NnNR0LZTGGbYaQd5GTPxRB4MSdoEQwt7kR6GRiururfuilWeLFnL7gBvK9
r9atbdHdUZzzLR/GQoaY+UkVUh93SzB/vHht6WBaPpl5JCGAui3qbVHNpnqBFZ2g
+vc7dNLudPEMzGziobSr0t/t9vp1AbOuf0vU0Se5WSUlpkMLgYmqQajQkO8T6k2A
MiMY+yCOaapht9ApkUw5bzSoFRoZIAyAz6LCfME3PWLF8BJb3lHGD2KjU6KeMatl
oOTikAwb7tRI1kykNog1FjulWc0pDDZCaewaPXzrK6AHPUhC27Ac6r8z142yQ5nM
pW0J0ig8Vu3Xx/GFILRHW8Oz+j/GfQIWGMpRrTfRHogRIFM7rG5DQPySsxedAhix
24pu0oq13sbiPoqmhGB7oeQgIeZSPeRUG7aPme0i9PeLhrL57rhqzbhb+PXdfyaE
+kG2+lzj3cvWTjl17fM4LrOmPRbFAJymPTm6mibVwCTKWbQXDNYtJ8f2YPC8Okpi
bTYPSayediRVR0PbeQd/mer4qkO4IN92TAbPRMELWAAnw2l9m+fXBAKumQJXe8ha
frEQiAmEXENcNKduPlCE1kN8oPJ5xR8Qy5SY60Mh7bcE1OgH+HLnwFZVqFsYg1n5
60TLKpsOYQ3sUaEJiIt9Uf8OwTGTilwcAwgajMnX6iDgyLC7MbHzWlGu+NigRIt8
81ZcJaVQN7QKux7dvKIJEIjRGjHSr43xBZxwaqT/f331MNhxohhBEKlA8euKIAWu
QLzPLY2T5LBRbznHL6ASSD1gowPGHYF3qJpwlOfMlWJKdssPQ/V4pRbQohe9uFu5
h/V8VZUeWe77bfDVfkD1CkdwMj5jzPD/peE7yodBrSka0L1MhjAOr3aquO9fp6cc
FtQtF451x8HvS4RkDFKIqYEGG6aIkGsYhcvI51LsldViEEpuMmz/xUeNsBSUQiWw
Z4SUVcEgajAcXzxYQ1TkDTrC8p0Z+WuuEoF5vua6rPlCA0ZB184gwG2NWw3pylj8
xFwU+inN8Mkcjy4y1e6xDv/cFwm7uUgRjbxIbeGVNPDXzkYZt3A4pzJ/Y6lwzYsM
8pqJ2zgeA0SDEPY6fyBh0eaHvxJp91qNjBetLk3AwNkzpHaMbY7F46b4tpB2/tuO
JZWA0FTQuWPeBG2BcdZa8kTEh7uQe9uQB8m4xcsAxyIP4LdND80xoOBHgWxZyUh/
ZKhWjruSerIMT8G07c0QCTROs8FBqD56mzThq608cY/cgu1Gy+TwPtbrqEKAzdwN
1ZX4KemgM570R4TIlUC5eABaXjVdDHWUhlN2PGK9WW2kOwmdvAnOE0iS06Xfpf/4
MpGrJ66EA1A7pydDBVOYdQAS/qIqSB9qJzKuXYDLuV4ZKzYpvlXEj4zSH41bSb4I
9T80Cg9MWFwvmN9r5Yi9vWB/c/R5xEIZl77Xgg5zWzq9TQClwptnXVExEaxSHazE
3ztG7EGI8i5MpQtB+5aEmYH4D8fmdgg2zY8AlPkzBWD34CWpYCf3XsPgbfgGhNUx
dR+gVJFTP8CqhhSG02lmP/k/B+UhSCNfEY6nIRfg5C0rV5/YR4BlnNn5DxWFCxlz
26eTm1F5tmI55mP/fKSWXlh9G6/WdZdFSOCIVA6Pnl7GeuXFZAA9t32bZgWkjBXZ
k0aE8eznToG6F47ofopBWHy3DoyvQfLdXMumuTrkigvwo2hTVuK/DBbcL4xGwyEf
HXVuteToG8Y5YWEAuHjhWzuA5E4cmV2yta+o33P+JLVNpihhjW4da79OLHn11i3K
29aIX4O4fvghZk6SpTxOfti96bzVkdvoIq9w/smoNXj+OX7wC21O1TgmgOOG/UUh
PtdF7cznNYAH/xADRmfsPEiIOgTaVCsYmfL1br1x/SdvLrCMwCoHTpr2ioN2JW1G
LWX60Fe/oiIRRkN5yVFz+PZlBQGV1xSnyZVymwubzztB/Sw33UCoj9yhPw7ew9VJ
751dW1yJM+mrJ2ZkFrG8IMXiPPvcESz7VQkC1jCQf6XiVqj0qRgtbY5SmGIQXH1P
eRoci3LlaIAVXKLPjXBUudzy85i+sc5Iae94Ujfdq6hIBGM82HTFcd/l4/l+rbny
16AUoyyfBZPOVFkDksbZflynv8jcmzjY6h7tH5+zDlEKBHvBeTu0Th0XClOZUvQD
/pQErVuEoz9QBKRW9HCtbMJa743tuahAUYmF4uOfDANx3bcgfavMCzImyXmUX1TP
L9mHdVEsIMWwAyQHhEF/YrZIqiMGil8alIpomFoQBGy0ta490hrxGGOVjT+cznc0
Az7U0HHoZwoZ1P8UgY+UkWq58RvTVEszZMi4u1mF90Jpa7f+UHJUycgKR01eBfnn
rz2vGzskJMfhQ1SX+eDUf+xpdTlhZ9YjP/2+2AN4TwVnsLOcDs79+xSdmj7tb1zU
ZTRKBb6Jx39u1OTgpfgEMurWwJit2gEaQgaTc4VJvHvoSIhFkf9eMvGxbkim8oKk
cZO6JU2+dwPEK04qup+Lhye7zuQ526jG+1jI1Jm1Z1jnRoValgTj7qUInkg5rAZ/
4sBYY4gmdF6tD+/Db5t3sxCdCD3wTVvTAmSC8+EbMbBlLDrBPFqtKLnCRwnh8TAE
RN3zexJxztjNzAxP6IuwB2Qvf7n9y0kUQsW49u0ORemK43WmOuxv4jR3KxwL5xnv
TzHxh+nmkFQfeyl9u0YIHlolKSesqzhJOlkcPfMQ0W3BqPUYMlj2MxOoF3uHx+tg
T+LMi8yKy1y/XsJJhSgF0sCZZHnuL5ItTOApkBm4FAYND4oVg7UBYxsnp0H6xxMv
x+/roy3xUu1BHPOVn+dG7MwB7OvWLNjiLrxQMM+U3JH+5DNxO5lbdMVfxgbXsJZF
IGw3RR/mMMp1TgjKs6dhnc88qcbUqHxxcnjnL1/b+HAEdnipIJxh3XVE/jITdyyk
ppWoHYN9diQtukKwmQB3QRHO3zPI6mlU9BAiJXzDfKgzQnvq00bkauxD2bEvkHFi
ne6PUESfxLFS5kwNMoNQZIoKqB3i2A9ajdZP5A+LPK5FtUK4CJFhsSdaWmbGsdOu
U2EhOMtPvYDaK6CFGKQ3V9YH4vDCuDjfZZwTP3gZgf3Rs7hPjpw0a7ARJZk6aSYH
3L+U3l8jNGDVUJeuMfMXBfL6id5eDhWQZOwWZMrALeBGedjEB+GDxAYZEeqCt5ow
w40/3OeKqDyR2vAQIhFjYzLpG/Nf9AofYjsJU5ZuebMk7Rq7dSkCK95BqqsGAMsr
//pHUSkX0a8x0H+kUcEpBaorLCiWCeYRYFcR91B4mjC9MFRo61c+DczaoQfCIhcj
CN1KPDizb3OpPww5PRqi9CJqyy1Fjz5NcqCNLO4/V+GzUhNoywbH8+g0m0IQFNsz
pxStzby5WKOY89EZhkTPxbQO49Ih/+R4Gz6+zk2YiNcgaQtNVTaX1WQ57ypJY3TP
bPk3kZFtxw5XKxd4qOF/c2VDiwuvgA1SlUtAkXMHItXSuwU1L7BAdqLW/Ypj8GfF
gtXtocuMnSf7E53iOC7a36H3KFnHkthQyH3B0CH1CUKTntdKuf3Rra8pbR6RjOd5
GcacYX6Leu0aPUD8fG4JSwn4OMHAs2x8B8tBLxwLv2tovEvgU/H6dMGHFCt0KIDW
ghVXxLQp5oM47ee+qBgfVvYrcTTvzAB6pwcLncrxvYoEQZm5KGxYBNk8Ujeaj5zG
Xb3yHQj7+pN2hkFl+aSxF6hs4CdXvOA0bngIYjf3serp04srj6AsYJRSopBWZyPQ
wht4D++aw/k9uaLK5LWpUG56iilVTN1EJwlZkDXZYeL1Nf3oTQZIJom5naAZM3BT
HdG+xabOxAoP9YqmR36VrJovVoK246JgvOMffX8o42b97vvgyNqmuj3RtdNymMyh
U8ovswgDABKONs5eARPJoJeGf4JcBUry6UXc7MAN4lmMStH+iY8qP7zHxze1vlsV
oBzY50KQd53A38dKqXhsq8ngZK40TPRZy2/XkPA2SxUIjNQrtvgygNte2yumqVuV
3hDqfRc8Lhtk4MwtVK+mlJQ2thoWY9m4Srn/rkjdTZPowdfvFCzghDaVWulu3gcG
kIgQ+UEU3ZBDGNZVjg0PnaulN/Jl+jDHBKRsAhzZGI+Dfi5eGJlCfk58ctYD/MNj
WoGiTii4mxY+3tr6wc8LlrfONo/luIO+1fXohAdON8PgEe/exGS+vCyQMbbBGlmV
1tuRlTTcOF/RJUkFpyfRxsDzYjEnLvrn9cZQhwraDON07r+hBj0asFst0T5sq5SX
uBogsXw+sbLGghn4UHjEVsTBt1QDKOfd5ZLiLT+LjKBOPU6ZHZMFjU4/PQap9z8G
5bXpv0nJTpazY6/KhW3UyUCb8nj0RbORCtQp07UWCQsM/Vj+0Xo1079Yeq7lf7qm
anTm66iTLKzUeW5q39n/1gCjnJmY3Y9QtjyRbYrt0L8N3rb3yqCol6iKtuHvRaRR
EZV1vw+dTpFVRZ+S8HA9yCQYUZ8N7DFHJTgVvCfSMKqyyALEBkjDNte5c6LOocP1
eaylLqIdj9jcS+y406llHWUMfVJQSeUoUZMb87uM9Yeaokx3Z/Lvust51mMybzhs
7ewh2vfYp4mRrX2Ucy5sOGQyHkQkQ6+qgJBZTUgBEwSY6Xq/MP2pEybLpkO4jxV1
2uTdY77qxjcnU3fpCRFqwGBDlBud27EMfa4Noi4fO3exO484+tnUSRqEYnWYEPvg
Pnj/tZEjhixKEd87KvK3mNvB7DG87BbKl3JvFC0xW41+lSFo2W2hQOanDBuz1hVe
bd6OdtjbbeJk6qzAAnR1YIlLbhaLJLZm+Oe+N9Qesw3sf5rLP7JrboUakyrjqrXG
HEnb+1pxCs4BmNlJtMv9VGT+iTsmYgThmQ+RBc/po/ZTkRDSqJmOf2rIfcnu1zje
wsIVQ3T+Qr2KBmwmmtrCaC6HZJkIX3+j02lBPMTz/UMCGte0OwujqN4KWzVBU1n/
bP0hYWx2BeCH0+1g0z80CeH477+VM1UXZTAMrMGRQXyRCXrOJCvq6cgYNXGKeiBb
ojbjzl2ywl2G0Gmz+dn6mm1Kly6qGIZgjQw59WSSXaB9YX9nWneU6dr/wENqzHAk
PeW76L2JMy82ebOXjZVhkGTaw1GVKHa8Kc1MxXtxoVug5e8pgm6rBmx8o5JFfHoH
wsFsZo3mDtJLr3GLfcaGUWik/ITP44HGHdy0EeA1qnfh8jPyko953Y1FL4T6fa2+
+jx6RxrZN2NCQwrTH6v0c+vYyUn9mMQ23WrrHSDqPqbVv1+EtNbnzf6NXVUKMu/+
+jh8bem7Eafx+og+rbD/zxKO7ozAbFPlKxkYziXeCeDW3kvo7MmIxiy+u6JReZqX
GCadxe535ZJ8IjFL11yzGEwSpfaPntxW1iSMvxfSg4JzSirCj7lgs4jejTny1drW
xC6R8PTFVupy6zd5V0XbueGIu06d99CdVwftglK9s+AIzOqrL7V+cqcx/iwIEBfQ
yHN3tB8ezeXw4YK+1x5A3zXaqk9w7QitvV0RiB+AgWDyJAyNT4GUnG9A1BnnSNB9
WQy+o+X5uep79ksFA5ZU/k01uRmsXV0MpVmoBwHdu9kMroti+OU3e/nhzqHFEHDB
mhIsj8NsEgH76ejmWMJwiOf69NEj9enDW+8uX+Fw34GeIYHMh79rUUJGN0cgxc8K
kCvyv4RTEjQyhAnEE0630w28hMwtmNNgv+zDZxcbKfraAm0bJJDtUwyC6wyA/zc5
xCZWiJw7/jj47DNt2RaYbDD5GHIJ1VKYbXLcn4SU+RzbImyquk/DagPSeW2eg/9p
6HhJ2zcHTBhWc3IH9xGOc7x8hl1MC2QKb4BXV1UWIm6FcMzADdUG4DTZSR9JREWg
gqohUfvkGgb0kRTL9rLAT0i3liqmqt334WC8aJLx3XDHJ7NXbNwrAGw9jIbIzPvG
jVJeCFzlb4JTaStVeBzM7iAqFdYE+ERv3Gq0zLkRFWrTbz2cRN0Clv1XDuP1Rqb9
QC/imrwAZcoyy66zS0p2key7CJSuVgpOcFJ1/XeENuImtkF3dnW+1HOik2K6o+zM
8KBf/MQx6hvgyx+WkX9UsWikBB8bH8EJZep5DtsbheknJ8kg2KSK9IIgtj1GXEcE
AxwtbH1dDrEdizKlAezTwv530tFqTB1bhhZQXgcbFfU6Cw8znmCQvpAWdLyT5Ckm
dx+7yOkhSSyR9ENZHGvFx0tA+Js5xtVx3ev2NUuOm7yGBa6r34oPUlcJ2EJC9Wqk
0yTYbY5S6RcB+c5NPogcBwMRXAe1miD6l8bRskDtIhuW/JCcplEkQdJpYPlUA0eH
ku6hFm+HexJ9Bw1WEBAZA2oGmdirzAvY7TqFfKwpUknMRt8+yadQTqjqwhwEVQW6
gwgqp3iPmSLuUJM4GX5Icz9vQl0RMmc7jBbIsrnPETgICSG3wvHH+gJmiZ6tBOfI
xILyb50l02Imy+h/u0elyxgyMAtBT6D2Sq1zhPiIgyu2VnlIqRhzijWpz/HpZSsT
auS4P/HxyrkOW17JrrEQpdRYVvqgtspz7RPWgkKT3vOUNUp/wGvJHu+4Z3S3K2or
/G1RXRNz8rRvaxJ7nMga809ufnR8dls+DJtPun9/KwjqUyM5urrhWZDzKQe4u3Kq
IdoJ3m592TPT3hrukm9rhloA9zOkq9Ho9HilHPFfbyciiYZ1MJ6DK+06mTJYI5R8
Yvxhm2WFSmqn0/Rj3NkiPVofPXAlfhxrOIeKoKgT+0x1P6S8SD1p9hWkv7HJYCpb
krYuZ7Y7OY+WCuI0lK9R1GJeNk7oi1EXgCjQYX/zTt3+2zYXv4pm0P4vIbJXVZA0
j47oHxN+9A0hjgiR/3/2Lt7oOkdrjcLvINUxXev8NwXyFNQvcol8DDlI8nhNck0U
il+WyB97fHUDYhURYCxA7YIL10VVFuKpPEDYQayfbkub0/QIObGotLbEXRWQFi0t
bWFRCyczZwEoTzA/9S9p8dGIgmOvdYX62YeQ8Y58MfJpL537t35W4LGkgTJNO6gG
Uh4HqiAkEhLydZE3PChfJPZ+uuLj4kNxQnvvzb75XydMx/7Yhux3tHiB4p/Dczlx
CS3CmvzTY2lStPh11eV6r+iYn/kcEpVPPP6zxGAyvFEGW5otrwxJnEyx61sMNiyp
/WvcQcf9L95RoBN6GhpVuPe5gH7Wov+Cl7w8CaZdRCk666Mn/bTsEyESCaK3/mLC
FO8y8cXvXO9XkPzIQjgJJATw8sqy2q/Thy/0FvVQac3Vt/6RGiYl2fx8HftFNn6r
yZhTW9fKMDspnjy9e0BIpvh4ltReTrFKxWlgeXBX2pGEACN5swPBZuxfUzC2l9Wd
burnR57Ai4kDiTf7DfvbCZF5XsEG/Rr+qbXuuJPBrfZ/6zWxUXEJnfK3QHVnDzp9
8h/K4eXm4gQVfZK1APfYHcHqjDQGKc5hJvesh4OKjKvdTLeIk5Hq3kpT8Tv2W4lQ
RSgHEMOymsPp7tuYNZkGwtkA7btiMfq18Vf652tqamdm05mfkNfl36vLF2KakaF0
9/ubUzJORcmcEqvZ2frbjENu935HDh4Y/8gbOMzhYOkJUQ13Byqm0jB/kzhCcHMS
SCKCs/JQ1QQdkH7Qw3PYP38JxwQTWI7Rp0V809HalEC3qG/G6GwjU3829cJ3xnA2
YXgHEjbpp73Wf2h8BRGXeS8jwS+Rfelz0ivmBXJSfEeblWW4fhqlGX4ApcNN9gkO
fbWGqeGWbHLyHkI3jC3wXX2FBo4vyTagBv10rSogpM5SfjhshFBY84CpsiUOhkpN
juorQV2yj7IggkWBEVOfoWFKMkrPtj3gdkp7DVIdHwRpRSG36rL7TvZUgf7NinE0
4/i571tW2qMNOMoVJw7KBErBQqdZ+TTFVmH2A386YxYKXRlBmpA1W+uTXa1Mj5gL
fOLGaveH2Bt4Kfm5oOiXYt0nr2FbzF3gNLE8nNzNIw3toOF8bdXT1R79iZV5nNCd
izPi4YnX3h+XEWBJZK0nOYyNkANQzwtvwsaeoo6Ro8aabcsJbCfbjtN9VpoErMXR
AawUaa9yqh8gG2YI5E5PyVGtaPmMbugChn2tIbAtksGH5vuCSfTwhkFBBjTxlTa0
ltLqCIb6yrXzDa4u4K0l6LkyTRNuJJht7fChBjrpngBuUnT8lfwCKZUuL6MJSgc3
cZ8NA/sRLlsej3/6GzN6K1qL9ueId0sM/kBIEEvhbhxFHMF9I+gfO7TWvoP4u1Rr
v0UUq2EqOrBtoOKBG1D/xzSZs2eJGk4b9vc1jx8eD1gkDxLQaYsANixkSF3nAsX0
9ARZK9hbptAROkdGhRDnToybmY8iN8RUdUojwKPX5ENVv435yzD5vgYk0/LX1QZf
/alw4WnUO+9gim7zo/72+1piMGUCePpASYzzyg6lqhcflnJhrbioUC3p2XE4EU0X
4U4yMeOC2ks9KmczJ6VA9IGyTbwInqD5nkFVKMg+OCYF6i4YzzuCp9Od9r7NJBI6
ZIaiLpWvN6323mfaVkKpnfOVGz/pL7AyGM4ohZNQdQGTWawPJDA+/ffSeE8znC2T
47I7Va+F2JIXJ2+TIc4foBHaR3H2U8FA9937GKO3JB3c3ZTV3d2i4FQssxZcfHNK
ND+NBxzemizfQYV367ZsC+SpdKydgadJpTJONdJXHWcvDiTUEMe+uhJqPWCI6PJE
VlXFuSRXKM/o9Ymuk90YS6WBHviuFACY83S4xN37r83xLHUvZh2K4m569BTozJ7S
sp+djRuY79p3ChPQMnyVAqZ/LrwHHzpv8H+uQQrRYmIZxS7jDgC8cPBc8y6vOciK
0/bsFGIhqmxt3LaH4AkXtWrxEj8BZ2XcTgr/NDswaWcVj5jyWwWKopjOiYsSCx18
Nv0PiN3wkXmSN53V5hdneQ6kJuWIcQNphzScaFKmk/x3CsZybMI34OdB0vSkh3O3
H8a4okBW246zUiMWLBsiwjpnGKHLCwQ5OzDWqPd4aYLgLoUVN0Xtbqf7dOl/htC1
XUyX3ClxHI5U8Cyc3zCglUWiAMnl/rvFS9zciDLMc21uz+2e1Y8g2M1wFsvFLuqM
0jG6JXkfn35FqRHggBSuBHxoyb/dwvQcBZJO7IklV7AinCm0aEx/WMzEPDQGe77A
TZKrj7MvEWomFBq3bRDerbqk1qi5aCYs+sHu8497vafDbMAhCM91hIvXOaPffKQi
s4cVDcxlSuqGc0YpB3YD/WahYNezx32VliMrmR08Ua5Cuwz5dvx+n76o47lO7LDX
3eibiTTr8wQsnkt47qohW58j8rO5fiOc9E9FY/0tH0s18MkdRAoJplVY/lHwmS51
8HyzvVhlUQuxAsHUFJZb8opHOHjlVWzRNxMZhMwofKA4JkHjK605v4pLi+cvXJLn
BawrFNdGfilxS6OZVT/82XZkIXyk4avEeFtKnwQ8sPrTetdiLVEH4BKqQprnWWl0
cn+k13HR87cytIf5dLWrz+s5XWGP7O+5nKOpgKlnCn5PdBCYZBNcr6/V8YcNPOQy
gZABJze0ykCalEqwCj9/8NrpnEwRMXGpPl3/8k+t1iaZu6lfEimsbz8i3dDINeuI
7f8Mi+yWFCAs4qeJZY0Q2Oox8keaCXcA75SHLq44tdUS9LW8C5OBKwvYH9zICMPP
ENY4LHE7qYLz6+6Ydby8T6CtWEPz/Vw2kXDD6JO5einmKuQ237+MiQpQ+GwkP9Hb
yNOlSv9D0xUe5d1VoHIWDS2BCN6GZ5oOYcCJggBW5Z7IDeAswEwFsLFQ3fkjM1Q2
+qpk90ExIxusH4tNREQ6XYX+YaF9gY3eNqkNObEfOtwUSII46NkJYzjc9TNlN/dI
IrM2JiyVu+JnAv98Kf0caHNu1qlI9ixsbTLrsoZKwiXm/58FIcx+0UWMcbiroYE2
CrZunvohymlVplTrBdjeu11t/e+dommde+keJBOpn5fXAqCTuGPlHoR5E+t/EmvL
R5E+mUgYRPTJ8aBGQlekmb+3QzaQcBzGm7gUaDtFnKLr2uTsQOjEqLfdewIe6nVg
kUZcno+O0vFW28K98KBlfwlYPoqZq6tQC/NAfCromz2xZcGD3Rrcf9+9gSFJRtdq
+ltqTIcBozOBSJuekBfT4KNNkHFoqk7xD+QmeRpiB+Mk1Z2Ip/REk4OtzjviJNed
RVc373Bl4o+IFRkahip3uG8oOzA6kFWcbq2RdYo4+ml/FHZ5bwSkL+H4RkPGcqIZ
13KaQ38aWyJptH8c4DQi/gIJlEIpyZLSTP5RMPy1gr+sNfIIWo8sVbiGVNDrfksJ
27lcTwks1mU2HVxmOBkX517yEa4W+FbVqZdwBrlTSBScSsYv5wuTx46N6glL/egI
0teD6eftt6dH1hbBEcfCAcNKsv3lRsoCP9wAECS9FNFemzHuWyIhEIi4Lh+C2o50
7EQahU6ng4tZrlUqAOp38tIicRRjMcCX2fYjkFCKi/2e9yZOhgth65r3TadsY1f4
JTICl0UBKre9incS7TvLhbGSJOF71gbLKwukfujYLkpBxCOSUhQWUJtOjdkHMf64
NmZDvsrjvncgjn0DqO/WfOOzo8q3ookmYs8B10SC5aoZn0fL+NkU9UhK0y6C9qA4
h8ZNowPGb+n85+OhkXP5w6scjF5Zp/OsU+TLaWbEt5+BUmnNWLczeFgdiv/AODMR
t7dDUKIb+elzdCyBRAEIHNgWip7ClKwHgvjjFJPHm7yD+ZLnRDLhLI41UBTyc/eY
Ojjs41TCL7nSrIw/JAt9cYjarXJeqrKUG751IDQ02AV8fPpiKAVpwRWuHvNYk2ZM
wWJO0MYW7PtVMGiL2bnCvCwEkITApxLfM1n7lfw711z2IMKidBmOxUdHwm0hio2U
lAPQjje6Trw0GwOtVCwXQFnh9Xx2IRWd9Vq/Gm+P3K/+o1EKeE8kTCEYz4nUVJBy
4HypUu1HoETxOoHbqSolCp7ikBW+2Qk6uNwokIJmVROICRGHhC5nkPbTSLjUS8Iw
GKdPbJ2K1jdjW1QzIP7+n0OzfpQFjXmiHXW7nclmNw9z67gEPTMRkVjYyeDGCyUr
YwNgZSXRkgqNpAMdycOJbRB4i/fiaqCXzVDsSg7NTn4RR8IbFQU2kZ6of3FTUtqp
GoJCjWwo30OC6FAchqOQ+R0p1bjg3k6AnxTKwN11e9QipY+SlvctlZFWndehlE6v
XPWjB3f0A3+W+TIerMzotfJt+A4Xc3qV+hBPvjPf2hnCQQN1dBVEtkeaAk2CKav1
9m+iLGI8v7HumQYPofSaVPMcYwjYMWLElRSWxfAieMpnVPPDUfdenDz8Da6SB7yo
cPv8GkEbpvaZPYKil/fToiU1P5MSsgdQFlpUX3c8O9gkZMTsmo8NFpBLUJ9xZQjY
0be5ID+gSqI0wBpRKAdUDz6aR8apyxXXkzaSIER/tyvLFcqbKGy1Tes8j+GCRW62
sgeRdrSXHieSRezgpWtYWJpW5tlfABuFx4f5RvVpW2Wjc9fT/VcX7/0xma0CwrVL
u66ddepDJC4pev81COPWoUu8bwIW9YOOstIJpw6rovUGSt2tB9OeIHwbSnufDKh1
hutk7S9wb8gSqXMauM15T6fL5ef2NGYbwenihLpVikOb7Y0Q+J9j0OyvJdSVsPKJ
Y3+qw+5UBTt6gBAK2E2jYYMdssr2ZldRyjzDV3BBUAY1Q7k2gJ/a9ARTH06NS38x
Bh93AuKITwzHAYBUh6G8ob7ahRTrAtrT4M9xOpd3u/JGC2mapkgFdoWOou7SL1ea
EWtexxZ8OzVM/gjy6bI45cLRkMLaO8jxs0jPKYD7ZGX9HQ2EVLHgLlS2d4okNZtN
3c/Clje919KCx5HBxBxZPWki8PF4rppJgdYv94nCeMb70uRcs2lX2d/vCfmvCXoQ
t26Sv/J7oogCR8zbBazKOYXyf68E6tux9gvt0s9diTuG3bnbms+nivsAAtvp2edS
1yOh0TPxs6QumZS6gEB4TWw9wxPEDg2xH7enRPDwNHEQTbB1XIZpB7Py6vqvp8rq
zs9fOB1WrY4vJLfZ6y68rdr3BNAKnQVH4EiDaLUG6+XukXtldihlu4kZFzQNKm46
+ymqYcLEz0NSmxdBe69ncK+DtZEW5Fa9G0iLolyJ9gu3X3g1yPgnVJrsUalCC5Rn
0P5TEbKj4i5BpinCiG7piQGES0WL+23BXKzuUNyk9/8K4GzoqI0cqr0cgYg7Kzrb
GBh6H8TAVbyz1t20ZtbkEV/sQkN5lil+G0N4fspAWiRJ/1q+Ck8BhllDV29AVfo9
+Rt3RDBYcDLXXcwZV1ICBmmiS3/jUydKfX/8aCbOfqfCgLYZVJIXxt3pZmiHYaqK
TQ+KdfeCH/zzrM1fFMxBt/SbJJiPGXs7hqYRmwf2sTO5UVZ+IUGuqOguchkT6j1V
UTqOG2sPU/rKV4zU9MwIQ9EO3st+lbnbYSGHnzDCR/SIOhQTaypXivcSkFnkWMKe
B8GKe1d61L5PE5526s2UW2eIqCpUdaTtLSp0gjLwXbomxcv9OOa3ECOFcKbRgYVc
TcKKQFylBCoG4ntx7BJK424KB053VSoCXU6H8NgCWiYhewd/WQj/XuAFjuqtFjFH
PCz5xHO3RgZc7yC4daI/EUnFWAag8rXfVbrDZdUGbyedLlarIX/e14+QWYvnd3r6
01iIMUGH1+OyHW3WfOCjYDgvnEuL1J2zxO2qgDY38YIJ/oBRl8VKbO1zWfu6ZuXX
+c1veuTrRI2ONRGsG+qZ2pQ16Qi0WVAeew2rtWhD66+inypqcmWGw5iH1sNCmc7k
1S+t9Y2jGTByx6DrhakXdCbj+WnAdF7t9VmS63gPOZowctPdizkdX36numZNYol+
ZhuXeqa8nxL9zvnF6rS3k72zOIl5D65XOMYKmCXT/3QoDkbBzku/ItcuTJxSkVAj
avrIOFV7ANzLDXVN4vUxwa//uLfJbEf94dNHwS2ZCi05pX7TssSaoPOd3eWSJo0D
jAk/no3MxDU/DvBlZ5dzv+KDAjRjB0s+GKxpYbIXperkrcr2I7ZOZlL6CT/NusN6
OUD7ToQnaEH33NLVsmxvvv02o3oLgI2TZdTQJ1rebK56jEW4st7alEQeVyaouMv0
DKNxYSBUdJw2sFygnsm9oYsAMKUqBcGzjv79gOautgDBhTrr161NoA5psbP6XMIh
daIaAgTNk1sBCZEvd74rlY6JQ8tuKG1XKUm4ZWPpNcpw21JZ0rSrb5oaI/bO/zFe
6+hp09YF2WhHmZFMf141AxENRrETUL39q0HncCzS61gKX03R9bZ6y+K42Egyj5g6
1VK5eTnzqI5vRpcbvmDTOKWuTrCWD8b3gNC4d8cUX/jowFpYpqeqXpJa9EVafaMI
SwVUz5ALkNmuzbC8ZcWt4us1qcB9v0aiK7dY2PhtBBBeeDCC2nAhgk5t61MB2QNM
3upTrHLCu21F0M3FJl/yGchUPwrEagX6JnvfEK8jcWVLSBe6UysY22VOcZQSnhfV
hM5g212BpDbLWdhBjOk6sW2mvdV+BUHlG7cjK8NrAGTEORHNjm3yprF4sD0nkjXA
QC1WNDYy7j3emDds96pxEofj8VbnY3NiJNVUmcq6TT9gizFQzO+8SyMKET7WWVPp
4CjI+3SCjNRk1eAszKO6NZTHu3ZdmdtByvO6ZZ1nCKu8dCzux/Oyo1LBXwHPfZlX
bQq8o+kXamD4wjZbA7vDFXhDOR+SO1K1bEkqTw7oNdkq0nHG3B93Dtxaj6kxo31G
fJuwWOD6ZsPgHDpTaAi0uD6mJwTP1cjm7DewIXTP308hVP3mdLioPWkMwnTN9oU0
577P1NO6aI09mzD/fAG4HWCT/ToZWRkjwTKZg8h7a9wP+RpLFcPmZnrL+vmxKBKD
HWPoUb2lE6lr3DW8eeFlPiooUEnXybtbGZWvD+SkAXhAgmHm6y0O1e0JHqLCnrFn
vo8S1yK1myqhqb3BU7V4sasJqvNxCBHnCo4MFNgSZmO4Blrpkhc2k3rmiTpD9Oo6
NmBzCa1GIlCFzie/wyuXBbmGJoe538XaYKssYI5qQ5xt5tTeqDlH2MEyZrrzAR4q
rbPjA7FoNh+UX5Md39OXI6f/3uPNYXXj2kTG1v7BAb1nkpuPOuz+zJ+H5RIqm8WC
rJqZyGftQpM4M7DsfJzuNMwAX25ymgPlvndRoAEdzR1DBq/Z8eQaQA31FxgeA3mB
Gbiju9lvqDygTGous3WO9T5FA5J+x4Mqx0fLmOpUlPmE+kmWverGEWLxl/JbLWyQ
acYhMlPQPN+2TY4CwaDgEwPRCBU7Sg6+gR8Vlj7KRfm/Be33La7ljqj7ZNq0gR/x
2oFMHy+00wOEXUpYl+G/u1VBtlVe1t/8qnMlrh1HiBNDS7dvNFTQQst/CB7JQdPP
V2LcxWatUG02jKWZ0Y+f/JX71vAnXT9TKmPB9wlPjdlI2prfNgoxrTEpyEVzEEBV
CNJanoKSN/TNk68MmGSg9CzdgJWXQZgUeQvs1t5Clmw6Z/xdrPqpMlxjRvxmgKrc
h11FpaPI67y9GKD6asRwbf+l6c7qLWSmY5eQLPs0JFQ3gwUQjnKFhh++3y+H5Gej
0StsuVoX+cOM8lMsTN7pOToR7kZKz3RRVatbieXXJYI8l/MxZZCQEje9sULJBtCw
UFp2p7UhMbTDNKC9/jKlP1GW/QVrhEuANXnBDYFfluKJYGioLwWNMdFooNcJiVWf
zzsnCO++fyLNtxUVmI5hBgaeycWzPk+Ivlyldp4x13DEfffy3EA8wy8jI8raQ4wh
QCJqRQ1/r0eepu/SoJRD3yg/tRJq22NSFLRE1bCDfJ8/1c6rBqOfkveeObzBcx/N
/bCA4aFmVoyZ2OQ3OfJdOBMusIMABXi8lij8f8kaz3DCbw7ReacudHzwk25MliNM
yQLwWQHu6Ye+r8hmN5e1xJMWfDPODahBs6/8sbCjp9XTNAeD9ccrM9dIk4+EBAcO
29orxKySEvmBDX47Mjc09ZYmKXOVeziMNp2Isp9JWopsN93mX4+z206c1jjPRzGb
sI0aE68NWmuNmnB0aJ21ug89AvE2nBm27hwFkPYqoeo3ieUcWHhYayVytGFoVM7C
DU/SZ3ijfju4q2W/bHOvvNHZmezBZGzlZxDz/iQa7AltPF0YD8JmTCglMfAeo8zp
H+ar7A3ONWMf+nsplTDzE61I1vetARSbakoTL1LE2JU2GfqF+VaVWJiim9dNucLU
GfFb1HAsA2ADqXXmzU+wPlxugSJ7MiPzhs3YcyeFfaUx6bMvTORJea/tpP5gReSI
cOJ47gKtTGxi3AH4WzJzdHQ8u8AqNwjml5EAi1Ma+mMvWqsTr9y/oIk02ELRi1ly
/gAP2w6cCpefbSKA9yqy31+GSaN9rehqsxGkRjX4Yl5rM5XGlgS9tZO9v6SUY0+F
k4rbmKBMdIKbq60StBMtn+AaGMaRbDdUI188p4mfA7FIZXBn6I85C6DlrObtbt98
SdXq/FZSUx6J1x/hiPsNiLQtol9R7KKn6g1YB9AYPLvymMs7TxYcptMJ65FlX2id
zcDaDw/oZ7vPzUI7Rzcxtt+TOf8Uvy0TFVLaBo1DjNBBOmAivNpOX0oHMOPrC2DW
uDKjt1V6H8sILmROjylYxq0nCFl28Q7RpmM0cximySd+yjIDYCGdw8obX/FLxzhA
KWjyQsHmiQi8kUhPisC0u5MLH066BFg5IhoQFnwJPVPQbeWgLQe8MGiri/xuvYp7
VMcUf/mmAiqfjtj+0bX080xJC89U9VZabyxEuLrkHdwK36jSZGCN05X5xZ9u7dBz
vjNcURk9rnRCCQu7FtXCkbnA4oKhNIXJxEGKBnxe2IC7Ah2CtfD1GRDCBYncgkKp
IG7IW4DRZy03exPO97FE3n+25MS5uB4hVkLr9+xKr8bRkseytbYaIFsqDr7u8FHK
aAlAiAoOZX7teojwLQktl7bR7IsV959j79v4wW4GXSqu9hwiqO7S26kp4Y8SoLBn
d9XEugn+8/EQ7JVfsc2BW8qTv9tM7MPvikas9T0M664hgR6wcguS4B7HNflhPGvP
z7iyxQEWv8ySNQ5hwcyXfd0JPabovwQLz1o5/QOpg1Uxu73Ejzkpa2RVQMDrdzcJ
thG4Aal7AL8MZey0D0agkU2KcCYjC3Lnm2FnKkojI+egangpV4hDPZhdpVHSb1cw
B/29dgUSqMTYAZqkadkn4sMFs8zbfuLBGCDZ4D9WOhVTvqRuFfvXO1bLZKJuSUWB
F+FPEesMizg192HaGNNSFhN3VjP/ZaDZT2a2SsOhXLD4PWl7MWNnQACvzX2Z2GhS
eC60vn83dK7U33PW77yr7nyp4BcU+wvQDolX8t4U0pI0WvSBoR0uRZWYs+VtYe/C
elm2RgxfhlRntTYlCAEDC9Q6yRWgcXBTEGHyN4t0QPCic91vVeiluTMu5fLDULxq
lFuwr5P75OHmGuiSKtoBAeQX7yhcusOUD2i8H/GImVOIlQ9sgZkw8QAitu14DiKS
8vNjD3Ct5uM/hgTcrbe7hJo+8LYvXe+Ktu1cM2u3mimgb834VPFpegCP1P6epa10
dSEZEeLF9bHxTj4zHn6Mmgztj/ZNGReyYwKHyvtv529jpJRtPEKF6l8zqOANhHRK
dd9L1KMsfZS7fmNXIbjJ0k6RGWUOolS/jhA2oDdCdIllKQ7ulaViO70K5lw5nBX/
gtrEpFZiPJf3yiqtOEuwRr09rN2+a6rYGi0887LKxA6HWz5Vqr4PavcLZb1kQwDm
khTySIUD8PNMtvmpKTF9o2QbUHtYtFUgPE90fCdRp43kenH8OdGDFkktROhE8Vo4
Xjs0kLnIUavSvkLN1rlsgCig/adke3vZiV8Skv74rATb/dhQkLFmcrHxXtmaA0np
4PqXjn7mqKLiikdgI2mINyM6dqkZFWgQ8FZx5G1WAu5wiDRA4AiMisZdN/sNTz63
684i1/v+1owhdxmYAgSeOAV/FTSZWvdvVEiH04wxpBYcIfdteTgEYtPHihSTi76w
cz1rkeijbE0xig0AIp6EqCBFYlqVsdqeDydS4pxi+ywZEayhOZjLdXNqXnxy8qlS
H5O9g50UvsVrLeuyS4uCp3m0+i1XCe4yvzzEm8ESAVmBowXHp7Yxq/+NLwC4Cy8c
Ji5LV1Wn7ieJMItyd1fQymYPRtLLzwbDHucjYgnhdO/z9khHL1Rwiqf5lup6sKxJ
H6+UYayE9xXvxL6xXHLbHKbKZdtyTh3wKLbm1xtHV8Tpvmj0GqH8LV4JTBGWtSxZ
UzMN15jskHCIg35vsX6KP6sAP/mAlQpCxpSsKvsG1Kk/VrXqq2gPOQ6rjowJlKX5
uPK6JX8gHOMycWtYqMx/QkN4impq1Lv/nqAzInA73HOK7dVSGeAr13AAGjdAR3/w
Fe43QQiZcOepVhUIRy079WwfDUDTK/9qPGs3mcMvr1ADfPu2Hw6Jjnci2ePpHsOX
lMDe8TEE6AIIzu9AWYuuijNKFEQlgd7JkEQOFIamewMNeq15ZLKQ6mjcJlG7xMcN
/sjXu8UagrTKmdFdqzvpibWxi/bGI9GqDXFystuMNtxFxRhQBN84oWxxweHq0jGR
dStVfl4WCVJ4vtOAa7oDnSfHMnTKVRhcVZrhXpztHzGPlcvlp8+u/IzdJVysj3Ux
Mbs+9humSix5q0LEvkkxJfeQQGdIwv1goUCqy9gs8qjy0z0bmCtBjP+valptHDlK
BAhsM0/pwmr3vVhyZkhunXgn2GNX+Ynof4OpBJT2a2fYd/nEms5/zkD40g3UCzis
TDUSSwYpTsx3kI7yAAFfe/RZf3YOEZ4Rf3Twm/mjvi7yaxMEVcsb3c3OEEhKTqoo
PcD0JGcZ3UU0/35YatPcalGc+pQxUMbnHIZUieeu+LOIv2VSMEMtgVIhJhMyMonl
Fe/fRw1TCbcEziMvuOZcEISksWMId7pFPx90H7skPbWHCwMKIiJWJhf3AxR/nnvQ
A+suOYfSfChqP3DSj3Y2rnBUcw6G0dNFc2nT7iLfEW0RAaLgzzegU+Sah2NcPeeB
63jyhyOU0RdSnJHH38HyTh7nmkJ4PYLHEBTgJTx+uaZFSgCmtIdWM5G0jJBWS+9J
BGvgaffeDv3cXc3r0/E9HSsqlYu1hZve8sXaG7Xo90a63+f2CrBiDv/t2bxBlOQH
riYD7VDFXU4ECJaIduSUsrP0criZlXCbeZ59rKYp+GLnHEOwo8D8Heh+7HHd/Zim
/Kc6OpftBOPpFPx8LCVD6NFpp/4j6jqMo0vh4YQKQubfv3dzDZDNTwmCYB0kVBxS
a0r3ChnWnFnO1SQ4b9XyAvYLPRaERM2z6qSLESX0vu3mQj7iO/mMKUAogMPT7f3e
a8JxYzKobcAE+MZ6DDPyYKgFZjfzN0FZYBjgt960pjJo9zQA6z6r9dVlyK+XvyPZ
WXdQRj19PKm0JawqpcmwYmeXt6F41j0Z+UlZsBQhwh6GLWHiN9c7AzIPdING35fs
AZXPU7tH0DstNbCsaWiDnbUXVQ7Ra4rGIvv8NL5GJmx4FtHBSXgonC+sQduQCecl
Vc8F46XUfJty7jE19/KEvUQJjKrJ+DGycbyzGwn/54HT+hXHHGAfCtGFmpSmRfiy
fJI3xMbtskOm/BD4zKDC5/rBZFzZL2b1KJ0p+7eck32YBqcZ17b+H8yG5WQto3Qo
NtHhtWFKD0zRMKk0Sj3qOmAxPHlcQwMgOdZKmEb8zMkKcOyLQ/tCGD149qko7NI0
CWrI/44hnNI+EsRjYH7SlADFcb1hEnkhdgUnpXMAsVh5coJTCUzQ1C7cInikPBgu
dmCOJDEPEZizFaSHzd62T8rYoykY2wPJgMIFBbGDF0bcFBHX5n2CUGmQakDZlsC4
7zUm2ydU4qFb9q/HL1LBvgDxZMYiVRxIzZJ2pCPhqgUnd2w3ShTbOnND3ikj2WbS
0JiGHIenZrpNCZsC7SP3X1oM6iiTQ+dnAlKGvzYEGWp5PxRD1IvTKbKyWQwExovA
GiSDR6rzOSm3qY/8gghtkWC4v30euLegvs9QFqgMr3/MvkuV/ay/YWmKiN558y8N
Ncx3sjpAWpwxSVS+7IyWUVv92KNxU9e++O0s3DK7LXM4Pwlc8/PJAX7BPbAo8LbY
uAVnSV691ZyTfObb57RwXIlyhDptdt7KxRD7VTD3uEHhFWGwzEqyMg3JmfRKY9T3
XIPh0x9cyL3zXQos/BBu3Na/eufFJ41PQYJTMIr1b7gMUOzz+tAAR1ZyMSYx4sER
NXio2t+XJ+JLl+vav5vV1mM2Owhld0bsQhH2pBpOIuUNALRstZeqaj23wFE0hdg0
UjiL2cw6VbhdsWGWuZgxrqgJqQ8moG5y7Xo4//zvxAnFhAsg7Tl4dOXVtMEu67hR
z+1NmITIq4WC7BOpffQHOLB4YA7gQo+Bgqxmv1w1cTvY3jjvb6oA+2rJVk67cdmx
rgIv729A/fZW74F3hKEwdtv9uq/gG85zPoxVILxZkQoWxXpnDRfvpgdWHk50bJPa
Fe/43e5Jqk1AE32NMWFxRItYcCDE1b9EJdqA7rKeUpRsJr1SdDfgqUO1VMO48OXY
P4vuyi6Hp1tu3DeZ9zdADOVg2Aaa7A7VMcw//p9YkwPn1EwM8bGoKKFyVrvBqse/
NJNdzkT6/4iAU/J/CTxZoa2Nkp0md9voYxnKsLsS0t31h/ecn15HFHj7I7fn56rD
2VH74JmUNTHVSbv9oTPIgGaukKzdiZEUnR6beN/S1W42SXKks1lAam6GzKb9UMTn
KUuX23ZHN48LMFYdrR5EvrtwHyVsnVV391FGywIGaiggMY/LPi6dqNJD5EbPJ0tw
5BoeJh0xO95NZ3plER9NHAalT9K2nwgsvAemfB8H7ZTCSI81JJMFu//SdXNBWh9d
KczNmnJiSBRu3/Lk4aQ77/l7bu9J+cdMxuskbPiK9QQ0tSIyfvWebpC53VEWp6tL
Ox9H+HcKXJxVWMdXQl6oPhFbw2WZiawtcDKu3It8PGSJxRWgWYMheg1XPcjxS8qb
ebLQ8iIkLTXQERLKI0VB5q9WnwJqK66LSs/ZwgsdiEhJG6RLHjGl3L7m1DQ6gfps
Z2UJiDYUx280QlDjOLopkeqN98g4ohB0YhRioTPs8NT9dfKEw+r14o7SyumqW+Z/
6HqhiH7KJJl+SLThSxNSL1jm+ap6LKdrlI2RJOxEEMITr84+xY7wdoRVFrk/a2lh
J841AsmFb+Nj3Up/OrZCaJv1r0jUXAfc6vjtiy9/lcWQcQD0wrWqMAXK5WzusuER
LP9s4gA8y1MWggTjRFxcs6uObTziTUsiE5BBqV653/gb10IoNKm3en+TAOl8/GZr
gEuC43hKM6S37uOI+RxhjBPnOnLD3nW2BFFurHuVEDBGgU1emR2YbqR1OF9g2yFq
eSM1ew1cZy3xMzKtOJ8iQff78UxcL+wWFbXpTYXztHeGIVXxsd7EnmkbujPAO/Lu
Z6eReyinjGN3BEZiywjgvQaFw5GUrT+Uds4YkH8++v1XQBR/L6IoUfCJlxfILh9Z
Hy0mtAjChGQ7ZR3lYWksikixNj1DSXpeCNdVj1/f9B5sPi0nB5JklLeL1cXp3Fic
9+tJT6lHy18nSqRyuV2Q7rITk3YJod0Oc4U/I/QcA6rAvVRH0Icyb8sJdp5IR/HM
at/R95FhVeFGgr8a1Mk9LX7nKcMD1XkHtp4SlmMDndw2nI5dO10F7uy27yfjHTBp
849WrPN+kP80CEiJs0dJ30EIwhoXvUntdwQqzV1DmiyFaj0EsNA0hsxumYexoDj/
C2xClhuglcfJwoMAwRi9PJ6VvgnEPTa0u2Xfg1iq+tM98MEnKXXyue7VhzKrqaVZ
k3VBpwnKfCPAuNpth+snmXmqEpoxNt9PXp2ljY5HJkV5fcg/6Duy8zZ4GRuRf+px
gphYQYlVqmMjCXKOILYVehEr2ZZ0OFjimWbSg2Oi288bLx7f749DTaG+cmsKGajJ
2S2hRylAnhT+KAuPs/WjU1gliRImhZw/P8Je8syjNodqzPPF76g5wd/Z1dYX3it8
UGUXnPxiIIvdGMBc7cT2k8xHKFRyze6n0I1TSDHDh5JHPZDFKNgI7eaaGBWlv6mj
cdoSe3oFN4WW0SrI1rZ0pb4ZnzaZWtPsP2ogoJmmBWJsuIpOFREg3HXoE5UAHWz3
hr7pPVdrOtqMWMAl7Yzp24FSGV5UAxZFdwIxO3th22892OOJZu39bUuIC762BDnO
8ah+2ClTzF+52/AHix55R0Hv/oio6X2URsRt/a2K7wjNMPcnvRWK52k2ZA76XlpV
W/Qh7RrIt9CdgkpmTaSsoRE6zxUNdQfQ3Gpi6kPNNVgjuo4zQ3qJzvpo/Cuf44Wc
7dboU6jC8O4OmXNIlcedUvoWph/1FilEKMjfFfSECZ2kkq4fpHU6Wz/Mp+3/o7aY
3HPVAOdtc6VGt0+VQ++0EIxoXcUcEO7nadlARw+d/BQG2ElK+dzPQcohZhWkkC9v
/wb0p9oaaUlb/4aEEoVIOcJiUahWasQ3kebMQnP30nWAcD9P+lA5CawPag3iBGcu
rBdtOqXbKIEkS/wJaCmPoW33d3Ra4NQf4SJcXFTXxpjC045j4k/sljfL3k2fpwP0
rFW0vVBZEG4bC1h0mbVbTK/GM0TYrb1hBAeJZJKpPkMieQZpUP9jdvU2K9IV+WFS
b18aAC06Q57UmPdphS47Nwavk5wcJ5bJDBWZkdPUjjPrONSnP+6ULZ3B87YYD3rd
ePfgrlvkvziUM7wD3EMu8gYCOIVabKhl8+yVlkLbStXBCEqLqca9jT+QRW+r8cGk
XyCGmrBGBEh3QmWI3jAzV6Dyfn4C8/ycIktWd19lb8pBjt9jk1ySmFXq8IdEf0Nr
C5Jl1ABCUtklTnQjUGqfqWO+NhS38WZD4czeV3GrOJw4sm886XHy+VGxblhcrOdo
d/Hg7UnE1iz3orMfSS5lOeE9SwUJVkQqBNqz6rL5O0tE26ibUWN6ckVWOr6D8ono
BF0h0FcxTvMBYzzY0ni3z9NplOrYAJ1dTA9n/0eAK3D55C1vG5JHh2v+SaFCOHHh
Vej7i70GUvemlalpFAWXqZSCwlTUeI+BR9NW31yY/zW2nZCaZGURinB5U7fF63tq
hcrhV+D2k7iW4cFpuB051J3a2iBRrFNzJ8Z0B+NtGAU+sQ/Y9Hlr7oD0VbX3IcHg
JBJyKlKDXaGdgaYA844rNFb6NnZVqPcG+3UaBIZ7E3eAV359rsbQvE8j0SQXd9Mf
kB61Mzn/kjQ/GtZnG3k/0ZGQm7AXMn3NGXtkodUP2/8s7sQnMIdKxzM9S84ElzkR
xXiOv4XWtV/jm8Zzb65NBD9mXpLi/FrKPgvDNb+2tinxlrfOOEzxM//2zCBlrDqc
XJ1nFsuI+uIPMaBGPaYot4bgKBlBdlaTaiaozuyd3NOlqSHhD7R0pffZPx1vFLgw
Ioprm3yXsr6maZQN8T1Sph8D+5EbLpL9+iyI7SPstwFOlag8O92inBVwwPl4qFWi
nxE2SsNmcWUZOGjrrVA7y1XvIXkVxZPDG4oyqnXBkjAVEzoC/kxZ/E7i/g+GUIIH
Gi1tu8M1p5k2JYkhQ4iPwxE6fLcWGVeO7Tt4TMbONkdHaTy+mE/EatB0RsuufKz+
QTsMH9fNx9R7PU4wyL4Tf2aIc3VxzjMYl93X/ZP/8Jc/FugO/gIOdgJpYVKufZ5q
wR6kyJZuuMa1ouacuh/9qXPOrn6zu+5J15Ve1T5UOrb0i9iek9CZ7wubd6MH7vKN
WZm7gWh+9mFZsRouJFsQ6kiTyJ3I3aHoxL8ZPqk8BifvSgUH7TLuqSG6YkGrkfHi
yOjfEfH/Co9ZxS54bqB8z/nj5gPXyXWWEk27u7+1w6gbde93wiPbAw2EcX6JZRJZ
+3M4ePnjeA0KasOPmD5z1sTZq0WzqXNcN5Ls9XVvPm+vkFc34iwq4pyLHxdoPonP
dhChxMYWN7wo0tVcfHc4KGKI30ADArVuISPayUyOdlvKiZWlm4g844SKVjIgSs1H
cBzRXT8o7rBGd+pN/wbXIe2oQdz8wN+o8qnDl6lMaBoiRPA5KyU+laGqb+qoQD8O
bTRypEEtXBOtIAEAavLu2BltWIOPJWJmEr+t65XwTqSwdruPvqnZFmYlWeICsuVI
R015g0FibhVKaxmHj7xh5mrLcMrxniTrQUp8P2IOMEd1XRpICi3OakwT3TytmCB5
sibvrK49I+4Oivg7+hmNz9HbBVJfyZX/fKmsmZOyTMpmHn3s8nkaOEdF79Q+64xw
D+jx6SgDOtvUjndKPaXABievVYTrNaTEjz8fLqDEBWAP9cRYdPVdQV1eUJJp3s6t
dKKjPFQdXNPRhicF+FPbrzeNgxvf4iAwnbUtBVnlWtPYnEW3gEffT41BMYijXSjg
u4A+K3CqlRX4Jii2e5hTOL5WGaHYmEZsNbttF9dWTncQDC2BXy+qo3HQ0AvYTFP9
w2BcGIgxASGPOjM5+mCEDJkPWySItdVJXDH4rmXtgHToMZAZC3ERKiZuaoecoNom
EDes4CZDXpJgbXNYWM0+GMVGNHoXqD6ywqtKojQp46e2GYl6pEehhl4/3I0704I1
/qvkYrrHuZD5uJ/4VCxZoEfmp3GYrQpVgQdj9dxx4Hsz/JCsgMiCdPkPb8RDv5HB
+kuEmzxImxEqEhueZIIu6KkwXtzZZ+W/GErVPhVloGP+16BtIN+l8bIx9mf1yRRB
DfF6DoNHNJuCalMTsxqSahbLQS3op40sboTaqoi5HaIaiZl59ifzStEyWEph6QVh
NRnLjdgPiLYRRSpnWLk0B48HXx2hln9tNxnPNfDjBwjAFTHU16r/rpvtXiJcVYDr
ZN/IsRPYFzNXBYVLgExQoZKvQ45jvGW8lz9mRXJZ1ssO+HA65MnPaEiQUETdDEoQ
qAn/1dWXxoweE50cpldQdarVYDbN4fyY9vgUZY1wYaLfqfmppCQ5JGx/EpzjW/5V
K+K1Co62CsJBeP9Gvt4CwrIMpqrA3CGUB4npX/vzKScynPf1VAINLGsIigLd8+4w
Y8vpE9uvhZpM3ld96z7qww6EGO7J6cqdE/zGW26RX9GZ/Gn9PJsaZf5lTIbB2KrY
xpnER9dw48pe9x5K4KYCZdf9Ov5Z3LPIbSaTSU0SN4uqkJmpob8WD4r1PJsO07WT
iLTqN1UFoKCdVcEvQ/Y11XfELhFRN6dkfATyOe3OI9Wnyd9b88t5oPsytpaLs1FS
kTgIInzSTymq9Oz38ISSWunI4Vd2DHVgzH0wz/9bOEZYAhY0O4Qj/uUtP8b0Oq+X
mogj+2VZudk5Tg12IUvCR2Iwsn+RrM0nEuaWBhtekkTLVH7floaNT88dzaRaYM8z
sEKWMykSglbVJ8nhOhqnBTaw1KdDJ8DHKFvFIhfAya5hoX+a3ObDOHWUehYWQE9U
CJjqsxzgA586GfURRzZLnVPZ2dXVCaPCxMMLICF9sKYVH6uaIIjMV30LKQ6skdhe
s8E6nytHvEeZUmI18K6cY6MBQEK5JYoooVRDO2k+j/8ujeQnq5lOABl0q6RruvM+
DOA116EdNnwonxafMuQah1yttSBR34BbhWWn0SvwU9ow6Se5DJngD2qvSbbCeBXl
SkCMt9mFOfsQwjHKBqeCZGNGFb6UMP+h4MBa6Ku8sBWAROdT7uNTzrlNkBok1ob8
IcNWs2WrnXJmGqbM3t0znjudmpKn/AdibL63wiaLrpQaFEpISMyG7XR8jWy/cONo
bKApWauxTm00aT1LehiJ/vgAq+7SiZowvaKiHSbPdbwULgj2YzSJSS0k15Ujt6O1
FWQKzuK2eL7YdMGOCZNkRi1YQYsU9BmvUgw8fvmLkEJNkKsxaRW05TNzjtfWfXXA
lldwCwFN1hDagVLysfaVAQfewnxyoIpDBFKOvDiuxyhZn6fZb5d87AN3W5pFKSER
aMI2Ju7qSLrg4l51OnsLVfszTf33FjEbrxYqMfFl/EDgrkR96t8omYXEqcwiDGR8
5+4CqsGgRKSCgWTvyPG/sw3hua5Pauy46ObLs8QCjSTGShAjXCOkTanEX85v7y/i
CYXvyU18gHhbmpadMJl4tsSY50xLvjUngRZIh6f/BwAuvgIJBjaxkW/bHik5WQWi
N/LW2r3H5CuHKyrp56Uf85+rYjfRZ+ljYXzMU/amxnNIxL2lQSBpPpJkYcwQEifC
bjcP48YguitE+3IyXdRBZ+qdgXLuTDCzL9NrmQy/p21gu9A8zVE0VfTNWkcLkGz8
1dzUqj+ay8bqsg+jj7nyD2XafH2d8P3TOwuq2brt+qe7l7z8r35OhYRLFXOeDW1s
9uJd/vDtuyET1ik1V6F2a0yHbbESqkRzm5cEWg0Uvs36YqWaw449KztWJqv0eV7A
01Nk840EPR72OktkCMgssV6o5h3m5WfMlKKzs8fr0kKtU0W1ZSyb6I9OeHBUV20E
N08rd85cQh5w6iW1BfYWycpFm3gskGCCOl/W/BjsFyhHLN0SS1RMjtZ895SS7GuC
7OJFm+rc3YpHuuXdCOtn/Czt5+g8Uw7NIgwVyoALr0306DAVvoqrL1dN6lhLxymL
sK8ZUzePJSzdzx8464VkjPL2HaIfBWM+pJ697HxOOnDyrqB7EMNW7C+yirWAMva2
7Sv/YAZ6yuTpwcVQPSZLqv3+VdaKvTkQRf3B0RiSbQmAeb975sVn3mOj6mOwjqhI
nfjRiziM9o8jZ8aC4YeacVs7f6T3hcsgVVtUO576PUY47M+x24hxPCK7xIhqtYqP
O3LFLRYcbb9keuAvzW5dW+NV109nMlhJ6CLfpV+R6EWJikXElLp6xAxTWA2bPOMi
Px4RywjVz7hj4BXOJ33myNAt9DW1BbqNzCgR+yTUEt5yEkY7FhVnjZ+eTvGOmiqA
navBKen7DkCB+7sfj8bBUkOF0NFcutazq5GuuADHz0fGNpqUdl02VyCaFAEkDia3
/YGquGoo7WN3LgSgHu/4sfDVG2ZqgOK5jETNDUvnyPRkEW56ns4Br085LZEn+6Lz
n4Ta30BLHkklnyvRaHFxmQ8yYjbbrTz3FR9Y7eYrHTDYspHA0KSMP+YaVvaz6Fs6
BO/Yt9u6s+HXIcyLztv5n8yQeqid/lrXtsUW9RHFiAZQOG9zediUanr4MgZeHt3J
+LuD47N+7ZUN2LXyozUS4UA4W4jZPsa0TMmRkgzTF/B9FpyM1OpsNn7W5hhPhJBW
1ew5a59pthKZoUbI8ux3rPmfrCgU43bL+4WjOjGqAh5UVBhQFhw3S8+dikbB25Cm
PPN2O+9CeXG1aQhECyxPU1bKAgX/iffL24WhfFZCGxbpJqPgkVKlVdskoDdo2ejM
GumooFF7loh+0NoNZDW6g+AGaxllyD06/m7vmVPysY8AzSmJGchl8wh8zOejJmfF
coWdEVcmV7icQMSwFvnQyuZK/JoGEWdTJdU+xlGZQaLhbwSNyYREO/8DELPc0NM6
cyEIrkPhCJn8bMaulRMVot7laRdqhVuu7dPS6s3G+pv5e9iqduzI+o0hi7EcH1Xi
9Iu0Szw0MbZ6Oo/VfK+spv5sapJpyxjCYoNxcxDYX0ujcZPaaeCTiEu0cdhyS/0u
EVQJUDx98NC3ECboIFi2zhYl8gr1Ffvb8ib2JRFl7xsmUIFTs2y+2Q241fkBL4z6
bOAcWovXrZe30TIPRc92DvDJ7BJtxlfQ6CqnWgsInamqnA+mRgm1b8DsGbKrifkm
cdUk+5jtF1d9WeQhbEr8si6XLkZFCaBjdZ4gWV/d7cs7reD2SnsPcq9a7mgQyOJA
ojb+ab8dnp7qJcad94FTWCkzW3AqQP3j3Hott6Kpyzfh06Ps6wuEUzszg3RB7Xhj
juxlcBYZN2KZO8Sji3sT+29pg97+VOhYE6vcD/9vEz13eNl7qvTfPRvGZIeuCCTy
QSVw/y0RbxpE17n/6/TGYItHauf4bkCGFqcZJM8b4XAm6VoIvV8s6fWdUk9OOYFc
bivRw0BLUPgH/Z4OFSrdYt6n53j6YJk/Afql/7KzJ59T6PfBIBo+yClejN59et1f
JPpcSN3dm44+zvurANmpEE9Dv8gm3UE+Jv9ayx3JjBVMbAVOPBH8/lJ20lCsXR+5
/6NpyFba/KVs8e5qk7CE715dSzMEuCxci24wsVNsiyk4xNTNcZwElClByf4CKbGL
GuG6Qng2fpcLdhthzHpWzToJsqHULpzoMBjdaC4x03rGmpLEaGj64ikw/LkuYjaE
XmTahbybK2Gc7BmqFenbamNfUe1DD5pos5QIU8ssxnTD5Z9GldmFGXlMoS2e7Eu+
YWWSkDmJQ4gxueU2fBBPnk+FPaGnFHlvdshZp7TeCoHQONQrtxChaxOADnotptaG
lZ0lI9ryWAnTmhmpeRruXkEoHyTizz7M08c4JylpJjFL+iUvofMY5j14aeK14pJq
8sctjDT/Juh5NdimGWBpjP2jA9HPe36EjyorhIW7JQbW4zzy5LbZd2LsqS3RVtcl
C6RldWdyJRhmVeV71UvgRKPTbzoe0H4GaXDW1sM0lM9g3oQaQSYYeB+UBuIgtdtr
0WeLZZsbMt7KXfas9C3DerKwiW7AWhL0ilPKb6GkmEkujL1aa+IfiqaOlzLkBXeh
R+1y14tqbIm8jPUtAW3QhAMuVP757SQvQ6UxsU/A7YJi6ji3lNQ7JYSBzFnPadB0
R+CoN21+WbRMPstIPZ95z0qTVSxcnuSIEA5mRtx9MLZjxC4KwazfW6l6ZxZgkbC7
MaFs0/qtp1P2LueM4kEOqzdanKhtCp2wdZOiRj/GldINKdJrJ6gQOaCA/vU2c4v8
Oy7n9mlLm0WRIUXwqklT3vpsbkcfccuFs3T1sqCPWDOxTg/9QQtEFqWRV8OWySgy
yXhyd7Srf+fcb26qFcgQjt9tcP6LW+vRq0J1WGV8acM4pJP36Bxy6XN7mCp8MVqZ
Kv1DohI43MNGrxZjie1FSv6JyHRJQ25+BUOE5vd0EpjqqvCDAY2n6vBDfIo8h8Tn
wlYUGNHxKLcpcQO/vwWZNjycpUU3vRTkz9omWDkblm+8oF8NfYMxYZgzyTWFAjcU
lKmo2IeV6wUce6QLogD8dOvfGW+6DKlo7sst5cQGNTm0tG8uB8yFdf6FIEEESDng
gBkPwrUCvkfNDhIGFC0yeY7dPN+b8rX33DdTaQDctkrB0LuGVmuDrZqKEJjSWhCk
mRHo6e7UCg59fOqDdMYXM/QyYzK7PazgoaznuP0sFLSXNR56h41Tkgd/a8F9FnxP
yKUnBqeFfNywWrooWchrjo/gvrzPZ5r+PHxvzk0qzZnzlc5+w4LLTQ0lsAU7PXEg
KVA1QCPTHi1u3V14BZCi2QXvt8qKzD8r9q0pt082/QTPBby51X9qdfdlw++14esW
DfY1X7eUtaPYMgVPUA49nnT4GWFU+dXcVNUeGndElVaRPJ+6QBFvNjmMq25dYm20
CBHYHOwCYrGxhm00C0x+DKT6gMJSqfXosrYwl3bFeeByTSrFEwl7UZEEc71XWbHH
mrADb+6OaN45nf6o+G6uhUVXTLRWab7gBvL8gtrGM+Te8GxkPvuZxL/pIQyw7kYN
QE7qQ5XWHzL6290MucrZO8SWYJlLaM5KbwZJs1JR20pxz3aW+pddKX1UvpXYh9qL
hKzt0Z+R9q6/ntTh2gBMSWuSe/Lgj4ERxZXVN2NUF5v1UB26nxbZU8Oz28GHqLK1
mpH0DNhFkP6x/W9hj7UhNhORO0dxpFDpUW8YL7Zp2l+lkMV1oEyN/sA7fWvBlkuC
g6BVjI9Lls7lShq9cjx8l4MpDxaNJdQUBvK4Gzqktxhq3t07luP695Z0fnJbWU7a
ychatcZOu/HcPC5HewK5XKbcHhTIrujcirawLpqn5nSZiFDJtLT+bpUr3O1G1w97
6xl7mYdQY7I/lKApomfVzo6Hi41C5cwEBk5NlWbRIpD2ry2ivjS4NVkEYcZ1DQKF
5B2yV8z09g0xj3wAo+nPqKv1ESsbV1s32Wcd4Lah2cnRdxnRw9Lm/yBzjxgTBmIA
/8+IZ5P7XOzXf2i3AS1AmiojyU1sPE6VMRqEI1ZTUEPmNwZNk6mWpunAYGBrLTgO
ie2x2GGkAjI4vo/wzgHjwtOkTUGqLuGcj12Unj30XouEI5brOJv3QHem2a+oHoje
T7wZ05e/dnD4BX4mHjElJuPJLFqqUADnQxgIRe+ohGGCQ7U0uyMGw+1awnGRUXyl
rgJ3AjzbRYee4paeRgUABZw2yIqbeudq1V222oT+nhdK7KLo4wgQYAzGJUHiYqXX
PByqD1GZmFpCDYF9HtV4jMpE80XJtLp80v1OtQxEOGyZMUxrT5rtQsktITeB6elF
aYiubG+SWUC6n4oDfXKycAxN7sPoELbM2IFlbyMJFREwhHVtbc1+yJXPejNMc6JO
E6ePTtLktOPdetoGbALoweq3F/q5FoYB4Ynx0gVN46cNJYjmfVYl1BeFEVVFp/LC
NDc9CVIM3GJ1SBGg/qTasKRH5GsmvT/GpbJ0HNGaI5afZrK1PrHDHEPuK0hX56uJ
OqL+bOYsAQdlLjDUAcNw9QmPR0eDN8mNmRIIdFxgPJB3pOpq0lXhBxAK5oR6PNZb
JY7oaPRKgyZQ6i56L9xart92hcOqxZ9tnV0KEy/TIQIWMwOur+0hDI29pgKmDIj2
y52r6z1DC9+D4fhERu4Yj4aE/6Ss6AeEXXJSqjLsR8OuYVtT7cX5ivPK3Eh3lPxT
d6OgikIZF1gKmLhDj9fKkpvYec2uPogDhrVipMkuUJl3w44e0q8IQ7ZGmxYS6oeH
pA2k4DJ7KLP7AnJabTtMBTbNkv6PNqj0Etf29WfkEjpzLZEo/zegibvDDnDufhya
sprOs/QLH+i5Myn49tVBqa/+Ii2dvMsUiQjRC9bWxwxpCRMJdNlZ/IFC5hsmJLdR
yqnZ4zz/nyzMZH1GeURlBRnlb2/4NW/fsjuDXyV9Gzz9gN09OaMTRUTLNQuY+oei
mJgYYBZYcyJK0u3bPmvbZ5XwFLk/ABj9ATMkAuTOaz9k6fNNV/0yzfWCFV9rekIO
kUInk0mDe7f0DDRQmsH4twMRGnQn0DqLZufhntCsauUx1aDkBupmvpA3joLzlkTY
JtA/ys+YC5q+GKeDTtZRq+MqjmfXvsOVoCdQM8AXcXjhHl+zcJhoq0oxufEyYwSw
5TK8+f1h3I6F7vE6N3i3HpmZBsi6DhoVLAMDQ2iq6d1kmgHFq2KNjwobUVy8e9aA
e+EFrm5j6zXE/7oEgzzaTBTxxu/JXgFq/r0v24ozMsnra5Msed49y7PkPe5nmRdI
sR1+MEHqRtV9o0ECROnUS7X9EPqG2HPHxRjayPXumLDYNIyA1hmBzN62iSgElRBV
arNiDKrFjjvfwPGrhEslKNbtXfbHK6FfWGf/JUp6UoG45LuZ+YO5ovMHVT2WTIP9
jTO/4rvYY7A6TjCIarDX0zDiUcVdtLNXWA/cYRW2ECQI7+CFHJs0KlLqwWZRi270
Tpu2b4a5l+4BO6Afh4HNmnt2MPelAsJNmpIqlvsPTytACcp3tj7yZwEbfRX5unLu
aKwobcB+ewP8/gs5H5hb0B++nbaMAor6D75vQLG43dQlfewjdP4FI7l4NXYoCioY
PyNZkiONJUOHOY4LOPy2IQg/R1aQNf4H4l3juoJaLl2PQrZgvM74HUjO3TiCH0dr
lONT5EXF8mwpeWiyiXNzdr0po0Jd+ADQQjFy/vfT9aiyFHrIp8YT8DGd0YWAznsO
DHpAKePjb2U192JtXZJJcgk1lxjGSy7AI2QLA4mfJ5nF3D9X8dZawGhUJU8G2UMG
DlvjDQqy8aqooTsjtM6RYzjLS5LkHG34olMFn2dwTc9rW1nnDoVSCaK/EPoZJ3ag
ojj+h6B9GnSVG4Mm8UsPBchAozT2rXZl/dF6Eor69vXkGRvPy6nGz+srBS801LJn
dYePoKKYb7Aq055jvCI1Dnmg8zIOhQoQh24Pr486uaDNDbwkdahTWezkI6GyFx7J
826EVvG9Uz21Onn39ubG0AhcNec3VC38FI/ahkZzJjOdB4hY3JkQJ/b9oXAslEvN
W3Nh6N6rq8c99pW9Ke4O7uu1TXuy49A4SD712kBXf+LGm7y72h9hQ9O9hxO9kxit
xcZphZU+cuZJ+6tRicV1D7C70ixg8ufvW1QGqGNAcu7ZWUmi8ei+Ca/UalqJ3y2M
S6SzKZzhR1VIgsHuJmX7XE0dZX9wFpXyyaIkmNoHc1+6nOS/POYUFcfus6Vt2Hbg
KOFL0LRhGuRgZKov07dDvdVLpaGexFisP+tkvMMoRbhBSvug9jBz+OMAgmx0Njzq
8iH/HQm8JTLy7Tb5Rt1tM0MSr1HkPXa3J/rtWCvmTfZoFVxYrvaL+m4+S/ppnZ8N
ad7R5JpfI85gYtHIQ3pz6qhqGiu8XB/WWudVsTGgwZab/qCXRgx7L4p7abyVAaF7
XOyf4q54NW4K5YZK6JkcZNEND/8B35h+5UKNy3BCTW1RM5uxbZ/ovLhvHxo8IDdy
dUnjL5vdt04ReNs3XwFIZ7bRajXA8Na9y3+pRUszK/bMdgwrtxP/gHDY+Qh6wqrY
KZ9Q6iikVDSkdDjaUMjiCUAAe+LVzocaT+EdCAXuSgJQyh8KfZu29aLYvYvwt6SV
wTgwHsMdHpbvVUz6dUuaYnnXbxNSPvaRFHjRfO5ZzdWZnXe2aRBvGluuimLO/Iwa
ILLzIdA1DFK4Hr6axgxme8kVrK3MX6MrVUx/EIhCxF3Q8UpCM8nIjSoqBfI8veX1
7z+ZLAv8Or99HfPdlfxRKtIfIKCCwMALSzoEOjgUpoIhmL51ClTUCL2/5aFI8X8m
hyLQHK7NaaRbRMH81bLmmw8981oaJroqU0edaLaFpVyrEDzObj9S0IBqCtLWOjf9
Nib0a0HlqXJ0APguA9q9xNVsO79yz2YuTxzorLa52n3Euv77ZLiPcZUCHkqbv9iI
jN0HdHPNqyVxzuicW3Qd2LYvOV+5LCwJ+CorCxDzZiyV3j4P5QodpHXXaUV8SWVd
6bAtI/sQs6t/TQC1Ts1kZfYMIGXoTI/ItjbUGPjOHwSlPwzYkLiH9HOZPXtil4Ur
wE9MZ4fw2lgYfILCBxF+o6ug98XUfJhrRxiEKxFMgKBHvH5G0acbvWlsDBWa5pix
xM3mXfEv4m2MITIk47+2EslDqTot0HoqkA9rXY0hsgUV4YWQkHfVC7sYmSFmjRee
LvcFzE6FhXg59r0CynhFb/z4vMb6KaFPdxfECg3AUKLSDVUiZp1CCwxEm+jz4l8j
W3cAIS8TnoWx0lHjdaf03Nge59ISlIIikMCtNNLlfnM332uJALQJEv5jni3454rP
RWHFkiAiMdSAF83U+zw7SL5rlLzbzNfoDtzXW4+Nin5RLVkj9R2pG9i6KsrO2RUA
LmaBZlcvpVzmofHvSOiimivoNx7Jt8dzC3aDCEKV1PJ59PpiftbD0n/vL2fAkWsq
wRXQRtLsg+y3lR2REwk0KILRlnUo8Rkc2V0hcGHtGBEmBP7sXeO0H2ljtR7RdBkV
wh2mHza65434Y6qqtIEpufzCzsQ6sJZhBGamZSdfBrWZTTWARXBTEBwdKdbHv+aK
JRueyolYzM2SEu5RjaR7UJ6z9oj3pHSIjj0HJ6E4tIKjU+6vQl3QW6HLsFQu3VUb
3oMaSn37qARDTkOBBxmdgYIFtIdJ6GYq7pMNnp5k8aS2+PO6dCx/Ke6rpspXUbII
PO1I0brLHIVNDKB3vBPzv5BnkLmmxPOaihdKo7cE3SWcVFHDM9BaJNmivK3BSz7E
+8jTtq94N7g1VFcVjyBpZcl+2n4cjtJhLUsIgURbILpulesH1Z+AUcT1oXxAXqlm
jiRA/b1D/FGaNvI+enFAzoJBaYkLKJpWXLtw+saOuF11LSJvkHmkIjDQSNMDl8vu
JAIDEJDXOAp1i6EwftSoQm6l59Nddjkl79ANUUecn9sYzth1qCHWdKfr48umLKlu
fUxckd5tZD8SCt1O9m/9fGzzVZfwHdTK8eEadqlByo3dQsSp8IbHzDj30H5/0JPw
+bnk1tWQ6vdjL+4+3ulxnbUZwEUEbvo7otxBddKxOZdWehF+BHVO4AIrNrhNMQtI
pjDBSwh1ZWT49r/knKadctsLskXLA1X7WMMbLTc7lFWinn1txgF8csUdRC/OnYEY
dhuNzlvW44lAhuVvRV67fXFCqW/Nd7kXbBXuEp9CT/aEMqAJt7QZur1tz/M9FU1i
ebrK7B41LQzXrozt11vkLjXdX2tK4LPCn0jIY0HdCJGFd07VfMk0SPPvWKdx3St4
yxzk/rY6lMbdwiHHQrMeKkNCa3BiG48Jr57hm6blFQ1IiyhQjZu+kves6mBCUhek
bXzIy6El4DJUmX96+JqhXvtyUMh0lpeNNCyn5wdhgnyS3bvPjEI6vAKoPp8sr9l/
HIabw5EltNtl6mRVxZnJxyXSDqDMOLQ7V1dqmG/RRQDaaupsP6x2SNFx5a0qw5ML
rwxQslO/rJD2W8pyGwfEBgY4S6QK2gH7gpvZJwIhuXAfZLMfAyHBkVXS4t/ZyzUP
dL+S8Qwuy2Uaf7w1QwkZxfDeJ5O/Exl/6roGjrvlG5Dxy7RT0QZOFglknkMHFK3a
iXKoBZYaVqDRQWd6cgjCSWiaM/Ko1cggOgzUvuC1uTt9T3aclA/1H0J45SAXxIGx
0ACFPJxS4x40FZon/hBzQ+FW9B5uZP/iNjWmKQhmvferCDxQgVhEIJSNetvdrd9O
2ROyB2gNkZe50VgZbOi88n43akpMcHUGfVnQ/DqdY2lJWuKvmL2xK9xwAaDLq4fI
qc5YplHkGz5RTqMW5g4tuf/N0xvzAk8pFMPvly4Mmvj4ZSUcRjmVX5xDV0mSghpw
bTERCzV0wJGeJjMp2GbwX45EptZ5QjuSej7REuBkOFGWPEBSpsb4sOAut+kNKo4W
IKdyGD1YMclQ7jjFuuFtXMaHp329vbKY3eyPOQ4z9WeFTdNTnPoQgd6L4lXt08F6
IxMS/il8162Yds6TDWI1RxLHYHx37x36LZY8kK8XAsVClCRYsP/vkS4+5f7VP8pG
sWz+leINROxerR/pCDfqXAiobU2RUpfLMU6v02XghN4OgAXEgsbQ3SxE1iC0Iq6S
EtqS8H/MpLlY4OOLvOVDhhzUcQQtDutBk9C7aeZsz8muMdIoZrHjXdywPtt8EsJ4
aVrDRpIzlIsQNxclPvxqlCaKTi4FedDnbdjtPQcUVdGBJWUS5j5gWkvEFWdIv/5Z
nL+6fqKLWKnxCGVrcR6H29HflTOcY05vIh/BfJw2qcyYJaugpU8y7xzBnqIfv4MV
xqafGGz89ujmIzbO6Pnbj+392lkEMNsq4ahDfRBO0w+SeTsw49PzYufLhiWf+vvu
DeqrBDr5PzPz/vxUDCg8gT8Rp1g7kC4IZsmQ3uXntX5g0uRvGBbO88iziCeX8TZH
Zr0a0O5hHAaqjQSkvrxNnhmb4GQqo4h7Be9BxDBXmphbzgJrb7W7aRblThaL/FbW
Kj7s216gjRDfwmUoQIaTSNxW/Cpo9XrNsHZHDKWQ+1yAFR/HXF4ntfpC5NwoyRlF
2quyasJNgYPeCh8e91Iwr+/+wFBQJ4MUUjEHDrS19f/cKOxEnN+R1gTfo+T+QFKF
kwEZkrTiI9Jur8YmQJTrdjuR+xqWVlotZaGrSLyAoQmsFKSh2MmLcYO4h5N0e6KB
2bZ4UIkslfuYgC3SAYTNImJ+zCAYCjpC9Z40VZHdIYTrA2wylmUieZayYA4BNILH
omLX8G4ZhpPhySDJ7ca4Xo6N1j1oeNXJhOzI7FHEvDSSgu6b7dQAWXXLHnjWhLsM
kqwleolvVbc0CMHtBGgjLwL9mfOGaAYI14kpceRTAXIrsqP42qajMrRTbkRKmMc4
hmAig5cb8i+n+2QqLxMYKLE43OaHilY1Yh+pOy17IzxT0LnOc6WqOl1DsRKNjMqn
PmxTH3R6cUC1ht1M1yorDViChV6ueIybSzKGsBL51O8GZExWoLX4tjeOeGyo5gwp
f/6EY8OL6FJor4tgbxt9qthAwLpRxb1BgEN+JqfDej254tPUKcC72b7gf3C7ZRL3
cnkCYdaX2OZszkRv4BzMBOGR9jLdFdxhScHmEqmiiwmx9dBcliMdKKU4jwTzkXKC
7aETSBBpFaaRYtzkxUSg3FPiiMZL4k3OWZ5zGspAEgRRrJ87lomHrAfDiOeTk6FM
dA2huK/f9orYdHeFsEQ7dQ7ipwSdKDIAPUdSOFz/woxzaxdAHTB+lTrH51c4w3jA
MtYB0fj/F/7EzewS9G/9u/ecDJkYIFgc0jzmFzk2xrvi6sdHVuoLl8vxmT0mRRHZ
DHp8zPcmR15Hiab4T+VF5UNKeTdMHM0ZjLsh6sJIZd20a/0BF3i2OEj59hScuG2+
c5Mo5SVL2m+K+xokykiIS8xQK11kTv0gwd79qz8HFoSG/oSs11Hu279tf/Puy0L8
/phoa0YMZjITtrpL3Xrz4db0N8LLD7G6ypp7VLAFY0XzKVTxty+j32WLH7bWcb5T
VvmgmZZpXzM3Xi/WFCFhNPmt8wK/HQb/OVaZ5i3smG8kIGs8J8Shrfaum3NZ3q/9
ywQi0x/YidBa0BK07RcRiVazI3OTYRDaqdOTeB6gI2sRY+V7jZSez8pqqauvUWzK
IkcIjrSqV3IyqSu5UpJ+BDT0SOOREbH3dkcUfhHuH/r+np6UmyL0qxf3MBeVWgZ9
PmqMEExi6BEAReMsmTO9nGe3mkYztetMqaLFHHUjWSGUDpRLsDT62UaRbT7twIvY
lL6RKdI2Mf4RfPtmz9ySx6w12Q1qb+5D2cBtv6hIM6QWrkG+//bv/x7a7tb67a/Z
UpDlZcs8W6th5Xt4Lhu0lUviHN2qEwbOFpLpehIaQUaQeCj7CI78P6e+wxyNGanj
DjpLDxW4NUS04G2BPgGyNNNB62leEI44RCXnv5Rqj6GUO/Z7qsN4NjM5c5HgSqNM
Tbtw0bQCHsV+nxHm6+uFFzIlNMlUgNUngOB01arg3YyNLRoj67C5xRgr15V+eHO1
8YMAVXnLMZg1tIMCLKKHZRUBUYvQYU4fhnwxWzwUN1E9hUpCVV1wHwOboL5cDY/P
096WkTYlHP+5nfQ4cFg82GboicosoO9Kilt/DTKBVFgg0y06tshCdNEQRnQczXdc
mnfY/aW2OH+Atfq1VfEy5WizW/2ocRbFit+XeT1W+ZT1twM39dhP1NdWJfjFXrCd
89vL1Cgi9BhRc1VkSUNnvdnaofU0ndtxQz0G1nUkKN+W7hPSxcURcCrGh6r62+wy
AzeKG0avYGscad9B6RHeGrbjYqmpm07Icmq1T4wrp6/aT9VxDvqIAFG+TdLamUYI
gbG4wuOF0ebWLmSArERPKdLIfqiuB2TclksAcIy8WkHxFx+jXfR0e6DW8Mk5JA0h
q31V0GFyc2OOKoCRQjiUiIJJAGljfJnjfc+3KQGdIZoortRddYyeX68unlvbsZoW
DsZXNhbQmAPCpQ1BqyX8ATuvNNdFiLUp5Uwr5tu6rTinzKKnPtltPPxc265Flmeg
iTYtOtw49fiyBufqnnqPSBPiFHl5HaKs6WqzldQsZt/tMvCg5WRSSxD5wOpqr1XJ
1ydiTl84/Ajftm14L6n40UERInqfUFpmKqZeVA+jzzLxW9t6vZ6SkloB1jDXxnh3
oYFkArzZf8MKzX+7htWkSd8Hq6ugg95nRs9yMh+RiOGCjmLvUSYBuHXh4noG9lnE
F1iYfI8nvjzwSUGdoRHFTVYylWj6WilpW+JAWrHilPCqsuibYHv6ObXhX3Qiz1Gi
mE9JgiQ+spq9wBZ9CuWyGBHZiLOAEvSOEqWTRaEjehE+Bph+ChEahXtOahm+Xb0Z
jgzpV6e4F/3B9LHdfZeYhr9KHPlEp/h5Bk1ZkSlaDxBHIux46m6l2jbHwzbKez3o
50E7HotlfNYNnwTZaun0eiHPTt/8Kjc4f/GWLRPetGcwpFzYxvW8SrTbK79wPsUQ
0uYdVMH6DK2owVqo6qSR7SMr35n9u9cEwVDULqAdc5wBw4GlKb+0rOkDylDngVoB
7UiigX7qh4idRHJsA4r+BgA+o3RluT236zUACmEOfkle1d6fGjIoljVR5QKgsTpM
1szNf4NA4zpPb28r3t3LLHe8BQV4tC9tC+Fm5soXfzpFNq6Lp4haJUWo41Q5o2aX
o/HX/Gk/132PuWqR01BOGSo4SO3C+OeKB0BgWrrMPALdtwfYYKci8ww/tsXJZ+ML
EYesmdDmVz1BPOMxlnb7zQKRsts7aZCeXSzWbBmGXhz6ZGRwnE30MYViAH6+yVoE
JOaBonsNLFJZkbRvBY6Xz6oNw3jmKPgjnrLhdsCkkNU1ZWpPkIaEdlRAiUew7qps
P7d25dENWFcL4ne8IJ3LANklxYlFIKYGfy5aBhBJQvvC7ONgvWIEg09HgNMFPoi7
jNiTiubT2gOSKw2Egkee+FN3CJ6ELUZauPffmU6PkXST7H8Ir2xr2Az/qDz6lBzx
bvK+ldUN3BXMMHBQYpHVthPMErR/NXn3DYUpISwMJ4E8EZcS8FDFwAgQoR/Ujsj5
isgIdyYBQezIcYIDVMQ2OD4Hik9DosWg1oNwiRrtN4nCgaZgnRBvsSElwtK3stuB
XnBpG+luxsE5h38mPNitYTGHWbv05Ya7WdS2eOS0sXaqdI3QcPR2s+Wgw3bbzdkj
4QEKbMea20vjxCo4yeRr4BCvdwPntVHSTJr2wXeMgQqXJrAkNuKi4CJLkW+QEPAx
ktfxu9gIkeTWiZIpqhio0TJOo1nUdhKHfBItPWctekFiZ/M7nEXjIu76C1JUAwAc
xarYpIPpxAQPvpjxV1vyPfl5P7RpkQtP9QBUa8OWS9P0BWETJzKF2HTWfUjCtGie
OwjRynbuMg4wZZdgZ0Gs3jGO+WYUB8GofJOwCrS0E0F7IfqkGWgS2iL6wvn418TN
IHMS1LpPABTei7SlqNQtZfMNY/6QGb6hSjQpMecxi95bXqO2gvvfg4PiZQkC0mrN
vy2KzGdS934Z2Zxcs+QvvacydL0JsLpoZwNg2sWECSZ4Zm3gngrWD0SHqTrXh73u
WRqfQxBRlZsSL7IHLXc+UDAMlsh2AJWwi0/gwco43SZiinV6bK5nO6gTJhRXiwEZ
jF05uPPyQN249duGxSmFVpOVoCQUms4h8VnzNSJOD0AgnlujWnn/Pg0QLVgkT9wy
3crDYAdxuG04y6qWSwMhO/EWdoD0PlMGyHUMib5zUxG2qVBQZPM2uslNL6C/SbVq
9Se/r66SyWhKormfHEc8sSShnl8FFsQxNHp1yTr6ByzxButMcMN+SlxywtvwjXuY
lGg7fQPW+v6v9mxNAkAx2LofFED9gKIGTHHna2pPUSxk1lHN5Zv1vRS9lbch+iZI
cSVcfUcz8amWwYN/eVHiSHRDrJ5ngOvsoVd6kwg1VLJh5H2QvV7HvI59m6Tm9A7Z
RxMSguuZxVzKTS2cd4lCUC8NWcgHjVcQS5kxOw4MTljbu4L57cR7SRuYOxNe5yVl
EyLkoOAxEO0ASl4M9c1SVFirqvjBw+iofY9JDbrTdmIuQHDkOzcm83bPuLq1Wv91
vHdZp2XY+Q1Y31Qvqcm2hXKgP1ED/MH6Dpy7o7B3kjoOD86RrZdSX7oRdGPWyrDD
5kgwNPiwkMDbilmo8OsUcpizqnTjQVNAVeZeHMMtNSwyskHJOswByrf+GAhDRbF7
LXzrN3w3vFvjaZxO+iB6JmRadRCl5rneWBOuWtJkot/uPBIBVeZqtWnm7LoFBfqR
g2XRIo4/VxDeZOZm7eYc1wDxCdXhMxcK2ueUqx2LbZxNr9ZDGz+xdIgBjo/w5XU/
XipUUjdDJecuKHb4yuoVzYJLBUc+KdAIdWbLXwHOvr/3dB9mkuhyD61xNv46oJOJ
GknaBjglY7WqXd/Ndy70m11Ns48df3dR4C9KBQzvA/2vxOc8mV/Gpm5IR4jIGvJH
R+XjXVgS77ZbrnjM8vd4QA+6brrBFJL1GGzs38AIpJLrUKZUFZV6lfH2Q5HwYO6S
cgbaUPJEKsiqmDkJwz6tEN3N/23UvGEvXc+rhb2IXz+yaFZkdiMa3CMxHjZnz4mR
XKQnEyR6FzVIKFK/ve9E5zGQ+UwFnh8JNRztjCgZt2ZYpYIwiIUAVGBCWOJ6cOMs
pjhyyF4NE6UatLwEa2herJg+gbQZ1jXKkdb3TcJut5MFWRQYAIVc7fWC/adW1uTU
ZDGlttAFQO91POPBMjKXHg3NeRMDo5nOJWy62WW7BrtzbwKIRN2u5p/hnKIy6O+t
+LYjdPdQPe+kFxZVx+Xer5g0mZjJ9UY3znjJ9qf627W9DRLYj8Yd8IJjJLZOWfwV
WT8i1xYZHB6b+7vxMo2bAClxwwcMi00v5ueC7jy3c6LmZtt7YVFcMXz1OpcX6o/h
/gOTEmHNhrLtcwk3FX6Lk5TD2qMhTg2klXkB70y6qByFfl3fV14xfcFj7Wk+MSTV
sa+AETof+PoNl8Es4FAJtFas+ywX9S8CcsCxM9OGcNnUlVtP3yGb35Vgiwc16mP9
Wu6Oq1G57y4fRAOi3b5eoUi4TwSDvLm9BMxUVT8CQ9zO0mr2zhQnTUfyW6C8zBGF
tXQHUH4B7/RwAz7B8Jh0QVD/CBefq2LsdVSUyFp7FBrxTMeJPMadApCoYE36TnFl
mJrntzX7jJisbnVLPqhEXRda4wMDDWv851kQOm9GZ8JFI6CVq9zl/BYQtAumQYTr
SRs9SqP0HeqAe3+x8byEZzYXqBtSjh8xX7SfvNhYYqB73F9Jj2hfGDyQ7wxReGi0
FnbijvyyJAY1sXRJe10Z9c2n/1o1+FTQvkkLYv2K7C4Tzorkg7xlE5QWIbkYztkH
VgXwh+ZpCobiZOWLvZeYvnT/gSe+o9fLsoFWAFbf9lPefKiGexFMHrOvCYdVdaEW
b75X98jt5M45lKSZCWHD1Q958Z2n3MZ5117meOTNJ/iF9saNXw8VbZSIQ0LmCim2
6b9he0o3YqQ3DLs3XAfuGwuWDOBdgkNDmdcGtaGXgSWUVgNbVxVrRGhCfsVvvG49
l7luWcHoVbByzMW9uANztSbvmulK3tyCKio4u6HZiR5vnXEiW6l7vLWUAzqKBcAq
lfgyl+0gF/MMH9xLLzHKtSIJqV2SwSvSJNOP3reY1SPlf0iZ5pVDXWnn+sEpBTQM
0cfo5Cf8UG1H3fZu8j3XOgoVbLmNs0J3WBLkEjh8slllXwDrwckVwIxP9Z3zB9V/
3FSujt3h5AiiO9Io96lgFVAZDDWEl2J0uROmu7kJ/aeKHFKRW6wdfs+4mGr5Zsru
PfZFO5VJ+HgQ6Wea70SGWR4+w+D9aam3NXIV3kXjSrjHpNmyVmtujF7DMgH96Sqt
jCV3Q0DgjO2mRQl981ImXaC+C5Hv+tNlTG3OMg06rcDW62DsGaVP788PtW6HQf7L
kkBrDrRkGu1vAhHZSy5GQA0z3LZ9iQs8iH92v1M+MUlT5ILFuOxiSf6HxV2viABW
9pfd8EX/OuVnN22cZl8Hra0z5xsy8MpTKBLQ4asWVuj4AEsxTv8Mbjd98hzVxURv
a8TjqLmKVG3dx0Vrrr7Rzm/AjiY332IKXYmDrVyCNdo+hawEVGSbsgmpqM4x8FRD
c8+TSSX9Yuil9bBCWpHUD30GYi4kPQ8ppHlGLt5bDi3Wi2xz0C27k4TR+n42DBFS
DOOWCffiQRR8MnkCN0fK/LIy0+GTTv2g2LM+Q9MRIQIQEeY6H4JXo6GQxpEdwmSP
gAGE5JSlNDEys5lBTfopAO1sGedlq+PZBfdZHjCy3GiNJQxYjZ0sxh94TNW4LZzE
Bm/FnnrIFBBilWDCO2O4xCwfLABXkaRQxA/UYFBAf+bncG96kaVTGf7lqJb4tN3I
CpBcyuFDZEeut33S0fbHYwhpLLqOcwGzI7iD/YEXSYCjrXE+1XI2f6OV1rQGzFxW
nqKfKkeUAhhy3sEOrRwSHqL6WnNe2SgEnqxMjyARGQPMzhMoPvXTs8JKrHW4OndO
HaG5YmDA2m76AsY72fX9XYO65H585SxyYFN29y3SCDjcdLEXvC6kQ3lZReq+u12v
L1ucXHYsZ1UyrbjThLDh/BccTgVzwtLcc9WR2UAhFw9qKvsQN5oBUJ5EEY9tgn2L
LLBnquOchcRwZqEHx4yx2w85NXH9kjLZX99n+Ow4wncfUa11RUQlV1wEYr/9m3ub
MJ+hoZYXJIYdTLBdHRQjPe14iDKqDKULan2tAqGnJif3JL0/kA0Ah7YSUPrBSJw/
VtwVP2CVAanSDY4UdBzqcZhfo5qfhuaXN0R7n9055rNLVWXzqIkCVn9O23tQv0ro
4+g1U75uzEe/t3us2SFfl/yXMhTFeY75INDUq1QOGEaMNtq7aoTyFPNDQUMeuPAE
Vv1RM4dheQyYCzPSgZ2hEyvLqZOniddcUZxmLBegvoZ6Wcv71HINXyEWynWXXxXM
NkZmnFPcK8zsa9yBUCN6ZvpF9YyPGCRgx8S524R2Og7RjEesLuuvfRbbyy6K7nnP
pI3WRdIvJO9HEV7xksyH4VfUol56hI6G87dEAvTnHNbEX//8VRUJwlM0k9JsM2t6
j2XedGxYtOI1G8yyE4iiydwcUzZhzE4CPZdEI1/2JN4Kr/uLESe0YmWIp60owXaf
5ZPgqwKNk+Yo6Z1G0rpCcIKCa8Ey+/qPGK32CyMc0hMhLmRTzKVddVoucfJhvDkL
R0H0ye8fKBGRbQeidWkVqiFkab6Le8/iMQC1lZriiPrCtZW8YrCEYHbrhTGNzawA
vTaicKaxEXFPHsSK7U1dOgkxp98g6EIHtv3vFqSEXo/TKJJa3XGLN6Oeg8BABPXY
yjUHaaX2rzizXrx4djT6/rLdFOUmPrCzJnMe46OBmZs3k7cYPRxQnZV9o/o8XmUb
msCkTI8BVp59Tck+pvhY3Hlb4RD1T1CLPshil3WVV+7P62FaCIbwdtus430V1GtC
glYf5rU0wzDj3F5WwvZc93G1196P4KD4XjqbVwIDbdJsUjJxP41NFTpIuZgDlRbs
/iX0LoyVMrLhG4HcZk9md7Yuw31bsUt9mhcNv9QVqTvHBxcHl9GFEK6t6GX2cGn7
N8vSsVAsXqxtAtFfNad+UGY41ZbzOSdRJDtEqrsGUGTS/1IS/mGzSdb3MyMXicX4
vrClmmnnsYaklgmCJnu8rtoWoWQeFjnOR+DjymEdQRujIMgdIH8pT2UiC4kxX6Qf
xiF3UQTq6aIht/iXUiU074WAT6OVvE0EXK+zLuPmK8mDL5/uFCpA+iwfwBtRjm7t
/oykGGc6J/RfTzBlDBySfF7oN6loV+r3Go9TMJ4cnxCShSC3wzZoeawyHVRWhuAq
hWd+0yBm7iwqubHhmy39NUPgVYb0iOI8V6pDG4gju4B2lkf+BKaSPGzDoCtoqkkO
r9KInu5vqj8ZfV0ev/lzel1dsDMunMGw5AZFnsV2ho1Wjze87iYflOIM9+7/rhvL
HkE84lqTsKRtjnqARx1pftbct9Q3pEDoPVavX5NoqoOdMRQOkT3vV80OvpHFrU8Y
nFtO4Wsa9OSSSNwsxW1AftXaKCFZhNkZZijlYvCXYQ+73O/j5lEa+m78ZPY/7YqS
BuxGoBthFdRn3W4l4z7DtdM8rdNmjO2IB5MW8b+YHabGpCbtq+WFnBHRc5szeiuR
AxlIpjDjt3xio/mIBjrXvlAI8cIXm1ffg4HZMCekhxLBChljRTBW7jooZ4cKXycj
zIT+KIfQZO0lfDuhWLYQrwuPDUuttIuX10u9LLJ35i84sDeeYVQho1/VbDcI+sQs
HG2ZP+gVRFR+EctNoAmo2i29ELP5oSZEloZnVFPqPZspCr9Gvw+1wSXnCwdTn6m1
Y5mz75TRgL4uLBDmqGalK/DQRyFnqkSIObWQxuK+N2xhgQIewEhIRHYwmsEXmjEO
lccqO0lI0PJMGsYZVGiLkF+Qc2FTSOPvdYtKdUaqqh+hNX7HqshkOqzvEzKfdtzZ
fa9a3vwf/JO31LIsK3gaa0rQq8L4Wu/w0v0ybV7D7JzzpJqIePvtvM3upAqSlXot
a8xUdLdZiQAd3paN/GpfhsFOj7/ElynQrrxtXXkE0afCBWxOaAFYpeMLnEeTNWsM
khUYuYbs+zJDIYGTOw9azHh0mIR4SqV6NkE6xpUrm4N0Rc9tHZQZbWHHDXG7G11e
OuKmtHfK1X+9aky3L/9FZ8fOioZ5Vy6Iogm11kMEV6tj6atBBFlgY2gOw41RMeX4
DtJqbNWM9lM2NhkIbPV/fdyQJrClMUebvcUmCAwfVm0HlGlRso2aduyj6TVjIIa0
qsGwXu2gsrrpz02dV5yp8Ej5GiBcdR5dv7y3ZwpGwSFwbk0A1FWj5GPj1AT57YfN
FzVFyK1ZMdeXDaWztGeG/v2U/tssQ9mpBd6uIs2JX7hE1hIiemS93ytgFqMfeTbT
/RRY18m2mt6lZx8kdKS9C7RytkT/PzdVQKTQX4rZjxz8o2jni4sxiUuQPmkXbrtf
r8sGsGD4lwfotQYXGwcVx6AFISeDtudhvt0Gmv/8rEhE9Spkef8V50owaplknvga
M0khvvNzjKvGrEZwwHtKvBDN7+xVyFevCDkxU/PZu/GWH9WtCf/LDZiyw68bI1VC
TsyP8Q9tLLm/B77scubDuV+vmvOUwKbjDDhEO9i/sjnJOJmeuRweRw7sPK1CU7v7
Ys1UiddT4zcDqko+tE6x7ohKIc3DslptiLjWX4jhyiI2uiFG/fSQllEOAzjhBzy+
XyKO0qKQ/T2fiUEkc8I0lQCm35iqop6p83MNzRvADG7TkO2lJHtRwZzJCWaz40Mb
JprTXiWEHmn0rGK9upMkkpEuTgfWqm3sE07+66TqgzkUyYKpbndVholttYx1aPO+
sKb1tNsLKaWCuIRhDk1je8A8j/LAFo3hYXy5lH8eeMOoFBrmcUUy87dCyPbZ2NKz
e3UVZzmsMVuJ6gV/DZjfgL1rGqEX4OZ6X21wGvpsZ9dvhF5VEC8CPWZ+D4YD9UrG
TW583Ingf9h33Mk2RQyoFcEij1q/ldNQLX88J4dSiF54qsNeAmVZXWvTMsrhLSkt
ayQGpat6qB8+wiQbg6hJiqlhKgyta7lpmrYH8axYpnvTtlgbK5qmqswO0N4L9ZMK
wlk0YdWodl+jA+wpbOEqYF3Hp/WqrdXfJGtO4HQ94fbkbR3wK1WM/OhVcdM7a8So
8zjUBs/VhG/mFcsAegpxY9lsMmuHo5kqss2HJxKDFrAqLt7rQ4g9kPsr8X0XhD+z
YT/n2hrzUqBX+Be+30xPkSL6RSSgQ0KLABrf8KZ79hmMGyPxd8AqTFjDncr+db17
zi5GrX/3ihFPqV1sP2kO4qjp6/ItE48V6FErHLPPQRYe6cZ7L8QeXWxa9FZFBUhk
mXgsPEh3xQczQ/wy4BDQCoSpJU1CCJDrzgrQLQhrazq7c4ft+qhitlPiRtPA29HT
9/Zdz/oDYQFOsywd9eMv8qKhhYYhzgHYfWq/eZ8isMQ3ak9m3WlY+ttNlbWIJ6Vq
3G+1zLMDVUPY3pqObAWbSQHlwaTdAlcfmMR8lUUDIrXIyPBFLu753YTJC7dLJZuC
3WxpMNjJVpwp8pKsu/wRORHvDi5rtZd4j2DH4hNit7TsWfH4dFd2nbWNGLaFi+Tj
+brx6yWhCFCE/kxFkCecIJYhyrmfUF29MzLeIMnN/TiUJPml3JM8fp2/Xr98Jxnn
z6o1mb+lCuQS+ZAXFMvqErXC/LXcWdMN96ncWCHfBgBFfWL37kiAnv0zWNA75ilp
cgXDCB4pVfcmepX3t76bgBNbDuq0VDYbN2dLF/ElftIEwL4fbciNQ/G98sA75rMx
HDMDS8RINMv+9Wya9vE5hYsSqVOloav0e42OoBLtcaC6aNWQUY3Ly5M41BREVy5U
VRCnjK8qglPqFMKzpKPNOd83qxNqKxXGqU8hZN0X+RDiMd0j5sw3lKQh4r2v/ekv
KY2EZ/NWQIGLf9b1GPwB03u3E4xRrFZ8hjednPpe04PYY1YLf7AG1OQNrz7gsAzB
tdDnGDjxADryy+eV035N63CJaJXr8L9khM4D23gei1cuee3QO3NX+Q9S0GW/05D9
fHDFk0RNlIZhwBW24/xTJO9CWpBa+t7j1muL53x2jhgJ7BDN6mJvd7Af213+K2WD
FtDGuEmfCY0CFrTurZ3Al/AXpeyFM4ewWDIXDdoAu8XlQomVXgJongLXKeKrkk03
A0wHCpC3B6PM0g2uOUFxMe0dPVx+0wN3SH8QsO5ilyXfNVfJKidc+KDm8Fybc08g
rCrsLJsFt8fB0c/yQNFZqy735mXMmYRXP3KJ8G2ZP0zVW08q/O+37fFMuRaYe9Gj
CUgVwc3pvxkp+79bcn2870iLPVmjx1b+B3KW7XlNCMR7Ji1BxmbgY7E6ctk0fvFo
dwGifZqpnH7Id3q2W23E98B+Sd+BBOKSq9OkVx+/BtPA3Xh4SLjG7LZQNTfnPpAI
UvP6a++BDol2CflXXchSoKLF41QRVDg8Du1CDF9WIJbIZQ4tYos4V1XGDPtFDeEk
zfer9RuyvKJZjtYdZtbFYQXFl9c2Vw8E20iV+ekkeTYGmhivf6FJwPEL0EMCPjmW
VcAepc89D4FQ031qPGMoLlO7XsytHKJPvt1UZllJqQw/MuGcAGd3nK/XCcz6OX8I
n0ihprPYqGHSFW9/g+oZly/LkJqVimdyu2+gmRhdOtQ5qDCVXtRkKyRmK1/hdEvX
Yt2HNlwXlq809NMT0Q+Liu3CdUh2g+/QPVhd5e1yzxEUU2g3u57W3vQxU2Pnb0gZ
MHfpKupiV4h8oXZXIQdA/f5OezxPhthOI6r25CpqYkunGHOlifCkCA/Eyi9LVegN
dlxjY9rC2N5cXtS68aZCorlJvNVnf02AUdSaCBvAlfomtEevj+H8x0Di8ToLYhjp
LB3D5t/LRimxCbe095gkUD7ul5SEpSVeNT8fMDwIjyKbnGfWVAVqZQQDVH9QrC/e
KCyMgw0UM62K3aBf1akDyTapGVcJ9LIihgTHQGiF9wDxgLUUkQ1a4R08tN947Hwp
mMYylg2z4C3wYO2AVCyZYYQa+P9b1lXKpT0eMzhtlrNFy/5Km8R/zScs3lr+px/k
V3+eSd9oM9uQYMZ2iDt2d7H6cFkvUYnHVVg0Ig+0986ZlmDyGiDx+RQn7uiuX05/
jm1DajFffccANDOWJHlxXWdPOBYZ6QwJ/Ea42Qxbg5aFK0OWO2WPn8ROz8i6wUFL
wZLVb/j7fvXKkLC1IvbrAG3ozfTq+FERwygIPMJtYVPpI21ACDlgYXHms52U+GR0
sLawI9xqN9UiVW7IPnozXcWSv5CPFlxh++EQTnfdpS1ydsFBRwZrOE30pviOQeyj
zQLzy3dTKyNfMLqlIHI2+hMoGygj5rvh5b96GcyL+qbbTXhAvvStkkuju8MB5Jaj
YGA1VWFJk2sQWV1/2B3nDLK1cq0UbTbh0ZhkLTFRvX67/98Y9CzkLP+6IPazT6W2
cy+vZQMAmSuuW/QkN1SVXtr/QGsxoeGHG82YEKYHJbYHUNvI10MkL9Q7Bnvqhyiw
mqB6Wb38+RD9LAWdJvYyPXyt7s809eRIvkbMptgD4d5/ekkoRNGJawH9/wTD5tVg
tR2cwS3FOZJy+AWTDOKJpFJuBlyQ+n4R56L1z4Qu9Z71FHPFRLEKGt20tr10G6P1
FLeEIVpFUbUNLcqG4tsVJjXTIDu7Aip8mhyzjqeFjZlaofjiNNBYSjYOrY0xQ05u
R8Jemr6zxrRA+AFVm2UwcvJGwCNV4AT02kcrL17izmkfQESwmtDQ+D1qOTMWyNuO
grYhJI35rI5+domZ0Pnw+AQgvq87FDE7aktCZTW+G3hdxRCtV84QJt68IUSV62fQ
lG5MA+bz/WVahq9d5Xtn4jHpgmxxAZNsp2gvIOjOYFA6BojPPJdcUTL4NkTDJ6p+
bQKpP8vphAZdpWx2tr4WT/Te3IiRFUCpvCKREwUqt2+f8KU3iNsDHYHvysI9QUnX
j47QESog9BPPTr4wI80Z8aQTunJLxFbRbo6mg2D7BaN9+JKLdRx+U4jBJ0ixJNYV
sBltJU2H7eviVTlRoNlhLiikolmfvo7+Q/CAX+vVWQ3+EMKU6nkGN8g4kDdRV5mg
n3dlRJdJx1+NKfHf4E/WzEubQYXhRZl/yydIm1Ol3rSJdyJn3suK2NRlU4EN7HEH
0Q1gVOm+E5itFGQ3gadRhZL54WOJoXnmQHg2vJl0fVAW0G7YpW85r97q0fk4g88D
Dg3aYp2AAzTUx7ea7lFuMY7nH2CAdl4nuqFJSdSwli9lA6OpRrRsCAVFilgw08fo
jA9JJ29ZOtbO2NlTIYTqzA1mGncIyi7wVsRude2DgP5XKwS0t3lEJ6WFL2+PTqLK
nz3jvZ4mlj5YVXMGPAd6fPdaVP9soz77DfbkZFeiY5hGfbGvFRwV6azPND6+ppSR
L8/6w5Jg+oS8awpKU2N45JDAFHNxG8fj7YfsgfZKHXzQaRxXZsveedjuJB0r4IJA
xFa4W7xHRnPqy9ggsdUUbW/qAa0C2gB2dNKhgYQpQ2/IDTUMLHZr0WG7DkL8cn/6
QQW5UVzbY1IuTbSR6npQs39QtlYc8XBrWU706+EAIHpebtdCRrfqmSxxHjCO4PXt
Ib1U82cPhdW8uNLj4GLB80QlZGoUwKGKN6zJ0xONvcqlvuK1F3xLESiJYi0dia/5
uFpbYe0W/j12ofEtfK3EGY2GrE9J6i9N55c0WwFB+t2GUmZ0xIW6H4DzhM6Q6Grl
HQtxtetBAuzAdkeQsCitQd6xxVR/7DPwZjbVKxrL7C8BtOHXpxlbsK/MGubAEfpT
RTE/BN4cCEQcr1T1cuIe6+2eJNVGpDXnADlNe8VbnVKsk1GxojxTPrh45EgDxJLL
Mo3BAbimGnHyTBDY4wuvtGZJZpw5kFBjOZBAlMWqm87OpURQpRGFXjzCWugQK/+4
juHHiqF5JB8ht91aOnM0QysFqLQSR6etGHmw7HSTViHM1Cdr9z1rJ12iboCRB1wH
U7Au/gUhYZTvagHmweZfWLYL55+m2ITXsIPcc2l9DByyXlLV2soViow9ic2MINt7
sAt49MZKaR6u0aPUgAK6MOLrRfE+ooyJMV+v64ui+/yR2afPcJA4xvny2epDi4PI
y3DIByVxd3c7m2u11zvc8unpaePkyS4crn5sbBFxHHMNspGEOvkwFeOENB7AbMdi
wzyATS0ktphDLNtnOI5VRkX2aeODFEdQ1dEhYYqSpow1QnRqsdkY3hXWZu9GR3z/
cQ+XGd0JqNH8zvgm8WcuuCd58wj3VKs4iBPwbBFYo11fCDOqSLNxKuzDKLdmi09y
4ApDLCkBwlTmOy3yz7fu6FmDsCzjJTg6eBCdJkLrWS4IhRcJ3w847h2UFMCUaWwF
IpHkDZKNirsINNmlBfQJqO0wzqwZlDiZJarGae8iEkjZfiSlE4loabrzso64EpXb
phGj2F2LIBNvF+SHp0RwWsRD2YtrzYBjMkz5IcY/dRhNKXM/44rlVi2RI8pznu4o
qfXIOsneEoBbzDTumfA8p7ybBKng7F9fANdqyhWLnctQb/H2JWBrb5S7bVVdtve3
jZbO3hOw6Ec+xAg6h3sFpl2Ec31UzFX67/s5pB6jV16si5NHcaEFI6rteZjFIdIn
LJz4eGCUx29AoSxBmYGjs8bZ8MvxO53oexAx5KSKFKF6lhJxx7l9mDB9rJwlPtxO
fH5W6DSiNX0ZR+lTlLP4xUGU+rtBRYXYK1tFOmffT/OyHdBYb1l9XRzlRUVPohNl
VhnI1gfg0sjBqhpNXJQm89MjC1U7HQxTLemD3aMVd+KqSf9bDepI0ksWL6Ne/Fau
dC9Ig1adQIURkwwj0lPUAvROyAtDtzecxJp96TslNdAxoLjYQvrNt04SGcBqmswe
YCwf9xydMATY5tFqTWOVIwGsdYeijOnbZLsF38U09pSed/IV8VK3TDpGnVPv6nBW
j18PekPRvAtGRZCTfHVdlTl+p0ra4c8wgJfhyexquXeHncTmZMZoExIaDT0wh6mv
FvZbyA5KBDxqxUGmoBJnZIELA1en4/OX+iaxc3lJXIZBekOM0WRebYfvEw9qWGGD
yprRhg7YSMVokvCRlBC6tA5CCFjlNfeipHghV2c3E4FnRL8XDAZw31r3qbNpqD6+
pJGiKUcUA6jF3ulUnU6Ue2h7uwM7JtBChJbRzVhssR3NvXBNdaJ4pIaFuYi6tICY
w+P/8MhKb2KDNn6vIVGsdbIWtpaqIVTMVbrDoBvMtHOeIA2S2kQwjbWiGhzotwCk
XPUDETLOPH872YrJA4Cva6Oobpq0xBvr3gcZfYbVPJVICmI1Wg18LyE4Rp6gGOyP
OCJ8CIPyBji689i+HcUZZRBDTkYWdEanQRjgIJG/5oAW1x3GMnF/cGeVnB+bqks3
tSUXhZ47nifwA+fYQ7OA29dubaKiU/ofQv9wpPc+X+m/DbMsYVZTA9RiXx6A6K7j
F2pJv/n2Hejej/LjvIhWo0+v1TH1jDA5PSIWBlDSl7Us7obte9Ck48jyotRjrO5L
nyuZVzwhubLqAYpdPoiMIjmdRcVjBnEnLzTejHThBzSNg6by7mY50FYXUpJrzC7H
ZOC7QRVhlAZICMYm4I84ccbB1EiMT39jCjrjpDAkbDLggN0mHFvxcgBu8UJXMdgn
X+T99Jr2OAbl590Is/U1ESvI+X7sF0mcb5TCy5pDPYjPiodk8wLEwd4pwlVRM0M9
idas3PMfoRgNTfuQA/8Ftzi7uxGKnHexY+M3kvGzPJoeACkZp5mDpFcRXVH5uA//
M2mgH+J1ukXVAp76dafkQdXTV2XT90mov54i1qNsH8W+TbmZcjtCB5rw5PFkJGdp
esUa+vXSBUAAd82CuKZiufoT9hiRmYumtxEcBqOkeMDsOlKCJhoxSnxSvlxKbpc3
M68+vwumtHEtsksKeird+I7gCnCyuc6RHNgifaSs8w2YlxQSmrxnL04gW+eDeZiZ
43g/0pPpGDQucTShhDzPle4akA3uqOusm2gCDmCga3pfdRXECuRvygz7PfpHNGP2
3TxIWoV17EgeL1cn6h+LsMWYQbx547WXXl9Ff4QH8453HU1kGMvz3Ua6u1YkbPne
zA+f01i10hTaJb7aOaMXZhlZjNPulAdrzmfFs6VCs7pUWqFGrCYTHgahYYcMHvNb
sdM0UedzEH4YBxfjCImjorc1M1oGjV/qw+BZ5Pj5I3aJG3zqSnL/a6DlpYGuV07Q
exSWynDPPj2Lj5yJZMkNOWkW61oSVE0iD3teoJKUEV4uAyChQgDZd+g6kd5QGFiD
Dri9r3vTQQLW4mbin0VAu/jR3yvXRnT0QoxgPVaGcudOrlViR4y1S3Ios8pqJe56
CWSVVTPgsffGy7fcigZM16Ydtl9U/NwcO3HXZbISLvhvKrxafTiYkJSlhBWobg2D
lk6+MORuq8wIrhBfAdyaGLPqG3hjLKDKc6KFDrJOgqgVoODzYNkdycva+sTuLeEX
/b705Pi7Biy6ajBxHT8lSc1X213jpchBpOi+5Ubgsm634vf3MyCjc4rtzf8qYIVB
uNpwToQiT0ELEPExzki+vfx7YW33u/4iWcWOJzjUzs+W6Eywr6RervCiL+1kPaZQ
omttDcZ1CrjGCM0jyQN57q0UvmoeeqVQuWrp2xDceFLKTuAF/Uhsi4BhAUbsnmCp
Qt9Y8ADx6zicmLm9HIEM7Jkvgrj5T2fw27ZB+WzZZNWs0ibWKft8AHhMZ1UQgbhh
FQp873DPGJsb/UrtZvTnAU3enzf35ZyS0356QlBvnT8o15m4CiKsQ68jf7AxFlBy
U4SM7RJZnJOaXxsy2euWG8AY+3q9XIgsC/EjcSixzQcPmvfpHuxbBsFeVnYQZ1W/
xRzIpTSR8s/T3+A3EBRWodo+LKDISiWzrDpHiOMnlX2aE5XMTnZr/aGEXtEA1lbY
6CgtGucIbXgT4/OHUR/s70fndWXRgwdU3jTN5pXykq8stPQbfNjacr72j+j4FoOd
8m1JlkbxZ+9NTYHRCSRnosKpEpX4FSgUw00JSTqnoHKtkD6ZX98Gch7+KiBwmRqW
rcwhcEs2hVT8rG7o8MI5PRKoOpMNBn5ZsYjBR4njm80zAqexgs/icCccOgTs3VeF
oxl3rO7Qh5VbS21hw+hAhNtpOEQnmnExUDqgCiJjrfwhV6YowdN1btvu8Nid/+mX
BY4SRkOBVzX1XyZawL0g6wmuyuqx7G97MZCx/fnx/ztS0jf3CaKq1S0I+1XwGhr8
cPw5VhYciXIHHOVijNdtIO+Jp1GGq1LChTqMPGdxaO8Vu19G/2k4OfzRe5zkYw2n
VksrjYPYvWSwAmQL+lFw16R3HqyxPSPeSpIvy+TQK1LX5R6W8fUt6yXoD8iI8lQk
3YplhtApG3PzM7j8lqYbQNcxCkX561Q6obR6/gkJfGeSsxNwSZagjVsrVHO9bZEg
V+q0h3R5x22MdCJE9UMe53V5HKXi7ItULds2fNM59FKrkPfukL+oPJtvDkFuqBev
PbE/2FEblaYGmFLH8WUEX3cIqNYijknz77lYY+XZ+5Tf6Lh7CHfPhmA5+wlk68f8
43MW2DkXn/P82Q1dis/b0zbLa4wzqupsmiYzAIhMX/UPYbwgtBrCY+oe4ze9R1ZT
BvM5eWubfiqIjn4b1vfTCKS7vpRd6I/FBY+VB41FmNpVIajWmDiV/MCe3A+ZGryD
s5GC5zUMSFRdybXhkvW5x+C7at5RLW6dj6X+fmwGIaE7pCG/LOhhNkp1JXt28Hx4
hO93FB+EvtgGy9DxrEuHOuWAtjFlxaOInfZWESdJHn1ppKh5iSkuvAyEhO6MSzxN
MtdLMufUFgUrpzZqgaIYxSuC57uG857fo+2QZaZ/xNU6PrdLNYUpshD9PSnE5me/
TmKZiwH08s/fcuAyoOvKu3+MEnohwWCqgTdM9v1u0gsRGOiFhVGYlLt7mJqoR7tG
mVbPuoJlThsFbgwi5EiAjPdT64scRgc5PeMfdK+GSc8cdb8i0+NNkgUhc0ehq+rZ
0AIzsjr36QsttLqrNyYlFWIk0ke8IHHK6aW0xnJOIIbUuWg55zYgHKtyPsDDpMku
Be1/hgieXwoPl4rsjP5Z8LSTkr/0ByhbvWV3vSSCgL56JmG1AaQRt1ZC6Dw09H2A
HRfv+rs6v8/bXK43yXrYwqzMdUN5BoUsalprRqIQyuGXV3JiJJAKST4m+XFS5jR+
PqfsAU+JXNFrUjD0/lsjV9Usb3jWWFys444bnvBMWtZjeyPQVdAkk2RfpWmxefcs
p2DYWBNsE+RF1PIURHPAuMrhSSs6mTiM079aKoPuF5fP72Ida5z1+vZiZ4HIeeyN
byvft5RydRUZk2cQ2XeJpXPqpdkQMEB2cJcpZUiFZYuy9SHa8tLNNUup5GyUVgLz
zjFVzjwpu/D0cd+YBg0JSCH73DUTWY8zKFIMufi2O8LP65+soKYFPr+xiDaHUbPZ
M6k0imY0L9axE4tn3/6PGw==
`protect END_PROTECTED
