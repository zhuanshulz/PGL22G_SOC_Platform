`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bltcvrEq2vKFvao7zE07eYB9NQ5py1dkC/aXKylTwXmq4EtB6g4cbo7G9kJquaw
V4mCxQVIETG2pKntEZm4UXhlo3Bfm/rHqPkgqlFy3Wz5JzXeCoI/l5tQD1GIEtnn
HL6sDMTIgZLemtKmGKb5RNX15veL/c1ZDWq3VjYNfFArdXNM48u6T9jf0RQy00oV
Q6ZPLvoP2E8ZN7Q3Qyqb9tVVPfVlSuIJpJzY3tNBwCwqYr1EGhQbztlCSZ4KAoq/
Pe1gQWX2fokt8tEV67/aw64OQ5GmtYgh3I/FEqe39jBmy1gwQzCnEUDsLO/HUtgu
B07rP1B1YIZNUuBa0BKSN++GJ2inpJhJyUpuSdvAq+WhwLHq9lql103xcK0gsGy0
forYJV3+4PKeEVTu5S++r+Y4FUWaK49BqeAutrvVBmT1tjD0KwMvxVYjoWgyXpb/
K9tAhTEdvCBl1YBbiaYm7sDesRRb1StVPQ+tvy/X55DYFE8p4u9lvcecJcguhZxg
IXgWmZmB0e1ElUIuDOZKrvHKpEjWgxlZclrBh+MSkkAQWHXRAGRsh1Kho5kYUrvb
yvaprw1vlrYz7QppbFnZgsBqPPsxiTdaLsgmpCjJMvspizq2dN40zzxti7dBkR+a
RK82/QMCl0TxMNMTdKigudmWE8gW7vK9v8Ao48XCF8rsU7rS1UPH27GEjMMMZTjd
Hlx++7z0QtQ1UYliNVWvvlcwzLn2h+n/Ht1+MCkdzgCl5HQoUBW2CwiTCnDSo89m
P7Z++97GTJV85AO7d0hoMQITTRHE/iHoJcjrVbbDbi+jNRUjjIfuVJuhASMFJFIo
fqA1/P8ENhoYELhJUioMi+vbVMAa3dZDLa1BLlxQg/yly5JwQMnFwbyXR2qTy98U
j8qN5/nBoTarJ7ZJ78DZp4j9hQzeyxnMOQkbQYUbQ7VJ8UoYehx2UC6z3i6lgexp
hCGTUubzZj+BRStmb+bE9vggy8RCeBRgwSzduQB/qTRdR1GrhMVnH5Pd4PjQe72B
VhBXiFqhOkzNX5D57yk09zppINm0XD/8d1iAlImFdaT2etEhKKPwtGoHC7RfVlYk
ZG1NT3YQ6NtDlasZM/LwOFLejX1/6hYsdl6HT0zDJu2oOuS5EArp0Yss7oCcIyUj
s42ZMJPnOkSn844td9K7tJGHneXLxWzbproXdM9uOtB3zGVZmkhrkg258TZ2mA4X
GH3klhm/qtJM9oV6/r6aM4BGcHvyUzl+mEg1zj20t2YwIiyAIXOcD7Wul2plWtWz
eyaMnDgRxmU/xnf1bYrstRPCw9AC8Qe5vijSM8fXJx1nEADNn9I5AiYOZdIkzXqN
dMnGt7zep+bvMrj5763Vv88q2n8pWUHnSn4pcnWfZlVEuR5cxVrrtsDaHnim9sVn
xvwCh02Ldgu64hbiAZ0dirCUSNQ1xZfHIj2uHPt5YuJy82BKVHJa+fwtr8Zb5tRL
`protect END_PROTECTED
