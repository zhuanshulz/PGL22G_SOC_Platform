`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U8/0Z7ha2YvaEsO3ObqyS9WTqWRlf4PjW02JCH/pJ83BnqfJIpXLkRDMi+y/H3o7
yz7JaQQko5b5m+B2OWAFh2szeEOPYslc1YXPrDx3G2nMstiDEs1g0g6mV7lxraL7
HJR21s9mtaWi2qmWWYycFwDnYM8kuAlo9Gf+qVizL8VPzY7B1ah0p94f6grTDrFm
QOyauc+AwuRRezAPpmSOf6yeshATMRPa29QmisEkMyPVXjWD5Btjgz1DYKSJ/5Fd
v29mzayGRHJtA1rpYc8I6Hg02aWa+pVpQk481DWSm4S/yRQXW5BdDZQDaJCAWLO0
slZLrQ2tCeFdqFleqtJqAt/D27wdQbM3GQ7W+Pr1H3b1zytgRMLNR7foiu9jOa9i
csudxvEHS18x1EJpeYdjeCLM6Y6ZigGRRWW4yUAlIKKz9STgan5Uh9tYX6cWkJEY
fB9O6/6GM/clt2EgPCuD9eSsCxyGBTl5dSh1KnZ2yWsAZqcvkpUbGAYZkG2r/3Kz
Ha/L6P5iUT5z21gJbHpitTy7f812S5aP+n6xpQUKas5AsvT85knoH776hkg3+RuP
Z41/cpLzMjfkcIPb8oSM8jqW7QH1IVx4bPajOzVG4ghNbZZF7GlV01yw1gfbV1gY
sxe2w8Nd0OqnvB2B2yyhTL6LE97FKydw9tmSoimuDPYL/k8skvPVLnHveAzaGjHs
BIi8ewn8ZxKK+uMG1oQ4kJp0jyoAzVcf9ESdx7GL8BnimGJ1nwNLXK6t2nlkmpV1
xemJEyX28WrAZvkJg79Ti0foXJF2goKqGHo4XVymOXKZTwjeIL/D37+Z95H5dyLa
Guujwrjt23bJyOPSeDRAwj81rLLNE51nMWCSnEpWKrwtoPnR4jyNpFZRHlG/QchL
iee1EB4ShjxWgZkMTu8mA5/uSWvfqa6wKo6GVTZtqcw3Q05AEDWL+AvngqkM9C+5
sYK29x3E4qktPHTH4hyqF7bAzQO0xnajHCDAKM11o9V3o+mhMMWLCKg42wP519vF
o1Z+K64KiRuFE0LBUxZ3zp01JfeZJd2rUIKxYa2JAzQvKeoZcc4DHrhynhXAaR1l
M80SaVIt9rR2zdaG+Y1hdgFpKCH0Kblt1CrSCpHU8zDdUWBLStgD0blNRa86t3xs
YDbyETK43X414HL6cu5fovbxQSKLhfGdfBPwFqBvKJ5aknvG0ucsZlFP082RTWd+
lxCnHkipKPcdc94rFihsB6x2daRNcjxXtZvAcAkuv4I2ODSfER9NsdT/LGSNqD4b
3I6a268Q6LoD6e8J78KZ76P53rCsfFKenSCaVFFDKLA5H+oXjodO8FTWeSickws9
LEuI6gevlzd7gQdbTayCz+VFKBAButjl4mt5TFtWVYBp4xbwJab4ZTB1nsnAXErO
ZHzwHWXv9wEp6HQb0JHewV4lYnKDLaE6qxlQ50f1CWvr38GjrBi68H0Jyrn0VGfU
yt6XQZvU+K6u58135XZsagfWI2jJM68NDqlaSnyovpGl0thrCZn1eEibRdXnqY4G
gPuroJaflvGRXKCJa4gqhO2p4tWKwr9/fAzPyTaJevHoBinUcBXwq+K0MG83cIeP
En7sXAePFf3wq9SFKqetbE2W9xQLPhjyt+0+q9aK10/LfSsFgg1R7KlGCkija+ya
Rt4ZvsvM13U9mFQYZ2vup3/e/vV93tcoQWXemXfLM3kazYikz0wJq82H4WIpj37B
HEHSaTC5/k2O5Q2D/i1J8jnVReokOM6sJdYKE0N+qaRZwxwFyy0hK8zJGbc2mwWI
VxnsWtuQZTVgkjxj2TWs7qGwgE1F6paSYr+oS/uiF02em3zi2LmumsTEMLY9og7a
onqUoWtExJsYJe0sp/RPKjAffdcVtjHHiayo/5mjYlzJvPdtrbfukZUpd2uOgIDv
2/IUBBjfE1QM7LwRLdO9A9vvxaHZ5/8WPujzXzDo4llhCdONrSKDadoVzACEo+pE
RHC9z3xKhGmCKAJLATZK4MduKJAl/aXPDZ0zeFV3JWu8gpxE+LtJJCYDqXIqTVXu
GwdhBxl1jsojVk8oPkE0psgWrc/uId37ExQB//Uxb5+/R5tRWoay27tfWiQUZKF2
9rZz64zb2+irYXBpS8/CZ0rFKPdrOesgyNCdAOlOW0OE0ENW67JufRheElGGDRMt
KPJQ2c0Xfkwf+q+jrzaQP1LCZwRZmQMSGbi6Hz9Lk0JBksgSmJ8xQIa+Bg8nHKk8
1AbVgjpucLT6xiAaNcetHaglCjpUVqQFSh1jGxeFCNR4p2Eeob3xrx/jn7kJKtTe
l66uk0CpUY5v4uir7Bm92bwnWvneat2cN8+IItdS8YHlxKn6CEVjC1+4bk2p08ZM
hvymT5brITJdW3LxZkT7rPubpGQTLMNl4jEMd+UuRlL4KIKm8q91FFBHpQCGsLEe
1LUknOcJHJKyJRN3T4vdE4K4dw0HjaWYL65hUmKI2XkgufZi0N4bOvpUZqTd1HoT
FeXrWbfANov39VR1vtDpmS8JcpVMvz/HXynHb8beQuMNJpclpDPk7V9ZbWN/hcZ8
6B5Mk3YYTUHNkqOcOICcQT4OXkS0xCmQiYINB7lvzSZKc7i1I7bItFE/4fRcCdxd
24v6e+6AuHfGksbsrl7c+z4MfZm2xUirydV3EZ2Vm9H/6p5INun3K/eSf88gwstw
GpN4P2TlH+9AxfMkp4ZS8TMxjIHSfMPmrIUpBtCcJ3+CepODtTctE/ZLD74kBnpU
UB3s2v+FKB6rD9+glbsd62hWg7GBfxGv1mnpEqDJvtVHLSLsKVMulPq2OFOhndlP
ZEbL4rfL9m7bZkxfFzPcIgSXlDn3CycTcohK873Hv3N3mxvdBEqZhi1FERxPRP/m
UuioVwOMyCpoND4H02weWd5NQUEtvv32/tFCsox6AT9BoqAFcW74Tw//xyvpMPNy
ForZ6tjhpuD0/hsm44x8Aym/Jsq/XJ2N85bzdOH/E1bj4j12R+wdQQShg5NOtsL8
P5VIKW8FTTYAXXNbJttm0mGr+q22zV/6zwc1rY9pmkUhdf5J2/rB9nx8HwZ7F/7g
O94jEb3B7gGEnYsOevVbkZ9g81H8UD4DX4/uCoaOMFtYGZxCTyMfnqWgnV9Dslok
w8o8KdQ+SD/I8FxYi345zvN/C5lywSHGrJl4YgH+vxhFSQ7ypYm2lMROH1KiNggU
/ue6GecDHQ+dLyAzJHns0vaQphAKv/xBbyFsYrtubhHrp8OeiIT3Lh9lstfGjZ0E
8u/ziKrmkVRnJMk2RTWM/aYzDxCXbLQecZLF5LYH4/tTajFuexEmUNDy9I82KCN5
uXqTCMPnaup7mfLNDeqtzdB55tfFmJ+CLOvpbjTs3A0zQgtVHz8zBjmy49TjVqhn
+eS8sq8Q8PMCMGRrv/mTViDk9f7boPJofDHJduP4dc96iWxyaUDMysrogkm8bVDy
uwLtOV8JYkMLIrllQ5GiKRIaLNIQOtT2hX5Rvq1wIXpR8+S7dmi8JSvJiBZTED7+
+6Z1mmTo5YqNSjN8A5Q4kBpUvbGFdkRryNV3JAJNKY1WSxEOV6rZjg4+3VuEB0og
`protect END_PROTECTED
