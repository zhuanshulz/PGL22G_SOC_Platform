`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNxVMbNkPKJogMX3RPzMiOWyh1MDFr8/JfQgsaHOjUUSyIe/uHCf+auDHNZSUX+L
n64Y/Y5XWQhfBQjHcEXZez1V5aSBwyUkYP+iLVnyDzAd9cOeRBThZR/MAzxDjW3X
rwnoKZx2agMoiXu2eyfg/1ByTwUp43sdgT5WBjYLZWaiXS4wl5tVgmzP7ooukceN
h970O0hEGbEqHy9CcNh2ogWZ+kwm7GGmO7oTtvxGhbA9EFU3tb34rVzBUc6Gu5E7
XDhlM+97XjWg4DS9JvwHA+cf0sf1ffIwteKCTRd/GDSi4eOyFY0429Ll33YdoxDc
eEdgF0AneTszmDuS2eTzizOfwUgMinQhF8PqB3VnPJVjXMav/YzCgV+pGJFQnexO
A6Qa30SYgPxbw4E7gIw87u0biSKmnfd3nF6i4qvXJHo8ciYcQEpxa5QTfWcOHOWl
F+Xw9P2a/o5DcDlUC8rrAVxSU/phhEzdA8Xhnrx33yLonwhYZlrHnpv2+jq/ypKi
I6kR4OolFUBai/3xVe9W+1GIoYrJ8kcpxc4B79JuhIEIOf54SZWsQoUDli1q+VlA
gCWEeHYi/FWClgVh9c2fJp+qHa6WMw2K6dAHqFF7M5RrNY1atcQV8zyI64XB7Jxc
sL25Nc8nbELlTcky33p922wKNp/lJeuogsK69Hai8dwUmgdAE5pPy5QchGW8Kzf4
+qU9NfjhWlQK0VflITY7YaENz4em7XYkOikmJfdG8aoScYOToO10Nzz4sz/uf5ZI
Re1Vki6BT3EV8rz2BDvHpg4o23rD+7vv7fjlCO0AX6nod06DNd0+Fif9qs3k3Wmg
7H4nqOn1Dt6ylCcSWQOFVxX5XvDT6MmDpR72nM2F3scSoMe1vzjn3GXU4Tpt+Xjz
ErCapOsEBOrzD1/W8nD5hvinAaUj8afCIqHgwR+CsGUDyTOsYuJ8B4MtiI9LcXeA
gU54AZ2zDsYS2GiAw41Dro5dypSVSjnNGMUht5S8ltFzlkkSEy8j1k7vo8VuvFUp
RuYwI0HR7dJgM+YsdT8qHEUhwFxwuK2pzyhgZdtH8Kb/J0u3qW0vDoSJrQAksYLe
6gJN+WO2bMoFju469dvKBHFW95UxCzWiyiXc2ahENVdIT5bF1+wvk2jC1tLsuaJk
c2VWNhLojnYamMDhQjoxxC616bs8M8jEo9WmcbekNjL3L1VQjMo+g+edec/VMYze
/kp2cWNZFuja+ZsIDF9MR2f9G2SECLwNrZdat21MvakwKqqV0PW03cZYNK7oyIwN
3ewMCYjaRioHz5uznhHgmTKQVde/6TJq6yxTwleY+//f18ovvDDnpPZTiSh55aHt
T6EZr4hyczaQJBpbNHU0Dm6/k/s13B4x877v0hwD5Bc43LaiLEMTHRuP6dUkYg44
0KMJLkd+gpmHn/CopFP06w+sllueWkB1HFauw2axLBUEFr91ZZgL/Xy6/BmQ+34D
78KtuZ3tUHhEDkCwQhs99Feq2NdKtBWv1bZ7z6dk0QlApyfYzP3REX04b7OSvJxR
roulfGkk70NWo19EO2I7NyNOcS9zrWh6SSlnCa0G/S1x74a4xKvDca36XYjY8jJD
V/qvbCCD+3aaweDIa7HnKS5GwSq4zry8vN03y0Q/5e/zDg4CCudd3gJjM/a8bGNz
G68T8+aJH/GGmTpB137yGw==
`protect END_PROTECTED
