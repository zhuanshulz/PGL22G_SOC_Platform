`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ugXKTgPXLA6NWGX2bSdwGgNTgo2ltOasIi0jAJI14IAwDfflHxm1w8MmvkILLBSh
S0j06Umk1VUgtzGON7N7SI54RxBc7ICLhLr1A1oMknE/AdoOOGhu0BXKWWkEABWE
lj2ka2k2q2mm/CuP2YV2eA72txhkXK8j2OnzZ0y9m3DfI22VRqxN5vgQ+TdGIVq7
Lhczh7spA17XjwFWQfBXstJZxdXcyw79Z+OSsJOOWM2upXuBxvgei3ZEdo7fuXIj
Vaf9eYrqNCeHDoHkKiSisjPhubAw9tdswNZgvyZK5rAnJnUU1FNMxWAUCNUV8QgQ
76zUW5VWOCq67RdwBm3lRpCO4ZkaTME0A00OHIIxp3wFd5Y3uxZRf1r3zw5HkdN4
/cnfZIM0/phL7/rgGiWe1LfYt/EUWHd+U4Fkz6ugJdZVPyx22t9g0jnOr/XwH5Fb
8i+nFsZuaia51FR7hMyvepIDPa9iB2RGt/fco0iAQQ2+ssd9rhKpZ3q4/DM7NEst
cSCb+sCgYAmu878lgbexfoXo88eIqm3ZtnHWubDEZJlEc5C46AbdGpkbRmybYhlw
tAnnrYzxLhZD6hK3gfdrJechIocWKxpx7ipaWjpkQunwS4X8SFMRcRObH+7UZej1
XIzcMKdTxhU2Y2Gff5gEhCFSuBy3M8bqLLyODpRjBMaMhFLetjI14/tTz3BvpxHg
WFvQbYY9BtBbzAD+LamstBy23Rs8lJNy2ocqefkpesyBTUnBIWGM8jfpSmP87U95
0G2qayVEKBlkpDQjIxzW2j21mK6UMwWOErTxrj7uURFvLrpSji1mCcc/wLFa5XhW
O9O5B67iXuSR7Z3fBC5QhJ1Wial4asAwtnf8mdcJte8zqSkXjoBV01GFHw2Ltc0D
TTcHd1zRAV3jgvYXWnonylOyKaJGb9rNyxdjeHVq21x9ja8/q1z8JSa9Ftf6SNLn
M6qmKEU+dD66mPgnT0Q+E+1DHJ8vR0HJHo8sO4gVB0OowJdTiGp8c+vqHlfHe7dz
LZQ1SltDRG1ritJJpxIBXPCw57HPrD9UnNLUGHlZyLUjjMeEaBwbZERamNqigBeg
RXf5e81hfT/FbtGQDXQTQPGhewpnSdoJPVge0OM2kMQL1Rgo8Od8GAhN+5aJOKus
/7yzGJbCBrySsG00ABe3FUVUVRUy5AYzLLz/Ox26ij6cVcn0YU6Wa1MOVnI6QT+U
P50niPQC3WlM1RJL/w2T2xBfou8y0sl4IzQjcVwfC+qW3ANOqE7P4hu/hflBv8KT
XPVxOmxmWTaqUJeJu5xsJPYj0Yal3t2/u1wxgAVoqPs5pw6Ge39viqcTQWfI9eMH
`protect END_PROTECTED
