`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldSunBzbtZoiMiMNjpFLeZruipQA2TXPNRoqhQypxWypWz84V4/73k5cDWmJo7V2
7yQZj35kl7XGt/Kwas6UZvxjS7noy5k6sBrB5rsno7vmVeS1KCHKLmxufmJxa6fX
4q+3V+WOrCVLZq+Enqh9mQ==
`protect END_PROTECTED
