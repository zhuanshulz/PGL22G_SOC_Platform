`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d3UH1er2sSHpq/uCZZaiEGRYxP8PHG5MeMx2sonjPf3bi4VgKtGoBCcYE90ECr7V
Y9kK9rN39/73yv1MSB4hUWB/RbONiPFaBlpd0L/e/gR/kDFtj/Ktzwy9xNrkE4BB
knYOICPudVCZoO9kbKC5cz4RkBdKDdpDXL4kiCf67HpHkqNjLN9B3jxGq/pUDXsw
RuEtPipe5akRonNLaniOn+s5heqz/XT9Gu0GRgXH1lCUrQnCCXGrclDQFNyVifls
lzFgJ9yJY5TD24RqriK+B75LNsnqvwWfGL+Z/K/e7drL5ufpUI5P+8p88A0pLpmc
YSNV0HER1teyqagrDaVHrBFgTcBR/XM+QPmLJ5VfBoOBPSVO8mSXPMAx2PNYGHHy
ppCzig5WkC3O6+FikoNX3ij5380f1A4BIyXtLKpiSyc7MLoSxjaOVeqAdfTkuzt0
2PjQysXg4cCkpxl+wJNLWdvytl0gDmb2DsN4g7c3TRAycvGINZ78D8dt9XK+ST05
LKmrgThCTy00NFG3UFw9sxqijnx5Sb2WpzC5Kh1x2Z4=
`protect END_PROTECTED
