`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fiHMVgw3IaTlkF2dt6bbUuC77gtakMBzK+VCbSdoUnD666tICda4hijrnRc8uskD
u2HA95lVhzB3zrZBSZKG1usvsYJmMbOKeKCi/LV21+8W3XoIL1ycime2SpRW9dTp
y4S7/NuZF8dPg2Y6yr9qEDm+P4KpG1cEm9ifE7G86V56xCgR9sKh/spgYVdbiCBK
pLSOOwjxMWr6lHIHT5p3Quv/HoceRcYl4ZljW5BYhZmH1NjoOStJivU3sX+1USHx
ubmaRra4kngziVvKJC6iAI/8Ow4HTWIZeMqAiaZ6BUh3U2KR7rk6ZAckeyFyKJlb
qPBR5+ZmQSM/YrX5HNqgX0pS82HJYsY88Li7YcQFNTPJEa1HV/+9adOECcI6ImS9
qyLQkJzOk8VeYhQai9IoqA==
`protect END_PROTECTED
