`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J51Vnskms9TikdNxKn49eUUiJiunZkSPDwpiwwHWKpXWsWJzu6wtDmppQYRwjFuz
iZZezZcAQHukTfAqbXy+5Pw3aK17l6zNAXRBTSewNbSeGtuy3FkTTtfn8MaI2xQc
TjRBlNJPe9FF4ByvOUWVTT3r6KjVLjhfSRXnLg57UHoDgQCCbbylFG2eRMLPE6Fc
DMvBPy2BmxrocPBYbVnykTieu40J2GGtZ2KIUiJ9EvohxZ3sCtx2wb7xT8gOjPcN
ZdkcbTI+rwT8C7F91qThPe0CppKEcMViK0kxM2EmwuvPGwfcxotZQyVL8rQ+gxTA
f/oWLcplWl9JmX9KxvR7CjOMUhq/8YyqX44fGJARdt9UneTnZM51ZYuj3zwpPGQ1
K4LRmN/xd2WTe5xjZWEp/Qr7YtSaUSi4FIuSV5RX5vyE46GTafU30Qqf5x4T0scU
U9t2YH5mvOb08Q1sEJRKjQ4iOGHkGt2flGsMHZRRahyUhR3VWswD2GGeCsL1TuRu
4soVNEhVuDZtHseHp/p+p5KWi7j2RGXK4ClJw7oyrD5/ai6nIJRQuwYJybU3CTwM
z0kaq9dtSVl7qOMfrgzwEe/FIrbTNRjZVVXIu7Bdgf7NeEeaBuUDXYrVZIa3Jdr2
wCcL3V/E0CJQVt+0veTNlsfvak8JtcxtVKpo0+ct6tZcFv7QyJApE105DOQg78cd
IxD2GWQITjInG+9vEmd/T7QNgahUmmoUHXe9eoBa6GTy5RhysDHxC6Ymiyp2Yt/y
9S+HbXDligDq4r1mKSlfRlqFZr0dRc/jPksE47CYnGjED8ofCoUKSEHaYLQehL+m
CE+sG+0EUHrh+YxalUV7F3/tmLPloZLzO/A74hO79lk=
`protect END_PROTECTED
