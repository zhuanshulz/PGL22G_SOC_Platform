`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eDFu5IHAVXMf8d3jpOoltB4XazyIoeJLZ2WKYiY8ZVTmPeqyKIDnPN8PWN7kjz4E
nnVmf4Q3Z8If4VFNJkDeMjuSuuP4qihm6rkCsHiiIitb9xDekXjO+wlVK6cOaRO5
bxpJkwtSBCN7QPADq47MwqSiMiIN6tjT99oDZtwNw2e4zWMRZdhHdlm7zTV6I82D
GhnFoU/ZsNZdDxSYuT6GdxcANC2Zuq3cw2LG+Ngi/2Wf54gmapWvhKvxv3qPYHKC
Smqq2x3zGHWu9Zz1dge4o0k2z0rUmc4L71V6I+0R3ErmCUWWwV8re0VYCJexTnHS
7FR+nNFZLnAS7S0dBR4M2ED7MVYPFoaHlJbibt8c2qSaJgOef4cPi0qooZOb8d7n
qQKsTTBq7j2R0Pssp+7Z6P2xfv0bx4kIUWtBT2ZvbIejsP/VJFSBY7GgXUKi0uBh
mjr0K7CswWw+bqQv5dapuVVcSaDiLmcEiicVvWYHVCtyK0o9WQAOB0otTQ3ldcMt
EubXgGdSUJx/zbO2gyIbIYKNdKnf+qYtfiVlEfw7DAKd0MgSXEPX2MBj9XaA878w
69VbtB0L2X5qX7GCrM7C5YdXiXo4iZwIqzmf5vrNXjJpCisVVWsnFbWYy08btZxI
`protect END_PROTECTED
