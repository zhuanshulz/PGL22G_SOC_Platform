`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IlUuv9Hh6awo+n9IhF5AmM6PyIToJUboj+o/Dda+O0IiJhfCyunR2FrofKbD3vt4
PliJ/b7mClvs+ZaK3A2n8cWqLHUzs3Qt/yxqf2UhU6ggw0aj5ueH0j94rLd4Ie6r
giZEX9f3Iez6Uf+xNMcY05ibrhNg1WusP9NemqfC6VtWjfY/iT4HGdAwEwkjlQ1R
p2g7Ht/5GBjExLVokvGplZMf20qUp4GcgSG5LN8va94vldBU2dLL39jPHOTZKExL
P2zoHEz6IVYRF/UZKGgz7N0/TZatezDS37I5mbn2CtS/MdQDkIcwMU5LEBgzSzmB
or7hgPUVPxDxjX+kPbjMdFE8lvpcLs/0lAyEom+mJsQiZzln7ilyxlu1muP5c9ep
4GCNDl9xr8OdJtvaSQuAwDYGfR2LkJHGe2Ueo6js8vXHXYDbf0eIDZUncOlOcxR6
HLnGfXToh5qbKwSIgMjdR6WFOLDodTlbuTWi5cJrnqRKObI+J721zB7geJj/h37u
zgbXwKJ4nS+bLq8btfgUBMu84AOTnM2iDQq7nM5y1+X1BUIMhVr9NiEyAFslTFz4
Q28mMXhe1EKtZuJwEwrZ4A==
`protect END_PROTECTED
