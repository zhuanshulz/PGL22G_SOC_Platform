`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ZKqwv13HaolSXulesy30vP20mEw3xP+9SuEAp0MacVRB1AAv/EHvbEJ2wjZC7xI
FM42VBbaVX6DV1X7O+fNVfKTzpC84f74b1vCm3UNb/wFYCkZLoDZxpfjWGROOXqV
pHWH0yIYVFzcEfPVWmoh+lkST8JeVoaXN3zMW9s2RqlMbw2x0VgNLiPQRyOB/214
Duz/En3pYrMTJum+YlLtQeM3nOHQt/Bm793PtQSDEOk04YmnHu19ZeIaavAVCHO4
m8BizLf3vXO9AJJyRnHrmQA8dOZDpbP/31k5uN0/oAiAPkEUjSWFpuSMu/g+Q1oF
eY1kaUFL6xjJvU9BjR/JIxNGXVVz9XTzZ8QdZlZCwnSl0Vc3liLRSxrCDnZiZCGl
oFio3b3OBLIpU8iz1n4iXGPCxM1qRzmQxi1h001wlLf4O14M3FYZCh92DuwC/eJw
st6W6y+6WyRUyVET9QMMgGQXlSF4Iqu1Uh5bf+uVTiuxivlY5encXfYJGw1+LFjA
aEaWTmokM22yg/SVrai9utEDFTw0wndn9rg6VzlZ9EI6TurNhIfIi+AbPJo5CBap
wuUTbYTKUI7eBFAT3WIBRNG6tUcIFGi/Up1c+W/ibo1hcZz+NScPVp3i+feHCXKd
lw4qhkx/hhTurAg53m+XekFK2PXVall6mhY/lKKT95xjCBkjEih5CT02ABTyf1JK
NOkeM+HuEQYXmx/DVxQliBi63GZYE7LT29OvtJKj4yuhuFJ4GMSGyD2ZPnADBRYb
7HE7+URcsjzt7aCNnDuYgYZTCe8TxjprQCgir55dXcaoT+2t3/uBZf8UN/nus73R
9ZeTOaE4gUFPKBryJmiEfDwGveUxWfj7Pmecge2EY3E=
`protect END_PROTECTED
