`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L/xOyBWWnirl+i24D9lQzwxX6Giq6okTHkg/Sfyyp0aGLFvaMp8v8UzTbAi7z0q3
i/ksHsgxldVm5XluCrChZM7E4XLR795Bngldu6iPVd82FxgbQCftVj/i4HdLJ9SD
iUKu2pmTyu/H4F8OnTW10vnZ/EDW7UgMOMAFv2K4Z/b7G2xQBDdfShWn2cO6IgXo
4f2cJOjjfq8U6L9o+ZSOHsX6H+NrXU/Gi2pVpWC9wsVDCV+2vPLKQYTHPMvfD+iC
muTOyObSNNpExY6SQkauHhvTRARe2KcRrmJh3C7TfjjAbPsnrFYeRhPA7myXQX1y
TXUa2b+1H/gy7brpXkj8vClSaNWEQfam99N5Vqrs4c7uYOyXQl4ZlIkGb/kxFihw
BOo/5y/VtJYOp6BB32l5nXOBEiwg8mAxw7rE1AfrQh0axd2pgYhDDQSYvT19BguC
Zl4PdPg7u471eq/Nrg93/Pzs4nQ+s8Bo+ke5G5WAys6jx391lrrKt2l3Ifr7zfG8
L/wK621LRBLejirobd7gFEHhVUG9/nBFA/TwFOGp5qSyhsoyh2pymsfdHKlEAppr
FaA+NrwjeR69Opbe+Fl1adY1VcCR440tT+ompwUNnEuwvMwbQlqM28TanvOQaHnZ
5ltTfvwcVRH+lRYHPT1kWjmS9lB/Af4xR8oy2WIxLIXwunxbECFeC/r8nUOHyU1k
c/mRlB0fuq3nBKfG8VCu//s1IF7qj5HYzUXeW1AjNeUrA+xGnXj/SgVp9r6VT+qR
35Y00YL88r4nQ4kn2ltVUeMIj1R5MTgF6qJ/X5uMv58ygo7og3VA2T88zvn1X5jd
wwJzwOtq4KwwJ/4ikOm+g7KmUJelJRBLKwTfUUKEHEayWKbqzY8Vq7+reCp3QAtG
hXQu+hSflERWNDRTOhPNKc0D661GnCbfGRNknmtksU86G5BKR8155766o6DluYG1
ABN1dtcJjV2sjCom3Rr0LUsGXPjDclqtk838oPfs+9MCPe0zWqbIji+Su+0pvTyu
KwuNEwoJ/T5F0l668NoU9vvW8I1juBdkE5xPQsMShps5C1UOI3Lm6ADPC6nh0Eng
D7l3rmPVbGQ2YwGYq8brLaIcP0zkqVgdZZnEts5oywBI79JeMCbZs0Q3DY11bXzQ
BBWUa8JsmBr7NcpG+dIcIBT3SecmSDNVCuKRn7LkA2BzhLSQKmNwAJiUHONMh0xn
4r4F4NXT/aISVuDfBYS/ki6vw8NHqILATWk/YW3Fydrpx2VsyEAvuQ2g4vMDjTJn
mTHfjl1//5OLewIuVaZBVPKA1W9gRGYOsP939CdrKPwolW81swIFeRhQOU4CfpVk
KJnMZZpUlW0Z6apTC8FnKru4E8FEx8xlDliVmgzkj75XSNLJpknAk8tIJ86OdFfA
dU0EWL/b30je+R0VxBwgLxBvY6XfD0iYEaVKVKhAHNdZLTrZqpMa60gm924+lRAS
USk6tEHyghhU0x0KQ275o+pD2AzenCyWOMcn8VSUhY+GYIrharlwf5/76luPLwPv
Ps2mjDenDwMIVvWrSaZ4IaIqCfgnk1GRxP83Nc5BfEhF8ZU7UnSTUhYGx3wsDcll
j/QLk1IXgJsqBvIVJTD4rP+eU2FIf1+IUfAHwTe5x0VrqFA6zmCtiAHglYw91y+A
QWRqG6czahSWw3KC/EuhkFyWU46GttecSetWAdVabv9vKqJJD9XotPmu4+sV963u
jUDT1x0O30rLydL/8tgSkylHOlXqK/V7GdWwpI0ScCm5pygIpB03PCMW8GGeHXRl
niF6c00Ox/3j2nBLparGbS3YwnvgLT9cVa19VOe13DDz4PrTwToYuzyV4f9u6Grc
gP59ZGtr3VnnQlNaM1SsEerqIFXaUUvbZB6pO0/3u9uEh2lz0ZswJjR+JtQQO/Pb
jZeiw4hLfSEbmSskRx80re/3csR2c4BuKfg9X7JTW3XVFyB4BapOSbQ970J6AoGq
yGj0QYnzjpSByeZ91U6J+WyvOQXBI1mhWiYSceTS6feEysm93bE9yfWaDVaQP4bX
QyYiSbTUNrGnvHyQafEtw/TZ5XJMfuKYGDLuOkD8dkyI9xYOb+vNyOZVn8RuKnnO
jUEWDabBU9moZQI4e/lwfTAy+0Gr/Jo+ZyPPpWhBkcv+2vsTJofwim2y8YmuOMeI
F/lyIG9zqZoSANqrmO8LzwIzilIJx7Pz4rQywFX7exG9Polhg8laSeP23nL1oKAx
clv5j2Z79xFzNt/s5aNxTvWr7oX+XZzVb0bls9mNLh0t1SJMCxORfmzoOEeCs/Qc
bbH/OJ68IMNLMk4Exq1xekPNZjJhIEjqWJieSHOB6zhKqPAkOSikzCKfMY9Ch8iG
/0MhbC6g7q5LTPhHJJa97vyZ48YsfA8CuOuy3b3zpnQpFSgfP+fkhQUhKnqXsI+h
oq1734vHe3wYWLt0T5bq/w05+Gnql3RPahuDYwTlzFrfJLIw3yyo/pVAYaSRXZxX
BCyj5v1SfPghTZJAs1cxOFKrjHuIWaAKcZyTIW3qgLRj40lxN6WI+Oe2buJ+kmYG
KsR3HxVoiJw1nCmm9REoeyURMvn1v7CpTPPEUbuAXf3Le4RwzM2tPDBmF/Hemhki
nKI+DozYQy1BpEGsw5snZ4+Ez96sWvOHoB8asWtRQa6yn1e1vxocOKxfuqDa9+Rn
8y+pSObRELaxXrl6Q7ZFGKuM4I+ZDhtDVHRJQtb7HTlSoyZccrcUYmd4InFGc8j6
EWXPcI0+m0Qi9aeQncHUdQpeGYROj2gEy/RRzMI34rWN1L5G/nyLO/KrI3wAUJKZ
EUUFpv+KFp4hEmsmO3yDbVo7ZmD1vRr4qIeoDinT/QHfgxXO/g2FyB95lQPQ8HUI
4E2U8OksREO3AIWxnEdVk+yise5dbzHvvbZ1FO3aAt5BsTpXhLPbWVzFwAzaZkAY
vCQqS1ixjkpceoGf3jO5tlsaCkojcPAXOfcelO6GR5dsANEeQtUDW3qyLQSyqztf
awPujaN8UkZ+2Vw4SNKDugPCOJw/QrIpTsqFnRLwI5/nZDl7UEp99KvGZMSsfpDr
Gq5iVHNpEVTbPrJgXqQ2En/yZh1zW2f/4rOz38HwrSHGmNt18WoV+dLMxZZbIaW9
6PJ44M/1ruW8+O/dMVX5nKeNv8O7+SngH3GxookNSFiCM8iI7mhAVLBAQjABgFp/
qXVirBaF0ME1y1p3+eVj+VUZr4j1ur5bgK/X3B+BqxCjxj22PtNk/Tw+gQQu/A/z
yVgjdSAXn0o8JqSk4RyapduFS1y1sCEyWZ3URKtQX0STVv2a6BNtGwn0ayIibDp4
g7l/5kLa68laVbm0h+ollCq3s8hpiQMFjLm5kX4q3P8KIcwD0zj/uJcyP+hmoazo
nTduZLStt1Q6S9jw/EKEuCYx9hg8weZy+jbNIsLu/BHVPXW/4qsbLA+fSAvkDBSZ
WE7oXIidoZECu+4IPNwDJEQz7NvZWqglwCFBWbcge/LFqpxO8tQgS0JuDW0R6twJ
t3vsu5UQ/2AodEPi8YF17PwLmUe0XeeuV3a7dlfOVafe0Xep3/wBwhMNOWnETThO
n7zZDQI59YGlM+qAz2hTHwcd7VQiXawbzwJdto15b4qL0cm29N8irC8Dfi7TeBBb
01yP5e/VeTaU1RnEvFReaIKJi+iMBNGXuzM3jFBk0Vctmbfvx3/v7haBA5+0qQfJ
YqGZWJjmYGFH8OgEX0qdxK8knAZbYDI0kMdm++S2fuFuA3qUqCU08yRKEhOgzBSf
1M4c1F93agvaQ4pkEgPn5BpY6ihn2Av2UQ6wDyUil+ozi2MxqIjjF43zFHqUhWwr
L9hnFdz6S7Kog60pxjcF5DpGdRBtiQjNsM0Fk9sWS1pF6Ezf1BRdhmGsXRa4exvs
OP8+kUqRDwlibSYOTV8ZDgSL6K8IEhCby+1YxR2oFJi7w66uGQ4Ru/vPhgxt6vLM
LgxgyDyfx8+nRqIsFOnnHxXNu8yzRxbvE0L/aKRk1unvhyXFXIXZOCm7BW2gzOuI
dXyNU0ZoorDyHN32aSy6qUTU+PnWsgVX1+n4P5aCsvnjaZAYFSWU7WkYin0iCtyQ
6n0iA2JGSP0SgSZBSF37wxnXnVU1t9G3x0ZTUxZyQxL1tEDYXRP9UspEA9H+NxFB
gpUQXaI1umpPs0bJDIJSV+6hbOMAlIjQWQbOSh1aKP16M3k0Boh2zX8o7vXmOwit
F988Pvv3lrXW85l1GowsLO8Koha68k/BtxRhqn1dJcoSAc0jV5nwDWaSKmQygV35
wO2764FnBVhQSLkNB3Js9th0LQeyvHowd9ew+9cf/1M=
`protect END_PROTECTED
