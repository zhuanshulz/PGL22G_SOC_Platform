`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnwrUeB1SFuCGTtGB17ate7zFYkq9dvFEvJkZxMdY5W4X4F8EWn7UxKm09Hcud70
acuAixMnYy34fbQLb2W3mXzyKLQHzIIbjTRWk9i740Nth0OCG6DJwxsQr4hbGFXb
VspNL+vhvjZ9DQvamPY9QgX/4wH2Tzubrp9j3aSAfONNggu2qmcxCTo0YuhE6L3l
I9qFnKL1SBPkJ4sYCKADgf1jlOpm3bUKqjMyxzYL/S3ZvxqpjKkX6fvpKITY9A54
f+F7ZcxSCFYiHchyX5GDbGORQdzWVkLWyMiizzuTTJ1FjXSLJYJw6SlPrgVw+HH1
zWA66UHN9XRcT6o/t9ivjk7u14R6jV67M/ONcquUK9yXqtRPk9Wq1BuRvwHW6/N+
0AY+/P6zwSVOJPXhdutSKsUZ3ilo4eIxmLbKAbZ7j/U0mQWrEqCYJHmTu2HD2xKD
SCgXRhFWPBr/IqMAjj5phvGrcxca+DrMJRZTRVgkeWNdIL2bOJyKnPSli4AzYhn8
3oamJh3XfmfdJnFT1omXkK/xY0IISMSCeb4y1husnigAfEkN1DKnpff9u+D61acC
3F9+OHIuGhKIbOI5YpB0qUn/Ndr7oYqFsGMi7us2ccfF2b4t98jt2kB7Zha3kwXO
`protect END_PROTECTED
