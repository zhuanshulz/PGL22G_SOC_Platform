`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKnj+MRIS64hBbeeKvV3xCMr2j5WdNtkX08iUbqeNDTjKikop5/mCgQ0XdR+25RJ
lrdhO7iQf3zwzGpz64T9zOtZWGXnOo9Xjc2tzWFmfjoHUjjN1Dwv7K8Far1z+qG2
miAYMAWikDb7vBDMpmExdnY8auD2j3lDaF4D3I7yVpyupalVd+6LUL4FyecWa1ar
cajDrw1bElb4n339fibIOab/oS1eng5AWy7gFnyNvhM13ZewwkV58BAghgsfYyZ5
eFqEfkqJy5JPhM5sWxGQF8rT8bYo9w0OBQ8GPv1TT8vyn9+l9IMoPkoSbnNh/CKD
QEK9TfQR71VFmX7vBI+bYDzhJuzS4lBzLxErM78TbJsqy/8qh2qqCIB/fdEVgWlB
wJ4gzxR3I8/nGPan4nS8n3zkDsUvLR+AcIyGEcm0whWfVewhVZKCDKXJvwqTjL2s
aFWeXWPxA2Je1nmWQlyNAHj1y2Usw2YsQFse4aADEZ/T9iHIP7+UK36OwTbC6/fT
bQOI0YI3yQMdUwBwyZsQEwrycsgWjNtnTICNPWHYwiiW6Kc5Lnxl2IuAACHD3CV9
psrLqhvZ6zifKqyqr3FmQNM3EvIrtMbJZltcjAa+b6Bl9l8ecwMVzE3eJlqCtWin
/yY+4aXPLQeX7oaGmeXccFtALN6khiJG8G+BQibee7DbsbufDYQjKzO/FFNWNKaS
V2YbG1THTUxh88hIpUyEgp0e+KyRyX2ydPnFT2YQ16bOSt7fMmwzCCLt5cv8VsUX
4u7N7WdsWcE0yQpN6eYvypuKcDVx6GUEdovTKWBj7wnuYbJlVeYOyaBtaicctfg0
cLBLBFiPRw6QXWKB8H8Aatm8MlOrSaOkHtC8MsYdXwRx+De784TT5Mc9eFkOYB6H
WYpOXKskr9uzRuExuVInGFcJSx5wqKrPpy9usOox7DESsS+nx4/dt8lrWUhyGKOb
KfYxT2oN+X6sGsCepWWekLqmc4fYKVi9yd1SZMrYDCEIp95QiFsrXuaoi0P6n5F+
FwFnYS5ckTOt7150mRbYgcus8+0gcogLuSQxlWFjstWjiYYK1xSH1ssMmDO+I0Bs
f5HgWzrBFBqZXYYcKExM7moPwszG7xjoP28RYaRCVikwyOPqFJWKFKTNov2Nekt7
jDTwzRMxOrNGSRoNNR1UBLQ40TWnRhBqROdxVR5szNMD8ysi+f65ONilnZ/kaoCi
LuUz0l7VRT5fUBZ5qYqCB2xOJ/frwYeTWgpGJ8nha9VTMjJTAOJqBkLWVGnX+dZy
1HitORRmG8iwdxvw9+zVDLGrgiQqOhUp4JjgaiPMnjDZhK2LNUTTpkLA2oX4zR/n
eKo2zfdBxLDjg734FpYyPJCOYdD+dgI6IadEaiGLqj7f1T2sYzaJEz8gDQ2T6/WT
XaxFcr+ZLbS7OhExp3DO5jJdoM+2mMJcCVKu4BxH275q8l6htCPs7QS30Bv5aqds
UCLwtNrb9lVWw1QWFi26bcR8DRi5jol2jM7NJIlm6/YiFK89lwDy5syI1jThoNer
cD1jIRrWvglTW33u5KvZffyd+t/4HZagkYULE09RYYRu9aEr5SXIMoGLgsQ0940I
TscIZFkpq9g1ITPvrypM03RPvrJFx7lYYVXSOoAg8JcYfXJaTRLyWVMcNUCnpaVQ
1oaIfFSBKxS+Yoq7Bknd6EleZBgNceD+So+OYWOEjHaiw64LkkOalDDROEO8ZQf+
8Xh+QODH4+1CoDS2pWbtvreWR0/652hv7uSC76p9MYvjDWziDB2ym9tscMvB8mjC
ThxCwzaEvvLp1vq5frI/SGtzWG1aLOrgkX/9MqKVpONOthfFQaTTPHOPQz57FByj
EjDiUr/6X7QFhVbyKqws1O1gKaXKJqeh9zy1NEX6ShkXqzK3J5lwRh+2Y/9AWliH
DMGQ2FVQhUpaoXzBz8se6YYY88v8UVeO8a/RxFXfxdyCz1CBvbq1Ww5lq9TqTKl6
kKF+20Htj3gAGgIaZ9W3n2LEYTLxwMWgCjHhhrDBETu+6x85b2oFIFPbSX4mp4LD
AmklkK1JrJNzb28EERArM/AlBCrdFGGVORcqbt4cZa21kQKKgQRnjMoBf8x+k9X3
BEMEsgVDXPbMvgQNnbwG0xe3KSLlPX+ASX9IIdjWgJhc4AYZQ45q6wbMW7RcsDG2
Lu0OGS4dvX61dRwZPVlrfWnox9l4LMcH2ZbLrZCc6GgT0+tZNSb/e4jAfiYIieVn
Mh63M57+J9/QHUSTjeAFgUUqjfPBjF2SWS40fh7jHY1ehX/x3V905obqMuB70NBz
wydmRTWkzlmudBVEou42McAf9/SX+aBdfshSCe4PQijIgQwWk6Txj/CayoqFHvWA
YalIMAyZtLo3Tk+gGWbY38yB5Dih3GfnNhau4Oo9j6v4TbCYRUGLb2UHFoP1MXRh
K/oI9VRl1PbVuhRhYOEe52+WylFgHDzUF0Kuq1bEdDbkKAclnrvZxAk4864NrS5E
IDhyuu/b8tOCW5AeDT36qEyTeX5kC7UQGrv2cLWhvcyvq06Y53A/BZEEXyYiaKKX
BhfyGrdS4kh/zLzBe7HzBcCTyH7RZ97rm5PEtVya3l2ocwSCpfs7XqfTEmQbAqT/
vt+O8O4CJ9vYTvsBAmHHjTlevpUOha+EW/lK+wpq/dqJFzfBjDrx2y/3FmBg75c/
2h0zlCobWpeYNEZaq8ahAP4pRJWppeScFdKwmItWNg7FxZz4wxWd/n9J5mc8iH6m
CRgtuvETacW0UQ6tZnPOfPfsBOFo2fArnE7CFvgp7yI6tO9FBsw2fbV2vNbR1e5F
`protect END_PROTECTED
