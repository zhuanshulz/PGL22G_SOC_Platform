`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftkRb3qAHf8pnlHOmjs7Gee4ReLIATrjM9mhshF4HfX1eokFVk6HIyluKQPOULhc
RNd48A4o6kjaNBRIJ1/jBDkS9Z31/oraU5Vizcae5z5s6BJ2FLeaL+snu2LfIL0s
3FLRoU2lQwGj3n2JdO20CeSMBxgl/1JWgkP+lq9vmXQFjqYK/Kk8ddRw5gZZw4SY
fPzkYshzWUL8CSzIrevIesOq5DmC5WHX1GCm66weEg0a3iWW4vL0jeBq0y8Eo1Wp
HGiompY1kQeY+1rJWmh6OlIkIndDf+i15zo1k2Vz8HrCzWuQhOob0U82ts05Md/D
qhEbx5wv9XVzncyZByh1Z4gtzoFgBGDBkmKmCPGh33GK5+9CIfKVmzlA08JUodpP
Z61RmOtRIjO9/tMFdcPmHTL9P5qBOXTfSe0MI2shv/17XseJp0d95FX3y/j8hihZ
3BhHtzqmNTTi8k7OIhNz9S6mu6qoCSGJWNz7U71htPG5PdvmEMX32GzVXdcRX2u4
B6D4poIMN2UQd66DrZjIc8RhVJ9ezXrMx4/SEyHVhPLhLh+P0ejk0mqMT0LJTEap
CdCdzCBa7wIH7rTjCt1wp24lqqmbLqoC13GPeMHoHvxuffxCOV64sXC1sgsCoBgK
jRm+TsIdnEP/6evrq+3uVWzFvZAg9XegtwjUisBu6G7Wv16gClWpDYafySk1p2CN
CHO7gK8Cn8sFeSpHzadlVTc6JsrdKBfHV4v7Pewe4wpi7zGZqd/dXXZogD5jH1ax
F3fwpLYSy9tmh7sjeacZnNtdYFkYt0UrqQsRtsAfZlQn3bZkNF/bKUX+6BBSwPel
+/EnMQnf6fSVf3TN8gxyAthVjkHHXwaJ96Nw243yVajomtqim4iF8YM3ngw89Rm1
TY0Y6lHJoQ5ybBTA7BPpXRvBXAGugi5GYnDkQ9nQt60LdkNhX7mcVJRgkbo8FDg1
5O0gkFP87aWZ/wtmmkBksHDTsz50u9mdrnItpgY6OTVIH6EPHjlGBYYw+UREZqf6
EQGgW4kEKkLBul7bXBprwu1q+pW2QWes7VNL3g5zQymMptmpjul1dcA0uCAfTb9e
5fdZ+elK/pTKCv0TwD++0G6DeUYHe7Gmz3wDk12fbw8+qii/hkL2ZnqeadW6vja4
OubqNRgjlSneuAvuqozzH+7yjVJ+YuNGaJSOcvEA10DxMRSlLPxIJNt3O48gYFPA
PXu+hWnQWbfYdwFxe9yvceXWpZYvpkdAeXh0OnUsMwt9TB2fZT6bKt5oL8QOnErc
5qjp8gJDxT0dc/4vffApxOPSbxQo9Hgn8JLlRWiVtyfoPD0qun68tIf0Cdl+xP+D
NOQohWS2kQFEEjpZ95gOEfGsyBCiFlBDvUYY8C+bl9mtjKY0AuarXqEAtwO2t/zN
BPZGpvBMovtxbabjF+yctzHxCU4wsVlmm5pDeZsE3VJE9VQBj9esl+r1xKvMvrJ3
/M8mFJlgWcAGpk84ESE2D9fN1dGC2Vf3yt0UcdiAEjG8Al+COtTnhAZBGo2Xlqp+
QhUTo3d2ExNjlKoFFVgqalrkBHm5WdKV/hVJ7pg3+0l7+gahdVr5esVnmKzdA4EK
qn3WOF4DuL+L4qZmjeEnw2/5jc4WNLK6HLgx44ZHKZuUjujHFMvh3UwMTbmvyqGY
1fJ1hjQ1fG4Poh+qiS9PJtgibkwkx6Q15MQverQPPZSoQBnKwMiPcpOzOawTeuYq
CxKBMX3tdorgfdP5kmweoY9twfU91il3J5Git/Blysfhf0Ji7BE6wA7NgjOA3nOH
vYE06pHItIP2W4UwWiCslB+AacJrYAyW1qDYCsdDxWvxU0rw1s3OVu5rJXbehrGI
Ks+ubw9NwWx7jXqpc0jDBuNOXfVa14XajQxNx+XyB+5BaCPUj0PR3+C0j4LjEBuJ
YO0KTwVoRJUr6qj/Czc4qBpb8rOEpFkRldAJiMoH1Uq/DrDIsy6At0At0S01dBld
1rvyTMqZVoyIbU5VZsWS06M9zcqxlfNU121pQEwPibyJXP/GTW93+qnqeLl/EKmr
zdrDLokM5HS05W2Ovemulrdnt2tDpm1CQzTCIlp8hJ5QBqgJtV8ZBENB9ug/fR3F
LcywHNgAFs6mxIYxqEKcGPuLPr93hAgVatQLL3mJ+UQL18/d0LKHMx1YskYX12fb
0NA1IB1i+nu21yMW2Jl2djVLJbZ023EM4nqtOWAQQTr2xa/toDVufP+nIZqEViz0
+m+/0ar2ob6WkDwj/CeEv7/tSajwD4FALLUOrvmQWW7mHDBWiSfz1HkSQ4XCx39M
Xzkb/LfRyrv2fifOJF7wcjGWWgTOZe59pMmTgNGAublqC3pZCMHBJ+XPTQEhGO4j
KMCPsrDcjUYLMXVLPNeirXYDMKk33JnbMRCCKblcSXan2cS6otme7AHyHeJ+d0dL
fXX3tc/5/h5rdI6nPkx0qveIAAcF3uxvtGqPw3CdkdgFSlGSQM1DDAqRug3Xp/jT
krYdgjJ5wCL0NtnuS5f3zic/EwQcfMA49VDSMdFq1UgvqQ7b7Q0Asm+iTINpvFVU
gnw/C9tlNvjxAf2obor6JSALhJ+Rxkzpo00upZYmSp5auBhXkTmFIP5ocA3B1zXL
qdUTs+x3pTirIM1FUtG4MzCLJxe4GsjHaokwUslFo8yDTk6a+9fwtiyyKRLMXHAi
rYR9XZsm8WZTMhgNx5Ie6HF0C8u+xv31utxB3+WKtBV3E4GY9dix32gpr1OQL8FX
t+GVGrSRNmCprelG3PpDLr1r8IOSxaMZn4pjHVXHfau7CqizlsiCpSpKCDUq5Lse
BtpgmWpgtxOOZJEf+toRWm8rkbcHTkA0eMjI/4Q3Fey0tdIbwU1FqYDmMl1ROHH7
zVPKSiWv3lMAYzwrKV3IsekjyEk1JSdipP/74LZ7zixElWuNl1TzFesfoBmsxIS6
cqex+Sh4aYn1XUgxEsStFz6w+to6sC05FMklKnIB6fsnywoFVwhps1ROoXIZc+hy
cnT9yF9AsolennwEyna+rLPIIO8PYskaBZcfnOSFoxFiV5b8aq9Je5b8RBeY4d9p
dn4Ngj7Lq2pqbmMmPJFAwisHeX5gK+oKxo/ZmxBHf9+LEAgO5y6m2JBLmzJbhIOh
Eo6q29LotpvSUcapANteI+uNmspWeKtNDEWc8vmF+/c7LXoCMqzZIXccpDnGIAWs
luJiqSOg3kAzZ3qR2AiuKCeHXkGDdl7IFw0D7aIVaab4PQZLdWhKztrJ7bG66oKZ
mPiSDyihiWdBFqvVm9WS7Sa96wIsE41Fm3qh+v/QZWm0OrFYN84TtdpsReeAPQnb
HhVZu/y6cRg3ii6tc9hPdlhRD1oouX/UDKBzFpsP80KOxQuNpalw6HY/0T8oVTk7
ykGUNjIR7DBlMLCk/1STV/FGOE9U/RUfDYKCBc7thb+AiXIbBOAXEAWpZ0orFGLA
IuwUsmZesaXnrH34zUkHTmYMfFO246Fwey7xQvXHsAF407vGDghz0uMQEsMG5rKb
5gbXyys5y7I2xJf8fl8zcfJ0N6KkfW2ClU2zSidhTLrBV3ItDOgNe0AYaGHmUPnM
RJCQ95embzwVot2OxELGRUxaEpyTHicOJa8EYcaKjv8OELjfaJbmfHLhJqDhyKLM
bmQYWcE61QxZwK/I5Rp4ZjV6YFSA+f7LDbtsobi6XzPX1Exydopqgf17E4Gnmz4K
InWv0eQZoJOhoVvb0DxUIb3pr5E3BjUjPJ11JNMnCR0gGNUPqW3vXthP9lcRzGhr
TyK73njfsrEIscBXYRJkDiG/kn7QqgX+/MYnnh/vG1mGaYWPJvT1F8kFU0CTKqK/
TReXgjXp42CqULwam5NtSk+lgVSmjMfwP5S9OVtkMbiwyrCwkU56EeH5OOkT1r60
LkVyu5f+Pj0gipafDeGTUACUWsE0paEST8BrN31rM1bwkXeUyGiSe5lC8ACV1vcU
/Utr5RpXgvx1PfOGpmHbNjTnX36l8mnN3tAw+DuQuhU2vQ52hNfKnu7wxGsdVXKr
AWCKJ3jpz3smjCkz7LTjSybQzC+BW2+tbXV6GOR/v5j8+Yi+jGtgC+WRkHOOx5BO
+vXBODTUO7vR7+aOn5ktAy+JeHqax00BrT6aauSNGyNXKQkDbg0gZU+Xs5waqFL/
wCd+7OEP/2ksRyX/j/WjNIGHvyf0W9BQItE9332YVxqT4bYPLlKs2YLvT8sZmppq
5M+iympCKO3FplPst2+N8F1Fi9HOVbpYqTpYLyTe0UW2mBcfw3ks5capoAPK31qy
RfKCmOB8+0UEYaSrRBSq60xzFe+jX3c/gr36vp+r7kZVCxJ8s/EcpRioTrnW3i0R
xAn2v/t37IbCbiDzqtCX/3lJGIOrw+KUdulGONpt7CWR6xcLWuFDgreoAxPcetAN
Via6jr/GFz7c6omqBOdxoZX4IP3uD4+HD4JXfu0RtDH+6vOtQ79Y36GtPwEZP/x2
Rhlqg8UXz/Q6TScSLZjb8v7CeX029D82ylJhjlyZ964x2dnOlsXKLtmitBxru3He
UcWrPSudWa/z1nNIy1Ec7P/mGs9DFSBYGxpxo/BFrBgpyPvifU6uqglt3+7R31Fw
avkaZVBWkdJFkt+kGZqTWqZycEIJyQAlTeINSniA/zTC7HeM2PdcoiHIrdRSjvLU
oVlAGRSIVlvTS9yYfo3LvBz1wbtnOUL3zH0mUR3FAOQ3PdRbyAiRwAPE0VwsAG6j
UDEYbY0mcL/I7+Z0jq626dxgayObdOKpCCBdxNAXwDb5Zd3KSf8TIQRauI8aB6og
oit+vqwwXRbELS4u2x1TOVm+5ftgkX7DfBgtNqbBjROVYQhxiLsum+JwqFrQX4AJ
UKjz2mB4VvIOsCtElwzwghOKnmsCCBkItuTGEj7TSSzt0gxzQXOOxtwlVilPPTLa
Ox4EYIBkAHpvS0w0Mw6EYCTMH/aWVPKdFbC/7DjGcI+tv/kCgYMOzG7J8U+3OerC
P35f1Vtzw2jSx5Dc73PCpzVybIepRs7qZLNHblo7T7QccwbEfzx/hmYS4fAUIZ6/
/nFionQaVOQghpfLjiluUf5Sl4S4RWPo0NeYXiGe/MZYC8woJjDZHZTLFcg0xQWS
q4JVjj8/Qh6ZIhVTqa4i73bf3JaqtEVWkaKlbQMwvL4McgYaI13eRrzUTT34VEQC
JVnv0mkYOAwgV/nWuRKpvxJ0hXwBeZx98sHr6XLdNz/aVE1rk3IK1kB9joSGmUHI
8Cc2RTXKER+hcZ8Ix2Z208tvjl1LbHEGr1W81wJdncoVdVI4lB8Kb0k6Fs4cIvxH
eHtJYEIBVEbmGJ1DrPCqL85/Q96Ra9cqB/KnYAq7cUk=
`protect END_PROTECTED
