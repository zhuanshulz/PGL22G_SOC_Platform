`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zOnfugCKKjgp+ozG/07ms9ZwwAJox3t5d3SNIfVKSKjCYSRKoeagXtSo1QLNDL5F
jiHa5p1UXKLH4DIQPRKPMdibs6cRzRmH4h2pVddrDoMlrOWfhBgHUwDmqR5vZ2Zy
lFGg0ncSYAFG30TbS22oNiD6+sySfoJI48CRKi9zby8xAYR3MlxgtQgGE5DtMLH2
QeUASqpBWuXfI+S71w1cRGxnwXp+s3+8KCyfdIlLNx1Qo3qA5x4I2MxO0/tiFAl5
qQ3IC4QCP2oS/ClB83VeCcYME9/lJJkpoaOJRR8aNyGhJY6kjhK8rmNdXY8OPPIe
v0ENsFfxCevbzAQ7jHHmtPhxVZN9DlKRBcj3gsB8bCGa12Jfh/vP1zjPAHmnTsiW
f5zCSt5s90V9dmmSqH5FJ1ccASecRWYsbUqGChyN98igi+XqplT9wzEfcpNI/1Ow
7lVriJbNZG1t+M7n2saH5i+NzXaFMgVz+yPsYwxYEy81BjiZwON8yOFDMdesb3kc
mqkLLzokJBpQehq9UKu/hyN9xmvjAY3KutfefV5AyI9Ps3YkglzLV2q09h5CYrU8
LNLuqTyhKs0QhUZTv0MgbzypVqw9zI3Se6qCx59kXyoJQ9U0M/8/kvNyEEptzI2v
`protect END_PROTECTED
