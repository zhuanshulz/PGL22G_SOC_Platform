`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0dZuk4GQio1vGdWwrLCawLxR/llNlUMrqliO5rUNJHuICXroDTAFzCGAcBDuw/5
CAvA9U2a6eblBM5Hg0Q1hIo6MlKNjiY2bO1GIcQo0FbfA1IB/M5XDSDcmf2NoJni
6e+Lx1vVz/TzTflA1PsF7d2ioKC0GhnvVZN3ywnQ5Y0rJU050t4pMwYwnKkUZe9Q
dO4tHOJSK8bYWGIdd00poeJgZZGHADN+wbR5Dk87Pyi6UBFHo3+/yXE6hc3nyEnw
vxMnNWlAwDMmehgajTHyYmqn1vD2Gk7cSUWhlanlHurrrNxU2nimx4w1ldly/k6v
kO7aHU/Uq7pnyiCZ+UVhR8S885cgw+X/5sFei9Kt9O3LFGnh85fu54ZX9j6jxUCX
IrfqSKpuLgzE+NkPVMhTCw==
`protect END_PROTECTED
