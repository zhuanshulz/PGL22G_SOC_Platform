`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hl2VJDsEVJmHQG2UKqJu9VrZTu49Z5NWTdZPSKFYpMggOKaHmmwW4qhjYbWJmQl+
t4qHToc5FiiCAh5uCvycGS7isH4GSZYcDQo3pf8JHhCWAJuq0hlXcKrYI0L6AGrh
UjTeR7ya19AO93UhCXusn5xRwmQh5H2O2YPfYLRGK+wkSmBdG/DsMTecu8Nwe7WC
1rMYkQ2IcjmUKJT0mAeykuUOmbbhKBIp1n6t6nIf1SXhtjC8uFW2gXLscANxrbcZ
qEQjnj3DjUQk3ph5z7kRZqe8LjQB6jTvtX+K1Z4Vuhkls/R83U1EbZeGAoNk518Y
p6fUD8HsLnMHNL35xyBAqe42oK2hgg53daaeNC293jbZhI0XY5wGa9ZOu1a/jK8v
NmHBxybDqStE6amdJuCvxjcQ0s1gm3hziiYBGaffltUf/mpkhx4ILXLrXEYa1lWp
Iw9FXjMr0Y6QGp+QHJj2fFByTfRj+At/5h7Y6pxphMrORcmR3hP9RxdvX1uTLlph
to5jD/DkjwUfNg35FTTspMiABZHu1WYO1d0QVbz1IJh31U4SPk7YwCTdgRdgzp7t
mCKiIuBbLajECHx0LfLuNw==
`protect END_PROTECTED
