`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHVQtu5Ig8+0tlx4rNJz5fh6qufDmaByLuol8HNB/gfWIfF1JC9rjHCxaDYZJ9/v
KXZo/TEcu9QS5+hpIr/6cLCsLLutX1ZyWPAhw0uEzckA5b8GNmAkjMMGP0sT1Q93
qz06FGtwE+TadqFZua7cxDzKMjvSz17ApvhZezECdQ5VNm2gLoJ0h+reeFv2qlwG
EWMtO/E20I40iS+vvIz3i9p4G0ruygxwjteTvCj4xs4u4sIXkPZLDHOFgTBxotDm
eu+hrAu1eu1frO92OxJKmC7/hpiPRCPNkL2Pce3dDJA3eB46O1nhvTljNgxSaXl4
djJHKfso3AnEptfq5hS1XE5x7bkiFti5ZsFG1dkSrrkO6pr3kLlEQYB6rNXLRhbS
2d7is/6XxoXSK6Gmkr4b8Ae1MUYJaXC5w7Ae/FCQVaJDUC7BMOR2wmf6183CBUiW
AxhmYVOli6xYjTgctTa2a7LT7rDvgTmcsHnCuQglIgzp2UNmdkUX8a0AH5roMGJW
JMgkJ10q4EwB5dj+19Kv38VcM1o7+LGcMGyPnU1nP07/DFoh8gx710Xadxv1e5Z3
Lw44R0F4QuTCCoSRBdn9MVqz3ElM1tTyih1P2ITjVekSCVEHBcpmMempPurskM17
+gcorSp7f/t8Rky0DELlUm7LYfA+63z/csByTq04miskrS/nAqVHRoDeJYje7Map
P/ZrBTKasgcwIEj5vrktDMJDy7guMsvkhw9EMJNXwMTocJ0S+eGq3TbdcYZdrziG
AgOqEVBJt42GJWUSuEvNs28nn5YfssmLLCODaAhd37zOyImuTG7WRbLmmGj5tjQO
gjFtpXYBiM2RteaZapZ9/2Se3jI2A51NmfLUOWjaRrnJuYPSf75cV6HOHrNQDC0+
puC11yeCgjJRn0T5r0X2iE1a4PwmvMctzWM16HT9AYxrsE8Xc/5FHy1ITxPgfXF8
hoDK1ZFfcVejA5n65eGArrJQ8VFPxqozlOBZTbbCmAg0K0T6MEUqnoV6RcK8Zyp2
2LGLXcFlXu7JukB4/DhWuixlWQKsAflEyUyAVW/YuN5xkRM418Hj+CaaSMuKRlnT
FnRE8nXhLEfaNNOQCXml6DuhdDTzbIEvR7ViaM2JHryehxOqdUOl7NymJTP7R8lI
zIwZ+1kZ5+qAoH5ra+XMH1OtUAqcDsONR/RqMmRSQDASv4i8TAiGdjl1mzdnWwHw
mjs474yBFnRyx6VsLLKUjSxyaYM1JhYJJVvV2vl+v8q5wQ8Q1RYf1irKhoDfa3M8
K3DSzmkqlVhAqUYzLEdDtqJOKUPfNnfnWPQeK9qOFW7kFhVZbvCSJ1SDzutYo9+H
9X9BcLfwIcbCcD2fLtDAxEeCACnHuPpt9sp6Pncr7LSHoec652hArMejlI5Mii+3
Yfu39Hbyb6g60QG4PrypSRZmGtstaT0TXCIz6q1KxJmlarzGN2vtt0rMR3COudth
0GGKVPODlh3qytUIaJJl3kxvHAsCJrTPTYy04egM/Gh6V5YFgA4I+ClhIL1B1q+q
KQzu5yvMhFnlSYjnX8+dtietfcMv9jo9jX+BuVI40D6zhm6k2+fqj29Qd+QgMJ0l
tJ3a0dF29xILBRIJlvpIymiYth7VVunsi0a/NP/mBBpaNR6MrmTszVVmUk9KB9ao
dEz9Icfan4mnWYk6awHOFi207JFizqdg5KcWyOm57hADwI51FOZNq5ZwwVBjUSLw
aCPivNWPEY6rcL5sayDKC6gLj/kxZDlYDxWO8DNqNsSuDWIEmBOatWHDlBnzh2d4
HGOBQ/v+iwu1HdGQem7IQErR4bxqduTU2tdc5Debmw0=
`protect END_PROTECTED
