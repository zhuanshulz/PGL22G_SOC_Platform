`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q9ggl2GOAcmQY+PoAQxDXrgt6MW9Vfrgi0PlVsn3u+ZYIPGpoEwRdjXr943jydXI
xDduxCr69b+qxRzTyLvo7tqfIwpR37SnKgcd/Oo8zhEvA1+Qxh6PCDXGqvYiUUYP
pADZq3cIr4jbwaPFIhC+/MreOwmgx959bhH9D7sGllKn/YOamiZB6B9PT9iObaqR
Gz9qm6Oxg4UgtD9PiidNl6UfL2gIY5o7B+RLF51mjPN+/IwDA5JNWxsk5hcx+TOV
YrSObA9mddVelnKiclSZqa1KTceOP7wT3b4s+9GtNLzMqy2Nm/HivjrPIBQ4E6M8
h6idCss6jk6Fp78BU+TR/0GbL4xJWcS/k7W/5d/BF9mbZrya55Atde+l7UNtq+J+
hDzwazm2vHoLKIOSiZQAhQ==
`protect END_PROTECTED
