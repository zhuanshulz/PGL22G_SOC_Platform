`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GP/A9hV9PuiMlcOoFKoZJQr4anp21XKGS7bfCUTgHwxsjAelfbM7CQPws1owdOCr
OcITGh4As85UF3Hl7eNlRCy+b57ij9WtlUbuQyxbrvWUVgcbS9zV6JP/HVWB22Ke
Dd8Ce17a1aY5AhTfGb6KOv5nKDWSvqOJbQw27I3dBvBptFKJHKNJIcCONUqfFiS/
gXhp7hGwdi4urENlxyvLkw6xEh5jxFJRkPP3770zkaJZyKu1OwvqWbchqLw21u1q
H/+yrbWFfhv/IwPkNq2CU6cyJAIAs5KrIl9XDe+WMDU=
`protect END_PROTECTED
