`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9eI5ZXRovBWoYKjwvL+2J/2H5Ic+Vdy1qhIYUeUP3YyasUB8pwABa+YiW3+KkX5X
sZsfZRThCOp5PuKRL9WrMZI6m4Zzs1hMGrnTwDUhObWQdglQCaUTCU9ks1JrtPka
ZozTxLP39c96lWSYfiKLllUe58F9qZLEzyYeAyyRjS3zEhEGNtufMuqVA7A1aXA0
LIPrELT9JIHB2r1j8qHiEbyWdvyDxX66AoGs329va2TV/IemnPeTmm1SRoepLYFn
6IkRcELCZ27eU0U6n4CZEDV1Xk51/gRcUYzFJYIIWghQTxKBAFIsHpzH7rGvzNCw
S1cGrh3ajshwpuEJ7oAyPF3QTsM0uf279eV67TGNHNCKMgFqjhd9gtesI5Nu8JMU
y34yk08IaCtoxUitn5iAh1HDm1GWjHGPuzrU72jOdzOx76QTZVqnuUKdjQ2B0luL
`protect END_PROTECTED
