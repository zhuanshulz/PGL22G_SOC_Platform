`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y9prPoFwE4OhTctdXIIaIs+RjpToWIEosc6NHQMEjLb3oWXVsIZHdsEpSu7lqtOB
IQa16X8wX4VKLt2u79HMmHUPnYRzPul2kDlALMVnnZFufNauDCIqJ9oiYB8PXnNz
ZdW/us3K9qJmQsIXepU6qVUzUSlChgLQPi/eaHqh/StHJwI/DY7BGXMzC0boCTPU
InKPr56i0ik6mv55InHG6Y8y875MO42kA/ix4XAAz7E4/nN/9HSjhIcTAxDp4+Ba
g/V7+8mKcQ7nYvrW0nspKvL2RseHJOm525Z2D0tzo1rWKFmKw7vDGqLt7g9pi7rg
Gz/TOsTq9jYTGAeIld0li02+ObUh9SVZOAVcevrhh6iQh8ykggXp1w2dhzgRvqCT
7tT9BpBBU7k/wb7YdsW0YpJ53rphAgdUxR0x0b/jwI/cRa+QS8Mw18M3tRFyEcoc
6ey7wLZNVlw83E2NwflazHa5X9iEmqUyj7mgLBXoTUKYrGi44QWAaUfbQjPLKbqb
vf3eaBUHJe48FfduV5igfsdkhjW0YSh2jyMcdoCNVtW+bh0m83Wox6BvOjTTN5q+
HIx65sT4jIFWawUFEGYD6w==
`protect END_PROTECTED
