`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3+OOhi82tZnQb5KLph8/rqMmsiBJAwbkyIXEoNL8JoFqOfmJRKGvVoHYaqhxDf5
eErRoa1yGg/eR8RIzx8OwjD3ScK5rmfZnOzQHm4AssKG0RFJOleypAV8wCSkFvAV
7MLx3WROoiGC7gLvsa/qjOWxO3rfHb4eHm2Fv7C8VeEuXRjrOS//VWHpyVohTw1e
k9tvB8MkoLQjvksdsYijjsRX4Y5u0xbImNGAi6+WRYPbpZa/1dwKn9OlWUelYTt1
XZ3iO5IVmwmuDvAKaUtcTeQazlDseNR3W9kVTtaQ0+Y+XdbcxTm5Jt9qCHv3dDyU
iNZ1ozXZXRVXqyvG59QIQwlTodRTIQPByNuv70weykiEbMrw88c28DPFksIOvZe6
ff6FfApA2+vsXKlmE52ryhS5tZ54dkgiv0ftGRCl/VJLlnn7D7lCtVzZCDiLWM1Z
qXaegCwKFkVJ5wUJoLn3RgjUuRHt1h7eWjtNLL+0Q+9TnpkEBWYEU9OUHeDTfFDN
88RC0y8sIauOdswzYZsYHmKQg6x9/2ZqEnpQSYpH6mMjepl+6Q0KDk4tjflxfrtX
P1MaHMI86XwvZTttEGGWuk4CmjZVzM3YHf8kjchUfn//a880LJcF9U+6/NhHCJ7h
bcgW/QxUO6MFEApdw+YlFhzLSlH6JxC422GaORuwJ0Nm+OMNnTvDVt2UE/i2hyfu
ongcd7cuU2kBleXA2dqCwAjNuGFfwqLbfLuBy2pRzqh52cxMDnbhfbK3U7QeYVO5
uy5xgDhiKRp1C6R/BLjrSVYw+g5vuuvnVANRf36538NV3mELlrGjnKoLeKQNqAuX
CTFTkW5J/oewXJq27Iy+cAGHf+3rW8V3Qp+Zcf2DRtLtUbhRsEo5/u8VSI8wMoHA
z9ydMUocv0dYvtLxUpGrlUe+XbDwM1ceun+Bf7tg2hk4McfiR0r/oQcNlvyB5MYK
Wz3YMnnvdqoOZak9pL4LLhs3wZggfvQ374H9rcNNRctWbl6Iq8tKZDZT+4Gph/v0
NS6Plqa5B7xNfO9+D5fDb4vGCbDzUMgl/CrPahQS1MVvDXfyVfxTyWNStz/49V5i
/c+tXmcDl8SQg9UkUVCmKGiDbqbS2cK8oIXJcCYiindI/IhvV2zn99z76Vc6r+Sb
T/UOft+yt5F4N7K68pAIpUYLaeup2f7BH7x7VIP0Cku48XIGCnHcdMHj+Z0YX1AC
hBBDfEphrmG1RYyB3/c56IoG940s1A/kuYvoQShI/guEJH7H+mXHrKiUS4a0blQt
ten7V7WKLpiDucfWfDv/A/7gZ+LBjybVaQspM1H+gVq5AmcDO5RoPB3Tr8Qn0G/6
WvuZMJdCdXaa0cEAWhkpJ7j85NBTp3QOIKizMTEesJZ3av7Hmg4Fb6WVucFj+lkw
bmTZhllEmOw62vVRfBXnhGimMOANThAom7UEjqQrQF9bM5traSQn8TiXOJZQsTX2
9VxsqCPVo8ZAAIi8NOrX1LW6tAmTvjQgEmt58BXfSKUIv4vQKyhVQJhcphxulIwn
xPWkYKTdE7jv9Kt9c83x+MvV1LiRsAPsgMAKejbTfhq+ATcNvPE9DIcK8UOOzv20
XrmZQTxYBBps8PZRZrPD7K7fBsbY0wUcel32UxAfwrd39CtZvCTU5DB2anmiTKRz
f97DH7PP+X+m6Ca0MumemVpP6L1xbuXD6sie52rJ1Iva2fLaULuByaVdimg6Gus1
5d2of/8a1/VbubS+ltDarE+4jc3RzMCeoE98dM3CzN7R3P5OwcqT/h6wKz+X70E8
da3+3jhkexC0aE7lG2u4Udhvu5N+t3Z+IY5Qm7UPEbeNQjhMl/hkNZerZ5pd3+W+
a0ocndGZDtNA/8gesFiQw7Mcodqd9rE9L9TJlk6KDTZq2TwWeDSxloS6pMGPGoBq
irMdiUQtvd/K4/INuXAy/Jwjiahqxv2O68E9Q4i5rmd7KrZxC1GRNV11gjmNYNjI
DPGuiUc8ChR4hDHWZ3YF7nOWrweCJWYSDX1A4XYSuKKjlSWO2zTFOqnAjSqA+JGj
ZDu8Y2wRSm4xbyW3zNDXk3gZ3l21gBcILPJy6WyYLRzoCSGcO7si8RTJLxgsxAZB
zStfXVUbV5PfY+oOClL3B2d391Tl3qQcKTHkRG+2Yn0kUunXffrvGzipMTFUw/KB
zBPeiWGX7OJa1k7BjF3tUtO8JrHzO/GWrsiPI8sZoeeW+cCe0yt11Xo1G4ZG7bPx
OkMnJmN2l2BDEjihP5jdzoNz+RG/RejL2d0IKTu8PluhMzyQmz8Ohd6dbP/1vn9Z
gr2oMTmVjoTt11Cezeg/QDm/lH2K1KkmWOjzPbFCVkhJ6EB9SPpfhJpEs3XBI8TP
0u3Jox46hwOhwyVtRoiY8QP4coCJy/L4WHBGW51+cNOqn8FlM0QQD4jAz3AeI3Ft
hREhT63EASCJnPEcqrli7DL/5e7SYWKlN3LMuUQGClbXypOtsAwKKavtJrxRT79+
3q/LoUTEWtL5ZXP7QJ6fuD5wnPZIRpzPIYuseHjJVqlGgPvpS2E9Y0NZkeZ1Hvlb
i1JaqHMpMDoNaGir3P/oe0KF/rluMJkkoJsq/pi2upsRCApLsXI3uXX20shXY3u7
vMqUQZWzcpyhq2jYu2MqID1sXRcXRg1ubUu6BMiMC/WvuHMp/6LL/lUTeqwzCpDc
OXTE7W9CX0JzlFX3Dp+WSstxfZV70WCLs1dhSzq7ZbQny87CqCNYWLBBp3+/Kz5N
QxdH5iFRKtpCIkzhWvMaVlJV5R3rDdt3ChOMfohY1PyxgLIW3Ysp9dairNMYR3GL
PyUwrwYCHSYO0j1VHI7Fxdcv5Im2Fy14REOZRsNWnFXUQevcikkJW0kYMJjnEYRI
KeDSyI/BT7BioSDW7nGbIMdhn+NSH2JlfVPIyqEwh8OdLtpeydUiIZk+7Hd314FM
mKMSExlCL0aQY52opj7j7iokJTzSbYR2Uel/vrog0KNje7IIPx5HhGexMV4sPNqU
jL5HVLASp+PpfycVGMeJ0fh7VIaCZYAmitx8Bco+60pla4pRtcw8rKahzoyZ0bYj
byBfUd83/FuMgp8pdVZNYTOjPb4C3es94Pvf3jyvoXofWcxLtZ/C0+yJjxj2MM1M
QJaV+nNjVPXZmVBk9J9P4H6kl0TZFAaaBpwf6evGKxoBDkBQTAOlxB4NYi6a0Asb
j0h03gQo1PpZawAVnlvBczEXP3QWXAALuWV/kwFRL8bv5Iv++SFbObyhGAAW1mPO
NuqmbSwHc/gdq3PoOEeOzY8OngpcQnEt1GX9A6LtVIP3xzCG1nLJkhh8eoyYtnxY
DDga0F8QNBeZKD6D5wjGpJyb/doeMBUWHFWpR7jOZ9vuVPtBWNADWgTMl2xmBHds
1ZhHwmBSmBURxN/rv5V0UqU0aUCvgIgkXSraJ/q37nY0i+rGsuL+EfIWHqBwWtfF
0IZX/nmgnzgf9nUxhRxAzzSdr3mHCsyvNq9oDVd6dQtisJit2l1vZrj++kzDH+rF
tdH+TE9entZDAPtHSAtmrOYJyylPtWc6HtVk86LcCv+1xqZB66fzP+sgiivFyE6J
JefrOAjv+mGDkiJUE9oNWXsAvWMV9GQpvLWhA4Gk2IxPaiOrSq7/8aLmy33hM1P0
CP2+PyyyaEGNdXOOELpUZGuC4/psXc9r7zxkzexplUCwJo2bzhCP2o/FjihreNTi
rKABPtSxf0IqjPPnNzZPbMfJxK15CGKibj4a5fjbTL0VB8b9E79xNjPiJN3pUACi
ehXl8F6QJP+oi99AXR1tP+pAOjYXFsKNzSY7wswMA/Xj2XOE2tkq5n+jOR58r5gL
gE4y0E2lftWK7h7zU9Nu5eTr4p3G0nYxpszo8frf6g9hkrnCGL2DXPJI3Hf/cEYt
bT9rEDAfuVofO2RQ/cLJO3kU9yB1IIbR3KoJIcYzUYva528rrb7urw2+Bz+3GEsc
gq8vJhDda6u/548XRBFBQgqzwbYJIUnGrI9tHBjWOEnqE8ivwA7dRIF3ewU0BP6Z
d0Unx9EXB8wXEOYdWSXZ/H+1gG3qwKd2G47TRa1Mp+Bfsn8w7BGCA//5NAAu77g6
O9yqcrYQCvJjWF5oNQnaoEpZ7qgZKzTTRZZszWO7JeRaKIHPIUiEo4Wjl7KAZn/H
kA+8Qfh328gDAfjkB0gA95YrrQlycGVI/sHTIWFYEFyQ7CaA8AIx5lbuOYx3341D
2BMz9WoszRgCtWHDu6z2cOtP82EcwabmRi28zSE1/Kz9GqB9hl5Sit6BTaDre8JA
ykit1HEwZYi7d+BeroUoKjADl10DgG958BLli002klwiW6gc5cUo6Uy3T8L6TtYU
FGRgtqx5hFgreXx21wzJOMRH7VzZydpqs5TTcBl5cMFO+4Ufo1ECXTxbnznBM4mJ
siUxjUWz17jwoZTZz2I1q1+S528ZMvOhqDZvcvyTyFsQq6ouJ3wUA4zTUZgKMq4g
/QtfAqIF1ATLfVbLf6A+n6LKT9DopkY3yhIozxlADMTQnIPSCA7YC/NUu51vcFgq
lpVQT+p9mwHR7UrxJGKfdXcbSz5vT2t+sjdFYN6jJ5bSxK6/UzSDb/5CzvIeSPFK
kfc6LQZV0/mNHH3ww68uR+XwG5zEUwxI7U+lP0uw4jYLCfpyteEr3KR4PPQBPb9O
aewSKywk+9QMaIvJfmj0gZ80H+ZpZ49oH0FMSkzc4ykZa8qV5lHjcM9BwuGcAcEt
4wp1M+mjora5Q1K3+Tw5FFWbv03mEhxxCrez7izgWGC/gyvaJ9VeTOoatjje2M76
P9wCA/fGjMlxyGYOzIzVh/cgS8/73wazBXOXRWtKIUVz4G2nluBYca6brdW7ccRV
R43frNRCLgKa4Yv7iJ9Fta1Ev0VUH8kx/hKn56VJvCJthphQ9+lc7cPB76m3tpbT
2XB7CycXCOJgVsTQCDV7YJc4myvO/QglpzFmPui4L9jv+TnX4g7EJQ6tmBN5Pp4H
P9EpCZSAAirDNSYnePAKzrBshfojXTfXUdJhfTy0tJfe3h0g5bPsjf76K8k+/Cjw
pY4H1yPshxv5cDeVduO9SWpeVnH/2/QV2Lkhdesc41CHraeSEHVLtm7n4dp4T1MC
4dg2ecbTBZCSiPvRHFYTqSl2FxBp+69sFw11BdBZs+J4SwSk5wjMohyF6vdavXnM
rJs5FkJF8/QGMTiBneg/pr4XcJhpy5UQTQRtXdjKB+BNReS3E+S/CZyouqAWuFEA
bpB4e4iVGeW3uyznkcnMGE5m5FrCGhqi2+VZfdZEYu81dCTO0fauaz7UTNWuMgW5
x+oScE+IvDEB32El6Ddp4viRB7ouONmYlQy1R7MosfnB1Epf+cwkSjeYgWbZzgDg
Tnk8m7MzEfB3tNYBnHMzYfV0JV1102KDGYzxCtV7HkXSRq/4JfgX6hDvG+pedQrg
QKVu+Y6Zf239va8gp7x+g/MkRo8tVC7YxE7dpJmw0cFGwWVT4GHpbsSxueizB/oO
lKxzQ1w1Ijg0PVi6adU3EYiECk4I+LS5FuB7TWFfwMQ9k/MJ/W0Wx8em2Gc/zudf
1QKt3//ue3xWwJC1I8xTVDHhj91wO82T3U7y0bPip43fhP1c65+HHQYiFybQsfuB
hVfm2eCcKKbGsVtLZDvkKLtCXPjkKNAOAVaPzOBBkzYpyU4c6jtXqCakRJn2rNhq
FBvnDHd/aT/sBX4OsNRXTZHBORxJdIIVEdtKyfvn4zIYQQ7i2h+X9W5eeEtcwYqA
uANkAMtRjp5UryrDuojBVhFvGhmEsgdXm1QwrLPCELVPG9417midbeeRN5zT+HBz
jrJk2UtPLN5KzXx0IKj/zPzrrgtWROnZEgoPB0+kFdCJXX1vOmpMaiMcClv0UHGB
RcwMlS7kJ5lnb5HPG3vo1VPQV//Oz6/9Gj3Zi3mQ5+lfunYxj043A+kHfMHbBG70
oFk0wUAACrsT7jF2AkEK22ml/1cCoAF76d7wzoi43Hk77CGmqWHDKCOAiEFHQgem
vE6qQpHQB8HlWH0JW5rOlSAviXTdsAoOz/RcqpoD3DY3Lhhgp/MfmMg4remP2mxi
NPEavHS4rKhIuaehHYY6f9TCEPuUrbAPBebSRelQSdQ5YDuxZWttolGKmfTUWLjM
6lucwUkHhX9NgwundKcw2/UjRAgzvZFSgXbdO38EkMlPviAAzqFcIuAmINs8/Rvz
LDOAcUUlkDvosX7cb3GPOARbr+4VpDWbnldqNjuZBzE+rVg9iT/gQzrUZVuwP8sc
Z/6uXO1TYXZcQ3xSiGKNhXgCL+EZA2S4T6/RYZAkvNDEFJcx84owm3jvTbAGFiHF
AcDHooCW5ZEYmlBrddVfiKsT3RYyzSXF85CS3g0gRI+zAyxvs6hdziL+YBi3N3cP
mpAMr1Iue3IfAX2C4ortThR79KDH9oiIkEyniDSa20/WwKkbmk+adqrk/w9ZC0HA
6m/gyCLWbeEgOzK5NZc1athObvilxr1MrOaCvH4If4GiroRNnoc/2ckHv17qVp2E
WK1iVDYNKE4tApOH5FKM3PxW3nI49t9XqvtEsk4VJhl/VbYhQFKkW66snevc5vOP
SwRVwKA8RURzbyAUMWDunZXOdxycxawdnis85mnx8sWnqNTD8nXcG8urrwqetgIW
fdDgIA/osCxFaqWoswJT9r7yntZHG5npcORAGcizRE2pFOIT941AZCY63IxhYRZI
06b+MX1/OUOvFUkQEyvfXzeCzA+ONngyJRASsJ8zaifAjLYDbard+IaEMHM0UEeZ
e7peBDl5H+b/bisk2S0Z/mrzUF5xNr/igSDng69Ln+aaNiuT8cep4fk2KhSSTSwg
/svBTXMl7Lhg2SQYEp7HPukMfzsQKiDA7ASYV957g9XykRQBRuYhrmmKL+6tnq8O
GsVfFwQA47ck+dYAppy36jhcdKEG6I/RaMjtm05bNRnAejOjh+kXEu3S//ts6c1d
PemDl/jmaWyMVtflZFEkzPJeTQvgiJZYg0yJSuDkp7utfN6wy/V+S6bnO2QVdPMD
kqIAC0Sn7aYyoPtThlDa+F3ujzIdm65aX9qq13aCW91O1VWgHtP0rq4w/XsBVlbm
O+PSAh/TMxDNlZUg2KSf5oS4ayeJPJVh7PsChUWrLxWjQ7MMArFJymaZN/Ff9wWi
BR2jRhbcQ0lbFbHpgPoy0+ViCJsTOQQpoZdc62wzulnSAyS3LOTL3mpayZ4r7kUW
ZT1Z6jCxyqjX97kAIk2p3AxyGHVWcwBaqjYwdTg+DrrIg3S1R/+3k9VSsEOP9ulr
PsKLt0qYUb650IlCWUy7BGlu6cfKOlQG5eO1F3kEchRxmj96/SxsAP/Y86koXu4g
G2FHSWER3/lF/ScvQN745xSQPiK1bqKkYxrHJjgvW63XDnLZTvIq+TVxu7HIZgTE
Qs/ddFyUYH+dmEvA1k17O/UQKLjLCSdOlaCbyNCc1HNXGS1/1x+LgVCzl98G3ydw
UbCwMi66QpzPyNKDNFbw3T9JeiYhiUceXwHPo3dkBFCrTqnyOVTbr1p3NnzayJ5D
CI0LFAy7i+wZde9i5lOQuDDcuoMe9FbOCbhX8mdj4lwbYE/sm9MHwVOZsYYGmTzL
tJuUKRLGNOm+aUZPEjKh10NFtusbsX3zKGsy3NrUR+0Ad8OUfubLUyEf5qRgna4u
eCZFQxDcJ3gmIU3Llr+EH1mY2LM+d3JcYZ//RILO1I+2AxyxT0ab+2VVNUtHysCv
V62y7lySFi1NQ9vORi8/2Z754qNiEqleYyfCkgksDlSSJbBZp7CVaCPMn7vNQXJ3
SWxP6iLvyJ1Ud85sHzm64j4HRwzTIP09toda1LcFOY2RWTdVIljqGEmWkgrTx5N9
XDkkkx1cxNMU/GBhssQs5Uo6TjeqAcueVXFSC6G0PGsadZd/R+qbIDEeK/A6FsO6
wCVZBuT1hxDY45Wo7kMFVecTrBqYLrW3dJmhZmmSYXVJO7p17pMYmMBPrICHyM76
ie7wrAkRLXHPPRJLXS3PPuoUbwQnmcV8+0bvgZ1hrAiBhbWWhSxOH4CGoF/PPvPp
yALYs7O7RQBYwshZ8PJsbfmQqR7uvrLl2zom6Jbi47S9EDIIG40xdElXSI7hzA8z
c1zWccmfdRaHMpeotXtsf+Uy+d91IJYCfEtjYJJzjYOqZzI89OhEtZmEH23OGSPO
+4TTSN6wwf3lYk2dB7lx24mzBARNmoTivv8KEJhRHov8UI2fI8fT1uo3a5ImTgaL
d5oGOH5kmv41ByWcoqsvmKVh2iFggff+ObSpA2mblixo6THQgzg8YkD0Id7DQ8Gr
dub9kFZUJlZRxZ/qFXKkbeDQCOHiYsjOZwnIKl+Pvb0z08xYWlNHLPdw9JeL7AcT
cBKyWQIZB7+YavlaLls0rxsBAQsMtfdyHPU9blTYJNaau9TPQguV6M1H1Mu1kJGq
RNFtyBjon8m5uY/JFyrJsbvMWgEcQPuXdcjP3FxjJa0vhBoEGFIpE9gP4KSMnNVt
buaRZ5LslAcejKvv6Ml77WPi9jLM/dTDHyAo2hV9yibknBi183idAtmr49DitbMe
iFrJnnpLasHi40xnlns+Yxlv3Z5pAhJpM9R1YIakRvS2/n3DgXKmKqPXAyOiLXr9
Z+HsIYrm2uB/EATJdAaVWpQC+axnbGOhqq4w8wQZWMGjZTnMczl3yRz49Bqqausu
T/CQgVUhV4bJ3hPexVQH5VzjZAw4RXSvXqU9eFQXy7991VZ5KqplMX7yvchXp1Zi
4DfPHftnXYJEN60SU8tmEBmM5L1zMVZwJlwjWzOm2s/OeZGQ7f+4ibKpD0CZ5yo0
Zq6TgvGZ26llrR3A7siwVpT57G3+Oqq3P3mSstOZSfgVumK0Lr6NE6UIuUXBPKyL
9sjJlBmq1QXv1CD4wG/RUV5jME7KfmOFkSuMsasBkQxXNSl7TWAAhOHVq6slCcfs
AEp7LU2kl6W1+6K8c2dqy05vPuX8Eyj2v45dx+FSJPDgfeoSk2AVYvZpjlxDawR1
I2OgYraqKoNASI6Jx3qeCmPzXeRL1ynd6nKmwFRAi1BERnFTY/SepE9SQWuZW2RE
Krhyp8DelMl96YhpLDdjzlYcB8h37c0+C8xcpgpgNGlOYQVPA1lYTiCIVkCSSLKz
g0fnPMadasHoqhJpCBr1TuuriOeSgNkKy73ico0ljRqgLBc/hg1XCVLnolW0AkMn
V+4UC5fiEVJxdqhgL2qePXsxTkao5oyOeSJcIZV8YrKX8BCntFDJIS/s2Mp30ita
zMzgXS+WaW3QGVjDp8/TN3UbhFeK3sMDvOZ4Dl4hDdlTCOrW4ljdT2U9XpAIVXnC
FzDz3dSwHPLPGvS+wVFmQH+sRc0BKqAKxm2gaOOciU2DxKOLVI40SERM72PR7H7c
QRDDIv/JSrUMtNsDIlfOpGscQgNQRfEC4E2YL449ri6fETQ32TvhOvXSSLgX0P9j
T8bHduHL1inocY83n/kPrKUk7Y2yXLkk8facXHnWr+itvYQY+p0MoQInuL7tnErN
TCthJD4pGK2vNlW1aAyMV8wLbYlUVVPOnvEiucEMmm6iYAPxAO0q93sYxIa7nK3N
2o/TjiXFfis7TVAIFErzH6Kv7sI350W9xDhjYq4MFPSpDSHNOC98ibXKclEppZiv
yhfYfrUr5JKNTlI+iRV5SJWibs4w1MckkSS70J1gn7p8RbIR6V3muOYJ4IWIc7bh
QKo5fCfJhprnYecTjRz69reeYwxGXr7POWNUYpHMB7PDt0PHaJSZzOSEayAjmVs3
2cucBKl6tLADN27Z0oA8WnpCJbePUKtTuPjLH9XAUxsxn1IfXZHy4B6GFePIzu4O
68C7VCf9QsVLKxRH68vGNForzVe+O8VKBaegg5qayBpIIkRDVDim+t7RP1V+XNHL
DpM8QObSSmB5cwQK0INH00LGJR6z2jkE7aH87syK7o6d3H2+aLhYYE2FgnxHIc2t
AMjjXHGQSeV7jaeb/Kyo6WfubR1XJd7mQvE2frpH7DfOleVMncVFTmOv0MeFZ7wp
7eer9w6oWCS4wnf3hWfBMuuoVcCti0PnnIW05BaOgfwCYKOOdtmPap7JvvpW5R9h
a5zYSoGbAmEvNIPUMdmAql7HGfTK9Zg7oREyi7GvTmsXQY2gN9ReGyU1sDosRQHe
qz6rBrBeH9BhL5yWcgcP3WKYIEniYlc7VN2eSHZVyaHgcTbGPf86OxTYFfKAiLTD
vv967siND55qjAygIrSidbP0WSOtSVYS3RR7mhpOh8ZG5QNtEZGrz1buawhbSII1
+6R+lQ+7T4psZ2ngzNea1npiAyt4DXnUnWxVtSbn+/RIcrYUsFWZAj4qtOKHohjv
fdi+o9NaCxxd4OioWmoGGuP5eNlnaknKNkBEVDrPu6l3lfpyXv+8AV/7KmCUTS5s
lV/hv4xUnjpFw+h2jNmge+qCyN2ZnyGgv51QHIDiUdyPXvK03FPq6PtbYyA6NTzm
zUx3Gslk03CaeSZJlR+EsWbez16W/Sp19oOapmZAb9iyPQ30eKYYN2Bh3s84BhF0
As1cvclw/Nuk/2fBv7qH2fUuZHkpXAicY18HHimIdp2XZ//4TfkUCNdAqg439aDi
gab6koAe8NpwWPseb8QrOD3Svf6SGaQTRVdE9sv9zXhMf5zyTfOGsn4os/7nnn8M
mvoyIOobEWL+tT3eZs4PIkfJAJURNozmy+32xONLNo9u3ZKzxpwijH+lnnRVh8yW
oH2qSi/0VMjCj+G8M4l1a7uhXq8atxEWHO+gi9cnQO42DCqNGdGjd+q2/gZN5IWG
iuD0jtexzFW4gdsKsDMckXAwFzKAMWEEpXED9hxu+MvZGaXVB7nqjPVlPLy5lFYx
Ydb//z/tJ4S1kGwMA0HPhlBMbF+RSoN0tm/AWjeaP4g3Lm7O9raJ9fTT4/SttFos
nttqvirt/4YR+CJHX//X991jKLEoTKA/BgGzg4TwU5ZrUzEM7azstMumg+YoZlUu
r1BsjuUW96pOK09cMbaip0LAptqvlSXgHYs2Z9dzElvxGQfjc9+4rtId+LXSXnDJ
oUOjckbo0xBcr5OIItv+scj0XLz3Z9ylz2saTzEw7DWjatlXCmyqOxP9j71Bdwzc
if8z9exP8LdZXbznzVA16D1vT+jCL/jL8msVPN8/boXEqd1ljS7EFYN6Qt5y/V/O
+EsY/rjPbsLzbLlB859OSJKZ2jUBc3yi2y/jQdXgOCSA7A2XJdlqJ3MaCeyTZPfd
KQxRGum8Z2jL+W+m5n4yIM1zmo0c26bfuIFaNUWlNdYZT5g1zeosdW8PvYB+PA0+
WG5n7i9B06SUjM33q0pNUy7SXiEMf+VZMM5R+p0FWiSekK3VH9mssRaEomwwJuX0
mNUa7f6MlbT37HGWcaldq3w4V3gQu3eiojsYtbd9j1UYfBQAuFtZkf+hpEIusVey
DlkMUoEUwfTpmUN+P2nSAg1WKakhyTanE87ZrjjoKrI/zj3NtVVB2Y5Qq8QsIhjV
9/XHPNchFOF2tIVXIwdd/hcUu2NZAKSVixc2lFHUVjNLDvY8hJHd5iLD7xi9PvWg
NMC6LHAlCTif0/TKoUjZaDfQA4GOpIaE6ySdK4jG0Kn6FpM01GRqEpSe77Rj1qtB
gHcah8BXOCHMZZEsCiv3uuE77dolCR8euEhR73aQanoJlSrtj5shmCZdI2WcFZwg
bFanM76JCX9iU3+eslimzqMwqB1lLjcjMc2b88ZCEtsp5V+IcZ6B7JLOLr4z8WA1
FZNFZoGChgbycRpVbWydiBu0BpN0lwOkV1W9Yh0M01m5ep9aXmnsDMyYq2ZV47ii
lGNS18FmLgaeQLPqyvkuw53hD97whnEyX2GLTA2MfdCvOf0HtwuuAaVQaItP4q7x
NC4az1WKah6Aqy35UFgKkhmofA8Iqp3U2Ptm2+a3DQ9bk/JFBueye4hY7+i8UjZa
nKBHSkJ8nrOzM8W3U3SAChcEg5iC/Oti7IbWBUx3cvorJVjjplfaN3ZTP/v6fSZm
oYRTLrBOXdsd1EzodvEaMWFUyN7oocNxpbm0PXQNRya6ryxFTeNZ5NEoUL07J2Yr
bbNmXVHJA5enptBHUD+OlWOPzDQ2nRbUGxf0GopVpzjXlB0OGSDCBcK5TPINnCbS
AvuYkb2rxQ129UsR+3OXHGnODil04HBND3+viQyzMm3/x9ScImDkUfLX1eqFhCer
IRkkW/1CLOO9lp/Vr4EFgbM83sioKZO6J6s5AR4lEiS9ZPZIVaKtAvuG8szjQLSi
hFpljLemFhgLERSP7GRxSWNZBpwvOHYDBbLkykSDugW9xOWD11epmbiS0EmJDmHG
1TpVebesEiRd1uujSNByREa6BS8Ygt3hkAuTH8HX5sRjy7Zk2oYmykaSmnEpUFys
9hii3mIHxqeebM9vSt6Inx2xEEVRPXn9kQrb5rvbwGLSPeNdubjJcHxPDhnWFuWh
zrOlhrAI27Mh2PoISwmpeU2RutQvGl73zm7T8xLBiXYRLvhZ3mYsa7n45PUSn9am
XuFuqcl1mz2nqSkNJnln3i8rWsv6SJARpyFGLK3YDvWs77CBNQ4r8LX90j95EXwH
eeuYKrXL9fsMjYsZJ+eQ7mqAGrj3CDVGi93liB7foSE24+6KLsPrAA0MgACU5ZfA
`protect END_PROTECTED
