`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yOgp4wd2KbKtrWhKYWMiUZqB/KKrbxmpr9H84txnD3lzktDe/J+dIVoOl7qSPfvp
RKAWNzXx5NbuFIvyahWpLYWSNCkjkAYQuQq5fPiz772ZYLaelhwCDlEQdE5k59Sr
I0pdutYKpB8x0i0hFSyXYxoCca5yWiCJjNElNDG1ORb27aIcxidLKCDvbcyclJ7+
coqbkvvBIpEkMFkRMQQHQ+yoFOfelrKk2+PPGbGDVtliBQZBYCi1N2fIK7+vMw3S
+PegBQxsey6aT38fxdSTaeo2W2+GG3diosmrkCYxs0mwJZmy2vzeBtw7N9l0pfPZ
MKKW0kelsWtboEMTKPJFpbccjc63P4kLxdxkGc5jHQ/vC+dD/72sEVGUikkmY1Zz
uLYQXjq695nqIKO3aC0oSwn02i7vUjkNCieBuE1N5oFCSSTZyRhpqjR9q+VEsfaV
2740HR3r+SDDa+cfKqVYqcawvw+YpDn+pEPVWcl1blb8aUJ1DnmS+KKs4T4jM8HC
QQX7hqd32mVXw7BW/acfpyLf1B+cAZVqZkLvv8mu0bgPZ2EW9WPsCE4KoVIex11P
3VbEX6gWcIIlYXzPMezJo26WeMyuOoIJpiP/H9lCcTJIcC3yGLeRtxAmCdOwVDtA
TwGhshyxeAvWYGAgeIZUZjL8lUmIknPmy6dSWShs+3BdZ7vfEPP8ocituU6O6Nkn
/SyegebDfdL1vvAkbJhBuIvJ6qJkniDiigFybPtRHiO1NNPhBhNxEeFulbv5vlAQ
BXhXFrvSmL7nX2QlpYjgnrYoUhWJYZB3Dhc1e28v28t3rXgr9ZR1GAMgLQHyYll1
RvZQX07OJyxcFNtRJ7z2s8rAo4jZqw2EIneuwj1hNz12120ajooifD0VNj1S3qq7
7coW4TSiVo1pNARjuoD6tiIIiXzTNKqyBrEl0NJtuFLcB6la5UQenc3h3tR1dR2k
VaKk7UM2pqWhzHe8t/RCV7iwCMWfi+5ykd2BK33pm8EF3yc2izHeYc+RukJfcHyt
kJB3aY0DJtYa9MqT0QWICbQ8VheUc5eK7sImCcEYaQ9fJTcrOu7M/guhllVQKIKE
`protect END_PROTECTED
