`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ImRL0czi/MTx93H+7YxZOI//gncVXBcVe7vpO1OmdQbG6MYGD7mzJZyf4FwA6z+X
g30qzOj1+WP+kVLN9RPi/h255/nTFmLggyJ2bHauJ3ME1aJi9J13cjmfbUflZTCw
xJMOCrkUxa2DLymlm5hOJSC9EDJpaIYQRDBsdZLJkU4Qh98kVXrBxFqgdtydAOwT
xfQZZ4/npQPnP5zN4RVQbr57gUceBZnUUDPoRkI5wOft8cc1LNldZ6sc15QPfspn
3p/HOZA9K/B6leTZz/8Ej4/Z6taPkhkA306b46r/ruEfR057Y56WEWieernGdJGM
aKQfPlINYga1u9LPMVctDB+A7re8vDCpn2BzlU/sVmMO7EaglWlvyB6g8V6QiBYq
QNwHJafndDAKsD2cArma30ALHBNKV/bEBWwG7ppdFuIawu6zkuhqIJdXafStt6mh
KmdCpTL4vb9P2HwkEEyF2FcpQHEMsz0MLzqkPW8tDK7Se2faUDrAe+gxA0uGVm53
VLYUI2mGP2R+wcRPP4YL+qX+0fcg6Zs9nJID0WvLExsNgKgAGb3mivpSTFjwAC/f
Mpbo/e1JsxvjVBTcmCMr3WO5HW1llSrHu/5jLl7BE26SqkoM9t5J4y4nUMTbYLIH
tI3vMIdVDohRNHriVE3A6z+TtMdkg0LxWT8rudeVM3qm/2fDonRZUdENNgP1hdkz
206yivzpCjHjfOlJo4fM/rtxb8Lefe7x3+O4GsZNU0PIFuDTC8MIvTIv2KfEVMzi
adSSlIDW0Z4I3oVDpPIIMnCNZe/CPVJqHculeq5KPONk3ouwHX2QVHCA9OM9reGp
sSI0/wtRX03AVs5/3CmMEW//IABUhK+yQsWvZWDnaAuvxmVU6A8FDUF6cxT2i+3U
FWZyGk6kXWzpg5/NCthxLGO11s8vFyuNIVO4gXwoAC9cKfXenmrtxVK8B9qmNCCq
q8NydWhKAlTf3wTympy1nTdsPQUbos5g4rmD+unLhOAwp5GzfgvbUEg+iO55UQgF
wKA/JLqUVtq43pSNE8CrG3J6KLgaIJrYhEYejPhr4y69cvX1wXz3tLyLzAnX72Lx
84LbfQw1UxY9V77TShFrnP7FFiaI7dvWgLxyJo0YipA8vzA8mNOOjoP2qRxzEACv
o2omIHbK/1Dnb98tcAEfsr00XOxyYIop97kHQj4KB/r+MB9AZk8et1LqppofkPzD
WHVTGGPS84HBnXziFbgqhmgshEV1U8AAV772GeebHlp/bJneX6s5yNdjQsgVt2KE
nl8vRMjZCPeDjbqe5CEiDniYhkexQR5vVGBpDUGWkySRgCI03tcM9Kr+7LMYh2Be
mxYUq+g8CJ7Eq9dvEjLUHYnzPau2BH+ELT0DWQEQ+IUaOC+0IA7EwtNpIYsvfaNW
xcjBVt9JYMLAmUZR5vVnpcLa3kEFQdtRXyz1FFO01OE2zyMNyoP0gFtj8M3tGRae
wbqVIAljLdJo70s0AysCsm/OUCwrHMMXe24tleMvPjzQ/m4eg1v4Gfva3CsM65qP
lxdc442WFzlHFszFx4gbOP/RBv4nA4n3pNIGDuUwn7VzTsJqNLgwmei3/5AZLTmH
jnsgzeD8JNmoFVYTtKXiTqDR8mF//ZCVpP5n0mMCXDo+5eUJ9HEtRAUX+SEe6nD7
ahfBOnx0lZvLLh+Zd/B/3aVllZUJ3b1Cegilgbm3hwn+0CaLHTCkveaf21BYyVMP
yY9lPtCXBf3lxW8n7WrbmX+nZqY848ZIRfPxRSLarIFkMMWSOlL4NL9caRLCbRAF
gbR1jZTN/YoliCy2YsLXx8jLkmkxxXOGpEv/k/iBnCiRMKaLRq9RNUOcWBHbrv8Q
gYerchvGrMnRlOUiLvPT1Y3O3LLmnUrlaVdcDwDBZiaNnFdfpH0HUlVbFfRI7kCZ
wQnwtOnzcwsr4KsxCb6e4HgC2+grbzO4l6NwgepKTFlKP/JuaPNaWPpK6dGXm8Iq
MCXJDTV64gvQJvhdht+nzJhaaTiDjFfhuVqsxPZEP5FCajPoB8bklOojP1uLcZnh
cWxXqL21dGWSYnsG74vKQVKghYzLDKlEw/nbCqfxJcd2VMeztk1fFzqMBJIdnH0c
MFCyKKBwxaJzNrzJCOkkzCCLx0hjMPC5wygywSI8uNsMsJZyMUc3epSSg/6dbjMD
yEl8aESvHtK3V9EEUBXGykDKD7JpDDqJQuXQ87onERf4m9k4oqYwKUckWDRm8Cjh
5cbbPkR0eAo5wnbYgl9N49A9cpmiQG8peOLov3+vSvmm2sJzy7Drk6KP9peC8IeT
oItxFEam1MGeXGt38VRSvlMr90hr8Z9G9WDN97GXIv81WTQbfmx2D/nkBsVbLV+I
SseToJ6DytKECrzYDr0zYtGXGX9QNxmM4IAXDPxSObeik10FYZNTTs+Bm0m+Fkh5
wqRYQtXUP72NYM1DMcRRGKAF0mFizBny7+eTfK5qFLtJKAJyiqRnULO9gbZxRrwf
3DevpWG3zdkxtZ5vh2qMlA==
`protect END_PROTECTED
