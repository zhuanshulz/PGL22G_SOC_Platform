`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7XFewMylD4+2fApWsHVK7/TSF2kEtwWa877afKzppyQNrkX813/+3v9nkcvrPiAL
9ZFNTl2hwDwIyTOKfy9YXFJYkJLQD+nGfxLsy0sszLXw3gzvVG2aJpNcsXE3krhS
YkG+BKWnR8A+ebA05xRYXmekWqMeSCGO54wykZKW+1iUiUC6qLm89yK3NLkP9pcf
p7hOgfaR9fGXNzcGT6m+0jIpBlrZ2YEY4qms+dZbZ/YDXO7TjJWR/3v+KBacEbFi
fGC9OZ2yEtGjIIgAhJaZikS7ZTEFjMJ9Z1GetOyDui68Ifli+uBwz8cHZuWZX9XL
jRbh/3/uCjkww+6Rbu387D6ZsLA6l5IYh3J5Ynqug6F6vV4dLvB+g23T9rCcm7ut
XWUm6EQ3hS4YgXQr6EXkXPUdxlidPy1Iyu/95PN/zyP/GR/i0r8nclfq5b2qOFfO
RB0o4RoDQBIo8oxPot56fZX3H7sE4l6L+yZzr1w2XsACa8fYM0kStYEm3c+FFqfH
dxPXEZdEHmWT2uaE9NR3Bw==
`protect END_PROTECTED
