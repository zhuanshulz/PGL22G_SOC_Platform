`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E7SuMR2/BLqnx78RZ/tnr7AYk9r2GUmrzm42c9B+neC6FWZwAfukhks89h8gp+sJ
aE1rFAFrF073OAHXk24LlbMu+Yak62XRynrU1pL+Gq9Ff319LM3azTz8AXbODbdE
xELCtk8KqZ4CVrs89NoiiKlXvoYk7JPGt6l7oHkCwr5K75mtEDC+y2dc8Xer7BAO
TRs6WSpZOdDFT1Bi49sH0H9Fn3CUPqaSiHRV+zXG6j9cD5nG5vMLf+1i2siszpQ+
8Oq6BCGgYHR6cpPhPnitp9XtEEWahrfd1BwKWt2G9aij51iHgcM6WMadEZZX0TMV
9v0voT8PsFJ61zhIihDBCw==
`protect END_PROTECTED
