`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JrteeKYuidVRbu7EKts50obSV3BuQbqbH2g3Q1FYAb0buT9Wn8ixXiYCZ5wxm23L
FZcI2ecyW+BIJgljp3qhdy4aPf962MI4X5cnP072afjWw74nvROePWIM5SxXUpaQ
aANrFIW0Q2x7uVGkvUg683A2pfp3F36gCJXmUd6nPCPRpBsPAYCUBGIJfAVxTvdv
SRED//Brk1e3ZLcbuHshZIyTB8su7oRnA73D5bXOHK/gJOKGbHnTSdhpyhtDHWPs
b4KOlrUA6B/jVlkUvD85BaUd3i7MFVVcirrKzwI2sGIRGJTVG12nD9wNWafDLWZv
aPm9LEubvsULpXIDvRB2jRiMuERXvyxZM9yB+vGdx4e8UhuRpN/gtC0oip1U+0tS
urTCcnYW7IXGew0AawCH2Z+zkWqhqk+PknIqBOSzXZd1np9U7eU9wtzlY+5C03H1
XfPah4zmhMEqEjHoxlpP779tu+CXztw4QWO/L6pBcNTAXhiJsgAAXtcL1n75WOcf
/JSfYK12aUFVflcnZjt5+44Px02JDIw/LbmioCPj6jHc3BLQcGzVx/C9vUSsyvNa
eizbzgC0z1fLYqQOXUwXNX1Zv9qwltwV/6VV4WCtiDZd9D8bChRJuXZDbwvJHcwx
k/OOnXE7YaNJC64bBD/fV9J6BBHYjIJPGZgokQY3lB73+iXPIdW4b5Vu7AOq0a0Q
AOE0Cgc5dgWYA2F0UD4VzJx+//mk17wUybfZtj5V6C49tDqqTRuqvPOokNXGA94f
v2KOvVSbePRWo17PdVfstQyacTPhCUwGQlSt+l9iwfYfqJF+1Z4tlYXODihgnb3u
aI1uA/ycNPm7cdiL3OTAitvA3k4sxy8Kcyxqlmfe9xBn7Kx7KyFgjO8/1shnKHGf
ruQ2086zd9+r3kQ/r50wx/NInax2Lc5tyn8CwdpmeN3ZQ+x1KTUe1EFaNUtD+bas
RGwRReyUOZj+I//9KhBOu6q+KRhL/0GhJurrH/jviC2brT1nYPKv14UxoKZw5CvD
OaTt7NeKIaruhVbjZXU9uTDdUnGVVcyXrHPvH9pRvPJ9jwcB3RE0NobUGLTRsoCA
O75SkrwUTm5nlQd+zVh5pVZSyGc3c8ZvLsbRa7fqi4ay/abwLjLgMrtFRvVeHVFV
Ah5JZyyP8Klpc5kRIemhPexA8ttSV4oJxfu2LBoYh2Ok8EiE/4vQEp+g6c6UvhZl
bunlaDeQhJa5Dkxs0XnTxV4BAh9ncIXezSIW9Z5vXBfYFh4FtmvIOGOklPu95Mm6
EOLFtpHuaXpVkUO/96B5+GeR/L2VRw00vIjkGjunH+dZZSqpfROg1ixz7zF45FHm
ZQ1cDL+LnLUafHzPPmLqncnT63V1lFK7puQj/YqskhNP2yQzcimysPtTtK655fmD
UIsA+3Xk3NcD5yayKiDboNgXqqQEZgwdAQVTN6iL2Q1b6xETaxQlA+gMDcnnhP+2
vl/+qIjoVIl+klXYNlfx03pd62C8E0zwoDX3XAXHnChZbAenRF0xsCGqBUcV8GJR
DGK/vriI5RLz6ke/CjViOlmH+ZgHjYPslP7yl17x1xiDcz//chrQevVKHoI+e+Lq
1Eb9JTvzdfGlQmNkSw2r4vrWu3Rq842ubJNXrKyPMp+3m1bHPL45b85kbnwklMUm
FqknUDIv3VNq7Xo2+a5o2Byo6kcpqw71u0XBmx2gN1QArq0VKsuHnA2KlDjgz2zS
`protect END_PROTECTED
