`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4CYUlBbRK7DFKRUWiwP9dC1DkXwr3uHoWKPTmDd2swc60GSRTDkFWbeDqHUHS9EG
xTxQMO2MFc2woGKrrCQg7DhxxN6m7hDD9BtWs28AqZ17jqtkfGncN4iAWVYmBn15
9V+65SPjgdOKTmSKpY8rO0AuynfsD+1lolJm+JDGPmHP+ux5N+ynP/P/kGVUbX/O
eQiEZ5VKF+ViERd4JBoFNwRjzNRlGdKiVOROqBagz3wDXeMg/9R+dmx8uA1eW8ay
Edckdetzg5CLP19l0Rtn0Q+TE0xNJDC2ZQsmrRjtN4ldlbQ//G6AaVubbVjJxB8C
10RUL9iVptP08B8LEB6f3sbJIfxyeh5R8VNsziSsQR97XbHi32pci3x84UAX9vlI
Iux874u9iUlBPOKE/ODgTwxIH1DNvZy/os29tFjA42Az2jKM6DI6My53wu1I8diB
RNKAUwYNOraVFtszPSzhr0KJF3rwMsRt7Rpnjs2QaTRpFDDvXDDRh9ebnA36tpZT
Y93xuYPKeOV0YESuDsk0P1UFzFFXacKLs4X0caLhxsJ2Vq2iQHhg6BiUjlNIcqFx
0W5Vt3Gho78UTz6jSj1nbA9IQU/CO5J5V+k8brq3bSlwjtxGTDxAeNyRxzIZstlc
YvUOV1vZ3g3LqWUOiKz3FzxNcZdCxvTOR4zvfd7nP7mWo4v0jK5UfbfDfrWh3zQe
jsrwxKysrubUTg63IElO3cCCLqu0tDf9s+9sjc/b84TG4wKBDiUdsKI6aQZZhsMP
Lwryou5/fZDmQm7s/lKkEBZFnmfh/+QUp9tw8XACzGfFbGYTp6TN/kaS0UG2Wrak
b75JQPNybPC5G931tVmRUS58eZDmRHbGvNniNd5xoruRSaZRsUQM9NQ9oqBg5iUC
eMszWQqIWEPLz7b5t3ujBFSYX3IAsmBQwHh9bQlOO8Ft4K5njThaj+z0dqzgi1bb
KOsPtaN0GokytRLbJJTw3rwbL8fCYfONNJn91/4lCRs6AG9sPg3liWLFcC2A0eP5
7PCu/g/xH8vpcGYIv3zQqYZ55IlnQL32pWKrrx/7HUJT0v+i3E2Iuk91PDLrX0p6
KGBtInI2C8JzYbOhFPofgsqCrz9N0OStjv+k6XnELdGlLUIHcBhmwXMIwEO4gQhy
XmZaV6weXzm06s+KDEJ3ynhqOBvsO5Z7WWk2VPeJ33LBHjXGv9SrAsjaxbuTtQ9m
nmN9ZwP7KjSOsrdNDgMmPRco0FSjT9iru7A9fv08TGiDk3gTfdOsqmEFXKF388Qo
q/5NeELFIbyNwQK96e2Cw8WFOIENdj+jCHJywnHtR5S+pPPCqqMfnHyDIvcJ65qV
7XoJdzTST3wvV/OuXAfePiujTRBcppvKmLplJh37HgqvFK5VsZ1Zf63aHSCUM0KZ
wrgzIGkxf1tgr0RgG3yFITmEsvtgrtKhmM15fnWbu4rmSNq52ffFFPxL/Bprjp+B
czBZh+ry9IgMcUdb9KyWNbkPJRp4yN/S5oVSh1zs2QnsQc0JPj66Pe7Oz1XkMKRw
n62EDvWw1qbFkcUviPUb5ntaSVzkCuICRG9IiKTpTm1od6RGKI1kUI6P+7HoouQ6
IRR9pRqNUCryEAFp/8nLLDyNx/0hWkBzMrsEHRDuASAfsVAZs2TNA7uQyj4VtFgk
EghG9bgfaxJNvzVWU0XAilxvQ+XQwCMqUfoeXz0OKY+2E4q+V/cvqtfSoLUx27q9
6rWgHYxdoNPbJ1fSaUUBuvz38BIXUQaeQ2s1eXSOLTAwOUxMwVqXed4YHpkAgQQI
l7oCe0C0Ov8n1nIBuJLSm2gYblkNX5bdwEFha2Gk1YvbIiu6Lf/LSe0RO38BBWMA
nn1hLIWng+rJL2U3xL56UEIGMPVzP2X+lnnbpR6OGclLPTX2Mwrm8IF4ANMMM5jN
FOXHZSG4eWIdOMvc3Rvq2J+Fung+gOyvvvIDpxX2T2Yo68wxN0te9VF5UzKX2mv8
XVjT7vod10OAGWGPZ7EWadgJjz3JGmE4aa6Cg+CB4HBaSJawforY98VPg21YoPLZ
U14i5P9qPre+vbIdXg5wUSKeuufX+Q5HCq4fMwen1yJBMD2AOwAC8ZYhSBxsG3lz
kBwTYsMwyvSCekofNtrBHyvn96m4Mg8Pd2XPinrEiW8pMXPfHZ//eZ5/SKEzWEtB
UhfcQaWHbyrofpIskcu1tMn+/SW/8ZPZNTmR6skaQp/kx1/2zf6atHdPC8NHQX+p
sBnzA0MnqykdV3KI0EJkSuQcpYsgoefqV4qtsSMKMpsv3/4M116lnKe4U6/smCqD
MPRHAFKIoTRhJ8N+YG1E+uTxSJutPP+s/egmTEPKmlvbEy7SrOJr4rO/cZPu2BZ7
kTfIDt/zCv2zKMwnaFEnCZ1Ejt9Nxjtk2QeS3ig87asU6RpEYU6Vwt+KkRCsuIOo
Mev1LiCEt/hVcrJ4pSiRmYut4Vvgh2YGx2UEgUFgta4XbcJM1x07g/ZTd7D4biCy
ZskkWuzoBlVficZznKfwLVjefRPlYAV005u90LO4KLTtaQOt0txFonQm7VM5NWEC
9twtqQ2qz+ymAcvR4ew4Zp3d4EZ5ZJRwzBj1PqM+RrY4yMtE3yJjZmtEewfWSwqj
F1LAcKA2//0E0gG/hlv3IxsXSzzkeLwAo61zD9SR3qthAmQl7RPeCxfGOYVAcdle
2iRPINLpzY4K8FdU9EJUQzsOkPXTUBqklt+IrW/h+0bctlUDn99jlluVAfGPs6cq
W0Nz9gqARxBr3sJbRzOyk8NTXWBy0BYOTcqa3GFVD4XXRHehTAgDMEFUdyh271j4
FSEnq1tI/YT6j78REuFhLhH1B1Q3jU9ptmgaErtA9S7S8fIldjcWA6JuewBow+iX
3Eb5NJfJtlocecNuZL8jc1LrdioJ9H81gkGKC1ZtY55BACvYUEh/YgF8SVv2WNPa
eijvXpqD7CDKd9baudW22hgmt+I/CM+3/2F4xNZ5qYkyOsoM8/mCR68qt2jc4OIK
tovptdYwYzR1fV24u4Gk5sYiwdkCkK9tGUaRr72J/M3ieDzvnhQyL0kQ6ay7SfFu
IZrxTnK6Z7W7/xjKAj5WaT3LFrgnDcBDkY7OIZxU0PPe611TyogJDvWBuzl3wNqu
i7tL2pAGYe58W5/XV04Iu2vmObpTj6LDTRUNppA6Wgr/tgBiAv3HLmcuxc+F+y4g
pqyNLhXF8vKIY9pBxktgkPTqfizOLRxnyPVKhtBQBxaGFuLjE7ovX/XFpspOQjXv
ALVOQ356JTNSMxXo8SqNlaES5zad3QcK1XyhCIuLOqvtTIAz6mbmBX8GYMOvhAO0
B+aAsXd4CF4GVPEfTuz6ykMqf6iuGNdr0PAexVcs+9MAG5c5zODKG/fQg1crPK9/
zs9VmqejGWrHUXwhQQ76zQwQ7sZB5SNM1LWkG3SivG0HJmq+mLN0Wa4Ozwaro3mX
VdLiquqiYwEp2t6SDrQ+2I6SYfi9Wc5kRD4mXeCiKVC/kv075MhA1DYNss/yz186
nA9FJPfLKkjLfJrWXlmiIR+SbJD1hW6eJG6MiCSxZCDq2KGEAH2y55HRRtfwQZ/Q
yiM31V7EMHQPgvQIpS/8PUfHmiJytl0CUqIVmH/SlMrywO4WhzGxDEsgsVMOVtqy
7RabxNcb32dbtmuSjtvxIwZbSxtSWNwgb9mnTO27iN8pe33SxxFMQlnt9jzev8Gi
/cHsFwOB83Di0XS6Tcg0PWaCda/uQcNK2gCiX+e/WxUM1pzB+oO0FA+EFr5vXyDi
r7lwGWQbn1WrfomBcZuBVs6fbJ1xz5izFxkr3NkWy7KFh97bF9m4vZi+QTH0hgto
CHRaU6DKwrOe6h8hoXKKxOvQ5vV8vkQEZkIZQTjUIJPbe21qxE2KY+fRjeZyjt7W
ffvKdG1+mGurSEMV0ZekKM/+1Ehe+1fgd/IVgTrAABQL1XlzpJSR0TSyqYPCU9eU
5ALBDRjtEX5dJWzz5s9OuiOFop4bx48cv6t3Q+b1g2rmScbtTVQsQTN+XQUcHPMn
1nj7uJ5INdOrgLH2tM38qHrpEgfk4BARPasLRd7Gp2sbRCqkDa1J70LFFHzPY1pV
bXxin2V284g7gVRMyW3ItoeR/tLalYvrna4ktVdn20CM3DURC3FhliqGNiIXoUhG
oFw9192OL+KOtcT0D+o7+YTOfkMveVgb60Y8uaSAMUM4OA3eLy7TTi6wRd0hSHr3
2Xhky4sqAp2hePahfshIVuwLaakplTyxOLZ1qVjQqiIranQov3LqHpNweak9iqrC
LNY3WMVQgDj+pBXSfEPlCzdmgbTNz+9L2CfFFVn1xYOnIIru8M5uCjGUXvDr6NEG
SxgIoe0rl/n0TUKQJ2KMLGpj2arGauQW64kFSpMTjdmYnROkL/BKMNjn/81noSGH
dTrb4xge687mdwN3V06//EM2KzHf/36gb4Mh9EweD8untm4bmq4xJWk3DrEHh2KT
I8NF+A+3NQa54ecYZx3IK5jflBWi6Nu6kFFHKCtjJV8XzWYVvACDR2szLHrsaOs2
yifr7MrPOCtpcuE5Gu9FSfKFS145HokY4G0cyMiRvlnV6jz1grgOCiplHIU3B9Lp
GHz3GNIiSDe8sSqwaTFNVK0MG55GFgX/6mx6RXNu0C17b/CPdqfw8tIH8IsFvqkg
WKfIUCNwwxqBCa6E4pjUAyHQy8koSScVLXOWAQlZfpoml3ZV1u7og16Qg3CSgifF
u9kLW7AYv4iB0uFRKk8pQv4f2VpPSEHkjzHu9BuD0mH5c+2HfFGWiRRZsPwgJMBk
/LFkr3c8hZekJ0lnHHhWVmh1XOsjxQmwe7R1b7k91UA3ig88mZxsrvldljL9sZoE
n0B6yJzZKGlKVZstHMjD4EmgmjvFlLashdVRYYczTDxxr0u58sZRheMxxAmgujQ9
B13FMIjJTaA0xj802rTBCO0JlsoAmBrJRWGLm1GdMnPOIBqtvjtH6Vt8sQMSlAjE
5UDKVaNtFEdVx8C1W4AQfxXHasBmnjumfNZfKIRuS2No906n178zniNpwQYT8rDE
PGsQxnCHxA0M2Pq03Q51//CgwN473wHG8PR9m8hN+P1cD0E14hTyEDZucw54Ift3
K0h5JtreXlJqN2xbNkevP/HAch1DYZvrTwWGPKNZTHt4bQG8opSUsVEsogCxgJM/
NmysP12i/JYQmbv5nAZA58gmgILRgvekU+82YCRtIpm4rqUW9OURN4ySnvyKCvRj
dZhUxoZBx/TlVewBuz3LFQ+h+9JDFeSqDCN9w0KEY8RKXEMzgHWA0H0FRHUOqiq/
TYgDj1bJvJfnlknWcqLUockW3WKOeb9sGFWPtIp1PUKVEdmFforKzCtCg+gM3PVN
WlfUXzuGNbCrBPXyxHpgraSamEbGKvKckeVtGcq+Ku/4bl/7Rby6/xTRLs8fcO/o
R8XzcnMJ8vRMVtGCDYcT7TvcqHfiJPa0rSGSU9lvWtiD1zmi2sBVBLLIwkwDo24Q
IKw1UAkttM10PbLJvu1xuvJfvuhQWvJHWmOzeBT/9FlKAK/23YDSiYz0Yp+huuZ/
lGTo2UH/vQh6pGQAibh7Yy8Qu/qK54t4ZViZgeUSCpnDfbibmCMURNCCx/4E0pa4
nDCYb2vxvATGxbpCfv7CKLoib+FnZe95ROSyYhTn8zeSKVCTYOsFsl5HMdWHJRxr
c8u1Meel4almRNR9I52g0fHfdYf2hPPWmuIUoRb5BRriAd5hjoHjPVqc9j0MdL4B
jXxAIaczP6ecKJVfDct+P/jZoauFw9LnmLZGfxTcoj3Tch52kcq0wqC2IMOnlDGu
w3aG5HHiz4dxC3d85jG3wrnUHCeVfECnBQ6emtW/nwsuK/0Px+jQHfwCQHHgbpAc
S/YWTahWxvGk1hf5UWm0ipQeSay0qlqKKY2IOou+DfY+npC1wFBFMVPgXTgKTDI2
dTpuly1si8kmXUp48gIebtNAEB4ZVdljYXktYrGXyaTMdBm7g41+GCPkiRKkgrXH
2bx+VnzY744Ylf+ZgzkawecJvzawU9irEqyspbYz638n+PrQdEyQjgsXX6Np5tAy
7zHn2m+hDnocKs/ecz+tt2qAPsnqkeUmMzcWUN9TVGWZd0iuLnr6mUzzI3Fnwyyi
HGWWkscxnBgfortq0sfDMkxtSceFoj02wkd3yGkIrqsXMls+NIoXZjXIrWe0AguK
crNds/eZTXdEfwx/MCMCEtT142RcB+qemjbGoqMKLtpdSmneb16idgg3NDaaYJo1
IqbIE/NvBsgMG5ii0bqvshxS2L62UdJWx76qjhqUznUuon5Botey0bqAwugOUmCs
8WFf/h8cf/VmPllGPjpaPqWXIhdKI6PvnuQVeUSQ4UOwvfBT1bDdYgFlpFSZmBNy
SjUYCEHKkOjGVK92w2fH1Xf/GLzRdMsmxJ23LptKK6wzLq5Mj4Ke27tlqGQ3Kwd6
oUFTtbcl5h8srswhZrW9DICM64irpz/YXHzle0ksE3hVLchEpDI5YjNrL6BENc3H
/aBWVYwYYqO5e7wIZnBdt6SOplQwxrol4/VJw3ZRCVJ+xCj6MtRu+mJQgia4xG/F
n9KEGDN3WtKzm9jNBASdgaP0eKcqPFoMqffLlWOor5iaZxflIMOd9J5WZf2dgkGp
O2LCGk47u8T8yC0wielFiyKwei/Iyjs8xKWMx3TPyAiCQP0kmFR0nzxRqKQ0Wk9e
6Gj4yEIK3JQhtocTHpWPdnkMFHzHlmNgPTJbzJ/QpswvIImBrPBUsmqKf2siGIX+
rkjNV/oJS8jDQLQslxAGJty1Z7ovxHoSmR7igpdKp8dI+sEcZ1EuYHZHgvIE7INV
xjZV8+58uI8ezjS/AthxONCqo0DbBK1KijlKQhV2s8ILorZ49AGR8847BCDsw+02
y2E+Hy6c1W2+4guupY9tNU2qBvCFC+p/m/4pBcNAHaJUyzDWtV+cW2Sy9aqQIogH
eGSHU/XLuptv2TggHlGirVsAvcGfXigfgUqmpn1IJXHgFgUJ41U/eETqSnl0iTkx
NwtTqR0g/6qb6JbK5XfB4JBw+MI+vvR2h0c4umJM/5cLnPbhB9e1uTz020s4qOwx
2qADaUjQcxxRr7T6yoqVw+aFAEHfj/1xPQemA9LrsOhJsDR337ZpHFyZxVeyrfeb
vCSo/ODKImbZjmfaQkJoo4eJtuQz03Gje0E5WreG4Y7zjHi8MSzFT1tNcc+kiMnO
3M1sgmLUytsrt0LiGrazp2hKpTubsEoJ4ApBC1LE8WlMzpFDkcGsdnK4fNgod8x/
bBag6LjilJ37PXiGSEa7fV658c1FvjmaB3gu7jg+slX46VIHraSyoStLdxsJzk9w
oKBOGJ8Wy4vqLcdgzD1dq/9xZMB+rwY7G+VzloWIZrttBAevhFBTaweYUFYF1Egb
BJENbH+TeQ0Cj8nrbk8gOScCTcM1o7r6RNF5hAWVOo74iufsFFiVHNjxiS05gFaJ
TxE9Bq3Jy9LgpKzv6u2vPt3l0MpBubV831YEdDvf0cdaR3wQt3sz2zYoiRUmUP8E
LSaDaCBCzwIoslkzoE1VHU2UjP7SFdBQ4DjGMJ5Gz1tUZnORmXgF79KXs3268TzS
RHZ58Ng39yPWjSD+8lXMcrkNpYPL1J8RYf+52SmOwgdz5IpmOKAfwAb7IDnUPo1h
P4kmXgSYRGaE3C9M0cKu6A6rfNsvMjCmFwa7314S/gwNabB1b2vJa+qe4UJmN+Y/
YlB2dPQtAooXYE5eMqozNvaX/eeqxv2tpyH33Kgf8lN/E+V2NMYebVxSmbeDDYHT
Z/ypkiRZpwB+DBUKtO+pPzz7S5Ai1tObe9/8hKlSnEkAQULSE2rKcYMQAKgsQreD
LCjIdrdyEWE4ZExfLC9iea8qCCnitLiYnXJXjLlKE9cSBCbYjj+BPpK+hS8BfGNA
7cf/HpM2J7xOUU4DAVjnyZrJt60TLtHnPbmE2i22Am8JtgjNnr3bF7Fa2p8OUHXp
qd/RovENIPuj/pu2S+b6nqbr7xdMBwfSTLnGFrkE4Jls4/4+BSTJuK5zM5cH17xz
TcIRaRC6Jp29Zo3icQiDrwUXd0dVqnm/S+zSDNsQ5R4lYSZvJbnzcvNukFDvwzkV
PA5i+i4Qn/tfKIS/6lbbRFW250JPmNvL77dnh1iHkjnH4wz4ZyTp9brM5dPIMLwI
K37Wy/XoI9cwZDK4tqsXQFVAiX/VhVe44vQx5K3TAWoJ6tVuiZV6D0l0nIklLJ5G
Izqw1LlZtNxuBwOxHklPWzmiL+tZAhT5g64bYQ+kWtW6OvqiEtW0EUUUMnxGJxj4
RxJE5umQBaxn0qkdjIvMj79cqOMOjpot8YBPu0f/GHSnfwLK8+HxCjSjjOBcW+aC
cFB2vWDYDh+IWYRLwS3rUi30wyyLZqPQEBfUU3VYxafVLJZzjcI/F6XwLMJ/vYoU
bOBP32wrY/WwM+OpqlrXor44EH/G83sxCytqKZDRb8FYC7OKtOiXNXDy9FSNDm1m
obfMLj7/iDu6MPTb5K0Z5Seq9ZeAzFmVtj0mUFp3OhdAuH+XnpSkfIwmabhPnjBe
92KPsZzmFUzz2EcGjZ/AcqyIuvMmKe19Q4/798zFwbArvCV6b4kiSDw9GT6uA1g1
I8nunMncOG2cUr6DmS5cMMlYO2WfD6zXyEJY/eJI2oCUiuz5XP1PC0K2CXpRFPfM
cl8uJKbUiCKsIVHH8ZPMDQXZG4bPJXYEFLKmA1nNH6jNC1/0/1M//e632JY9nRah
zzFd1J0FXwGsiZW0hONAGKeyIcx17MaXhjNMfRoKQ2CTQP+mKl0L353WskfV1cRF
7ophviPgePjvtNEWXfsRCgU3dNnLqmqpgOTtBhJY1/TD+eH/hf6JcE50LEOGNBUO
bAm5PhO56DP5KVgCaNv3MJuBaw5pwgatxNnFTK63pZ8i2QuDKstK+/QRUUnWt3q2
Nmoa/MTJFjx7xxol1OGDEZW+6kpSg6Vt2JcKVI5uPEkHrakaokWZ6d+izBktRnkZ
uG/lJINsdBB3OMvaOZBRsEadu1z8ChJSgm0TBGu+cBQtuH1bPIzmrwoToPUPTYRB
3ES2quUTDA45+Ym12zf3PzSz8feht9Vq3SdvuUDzHVYGHaAhCNdb0OPjlSWOigAS
sGV0ZtYZxMaFrE88vqNE0XKnX5UTAirxq45JOT64zcAhzYUrgYKWY7lLeQAYNQv8
xqyRaA6ewR10xg3/pQ85OsOKRTpiWMv/ja6CJLHRaTgyUhqIV9E06NJqs8nXBYc8
IGY+9qkSxNKcFwf253z8D7/F2scqNFwNnUnot5Uc+9WAxkXUNJuxzy0EiAg05Ejc
15nkknv3U/LI+AA8PzUomldyFOn8RhXHnKZVKFkVyew6dYonvpmFJE6IIO2SgqcD
BIahLgBme56VPj+3jssTgtbYsM8AZLhlFJOLzeG6vgBzBOVJJnuULkTiaODqqmPK
jNOj9x2hPgDyaQYyKllVIrPrD+ZUaVkOpEpKgne5f5tIeRF4EbfgV/otYvjN/i6u
DrDpzjkv/pW0Ex1q5shHfnWgxVfe5wjOGyJb8Hhp9fwPoCOmrZ6gst2V75hwcrmi
Mmscg6Gru8p1qCVxwpn+93eByHFUOfWqBnv1jFDxKI6SKS5vyfb9NhA98W9gNOiS
QuhOQPScigczGUOLw4SzdW2pwJsv3vLvi0wPS9nq9GqzoBZSsX1aMR+hCkLu349S
YGw5bKK4BebRt3WpKhO2eOEGhSC6RoIBLdhZQvf/BSl0i6/j+NnMJalqvP1U6zTz
csaGPGyX3Nj8aPizC1xpLGyTOSJik5yBvIGH3veRTUZ0qWK1suHRqVYCjeqp2XV9
swb+h3jWrLBvCqhRll0PCpdTlaO4iMFa7o88bGSmVsPrjSXqBt3X/ZhfyfBRsLce
OOMCMN1L3ILhVxayIT0Ay3JCYimYd+ElVPTvsfwS+g8IrBiGUKQFPAUSJ+KP3Uxe
vTFpqPteZhULuJd8GMCAaaTEviIz54rJD1Sw61XFNxobYEp6gL753+NrHNtT+vnx
wiYAQAy2DKOipm1k81kUpkIgygfgaTuKy+DDlwYlTPVm08clnHxuC3M2gDU23Ljo
ETXBf5rLHFMDXjN4NDpzszcknNSzd4+XEqEppRFmzEZ5dbN/E01VDvFsmgvVE9OD
ZH1JtmBM93fFuy0rI28qvPJ4+hj4pcSp471AbPqHK7sF8MlVsuj+o1Y/ONQ8KFGo
HOFW+/UiJyyVcj7vD9jMDbGhm11RbxifUWsXPAOcRoMAhSVjYOl8yDxSL0Q7AIBU
WOkWwqqc1/PmkqLQQAo7HEwfbH3mQspi82E/OxNQ49CNucYW/HeSQrmcymbOQU2Y
iZiQpkF9mFo7FtSShzp7lttM49LrGHvTXydW0CaBNv9+vu7MsSilqL7pmDVJ5p+z
4Zhza5xCNzsI22eE0aDNQhhLcZTSYoL6U+iktR+UDsoGRt8NmL5bw3neuqwQNoVR
+Wqd408163mFyNzQ/Emo4D2Y4n1ckCHom6sXRO4KJgHtGE4UasEysPfiplcnyVhZ
CWQ0oBM3oDPpob6J6BVj3mNyqfC0JGsjyf9/4/lwBoo=
`protect END_PROTECTED
