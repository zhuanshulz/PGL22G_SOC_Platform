`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Z06UsfxK9X5q2Rg1bCm/8DQBwgJ0Inm7GBZSvHnc9RFHp9hO7F5cSk5CJE1Ptwz
qvP8iq8FC5/lV88CC/Siff+nvFn6Hi/LCbk1DZQfO4eNnN/SwCAmNcU5c+z5Z4K4
Ka6GobKpX+DX0SWd5DohZnl4N31DgwVM6In7h7F4OoOxwWS8xsgjgdv7vIQ46dSH
8Lbb7A0tJvtV2+z8She+CRX+ExSTDAzmTWDRhwIk9qtqFVjj3iSQJJQTiBz7WMgz
typh9Tbhl5VjY/3xSgpqgrJfRpjfAgq9vg7fTrNngG5DK18DGajcgwN6sY7+G8aD
KXY4GHuzfcSY0nrdLF4fc1u5SbeTK8meZy1kvo6WvHiTOxAuYooy78HZ5cyt3j1h
GRsU7Lfli6zmARI8c8SfP4n7BW/3ALqIKILKwp3GRZD1zerqiLY/If/lPPIY+TRv
vSbnL1ER5Fk6DeKl3F2wMYS1+qIyb9cKbmHJlnTtrxYhoPvN63CEREcGwYPKvFNi
bOKvP3pj3iEGgHsJHHhBQlk9Mw8VVd/mya11eGYbPsJLynDOkHkBriGM9EBFHvvD
oeEwGvM50FN2vN4LmMpmPwQtYjLxtZzJhC4RifbnYT4fticfRuePttCb7MRY/2DG
B1UhUXFkeMtnORElLN9Rqhz03lDiXtqb11R0ksw6d4xxMO0PK6Nhef8eBpzrWpWF
q+498csLsicO0tUNmOTO+eXGH7SafQgNnfH4I7xsnsJNeKlFY8MVjQwK3dajLowC
T7x8iKKt312SMtaqVvt33WiASiLbXqjurFX5rCigWLrReYP3aeh6aA6g0xtnPe4G
y9tybSlNxVOBAe/OZnpUAhD2c4tb+hAtgMVbxPyrMsmTb4wdclBRPXzZ1BFJG82C
+tR2s0/Yq7jizAYdW0zLORZUgLGvD3h1s4gGsOep3mW684xzhW1iZplYhtOykQWp
OrLUFzij6feWMVUOq7wjO8z+XA+4JR1f9KofXr6sEVvduSvEM5uNuewqW9tktAHl
F4sC3EQePqc62iPsfZ3U8h6JFxIweG4+5RkBEdc5upBuPGU3WuLlnIAXF8x7kva1
+5gcKJNMEbM/mpGpjT2f5sWWpZyX/limlZNEEj1hFDUdU4LN5R2IhLrkdZrETnUo
USpM4+pTL8zTpDYBREAobbXFL7bLqS5xlu731Rl0ig9DnJ+CwznE2ZCEb8J6K2zT
zaJPHn9llVCriGkkJ9iY9Mu7/U60/M+1PX+ohJ2BCXxkcT1PHC1h2KsR+DifAE9w
rC3+uUX4z6e44IH+3qjNehIZuKmD/WJZTRoMqdHV3vZkBPyjkY/gWAJJiq7IDLUV
WWmkfhHaoXIDVhKfvbAWR5CoxQhJt9hqZnYqrb6UVrz9XA4JGRuBoHFttmImX5op
TxgioempJaUFN5sj7xz9Qz2vja6AEmlBuPtCYqbiDpDnUkMMNy3nCivoodmAmVVI
eSe/3hEfbC7IylFpgShXeBqtt/CoD3j+jNGIy0kdrPr4U6rEKxRmOSF7ZWb8/g8e
loFzbMJaM11ODeDeNtLODVd7RPM7JcU45HA7gHD82NAbuX6UOUoposRupYtlFtr8
YWFMIfgqTuXkDdR+O61KcD4BQBM74gHdfjpsVLhVPA2ICOeStWcNarV1etLYRVcf
eb8a3s0ZzGIMVunHnct/5vRmYCEu0Eb85BOoUqrWljoZIUpRjTbCXK7WQwc5ypT8
qZXLUgNQn/F0kmdV2f/U2suJjBQUmBBLFezM6Ulm+oseU7RRDqpBABiyxpZH/WYw
9pTnM4/GsCeenD9yUo6yNww07HC2KGbLuE9RX3Jc2XXatJZIej56mw0J6eNs0/4L
ypXZxwwoJoBAzSozDIjAO/gjliZeShWrs53x5zBphCZcx2gaBSneSAFXIa4cI9J7
cj+fhDBaZmdQax29Z5T7YHQxxTIE9J7RvUu7rOy+s0OvUnomCWtfY6XcgYgaLlDS
FxJXMHoW7xrUJUQiS745zgQ8SUh67mA3HZI0hL+ZpePW2nV75aJW+o4MLqKsqx2d
BVhj+eiw3JDE+TmRY7rEAQVYRWH+IxaCL4clo4zR/8RtNFxCeuHbwavuZVcOQ8v8
GGPLn7UG7ZEbrS4FVIhNwP6JOVl9ETyIQao3V+9MyreIKvwaeCgRrFkzv3so2rqQ
np3x3WHyil9HQBh9AWFdBpLU4hGsFooXO+FxTMlujLrhQoqLf556X3yODmHkjfxB
yhaYJq4YZib349EPVr5RSpH2GRlauYBjJw5mGMiN7nQp+XpOnePETQVH5cbzjsv6
Y8kceJTo2U/sXHAMYIEQu/SGdetfFoX8idjmiqNJ3sTx1uryz/ZEZ0a5AokX0XMc
bYndDauNIW4ltUBB/4Z/Yq1RxEKI5JmK7OsHdOioApz/9zFxOI8hmn8UcHyiVdb/
JkT/vqRbtHIq+zAS9zd1B2uvXqHU70lRjKGflU3p1Wdu90l3i71Z8C+jSb2HlBMd
6y5mOhS90fAFqG/7H/nUekA2BvHqkowxM6F9WnWLury1RJkhGoHqouoxsxwZzMvl
pPi48qYVTnqvW5DG5mX5UEh6uc1eKEAClputmTi9Mm7PDWXFxO02RMXJZEAaCaWM
zwYY13G++/xQjt4HqTpPMhmernm4m/gTH0Hjrb1rE9GlY4qagbT9+bjtKgi4OUsb
fL0feJFkRORinIHrZAPV4WlN7NJFC7y59fWzyaiwsH17mijFamAFCZdIbn1P74Lb
frHXCldIbZGAFPSwZXoBtN65tenWcKaBN3iCdTRwzfPF48ste19I6QcQ5j/p/Q90
DNtIM4VHz4gZLK3yNRcIWzp05frIdwdYpqutIPdf6aKze/hsx1vvnevWsIWCRzeP
lLFzkG2O6rWAeonGA52sXBbqHHrljTbRyvzWUoyIv2hOJQzVUqQecC3vVohD8tGE
BvsdlEjDCqKasEbJXbe78xeHTQZAcN3WxJ5wXRiLyPo=
`protect END_PROTECTED
