`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gnCWL+Tro/VzLohMmsZc2LPQqvgPJssjlV9hBE7I2TtNkMxgrPYX2pHw/QInXm0Z
GDSw9ClaUMmgkRfbwSOlyS25lbFyEZpb9KglyF/dKNEn0nWfzcGwbciI5dCWzAxu
ve8SUer8Os60m7pBtsid9cO65iDWNywG9jtaPmDQjfKGXxCeW6hNmFulch7u6akJ
pNMh234FBKGin3d6iXipKQS29vHts+Db7csqXyjlpqmbN0IG5UtXQyq58lbT6Igz
yEdqGI/8VeRyMlLraG1XrT2xQqYlkOVIoa3pa4SupksUU4oN+VmaWCtkQVmaeQGn
VLu70JESJiwjdjSTsIexZaS/raGsZmDTxnUJdudYLRXPJ6FvzmcrqSTlxOMgdS8r
NFWVgtnIs56Wx49Vt7lNvl7F8FUv5ObimTclzTkvXhS3WjfxjvYaWBoWAsQHAwuw
kfJXRuobDAcr3rjvaaXiJPmsLfZx3X7thMJfeAIM31yVhraKwnmtdTTeHdAPFK6M
BnamC++ueVXMy0i/O0OVawdWH8EuLFUZdOeAJbdk6KjJY13MzpuSMHPPrJ0VJ7qO
e9DrZhwSGH95EO4z/QqqWZ/H2aDb8vFec+dh4/F8/Jsr8npJERf+tjgpkBH7PqF2
DyR7Fpz1LjUPgR36dJDTlufXgp+im9P7rxgb14hWz2LUp11oxn2ykbENuHEQUqlj
WZLEatLgWfDRGf0zmUrkDMnlBM7VLRG2adaMppPLrr7tEyZ1pN47g6OtmOAJhgWU
RAmHRGd359F6OO2jIJM53vSqcyyCzKRSkQqpeZE9KegF2X/M/MQrf8gp/vvlFbBv
/R6mS+cVgbvHj8aBMOyEsGann4UsL3qxmXh+EdNEfEOAM6ET7MyhBMfYjvOMZ5n6
ksUXUDzk6xbiNotHY0zuTh3NPzvFIE+LDkjFL4iVIm4UKZFxthHiI0sjQDliSxKS
iQfpvaNBfTJsKUf3zcXBCViUlLGnxXJy9Zc0q6Y0/+WDjaLaslhxwyQFY1llsaZV
vwd2m6XCVycqxegmgkrSbnXyzrA+qMa/XNf3EyP6IdrfTmPXbdyt/iAi9rJLQWGi
UEpshN2s6I/lPMzjXL33AjSAgwjjb7JMMpsax6v6uJymtb7tCNrjp4rDdPobLZCX
YPNC77XL8bdSMktmxAPIK39Fym2Z5V2qucQYxwFcjixHEnmk3zdBJfm8Rqociv+p
mQeeu4haq2ecGF6Xf6DpIh3AfEl9w/j2fzr0L+5UJzhPeqpiXg54rUlr2RHAHnyf
MK+J8x6ZyEWNoa0l+6JgocoDavF5YNpPiDudSPRBIWz6GyICs8by7aYInRgkdnPd
nxzFqHQ86dqzxqLDdyqY1vFSPqqgA1KOOtL1WlB7WyXmfV+3/YtQ206Kz+p4uNH4
Sq2IB1MYzSZC0J/WbcSuD98abT8dXl9JxfXmCSRtorUBct4z4j1+4WD8vaxAbYy1
FcglV/lL9ozxAmS9PLUm3jwbSp1JvNipjZsscELY4YvNAgdvflWibit2vkTjdhGf
Mi9wkksVJF2JoroJCTxXmGoi59n4o2gjfW9bY8tWt2YhU118bPlyQeoN1kMPXiuK
a5im+j/zB8BF38W4GfR99c+ZUFHnGmnfjCGjUyOyQrhkLsnxF1Z2ci9zuOTukfYK
dkXYT0SlRcoWjBEIMgMcAsbBhv1SC0J7WAcFWKDRVpSIfqpxToaZBzaF779Tob0R
S7Lb+phiT6bYtNjnp+mtOVcORWkunKFS+wbRV/BcZqdqD/mpAmlKH+N4L5JdNO4G
zDzmWxfS6c7nTrHemkb95nOipBiOJfkT9xgLCQ7oHmXzLFv55kPi/15sCKwoDDj+
zf2tQH2VtJrDiS74Y3rMd3C+ZCzBB7HU13HKGCE6v56237gj7agJXwUb2tHtKAjU
FwSl2TTMJU4Tn2/6y8DWSvDbc3EaGdYxZvSdgEhZBmB2C4rVMiJc6j0JVx2Ai6Xa
hQpwWTrL19PX5EHU2pCp6xnDHYod3Jtx4BT4EVzDS0HMlmPoh31I3p1DT/JzbZox
TIaA8LxS+hwBz2+fNTytbiWhyXFdQXqijnMHdSHZ5ld/lmfXNyXsoUtPXVSnNoyv
5fq8AuxqEHfKhP+i9pHVLPHKlSFxK2trAf4BdZESmbDUOMK19T7ZRIIDkovP/48L
3V1IaSRPOcvxDFIeAzXZWu44pVTB97twAz2n9HpNvpNcEwCe1Dj6UO2IvxBAvn0s
2JUCOwUZQgGsikLZxRPsUXLhX6uMwt5vLIWqnRlhMTnGXs0Q+Xnv1qvO3VVmBzIV
W3hlMZt5+mVE+3+A2cjpTyOxYY8mWBoRbBLA8+zcv254wURJ0sw2PCmtZT1n2Xau
hXhOq+2x+LkN8r94XAdhGcJ+0XLJa98G/ZXN5C6xIdokbCSBeVGPvwtdYufp/TLc
vw5agk33wdo9c/WVk5xJxJUTNw5ZcypVvyHlYFg2ndjZrrc1SWC7PgRmk5NB/5+v
+O90XE3D0b4Xnjt7UDFuTBshmi8wtqSQzBn1I46kd1m/Cx3wF72/RTOy5blJZ2kR
KX6kzIHmOElLVijbS2mmY2NpIJt2Ic5cjlFi+eFVyW5eQFu/2MxYgkXPBDBGtzCg
uq3/zXgIm8qiEZYD72PFM2g4G9wdsVT8WSmcaBmFNijOoHJcDfClmUQ7BlPVp8a8
eKFuPUsbM1hftdJjurO/GVqw25K3ZBJUGd9xYoslhdXvF2DbuKJnrt3PF0xahHGF
yYtsiNTDCckAZxAK9CSZLtaF7R3ipsrYMgfHCWHMQz+NjINKLEsnMPdYc8W1x51H
/a32UPu/oRwkbSNp+y/how5X05A/qL3XqokGFcbqRwnowBKj8B0sM2jeoDFvBYSU
EURLDQAr5uB6gVP7LXSkJgka1F9E8qF1xEB38GHub8/XEwSSPYCwQTgAsAPNQtAr
hNm/ejACUl9OWACNCCQLTxYlUhtJyR8PvS3LIfKrM1z3wQu2+5rbQLlGzoyvxDq4
Di0J+B0k6rDRpQGMPWCzgjtiiDwAdF9pE2bQFTZZ65vILnnWISGFbupy276g6WOA
omCsh4cXJHTa6ZkYwnw+jNqqEYalvE/CWRXYR2UVdtcxTvBGKzklKC08qVcegz0L
ax75CQPckZHvZMIsBps4ABMMUp9v6jWbAp7Ur0KMI9TKLfUwWgAQLwwYB+JO9U92
7DuPYgiUWxcTIQk/46YP4voFi3s3/rI3ix6mA4vXikT5u7kkvITLpua6OOYjLb4R
5ZJBro2XnxxNYTQRSaXvF/WJTgw1onDvUX3PaTLckSsYy1RVR3C1OEuk443f/540
gc5IU/IIJpJbm9DSCKlUVHrd8Px9BLg/zU4Aw45XA5qsrvfOBbC0II0JE6phlQyT
QStMPWXQ20zOaNIx+xB320f7jIR85rKEjWuXlzuArji5q1Gn3MKvN/36tsnS3DNH
Ra3mr2m5Cuce+/vvaXw08PNOrTFl+M3QlqPa+CkOaTL451Y/MN4nyphCWHeMLTaF
3P9foiUJxu1qKTN2O4BdQuY70kdwqyRyJeOkNQ42uRTA/35YHXBw2Znz+oquF+mY
jpBBtzjZlu2z43iunvIv4aJkP2x3lavNUGCLWetdpUiYHoPrwfoONQNzJ6oLWk4d
2vbsipi45rj/tom9wHHLzjq20W6zxkjmsPddwFX4JnEpxfrGIR1+P4xa4V3Su+uK
gtPzr7tiZXOZG2MKD0ei+diysSh4l8FDF44teekOW53mf4PAQs+sp28n3CtTvJ9I
ku9asqYiCJsJfW2vl2N1G2Chg2ThWSYbGXIABC5aSj6VYF9ry0eYFL1cZDpF26Xq
Q/xg2fjcHQh5Dpkw9JBOd6tA/Orlup4LSsIa0e9TEJbQ+u40lr416FV1jj55lIaH
`protect END_PROTECTED
