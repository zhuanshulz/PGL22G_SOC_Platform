`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LxCZOEGFfGGN2XPdd8dQlxeXMuYuN7JM4J63rxbsqgr0L5hIsOn7exziUgmEreXn
HaOEB3sMnBDe5OpCbXxuKZmfys1AqJL8mov6jWrwqV+NcXMD9CP5CabLQEilp0eZ
6KULm9ZM0IPmE4LZ+qWL62oJ+o/+KBo4nLCXf22SupIk6ksMnK3wFmSmpxOJKKfl
+FtGiPxZPFpvfdul1P/HfDoCLdSI0qy0woBProqwK4ViolFW3Upik25bvcAOAwGh
4EDz4MVi+q9OSG47EtLgUR723T359b1H+2CjqHXF6nF7LG79rwN34wrobfuS99rq
28srzYtnkUJbe587kauNNVdusjVtYLLfgjM6+feDZHEk7eMx2tnZyRRmUFkAkkCt
lLjYsulaB1Vo+d7QsSLq964Yv3J8HPM2mNGOOjmW5oDlCjKyd0xzV4HgcfzAsOwu
jceAR0xUwwZIu1w0NEozkjriGBIK9GVQwhMPEPWjry/ki/ZZh02pGI59x63rrgkE
8iMjGzMRVYzNZ80BfzyLj7n9WeFg5wYnaIRHD9tpu2Lk3rShrWm82InhgI32z0yG
IgVHz1qLGglmVvYqs96jK1Tp/Q57JdQCSJ/ilOqKKTGVLdWlhdmddgM7Z8ZeCQW7
Ej7mucIrF+DoF2aTDmWAIcTWD1SBar4le7w/WykBI3a8OcXfquueO5+hXOpfC5Pa
pcfVyJQLukTufVx/KTtVfW7MZnEySU9Op+YbZMiE+zdpEiWcZ7a39mbCltUaWO9g
yDCpHl5JeF22FXxcsarPoHWY3oEs2/Px29QNLiRzbz4=
`protect END_PROTECTED
