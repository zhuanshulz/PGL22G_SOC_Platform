`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fL3iyB5nmywilEnSrtx5LsnzYdW98ebnrISL0IyPrKamCPx9LjYMsCXNoahvxwnF
M/g0xR/L6EZrapKunPWcC40nLH5vTQlP4oLLEThC9QvbiHEFEQ30uy5wYsbHG+7L
Kq3SOxuZIJZuwT5zXD1oJr0Dyda4dTTazkkcGCd8tP0VmZ1amM0I+V3IF2NrhYHw
Q8Q1fxEkDgEImqcppXskmKY4QW3zTqarptXpNcVdZzJrHUsQHNlm3zdV+MpfDLqT
2B0ovRphmHhwkRZU4f/WGzecaf6q8xizLcz7DbcRm8CZInacb3gWckhOMoiKxIFz
z66Swi+hgJjxLffRsceErgj41gr5tRS4sk6gky7cMPA4DaNLeyczhrMieP28nV6O
XcfQKk3n6lnYNzcNnJSZy1qa5mO0t/gQjxFHTcqdJK7GOezOsU/tIy2Pq4bxP7NP
whCY5s9fBQX3E7Q45ukkJBUwX7CftJAc4RhfKaMuASMXCKj9xtgiPUo+RFbMj9I4
RtbGzDrwUcmzE209FEBr1Jsnhi3di6itY4LpiYPVdEDADvtvfvlErB1yLsDW8sos
Zqz0oYDo6mHfoMO4evwsi8EF8XfcEyO+WTInRwSZzaO8J9QfeJls6KhAl4yCE71F
QQONY/D2+VvidOBkQcM0TpeMKpdsANqQMZFhoQRI2di/s9QpchYagfseMVhcg7p3
3dInLAxH3KcWbJkcWW7nEDZyCet0p1fBLNAX00rPe3s1YyhY7jBqEyBX2zHkzCeY
PZfzBv4gt85AcFc4qLiRWpw4uDTLeHOFpsSgpfAKHQxHj9DQcmgfRVRx7e6vSyXk
7tpCUi28Tbnl9dZgPqDdnKE+6bKTn3m4x9G99xz7h7UmCjxN0pDMOhFXjPIuD6xg
6BuATtTHU/znuU7ALnc1Z5djR0QnbsmOmLfATpm9qDll70yYfqOahFJ/YbN+5JZa
TdDpFL9r/noDJEO1q0yYVVeurUNGqkLLVsVAMn77gaSS+2HVuRRrw/v3O6L9PMnb
KCLEkgjdHJyEQbNNovTxEIFEnsvcQiQQrhEwNX035Mdb45sB1mIc8cujY4s6URmB
HdpBFqz74F19QZskaKTgWlTrcEph5FsSHYQN2Qg2jgplrZ+R4dt1DTiys9MWeB2n
ekEhBiB6tn0tk7lBSQBNe76TcmWXZT8c0qfbuQTc89VBrT6F+YWj2eHTJtoTC7GC
JPk0PFvrgQaNRHgvleN2vakDVkUeEFEOhoEzymVoPztQDT13lzjgd8apHosueANq
ky2lTcKcer+JrS5ctGlH+5XAOHmy7tpVGVbPSMirhZdsTWsWszYPisvU4pe/klIp
NrtGw7lhtx7Y2HSOrnSeGLSWQlLSkblPDI4CrkT8/NjN+0R9Vogf3KNWO8KhwZlm
JKodeBxZMolB7RCCONTMAIGXyqzdtQ4in9ou3SywHp736G8P266RqN8YtoJXh5hD
4ktxM9OPYeeuBkO7b+bTXRqL5mL+eoNkocSTpf8Jt9KhGXu0qX3M0HR/j1zuwNoC
I/T21t1dkPVuC2tHdjJlTpfOcGrcidueUgSj2zmtvTqxcUHRSq1VmjkBSltYsIyg
cpQxLY5F0R2BOoKc90XHtvciamdBg4/qHPPPT6zfqNkkT1sbjMjapuGH928Zf4AI
JxU4/xdqC2QV1aWt8ws74jEuFafBUD2kCRAKb88tcEg3vclmTBwTYMXXfLXwP2rm
Pptks3W/kA7FiXwMHkmDEFamNS5D4zSoYwzgGT+IFJDh2s/i0LrfZEfz4Xj6/x4e
85MCmskCRnMdC4NNm0vJXohmKvbYdRrO5OnsAt7Z3a9SZwlUipJeWnrM0twpdjbJ
UrPOrJBnxDs/Z2CUYfzFzaU6IiXqXGDSBBj2fIMgQMqw0PWL8F7Za/elUeBe79fk
sfD6aV0n7ugb8j2qgUKjLInh/3pFHMDG0PYqMZ4+Ky94O5qrFEwZc7Tr9AO2jCjm
CxSmWp6Qz1GMZrj/cmjSiUdCoHPmZIIJ7xmf8lbtbxaaZB/7QB6SZ3sRau0H7PdC
KSZp5T70BkHbEtlfjViGs2mLCM/f0TiiuTiSmwrKY0yS7vuAWfBkhTjItCGriCTm
llCiF9tHiB96OuGzduZyptj9JPpHhTdb6Q/y9I5ftPTrnkqAZUbLyWtIiQP9v+3o
r5so+SAJmXc6grRh4ECMvmUsr1EgW7ztkr6KGM9gdVoQrKq5KNDBRKZJwidwpwag
O24LG0JfDeYKG/Qt2hEhcvIoiMRH2T+Xszib01qWqFQALRXGmqUNyRJp0W1A58GE
DbzbZIYqI3CHNXEFY5gTFj7OjiH7gh1C1ncaL7ctwkAIHEty2fxb6tiSjHKq+/mm
I/4fyEQQgBBVKUb7jdziJwATP5iw4ZQqsJ7uC8rHoW7U9yv1zYySB+Hvx+0jT10c
ldhSXrptBXhA1YN98bxiZC6NWiRp4+kqkmZNYlmMtzU4gyjiuHBrWp2V4Lp6UCfx
ycoNsCB56WiJUgzFU6vz9qNdxBKkGRAJZZ8fVKV9YZWytaUXpmtQx1Vm4kKorEFP
jdQY00HpbMEcB+eNaVA9PalWUktImTdc116sNbSOaV8GQF5JyBEdYVh3cBhLOpmq
8DxF/4pmntq9rPijeaWI/XICChKRMwKF1Wcgglo81GhG0nSlY3FQ6vRF7shTcG+y
WOmbqj3UNAM6/mpC3XyEsgTldqLoIUBVptb4sIGXBDS0BQVhr2TN2RvkbG7PXnHR
ue4al/mD/zsalyC1ea3dmCF3PuNvwgm48Hb/cKpNufxO8AAnXvmhvs3HyjmfmGty
vupOc+/AaS5hb8erHkmQO9QEo8gFaJuHHacsiXaXkv5QqeZP9dgfwM+eR0+McpSK
LprhZ3Mu+8WxNbAjzQMTEoa2Suc0RrZfHQPO03XnJZqIQ9QrOb4rC7xhZXTa9lBR
FC243B8YveV+LCKhvn1Y86UHkeFP/RvdZSLQJgJq0K9mqLTLZDWQ4GpcB9l2shP7
4GJ6V0nBNrgpwKnjFlxcZN4mipqD4P5FswMlwGXn8X4wKkD8iKdvKbZrm0Oy1Y5y
qBwUKTf6TPHhIK1GnvrRjSzhLYtBcWQ71bRgIEsQIoxwMFTZ6l5MsKONup0LTzPM
k48ODR6KuDXN1D+OP7MrHIGLxaGM/Auqft9j0ZfRCD0IUkCaQaOZ7FcsW6tA2f9E
o3zEy/m1rlQwiqGILX/KqV4hxTBMOBgQjZevxzoYwsUaVc8054AYNhEhFRjXaqvC
9xHl895Phd4UTLnVh4/Ff+CRWZ70VtAcxna8AhG6L3CWqb3Aq02xu/HSf64Km/uk
hsNMwFV1jvigGgr5JsomL04+KTcklLdjzqEMo4WbTiEV38eK6xfM1hyOxpIE8TEj
FgXQEODn/p+1hwcf2io/9xiyr2xf3JKKb5Z1HVGsi/ATshtW6AMVpz5BjFLXZz2R
P4/6i1aXxAu62YLMjqxtN9Jrn9vQBVLNb8uVyAsZoqJKzWKqY9C/kcTR1xbwv0AO
LQYCsc+7DJPMHth7BUNAWSDlRI52Dp2tN/umm5nC8Mdw7f5UmgeD2CiBJVOrOMUW
l6mTXtDIGV1Aifnvhaf9bWi4Fb3+e28BNzGQpf53egjP/MF3xhBCnFbRm4wZiTQO
49C4elTB1W9vFVMByGolKfZnGgrpakf0GANfHl5WoZO0F5W5eAkiErid3mTnM42D
AP0mBYblYXryyXQTFNfe8m5RPqv2ppkCWZ69rSnTXc+Nq7dvu+qjnEHLjwJIQ8aH
hN+av+Woapjsltelf3RhQUVC8zoOSUDDdILcMKXwlvDL3S5P6svvUAwtIFCHx5hn
J/ZW2yA9SL+xJOlMiknHYBmO2tnnglMUBPgtjM4Azd5Z1rJA0jxUSRYFMxB+lpP4
Uv4cybrJWabub/X7wXvIV3qEUv9bidI/e3yjJecLPstQ+j5UA3dq78hlaCk0/Tak
TYqpZyxzEAc6pEn81aB/lyhtRZrGNcnUuXl2kxROKjww5WMwYojGks7W0+UYutM6
frl590y93qguSiRyoPHxZq03evpvtTDd9/7OPm8qculcnlN+z6g4edDvJwsvzFiM
t4cW5qlLjizRsIXqW2wE0nAoj4pQwZcEvM9FJsH3IbTmM4FXGlzwhfc3knf7oZyZ
1rPoETGngVK7l+GCQWyNlQj0sjbeB2Aodg5fGgWIbNtA094wG7smhvqcGBTOeypH
W3ne/av3BUQ/Ly7rioJc/I4ec8JoYCnJBwSG7sTvT9vy00jOdijYpNstTxJKoanX
MPPxe01ks7qfpzaXq1LuoXE2y9xZvXVPCquxfbuxeBxcVR11f0R452OlFWw28GMW
amP8cq2Ve5nGBLGvOV0j/XRyt9iT+2H8RF/VBli/q75yE+5Yy/IOQJDdxiIWUFWL
Pl1Mqw3sTExBfbfl4gz2LhAgKSsT9I3xOG+WZHpd1RkpC5EIhSjSujQ2B+e1oBCN
sI9h9i8ecJYsm7XVreJfMVCqgwbzDWQZEnO3Fmuz/sfMpxn4CcKzTbLeLPPE1Eb3
WaKnVYf1QPG+gSBim0obNUGjSl5gN8GKN0tN9JUlVvvbNwjUVfkBW9gZ2viCE6Gz
0RB70RhzuyswJzB6HrdWUTvVK8wp8Fx8L/2rT2ZzJvmdXUgb/KDB9XQ4KS1qbJGk
TZvRKyoEeaLRn/Bl6MnY7OYvR/s7naeF7BhcmhjkKy+l6gDgIj/e6NanbIKISaPk
k+64vZ4E+ixgzFQdLm0C/2GStVE87Uj7Kk00Wf6GhU9CZrlgMS/R6xwNZYdmoyH/
K2TIXM3dT054jDx0RSL+lo6gzxRnD5H8OTglBSAyPnF1DWnZdhOdvJ2qKFCFx0dM
qDsglZcWo98k/rbrUABUvcRV+QtFPgR08jKtpL+mA1ELNPL41KY6J3K1Lg+Q0pUJ
uPp/AM1woSjiSA8h6NcgZ/fcekUWDBlsT/Dp8V+U6GwhLzgoZ6aSD3MakkcuHb60
mBDUR1lova+JwJKnD0iBvTcCUNSSQKBuUaWY7DgXYg1aSyuNe6O9EMz/hpdiYfGV
0ZfOHygeLMM+iUDyTNo7vg==
`protect END_PROTECTED
