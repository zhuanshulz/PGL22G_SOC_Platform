`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H67zgsQ4YkQyZWpMWs2To/YsLKYmGkngT0bKJowJFeR+He1uXsue6kv9tykBauEG
FiMkJnHqQEgXRPEAYO9Va7ttAgoHo7XDqeIK7dIjJiyjvRO5Gnu/AuXUSuMGKZNP
S/2+7c1us55VCWoScnuu2z1lPh75CK2Gvnv9szV7jg+mVfARzuji4XQlSIDav91Z
9CGKNUhPXnAtgzVHK8XpOwUEfL8cr5xKSJinPxqZhI7sbSckncJ05BvMLI6POz5v
eGWeNtxf9hq/2zPwC0hIF75vZk9hxQcZ28Yft7jBdbj0ll4T48zHVyHCKMW8w0+Z
hPtlgXItDkPX03DkZwvVxgd/UD6Zg1b9klAtfK1SbOwklnRMNVu7Ka08QYEGBKOw
oqgQa8lPdWKW6+nSQIEEiXIAuknMWKNDMRCpVguckIBeqoU34oFoWDhdQPab18NW
oRoOH61rHJs5akyOXqjRw33VUPF79OyayAURmu0KNQ1M7VRf+l5IH1mXYAlZcsKp
jjr7E1sRXB34thXm0egGb2TK26NEAtgfL6sf0BJY0ygBg7Vh3Otj1EyQpnwL+8AK
jO11w6NYRPsWaUPE0ebsBtsOvArtmZ+4GzFdNicRSb+N6oAApYhVp6hLk+aPgulw
6eHFv/mKjcIVI/Er8FsAEAyBkyEfwwI/nQQpAK1CZGv8NKXmWumMtu0xIaz9swaX
Jwyc9pkZnJM/4Be124JQ8XGFQb4NjIhnKf3vJpOVQ5tfScwLua1uHfDobijh+Iec
NgtqpsI4w5UKdLluFh6uFw0rpcoD796TBIAF7fENzQY=
`protect END_PROTECTED
