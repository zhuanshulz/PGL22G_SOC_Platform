`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1grPgEkJK1+nkfuiv4nTgEreQWZ49UZCXcCPN1B3dbojpqlDDjZToZvxucVh49J8
fIEGspDuMpGNsKhsQnDXkKSRYsPVb61AUIlbj0iTEOn+yhqhkgxQzDTZX9cuupY5
A9pGiXFZbJjq4Kk56R+go1FO6TCZNHe9v5N+tQMo9V4K70gsvTI1IBof9kcFBhTR
CvbtilgHpJlQUehdgLT6jcsZobZhV1Gw1d+St95IdzjXcFg6pl104EbwuJS14soT
P0+XYdtteUeoCPRJvPpG0n5sJ3Uh64t/x2fmBklnodm4rELHAn7Mo1V6D+oQO8ss
CV4kXfpO+cuWiQgcPfIEB5N3xoDNniwTWej2Z3lv8EkOrRjSkPVnvrXvPt5/hOTQ
bCzViUhpSLXFCCtUFjs8mMvPu7DE0fSW5zqYpuWgU6Vk8zLd2ZlqIegpjwq7dClx
TlVx6C00NxMy4IpzLCRHujrD482KYf12h61B1F8J64ueqMyDtPMkapLnv/ZLnY38
sodv6VmPHqsAPPqlQh/N31H7TyLa2SQl1jAesZGdtvIsWiJAiNUX+ShtUIGMUH9A
nzjEB4YQ7rsWwWoTqfJ9w2ZlXmx4o+Zz+s769V95F/6DUwUSNuxr4Y9xYBeLycdi
jCrxnEiMbAtdFAgXJRte/Kvx0iPzOHw/1L/AHTn+F2ovfF41uR1eYd7E/UczpQsz
AjN9ClNG5YWJapBGuxKlgDoL37MBBJjCSZc76I95W2Wd5u5nHySDOPVi7PxifDKO
IoS9oEyN3QTLj3I7EjuvzVfJhGl2vlypyaK64gjEgUGDHzeP0zCSCDT7KnjqYUV3
RZ42jG1n4mkF57AHiOWos70QSz1wDICxxiYssFI4Fu7oqsUh5ijuOf5unwd+W5FC
Poo+PFqB7b/NwWWvgm7PbF8NYviknJRsukvchSNjoueRCLl22VA8l4nl3/hByEPC
FjEMfPy/TqOdnaSa1PP5Opwruww6JmWp9AXVnSYb3O1aZhGjqAki6ROKvGNc2hMJ
iFhdOrLygbr36KYppoJuwM5u9N6fdsNyoiiJG4jrZlaK3zAzLo2MzbmgaRMU35cZ
BelVBJ4mmz/91Wj28HVPr8K0rAXCWrLbmkGKuVo2xhl9GGHTqfKK7Bnzqi9OMJ4X
ZJXMweCQ0yrwqx53D5EyJkgHqmbUVDxptiG2ymgOTF9RECOAKtdkovLE3CEyOtPR
/X6yoZoARUhW11X9HbE3IrarNs5J6iuAZAFe4wazilQZprmZ+PuS4ttDqngdQljm
LB4NET/jnyJ85XTSpJjJFkbFgycNwUsPAl2LGXoqZK1Vt49XQNkH3XfmtOjzwnNQ
XoIw2cYh0bonUoo25Vk7MEvfUJ1VZA3WEQapdZYs7Z4VAewNiHN9qGEu6uyIWtea
ZtkgV/B72XVUa0XfM3Tk0voanIwa+aYFHx3C26TV5Fwz2oADvu1RzYTZzt0g6CsK
U+TYWXiWwep7gK+njxScYkXcxX0Zt3/19M1Ut7MMfo7ZGsD3yRb0OEDh17Pny8+V
XKVRx08Y1/OXu0nJzwjgNZE/C7k4eh6Q78DGOvCcZmMNj0q96WRI6TDHLJAsg5a+
HB9+9ZozDv0ocQrQMNwZt55czyxl/d7N768xzpzkkVmAv9t39W/V3dVLaNg0LKQJ
Md5Ow3U6R3boh8Y08EkbcoL1uYhJJONxWH/hfZz5mjjThVStUrR4OdAA73KNkYyU
WNVEWwo2a6WnuogCVwY4diNhRUqqy4W/QVd62XNi0efcHJo5Ds8lfIlh1wBsovqz
c4qiR34FtCluineyFzyi9zn/BbYZjdVgOzK/RX6HGir5x8DPM2g9GK2NHj1yWaRd
wlYWuBCpCybpckquJ0h7egbCLcxi06ciZBYfYoyQk24Lmc8oJRm3vIBlvQYjEAIb
AIbdE2ruTR8kK5IhSAAFxhmPP6q7ixVqlU5hgXEGKyFAegtj6mT/QWGg3sHqwrFD
zwUOH1k0f3mzNwQ6HyUmI2Ckr+BoC1fKvpkOdyTE5PU6aBkUM2GHuEYqfGOxzuyA
0jyGYVZ7AiSNtubLz1qvB+vO94B/U2kXY16AYuqqgCTuNyp2JsBU5RDBHK1Orl60
p/TdAxz2/RXtuPCYS8hiP58VQkIB0uWnjgMbqqk9dwdIYF6uZjJasm/dIvT21cAw
oZ1Rendr5bNjlNjQA5f3TzszBu2/eXvYkApX33O6EpMFLBYMdp7V10xSyRI4EHmc
UUs1pau7M5y7rbMedJ7w1p+STWkzlFPGNLwNXL5LXz4t4C4Ah6MLDua5cHA22llp
VI5lttef850VbQZOVBrW3Gsu5ac1N/n38pcZkV8HD3VTW5AC5C1BqoEFBnkeNK+z
MKHGrUrvSMsxunwla8aQ8WM+oBL1Om6hz8DRxWiFCCKhhOdAL3m5LH5q3eVaMyho
EoJoOIlVV4qfQMWtbmiiVsgkOPCk0rtqb5/I7S3qWMP4QAYDNfjpN/cHFoc9yG/i
TH2iamUKHq8sfCqudo0HyUdeIzNDcyenDy1epM216rbbREpwIQh1FYDdat9orGoW
5vjJgV3nDSibqQN8+xUryQTUP54tB4zPnL3XJYhhwF8mCgP47LoMXsEVE1uQHhO2
fz3NPKodx90nNU8wbIU5pbPnXwbQFOedxdcmiU4xIVFxh/yJMVSD+ZeFgEQiwOBl
iao6/zkirqjhiqcShM0ZgRLZNafcFXnmJ15/IjKRg+bQNZkMgZfpprEMgJq4pUaC
NDBKJE9Qmv9pwpdpshPoLqaVbizlFreQQtVQ4QQdYM6nQvNYkoN0+8ehPQbSWHAY
Jd8OkuFgDAMZaAIAltavavXjSST10Nt+ahK5pM5xNtBUKGKKwa2dPVr7ynB8w2Hp
6FG9Y5oF/jELPergbPq49jtFtnV42IGyel1hvuGTn0HTTSk/6KDbfEIDkBNcL4sT
OcdCidUMzboP4NUSIxWfkSoEuLd+wBaGeTi67diHF0Qte6nc/euagq9DFzTXK2Nv
RqtvuWbc5vv91GDe6QpVoGucwCUYb0jT3kwtg7jfz6vmcSD2YwtSDHYl80w1ZHSr
dLToIFvMkRRufmzRZxTwl2PcbybNY8UKkiBLTqPxFb3+sexPRp1fe4L6YJdPkidB
JTUr7ncmo5nK+POUSeCamidN3W0RQESfP6Gscir/xhS4sr1YjzlqphudxPw37m9q
rtTqUa+0/0DdH1UVVfBpadYir4rBJzhYWP+F+4mukZLfqhPk2EW3sqUBje1pfggS
CiBugVzzPk5Dj9sj4JotmECK+2Rvnvh5JZNvkNFVWdIyHdSWizU2piH4Zo2kdEBr
yMlMpIUfeZGdRNeEzM5gm2ftv4gYlyfQg3wWSdOo4ReO9I7ZezF3/0xItOvR/WYL
E9unV+mVBR8TfieZuLlj+To1xIXm2QjeoFF41na6f0ZmA8G4buvOqo0p/rbrAkSc
asYd1yUyuZPvV7Fxxb/l5Y5cSQ/MFu8CWe6Sn9qMVl8cD6Kq+mpCtIkuuSNkQs4h
Mb96yo/u0RAI/UABZ6d15Wmiz/g+uG4tgOOZCuSw3AjGm0vU2yNjhg25PzuiUJPZ
xl3QRRiz5mli7LoEqLgq/mFSnILwocho8mAMwK7bnu7Gw2QwGaNAi4DBQ0f6Hn3P
ZxtD/OrP1ZS9PFMmSf/gZdiyTNmnvYIAUYcmbYvUTWGQF6PKYLhHyVm0h+2OXIM1
ylJwvvZKpII92Jo0sDSG/FGfvmsz9UIt2QgbS4gawZrwpUbgEoQ6UybgxAgLMxin
wJsDnhCQQZ522kTbBzeaio5LTFBa8AShptiBAB7QLrcwE4YFIXsX0XhuhzOcr9A3
/6823PxKAAhAJ37qt35NDzRsyUdMTHE9+5su/nRd1cpMQG9MPHOcq13j/oYHl0xW
nEPNmQAo1mjiChn0iptsoxDx5btWhqTk1wwoaYUrnqWUYOrKkaxf+7hqGQKdvH0p
JkDE6rYS4f56d1tO4H4SR96fcmtFoEj2qpl6SqtjxW6GrDEJza6AcD6qPrdevFi6
EeqKseMbS++fFVQfJ/WDqIu5Ji+gOnHRymTOz6R8CsTbGGRWAEeLFxdcELFcnVT+
65tX9ZVROtNKY3O5bAB0Z5c+8BAL2Vdg4y6JpNlr6BjoDmu3rh8tHYPx45ECuDS4
0k57FrtxXsopMEbPHZ6qAsjXRwzRcThENVGBraW3rEDun/xkhk4JjHWTJsTuF836
hZBsSPSca4gqhKxyTV8LRtolxgF1ZeZCiy4hpnoma3n0m+KRpiYRLTmKeKBlYUUC
fBMnG22EDIbP74tQGpYNK+412J6BYCz/MGnjHxd/axNUAPVxPP48Sf3PVyr8TrMP
G8Y/8+ZMx70nXK2q+hvBSpzRTQmGnjFnEHYSGT7K/RTsuV2dky5rw3Z93o7/zGXG
dm4mUmblMzNFrBKi9S9W2TSnWZwaHf9Ezqu5uDHfbahPsN5XvTgLtH3t40mTpsAF
FrPusUYOw4D1lwlNItSX7b99C4xnq75r8AXi2dNpjStysrpVegRlCYehI6Y2Y/UN
Cinr3sSCpzWxROiusrWF2uj5AwVRi7bbmcotUI/6mSvm1YiQ+VgHz34NwyYwG2fU
k+FmSkWfoi4/64UCWM/9IIdWZFeWm7UX7wYBiJfyYvpCue+7+jtqHCfA6GIsQW+k
VqjFVrNXrQ7GcuVq8KV0A3ITdQ5M8VHv9ctd7hgwi8MO0VvBxOqnIG4rc1+kLz6Q
vkV7gpr1psyenUiZ9OwMH3kLs8oDHl/sw5ZAP7GuPBJMQktWW/Paa91CneZCfBox
CxZ4Q9i3or3YZZf3qHgMYP08S8Gf0fJGhtMNbuUMezog74PVX75O4BWhnHq9uH8E
2oZ8EUnfy+HIRZw/1FL1KeMj2kuVsq3gwrG8gECKkjuek6HP5kMSbsGfalmPtdE9
PNUMNwhAKlWZeaCGQmivE4O9/u/zPkdSfeFsUJ5DckJwxHpEQDD5usVxq6+xyrSy
jngboILmEHsWHhiyvr3ke7lTmkAe54jjU9h7J1vTGoNPtqdi0p+RErKFXWeRknaR
v32/pRN8FxBCBrVNb3bVpMOBsn7IrpUF/Bx+MxrSKhuSETIv/D4jeaCzQJ7f+68h
vHn77szObys452SDSQo2eQe1eIOHApj464gknwdZuGPCthGJiz3bBZU7vLuZNmTM
SpfWHumhw/3LXYkRPKSLoaVpAgY1iMKbLzICupdDNmdlapxLM2b0Wt7GLwfd44pF
Aeb8ICb6y9DBIsGVl/nurfciIkOgjJCZzL1eD2qul/+rGrRx6YGIjTKVlDW2cmWu
oWgsSZWPCniEg1l+DnAe5egf02Ah+1qo4A1cnd6i8GPJ3IHemEKbTERmbfxi3UT4
hXzivCmDYoXCR3g01e+FlynzD5Xj4gcZh6dn0qlIY6ksHbzjgE6EuTxjgyw2kFLF
BP5WKV+TJ3kp47LXOlzcJ+JwdGx5z72GKoocPcIOMtdIPZDTquQWh67K/rhfaojP
UpYhN0zPZ/VMJK51XLsAeBCzLiZa9eSTtwwmdhl1r3SO7sVpXCndL0tiokmpdXy2
i2ZOKQhaAzEWrCwD1hkir7rZYx3W2HNP5NlqhU/a5GK/T3V+8je/tdDq4tOLwZ6d
uEPvLWqt2amXg1jVu7s2l/O4TMUS8wV5GFygBLnx2p7kcYen6OVbLfHjLuZyJSqD
kMPCiMHYGKgNRbKuXbnUUbOXTlCiZv2GGYpBXso0qkkq4iKNLf2342eigeZ6J8dO
XGsPVTGtxjmwaUym9ZvhSa8Czgaq3bFSsqWpb1oBqsnzByrzarKCqUmwytxeJSHV
WMJ5IHexANb3W+6T6IWA38KnosPE6VcXkKfgrTnZ/Bz093LwC8+1d2ttHQYURYJS
C0K7+JTqkG5nzD9Gfu0rAVT9m2as5Si1KP8FIEbYGpxcQGEpeqIz3Hmva/TBqpr+
cqGKptgw+R6DCfHWU9kTM0M3l/kVv8ydm8zxTRNPo+t12P3q1OjIUh5FQJVXMxbH
rawLVIadjp86t9xTisheCeyd6eDWOkM7SlsPZanLLHNg6GB3WMFmUo6QPUxcKLuo
FJdGQIwJwGJjELhWLswDWCoVleEezhOFRsiZwoJJ8pM=
`protect END_PROTECTED
