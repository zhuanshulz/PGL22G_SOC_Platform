`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7FdiKoGEHscviLrWzthnJxFhDxtto4nEetR30YNERmukapJTd7K2SATcU1/R7cY
kC6Y48L+zKYFYrD1p5W4iPbUSzCYJfpUDUfMdQChaS0HMFIsx6WTupkfRNvaOspL
LXfaUKPfjFIrqj/3q4cH7TxhvlJDRQOlhWKmNHYbj4BpJY4CxohQjp4rlwUk0rtd
3i5U7I83krq7BIqugKHwRksCbznWPXcisIf2vb/3zZ+YGh9pL5ztZO7xzZtdpTx0
e+2eH7KIaZq2qM2GWiFaIvmAw9h4yK8xUVyi7JcFkkkxxKQ8karavGNSLyhBI4Ws
gNF3teMS6mdYLAQjl+ALreUtou3uMCXPUukbKzuAOaAyVPsoPYdNPAcT485NPhAm
QUK23Th5EKQFas+fDHfW2xPibmpBHZaVTPahb33tHQlp/bdMpiiNmcklF7VcXW92
EiUknBL/rwVTwpro5HPMJWZzKKkXGmmR5BF3epLkAT8jQj8eVTfXdRUUU9AUAauJ
zv40yuMUXtkugK76znzOKbBMHQr6+fRPNfgGME+a4dHEFNgU8HK7+Bslo6HoDrth
M0V+CD0hbu2U71nSlwvP65fbXoqOSAOFJHFuHjXXfWFyo3SfAiPjZZ9WymPr/uWo
Vu/ltyJaPsBW1Zek9Gly8szcUPFJ2pR2uM+12Wxu4lAbXj6o9oqTwJx8I2IvENm6
KJK5M6XuKYGQ08Fth2SU1gRNFMe0LO8RU34GirVrBXa+JbeayDklFpBeTlv4gfM8
/KQxJRX1vjsE2xZXF09FBEF8AuSiYJBfo/Ah8gBOUHP0mSKUwyZyMHaua7sLNN8L
l2vqzDyDX+ndIps1B0mqsRiBK+ucQAf2k+Y44EmEGv/1YoTgHQnBgY7ZJxktOkXZ
H/NoUiG1PhPD2nw+bqd5XZEwGJ0Hrubkw8lw+q9PwOYgqW0i3I9yjk2gAqySgE2R
4IEOHJg4N6TPk/meu+zJNp+tN/X+0DvHgdiIY5xZixe/N8ZYmOXEtPsMmEwMOApN
rCLyqaUevwCP0YInJy9cLI2J+kZhJD707TRw3khYpXFfQVhgER6LSGGtPzUELhuq
gsZVzer+j46nlWZwOs5xkV9qfhl526EOpVheHam84twjKgW1Jt6X3Z+jrHUf6br3
d+SKVkl9KdctcbgZYKjdk+C/MRFMJsK0zhCkXaBvi3vo4gciVLU4rpgV4Uvlezac
+FfgaPgM8Rq2jZqN8PwLpsc+ogB7Xa2gR6jUUFn4heJ5m1tviJ1pmz2+6bq3VtsW
pMGkpDtwva6DGy2phPNLMV92OFqZo0BLUEp7RoMMK7J3bffzFOiPdEnS4RicqfDa
aZWVLHNm/wnwrby6UlwmR9MepUZP+VK0IfJgjATpCnjSj8C7KQfezUV3PHl4RiKJ
gFg62/TqkLVfh82FOYvL7+gmLxWncILI56oPq9664Du5K6NVH/aZbLksFeVCnbWR
94ap4H/QhZaNrTjDX7Q4SagNYf49VMoRAIuDwOxDaIYTEwsxzhYuc7nfbxzK6gIG
69vXTHzqZI4ZLfwMI0d6jYw3SHkvXtR4Q8QjtZ6s+JIjF2sKI2kohH4a0Yge8gRs
P6uXFPABXNaer1f1JKpe3pKwrFj7QBOHxtv+WNFfPtMDDhouC0w4WvdMoRUy5QAg
fnYLww/94Ca10gAi3PxmepJhpVUwFqk2SAaZdWFt1WgaeAkZ5hfljqwvbsTZJWCR
CgS79dlbvMkga9mKT40Q3o8Vo5U0cxrBkSMnuTkKlDn4ECEABV/U5Mb+nztJThzR
Ow7z4OcSfVk7KjF6brjm0Glkd7rwQzQ+8jna0m5THuahygmeCByoqJzadB61bG4r
PIH7zxJbCw3yQvofUQX2ngSFAfzNBqUZnvbKCq1N3d4sq8PLzUHKVaNHeQ53tjB+
GhJYGGAgpFpV2cK7QSTHG8iYUYvD3b71xVJ1VQZE/z3ZHBW/LhrqEPbFTYCtFZBi
LpA+iViUpjqy24xMj4yZdnYlCYNBF336oHOhNzNgN9vdjzHjO+RZNqvNUuZ0rly0
0jKzn81oDDUkLYo597qDX6r0hmB4+91nn3V1GWTj7WKsuHrM6/47pIjBMk5egIAF
H5C6Oh+p13XOWWs19RQ90+yigHqv0/CUWHVtutUsyDvTSJOmO4af9/lByzg0nePR
C9LXDwDyPqKgG8OKvcrbgQ==
`protect END_PROTECTED
