`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SrRR77L1+cSn3cacqMasNcOLkU9hWd/iKSaH9Fpc8dRG21GCtWbOghmXvNJ8zOS4
3W6Hpx84hY9JrM4YKCX1RJCLa/Dlvrz3dNs3RXC/UcHmkA4T9kNfNkQMR+7jIc6M
a5qeWZMNc/WBOSZYVsEQoCIVJinauZH9yKx8FO2zDdqcuCyCqpODX34AD2ESs1+d
0mPjrFROVTgDqzf5Gb+1Z/MK1q+G6eAhusznjj1TTcCujX+QLpWSOrmTx5HsdE5N
+sW0WWCf7BrkvhzHHVPxUikT0BzPJIao8Epr9ob8e39eyeg+cxFXi60rbCU2JrcD
GySwlsGTJ2LtRMuPlXuCVSaklmMB6dsCJ2BLLzS3nDKTcY6v+GxPMiJvI6zP42Y0
PbLEbxA8wRpEDFIguh5G14HeZ5gdP99FbuJztdqw3GHHy0hciziWgeiOIhzjb+K7
qmEmQfHqStYjcMSsQG98NhinGYhmCZJpPh5slj0zDdM5fpUNjbO7NT9x2O2KhV/6
IMCJqL8wFFm+DBaWABwsxd16UTD21gvqKqiaHFVKuTMnVBctsOSui8eYqWaDNHgw
hGNW6/gI6026c2D5eMoI9AsgNKYZVvlEchKKFFdtmLi7l+iWSZAU2fj3J6/cR03U
5vH+bZl8ywKmkcMvS/aIO0PoYc3DqsUbChP4KK+b2pRmO9XMPh85iqPv/OvsN0zn
yd8/Bed00w8Qnuc6mBey+PVeI4XAaKclmfy8vjaNpSkK1rKMov/kvp89ejWsNlGs
Wva2VWOAS9LvCxg3z2k0qdzAh1NRAoeez8jrDT+GHid2Ivdueo5JjqYpn3XtOEwv
l05SUiUm9KowRkmxncI5o5nbpw67hIX2X72Hhtz4hpQnktqFxKTwLuR3Hk7dJDfk
w8pLDDm47mAgLzNJ1v13jI+vty3gslZBeMvpYIIl1VYJdfJ+lKRaXwyF8Fo6i/R1
XKX8bUbdK/zqfhHhzmETQJMHDlS9pOoy+g97k0skhAWZUB+pU4rX7csE7ksTCMb9
sVRUIgZl5+yH9Au53mOlKEXibHq+36A4exJnMWmmy2lxU+mJl8dRTwlxfaC6y6F0
dg1bLwj+8QINF+7QgJPfbFltVLibK0jFYZuaZ2RyIPoXqXfKzmB6rsNphNrxw6NT
Rkpof3HRV8hq1405DH1q6qpBrBTvk/pAr/4WZM/b6dSM8sCJf45edoWIodPK2CmW
atSz7L2HgcEXgzlHPpxD2ae8LKtOAokBwbkNjMrY5G+qb/87CTeaTg7EYo65SqKa
U1dqMUxNo/rNDLXz9QIdccpwAf0AzkVSrKAIVPJ5T4c7PvMuyC4z6VJIi5QvLrmF
FhFCW5J3m3fa+R1z/G3lqvuryO9lNOrhrVJTh2kH1e65+XF0GKK4NPh4DVnGjQys
4h84YgP8aJuaLY0ie+fhF7YNHopNHbpFYjaubG+0NIJW8V1ucZRjImBS5NRWSC0t
QCF+h3TugvMtWfbkNogNYq4GHQk/sewNsqF8/QTHrju2p6U0TsKn9Y85pu9LjHO6
q2l4s5cAerUEzbw6QLzaVAXH4gzYYKhD1rIn94HtnZiCG+i5fh+2Xh2Rg6r1k1Tx
BA7vH0BdJCL+TIq6Iohsws+QH1TZ4YOUbRjLvkcHQTxmo+z1VOOtHqgNlGYMeCr4
r+valdoid4p+A+wBiDbHPHRXyOaW9wTLySJHJG4mphXmA+yLJfk4DhTNHDfexe+f
gY6OrB2J69zz805zeT7wrdFnz7WtPA+U4jigfsBWBknwhiGBkcQspjey+PMGqRkY
DHYTs4hU20bxi78xOPJxjVvE/KEx0Nra0AD/vRtiCzYdpCC9ZQp/SSjEFzYGz3kk
3bE4hOA0CBmuWiCibv775NppRQIWtULvVhdeRV4ghGP9Hv8hQvAhGGSphDqzN+Uy
o4bNCPpTSjJWIUHq3NF0cRHLcuTtvwIf7KGD2Bp0pa+GruqJnNIo969z0bLv02JQ
89jUbFdl8SAZ3KsTB4cpr9/SmZKMBE60qGUTzvaBdvrpBtOKiHswJ9EEARnTNGLs
z0gzI00BRZuOmfGdwvad0Sf+efXkcYrWe4ZqdcZT8ANIbbj44oXfd7it9TjozV0W
fAkT+M6PtQ5oM98lNNs/tu0hCNyHKzAVCg2B4BP7740H2t7yfrCrbJLYBfpyg+Sl
uy4JtIS9mtch26DaR1mr5AKTIXHeRznHpxFnZ7HhYRiluQqwkkSnRBIUXfz/EYjj
2zEL+lLKUscZvAG7maYtTrrYrEWzN0/GUV1SYuK4fonRR2hOzsZ9CAgDmO2E7hI/
qjp2SQlIIB/7kkdIW159xpjCXVdqwLsCA5F5OXMIxp+OnS22Fjr6bl0SL4ti97VS
2f1brWltMTvKjSrGCUDtEJoEt1OpjDqXbjacDptOM50WlvHZZDomLAR305HWs8d/
0TweVVrVMQc1Ac63rAyrXhIbhQ/I6rsZfIk0IHU7ibcf4jcxWJvG+vdnkHg5aXQ6
vyec+VeuV2kkLtcuuRy0GgDN4pxq6HV3IK8F6hnjf5RWGiG1lAPRwNiyWAMNAGFf
Zu2yp5Uihfq+AE5I9eqH3vJMmT4T1vmpGkeq7K+4PHznezeALISEaeWYz8Xc+Xv2
IZ0LKW+qRbIKWaXYLCufxjSsb3gBkeFys74TK7RVzgjkEH8U3/AW8sJz7a3d/vdq
kmSSbNlPOdXX4UloU0s9x9gC15a3ETxVM4B7cUfQiB80uuLl/DTb30znn95Mi70Y
5b0Wh5T3TIlpY/yj5ftUsD5aFsvnvLF2nRvHY/VmYj0Za2EuA/szU3L99u57dv+X
cj4b1HcYACryNnpPdswusLCgPnqpbXGjSTZ73At8J89T5WupxUeOMCgYkgGZSGYv
VmZtusTsP4s66R3uwcPJ9dDstmuxdEub+W1DiUlmzTpRxeebapZkj1GOJFDRsmFz
lZFrmeGzHBRc/7Z0KBaeXRh38IDGmexwKCskIFDsSZG2hHhaJDz5P81dlnQwIzwq
4JuEz5phgvAIN/fKeHA6gXOz2Eo6k4Q11ERWlflFUKrcSHAfCeF2P5IXsqtYhgHC
+pIOswFyQ0Wl7Igd42CRHGSGeDDPXOADsYHL4y8s38OQZ+tw5RD2RU8GPhtGljVb
I1+lURcn0WLvVQEE7XJ5I4yzRn1J2m6150VFFAT/KJhCCn260ygo44CL30X4GA57
oHSUvnxMBwVSlc+u0aO+j06kvM8soHJPA7BgJaEJc1YzqqIR5OPE31AS65DNnMzf
IiltcqQnxt2SujIiSEKxPW5Dufr9E8YlHq/krBw5h8qbzSWVfaYszcV6VTfTxoFK
3tp4dOfXTqm4bphIk40WKHaflHmxNTQeKTBHd8w6kwiBcpx1kuoI+D15QqtpEs4G
AFlUWOQhNaOOrwab0Q+2nQbNLA+AZZYv94gMAxEwUndiY7/yEUY3Yu06yd2m0VOY
rIdKJpTrJ7ETo8vnX79jbEELaY1ByRsG5APJgG3S1Q9aRDhC/gGSCAp4SRKChEgr
hnTnMmTPuh+qeaXjJf3ti6d6GAkhg3XwpkGsPFRO7xagKNQJHipGXbYQ2Ecxquix
Sw7O9j2jiHWPQRRmUSgQ16nmcBYZXwPnYRtSsuGxre1eqomQfUZrkgsUHpir7r9F
0FmuHO+oNrRPrh/szRwbcaG3F+k2jTyY88ZwQWns3w8QiRZe5CruBcV6IYGY66kk
qnLEKktnWdL2hR0Jm7AKDqsxLGaxqzAnmLUfPSm52I2/RB+SLuPQrInEaGlqiftM
ERx8C4Ytt38G7SMaSJvn49ITAR6i2wtwpcDOUB5rdRr9yhoZ/MFyA1lIxhgfGn62
wk4GzlXytFyP3ub03hTQ9dc3lE4FjmlUZ+BxNo0I/dXU8AqdOV3ue3jIorO2RCJt
JgRTJNizoHgqdkqe4cJaBdMAGW0v1rRGyGiY+8ExWHhcm9+0H1/wo9WHbXVPxhSz
AZKKgovlRb8jA+wUSKRC/Vwjp9oBqbRSvVfeeHjGxd6sClD5UbayKo9/CCQhr/E3
1pJyFLjLNu4nCQzx4C3g0lp+Zz+v/quPWyLH19ZeGW0IpL+dBfBW2gsXwT+DhwBN
7SaYf59C0JBLH7CgoPJpr+iMGQe6uX0wAZSyA5ml/Cz4+jueorDlPdQYrhh7t+9r
xDELhzvLa9wHQPZi4FtZ67MMnO2l2jth3hx1P+PbMpKD5wJeeuosRNLlAjNNvZVb
TyNMkUVUhjR1z+SI3rs2VyV2dP4LIinTzkg0CDpp2nu8FNxc4bmC5XvYIhZRK9z1
MjIjL0tKgvPKtxaZYWq6qnH8b12yMAAHDRPpxkkuJt102gzlm0dR0mKSorl1wdF5
Xkav5QiQpLzfgvAkrXGzobhu/qFc/tJ1VcemvEKtMBy/FtqNGvY3k6OqATSZYkCG
ePbk+n8tzH3aTfgf2XEaJ16xn1W+cPMrcFUYo42SWOBQ2k+8P7ydJR2xBhCB/ISQ
1YGGg/O2GYFoh4FEuhljsBp8p5AYiAzRpOQhyX7D2Z42x4ITqzb/es1Vi2wj5tpH
mJF6zQsVWCaWxDExLOwhdpszW7RN0HoJeHduDwobcuNVV2YPpZibflT04fn1C//4
PcbntlZqd51HtafMoq5hwfvmcDysGrYLd6kFotlDF5Un0GHxqgE0qLuKwy4Sn+is
DoE7NQJliLYQCHSpBKNlQBp3oHTrvtqiZ2Y8qsTmaFxxp7LwdQZpsDmCxz3DiLUn
XZ2QCADxglY+9feIlLdsly7YSawSFNMJLCujfKC6nTLlEMCtY/H2ol2SokOoyCTH
Zr2r7ZoTjHdYlbwNnuFSYFv1wqi+UCIBYjvJ3bZHf6q2SZceCddlwM2mg402SGzF
XDXKHSH8XDRhbsdRVobEN2MGw0wv1RRx6IVUSRpLFJ1+TTGL56u0/0sCf25hfP+B
Y+ZUjs8AJpiQUbeXFMOvmlCp6Nk4PKwv2LazCyssePWzm5uO6ahBnMRALg7a4STY
3VOdbzf3C+LSb4iomtrNgJhG0r1hMnkj8wlCEv4x1XF6IRkNnaclMb7InzWZApE2
C8yDY5N3XyJcbfjrt/9Rf/RXCGkTmQPgEVYpm/bKd+78coedIMmMbfBx7V2Bt+J/
gwL6/tRGUAIS8vL9O2PCal6C9Sns6UFtVcQv8/C0YRbQx3+3XoIn01zGb3+0Fx9x
RF+l+PlvBiAYG29SXutsAGCrOpsFyFEeHWcU/2EE4y2XqxFa5bqIN4u6kvjKLLOk
gP5aNZPPj9qTSvDVBCS+xVYpSr9zvKQlXt+3UHrM8wprLVNHicPXbZLTb5AP+VOo
hef6ASqQd7/WFi8COpChAFlKWAANqHcr9IljXV9PO6mZw3Fc1XBwXrmL130wretv
U5Gy16YxL04w+3fNkdl+QTpstMGSk5bspcBknLGK9hF1y0sTQ2nwtkHDDq8iHt99
Nr6mkW0pl8NR25gIduR5RZWF6Aa70Fpm39prwoM17n660s7yjeBYjgnHbud4o7+T
G0bh1uRvM3m41CEN2C9H58CUV1sZ9cpbsvDac6ztxN3nBt5ou7zn6q/ER58souP0
HhUz04CWW56zFHNy3S3I/FSpQ7MpfIVR0cfsAjOBPiba5wm4kYIFoKpK2a0D6xSy
iKBmgDsF5rNzgSfLSSsVDm2pGejLHmbwpwenXjlI/LKRD8wDHe/sZE+lvx+sgCGs
Mhkqddjy8I4UwQmH7GWq4qsXhqnV1CWjzz72sxvo8iuiIR0pKtQ9/JSdMM9Of7fI
wNRJGJOvjT8AaE27mUcoxcP4G8G5qz47cRSVPGLi5jk0iwr0l0OXy0tyUsvJyhjP
6N6JUCqxBPZ6iUwbaNqcQFgg24F64+ajpaNXjk+SKVQ49aMhYefN7Jqug/2K6uEA
Fq9yzgTWtpUcf7Dcp5PFbP2YiN8Vx7bpDpnNdqmA7AoGELHXGlB+CP5/2P1b8vKA
WXFrvbPQLCRlAaVbynCGIRUpSFClRNfcWwQChz9st4MhdKLGZIZKxxpD2GKv5Dyb
yw5pMOBGIythn2ySCKQkQscUNrIY6qDrlMpKlHJbHZ6yDrOJp1AZcG8VJVL3x2yu
wBA88CjqcPe3na0QREMLW1fPBQ9QhgpqiA7QFGiFiG1PL/NhCnwFZg3LHh1xds5a
hzx4uudLosjhFKfDUU4Is2NvSuD9T2KqKJKDNg1oIqOXybNCMWRyF7qVpZK302Pf
PG4zy8hZoRosTRh6nQYfJVzsZX9SyEE2qTbMRUQFboR4iPI5661vYiuSHK9LI7KR
2A7cXBH00ipmJqEjAKerRo4Q64RDHUbRmco5geV++Gz0Pi+ycEsK5eqqEwxIviXl
4h0apaPs4C6LibnhGkq8ZmXp+vAg6Qmue5DJTs/yf4RuAcXUT5pV24TUUmHRn/Et
QYM4z9xF9xXusuOTI6E9xZTaMfjVV1u20FR985NQIahriDggx/K8YyWLiaCm0djk
mf5HFJ+a7M2nFXYfGCvmmGr6ThhxU64cRAFySH48BKidpm3vNzH1MCD7pVN2rG75
eaUTjooDpIJZXEx+e8uRbrIOH91jk/IFAlr4nAxaaeliIBKVqWCFKEMwT4c7B1jJ
e4o7tSHuHuN0fTWX8Sooy4HBQtDAI4jFuZPrxkpwSn+EczVS1HhA9Q2k0E59RRWt
tJ3VdRV3K5C9YBs+ndjFDM4/Moi1M4thu10hyEEvzKd4QGXguRFYjXVHCl71RtLZ
1DHd3LurGeQngVhW2VkngKc/nTJY1y/j3CirFoEj7wjsAf9ovx5qpjc4LmevNRF7
2ZdBm9lW+NZJwVDn8x1b2SlgaNDgdkwIDdihlAqe8CWLjyJd43CP0fJeHxndfvqk
k5UqFfyl6rhl3EqBlsGWba7HqVmIk4i82JyD3voWCSe1Cs2+vzf7F9z6V5Dn/aZh
wgGOpZR1IYN2tgCxYJRj+Di3nUQYSqbUymHNSdAqP8CplyaxMr+x7XjRTM81S8vB
VemwtWmAN8W0rklqRNh1wA7IM/cdQC6f4CTWj3e0iPxKFVouCWekj2xoIgZCcfJM
tef7naBxKuv4M/+XrV77K3vyYDwxetaZLoRnQIMNwQFEDhyI1m/vBnZEsd8B/60N
Pr/tnPgOe7oHUMmdnY3ScUHiG957DbgEEsoB5e/+1vPsMB0mL1nEiiVOHLswAdak
slgH0bvPangKKG0g9+mY2HTVWCS5HYKKZVUS885gZ+IY9FzaohCUnlZwXl2S1t47
GJEYWmcYiXNZioqNkG0chKtC7o+HcA4lzWTbFIWEzG14H6jN2jkm8zLckASTbftI
Op2tQX3icQT0HivgpZi44ZISkjAr4dzZoyoyujM5J295qgQEGLKj8vyIrHnPaJds
WDL1CWN7Gf8sHBKIkDq5R2i+Dd6MAiSDZ3SlrjXUWqNoSCf9Oe+OD+i4W3FBW0vd
qgtnEdF2CMzRAAkUs/2cKoj68m6iZRVJKyEzJO6flw0Gt+PT87NRIXH/pDqsRE2j
iA+3TxmDisyDgHuhWXfTDpUF/Flzocpri+KS0SGiW27hvTmY4ix3nNnH9sg83kmM
BdUQ5SSl1DJxguOOsR7hrDXy1BYdyT4zYQn0ekAveoBaadivqdG0Fmc0ShIlmzDF
6HZ5xqLbFbYPmuPDFTeNLFCeSG0S3qjv9LBK83rPkK+Oi/IuHrO4AivrlhA0xOl+
r3xiNE34XcpxFEHYkpiP++NlrlxDwVaKBTTFJjBj3XqK1aHPW6oiGDCeL2Xh/AVi
73kvoyDh3J497zcVn4DpAo3UcLUqgUMDxc325jn8pQ1gtlYZ3fEtPeFJvrsNW5id
WZVz0CtbdN8Ko8unn3u93TVmUI9sCg5wIv1IyW4nHifSFYcm77QVchesjkrMUpMf
+RAbAf+gjzcLFg2oxcFSuPIVMm3EDEt4ffzZPcNq/Rhm50cX2hkemphSFH3zD0NF
wmfw2RUAvgIls4NXxqzbEcZjPWELlJmaNMXOm2T56VaD+3PnmbFB0YdHxoPO2scf
I7jOmZypa7UBAtnHeyo348plMnlsIp00uP+zKYu+bKY2xKx1BiIffH/ytVeRryn5
QR5sxt5kK513+QijelPUPqXxPEuTmRwLmGCVOaHf/vKJtZ6f0Mnfz8lS0HLG+xYj
IGj0j/h7B3DQCXbUjgRDSwPtFNo0bLICc46j3XkZnaB1Y85wgSha3LBbobsTtVC6
KftTqt94HZ79XpZoWufV199U7Rcx6cW+LXi/n2044tAjVcEoFewNOyXkKgu47Yc0
HkM6g1FfjyOuCS5ThQrmYFX8aeFordktsqlryNwi/0hM6PAmAs7giSXNlgb9l5r4
Sf+XwsM/PX+a9Cdd3H0PM6Z1PqVn6FUj2D6SKBFoDQc+QZV1UEQSd+rk7qAnE7x6
sAe86N0N6iw2ST/r13+xMsRMoOocqQwFw720fSw9hSBunBIoL5VDF5w6op9Tjg+d
Z3UKC80DJJc3KPsmk1a/G2oLl+eHxgF8Gc1kIp//F+ZYEFDIJcaSAEXV2wbZTDjF
Dr0cMMWOUUFRDiJh6R2m4TwMRNSUWyzr4ScrX1MfyzsIDL3l063+HpGOTk06C//U
+tjNGCeMHlAPtdXi9gFZHUTsG9Vm4Dmcj9iyVpQ8CpXUr/v1O5fZZXuELSAMdHNA
Jude2dZJpUuz0eS7J7zFSEm3KMeU+szO2Nz7hRvtB42Damxu+eDF1Km/ZJVJGjoc
hwc6XI3Fy2zhaaPXvDE+tZm64L6sUZX0o80xPM2/+32lz8HyJ7ZVARjnIhVuzJ7q
UHAtfi6dR3AYBE9LRe4TGkPTKxbgAiIrGbM1tWGbowrZnHr7HND16nfsEqLhh2F0
0mlcHdOGk3v47D5VMHp7nHv53tfiqo9eHnNVFAppPD+udNwxu9cR+pMfbgyfjRCM
3rfu9WFpijrbd9NS/zRV4reT1tn9Co3/NKIm95LVe4d2SIS5DL7LM64NTnrOYcXX
pksM4GwXfLfIAn/Sz4cHqwK1Pm2KZmk6xmIkUVYimyjiG3Uwrmc7xymsrmZjtkYn
M37jhtqPvGo/hlkmrzyfbBPIw37QBZAKQWLdSljNqJi3IFy+uxCpHr/bLkuAjneR
SPgFA80aF+threVz8fMlObx6H83iu6exg6Ox+TA4EkVkoWKHsXJYcOgmQTb1FFUt
FkBrRJlLQakzNRuflT8rWY6d4Ey8NrjyrwqAydW69R9H1oRt60R4O1KN7OPYClJl
ywjV/jO7IxUf5L7SQ+27Z/utiyIFbrsUb2yJ6INgQ14EJLMx1tCmR/qcs3+ojNm7
wR8+0Jqu68EBwgWCvn41yQrCowWyyHzPi4RzOVV0Heel4FDgYkX9CKvQkFMj26lN
34RSn5PUX8NoazoJCbU9CMpliFZdUqs5dy5VrlubGyxEjn6NwsicurluOeKQ4T71
CwIMumaqdWxRTBFZLQvPPqays77N0aYpBCLbHls96MBXMmbeguFJP/iHaJthXcpc
Dvr3Bl99Moj/xFvHh8/VKF40VN1j/ocG9is5zLsp3OHiOAeTcVdGH+w1N2/bkfbg
uDJwZh5lzsrbX4aZpjB+y2GEfQTnnRwrNK7xuVQu+T7lEsVQe+zNPbFtYYQAAD6Q
g8OYMuJOpN0r7+97mQ147oLHOgjyAZU3i3V0olyZPMx04Odm+rVsNXF1n2QMjAqw
mHnmq+5jDo79oIGCS1w9NX98zWuv73g7AebzhwNl1DgiZM2gj1L99HDA5zsHVweL
xwm+nMXzymSWGotS2pp3ZJHBI+BTrxdg5anQVTMkL/LVTCwi/cD5liCfzGwk9ynO
4abCFFuudLdh+31EjOwaozotp7ca+wX3zABW6wpstU4tSK2mu4yJImfDD+xEYH3f
lcZXIjzLgJOlzkN+ZI7KCAJtgqKx71YmxAgDOZU4nYNSfkqf5SUUASv/8FweH6HY
i0IsT9HTHA/N9+xcj0XICp0OS9tJT38TbtWM+6poYrOHgwvpkAGf495g5DF4Y9O8
bIzDc4sTaw5SUeDYPvOBktpeV3t40mQ0Ztgdz3AKnKLeYSgCkn82bGnLrkLdmGgE
hzqGQty84la+mqeXhp0EbDZvdhYSkqgDrdwN5ff9ToVCRhZZlWEHoPhpdqWqp3F1
EEY+Rf66M9zUnkWRRAQmyoGksnGxCGBLhCOB8TxLGeCvKus1wpNp+8mj2VhWzlBv
GZ73sqjdqoUZ9gPclHpDAO64e8+rPr3Xdxw1edbNPDs0fMpXHYVLFFosqTWWBWh9
A/QPrhxMv7oQ3N7+39S74iA9rpIPiUtbGc5DKV81ncYG3OChuEJQr0pl7e4N14O2
vlxrW9ePRrN/dyW8E+ck2Eg7OfAI+d2BGvrCfaFWyOSUc9vuGQT/hKqzgxszIZc0
e4iTuDsxmJ1yGNdhuwbBmCY4pgajSbJoXnFuqEnt22uYwXXPPjHcs8TjwFU8fkbB
A4qp2ozr13Pmh7pj19eGPao2odZh4GM/zq+FJQBdcUUskcP9u0/GMuplAi0X+cIj
/KSbIKXIr/pMSU3vqqZMzGz9qI9IwDmhZ5DoF7isi71H6R3SUAuePjzonVbpT5By
cPOxkvHFSHPVc6HqPwgFMCrq/AkgL6mQheYy6aJOyw8b+XwpZ26r4BuVuqVxq1ns
beZ5Z3dqUBtp+h8+h+c6swNSZUA7AdsYJZo/5wzR6Dla+AWc58f6tGHZUG9Wdlsk
X/9QANmgo3kFTDtMcUhfYxz72daGc2xK1gVmtp3WH8R8D5B2zvKop9N1vsB3biIX
ZO6dVyaBshsRHF7wW4h4JSTyJRAfraK0zucCjZ1f+higRE3XCZlc6TOavgIuKrj/
Ka2STz7/B/yXsnidD1cIXuN974nRz1VJZixKdej7PCgNMN4ilM6HQ+gLYpI0iK+v
5PpCBKs45MyrXXhE76JTh0IpKTyu2BIp3ekH1Tvevs2ndEo2IHAwedidPX3LfPHX
T0BLptu1aofWwpUF301PgRoc+twlJwQQ1AiyMVI2OuEH987WmTakRyF53k/rUOYT
9naf9+1SL9B7fbW5NWm2+FgfxKL0PJnPYcaF0AGY1f4YmIFPnaN4PUWyY2ORIjTj
XjU3FX1PyE6aHQL3b59TxxgvkOS0LFk692N57aWxVcSvLm51wtnO+5vM74pNGI31
tmbjnSG2+x2/GJ/lxYmHwS+n+l1A9r81JC2rBRr41N2dwdYIsOUULOy5H6NSLq2v
kk7Sm2gVBXpJtdvJwv1aRcu08gb5gfYDjnX1cMUE7OGwO4c5EiXG98ur5JiqmmI2
Zzrh71zeVsFH++TRfStED76wG6azCuE3bgW0mBta8DRRF03fB4p8amPeeI3FzrPR
cVbS5rqF2oGZd85q6wjyA6zw8ArOifSxGUi4Z4OOGPsNJwGWEOq1zXBNwVtY5h4U
UIcv678gVwbQwm/KOLdUffsdpzrdwz850TRGmyiuLFz7uJ9USgltM6PMVD3pCtV+
uv/lKRrd2P1jQ+6jYBU0IP1ZZTFdZABHgP00HrQug5ytQG78fdpyDlMx+5xPF+zM
78Iysu73XCfRcz4svYUHtjWrIJd7cH12pC6I0u7QJxP4fdaSf7NYNoss+/CrJFx3
I0dbz/J1/bdWW/shyJk8aeMCVwIN0uoI/TQqiC21AJkEVd8CX+zscmJfmRng9JZW
K1+s9vGas1gJwmXD7gsgP/lTfqxf1UkvIHV5Rmnw/ujSOh2hN8CvrPQdItuk2cVu
1qrZRxtPXAW0GW448LHO25/KXw82oG9jCl7gUj9EpyCLOA0bwPpjEIGFm/lK2zbR
5Gg13l6rDclPyRPTFY5GSvwuGZisbAXjNUcyn7KDqZyA3RVDhx8DGdZxgv2V75w5
H/ykucKojkEFmwg4cR2mMIluy3tZzNNaNiNyfZpqRQoyChg1sNpdCiVEWqKTzbCg
m1Vnb4GZ1FDgPy7war9aiDSqufz7REtjp424rGHKV0za953jtmG+qSPCFU4euGbc
OhunpYlP2idce4VGKhXquuPRt8Q81oR2kIZO1bS6VCFZeXH5b+BD528EOaEn6Avf
kqZKq9ttzR/OFsxhgO9Ffh8MPLhnaWCc84nDfI+QZ8nmP3ExJ+kmCXQzzG5A0yuS
+SXOeUCwGQHxBOvYqASL+D3NwJ40ZYCd82J+8ZrvcUAoKLVhMCWYT4YCxODiwuXw
4dj9lN/8bgxYycC1vOkYZuJZgqI8RUIRr/eeR0Uzt6LV5bNHC1HhgVvQWO39K665
FX2ZFbKM7V66BWTiLPVwCHTCpG0FDWqTAn7Wmqpt/aJt6krssrtpCDc4n0YykKlq
PyRJmTdmfk3bppRqPcY47H16gybM0ik3z6LZmjAHsoMnaOA+599gomR2gJNtTlsG
/Xafhq8fYrDE6Kdhb3+7veK9j+qscPiMCkawLzQo2qHTmikaAXdzNnl2f/9gIRFY
MMs1KMrJD4zyFF7JsqrHyAuId3EZkpfySFC/LBHfcLPTzoOQkuQOrQdGty3iSxdy
QRv8R/ZXVhz2NfrREEeLL8EUcoEReJnCZRslA0Dq6ygxv+KPr0yC5Apn1McBLqca
qVdwf20Ce8/zRmBpY0QQbE+wvBfUcfqt2VAlTK7fjU9AzUY2/D91z2xi/RoUnUyA
zzD6IJPBfm0jIigRvu8qcvtssiDg6b/tY01KlxaUcK3FaoGpGftL1IzDk0Kkk3Tx
`protect END_PROTECTED
