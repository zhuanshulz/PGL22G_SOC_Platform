`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ay7LNhmzJ3sVwRjwlTuGSHGs4ipOi6Y0T30oWCawYv4AbzgPjfZmYX7sMYjls8A
Xr1Mhe/hev3X+FB6wIsK+xOxFAefdLByNwJk9M0hVpo7IcqD8CHAFRvXr12pPuPw
tyq1CgUifSWuCTZobmeT3Co5gkeWrxe4X9RhRfXWucAFzHxT8PNkdjFSChaFFF3c
qO4GgmhvpCZrtzFcIox1K/FXjESoUMRrqDEDHSs1otmGQyauQCao5qz4wzOfZ+4u
UaRLhV3Uhfh9sbI0OPhOm2d+uOShjcP5lgTQBdaWF90GCWtAKQ/py+qLQPEmBygV
F2ob1owbjC6e+otQ4wdMDP2Ov/Or0NfiNadqVJr6RMywsRcixkT0lNFZaEsQC8FT
bFcpLHP8sLrIMGcFNui+qasD/KlJP3NfMgQ2xoQqt+8=
`protect END_PROTECTED
