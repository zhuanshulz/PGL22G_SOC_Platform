`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TUq+89d853DzAG/cTG4zOZZnThIElKXho7nXrYF95Ir6nBv4ydaK/eRnCjoGso2i
GcVi1VrsGbiDNcrVSVrIFnwhTfB/Hmf+E7qxO5yzURoy2xFhw/MQo1w1uXeuARkA
ardTv1gf87S/hiWkB+OAk4xBJ8jA2SPdREK915ppSyi0iig8vMyngLxVVEk5LsXf
LTqrswyW0ExP/ueXF2hgFwKNs047NXtkNiUYgPhlGGJCQHlD+fQYDml3vANe0tn6
HFAb+rhvifb/fBftKtnHHzgJhI3mM1CuCvhHWUTCRMAtUYW6lEUotJVUvv972brX
Z2UeEBFGsIVjq85FgMTHU25hlgLZD4JAU8I/uZrKBsBVOT2honas9NJ02dczQy5O
fOIoDDc5J5U8zSUfRieNlh79Hu4kdEyUMSFV9BILxYXiD61jgMVoJ7R7t+RN5udo
yhIsGLGxXmdQ69c0XDmmF/nWpX0Ilz0kUqTnVDXarJ/hrtoUVhNwtqMa5iMxhAdP
Rz1dSGyPPDKEtlsqSoCpq3fuskFhaJPtuQRDNvXe/MjKMcgVECxR5f0jS9CMnRid
4EWWcUnNz3JGR+gx47FJyAlxCnopCCl8ejpEdUNH+8GfwkdeZOsKqioCGm3iXus0
YWONF1Qr2BeJ98fX6sd4DXaWT+zYTUennDhtMuC7oa0XTPW44YagFeOH2eeKIUl7
VhNnPqe/h3SVzLr7xQ+V7THUj/9KOCGjRboQ7/tZTAnFIPocKj/8k9xR23rIWQ8G
LFCXWj3SQlHwZhH+f/yYw0bsoUGkO+ht+bOywXYbDKcyEYQ9KufeUKpZC7q6XQiF
0sROvd08oN9+L/kguWtTvsEAE8k80JYyAy4XNGBagVmXOAxdjTx5IgEmummhc5PS
GhCUP5OItkr85Fqq5EAH3mlhAh9Dq6vvws5U7W61+w32rnKKXGi1nwkSmeswUQ6d
O82qMyMApk9yTVPmlrKk7EMqB2K6lOwN3s7LH8vt6iKVeKnUyGAop6KfLB2o3x9e
6JWjl9Dqf9JMJsQzVj0XEKNhX5blt3dSLJE2kRusgr07oa8WF68ANQOESbQGU6Up
2RUTHpTbzSlrjOR7gOUVfQ1u/cjpiSv7pME//I7ShZti2rC1K/DaceqM0PMT/o87
iGBVx4Z3neYE7z1K06qGfh5DCWxxJIB7uAuGMBTALyxCcYGKScFmcJWXfLyIkjtY
b/SMCuPLjzYPXZ7kV+VMuMO81v7EKgAVG2wfDjAZov3dZxGuPgceNmHAcGIQf8pS
ZA3hkQv4FR9Wc45z7wNs2VDzjyE+ja5iGePgnecQatJVTutDRICEmil3tK9/2XPz
B7IPewazWIS+v19Bkq6ajbRqxofpeY8TraBK7x/dgqMRmbNFDOQIw9jjzgBPHRx3
vkiAFQ5hpmxEVPUkI8LeDxLJCM5zO25xZU1/yg+PBjF4p881dtWqbvAS5sQoU282
Nd4r+897Uyi+gd/xmhmDhTq2oLVQ4fOt5UbmPIDPhWaL2oKZ7tq1rx4/VO8LDCGq
KU99WAL/SkmauWMkv2STLT/bE9DVkO4ihwWbkpIaj0mEodk1ujWoGvxpTL6UIF8b
QUcxaG8dxhAF0OXlYmhkN3vi+ZaYD0dzam5+Zt6PfRy0NF0Yg5GQdqCdzFlqp/82
I/YrAydpKE3MWbTURLQWcBiIExq0LcavNyzS7ZSc0MsIScxqFG7R5xZAACNtstUy
rzoh02J7jwPGDLVn2Qq3D0bBnuzfIQiGeKCG2ShRGaZ/BW0MADQ7lMtcqi17Kx2j
8bjtFgyRU+yWTAcSDfgE74wn5a+v4xAu9Et+u4/IZW7OKoGXDg+zGlzdoKD5QJ/Z
CXqoIat7oa/u2V/QbpwSyZXp7qIv6ah3ATF1+E3kyCUALX2hGEyzOr0q9VF5fYev
cneRMpVD6fG+k2oHwsVuyCyLFsBG534VJRRNzHsIRyN2g2zxXpvO10Os3o/3M80G
6teoUAh/TmM0wfcmCE0l7wMNTawadj9tp0BHJUUVFisL0QRtzrjnNlUk5mZ+ldYw
tFd5gBm0TCQt5+Eb2hvawSIVEmibNkBZ9O9tBr0USY2kkNELut1LE572pS5E5GI/
GYtd7zKLJ5YiuTY1CkoWfFqIZrvis/NoG8cN9IEb9mJclhMawL9wjiocmW0mJXXX
6Wij/ZJyhNfaFnL5ZNxGmMpHzyKS4HUkTYKaKXLuzVRP30zxUFrKVKMsylKMMt6X
mKcSP/tuRBiz57Cuuw24HE+fqzYjBwIDOQjPdec/hXHK6quuMHssd6BULPh7DzXC
aZ3wM4vRtBdZ1A0jdOEDrU35jylbkO/B8g/pfuDezQKvpxDdhmwZa3Vycm+UbVbi
8srKlBWwZWGHfP5KOPGbkY5RNooBFqtijOzxOB7GIobtHJ1cRgllGE2OW4Fel8Zm
omPvoXB4BaVM+ZUKaJbkxIEDLIIOpI9XdTK+83Xi4a2fK2gJX9YKESokLRHwWT4z
2vcyJQ8S2uZ53ZBLl+b+guqmI90j5ejGh5KjEBmSR3mKxbRmyKK+vatjCBs2iulK
BrrWYfWLeW11Me+ZCqp20gQ8a0Az1DA9MFxS9gOA98OpUGG3FOGhubN6FRPVWSIT
IgxgspEga1jWjd6yLCLnl369KOVqBJov9Fm49LZccdnJszsF4CzIkycDkVzwrMm5
DvgiD3M+j/yM4WTOV5RbLjdANrTv7Q1xvZScYXTJdfWwa0dcPsWqy5wkev5VLkMh
9A23acpKt3QLrIKL6srcf1n+cc5ww5UN8w7RbIrDuC1+MF/1LmDVYkJD2sqhyzD9
touEY1JuRC29MOZwpDa+Kh3oh49SFR6+bK7gIr9cVHSD0NUYOqxkxDGpZkzXihpR
CqS3pCeuoEwb0K5sNuUDzMZ0zJ2Sn2Q0hotLXIB1bT/cIP3R+LJluf9YyKPxVNfC
IwTPndbFC4wSZLsUOhAowmnCk4svBcOh8Hokk8YdeSXS/g6wsIjCu/bw5tdhqy/K
C9Kn6lLH3JZGT7JrDMicpWDeW29HS8hDA8fkZPLAjJxvskTQHsxYdy6yOQlO03Ix
zjVkHDeLAQ30swpS7Lxt1HYtk2CSWtp42QW5wQG6ske7MnMcM3uKs7z+3L0jIxgQ
7hGKrZh7QsynQ5+60LhC39kXCuRFCwBteGHs6S2ICaXsy9AVyBg9F17Xd/qBe4U7
7iUvT7LTHnzQ7FdWLKCC7XAwz0JW0wTiMQlL761oh6NqErN84sfeHs9JVBO8fDdU
5BywBs3dVvPDOQXmCjlo4IQ8h6rFlzmqgqCWQKpV3mrVHLwH+i3IcJ5hvodzxYIo
eITiBT7UQj3p8t6M8Td6GnbJ2mhWDspoQyUUQp/AAcS82PJ+nWaVquR3MD8j32/z
hfg2JuF+9NKQU/xa4V9g+/ut1n8SIS3v1y1xKnxybk1n0hkNW3kHl+/FyLulAKTp
W7uUTHZgd6SuXhSQXVNxbsHBmgPDa+CyWPvCOFrXZsbBOua91gzSEvQbDTruwYjy
DpMdbfVuOigL65RkjuqI6VxaiUSW4VGvvrGVWRN57uZRUdQ7soeyqVHcTJULX053
QiPyNc1E4aWpvsdAUr/ljqb4buixzYPTpvXH+UFTYL+gWA6Ndk9OkHDuLbEryDFZ
JT/2D+lYJ78rbYeqniPRTTvazAD6Nyuscmjm/QUu/f4W4xyfSYSuR/tGg6Kfhz0n
ceFQ31T735r4MbM8YYXtpAKpdSSnnqUuf7YiCN9Acf55LlRgb/vtL8eAYVYb7Zrg
qHnE8K7T6ExTXuSz11FkwjrkYPMK74isMziS4G+RkoW0AttTxABZECU81ZmMp1eX
N0Or6G1jSjwm+xfNF0gYYQjTYgPGlO7D3b/f5Mk3MzfhISTTq1OKSXfWGjuc5BbR
zkmYJo9oULl4U6irqc80jIaYuTpuKfcHef0BSnSRLb6ntC+R0sNF9ks2SxiV8hRB
EZyAJJMHQx0L2JCmQZUJuuciBZdPI83z8sAN7jIksRJlW4difj4BBWsaZlx9RuA9
Zu1PMjFtDNdKZY9o30tq9eCLoQWLeUzGS6rYGVHtrGUV9WV0Eh9wq4/JYAl4tp3F
wjyxx9NRbOMYKbvL40JyPwXtaSxPe+hMexn/Ntp568b2PNLEMiLGzNEphz83r0tE
s9N+iPRl5wtNcGma+rA9ppoo6EBfdLf4RwZ5QMOGZVveGKAw9UxbzoOvFQgnV81s
urabNgnFr/YxjdeR0bDrq+EBvnnMcnIVbRbGdy0LEeA3tXbZ5XRPQUw+LX1Qf/zG
kFfh+xsxH8yuZ8z8IicQthQG6enEHkXS/D8e/RRbjQXvisJFQfHtp2f9L5AP1HA+
GMmQ3pPhWJV0Be1E7Nig/6UIxSXN81Sc2q6ug5rBmnoQCzOGVnOrGbb+EYrfeSn/
rr57/DeLe0PoniyPwNPgWAKFAa4lpDBK8fhe1pw+sdwPgrLMpuMSVY78Ico0HoNH
9DCJsDA/toXGv0vAsRliz1h4PMjOwGhu/kkXJTdhNB01tm6qcf/sgdmwkQsNchoA
yEdCsj0VXw38PRFj5cg9E2TX8q9ymogD4dDxto/+OGorOCH9SJ1W51kb+LxHb00G
caUjZr+cXndeM0kuUGAvHzB1fMPQmfYIwipZQYF2raG2BTy4rRG+aUuu8wcuCpcC
NIDDlup7wijgNzQO4a0JDndhfxmLbBBvsCjxu0srafa3Y3qfb0cHpjoMwNl+MHnX
7/gWQzzOVr7DstdXiPW1vuqpevdS7rs1BV5PyEQJjOabg/rcZRKLfW7WUUy7Ap0Q
2Ou734z3T4m3fifnuUqwFU//RP/8nqyC6QWnm+kOLPsopgxKHWWdwLlyYdynV1NQ
fpg2YHshc2h4npCWKqqiqiZIjH1JbSnDJiZcE/m1MjvqbINcvhxBfSIQwNy0+qAl
jfcaijuD8sM4fXiA+lGb66FbaeV7qevqUeUezpaMeABUyP1Ktgjf5C+XipILtrFj
TAjzuKahhd4SNzHIyoTuExPPh30Ow0IxYn43XgdQA9EBDEqpoaiaLRuTxY+SjfhU
UTdrG4oQZtfqebIkawgnxC/bzDCgpnwWzKUXMXirX3JNNiWJEuAF9lNSZoeKmOuG
dTA5KsLDadKcJhauouT5dX6AZn2Jr3iu37JL+yPwFijYVuhNb2AVTZC2g/ob7V6t
T//yrNx4on9JwoF0EAIzHW0FwnFo7A/hnchMbAssp3GwjCadj5cUfH7DzgBCAug9
80JhxbeS8kXTK52PSJGNwb/wlAPRxq6QJSejpEZNYKPGW0BD1WWxoaQMWQ5Iwq93
v1pn+Z+v6KxEIIZ2FaEd6vHxGaFuIFMb9W0tzV84jhr6fuY9YxycK8r9j6espMcL
019n4xAboZJguHTwvqMj8cMK/fbdgEwgfftee1SLWgwQotHUzMiDejuo6Bc0RfHN
bzFl1OSn2KW30t36c1McN6CBOUN+Jmoh660IYkz8om+4PATrEfpRqAE7aFTRUUUs
SZRwQ0AyMYP6xouQUWZzvgJVp8/vkYfI83/7KslfVI8euw+K7rlwR/CwGOWY7Gyo
qEswY3H8DSNDtQSXg82XYK+AOAldmDklkXIFWF4gOYDT7z00xNCW5OuXwyO+9Lnu
I7dpUo6S0y0hqSl/GflHfcGYZZ8716XDIVWCG4st7YV/LFrTli2nXKuoaURXHg8G
ZN8jDTGdfKvGB330BFvlAC9+EblwN5F5hbYXaCZpNhOpDMnJrbLcudUUDwmgBy/+
HmJZwaBEpoVM4CISQ9ZEd7sn1XqiUftUzVHvjTtzY5KDelOlEhe4CN/EPAA4+nXD
0Q4phcaec/VlUZqhmPhZ6GY9jL21Iwq70EYtwnBtQu8s/5wosLtJs+HOeaoK1Eje
zkL3HYUsalae+IUxZZuF+27cW9utXY8vQyP/XPHfffO6uEBCtRTnt14T5T3Mx0MS
kpQzsS0qb3UaI+OSclz1+WFYMMppWrZWrWCLOqLgbcClv/Xt6bg4bj5swrFxjFmz
2VKO0fFTUwdeGTDjquAT51Cqxd/OM4wf83Qe6nFnuiJeof2GM/zy9rymespxtsjg
BZK2bAoHuyfKdtx3gbYkybBYB0/BI3rtsxRi9YsR/FglJoNWIyPlFAVv0urXNmZl
oRtDz6bjksPvyg/TSFtZdVVUrqfIsxTIALci0c4Fa+1qsTUEoKmgTPRA3fIq4NDJ
+IRZqqvlZWeCogIIY6HE+KEYAs5cvjZ/qy3X7sh/rcH11zUUdh9l2Xc85EO5IVlA
wxbIJ5AEe3XuTCJVtuG4PPnWPs+P1IjdwyzNkGCiEud7j66v/W41XDVeCOLz4R0R
CO4lFS0r5qGqSSl4hTpNXG0VvL++IORmpTh/OMfgSUQL9GgZOYH1XKgAqQQ4d10L
8jFK0fGQSFhcdztJMhrrXEclGaIjHkZRsgOV4Kl+fvCf14PfTcGWpbrDiNWejjiu
9twHlQlOZEQZGNHs+9yzOeLbhYEooBkE4PtFNUNtff7sPXJk4uBSDCfD/y5F3V/E
ZEcJK6/2ypyGt/rqu9kBHYWvQUXlNWmtJcKBPR9egfyONwWorhRJ+idhh1e+MlX2
cSIkKvj8p7L72T43Oc7Y+WK+jIcTfjg+L+uCMhIhhJW95PBEAQU5b2cxa+vPzPLe
JQDGxyXxRejyl9Ty3DxwEbOyEomR2DvLKt42VGg67bnn3V/vXsjs9O1HUtAWR+iO
vszgvZKLXKvcZFZ9K0aRgBmi5U8LBPdGOS7H7PwaNHFz0ZGLfxnwJUfFMW1I7ZQb
QCtkcihhNwIqn2RFdWzmmcQwYxosSa6jxxZfvtw79+CC+XLSr9x3U6WmL2p9H++d
az0byGBTIboo3EuuV6U/39Qwidgz79r10oO3hrFtsLkzD+BFrWH9dBbGcfert2rs
7fv8xZjPd7L5RqxqRAPfiCKNlHoFZTvjvbQAmEAZXZBaeZHSP0uG6YbPaStcknLP
kGgvjHOjbLc+JQbOgI6BmcRNtBuiPVo2V3YQtyD+B00KZKetyvNmP3+8fHbmH/aB
Mfi6Uyv/ikMvImQn8MJ7WcQLKfV4vAopvh5qf0AzRhnzUtoCYTBZltNKar17Z0c9
wyi4D43gbSD31YJwdt5a/6tSWJj5vweNgvWWp4ibbvftwycGuWJbL2nm68PhbMAu
1nlg9Owy7aZBfJNvtPDuUptJM/EAINDcP/jRxVm9Hft421Ll7w7QjLb46q3IgDVn
qWlvQM/vkKtE+1STys/zDyuwvgd811EGYxv1zw1yPnllN63hGa6+ENbgc1illwEG
h2++6neX+w3LCcM9BhydVi3LqGKWwDJt6cfRs4scJCh47KyyuvUPhb5cRD8Dvk9f
3CQIKOxQ1Zw1lv8iD2Py5OIdDm9kk2Qj/emoNN9NrvZ0FqBEbIhwBNhiwJlVAMAZ
+yJTkcYTkxRu/fpUJI8RVuwQC0KnRGswD+zZoJtEETsKYWO0G/Dc1q0jZHgshN1k
crzJP4cw6kcqf4A8ORtmjUoCldez7uEVjMv9jUBp2ddcYE7NcDSLZGsyGtxDy+bo
wTE23LKnXB+uxdq29tc49e3cfX8ei08IHrM2ikU2SPE5Dcw0WfTxRB/eVwHV1Cha
PGEP9FD7lxTkWLu69xLsBZKDFwEpcCEDXgdHlpKqiVy0nH3PaTkn9w/Cn3a3oBoM
VBI9AWTZAzP8ZIgDLv27Y4vdpEI2MnN98WzcYoEJgajubZFVZpktWeXp1jKtgrf9
B7GY057TO0vrS05ichDpic76W31WojiIyUe4DkHAw+UeSmRP27g15c6eC5zWRByC
mOQXnOBwLZ8J97RUedLdwtsey37og/UUMtPBGWOeCFAPSzHw0vzctSzFoWsakECo
mz2TUDKPYnONr27HCjCN6ebx/3u+wHme2fav6RSALtnjbi19aDuwi20UtsiP0qEc
frlitQUm+yYqmoKaKOwgDA9SSe9jxHCh0gpOtfU/mDY+0fWOKfloHfSVI42t/UUz
XlMM3hD19bQs3/9tc+mcb1Om13mxrZT3M8dJqUVE1NaU9eXN0suYDk1ZCI+usUgC
59/qH4/IDjG1r8EYNEGL+0XiJ9+fbn0RFk980oUKgkFukhtkrX0bIgF7C/+sFF7z
pKwLd49MxFVdsoJcO/TJE97kXc9MqgWv7mO1wCtfalMM7tMkQDxbZctTRGF5fBeh
Wyvmidw6g6lZ6OLh7v1VXHx+W6bPWAJ+8OlgmyOkphdnXU24rSFNgEFkJeNVZWSg
IJjj63m/GTJQGh9dQsrn70aerPWTzky/2qRzr3GTHz7dnARTInvualzyfuFddUDj
vUH0aN1b9Q5LYYWcxH1DyhBy/g8nDvA2LnLm0TQRJ3AricPJqeIPgyxpaO5vGzsy
yd2K05qq4PCmXBZ5V7604GCz9RWl+W89v4qVhjD2rfVCJqHSIARCf3BrBI6eJ3qY
KOlukI6SDFNlkjwcfMPFnDsMp1wvh7lrRFDeg1i+PmQJ5kma6tDBH+e9Jlw/++9e
tfyshATWHdcL1ddTfj96PnsW3DAvY7qyYDHbKGby5e1Nbdlv8cz/S3U3BG1v5PgD
FeEk+L1fBsAVF71LdtVIE9TPWoMclWrer0aPKsVxkL3l+BDvKi7v6zPheT9RIai4
4FUQHuVET6zoHtn32O37/K/6uI5HBRiq2nCeQZP8p/leEFyb3Q8YP+Zs8Men5+56
zEbAELqmKsZ/Un3VvSaJpECAou7wwe0BpeaguCGg0/JbUEbIx/Ni35Ga/4yuGfdG
0uWhF1I2/TL4AVvLBc/XydOQ1WDq9u9q65i+OYAyEHBAZ+myBGXeXlhVOvxO5YCB
CdVJsHR3Yqd3SxAIeti+wGmAjJUBnWKxkQ3lmw7r5eKTbgG6ziLZ88v+uMlJJtMz
LCWmB3XbrGrMxi+1xn7CKPF1WY/RpLqXWTSTNglWmschmJn/VO+NGo/cEMegZyBA
kVaZZJlC4c+I4HEVs09/uKqC6jo/YvM5mJqbkkDDG/yYvTFUMuobQ2m5PG4e6M+S
e8J/Fl7C6yshqLDRbjMCaqLMTchtNujoOLYgQCVdjVYpEVw7/3C11aLNqCCQt/WA
AXBa7wyg4/7LpoafAYx9v9XbMG2VVPHqJ20h4iD0QKSGFUkA44uNkE5f8YwEUDFS
7b2XQ5qE2ErCAZCUoHbHVtCF5/CqJPSA200z+YK9w2lyHaauN00x5Ee99ZCU7eGt
Rd4fpmd0qTTLsvOOiV7gAMJhzRpdNhMQm3RR8GPp1u9+al0Vdet4bMODvO9D86do
Y1v5BkKFlQ/oSsrEr9fPjiQuzRiudSwu7zDCBvac7ai+b/9FCgNtLJOB6wZzHl0y
aI/Fbr6MXtXuCsKRrcnDp7MP71UG+buBrJbA+lLT1HadaZ7HrHSD6h5EVvZbwqZ4
I95tN5da8b269RjKqcHNuoSy1zy/PxLyW6Ks8U2iZW52kMDq02K+BVvKKWUaA26R
WgNj6agYZi6+yrfqCBjorAwL028FBcdXNxvGarswu48Dx/IBPe+vorvFC5Eilk6Q
EsMmeSFkq2r2V/6abOMSLjeL1gkABpsUI79LhDTBmcJi0p+4LxE3P2VI6tWF8oLv
N5VIUK0L5FA9WCfvCj5u4dRelACST9+Wrqbb7HRIEKGVuR/4MPxU5hIYCKIvwl4s
NW6XIgt8eH/JQG3w2/FzZmaTxf6R40AjrotC4I4j/QOLA3mewZIa29xZ9N0xy0wm
ffl4k5igm+12SKUJF6COBxNh5/WQcUMqnfs70ayX7Ry25F/gFdY+l/0gUqDMr8Jq
DDGVmm0d5IUmgHzFh1E8ikQc8EsHGrtCl+8n9J5SdQK2y3KdZJxhZLlAyO840NMb
KZAcDWqisYGNNRi/Hq4Ql57qooj4bu4j5qLzQjzTm0ggbFbuSPq6+YXAGBMWZfCN
OdHzc/YRt4zYfQ8+9tnocivn8KUtsOfT1SsFji5Z1KBWdHrOXj/Zlx5EbpN1dCiI
4WxeFZubgru0OJjq6eJmc3HErV1cnd6nXzjpVwMaAF2i4wEO3hAy2NWfHJU5rXcx
ShG/+ocUY+qYeIrnQqvHVBKzDwvqLH7VYsnsqthJrknpA+cqYCapKNM/vbBkc/5R
yaVe4pVibkTdFg0n1qvsQMtWLCjXIRr+L0CCdhBEt6NHgNz1Yiuu3m+vjfNObMxM
y5xiQp6rASMSY3HXGP3JJ/ejXZbAibzMhWr8/s++q3BK+k+lNR5pAahufPajiRdp
Iu75OXy1vcN52bAlKolo80EwrVW+7Yr9u0KB3FU1CiM/lfzydwjKhSICxX47BuRh
xtppKx96MmliIm+UgkhA4PgkI0zzPVfx5xuDqVrJnSs7UF8RMvTom4eMPuhqtnM6
rGmjvU3rACckkWEnkgWZNrmlSFMAAO7Kl6btsJxG0r2Bil/C03sh2tGU1tXx8YbS
5B20ASKwy8brsMeuR5ZTN89e35SNzAyQ8ZZj5v9OafLMnsLgKvR1bIkwt41Y1X+C
Uco1meQYHYIKTg8LQVoQYhV4a4bKgfC6YD6/YqNy7EtGqosd4BkL6ss5iQVWnvCZ
01Y9R9vbZMeX4gD+eD6/GwXhjf7MFVvqK3O6FNPZcI0+WkDVlBtdXO1RP2f8PW14
EQyLs6nkJAveZHLeDI6CIjUlnXhTQINL3L79KPjqYSDL3arZH0JBXTn/xdk1JYE6
wo2nuQMJK2oas57hgrC8KvW9LXd5tWMJ99W1vuQEUMoHXkx4uPojoCyCmpKH2Fbn
ZVXXf3eL2otmSefh7PkwmrBmC83277aethv14UrCJSTHL7d+Rf8zRJx0vCHpW4m6
LU9u+deulhP0/ZTVrfrVdx0Hh0TWTF03L7qzkwgEbq61i+jG7VzvicMSXV2oYuRC
jgp4ci/3ClrlRpv0AqgaFdV7v95TdIOnbSTyekYwInLiUYP6oJ8qAKZjIDGLs4tq
q1hWMyGKV7Ou469kC7JZ+OxdB52ko7hjKvw0d/G3lYRZP1wNnkc2yT7v2fVGDxQ9
caHFPWypj93x8m/jRUC5pnDfAkqB9Ea1QLOKS31hPNpka7U6XTXUAugXs0v3CW2b
JufaxxzDWzQCFSsFhWEIZMnYWEZlWpmCJ001rV/z27uVMmuoGDMqcR8Y8y6bRMTW
5Sx3Chpn7X9s8ZOWluMOLoYwpQQbW2XXJCWBrqgs3pPZ55FzzMNmydx5egGv18dk
KEN94zq7bepqVyF/Tng91MMMjbIa84vxh8sQFoipJzZCt7wNfrCWY5rt7Q9F6SqX
xh2tmfQnK9Iey5/Pkh9qDgXCuhOGdT7P5GWXOSQGL/MogaGzYTGvgGbGvLNXCzVJ
ZqOEv9lMmhuW7Gzm5VkhkpgPX9UU441lcUdslWWN02Wvjp48XXuqzcdMH3HAigl1
ilcfn1UH0lJaaPyckd/X8n/dOzUCJcOf1rcDriP6IYrRrHTAxSLrnsmuT8vuJMfY
HhsSgX5IZ3pFsOdHO1QwqTpwwXvRksnOPNi2L38u/PIscc3oKqi9OaaLvWdAhm9a
4L0FUabXRFIJG//W2gxjywonZvQHno+ddpvCJZp+dC2HDcGDJniDg+5vaV1FS5z3
h9bAAXnTJ+yAU8My9VhDvknDU0L4KPOUHKuPE0XkIhDSArej8UFcKCpbx9BCMvdH
8Uvm8wRLn7k6TghO+kZfbOioJsYeHxDJwlOHr2MEoS78f3INZkpLVFELDbd8cKrd
+2sPUZQYxoDzwHAVcULx/S5EF2dxjOwomG234kpfM2bxbDsULKYfw22ftN4dqx46
tINjpZnbV2Ow+zDigryA4DnYWPh5JhDhdAsmko95dOABaGvLdmo2EFYXd896Ly5D
jMwDNecVI62++ANAlRC9eyL8CvpAP3S7tk8Tj/S5ioM+LGPJX38nH9W3UIyazSB4
nD/YBnZi5kNuvty+dPWhsPYqTi1A+s4Nocm76VwUFgnaNqFDSRP5DbGR9Uuh8Y8m
WgLY5uHjtJI0SEuywcVDAVP6Gs6BaFYc+9OqTjVkwbGEf+7OOHO2jM92QxWWdkG4
+n/jwNSEBcfX30YbPApLUx9DCEnTJ5xGmPGqqvUnAuZyH3hXmZyatTxLpZ6ejzQ5
s8jg9to79QNt1o361kSRt3hMqfri61JEk0czOgCa/4xiopZxy9kHJk3YCM+Th4O8
AEAgD/1MdYaZNzfFMrew30T+hCzmJH8k8SNR2AdRyD3U6IxSAxEkjcElIrkwyH1o
Y+Pf+YcoKt3QSy/x1BJkrDOE0A/Wo5w5ncvhL6n2yF26Cx8agkk+tpeQxEbyHjma
Ww1FKymFMjEWxmg+Arlk/D3JVXTYfTDd+x86lr/rngzTRsO6IaucNYlfxjQHD3cW
77Txr1ZeL1koYx74XNKx+6omS2GAIOCqBpnYqGR4GbfFs8TFJfhGWMpWkjQnkcr4
NWDgwteRWMCa5EvYTMm0Ek3G3fp2DATdMTyYYCvkgjoLSLjH6OVOJrKjegKnTjaU
M+bPeo98k7OrxcfSnwMVCtbrAADXjVHjPPGfVher3AdJbonRA9+Y02bgmE99wzt7
WfWXBvq1YVbLJaHuziBvZ9HQx8vdFOhMGrMgy/dU9LWJXOn82TzEVVMph1o7zJe3
o5QjbCH+ma3NZIzSNg3FoSoaVuHjptj56nU8ujzUIlZvQxAZjvNbA0GDj9XVW8x8
3itJPnZXP+gs0Ej6fqsr6RVJXxTJPPeROxvYP9s58H0GSIkAwgOZVL1Pyz3hlSme
bd/dcTQTgtZvvjjHtbxuF1cNEwj0m75ha8pTbxT9jr1+j6GSBgW10wQlINiHDNGF
Gao4GT2a6Fs/UoAEbXWYhbmzORSbLREMvUcWszaerl+rAU6kDnv9rnQrhrAQtaCk
CSwXwz+R0gUxa9XVF8+pyJMSX4mQfQ0ctocIlNp9mDnSTrg3dCNPEHg2t6xbaOhB
IS6Evv+5pTRBLIGYF/g5dXjgPxgKpJtCh8DQW7lIgz/tKrflnfMHAj/BbEkkV+YX
iRtdl9fxmjOY+MsuK8yJLP4gOLVt39WlikqOKBI4Z+FnZY0MYzCaiXFJBkU6s2Ks
EfLTJ2En5FncovI1PWakZRp6phHiaOeoPi+iQZM3Sayacfr+ChFOnRvodwV3l6e1
xx1+kU+OafWgeN/q66KvYgS7KAsig8M0VXF+aBt//q58CkqPPsSi0NxqFSvtP2yY
c5DOlDSgXGehLJ9qbv6OHQmLDJYjj/WDtSENNQXTfbUAMJ2kUykrh2uoqwRA0L25
qau0G167UCr9o9gEz+eK5orht5IkB+AIgao9UeniIgTqmmxMbfK5XSBrQXJ2d3cJ
hcZCm3p8/+9Z3udN7NRrTrJ4vL9xNDIUeaL5+PNKBWmOVePgMhgSkrEnEivbCMy/
5LF0bn3dYgdbfLl84IZz2W9zXWWSmayFoOuhHqG+t4DGAPau0BIusEfIOyzpkWDU
YV/ggs9csvGSd6mLqVKeFUiHdkxVlSofTl3ykdnjUoT096Tw4BqgiXWw2EwXwDaM
TLvlPj4f8LoUG4gEGQf0wXIBU6ZFeJJKUhb6m9nsQzt9heaM2JpZ4aZREfAuCD6z
vGVOcEKetvBHqqCaA/6k7+aMpDEcZavPrHj2C+UUUCzHGJc7o5LYGt6SJ/cmLdK8
CLtZs+4zdctT6OSdLRWl3kqnxcv6F39N7d2FVPYXegYZM0KL46i4egUqtvDaZJ46
2OdQ3C9FS7IsDDAk3QhnCkAqcqatVdLbUM9tkNAL9cBJLTrsAR3+yDQ3WqkftQ/3
j5hol68FDfTKLczn1cRnAGwLUblgbX05cpDRh5bKU26xS5lZ99wz+U1CWWe1hLhm
5Lk7rb/Mt3mexQPKtkpQ8BYo9T4jdKGm1Qhaohv7P/z/4Mro8bWCVxbwSXrMnHa4
oD+Hq4g+l8KoPQRkr1HnC8MdAET18q8x3/1u1+tZRRbKRENqsvMkSysrkKrAvR23
urqDoYa67K2gm2aK/uKtig4s4b1ansFw6qhyYNU7S1m6yC8uZdJuE05BgtfJElsC
dfU6xEmkcgqis3YJ9LmqlpxEGMqiDsxBMEkV6gBOaVKI8V3XPDFgNF8bZpU7Md+r
tE26rxf5uLq/8AlyZaXyu64aPSX8pTc8G1VEy8ryfY5KKoyIIXg/Y2bX5netBR9W
OYlcqcS24miqZRkUzpi98u8R/UL3tOUVJyX76TFwHwmRpYFW/o2S+6YR2T4QQEWa
d0hsYHvosmFq4lOq/pjPOX1ixD4pEq3dx8Ez/S6+IUIaXAdOBBio/BEBo+XrDTy5
w+vIHD7UjhpVU0YV1fTPWYNZoA5gktYhb8YXnwklnDzpol5lZmbFLPRre3jLyqj7
+TLH66RTKgLL8sROYbgMQD/pmMfTGJJ5VsQhovSDWZ2r4kypzwO04DBObSWuwHT2
+UCxQ2iW7E2pqOM14EbAZRHB1o3jB4VdwMQBYXGdskpOrT97M3GB0KYAOz4nD049
t+t2BFaMNkuYzjlF7UiBquCImV0NNe6OWKix1AAZFCwzMcYkt6i/sfglR9HsW7Jp
Km0o7dJAcjsnUz/J5sIgVjPKVqbhlrf2KL7YYSBH06/mgiu4shPqJQGEdexacG/k
JUDD//avyExKOta9ZgkFRnwtsOdfZe4EwaN1ZvLMQOC9p90PNCfiC3Bk1tSubT1Q
qBXuRh27dr5twtZLjRWLFo+TojLSEm2Nx/rC3Pu8DZpzfE/eobdvym9qKAgSAlyz
D9VXsAqkVTHzuh6WGxfZX45jxew7oIygt5A5rF4BmZJJbda8ywgSwduaMsO+L2wW
DM85eRSqg/CnmFeq1Dur7Rd0rlC38MLPrCswcUaroz19GkXowzr/c92JspHGrQ7X
0kAJBNNMDsA9y6Od14vIu3+KgtU0T8aD8n6SKwpInTLdfm99fiLhceo3b9UxjCUS
SjSSGWl9WMenm9OduG4LHrocVGCs526ujg8EqR8llM5ECdvvBKECEQHmF8mK+R2Y
A6Qcgdp5hlbqrivp9fcZ7l4I6i2GYLIW5oUK8MPcsKxtTKhKke1bJ/yydIANZO23
GwiMn7hjg7ZHUWAoieaBw/ZKbenSIj1HjooDe77aAvSYgh0/RgYfp+w2zsz+YfIn
YRFlPYvrwulS+TXr9VjZH877AM1BX8U2xOSydXyIyxtqmbYHTEXinjZBdGS8Vw8B
+Ig1WMgKmK3qDfpk5NxuO32Un4jLTZHorr0seXUTplcoMyQg+HCM9kahNaNvkFvQ
ruR5AENEcW5HUcuRIUa+tN6vrvJgCsrlMU9B5Ho/59SGj7NEePp8gjCzXO6Sn8Xz
bD8PGqbEGi4zUPovA9RqbzIUUuCZY6uP1kF9Wwnm0rEtWRakhMctARCkwRGTZ/Fa
VqiXoq/+EpxPJbbZeZG/IjLS25bjsIhfPtoOsGp3mWLahmqge8UUSsurIdTi1cQK
lZ/L56/2S+6ZmULbeaqkWeYGVczkyOZ/mtglhwALADUqWAistEhgwjQHBkT+YnUy
Xvdz8kwW2eiu5xTxB3th+D/axdxGisUkbQoj+v+Iykfgg/PSI+LAVhKpcSctA0wx
PEHqWx7aJFzumV2xsAeOAPt7rkoqyOEDbq9/tIsL/UjUK21VaSW28nSDFaDPFJ+c
6CRzyvD0Ul6D/1JqU77EVlsY+kqog0CVxfNRZSoWhVn6JS+DjsbhtE7dqaozGcMJ
AqhtInlP5ecyn5f9xSbLXKArb4DO/QOd6kR2dBrBXOktf2DT8murLHRh1fEo3sZe
NoYQ/XBw7FIhpDVUAgWDIusphmdZ6XGhzJeR4pbhi2gWTU1ASP41h5/iq0o+YHkf
4Sl0JF9rEFEASVMRrFyb7MDIylW/2fecAMSuH2Xqos0SHUgvWHJu1kUUu6GPqdKg
Bu5Rusx3hOCgF4bb+aLOLngBVlaqOvzesrgTNtwkH8BxxYE5iybNv2SD0nhk+8+p
cmsowl/uqjxN016KXm+xKMs5Yf9KBnzCwvwUIhTFjSPrrsZUNgaT9QwZDTWwOCMH
x/EmRuywRxtlFDJp/d8evKzZdvOuzDsqG0Mv+pi64PjMUtDFktRdmkzUiAXHSm4G
3sIa6H958qFTBCGlVb4XXTHxoZB7JG/LNdqaN7HsPPIbCntcPNFOZl2yvO0qXI33
od4U2dNM0DAoRwh0otqhwaMGDkrxs26WCwFchbdOsavdwsN6PVIb70OSRqgJkTSK
7Xxbdyihi+6U9agqmYgvI27uMxs/mQqNg49EHphutRPEOP5B9kg3GdDQShkIrI6X
4pnXduqai8FmwgJyukey3Ztr6m0gQXrDFF1flCNx+p7ZeyvcxO7l4Smy+zhlE148
zEVav+58CVbDUZjL6hW/3FfLPPXAjj9hrT3tuQtVAl/Kq5VyMHLZr8GqY9byJC0E
z/YeEJtp6AGSbZX+HBGIJjvcpWsqbBCVwE998D+RhbbZyqoxPV26rhXEX1yRdSBe
Ly4eeWE2vP0CA3MRqY8Mpnv0HTVisC6i6eZoWMhDA5X32F3Q1kx5UmDaJ49wPnRy
Ff+++IY2Hm0t7tfZJ9Np6kDZoly69IT1XJqFXAVro1jE7Si3pG4vI7RrdjJTSnu9
lPLlOiAEwtl2EEyPJ+A3Ye9F609qaBJFLkMWXiAO4z8dgsMc9fcTUGcZ1o5Cp+hi
IlVo8RlL7Zlur+AV3ZVBSvuLj1q1jLoLKaKH1aFhCVgF3NszAGQFIeD7ZSXsezFG
68WB0iYHvh6csFjbvhaHdWP/hR2yXiBFZ6KMrzOPVnZuFnOxXtFcT3W10lP2bbIz
zHqIgo11Ydc2HxDgHKJMzel4h+4jSF0YAEvygSxOcJFCN1tmHzW5aDDBjL5Os5ny
hAtv/rTSpMXulsBuOJPAe8wva5FNB5wYXWDZKUZVwOT6jjNTCRG7OwpWW+vh1OCe
EB4pDR2XwwKoycRmejNcV9y8o1544d77ITuiPlDsmEk85j5LOUgPgeekaQsLOnnq
3qtXWMHJadyoGo2t61lUpGWKMl5sYRjGbUUi146390UdeuFpUeVEJ0FZmAg7MxSy
GQUAlSUE8oZYDLCJ6oex8DQD75PHsPU5yj4C7GF/26IceOsbKrnFz/hwMHpY4fGr
1lyBkuWuJ+KbgEcjvlfLpBhR0MXT+G3ZISnkRRkzN1koPYULQRgUQCSAZiQ39P0g
4b9siWYO6a5Rxz7//7zkV/QsrCfVUsmgkyLO2mKF25LwE2RGsnl8ArjEXCsYz0Wx
Dr8b7WWo71eDzhy0kVjQz/xlyupfljJlAxFET+7d/B+vHEPt1ElU6eGeZOP5Pzbk
5717TfJnjD2oksIVHr/WV0hewYy88Cmg3N1CbeYohmzqU5Yhj9s56RTrh6zM8HzK
W/xxHQyR8iYxei/w2v5kgWTYDHHF6/elQJrkKOiTkLzBoKDn3m4sT5RdIxRDZ9Fv
gTaR02eXLrzeyKfae8KCW1yJdhTAmwEKMBOkVmlR0qdtjMfz4YztEMW+tFclZJhI
KXB9V6X+xmgGrenjegrXMNB2KMW0n+++VHfgvlH7Z9cWDg4fXAAQCjoQkj3ec1zY
fgwJvrfT38Fgt3WBNL24wp0ezBnmPE/jdEUKUqM5aJmHE7XmzLOqNSldZtABzWlF
N1EtJsT+8kXx/IUTjeZSZnL8S16ZvdOXuPFkDQ1NvCZpIFIDrw8UKHVqWu2hAmSl
cQi4hJ8JuhY9veA1aNYvgvhIdC/+lPHYnV5HbOu3Lfo2YW9UGhb7eh4KIob7CDr6
2gLTEnCwxXo3WQhN7bflK6/HCp1jra1emQHSD9YJsOuicar0pz7nIvF3dvaT9uwu
GnodbUsrD1Mj7dyeTNpx3IPko4PP+CNQpclsnjEimuhltjzuHOh929S2rqDD94kN
bwzeFIXTU1KvpCVPLMI3cbiX4xBrC38qDMyt0E2rTKOk+Pc8tZJ0OYyw45C6WfIL
cZn7VPQlYW1dOZLQZPoL+fzvtVqRIQStotEo/6LFHZaDc5Z9ss0fTunA20S61zVI
rxslCO8Slzkoshdti2SZ/iZVa8B0Ia4Aiv2olMsDHcxSVjDmT9o8dAs22DZ91JYV
OAtPtuMVGwer3fjr3N9KRqgXMUxEoyG41L7ldv9P9guFjPSBCbiVWpBgZhOxs0Az
BiC88BMYjQfY1wo7NaNfpxNalQBj0NydnibQ5M/5f8vevXZm55o2yQc/N9zPQ0E4
Zg1YK2aqeCtcsolxaQcknTpecztVUsu1Khen8zZE+AMXGGocqx6rhHtMHAIJ4ffV
sQR5EuO61zM24z2BWy/oKklPxjfqdkmzHDiOCmrYavLGTGIT1VMjYBgH8l7Zm/2D
IFIf4DM87EgzwRwBzN76MLzeuVCQVwwjDM9CGJYxa5qM0runsyBtrfZoVRSyqBO4
FY64MlvTZ5FAYKSpx8oB3EwcO1M2RBbWlbCMK7Son6ZQuS9k47+kl4tcsKN2Ri+L
ouNMffHeLMQ+/iHUoAvJa467NS3JteJAF/iibjVkUVwPZbwj1evKFFFOVYX62ix3
uEl1p5rqRVFCIwd6Iu5D1V2zsFGrDxsNk0e03yht5Z+zxpdN9iw0N9OVTGWLxQZs
IGH3EdFKwLbtvK99/EBe8p+c8oSrvj5cU8rIB+i+qLzoN1kQNjsJZYmob/NmqoHq
zwdJHTvmraZIqzVuJp+kd8UD/eGhe176GzdTY7HQ/7opLQxVNFNEdPa9o63rqZIq
FUab5oke1/B4zttNGuwd2d1FooC7vqQ4ApXoyLPDmLb6EYxTapWeEl9yaUyGHTkq
kh/icR2KNXt+ERAtqyBV3i9lgbjaVdMex2S4jUTzVdR5IABglmeayeCkQf0zn7QJ
zDKgLyxiVIg6HGIaxxKjlIkdE+5Vot+nb0iQacVyQbVlWbboYvMYJCg2mI/UyLXw
TJ2Yk/PqWWBzFB8KPLHW7DzbCC6LoSb7JfFSU/lJGYVudNFTQ9sdKpXhcnYOdy5Z
u7AhmIHfhB9wKUsvJknm9+8+Uaa5PoE17ZFbbR2HtfAwp4Gj+RmRi6hCRYvbrCox
t12MnTvynYK0d3h9E0ucsbH6H9aiDY2ybOFgHDQv6UA9OMmVdggMKTjJWkjYWke1
CRbGMsHD1hGsVLgzkoAA9E5aKF4QYA+p+eaQL2wzXj6lqCJHM10CzbPORWUIx4qc
MxVR/rVb/Y/904dS5rKwGJjMRusLl18toOgdJKUE4Pmt9YdFUU8Yy5kNHfO2IohZ
AJnbKchjM1pyKnhH64rmK+bLXKWvnf0NTdpCvgX4aMeD8jk63/3XZXqYDQIScJ2H
m8gBtqJXSKQp1UkDlHXtTfv5y5HmKdn60f2FQllQs5tsaEgxeZmOnWux3nylTgTy
HmUtbfn/kIoQPy0aIs51+3z4lYthKePTv5Gyixs+Vfda/1QOYxES+XaX+5PBpw7q
YvEkTX5VOozpMEGcc4Q9M+jWEEIWpjgk9sMl9JaBnWYWeIVAmGKqR3VOgdFDbv8F
tvOmzjjktTzC2RpELUoTHXIWNWSH9zWjMGSbRJjpJMyZ8e2Ni/xaeWtjEsV0d5od
EJcvEvNs09QluqsH9d3I2WQ3myDXaIfEbwrrnIs/PopB+BQVacc/ThySFLV7neJv
LHT4gfOsdgWd1FWH9ORPUYQZCP5Kawd6KLGgNwjFSkqMdtD5shlX8oQz+n/RuzdB
ovGoAG9kK5QY/H9pIgcc/5/cpMO/CmuueuHu/16DAhOiYdYXwMrOr9ekgCMeDO7E
ob3GON9iFX0uQDn1LFfvgqDHYO/AF2Y7OMqgEqbmJSCHwibLaFKdGC0xcLEyJpqq
sfet/A9uz8v5tmVfhtc9ACrLt60aNqjbD20jcBwD1neE192uF3EE7kI7/TilJBfL
QFMddi7ls0kRM4Y2wdhIY0iKWLWtYRnmCWwZ+GL63GM976z6rbEdG0AUcHVQwi2F
94KkAN3xQCcAco1qzb3oJ9sKZPI1QTAr/HcAbd3AEr/FM5PT4h9KkWScFG9T+t/8
e4WDB4vFCo+D0+QdhnCMawQ8eyXWRZh9FB+ixsV3EUwvHQU1xjYilCyWHQ9c1dg2
N4MgrcTyxH+9eYz4UWT1ulElQeBIgBdGyXrC8VT59dP5Oob+BX8451Iwl9C//lO8
PiI9blJoovHwtiX1KFT5MN1hjFDUztJlm1o5CHZSG4rcxgC7YnasHidrDOtYXxnr
gEQ8oqXy2U/eLFyvqUf+JQFsVkcfHHEpeiE9GuyHtcobfPuWjgsw7O5KkheYzBrg
YKrQSLjmkYvnGGb+I79OBOpbUbv1HwGZmj4St9/Vxu+QuNC7Auv9IIFjNd9DVaYO
nBrwxjzDPDEqCBpgEuT2tHIPOEC3OLxCLFCbw/KKoBZoT4EIjK/F8EhQzU8s5xmm
MZB1v8WHWZYY/QPwAriXm/ilxiOC808U5lig8WoXlIigGn+bcwOpS+DW6IkgxV7I
GwgvaxkRx8/9RfJrig9RDLmhlAVRvA/etfMTNVNi21Zpp4at4pijatKnSBLJxaQm
M/dWgtYXUmDZDNsC30I8KJVC8fEUT6kzF01L23T7HtOWVohUC/PIBKRPWdGkDOYM
KGgtCDgXhGV0OTXzhnNKUFUIpV8gf7E9saSyCGNsNz/aAN7Vc70Ds25jbtr0ed1l
mrkRqQzisQhrms/NaKIWdsl4RcmGfqD6bM9eYu43U75NT0trKLQd2sbUlvFg8X/i
Qb7ASfffQs+ReCNBaGnjoPL7m/hecvacxG6rDCSmlClhq6vPSv+icVjofHjZXagc
3IqqohQCZZ7Fri9waCaYdD3HdExqQpoEOBlI4bB5B5B6//90QZQDwZXg4VjqVL6N
az59qSVD1YVTqG1YoLdWfLhzSQMLfsIwUWbRhC/GK5xJ4h7FHhOYTjXjHx+Z9IjL
Ity8+cEClxOEog+q9ICWz3VK8hYocjMtFSlzNLclThNUq/I4FmyYbQ/DTte9Abto
J2+5OralQTglC8Hjcdc5DHxJYu0eS/eGoZkpI0MESdCl4uRRgZV7I8XPRJaGvIp4
IOllQwoVrloWCRvxSyEnxtP7kd9ZZJGs/SgZcOxY9H56ll6BOKtCuYELRRSUGT07
SqBxxuZ8FrudIvKB9gN8xxQDjJ06mBJghTzRL6lyPsJEIcP3PPr92Oeo+Maao4mz
CUwytkqYBmdiCWOYiOyHHDQL8DVvJuj4YiWOCIgW8DQuatmpmcz1P32p1IGvAiVA
U2/3Aus01CG0w10GKzae1bbkwaeJIm/L4emf0OgOIUnmpOYQaM86gGqVqS8psQ46
iApSOS2cNcTpFfmiRuzhXzjdhjNodcRDG566PFcXE1mmL3/OxOhQAqfWmEgUxJMi
OG7V8nqtLrGpyI324WwYFKaSxR3OS6SyoH6XryGEz1gTRVZ1qrdsC+CKwsGUQ/Vv
s8hdMZilwhl6OQQzgdNPNNQ8pzMzZtHdi2Ylc5v3D+WLGZzcBkTnjn4BH+GhNOAw
9EldovdURt80CL3x3SJfVdh+/VenlTvpNT/Orw2sjVXvb+p3DpjGFQO9AO+xWxPf
gkkLqW+TxL9ZFEr1uRWR4hDIc0QYza+rupNztLpOb3iEAxl/oQIHaen7LgmNo58C
rf4vd3k/cQ4XxLqc9HpspeFIY9M6VRMnaiFGYIMIl4pbPeXuhdcKEsDLdz26cPDh
/54sm6XCkKynQ0zfHVM+snBmQWm68m6RLlXFSAPlcd+yp+nUTqZA7EfqInsVK0oo
bLRG5Z+Cmp/bGdroe58vmeo+dkBAkTYwHC9bElc0jrv6GTPTFcg0Nl3UJ6SgiYFs
u2XApiLEoQrIrLaDYA02zM4d3oD16GD9j/ZrOef0C9n8rGeg+DEugsZEW/2y1n+9
fJ0O2zHDd2QFZJAAEsncQe8xABr+aCpmRQRqk7GtsS216oE/VSZbtqvJyBfT7D50
jnBdKa+TVYE+osy98+1hgJcfPX175posnlnq2jbrB58dqF8XDWTfKj5T2eOYQRCa
9uqa4aXl/GIRg1YuNiWs7FeuUDfrYUOZZ8W58CQ2lJ+Rl+Dhlzz1DbB8deIJUptj
OITfEMWi6tkRmDuAdAATh2M2iZ5rCrwXB5NLavIdXgww8k6bidB3W6xm8sfnoNbT
mCwgNp3plwo/mGrvIjiezGoyeKAJ+WuKF/2OqybDZEEtxI9dLawSnvKDIsBc+XAx
r/ALWv83KJpK8wYLcr0Nfri2mANuFhTwoOL1daacf5wpcmaYE5VGjZiFuX4IeJBn
QADYPogY+CeaHR/EdOs6eQCzj9+kia0AoqkoE8ArySqLiQQY4v0ztiIwEbkMue78
sPE2KQkNmclwnKQj9goO1uFn52R2nnMikNW5haBSfoqgu+MhzFr/+oENbRCFdYiy
+0co+vjfQ+Xnp4c9hCDJAM5K+4LFBRECjq9RNFoAHU6y8LPw+9/woMWIRV1PbHl2
n1A0Op9RtYgJsBTQt90Kjx/2jBybmtMBFCN+WI3xLqEWilcIbSsKFTtMxx0KFhc0
YsbocOq/fj/u01S4UeeBmIqdnh1gC4ScKMtxIJtUo8fIiSJxDvTWFkQsme3/1qtZ
beveEznTSNxnFwozLT0TVula+fDljAwBwK8yxFXIDRiYvKYTWmQkT8CGLENQSs57
6ehpGWq9u9pZ/p+Pxpp8DRKE/cQKy41zidQ7I6vBiJ+vdCBscmQbPhoVW+0t5cuU
79iqH+r8ElDWHjwlmBZtw+Z6YOuZdr/3tlRAs62YAnCYw4OUE75GEcYXAWKIqyn9
nCQkxSOsmIJ1HW9eefuoERrWqSS125qhwS2srr2kbeykXilbC46T2rpMquYVaTTl
yi+wXyz0UAQonR5Rb70MNrzlpX/3bRzkz016f5Me6jWGnvAUywlN8hd/D+PWzCbP
IAG9gwZbB/hzm1sG9DGJMaNYzDcOT7Ag03EkioezV5p/vAzIXz9EwvdV6CnHNR0i
9r9i1tc/kuo5qQE66aXKMcWcWzcxQJHBWXv+VHkn1HN/5mscbtNu0d9amulYGzsB
Dp2WjDsjX6ko5T7FKAobwQm0/E6dQfQwFBWMFKXrFHpZxZJUgbnSt9uWQ+A1VzMv
8z89JqCpGiwV0P0EOg7yc98pmt3YLB61hH59NWPT9rucI/aej1sUk6LrmsGKvJxP
k1jq3L1JAcCdFLXU/RG0SpXqIqti7vDPf+87xUhW2zgXls3v2qxzVNqub9bSoWL8
1SjiHi3MMzWGs06D4yzZQKPelxleH9O3AGrZ09u0xAPebsWG4FOl40LOEx2Syuyb
NT2US5ievceRXYGIocY5EJrOGF9st3s05QPH4QDquuLwC0l4pJrZfuxyQ5FDfSMO
ynBpyNifJZ8KNUYW2Up0hjDkqKK+QV5OPzWSCFdPDxIWxESQ35eNywkAxTPD85mN
m9js/ZxRdd5guXBZIFy1beTAlCdbrRdz3UN0Aki64eQ+pukHoe+mi8KytrFVSkSF
C4UpZwEVI+Wgu17ZEtQVRrEkseWCgsjx4uloDgCuxjWYWi0syz+gim7JFSQIYM13
9RIurYMwM/KbiOiyqvR8F3KUUwCUOpmDHu4a0E3ZwQQVuseLhRNOuAWIv5B9vau2
QVPsc22uYBCa59fvCKpW0yA9j0O50ghop54DL7UvBMWeZg1Vr5EpEZkbddhJgOfv
fk7kqs/bCrVW6zRPzzLDrM9Zu/1KZBwAbmMoF/zQQM8S0iR+xrzACnErfg4mqr0K
OjPYpnsKOOyB+MzTgnjxp3dJz+B36jsmqMbfGNSFFRDFBEfIWqkAxyQizTFhi8Pu
DO95uBqlxNIyD5o+zA80r36hcpQK2itezJQ4o0Lm223W0krDhnpH2F+zoKqk+Muq
A3LvW/hOobAbHF2tUgGkG1L4jroni9x9TUTAqDOL7RWjquA8uZfOuEDsbMz6vzh/
ukLi9yGaWKP+Ki3a4Hx7wK1OkiYSz642lMIFAwxLyHjpg3zJL0d7fsGpCeVcLBAB
0LRrkbrx2MdJAWeehTMzRehYSYmd/V4SyKxpKQk/VpRbstCoWh/e3C0T60FNhdyD
UNHdnkc1rqJpATFPKBNlyq/mm3EkEiznXru/Z1FJ4+uey9uNMr6PGF3Z6E8wDtqB
Hwf+zLyI2wVZvaw6OJe5CuQcWmWkzNKIxMI8to9i8rVXOif9hxLIe06Mvb9VbjGa
MCIBUZ0p2JUj4pYHLHU1AhjBM7AArU9j6+JAh5P5rmLw7NezNVZ1+kWU3wg6PCV2
JnHvJAh4WXNwMK83op81S8e/U0MZtmKiWQb45b3/0EMkhgr1/LtN9ooE9QzA69sf
zAkCXyb+5+Tawtjv7l1s8JDVXgcqholx+sfdXL1P/7slBPnVaQabbftjnGCPXTsa
nqSGMJsK0ClRq5rrMSsDn5OhrV55Gir6AAniF4inon+KDrT8vOan9RAqK9vvFlUh
vQPTSHdXTz6wbKmsBaEbZ+lwJwJcm/0zoPFOY2RcKytTe8xozT3R7n7Oe5Wl6yfS
VC1BhOVNKpSrKkqigo2ZzE4Y86gSF23CO5wUV9iNH9IJMQQjoVsRKYOV+ZD1UyvC
OvvCSCrpedQPpn7+yT3HAfrqgoNY5ahF/x/Og9Y0vvGkKGlBlTkclf7WFBOzT3OH
6Xvom3bx+/oYGiFDGyRxAS8A2iAIv62ZURssItKsSfYPYFO8sDXJSW9bmVwXnCrz
FfeBHjQP7Xbbd84XOkLTa8Cr3y8VTDuGk4Lw4cSaw49UgvDp/Ei3JIQ3UmCi+g0m
Cd4hbKvg++3FlgFPVtbgRvgxLTe4f5KQ0jNcg82xvahOrItCZR497ZuH5KWBSHqF
bChj15wMFu6hTtyZC8qL01T1cHhIEbpFfkphrJHsB7+yZqwhtJ/oUAILdMMHMpqk
2EkZvqr7VVhFLIOe3aNw6xEl/2NapD2bFXJpCcclxEE7uw9XmiRUo+hnQCaanZYK
aQfEBnCFpsFotxYCKYeNwoM2HLqhOWVAOHIkBdPVEouZpv129s1pHSz2qvYETOgM
iYqYAywQ2Vg5+jZGKazKJGMkE1rb0+ZoL4MDgjFEca69zR5Kc7cJpccHMuxlhVzn
/3gKNhrtAsUYRYYC/XyHSvpdFQ2zhaBQTjc3xAIwsNH/3FToF9qqBw+cJq+rtfhy
DZVnizKsvREe3ICts31fU66gSQdQrnJK0fgHj5zg7Zd1GAhNzsllFtC0Yj/2H6fu
x76aZlfkSFWQhFgfjl5QVH4CNAIYayfVfV4VAfrf2LkV1CgwFGaEBGuD0FwvTJiK
vXLZp93i3enTVm/9yj0nMflezYKSYxAXvi3TyHT0K3YRzS1hoLHnUbnXNH5lGhX/
krK4M/LcEVdad23k7z7E8pXJHEoZ6LcEO6yuUazB5ViZyGTOIn5d8CjW0B2cATMo
QKJsj3+jDGEDx4n+uaij18uk2FWdbW61sYEpp3k+KsBnjVZXqpCxvg+01jGGX0F+
ull7ipK/sWhs6plWLY8arA87zM4mRhqnCZFTyJaYb1fud58r+A0pMHiOSzk3EnNt
i3LwHN9j5Rs3TB9qnRiRLfyjm/9U42uxowCsPgY3Ek+ECuva7beLC+UqSIlbPit8
1h3rEq4YDXzl2OcMnpJSGC54tG6L3aSulOgZg2r7YSj3Ml/53m36dFk63MbtxTyb
Ciq3iU00BYJbqncnEOya94EDWQCWWuTdI53aCNv+ln4cgPcIOb1i7ixdN6zCHIy8
W78A6oP4JCsQkUNAW1N/BPfmi87iponCEqBuD6pm/azEwqZYQcDDksAUgXq1KUcf
khFxRP7XJK17cAbwc3bCGBP/79Lq/QE1CkeNomeiQ0nWPK1wdnthkylzha/0Ef5R
gSrj69hAITxMv+thhwr6Ho1yvekVqBgW2IPbIl4odyjy8zrEmNv/NM7I5LHgR750
SLlZstEgEuQmbFuTYrURFNeqKCYiRl7WhVPnvRYPKHvP0M6HaZ+cKvJ0TC40uoi2
uhTT0LSDhj4rJ8dP8006cwwTefXFcBhafG5JcB8kXHNRhX2r/9vMLceBHrRkjb7J
H9lPpBufQx3ncXGDkyUEH3hhUka9sNA5ht3DTUkNGBmpfLGNpt5yskOzn6Y+eqLZ
wRmWyyhwUepD4kYzkbY4NPYfDl+oT+DSvrbDOtR5w5hJYR7SqMZVHpJ0HkcharsS
/TBqKMIx/TZCb7kcyVKKikdqfwMbC2TT8kwNHimzp/ffHaHfeGxzurJs4QpJ4tFf
KiXm4QcBJvdxlsl9duHeTG24ztz9VOf4bZIaa37RuGvSNXgI5XUNeuyXuoQxKxTG
sL2/HBf2wUbbStIaJUK76YnKB3QSEFXCPS6vehMkUjXMoSYwczrkQ0jNuUZpVSRi
dzvKaoyi7ZiuC7fPse3A1hfU3O7yd7N6XxvhEI749M0wcQWd/LSFLiBbMShClZB5
iV1p29tDmTkhcH96TJV+4hskTNI3RafAAKYmbgUFSysCILNt2xyUbwhk2mEBV9Ww
2tfjvTDv+Npd4eiF0+8mbx1lxuQ+vxQs+2ag6g96L1P9Sy+90MoYtDg0cJJSs2Jp
SqZzrXFVMMxyVMKdDMe+0auZ4SC07gNVMUks00UG0g1htmMSiH6SYtX+kQ/KPsdJ
NZDk1NwZhmmRVP2I6rOpAS9qk+HlDd2mLPLa21UXyKjnvoJDM6E2Zm4iZgfbnNQM
O6YM/TuAns90GeqweS2PicxS+6CSMyX2vA/XYATEwlAYBoZ30UgEcjMOeIPov3DV
tENmbDFPozABglXlOEhq0357N4twsjbqZJKskdGoOLZCpGbE0IMR+PLErdM3DlRC
ftbf09cifrCBpOrd2LLOzPSyesqdsrAioxFj3vsd7neo5E8CCzlJkeWMCUZyapRD
qt9luCe0/FWaIsDwxnWpWNyxwrh88R2H8ZS57f8JhZSNJmzaVUpBQcHyUqLZBjcb
CgRMTvVeE6mwP3EgrLKRoOJC2AI5doYxSm/YkfN2HXTgnHn6vx/n5Qzx6JqUAK5l
2uP+iSA8bLsLummrKJr0DyAxDeWTlg9BCsIxyBV62JRjObWz5tO336cKq4xIMv8T
IFl21pgRdn2TRdprBqYvKm0q+xZ2uYyqbKBV/H6U5PShE01utFJgpxs9TyPi+SBH
9kZrhmYXUO9Nx5eFqig7Ly/paehiJRKf9El+57kAQQ9YCXFzV5V+hEZlR6vIUpbX
s4eq2OzePfEZ0gGJ1jeLw472ONwok5sNNWlSoRWqMybDNJg10kENkzCcwdCiWqDg
riDzAPG61WQS3eXWdeDnXEpbl5D51E1dOjQX2tqNo0OFdaYvtkIKoQgSjGucdxtK
f0hwQa3/gq+iIP+wXAGOPRvxeIKDaj9i8qq/grljwU4UsSNs0h1SZT68UMfV1hFZ
ttukwXBewdSoZspXxVa7At0Vrq9xoaCeN0ONht6qNvMMlU5LHzMJFONjtjBRkiiz
0IHavhoXYC8E2qjB+tf5CShLWrRFtRwUJTgCaxam9xGQ6WgxlCye8bJf49ey6OCX
JHXFmFHExpWjxYb+fnl+dID/VrdFk+pEbjBFnFTtddxULZjK+jKGot/CoGnWPDaX
+IsfR0FCsBSLiAKAl+8sc2aOh/+Q9cTItHyAc9q/KwLzwfygyo9kevx6lcSKtIMJ
j1dU9LOaNYZewoPRZMGzej63H1Rh8f+Y9RhYNRjaRaxgx/Zw2IduMP/XChhFPTm1
Yp6ob2oNas0vmEZqsjFDoK0zdCxSq+xloZGvi8aICO8ao5HA4QQtwW4LzJcF0YPY
h+rBXhvntjcTVZoWmth3LjT6Gm/CDVeMcuSx2NXsEaacWKt2GqKgrDuVe79aatFd
xMVde+3XQqWjPjFYv0GoeH0SGO9VGV/dkVOAqKPfEn77cL3C7GjYIkFckYcQWDcu
NB3bfAEtVB72fyPdQVu7eDkURxhOtacAIMXsBmhiHYRNX1g6JEkI9bSmBbWn3Z0q
T8rtug1a5hoQ2sGz3S9fgFZTxMUc+xiUVP9vQgZ7IBgKafsP3wIkEFxQfPGBwp7y
GzgwtN3gGt31FI83vxyEj6wkCDmKpyNIAfu+7XqjXOwntCb604Xxnh6DwNBv1njG
h0cJ7DIu7SlAgXOWfIdJhp+KE66TIktpBKOqz2JJMNL1ScE/5SXBGd3PD31EV0J2
R1DWR7/m6zweCbVhiVdtrl+iKfuITr637nmufpCTXs1yJgt2CK35MiaZnhBOH9Lj
Uy5lQU1K4kYBxtwo3UQGWnWV3uk3PKyI8ue9o1tJpAf8tbfdWPEzP3YX9Ds+ASRq
HibSajzmAlDHnpGwKB30d/mI+EbzN8a2co8vwaycuFil63qYHqnz2cRjAqLBvpPg
FP3qZdrI0nyVqxzzrU09k2CRJhkUuU5n4e5pOO33GyZT+tH0fRxy9vWlwidl59Eb
iy3/Avrmo//as/JNMiBa1UJ4PUD+2msakaC4LyG8NSV2MKaZp9MoIB8Gd816WDyh
3gt433+fW9Y/AumtrVz4Ft6K1s9n5c4nrGVy2PXFU4e9YgY4QwinKf4+vTWiPxRJ
1oNcW6NwRzE6IyPQRP3TId96dUD2xsoZK2UYnlDNLEJWgh/svsRlq6zJRA7GFcmJ
+hKdHTYaw8ZSzhKPGL3tB5pc6De/m317XToZEQHW0mlMCaetLKjLkF+qs26VLcsl
//tZJYEAKc8OkfWI0m1JV18LqwCGTtDNGn5CjLoX97B6p+ShmWeJNW6ZrjrhOtyg
HrfHjgP3XrASwumYGgxxh+tAdnyPFavmMrM7FFY3AFsV1RFXvnoGRVPxPLng9Qfo
MSboypiv4/svyWt1arFcz8rM8ID6o21txpYvH1Lom49y8OoFheOcI+5Je+5A6zrM
OhCCnkELGQdVjjOB4jd5LN6hB9LfSZUOooQilo78+eLekYnFsTJXb7HOjr4jCf7B
b8tnuT6jHD5jM+NkmzbPOgVe0657EbSUoyNhT223M9noV09E02+1pONF+Nz570I2
G25908qCxntYlSQUl6tnQulh0AqHigKebgW5hdVWlVd1UxSwcGFtQhuaMG74Njw7
e4/uYNcupUO1ysWS1A4BCquOaDk22ki5ebGaKuqOOKMCPPBB3gV/LuJxzBGYVYrn
b31DLX3EFCQr1hCaP2TB1UJAFN5H/5+HgPdPqlh0iFvAPODo+nA/cqmJaAVi1uSC
SEFB81hzheIjmUSuq3w8IaaejmpjL2v7h05Dwqeaa0ZxqoGcyOWLJIft9ssVLv4/
jYZ53rFFjXQ678DuT6xHKDMi8pYfXpWSKjraaeG/R5Pbu8EHEHgMLvaIdOwxZPss
bwBs4Khxg0KYHeZPct+EHMeyAzE8Oj0BKFRfD7dpHhvsmsKyoDscikBPpjYHHWpu
6c9IPvqVPlvrjUOp6pXhGSRWczyhVl9S2gUu+JZYAaW456KPJPVu+Tb436efra/9
U2LIa7cN6lGUHWpilGX0Nk68M8jh1OVwcnSERZUMluk31z9yk9a3FdFEQ5ztB0hC
SYnO0ZfAYPyp3reE/NFGS4mqvEZXq/urZNN7j1jH4hcyrwNycm9PBARp4Uq9Vuzn
mtI2KcvBkGCZM9/3k0FL+2lFLgGg5154+9QoR3WgUFbGRXz9+Z3eNECSizvFfqns
wONAm69be78rZjgePm1GhMZdqfPNUeY+J2ZWZdQHJqobojqEeZTO6XQqKBTjjye8
5jrLo39y8i3T6v/I4VDmxFZfS9LlqEjw6scsz8U5ZKRZU1KpUFGKG52YVaNufUqt
cieuL+dUWYstSL9xUPKXE2PqXwANqb53ARYrmGryZBc4iK29U9Lk5CKX7bHFYr1D
1XyzuobsXutsQE5fMqcn3fR+wXgnS2F5/bltex+Py43GQUTdMb3eqXafdfXmT2bE
KOkfe6byL3lKPB5rwSXi4tHerY9uWENmlzdEQQwujOvSdxRNJu4CcnREzkN5DFud
4Ps4U626QwAi3ZRsW9EZI64lOhZIr4KImB/U4/cUObm4MEETIcUO4hcIcGhJDjFQ
0MPPeN4n33qJ29RUVHrVkWY8jvNlHvxklR+RffKdMAKGWFEvzG1quYf/q9HWd7of
ZkwrpWPwL5DcP2A6PSTRKxnfo6rSbSZHelkyi6O1aIycNZ3Ohy5SIZHFBrqbPLuF
GGLeEEskiXhfmjFxIp2D8JZ1mXhYrn6W2qYTMnAJHM/UJEqT5l/5v7kuo53A3ssC
9xiUjZjV4F5aTbfF1J+2AJJbtX8MgB6uwVuANZbK0CbLbSjRbE+e/WNaLRXyVEda
Z050c6TfFrdQQ61jcrJ41aYbGoaYOW9nO1ynmxQL+mZcS71sCLVLjtAL3k6XjgiE
6qwFngPQ7HTZBx9WdKW/6pX3yUYeaxzM08Aj6jdo+HPex1grIrUhQ4+fvT+R9d6h
q5OThArP4xZE5DJhOPyjYo8fwfZ+4uWcZ2IEjInnHLs4jdcq7uux/lVBw/eGm/uv
BaIhGILf6UP3EXfo+r5l6Vfaf3oxb62zKXHMpy79XUOLkA+MKOy+7pZFVioHLlfB
IfVtfbTneSgGCtP6TAumBEusJqGTJo/0uqqj+Sj5w21+ChZyF3DBfGiIfInEzqMv
lwYg8MwWpuwDdHZ/xkINN9s5cTTYUE5YAj0zZbMRx7CLBLcdqs+ZI0+/MnpBpgKN
JtCzwnVjgwKj+sNvSyhK9k6zSf45UC0r3DvRxtY8n5h3qZM6zz2nzJI6m/jXLA7Q
CVnzK+SXGgwLQoTtvqgzkSTgwESW2Yj2bYVtjyVBAdaxMurxxXyhAHNa0l/nnQBx
W1xwzC4BsdQyfleNVgJ7r3kOHLHt0gJdK/lIkygK56aazpzcVz0awk1YuYRloqaQ
2r3DdGRJxXD9H1WD1jRbLgYpd+n/kH5es+0mzwpectq5+TyqoeEtKSaR4DzTDt49
IABqeACDGcDDlmur/Ig3BsfqaGkN6chalkTRrYZ8ATBwIBcgt56yrXbZBCqHH1DF
bS056W1kHyA5DOs7NIHwBktpzjQ1dsVB98QjZoS05YTkeWStDoPPIuJnYxzDdEg+
fvuriLoENXIzoRep6gYEz3t2L9Kk9jjblIso+C8Z1yK1j4N2GcFSGVyNUlRtM6bP
a4N1RZQyUjNf6IdQlsU9Szbze1cJ+R44d89KvoRU50LQOyl6/7ZmxEmvQqFZn9hz
V213dXbgnlYs+qffhxstbFtQukqYEV/hoZQgOh/s4m+3t7FX/CUz2APGffjWaICk
sLVeurF+dbdyvz1o5CEBhKcC5sBmYaBdcVaJ9gpP+CSyx9aojsts+1YsnoCWtqNI
g9KMqlNRWKOwUcfhDhVuNe3PaCni5Lb+IUg3+cwLKgP92s2IsLt7YGwFkKPU3kaR
4LmnFLERVKipZKmwZE3SSHu+ZGc5UZKP/gm1mJWbtXD6z9+ZBfF7m2NaiwgULPTe
fxSchFZDiHDV2N1skgKxA8fVIVAOw0D2NSUKj7YaZqh1lVBSyLXOac/gEuHgN1e3
abt7BG5mFxm8R8H8d7Umz06bx+2TgLw/xiD32QifmVd+z13M6/w2kAHhLv2UC8VM
nZo/7SQHUpAD5GcRVXyNnkg9+A74jvoUNQKN4hPeBdAlMG+xi0iE0ysNAB3vXCQC
NE4J0j39TYWUQjNLxKjkvLiBEj8NgHd/AHKCVXrS7zUdmnuif5xvSO8FkCz507P+
fVCf6lVKYOeq1US+u4z0Zpbry/XShm/QH48u5I8CNYYcuuvIDGgZ78XAkkKXQQSl
XtfSMcwL/rY5T2PqMuwgn/Dy5u0YbuMysBqa0d6hbJWwtFE+n3d+0kFdV3xx7HtP
st9KE6FVALBxcri04FkMuM4O3affQhY2E40beUxbdaQe9aOiqfFMbppTQ+a8gKSU
kadKbCft3LhKjXbvGj0BQ92yGgC5jKP500EU1RWBjR1eL46jWNhIiCv6zEfSUgFV
qthts7gwWox72JCsd5j3Zx9I4s6wIL/8dESvDtd7H83uhuhiWjLER+4WZ2rg7U7x
WdIqg99yRtyBV2HxIyrhLY7SEVMt2KgLFSIeXpNiEtcuGTzsZZHZTcgNDdgBPR6o
EVUSI9/zHi8rGATe6PAmZkJ9By60SBCiN4rZWRMbjGsjjln4Ydn3UFZaZOvVc6ot
+q/NsRCEktiju81vXFoMSImmo+V/7MQ1Ko8UuNe45/7X8eTg7UjXNCrgqWFhC9+N
wv3YAo5YHEtSVbYCifMBhXfTUx0p0dBI335V1ma2rjgU1/y8a9dJrVuFf2DZ7iBS
oU0aP9n7rLPXG3aciyTL2RjyYL6zwXWXWX68GgyT0OJjaNlXnoidunZHtdQtqN6Z
HB9+V+f2NNJaPK3HyLcb5TIdiTdGauKTVib+jJCUbH4kW4aOADPUN9hvrzfi5zsz
RjARmiKzQBRPt/ic6fx7ur2/ETwIwD8dVfucamr+IZnSHf1FxfGV+gq4q244nWKC
9kD5o97QdVyn1DI7G1CC4zdgKuUCV7HhYQe7CJKBNEK694HeZEa+JWj9AW3z+k4A
s4S5NIas5HFMRgORiAAJrMPDsdwhXIWVIIBKUxOq+XkTtw1YFBHTnj+AcFXRn0kN
EuuywS8PSjdwdUzIe0Wh3Uv3fCeLhMtv1GZaiha2bqys4AW8byYpX1pNKKRACUBa
m32yNzUEBgRH8f+lVc70jRR2TyY/TI5pcnDjKM1ml1zdWsLeuxkWHCEMRZ1lKr6y
GKWhbYqjlLgS0YW+zrJf3azIGC/Hgtto3e/QIdOwSscRIilX0qQ1+hEgMJxcAzKO
Oc/gOx/lqpiPAZuIdwz3Kk4CB0rzh4OPlfS6PmDErGYpCA90QJ0EpyXNjdgVT3q0
VMpkvhxuMIhEoC/sGAQIRSk7AVoG1Q+1pdOgG1HXbA6IdEONEvxyiYkdfsJXjQOa
zEF7a+omEaWm1ak6sElj+5UAr6gZu/exJ/QkULYXo6Q1oQm6NXjYoRo3d0CH2/bo
8dL9QHRiR0DJ6hIXAAYubHufjENndwTXkWKG+7DyrHAjXtH1pS5Oa40CBEOShW9J
XEWxyfWSmL7VN2FhQg+FOJpAB9tsHA6nmkqqNkzWcMa4JsEjZHhw9E4d832+Kbdn
n87e89Kt17c7BP6vkwc4ecVCclifmSzB8GAgnpnCoIhQZh1jcP5IyH1ZSrysO5BL
71KOZqIJiOmmMQgpK91SyRTNFt9qyensV02kmEsJDdkyR6yvzv7foJs+qcilOHIz
nYYvdqJfTRA3Wtmt4ODVPUosrF1A/KETDfQnL4sabaeRbFr6pmMtvOWYhEgCSNTQ
5xtoCPPd///EdIUqtYBCJsNYzKxIDomFTrLn0SlZGlDEgpZDfGrY/EeVnbXtWCHe
7TkQeu2tuaiHEXK4RJTRD8b9vsId3oOvXKVNwxRUPN+5WyQI2vNQ14PPcu/vVl4Y
xboHo3ze2bXtwnIDcmUva+b8v4J/ZYQXcijjM2QlvbKDcAXkn9kSxO3XX5oYUv9e
Qe1RWdBGKpEs9R5m54N8VrruS7PrFp944fgNMdykv/jdbKqjtKkW8vr6h+v60D7P
yEt9yrIeGLc0eO703C9hS5RVBIbAVShpdOsraaibfwtOlTUSVmAtBR9VFrF2BpeG
rEwX9GMiK+7vbuCq2hLLQDlSu+Ws9E17z+pwDX8ZSCTgi20nVtwVzrO6sFAMsN7J
JlQcnY4sgglJf6MrCHIkoG+X9mn+OJD6ubyYKYdx0e4gEaaEkf+pxMMN6bkMvQ0m
nH4mJn8jS3hh6+EfeLpjAfDPLTO28+gnAXfFWSDTTxaWNr65wX+u1ekyhxzUQ+Jq
zKfxklEMmd3LI2koYCYvbDCaaw5kuh+OdA/XZSnXkXfQe4q2ZI0aJgu/hIzETjgP
0toZWMy4NZI3Tx7HPSqTE2aE0O0b3F2hVVGPgHt6hNXl7xBhVXLwETXKP0+XJXJb
3r9rMEGT0biBjXY/JBMDskYDA9ufsqGeI0xM4QRajmUrg/gpBEOYprbvY/oYeM8D
+t5RbFixmUZPP8maVBR30SyfTmfoDSFYYcRTSqK7lDVtlVHxTcovArKTjuL6IkGu
UezJKunVqOw81N9K0mu/hj+qcgiRMc2ucWpxTRYqcCBFqeUYAijjYGwxqjMP5d4W
DgvtSn8wYtbCT1urNr/1JJAdC2H91+uCZ2SSr7rDYrAO5CRvcCVvxhVr0wBzShsi
6kZ1xiLHc1UoHLf1oVtaP9iL/O1VDt2OjIgfPp1AVK/325USnQAZFe5Mn+KrfjE8
FByOiFVh9K67T2DUlO8IrTVEsmPpYfcaOsdsudulH8v6wAS+5nCkgj/HWQw49mRo
UElUJunWtQil2lKXFxNUdK8qUydWe1Roo7f/fgmX8lstPQkeh1yUj+m0A7fWCAwj
lcRy8NeszmVZ/Ls5BpBDsTsrM2/zmVbMpKzJL1oIWWtOiHQiwEqdmxSPWsfBub6F
8/P7AOBizd6wZN2s0AAcuqixgf6CWwtTpWBrWfWAEzQBp7sV1NbZERi1ydtdv+hx
9tMUXmMtxaFOyqCdUfS+UbahU+AJtKymulxkBytAnAzcIzsUax2VW04rrRbag4vb
E7hA1s3lVpASCPqLmwJO7uBtWwdkOVU7nWIKE+hWvSz5XMewA7zndfJPGh+DXSYP
1Y+eMS7sEfYDjzOumoPiEPFFAa2R0rVf64hkGP+vhjJ7ZK2e5brzJhSYAj1BDopQ
lkb2v756LrLWS66qFA35pWc8t5L3dXJhyEcTHMNoKFMzpq0X8jbg/xFJ3psDAR12
lkYVPI2ZRoVQXDm1ZCftMBmhuR+RlD6udN+Z2Vovd7uK8pcGH/pT+FlLsoMoU//V
v6QgJQR64P3tOF2P9UEkCvn3GTy7/3J8P3mRuSYrrzE7PMrZ4ClTM2c5uUUFqa+A
2tHaZE1Bk4EB2cvam2OAX2rT06RF0SmSqZftIdY0Y9V+ggnmwMhIRHW8mSR3ZLwW
sPBX+HDz/GkUq7tBHcpYSAIkJor4+cvpbr4NgMRIALALqDuNOYsGF4vy5O8EbNGq
dLX+BqZ5hoGlwsOjjkf5XpCQt6rKtxaPb+BsNV9fQxzNOrmXr+KCtadQWQUAofI1
WbwmzKX0irxVVu3xl2fStkhZ7YA/7gxVPhY0QEQS0RaFxTSSnlQu5HRC0EiiANWQ
jQP5l/MEmhI5dkGn6kl5rHMYdoIAra28Y8sNq2080tSwhAwoIZH/uvo4pTVMpGQi
z0EYbMHoQQNQg+yYyJLpp5W8D8TO5lEZcW9oEvtTLyfx/FZKH6zfD3Qu6NMGRT9G
SO4olhZGAMkeFdc/7noe2fgcg9pZzkhqEKdFmyW0qXkAghHS9Yv6TqHXnC2jrv0B
MO9qemXJM7TDRX/USPdm6yQ+CbGnKz2Cdt8gFXrP4Y2IFt8/PymrpaFjoVwHhujk
vsChzEIJAK5M6dFxmWIXQARb+oJ46+VHuatTPIU+EtOCprwJQBwsGbkMis74NO2F
Lu6b6kY4R9VYLtkQFr5R9A8vwTh136EzgUjO6wfs2oFpKD8bd8fdYLypeo9YqFGi
qR1KFCZKFbivaqUb97yzL48+RhHUgoo70zBcPdxDsZa0qXx/qaDBPu48w+1Nvayd
cbNNjtoLH30taiaTRpwPSlPZgw5u/JEBIUyIs7U7hEFQaml7TLK2aRllF/E9F573
PGUA6ZIAP2ZM9Uxebc9IKs3C2bkenCPOpBWdhgNktf4q0QaLx7tkwErdhxuoQrtS
AV3u6wDPHkgZzVfcyWy5DUp3MLMsUXxO0JI97lCb7XC2IzIbWeqVR1hKEKRn+g20
cCrhK1l5KZ044kCx3rujm+On0mkU0Rqm3VquStioNiebGge+gIP/mwAjdQNkt5is
UWkqlNaqzijQ0bipelfi4sVVijzU/ooYAIClsMRwkTOnM7nDzJ5ZmZZamsrWPSAP
PUkcwB56HvoIqfsVAW5pQdbaw1TQ7aOq3E4trDzLSRy4gNLOsYH/lN3wskiH48qm
Yfk/ePFheJXCCva8hxsn4HJkfSOTLzY24bP4Grzl+BKvW59ZbN0kyffogGG/JzDI
+8RrQ5m3SfKpptCtrbqyBnBcXB4upB4FzHjN2lPhrHW30N5mibZ+4drfO1Pgdh64
iObGSgvRjsLMR/GbHgoF4J0PrP+VpBEE1XbxNkXMmq7s+NQs6K04G61mTNPYuXhW
+2CTsxeJ/9okA/670U3UgdJBGp4wGUXIYedFA8jvMrb5WVBjtb0GnjK7Ex5dxIwh
biYSBo/QQgwT4hzxu3r/pGCe+c5TcXs6J+QLTcdovVwEAgrgXiu/Jp3F2OY/BuhQ
sLSCelyvJa6h3cYELvxyJnL4f8olFT7Z8rX2nXO/b5kRwtmWBZ5yMa1EZrRoIPif
y0N5ZVcVvlcZR48+MaCi/mxY+UIk9wUA9/yNElRVBs04lm4r0SaheuZ+1iSRKjkx
s3vOMmOeLz0q1Dr0WhrnV1nSyCFA2fNzD4Pr9P9n3iTTqskeH28X4fMLEz+wsSq/
qt0nLNB4VwYxEJjmAzbUHv5PRlI8hoENeWsT6kzFPsOsUs1vDGLqO89FsuAlQLt/
5kOfrTNWTAjYSKORIHVidfPNpsn461SD2WDIIMUUZyaqj1L6cX4lpUEg2O1mElly
JEHD5nLB55dkcLag9tHnLGsAg7W3kQHjASD1CG7JJssUu31khGVEQqPAGYv/zvfD
sYdTYbbGOJDTUhwfOaVKaoVzrE10LypPF7o1ORnX2dD6gz/6J2wu0jvWRkEa4FGc
ZKwOoB6VyHMlNTMKIvdCbnIHsiOprR6dFGDDSLFL6j2KMUNjnnhauA+a0spcX3M+
v7aObg04o79RgAlURXu8R2KIU3kX5/nlwK4KhRrFvLO6fAwQ1boWg9pKoeM+RcLe
pAF+PWFcrYRuJWB9DjtZBHkyc7oBYl6NUJMMt2wfcLpV2WW9lvymnw2d3/r19q0w
YrXNh1ez58AdFB52QUhSviAY1qfUb17ZfJDiK4WVBgD5DFlXr3gpvlHmNCBJulP5
FUG178vkL6Wj+O5v6BUSl0GMRvgoSwwCbcRVcnDPNZitRtK5qExNezycTR8NfU5E
/ZQj1WAccOq/MsqORosczr4AGzdhQD/4vNiRmIVsCNNZyrUBX2sGUk3PJluQCW6+
8tzTYIXwTCnIcjm8Oa2LBoeEO2VzJbIRtapT5arxBy4jS7Z0g8gkOuF63r1BSnmd
MW2xX4AnExFskYnpInrL4CubaARNy6hUiSGsm1Q1ISVv8ZL/xKyMmozXephvdymj
HjMPxqejYl/hBTJmP8WM+ett26M7V4k1nhOnHW8HH5DjlvzpqMyVJD5d8Q8TpMhl
B95CTmRfZRONW/sFp7x4G2fRWHyvJRTwCw9JctfQ/oGorFtEBVga4tphNqKsJlaK
NjAhtzBvJIqE65buWyEKSO23T3/rCV1KdcxFSht4IQKoXZrc1wsWL2BAe/eonXHB
IVg6zr1ocDpGS/vWaEP17v7taPjEdquXY6YQ8Y/1Gdr0QPe8uopUdO+PJOEQs7E+
/YQOUnPWnSe6TU1TkWYf636bNAcjUks0r48lBdnJCANhvEOQuiRY5xbDcA5bJu1Y
duage0B8pbSJlyQMTfjw2L/wlvlaStfFfVgbQCebGHpVUt+3RHatgZfsdr2RsR0q
zmbS7RoG32UR1IYBR5uEb4sJkC7MGuVxunUOiJXvUMXtDR6oz6vz9/UWdGxA2yz2
lJoZ47nQdrTG8JWR1aty5uBsfO9v85YpM7gagxB/DTBaoTvnSxQLv0blaaT/x8oC
fXSnz91HyJhoFrR462BcON5XFW+vsxw2hfv+Av7d4GeRInNB3SOkCpe5qeTTny2F
eXA7iZtyIN2B3gn5IEjvhD/IqjvOuZwbczmzhENIHXMZDsZXPCaXT+YMBh68QHjb
axTSkRGCIpytWZak0yUbE87SCjWKSuQVmd9n5ogp3waXg4qUiJu0BBSpJiKLPK0A
PvHbFLmDR7lzvDkxCw2E3MyMcoAUVL7VL/gHwso/I7YFNd9+y8zeVFsENFjkbHLp
O45MdcdzAI7F1tf3b6VLWf4lPyAa0+/bFbBvSkGVaH03Jq04wCQvrOzxwYJk02QW
tA7BuTiBslI42BVWOsHnFtUNByLIl7+kPCIIZ33zwzX5EAf747dVLkWeLRL6Y1kS
lnv9ohJtetGzd8fMvtKaasdKsfeyCkBSOsj1r8dOG5CY8/J+Jp6+HSxNEAbbLbCj
uEtFa7Wfp/sKEh7sHetmOc1krnvcszgggvwK1xa1OHzspMr8Dmabde8ULGKPOx7g
Sza5a2/QRuYohiV0SxZ5LCEcHtix11L0SN8whpyxw3ylIVo+o4Jx5xT/9+i1rFee
5WIp0rmOkR2t0jrPtZG0hAziBrJbpqFBLXAyc42Z+3yAFpSkr6FZQSLHn2CwrCiH
mfU+fKP/GiKJgFRL46lX1fGSkSnsFoGhm2qChJC0eeh62lRDphMmuWk5nCzWcNrf
Z8soeTEMhg29d3F3GlFmiegfO0OXxigQb2BDrHigcD0PF+fTHnLyAsVXmXh5tG9u
xJl45zl09B9rXv/5UiqcaNohtWQgUJrLpXEw1hzfZV7ykcXIviz3grc816vQ+pb5
L1eDf1+iQqotmSQdDKAhG8/5C3lGTh46zecUehUH1ZeCAzAr0gN3hRt12LFfglDB
wkstgw0Yw6hZIo26pUS3dAJI0edfP2uCHYxDOczodyJRsm8xZKZEglXKSoAHZ4rH
PwDqIQks7kAqXeFt02Id3CouxFmX2K1XveXgct1mJ74/mGP2IX7d5Zb/QrcypMx3
su6wzaQ+QnnUz4QqE+HYeCP701PNFWLT58Wpo2aK6YhY3fQ4IMGNafsRrF5ZZhs/
ku8u+BgEkEwSldU9v1JaKVJb1OawOAPqENVybp+XDuE5KJ8csOKd62xr0RFwrWDQ
Zoo4aEFfsr5+CopAUCsq1tVAH+7BQwK7vkHK0t7pGV2PGjl3kQLEgaqQFtWbOp+Y
6uxJfY/8HC66QnII2PQS7fVRu/GvjjLzt5XpRUbqN1RsWdhO76WedxZLMmqn5O1r
cYj+s6wA3Jfe3jrY+N9li+rvXtSppUQFGWn9ZNXsw8xEIYVuvm6brnScvZiZGMgK
p0bXfevOd3Xzh5F7i7ivVojNU7EFFe2O2aRrQ0VxwixPMP2rVrV6/geIMwG/2hNw
F72rD/utOQRvHLbI0HDpyk/u+ixAi8s4yyLvojU8BDYEda/x8GcoG+1oTQWjizVq
Og2VhNahN2qm8UP5auwt8baXTXK7mzAmgGIALzSqmDU6+smL2FQbmH+//OuBk3uo
9JOQNsP/erog1sVKSjgiT0AQZMbnGb/INV0/1nec0pB2zfbvaqAU1bq102P2id79
x1qQu3ahoHU1bbLh6Bs8T4YCXfF8HRTWH26lTyNPP7ZPZoL40b2QaPhdVq4DOFAZ
sdLoT26tLb5pob6guTOP2VndVS1M8zFoeFqFZJYWbBS5rrpDFwHFW2iahGSW1c76
nwBK6dX0+Dw2u/ftMFG2puRbB5lpv8D2KPldis+zaZUk5okhlSpdBgzyRpgqhaBI
XxbpbJll/qs58xXs6yn23bMgNP9Jir/tbhAbSMztBcLPYnRp31hP+LvpPyhyTD2r
4N4KcTcnbTZpfwJJ8kUSb7ImjgRc8lrFN9yDj7PuuTtzBOhIqh1L8dYm1++Pvi82
TEjWnboICAMfDixTmSEt9vlIKjw4CGxlKVjCu6MwmlGC4bUSILeF/fU1uDKGxp3y
G+j0LECp6Mk8BlnwDeupsOkbH7rieDQ3uSoa1hwwagjdrhxhMMfEtzuXaUPINgWv
u4tXofGfIhx41iZRTSAiyRnRf3YFw69zbWaKg3UgGETeG9S1XuRp2ETXgiBa6Dcl
0ObWqmrhkY30v/ln2K4TjWKrEJeKQ8nBeLVMClJ3ogMZmJm1/i9oIsNE25eo8TP7
te4PQ+SneA7FBOaci0roDFdaYvmyvQ2PB1BVGgonHYmYQSAFN36gqEWOKn+IgC57
btdtpBp9yLwGJ5vj5osd0DAW7W4hW7d/p3UTMnT6IEqzdGUim1jXslDxRiEEwStz
HOCxmnven7vHeTRLYJSmc6Nb0m5XB/W7+yXBDwD1n9xh+IJIxtNOXoeMzznKJDqg
S5TCw52e8dPImTT4yAKXShHW4mbRrFwrGhkiWUUMZUwOguewKl+cynzi6CD1An9e
p9GQgr5l9YFVqxZFRjQlECb/KYm5qxCMDMo9WEVHUXDfrr4pLsR+L7QevhNFLzNY
AsxE8w/5wZXsNrY7R5SgI6gOA+5riqe/Uu4jB8vSYG9mFAECfGLHCd2pb7rbUi7k
udDmWJeyD/FFHuJ6ugAKuEhJrp8j8TnlaazrQjHt3I8J1IuKzqB43YMnkO7Tomfd
7PC/tbv7zlQjxeaCT9W33f8nKubYAyBIArPv33uedYwUUYzeYQ/10LIktoli76F+
b/4IILcBkRFSgBJ57J6hXzj6fZ8ooUqEVt4Ac73qC7U2astFYe2PFasrbDjEej9v
17L2t9KFW5RSTm4KTMXNBtLI2RUmpwpl9W31dADmbG8KBlTnhTWhJXVAPr9ix9Y6
FtyZGC11wwH6wAwo8eemLsPl3qOWRjESVsN8mk502I3PSwtu5iiOS6GbcV71/+vZ
XZ156Kbv9M98xfHsaQ+CXI8NVc5Oh6tDuJoLVYDh2aT/6qgj3EbYNTvGmtDuY/h/
do9HQRXiKEuU5glAYL0q/CZEPDGW6CSkJCzqyJrRNd59HAZVu8qJPf3AcTV1UqfW
YudI71lSN8XDramYlFYL9xgCVl8SzCZjE0itRVRxGopsxx7j2tlc7z37ZCr2lgVZ
Rrml8BzQ5dHs2qiSCMzATiYlFJbb++ZvTHlLzS/+5wCFvmwfYodeAo0OsNW3K2Tj
H+/evUCshtLAfeqmjRFgyk/J+JG4SZ6OSDsT1TEVGPWBHsH8Voyh+ZGOdy115ypB
NCrSSUhUA5Zlqoswj3koSNDvenJr9Jddq2MyGzdhBpjlbj2o0snibkAGXNlf8tYt
OX2rtNdtckk/FLrfQw+OuR8JSBobUpRWzMxEkRmS1tDCpZMA0qEqjIdfSj8QaLfG
yVVPLY8ist9xYZjzAWX+7FRE5Dfx3Q75inY3ekGgaVqL7koIGLLEq2EOs7n2Nmw7
HblqK+8ZfMbgY1T/1NB67PHzkumGNL5WbBIse0j7jOseZRzoSEDsA4q2CCQUwaRY
SaBGlB0INMN5sjBweYAOcmYOKi+YU/8PADhBq10pT4f5kejXypOUuyG1g/lAP5Ut
fl7o2vVCvcggUq08Q5qamf/pRmjNUYETPclVOviY9/ygxEoRozsP3iEyUxe7QHe5
IXT9Ug1bSjvSzrBGimLfJP9MtP7HEVvC/RuV0pZBpft7ykC9h9JQbbLgs6bp3as6
L8xmCXixuOM32LRoST4HQU55mOX9kiUMeq0rY0jeLTnIXmd6VLHhwkgwaG0Jwcfh
0aqzfqAoqR2CDbafXgr/Xo4tY/DfCkA9fZP837QirrGRYLTyokDJVD7I7JZl0ClB
ot4iMd2EuidJex9uydxsDqTHnzI95bt/UdamjXsw+34CA4z39vi5ufELg+4o8C9f
3qSur356QUrTvTSSxEfLRbJ15pR9epESeztHeAVSJ+L2ji4cJRbQrh3U633zWRqV
aUkbhJ22WCx4VvDgAYLQLeimv5hWBmzWhfJl7s8oC3ZWekf7Jyu3470CvNVPsgwt
t76AsScAfmydJFkO03Y3ZtRo2Sr2BtJmG3cH1M77Nm1n9BRcp9ibOoIR/xPCx1Xg
m6SRl0v22LE8XdGqnMv45GJmT+vKrbnhrorgU0HfsiWw64I2LaXTDBWYhRCW9CBD
oBf5pPJsazmbCP38Bzj115sZnEhmClmIJv6Ro4rmHgnAY/+VvJQQMA7VjHkBeUtq
blcYWjyAcHW5FdFQTI3qLypAHbylEKt057fbGUgF/XB4NtEQZJPHpQgxxAaIDrvB
hN1ZNa3eWZxVsn91c6HXWVLDQ4mWTOfeluMmJzGVsTubT2Uvh89kpwO39HhqfiiE
F9OYdz/hf9DP+gwGYAwWHlSQ5GJkEppBj8xZOErxAA8z3gn4GPEoxvEUwICJozlj
pLn6MKgu5xz3Fl+gQX9lOzc9oU/+A0rFK6CUF5GhdJdg7PbCAVJI5a5TqT5utYmF
D3x/k3UN9VSJ346Ie+BBcSmciOQlY1VZHgg4c+1AIuCDocSw5Bqp97G+BA5ijOk4
nbZjRTs7HpUHUbxZjhrnqdJSkJZUfnYzh4OjfsRqcGJEQHTfq3o6hu3caTgQptpT
yAKUlyvMKkBxaG9CjfJeBbOXTOqLP/3heZzBZgqcGvyLh81zUESq8CP0TDfAvEJ7
MjL2HEalHd470hCLGYZV3Y0qH+GQ4VKcWr0GErya7ZvoREfrvFHc4YOQ2/H/vInW
KQUES4w7lfqaxxx09C4q3HEHv8H9w6bg2ZggCWLbGrkJp6d4nL11BHzmtnUVCsGw
a4FvryWMYQlOZHexVxzPd0+Ib2M8gQslR+P4WJjbd0KLHDy/H27HrSialQluaase
Vh8/YIrwZXFndAPzzuzExe8EkiuyqnZ3E/1sErkD6w3agd9UwywNr67IifsnTx5K
1E5OZ8cQ3Z6AvfCpvk1Ag8tCdGrsqMDWnvuZRM7fX0mk/7E6d2OfX9/obKcpXo6b
Ydc05dpb+GL94g2UJHK7P02NtXcBDzOcbNan49aAyckHHnzQLhOiU9yAjwT8qLqW
XLbQQQuWPqrQk5GHPZejsNLRw/7KF9Pwq4IniOUJHXib7sp0qClStkPk6OxQqE+M
ud8mmpS3ejexwDsHAWEcZ0oLaekC6Ukvp3TguRhaBVRxAejqVQesBlAVLGHVitSz
M3+OLE7gU0/bvJnni+JUPJ+qa8cIRe3gUcgvt0vky77JYCaBGUCtsNq7aJE+n9JT
OCIzXdCQ4jCzSCnHIq11ag+U0lOSxO0Ew61GuSUG/MKQYvOfCRFMVs/53jQ7AJ3D
H7fxQWP3Am2HrzEBaYZWaLRjot2fNQeQIgmk5RxkF+9e0PkNV5FbXU8HuOuLV4Uq
bU9iGMiC5ZLyMRE3vqikVDKtftvEA4RTD7VN1BIUjbZTxUHnBHQA5kT/vKAnN3vb
IrDRb+xmpeXBzMfbc5qnlqvvxxaPseyPyOeUAsyWO/0mlMJgYl553WewdKj+FST+
CBkagFbKedoDtHFid7EfqThzAdonW5Qwqv32GPDKhVz0hHhGC6jZMU19TcCYwPhR
Dv3XzLTjm4D/Lhl9RXzZZe0+HovBmkNLLdXIjd0hKyU8DhXalD0FM7064uYqnKUn
neyBcgBDTbLYCWEoA7RqOCwcGBKWQ8vwWIBwK2qJDb6ea/FwZtcMzzIrLlqqmdB8
B5Fbt3/2gsfkqiEBN8QBQy61v7n9NFSBCRA4Oq5Wtv8VvXXe1pjoz1GSPDRcA8Qu
R6wJo87XDWKTGdDYjEbl65CUSabKZBeSZoQfDV8/DPozexVxErf7+7tmXipInAnM
IQMfWm/BFWYk+KNLbzFNQqsCRl2uFReqBDCXQJrL7a5+4NywzKwexXqDeGcFTdzv
aAhTiQCsLWvq0nwTI2BsrikHz2YeapOuHzg1hLrZFkJX8G+qzwTKC2G4wlImIefG
665TyymzFwv/2LtbUqReDFvW6Kj7IDpCsHTWhtGrCfmZtqVki1wlXy2SZje7Zjec
OdkPPFCzHS0AVmCmWBZ7Iu8vqbZ0CAPNH+HLLVvwVNIB8gPQaMjiX8Owk5Xz6c+Z
ID/4GCsk1+lfp218QRjJcKmczJwuwdjUq0mvKJthvxJp3TdXD3AzN6HCWpem++xa
uyf/mA5IPZs9DQ9kFIcWW6I1/e55W3PGdvY3z3rOtZEtPjC6KU/K5HQTCvzl73sa
s4p8Xdd8PRch/Gh3dC8u5U3uqJE9HRi/PWhHssVUrUmYyZPChc0jN6vvm1VULcnh
YGT9LSVoiWPou2Ry329k90MMWtXa1i4+k623/l02vA3QWkcZ6bQ+Te+jilwcsNDV
8LxtyyHr4HkVqP5VWEr3HN7OLrpApTBFH86Ia71SEq9XqzHBP5tp46yZJQc4ZUF7
hTBBjFeUnOioNjK4iw/V9MgRX32VqGn8cHRfqhwb1tfxo9swUfpbPmts1f2ToDVD
NvxA9fy/GgivCeY3rmIByqa84WvqV+iUPDKlk5Ae/q5lRYQ7CTB6IyK1FGqYAqXT
MtMAR0FpljylDa/DD8IAriMxc9y0PYAJa4bVER59kAfyuXSxzsSWxJ3R6xBibBt1
ms/FekyPSMzX8OMbrj5Ojp3ZtDBtdeZy5IESNh/GtuDjCn8rsXnB5EApIVogEKq0
HZuTis5HjsLOHtJNF+c7StQkhUTkI8EAMijOGtRL+BxGnlKMnZkBMI7kC/ngb4ZA
9SRfWtDFaAkRY/XJS43UuRs9Fl9RpcAOs7AFln25vDLtVwXB9SM/HrpG0OTeJ+N2
y5hj+PwlNV+LIjgcMgvjm9gDjjaL5OUUKz/ixWLDFQ6LzKTpnKB0ymkKh1HO7koY
go5u8dxzY41JQz2xPci1VKwcadhT679qyEbX4nxN5mYDuaRazW6wUEtd49BZc8b9
0agiKVGOk1ZgVjmw49gNwpOg8vrgkjcGsL5aOCCGzsd7svqrfNeBmxzanlqgY+bw
4vUXltjbwtjEJWNE5Srf8WvkZfUnHU1um3sU5qa6a/W379mZhxT22wQU3/MIA5Yo
Fx4X6oBCv6BG8iaGZo0IjiiKulSukzmJHF9LMt/qv79k/nGIwceNyFmTeUAdz1lR
6zgCt0HLACr2T0lVO18gEjVe8hRwj0sAvaPNHYbmuZtGkx8rpezWVq2iDAgJliWy
6toFGjyK1hiiFDFtXlz7k/9zBS0g0llhbViCzg8FZW1oB4KjJPnQQX08COkOVgv2
vi1Fguw4kq4cRDVbtswvBNzHvnMyUTdnHvMgsfN2ylKjcQc1p6rn4Two7GVMOyx/
vpyQHZZYnIAcCjsJQQBmlDrbZSt7kmk8rYrFTd9feAY53yzT24Wm98Ov9XzuXDi+
qxQe8FoWD9VuKwk7k9AxShyx0SJ1QGG14QKTR3oM1feTyxQfGMiOxX436Gj0pO7t
pKVPl2tTalrnDLkvNweYBoKfKxTTUyrfjXx9l/f3drV2TnOistkgIzrW8R2sN7Gf
pqGNCtvfPpyXpK8wGB/3TZnmux+ba+kOU8Ax6pgVn5hBH9tg3Fzv+Ea3aZzxKhsY
0m/FAMZiruTQ6wKI0Q5jR6xdlwcd8vkzcNQD93HNefez41LpykQT+B4toJdjiIUa
ljjSnbvJBCZdEu0JhX3pV9irpIzIStky8e8PN1lDKHo+C5neWTYQhIJFJFEPdP6C
6FmW/bEDkdZ84fcHIm0voPkPW2ExqmEYx2yDcAj81IaAHrWNCWTvxJSQp3b8/9nm
XvbR8Z7DdKyPRTSrA85l5//X49YTCUrLSuafBQkpaafdU+Ug7w6BJNVbwVXZ8sgu
lNpGlDpziaWZ6bmOdbq9egeeiCGjTAHm4xBaHGhKURh4VWLc6ood/zKOMF24c9Mz
TpOiZnLJVpqxxBifxaDJER4PD93OhlnTTZ2V38LVG83MUDKh6Xy9vYpGfM7Mg9qA
vYfKvnu85+3nUVd5NLIG6KmA8oRZ3EQaGtMI/9L10ZZKMHs240Mza4KzPy8Ro0SN
+KOj2zvb9En+JMhbDibssw9dw61rjoY3T7PwEsur5EAWIMPoSDqfan+KSHfX3Z1X
0JJ06Ma1eHxW4jtB+QmxTglPbgEx18JzWTmbgtRgm3TzC1vhQRJJkrFJVFwquryw
j+/jkGAs2ecox8oDvyiIsEhshkuy7a8rEE3VQMw+IeiCYTshpak6tQu0Vsp2yzF+
lw3RAKxjIwbzDD5PyIRO2gFMO/fiTl6jnXjp3jJmuQ+pYqU3iUj+XY+TqLOtk/z3
1y3n50I3IOudVtCXi8hETI0E280KszbsO22KzTwOPKnS4qCc2RvChMNKn9wU9Vbo
ZBYum2q+naAqvjPBYqrIfO5SoZCqUy6z7fO8BUW7ICR6IJjruZAPdtcnGP1HzaFG
iWPvXcRS5tMq0IN25oMvHDTm7OdIS/96zIknFCFkBpmrioNwUdMdZeLqAFpPXpCl
4SdWAK+Iz743tsxdMg2NmVDOSnTk05i9mco/oY7hDL9UtgpL/DDXkME3DZj2X1Zf
tU19OIsMsyf0hoXczJXVTmXDwbTaVQHLwF210wjRIpmpjaDSQ9mP530TYYvFER4b
JcSAH8bw2IYAbOsWTK+z9blXznK5T3g4KfRFc9BjZPf+kHfqhmNbh1NvRGsgq8GT
O8R4/3P4La63K+jNYq7M2vAJTB/NSfRNEfRm9bWM5ZCxiCCoyzf0MEe0NqJoXFja
qoG98sBaf5JGUNNXKQeOGnzrTBnAnH8QzMzGrn6ViZNy84luaLc94bnM737cZqo2
zl1dq0eHsufpfQW3ufXVwVUkJx9ZBSU7Cawsp4P2i8VyUEwGJYael5teHCUfnMC9
pb/yC3Zk2LoLhqrjS4OHnACw3ErTSevf9d8k2shEQaTcHwuA3CauU/ah89TlM2LF
L0uqi9Pz+0zNZo55LCeI90+Jbcxx4Ql4O+JNBZpuEDskPqvumlPFIrJVkvSzVQM0
EL1XsFcmSkb+Ni34HYAPLMLSIf8Ra+gRWduQf4gLX7/xWBWh+lu0exU9C+OkOUYp
2A02RHXeQeQPrpGM3fbMcwyV5Mk3tE7nIsYv2yWdIgSemtDf7Bub/7kkJCj85xvK
e0+OGGwXNWJHJ0zRTMuxg/bLdHc9AFTG5yroxSN0eHGesyWToSIlmTFcjP2Ke/uD
YZm6GGmEIyDNKkPwJ3x0NaTbSqLLLjsZm34dyucC7trH1dD9MR9VsYbtgrp+cR05
Xx4rsoAkLJct43Rt8ESsvk7WsYEFQ6Y+R+GSd4Q1hMMx0TIPW7t7JHjogw79iofg
hkNoaFsfRIccw/aiLb57CPXvWPSCdwkJOe1UYaEK0ZgLu5XrJo+PazG5Gl1gW91S
5DcnrQR93Qp5ws++bD3rqKkeae0yl9vYmc9e/eaXhiqgqJCGVMwq8V4IhMaObIaH
JMlzt+ehOOIdx4cW87JuPdR+PlQl5IUXjFk47sRcH85qImAY3jAqei/B2amUt09h
DhqjBFuzyd7XhsojVsDOo2tPRCjcgpuuAMDFSkMrBae+4q7+QZHsxWIq1dseL/50
SdijMkBrFIFv37/U9ehUzg5JgccvVtUSDDmwl4CJ8yKIq13bchE+1VUQG9E0I1+f
M04e4eel4zid7UwPPtayqu0iMbz91aCBhZnvnN1h51TtNs3t38v0svtqCbJFtMv3
DjhNUXT8uIroDrCM/s5KQCFVRTntajkLdF4yQbM6Gs5HzcWmSkB8rPc81Ctl522G
q8laIIiD9bq3LNk7R86nIh/Kd4QDB+ArRXjUvGgXFsPqSKW41TIwlBdatDzG1YeP
6UO3XHhSpxlVc4Py7+WhLzAn90GMaLQgO2d9Vci2g06eft405RozGNSJtxKuHamJ
hKb/0AlmBqc10d0OKDstxsbgck28m5xyg2KigcNrHGTLSyZPeZcF+peXqrBwIf7v
3kun/l1Cm8b0YWd5Wvs7wLPP+Oj8z871yegCBeHtaNMMnyUJ0VmGxg87eVaTq+Rf
LG5iqvIqtreGZmf+X5gSo6roG5S9YvmIzxnIC4w+opQ9Z+cunkAvWANtTKo2rmdG
b+BujZLmvArHLfWQrsqLthdK17mrq+7FzpuDEYQ4cNZfExyr71MQjHKKpeJgRouw
87HonRqNdzj4+gQLHffVK0MXxp30CHzuKLYnWaYu2yEwtfoJaIdObdiNNR0RsNak
U5jr6MvXKFXXaPRbtIKI5tiwVd06tO8ECet52KCpXu+gDZYju6UB3XPypj3jC7xm
lWKhnTahuxNWfF+9k2xAAPhKaUrFVy8LeeaAOPpfWeFhmO1x7qrsIzI0rqBwyq+R
yiL30Yfzzy0uoyNc6i/cESJ6LdHJ1qqsS1+VqYosNgjerzVp6pwJF55pCY5m9Eub
JUziJMWi4NeSFmBMbsm+oa4q9tCmpStmyKdYJctlQRphO5BS+7ZTs1sDtijEf+ah
Fm9qC+j3iGbe0M80IOWyTjLZCE9tA1y8rzJ32EWI3KengMMBx9xz/WoxicZkqcxI
jQbr9fc7gG1OEs4N8HE0iGZ68rmMaGRH/ChWivUhtmiV1sFbCM8y9/n99zOcMOh5
7VlNESAZMM3FtejtjG5U+rOtbC/l6lkAJolNIhs/68rrRRsWuG8ELE06IdfbHSpJ
kPebI3oUvOiK6DTd3Ubwo71765aPlIYiL2olIlbecLKdLAi7oPqBdChIFxu0lNx1
ovuyc69pdX3Y43iOkklFReBXKnkXSzBVbFAbeyji3iLef2a3AB3dgNMC5tdm9yox
J1Qcyt+VlT0s0qP/NSwW0PCqQomMj5x13yYuMEXP2lXyJbDNxoVhnIl75p9aMxrb
AHeIMV7VOgnUT+tHhP4CXkHTOZeWdztq93SgHNFXewvthRiJwGQh3cKZsovvzgI1
DQ8f7/uHiM/b/t58W/WFEcC2Ju2PGRwjrly2xDMcK2NkMQIcwFFfy4FZ8MSt+96j
hNcV8w25/xdQk9lGcSz+8Gystb/U8PKaKx8dzGabaUW1TyIxc7DQowJj/gjKFI7x
x1qO3Mm1rjB05AsN/pTDcU0xuvbjV2D7mapSoRUoF1++8DvpQxsLuBbMPOsiSlqH
1CsMdfbk/TSUtHRytP5X4RA5C/1+RoBGH4owKNr7ZRpAEkQ9rC89yY5uxrf71PrO
EKs240XldUJeWyTgo/lOUk5HqTYrzA1/DgBzs+dZgaA0Chtfg30OV1cjr3TlIt+G
HEWTWGkWheX8lCCkNZsVU9eeoOI0TwW3FHOZi97236V1oTVecBI+JVJ1Co12psRP
Vr6XCaXYFjloJZ03A6vS9kv9xVHJjDy9dfJveibmdK6N/i8Iu2eWO9yg/qBxDPKN
xq1LNZU3mhqOX8qCURK+0cNacCKp+TSLFbPKbi/YoBuLtGI48jXUOnXdkKAIsxdc
NePYV7FQGO069RR2HLDxS/0TbiCTI5xAL6iGwWwJRi4gEJ2hP2KRTJFif6oEcvKW
KR/dFUkn8cFpLjoukz+pbxst0Eu+88hZIDY4OOzoGSuAwaSs0zNf3pjtRUtiE5Gs
R9N2sDK3484otqTIuwwRmHV41iUrNRMPfhFHVYJoLJcBuaH/y7A7GHXyWuACJv4F
kaeItBoYZcCya8Mz6tINCR0NChCGg9nIkjQU4+r/uLyRLYF2API+ID7uMLbWeh9/
qHCIByS813Z36I0HGBkcdSauYboOVMrCHNPLGAj44DS+ahhVXO0GRxbylg/jt5xV
Lpj1rEYLDiMTctA+9q7O6RBUhTkxbWDU2KKJ4fee1cZziDidrB3CaoIi0pQJCUyC
KYL8xoVxLRVJejPYH6/Tvc05jd5QvrQAen+3yHuItiDHrZ+cRd+xTus8aNycBzkq
tODA5gyyT4TERfcSsyLpcENAQlE1dNGBSp5WlU/GfkHw+6lgdmsHOm7C4F39FVKe
vl0Wce7f2jbUJiibs0IndG4QpPUohQzbUM+18+psiG9XFSGC4Q8+/XHBtMIZFSu4
t6NaY6TRPSjTQsaYb9S3A5rxlEy84LrzTWI7AXwDqHvOCxjXNThQpA69JI0EsXeL
w89Vq6Z1NQk+BXyTI1Yfb9NAHGufJUd7g1h9YVWD8YpYP96ITltswRiDTyMtVKPr
7zk/3OXeZ7xJFIlIDGGLvwYzcXZcXIOMgSvKxY6+sPFq3aRAIDSaqB10fQNFFxGl
vFRCVrtkCyBwOUWpaMIEggdIHS4APRT7WclP/qHlrxjq6BYcXDXlA9WMzL55cztL
csVf5NhfDvgDhYln4DDG/584TpAurbBIx0qhmycfeKWVrDGCzU5EMvTW1JhCdW8+
zvLmdhAntmIFXYQn2uv47eVtcA8iCx9j9u/GUXrt9qcIg8oavsq+U8GoZvOwi9Ad
jBOV4He6meie2+RW0krDc45N2EHkijHa6p8nvOuk3v7shjgOudl5MtbrLwfQ2FwC
+0MYYnRjhu8Kf20l2LlpVpsKQ73zCBqIuW78vrvOocZ3ojSV5IkO1STJegzHW8GB
/PG/BCy89ht25BzNnsTXdGOalnKmwkXqHymmMuafpETqHFRU6r1mhq0LK16RH6OS
R2/fJeAp2uoNLQ0XeTS9y7DIVT4CKHc0K0Yk+cQ/Lv8bmTXo9mnWTLg8O9/ammXq
x3v+IMcJr+yX6Sj8KXQ2kl5FnyOi3OoZZxoyZDoFBQxMfDoFLyoneWkmft8LFkcx
PmR5ZreqsI8jjWjoJbh9VZqKrK4rNLewoqU+yS9EFtGO2Y/6WY9ZixvXFDxyKzLb
Gl46S/irf8XI+5Qqe5yOwwK3Mr0MJZfaI2m+B267XsdrLnBohrKMAF7+tG2l0q9X
BJjidal/uFyJp3GtzC+X5tI4y8unAhGtKj36qCSgOqSleH9qHjHZuKNz6w57iwi/
4qwmDREBzG3lEJErkfqiTAe9hJx4iV4SWNGvbm7qT5ZIJ2SlZCE3WwhvuqTinwaD
VCe54d0vBxxI6HJhk++f+2bwmjQmOJeLjxXtocAdN32kTWefXKSOAmyFoxGGHAyB
xmQeoZXzvJSEWGcYWNGj2NfIFTFFxw/Rv+FGEkdyPkjaA/ya5E+/GpNivQmM30QK
5N/hd7Z7B3dJ42iHVu97lKPSGJyJmF3Z07ErL5/A8RtHoMbub48BVbau6/oojVo+
hdIRf0fuFwJFE0dfLjUkoCVJZPDJGJR10rNEb6FVXf+xiINUb0J8MkClw5edRYiT
/eaeFLRiNKs6Dw3q0noSXBfrzmVcBUhf5cvi3YpNNEyz2yroiStHM0ylDF/rKdBo
kbTRxYFyOQrXhsTzo3/9KuiMZNgHBJEU/dNF11F9g5R+iDWIOrmllaXdfUpU7ava
hpnz4xTgOy9cbxMUxdLkBQEsxgPnpTTs4de1JYUUvTUGwWS5EhHWTGApuSS1C13j
BzOqnRcobVVUgF3JvTXkpce83YPeklhhW1LkqsejgDQnCHKZToVB8LJzSZOHrT3K
MdrKGStZF81EsslJuBo+PUcnPrQoWKAJdCwr3zjoUZWCclG54EaBZAc3x2sC/xCL
4uaiEEyyh+JoE2JEQKogBxhScc/9L5x5HsXA8SWHJq5w7qY+FYuimLyNYe2+gs0U
//97++oGQVNYBnV5DAWpS4DxXsgSvt8bWeZJI4fnvBTPSmjugU9y9nDQuPTuBhPE
LLAfMAzia1WO8fXyisu1sISw5algErzp+LV+MIolSqLbgU09EL8JF3hYZ6IRQcVP
ZqHL6f/1SEE+jF9vff6T/4jjA53vwIR6yLXhMOeyUtq0kVN7e0SPBmU/XGJXAijX
JeB9I38jGwLgZM35P5Ux+2ZryKNW1sWexNIubGGzx6ynbqFeYye0Eyp1xw9dlTLu
NATIeBQyDq6TNUmjAVlSzpalUmL/9+8Xzf+KluUBqWSdw0KpCqGWKBJHkg7P15hJ
ztJ13BnvsidAe64sBw4M0tGdeIloPDhpW8OrtKADzC2lgT4sWRd/+/PtIEwXJeR6
TZegfHshI6GxK+hVPJYP8NIY5faLQ19MfPtSqwxJbncSTVmAbNsOtD79ihLVYPP4
7z6pZJnhUlsxyBLKfdAvIfYh6i56A2xFxhpFXfXjjVzg5KBcq/JK/b9O4ThCqnaB
gteyvBErfK6XM2/NCAbE9FJERNh5oVlAe27LjY8kJ1r9L0bosWiPUy+80XPxyl/m
oPPCnrwMaEhnhBnbzq5sGF8iuJveBdae2FEx+BvtodtNx8PQN7jdYO2DiNfABIyS
2TZKutPlN+iOvuVCZmouhvgYHy9gxZJEpdq4uwBuD300F1oJI50UhavffkzXZZwK
iNaVmoUJzOkoZXtD2/QBI+5HzgYcLAnEyG/ObnQBGQcL+S/4ZBbnmJgiH0P+CEaq
MA/guwL++V8jbW20OuTVtKdHhuj+xS0f8UXVNlE9s9of049KJ0+0xQ5NZEQOo3oy
nsGEeOs+Z7Cqd+RAGCNhpqC/fdGuYjC0t9BRtOfvP8yv26Gs35uiLqM5oy22CA9y
6RU4FbR2ugeZGg9aQCrBXkRSf/VmARxfoVJ5VaMyVgWacY0jT8Zvkkxg5KcSUXZb
v50OYbszstwPxd4NXSyXuo+cit95EE8r/iaGdOlanihNnKtZuLfyvUgg63SPN4ST
e57a6ghlwqS/OHJqc8hhWyk0OfgBmJicVexn+X/2sfaOYdHWc2XHINktj02uNDGE
DQ9wSzdKB5fUK4xKvFWm3r3p8QMEKLVnKYnxORxFYYRXST7C2whusCrMgik9l+Rf
Yo8cP/pltwh13+Zqg8kccLLL5Uhr/8V5f55uMW3UyHiP83ht17C7zspAi8cLZZky
TkdItDm0Bo/0WTt6vzc3SH3/dr2bys8X1my63uGem6B5hV7uBBr4ChC0MNdu/gjv
kHseZJtJ0Mau22rDT4gAkRSnAx4xecchwyeB6HwKODjiEPD5/F+isDiXxT5Tj07z
KU5404cf5NAR4RZyocHo+3l+I1+//w38ckhmgPrAYSVqyLCQVUHC4tICexJttG/J
lwikkvLYqZ6HvqloLAdABJwVq5KJ3U09tfeQXJNVjQmBvaOFXTtPhNBZRed+y0Cq
mKk+TMgxj6go7QNDIGlVSAaakgLA6fvX0PTvDXVIIfLgkZXzLXMuZqd7cyRBoXvn
AjBmaPIK59IzVYhJJ8qIdvAEh4NrOdczn6MQO+HTRHBlu9lce/AG2UzEIkC8itSS
Is3h/nQLYWmnlpSG+tw+9zAnFQmrjH7HePKxpnv1jer7IVYC3XMmbS9atXXD93tF
QIao89WnwafqAi3moi3Pw8SMi28jYRvTe1H198w1MZKkUuQmKf+zb+11oJsAKred
t4YYd8wjUagB1sWJcEnGll2jBoq1pEfjW1nJtwsh06CIxe2rdnSvq3Ix73LLkw6j
gDmonRmfKxJpVbYDVdMjrNF9F5WzZMM4i7cqV2WrHmG+3BKq9xlqj8oWO2ZSPbPT
RXZUnkB8tmgnh78lW6xUs/F+/GG/PY/MrLPl08oEwicEmPJzdFcjM6DBzKWaYGc+
77fzx5KLyB5Nv/ixTENuVbq1kqA+odXnDTBpbMzcgPa+nSUt2Q2qIGmkiEMSv2wA
CGJEm8C73lHNn53x5qkJdPcvmVS0pSb4i8/WUJ401Lk27nA5NDJX3fASUmtQ59VH
1vUiNy9JN/Nfk3oOQ+4wW+GqIYV/SROuh9Jlz9pV/gPXR2Mhz9kEYEXAs70t79Yz
39wWkvVMn2umTgpefVAlJ24yUHy76cpZRzhGU3U/Og+8xjIRRwnt/1WwqS2C4ULL
34qnuLnhr5m5G84Sg2+Jg+1L5D3zVFJ6z98JcN61FtbyLxsVulBvHx/XxCVzzRY2
x4WIQkTGb23Q+ollaCM4vm4Omg+WjwGyakdARPJedPvn7LnFGQ6FG/M04ahS0kDQ
/4LS8LZTX2BFLyLZiqDf6EPoe0A3lJpVN+rdOtS8UJqLPT+6CFtcvlUNjOEYE/VW
2ZbUokBrxMI0kf9w4/AknmJwzs5fi513wPJ6T6fD+/wxjrN82Tc8I+Wy5E+IDGG0
rK560VbqsY6MLoG0TaaWkm0aGj6iCKyEOnWTsrozSspvZulTrMT6F2IEdQ6bVv3z
NwwTqaymrRN+uUeQ14k5VlJkJXeVV8MkNEzoCNy6Qjp5pDV2c2s95tpaPd9m9+tY
Y0XZAEGB2bWy6jCkoNFuqgPhUS9268hPs2qdszU217GqvfK+inPuoRfXO7qu+kvb
0TgtKhTAbYOBmsUsnPANesxa3SAT/VGqraYcFxZ62L0szOqSkb5h6dVYilP8SVIw
sGdDZtu82YBWS6FdiMwsCZgcQSSPfNeMgGbGv9znprnqkUFqCQEmqmJtIy+hPvrg
aoF/qDlw0l+n2AvIp98p7QyxkduVwYADEEpwS4llAxEbBR5nC6hqJKT6rNQHChCn
5lfPRQ+4bMCtftlByyPAvuYdPku2FrU/W4LGC4Ke3RC5KfBhff8rVKQfNLMrI+LL
uHfofiRWbsiMUbYkHLmBpzuTc58Elud4Gvf1lW8oCPDE2lICW4zk12qddz87xG0H
fa2yNt5aD/8guoZWo5DzYIaQJDJCOObEY8XZoQgDdTGe2+czwLDCLIGrvCBBkxu/
8yf914NBOPV4VPw9K3R/vDBcvfCqQBhG6wdJiKytc1PWb88uzBZQXSZj0y9AHU14
s8N0zxuUkBlNZpAV8wqP8voseyIh55M12rDvqKTjHFBBioJtXYByw6CDT40iKvGh
mXjvBKw4HUC50VOq4/z7eIYhHzI/FqH5kVLytCk47Oy/8SjpTid6mesoonpCtWO7
hsDIhxZMs3IvmOwxFewApwBW/t5+iT9XAZFXFjwUr4U+SxsudDsAhD/M9ZvcKEAK
Tu8t8eDWLBiEk2omcmZi5+Fy8wX7jMMElWC7UOhKRWykDWxWenVixbTMsn9Aw/8I
FJdluN/IsUpIS0BxhRmRHhhh+SFE7/XQiU4njwIPL3wPxQDIJKyGXtVxPTMp5Z2H
p03lquK3790cuSBPydkl/eC9+5IEXOO94CLpQaN7MXihj84G1UhMc6YDjG0dNceG
R5l7Kr8KRp09w8evACaUExY9TDVpR1E9w96SUQiKZ/+AsF+tWBOR6MSdOx30uu2c
OA7YFYkHclsVwVuhOTX2GLswvoffisryi0CoRlKeLc83nrJUVVafRlx2Kw9TJAgT
Vgxy29jiGu6DEesLQr10J0GH3+yP82uaSnmNbObxKK8TCF14ZUikctOBJItI43FZ
AAAYxruLQ4SgbRZO7rfVkRaPeefg/QVnn2eiAYH20DcEo72ULsZNjl9SDw0aKaIW
HI6/p//qwIDYcBysuwSzYV6UdJVBYeDIRuQ1HcDRo5H2f48tcUG7ant4AUuhec6s
/fy9vkS/NCbxqI61l9Nrwm6JABgHrUw546EWxC98JxMOUVJYHRduqkUjOBGilPRl
btsTvQdVw3SXIKXV1B5bZtBNWxRiRe5NQwoiVc3EYEcfhYtrXbXZ/wjydgbH4Xhz
68iEkQ0kJOM4I74QoPlw5miyKDl+04q9NeX1ijDPaUbY2+oQqEM4wF6qJAu2SW/9
XLbeLlqEe2dGkpp8C7S2iCl9i+E02B8pRJiyYGgCj60sVIiWg4VuJhyIINsgcDUM
8dwXEgFGdsQDqCBoRcTieBjsuNIrdm303E99DRGiGVqhcZacBxnXW/RTovY/EMNH
5MONxxUB+8GO5gd1VRjHE+Uytojsc377FCeMm7gkPL5jmTV1rXgawKHnwspVH5wV
/fSR+U1LFGPLah9uyQX5ECSMGNfqc+hBZBlZxMFnoxqoAw+pGmZZHjCcYJwCzF/p
R6QGD2NrKHujendxqvb0ePKnsKFpIcMxhN7JvAblYXeAIRVq03Yji9gVRxzjYCKb
PULlsgCxC4WPIPpSxCNt+z0GB7nOtfQ75tZKvB5o+SBVFSyFnA4EPJsV4d35Ttea
swL32jRoYLjRi5yZBwEccuSBDc3mjk2A6TPk8zaKe/aybRkxKfrFuhDU5S8MqekG
sz6NSTcpXSLHAHyITE5P1Ql2EfdPuRjjKSpqw+ZHsttXL9iU/zcgiXomGCOSTJNd
mrxB/t5aiXIsk5UiYT12vXlOfGFTDZj/7L4BhS99PhYMcGUEI4dYECVXD4A1K9T6
qhMKfTE6WiNPDhzcGf2in4fJuNoMOuyW553oCXp5WAoQTDWh9ThNUi94BlCLR9/x
nkICtjP+Laoktq3irzVXmm/hsnewz3o4fKGiDR4Jdo+AwUnHYtk3iSo3Zn3/ZnMD
Vxoz4R2+3z8bEJB60qxC/6nVs56/O4iyc7sf4xmm+h1j+Kjw8Fqhid9o7GU2PQQl
ttq7u41GAltcMLzEN5okekbOeCFjeoojUw77OvgMQLvzqCAkYSQKOA+U7kXnb1f8
X1zkihTModKcL5joRWvXxlIyYup2I5BYNTJW6ZQeh6HTmXBIUs+7/m/1bSWQiB7Z
dkw5EM8M50TRjE2czk8sle1WMQ7zFOpT+K9im6u8bcUUlAQaxOUqJiCJbjlM/8dN
znX/Sgvu2mUOXvI8mf0Di7FqUKbAgGgbFRorYaXerjS+TG4MjPTEuUf7Qyjmot2D
+eJ8RvxSToW8ERt78e0qL+3z3aucZEu8Vo8PXV/Cubc3rBXnCVY8Gb4T2EVr1SHb
nY1TdnBDDeo5PBecOqhmW66pCVUhXPkDRM4lB0OTIIUZRIhE5MC92fJhK5cg7ReQ
w7APDxna+aQRs/5vG46XVGa90Jn8zeG045ab+1rmnI9RYMRFEjVKdkqhUHHRj/dO
mjZTVlsGBWQ3YGB2oo16rupbNqB8O7F/74I/g6JNSkRR2C7xxAa7jb/toCgGbGzI
asfOJIVCen1XnPSb3FMGq+QTsvBavHIC90H9wbKXJnwxJw+Nn0Vp8qY4hfnUzxNW
hHgeQeuqR5zKx0n3uiPt/ZL0RASWNeWgwPsz3bOW6Rcbn8az7CgG5za8jHccNdLl
6aQaD1/AtrsYyfOEj6wdiaAxSEUn8sVOQdIoWR0nzU1LDZaHzVDn7CeKIQ8JOESN
eXZ9DrjJtRg4PwNAuQ9Wbd1ecPYPLztfKUiZdxKsYYOfViJ4dIugsw1Ebz4/yx6Q
kKBTgjkBEEIxKafKfxz5n1A0QCntwMBJGtqhcLe6i2YKSZmTtA1Vn21yDj9DRkXq
dKkhAfNW6JylNTIRMcjezQzncxueT0KWk+7AJRlTp3eKaIuoC9Nyyjkn0pchhJnT
GsnQy3kcWBcYpiKfkdF2A9NMXRJyrtqe3wAvn/mHHZs2eJEkUm7gfJo3gpBouolp
b18D2dO1UFNFJ3ZH1iCqUGUKLzzYIeF6MuJQR1ZDwKS0y/EHTS91aRiiX/RFCvDv
lrf/H5cP2X3XBBpWH2clJgnF9gzW6AQmQYT5+9PC3tDO1T8ASJE4+Wwj/v5I9SeQ
UwczClfQWoizRUJb2Qc8aZav4DduV6AjSxwWmEfGw2+1wyuN9eUljZ2/DAOVzOVw
n8HtmcvZ+KgCwoF/0UQE3EAncA2wEtZENJ3hwfPh/HBT1n6tJr3FoPm7eCEslpWD
7xqayAIP+PnWpvxFn+IgQ4BAcTsLKL9GGQ/GS7k1oQQuV2M3RVOENpIRGm3IygF9
i9S1BktMw6Gs3qEtcBmqhmFB0Zo44yfYukNJ5kPRnpb8qXh3hA9TJ7smGsi9Ds91
7HUnmhKKPEWUUsz5GDO9S8MsUgkQpNncFLXXbD3PdhFb/UdJaGmPnu02y8b5AB65
DmTNlLBJlf6sNMXWjMCI/oqItLWcpR0d4HhSspq82Tx+xpiaNsH0FEY3ksy6ckJn
NWfvtUNX+uFDXLk7mcOtY+dtUteH0ziE+4sI9lztGRP+eH+n2k3LE1+iu3zqjWkF
w1DO9ByQIc6JeicHXLFnPDWUkfL/iLOG/uy/TWZZHnoMBH4i8IHEOMev5TZYeu8+
dlw9/4xGenPR/0YtVVhVDgAODi2HCPwv/B7yoh4I+xmpXeC5N0+tOob4EIVukMKU
gjh2gtWgBjbt6Y9LfpSgpWAqitSknp61gTGOIa1u9b8tp0kwV2gocFlnbvOmQ2pF
6snFr8s1yNXQDx5sBG1qs+zOfWwPAvJRg/9w1RGtidVR6MTJiQR/lTPP55la3lzg
Qko6CzWa4Rjki9q2zyPa9b9yv7wSrdeF7/8PxcWjotr7qyL1ExePRJDjL23ea/Gf
B18ua0/Z8012MWqdQxyeCdPz7j2f4QXKlJXQ0U9x8IpWLN7VpG3t6lhg6Yg1VIPn
Eg482oga1NdXo6rDUfsbIVDOe86ULnJR70hfOe0z11RNsQsAb4MgcEjBTZBFv5bV
GgH5DflIrtmuVRCIX9aE/g4BKwzn6OOdMJW+bbc9oAUnf2sQUZ7RPukEM+5YhgCG
Rq1yTwJsJVbnK2+JhRp8LGyXw0DWszaxWISIqE3wLXA76TH/+Gijk6BWxD2yNDd2
nFnrFVLiHQGpn00SxpC/W8y0bKacpJdi8+JZRdXy+3Gs4J3mBlD96pFeXltJbDbS
08xftdP2JFfnmX2KwKXomFFuAxWOtcqu3U3hIuNde1jja8It4ZbHx0Vb4dVVPjTL
pQVEGZQtmKdIzNdRjnG/Lqp8x493klB+NXc9Ogmle3AiboXQwCBQ/jOwMb/QLMa2
7sp48wJcwsUAcYOwnsYUSLIUNzJ7ZJKK80xgRMpRj0nC75UViKaZELv6xweuTnP2
MJo2Sw+qeTPv0zRqERcMnHv69qKxX55RVQJKMz7s9zf5AVwWWTc3V1A3XCwWF777
zoiGsBoBD4wsHxgz52PWVw16m/XsI/9yCCyY2hmXvOtiquwLosaqEQ7O67ttAag8
SwmVJq2oWdsfdQtyb+t6H4lmMlPtsEGz8G4aU/0PDriiMDCd4PmVYDEE+vF6ZIdM
OXItRaEyAPvm7RLgPr8AF15ptOUOAr+XgHKPoePDpw5uDdIfHhPSKXtx4bRClkp5
8FyuPeLS+47pgMwlEZ30STGdkP8kkz5WiAaw3iCXGuZAy2mFYL5sSYi+W1JXP6we
SGLcd7hchT/BatAbkNTjjAon34IBY2xXGoGElsHsc3MnvlARbUGHsv96thyJnH4J
mvN2kQhzTfsnzc8q/uyxJZc1beYvIPW7/USaZSbKOI7WtfSZMq82TL7DGYb/fBi7
2p7DeMvFgbtZQAUC6P1zXX6GhhrcGtl/ZFbHsVGhY+jTqwjEtpV1ivaE9nsyUmyq
+JW1sjQQiBFLwEL28McMxG6d/pt7O9sMP2KT7dD9/lbb2BEs78/ao/W6OrQl788B
vuu7ZeBjq94NXGhqdohfcBxCtVyM2vncw/T9HufuUJ3ft1GqJRQ5gMTZ469vA1A/
2EzkIUHB+MJa5MoIraLfL3J376RuAm97/UF8FVRaoGMfFh334OCis37OUcBliPPR
g3Kge9venu9MpiVOY70PsbzFoCxOu1sNlQA5+uqaC0c3G+YCj+Xuu2DWPmIW4qiO
HqxZAs2r1BTqTWRuGGtGlY/N9S+NqKak6zy+jTVtcR+mefyhBESUJiolFTaujRtk
+xBlRDv4LWkHyugf7x5zM2b/F+ZA/5xj9mgiCOFaT0K3O2tKhLdxPuWwmCYhmsxe
+5jKGXOvKVu+0w9FlIniT327ML4IeC63Z2CQC75GTvxpjwges0ggEuUgiiIXROVL
lEpb1eT7/GQBdoKjt4l/E8VAjGy6tR7F0mKw5g/Wamu/Ak4BtCU4MReGQoTUOL0K
0crPgrSLj2vvpIF42oy4KWMmXSVGcZICeXkdC1QBSTShommU4JgDww09hH7BdlZI
idYAwKNQr1tVa/NOd90rrKLBRr6AuGYXEY7XaD0o5XdlyPt9poztIG+E9Rm3SUcp
xA9CgjvYKIZfJTUZ9idfz8CXuKUMZa6kPaGLrArT4hyB6/V8zxHGzwWXzxPAfM+T
IAVnW3xd4qqZiv0F3tLO5SB57hkAk0xoPNVymZ3khfI0nkopZzlY2RM9J3t7kYQv
l3XvhA45oqQmGs7KXBIkxn9Ee5gjLdscp8+lQQPfU7dYAuAFR2FkNFjpVLm45i5h
91eBwwiCy2Tdf6+0lB2hZd5KFX3deLePaiKQ+qbALIJ9PW4Lh5JPAbxGE/yAnv2K
Cmk2PCtHAzRqj5idynqRhBaYaWSGWDIZF1ZAh5CkFpduSDjymeScLLjo81NWTFRD
pKbIz3QOqijB7QunO6/LFJMhqYU69qdBXoz3n2Rm2V1Oxuy0OGWpIudpvcW/1TKU
pMj8VDoD9dg2RQvliuARB/iHaFrPNUExuO/Yl+uPRqUWAEEOB9kMOCSBjzm40rxN
1sskzlgardUHABUnNk2X82ARlE2fd1qy9R3cqzbATuXFoY+w1aqq49t427mZc+p/
QZIRBQl6rnZPfOC8r55rPOEYfapgdQ1U08OovhVhtL4Vfdfk5VdBLK27eL8zn/Gn
S4a9uAOKv5QsrTw1Te7OVZfQo05PPSxryFDLVdQr48ptvB7KrzEbWcwqJAlMfY5P
yEafwTN8dbkKgSJlaNQNazNf2t5XSrcGCRQXyCvdeDx+ckbWgaGwHwJR74J57lIB
6fbY0yiplSklnUwuMS6yzvY4S+bnv2Pq8tdbLYn8y5caZBdfCsGQwdiLvzXiw8+Q
2Kdk/dkG+OsgrdWKAARVocT/KF8HXKb8YXYz05yWL6NtMZucWR+DO5XVTrYPfgDH
WiaDZJWl6e+p0dstAnTvzJ2kWZpp5i3E8N7fH467GOG3sAlDfgy6RokufyI9KfPw
x53PHJnwx37ZQ5EDKaEJyloeLfnwGpmHvdz0b5fcBbcOaHDONIxdKkoD5YXhjxWh
KYD0xc3XFcJw3LFyLitPRbKyvL715xWmb6Iqi90GwJTWQYbCuEAVf08t9F8fUUki
w4NRjG6wkP0W8hhTwyfW6284QUWL2fd3C2a9JuBHSgKzXo7+QMEb4nz5BUOi5GEM
ccOIGLdYFQrWmeQ1QHyLpYaTm+0nlA9cQaIjy+zt+s0HOPJPZNZkjY3fcQTd56Bd
YcorL6RRj7/wnjWlPPExoCX2FeI7v3Fdnc2RGLIZPIz6PZYUCTAdYmMQ5WaH1pab
SW4w2vcDmKFXntWUT79vF9SY/pg68RhrayNGbj33PK33Zig75BUhvsIF+aXcPPiz
jOGt3oRuMVowJ+Pw+idO1uVFpU3egLzGZvU9z8c9BGOO1zI7bf2XWLi7MCKiFNZO
44rsYNn3CREKXJCsrHuUt3Afo4GRFsVZF9naE17aynHY2TMjd6I0b+7aOJHY+DiB
qdkSVQTKeySMWDX4WO/RmSCtAly6rSoerWgbufCBXW9mB87iBqCvxCUD+N/UILMH
vX0dqxZsVtq1TY2N1onTDnb0hUh6a5BbVVJ3k76/MAU+5bTEbXzp/R+kM+tr6aKG
hwItdXa6n+5GzWnah/oypFNyRJaVKwX2t5/RQIdtCELxEq37zg71XEjIsJ1nO+dA
7qw8DcZXv1fcy4apCvLiLWkInw9rQnZGTkgSZu24VY353Szkv49tZ8WsxIVAcEfG
PYwlTTVukOqroActDW95HCF6ZbSolLNiHGu0oHyu7/s/SpOvvthWstHS0qfbAWHl
KKzEn18Jmusg5ht/IC6oBXsWn7tmSxVSz7KqYYOOy2+jfAroBPACoSWHv9SWSasA
oBkHsmVjnSxVhkm/ZgG9Lgk9RYSmjmnH+J2dboiWUsCOBTUkey2UvyHF+07rzU9O
HZC7+vcDkEz+v2KEUvPmeSI0mCjP5iCL+TTJCA0ihcinp0rJjfITa4wb7DwgkTVs
KNvTP6uK9c0PEkgSfm943IXJzFHPblZruujQTx2UaRFfsQuk9AblG5tfGve2Lxv/
5DAwEZTJboj5Z15drxsUcgigcq2Ye/4kkFPY4Vwbp526pnlTwNV7FSuObvLCkbH5
WXOj2JV2atHq+TmwmdTc6SxJhAnar571w7FMmCspmCfxu0GczhQiHU2cQHDWEoEv
n2G8Q4AeYyp0REQWT+UuyjMLwPNIQGj8qzkc6gvdnlNyvcPnY6Wkjjgb8P3gzg3k
vldjSGCg4yw/M65IGsxF4+WZCWL14Z6EojPXnOCyd6V6tpSWr+gRv44C0NjnJo3t
B3DPoUShvFMxL+ObIa1LtGaFMX74mSbACmEZ2H/4J8YaiaAwIn7G3h0a/FyqB684
pkQFtIu8MadFSTGlvPksrC8Oywml6zz/61PnNQJX6vFeyTnvtqq1rZ7+frgAtCDh
8tMo14AAuTU8fXD8kV/HqVqaTEbYmWJt9Jlg1jl40DdzM1+TDOHguVe3KPSj99dp
ORLdaZlhJTTmGO99Lcg+OC/+10VVaO+N9uJBC8t1n6lhLwU7pSh4qNa1V4IH+EKB
hChHryZv7jFDcp2dAAjTqbdVmVOEE9Idy10ykTLJsQpNsG5l8bS16phiQq+I+QGE
7TR/+SfZ1++QOMB92EYesO1w0j99oAQypX1wZyU1ky1N2TTYHB4WhQJW30CK8xhR
Ty1bn4LfQKemNTtdxu67t7ObrdDh8Y11GaxfqnkQG+7izh3aUcvyeBgAbkjT/pf/
8KGRSc8gGlyQq2uK6zCMfHGiJg1I2jxKbzF2vy5mmaXVYDZDGSd940Y/xD1dCiPh
LvojzuZB+u3kTJUyzN5jGBJ1M3n6apYLV5Pdtt01ZooX0tGuppWV01OS1/VL5qlx
Vw06hj4Kz2kpl1GGhWKgTec2HgNBPlRQ02mo34uKq6mRtQUzsEUOJx30gCwMVw1i
7VYGPntgkEya+vdht7CUdgJKdBMSut96I/xwhFWbfgDO/HHK2p6WWAmtpgEhj0RG
0KFEFeFwgSjPX+t5VA7ldxlkDoAPdYK0kQ/fn/Q5R6cJt91AjvTelWNfZVcUPxXz
l+xXVtS2gL2lAMltCpp9YoEQPmeVLcoZ40M8lQDvbkc4euRBs+f5sROjhYKsGhMy
JS4AlIXs0GJPYb2UO7i+iV99QRp7TD0W0QecWGTYzH862l8OycY6WM0I/IQ8hLnS
sCJ2bvaBBi/o0mvGhEzrT8Q5Dg15iOt6PHWHLK1EOx09cTwBKRk69M4fdA/6ltKy
HgjFUN+Uo3m5g3ESVZ4VukLXezzjTvI2qPuK9XMATBG8OoJ5xqeyFF2G5v92OFyv
MnMtArdPhFGOseWDKB9Aq56fYGZknwj37gfBLUleXGfoEowRZpzGwZxsZSxVgpOI
jTmGeYtpRnsIuUdmbq0OsuwbVmz43WoRhEf0sMP4NXMWJncpGTvQOfWO6y1GQU6V
CVhHGXt0CBEBNFV4Go1ueh2jzD3sFMo9Rp8dhnNiKDDk1xok3FM94zaiuGAvBHsT
TWNmkylNk8oyFvNdjP9LA0q2uoMKoKtmBLf9I10ot1gNpqzhYxflP0CfZZbHwII2
e+8wVelTIQIpfrOM2iM599pq62vyGaF5JQ6QVf9k2B7/g6EWDqF9kiUIsCSt3yZ3
WRJHth4UT7vic3x08ePcD2EXPFgQYZY7zxvxPHmBm3P8aIYsY+ojr+8cb4Dnambv
57cHYmwnD2PMP0QaO3KknCurC3TopO6m5k17FaZwbzlabwBv0MN5iNiBmuONSnvF
A4Z/sooaKXiQQTa2iAigbvmhsUYB+qEEOibSIoCXOdsqDvZWhrI4ydIH+28pJxqV
u1w7vrPcXya6LLV2/wZx0aqnXXQPDKIoRUWbKPqT/hY9M6bB9hWT9yKBNC+KkoiJ
Q1QQkZ6NNQiin1hT5RD4wK510iUx0e0PVLR+dgtOUxX+8my8z7vWXlOhghyBkyNz
z/7+b1y5+JvPLRaz0J7u3wd+S6VbUhhm+TMNl4GIMexeUKhS0oZMsA6ns+1Zx+lj
eYT8mM/+FVkKk4V1dfYdAlMrjOCuNaiOyN/fLSl4y4oZmgXDoC5AU9CY0j40nkR2
D5mw3rWrSepfiUpaR7wTpYltH226xtudVgga179rUTH/3njRnZARluUryYNTPP/5
fOfD1GCuCHOCWJJxoWcsM65m7qhjobyDXExoWZSZUpukDZ1jFavOsG2ZPSFpsLA9
/85eKkofv/Z+XKKGEhhjzs32cXBma60oC9t2sZnBj/c96+itSUrbuOFo0x9CEOGs
pyfWLcREe/dgmT3g53VRBUE+ZiNX/DO44wrlwQpSjdlVU2tcE3sG6cS5bT/KpvpP
D5PYPaPRcbN+4ROul9DTE3GrySxVNN12qpegwpVDCMXAxdYcLStjF6uZinASo98D
aqpTH9uXhKxAFFk9vuIA3EOAH+N13IpHpAF9WPxHhbBPuuSJZI22bXn7afCr1jyW
YBIOROAmqYelamq380xYcCkbZaP39BAKs+GjTtfeNktm20qyC5u6rFQ7BmuxpAG/
BxtM4j4czSlDmJQWYe6xhyHiSRXiifSTpTNMMt8migJrRHxNQh/xKTTzpNuVvwUH
HD59k0ppvObuGg4EOrW7Qm+c59g4MF66tkyr4ev5PRbiRLIZTxO/OwvQ4gCbAaTK
lZKxdKfZFf2KCmIs3j/8FzB6YbX3n39ysyRQP2rFwrGoeAxZO3oDIMgALTKZoEv4
hn8ZjDCmkH0j/OaC4S3QGEhH9M2hHo+C9IP8R9TPEhoR+nJEvQuWLhDaYqMSkWcf
64J/GSvBSK0nM0bjs5tI1U/y4ogKZVG3sX3i11ggc4QGXueAg3XwRMUnmypoGRyW
2AuyGVauxaWgBuUn7HRJOMcLz+ZYAvb8SrHBtIMjFPTUkuz+TgemImav7851+1/n
F0zas3s+SI4vyY9+7ed9Eb1VEVMGayPQupriu8R6b3CJHlkkW9OBG5PtZuqOkqQL
IbNP+yIKjCMimLB/Whl+xnN7iV5wBW+FCp7MgtBLayWHxEK35xnRyLmBcFQu9LoI
XAIDlPXupfkY/fr413NxHLdTkN7+9KF/RkjCf1TxPhbRnPGWAErLnWEs+OvNnL4B
/QAHkfrvcBfLejZxuj+34x6zAu7TgHsBnOmS8wyFxORvfbEJexNeFrN2aMypT/fF
Ft21Pi7tj7xxSTAcmQZhWe1wxI6NRjNtEwPhp/LiJncPrkHYl7D5r3PekCOTbo0J
c0LSJdvF/XoozsXYKfsZRaEioh0/pVJAi+WBoVwyrIkPk23w0R7x76pg6P+Z+W9a
9g5oRBXXpuxCC8HHTFqGJqgN1VANblVJrph6uUvCCPK0eVvEOiWslE6vqrJMHjHw
zcLtUdF+CijGSrdyjptrPadBJoJuryMog63mBnxIHA/PZ1XjPEwZ3LTeVZQ0cTef
i0vtGJEVTojanAx+BoCwwGLewIa6rDzg4Lvsf0WW1iFKUz8RvEO4qNmB+gvJ7fIi
rUYW62MmLkxRU0jBd+1ZvCFSZUz1q12221+KDn+QWsRMfXD5zJu09ZaZQs7ajTbM
EirKOPcYLbKS2JOhOZM55FilnUs9JRXnY9cP1B8PKfOxQwdbzn5H5Wces/bft4tx
EUMgpmiifIjPgNyY0Ax8u/Z3KvQId2yZSE0QklKoeo+Bu3U1NlRhpHcoxi3EYvxg
ECwVClugnpdc4e+sHkdnNcO+6lj0qazgwF3sZ1BE9aBg7947nLeM1MEPVC5CfolX
1GzCZzghPyLbj29k7YlGogIRvdj0xqmblJgfdXERHtK68d4hSGo+fsIZwpTCwQaW
IHXRnZjR+SsQsxJHblpmCWMIONJpIJmLPB2hrnjTPvMEjCN2hWKyLgLCisK184em
odxyHy1anQZMYAPGQDz2u0Bnj1pnOXVPSk22tVTQW2HLZsy3P5+/qLsdtFBHvlcm
BA3qbFbyT1p5zAQkzHYSA6VsEEPAGxDDb8rc/0WNkxMZeI8rwzEN4boqlmvRZkHX
YVgDjuaEcdBi0grNPOK+sFfHzlC+33IdT8v8sybi8Qan5M/U7olyKNZ7OvNIqbN6
Vktdk11nlQgQY0hfY5c849XURBk41gkn+sLCTxc4uRgNT2mXV1Tk4qFmEiTPLNIb
F7anGpZnWdEFLphYP6K/G1a6lT/OdNNaBJJxkQ3OcniC1S9LegbBDZFWD/dPn4AL
WisBOMdOOhI/9VeQtMIEJw9fW7EG7QaQhlXnMMUkA1QPY+Icd+YO8yN1obARAHaM
EMsapoNaqlZ1UGopXBBkZ7FA54+C1dZDxuS+ws3bgfr7Xrq00LCceF/bAY27vvAy
LxLdBh7owgr3HPaxWjWldpb1DrX//UOhgraY/0x/lvdzkS05q8feWlsfRPJWUA7j
0moe/bDBE9U0uHowGwkj9IxrE2fbsRJyHcs8LSPvM7ZO9zThXk2Asl5U367mEbQA
O+rHYFSIcVXtkVy4y9tbE0V6fWHc1zMCMIo3zDxSldcC5JCvncNFC5NoNWta+es0
7cnsGYMwCj7LEvfzBjaCzEGENJaKvr2W1p8+11vBGCWzuyld6TsOAvk5PK7eDbRX
whwleMb1EAZYcU6HyqSbKxAU63D/lCHieUGMXS0a55RHUyLEy0lAr2HBLB/sJogs
icKYtbrKru0v8N7ZWDNgNzfVJ+pjkEgyjixJBMlgstAT9xyRd/edGUAcGOFZhZ9V
C76cEKoG0fn8aA0RTOc5jUWN4X+Skt/c0/+IoCSHSKLF02e3yWJpthmuW64T2+Fr
asAOhY1fUtLaEILcSbTDygrJPppk+Nsd6LDWx0OX9VePM0Z8PU1qDlMA//itlZd+
xZrjjdD8K8ZmR9H5Sra6PNoOzPwVMBjAfq7io1PfpNd+BIJySCvdJ+Clls79tKh7
91h+K/4InHmVRiGOy+Gkz1j9+qiZj1yJ5RYqiLSK5ERjdqhEvoQp8cBxaGI2PSpn
eymmXMST0RJg602nRYO70EyzSqTvUE32R5Jrt2N5xPOdot6Um71ZLMVEIJR29ZDD
16ivLZJOu8EzAHYG7ZHtjBwvvrG469n0CwgCUYl1bdFv0Itn2wzkRe3fWkYY3KnC
2qt+pDykGhM7AqzsNhWLfNIXw3Cjbbd8sAAWzJgR3WgFxY5diemXaiVYZ8PtxxuB
qp1RNcvrRCdTvIaoDS4N2NHbDaAXTnfPuwJJn6ElZVoMBgkbarAvcL67Lm9VjH7x
DrsPANDEUMzhoogZUCEUpO7cRS6CAnNF73PF2OlZCLSSevKIriF54kloLdUzNJ/A
AwdSsoUkv8yQ4NEkuI2QkJJorCR5torCBjZ2d+s9VL5rHXsNzO+qtRIYlGMcLnh+
Ns354G4WfaATnOhPQe2nhTU7b5VxNYU+Ca1GL/Lid2q8wADcOLLaVI9uYUOh0se1
1KWKS3QOorWTc669+IQaBrW8doxeoLKYU35SAKTpFUVU5ZSv64KDG2kQ5BHWEVdq
vdVx3Y2YIbZyoBXhFfsAD/X2ned5FY64UwUgkZ5Ghw9LvU9eGfnxVtJHdF/u4zge
pT3FN2a7ieev0IbDqQLH4Wi/k6Ma/FUMM4UAVktnzQgPioxSrApc875AjRlryvzV
oNKRRSVMVc5R1TUzo7YKkCVEz+6/K4p9371Il2BTunYnxozA5Lft8Gu7muLzYsPj
Q0lAKcU+G+rGPhfIofYU6Hk9bgH6arfK28C4A4dcJeTPmx3bEgUQYI1RYTtsgln6
rOX0vJz9ZpE5jFn8bgPMf3mu/XEW2Uu6WYoZg4OC0/Oxb+tejTIv5BIs4nKBuIpJ
LhjiVuOfBeLFV4mXfVI9dd8pa8NSIaIMIfF9B6G3i2I6KFWFMLkr8YUFs37/HmIY
wjUIj6V4mwC+Wq1Zt9JdDWJPyZwTIMq05RIcZdZN810ktJV3qeFmGiGuPGfPAQ+6
9b3qDev5YZCWyUVmfzBuPk7NIKvWgJ6qhU09diKhG/ms4JhWFmf5agFdsbfE5oXJ
OFjDKZ+HX8xk7NTs29p7/OviFRM4UegSjw3lxSQNR18FCekZs+mim2ZrX0s51hLI
Y6EpH8OJovCwslqezGavoHl5vsP08aR9NSOUb7uc5h1xvN+FwkVG5LIxo+dnNMqu
9S1KqpidTGFjtSTgldKgqhAhRsJv2xVIt9uum06bPDD6bH2Cbg+Z0pnxM3FibpPP
GUV3ta/c7neQGU3UqzxgysLWKcwRrKBYmdLrTqbURnV2TlkKpF4zkw4BqC40XgE5
TkTiSTAXBMgx/MqMfNZjzKobIdnRX8GJylPHc3u8k0ZVz6CHq8fKaVaLTX8lEXoU
PM4AffLFGel3uyW+0tvTyt6jbpKVNDQy6jIeNuvkBrkmZ37mXm9XYR+uQXMEOqGo
zSDSnwlTIQBjSW31o6ExVMUj7Ak2Y+ySDI/RGmZ09gxmbWRhxs78fTru3G4wXlLn
F4Xgl6jyI2F4REMQ5NZekRL37IIk7mC9mzZRkpVYi8b6zJvoqBqyLTxbJd93W+1s
q6+MIZ3GvrZSByWpGBzx/5gL5P9jEESXV5Mo9HjN4V4Dp1zY3wISz/lLEPDFcvxM
46xbt5P0cNDGpUUg6VObfoRjcEJ9syizZ9iPPpgoJk0pO0nycPyRsDneffvV/n50
9d2mWU/6EKfh1DZvlytrIk4jvDrAgsdaxV9ENY+yMD74s9Uwv7QHuBHF3HaOBq+h
FxTIow0LspGFda0VSx/djEVZuscEoMsc3CNSCkZ7Vt6wF0VnkIHADVAqvNWAr6BF
7VOU4IcAOtnE3iXlReRf9cE8vY4hLo4Bq3NADSPIjCCBnmudIYCSZXd037eR4OIT
WQ987XJ1FHoe0tR3sHZHNcqq/f/0GzT7BfqDCHN6SX5akbVtJ7soNku1ZB+5so1e
xOh02PZqsGxpUPtJ8ACGVi4iM/+YMcqXqskxNDIAIXEekSIkRL2qQkF2U/KN47wf
G17m22bRLtgDYFw5Q9JTZ05u57esYI3fVNqTtoHObWw2idw7EEIHzCN2mDTmRXkE
z7t0gF64EOlk2ofkb7EpWYe9KDkstdYC4xWNUtuZ0kULXnSLV7rjJS8zGt+CZp9x
+z8p//vZWgxfpI8SZL68C6He/wSkFAxCh+cd5buq++x4T6MoUTEil+YdBUSN6wSB
g8BVIJkPsyqQDfIIVKIMfohlMDcRCrHJJEW7wcGW0db5oHN2QtqYp0ryLpBZWZth
0BDE3dGBg8sw8FLJz/p6dI2C885QPiLTSKUBKyKCfW8CAAAzHy3+VqmYEBNQ35Fs
+xw3h9REBaq5884jeqbj8/xbs8mAYQcqgqMVlFcKe4W8lt6dRxzDRnahESo7PubK
/1+l7TToWCnBmM1Nq4wcZUWt10+ZnFSW5fODVJON8oOZ7l2VKRy4+6lO94sRz/9i
m1bN7Iqt8GmjJbbKGJ2S5ID+NBYJy6iHQ4UMI7FSlbYO5eMSclGBmKvOo5ZMv7F4
akt8y3LCeCytJ+mhgCtp8qyiSEEwldAuncSZBms7KZRuLUKQ9EyDQSkXjs4a7hG9
RWDjxp7QKg/bpf4lodki4EI/vjRUu6oYmiL1Sa3q0D4zNmA/IcHGhPeDcD9QvabS
sxRYDCdnGQB+aHQqyAbptLxBW34KGRoBQRO4cgZyoCByxdlF/1ob8GvOHXVG0oF7
k4VCV1jM7engwjqALKGRQWI758vHgSVEiI9TnV4pCB7ttleulzQFt6kZcpgG+Fb3
lLt0nYZylcg4Qf+jovPi28AfEuFzDXBAH4e0cfnhPKHjGKFJdXPZ5dfwgFRMZqr8
qnm8o2ETQ7EGICZypJ5eXdxPMziz4heHrU3gg/ef5UtYfcGBMKOAMLQmXte/I/Lk
oq8ZvB7i2HPqs1geeEM2iAwmpUqSH8ZJga1e0S1/dXkhb0r1BaYj/g5atzrvm/t7
A/cqHPVBrotpbZFruocFZMtQBpWfqnWc0be4Ze6fnYVY6eUx1DhxOUE2iHxaYo/C
I3XhFZKH+uJP+cKfvQeAuj2acp8q7DvjdwegIqbNY3tCVAb5WFDIYO1u3LAfeFVC
wUo6bjBtvfUnsdzcel1FfKUrtgJbRQcGB9vxwxw+UtWR/s1i6WOYGVxydsBO9hem
iWSXMhox1KVKNP8kXJFDhzYayYeO1U7tTqz2hYHFWZvZ8vXp9sdF9VW6kpYDbiTH
2s8GUYjVMhYJWNXsbcgnzXK5EbY8xF0vNmasm20Z59JIsHPCYsa0OBNoQEo8/cII
z/KtezFRzld6ajg7DiwTUtzRMS3Yq75vr8Nyer1wXx58MiVi3EMa4lAEH5Ga478S
0IvNfEpGQlRh//7RjB8x1JnlV53NsaRoRIDyLzKuGa007kDJvbzXg9+SqbOvL/vC
qls1e18FQv6dl3oj4OBlkJVcXFh+tszLutMxRxXEFDBhzzkFBdD4B80zc5bHhXzt
wh6EV5QQXl7BM9m3R2NgDq/qGKf4PXgoHoW8uBUkIKm5VtTdmobwDQYoxlJ3M3af
mIyqJTSsXuugbMqYWNxagWEqcE2eUpY+4eabXHO+/IJp543A3s6+B7KfqmvXL2wt
hAqZNxut/7FRam7wx94uB7mNjv/LhLt+QWacjXYqg1fMpTjxbyzIKWVck0+hUxP1
PZgEkf6/dPG9oT6vTauXvnjCWEU7+uCH2lLJwfj7WCKBQW0d060f2kdPeWSdx5ZF
cimaqcBeF8JcYSAw7OgAQkZcNZzE8yVs+BCPivmjA5l55TK+WGVdp14A3bHjN+2N
+8DtInUFzwPA6cQY1AhC0HFr81DXDevFgLqVp4rcvU151B2jhOQ9st1MaUyc2Qjt
4OeLWlOj7T2MMSv0KgAWYoq4sOi6bgHnhPrKABctyuYKJ87QzgU1n04xVovTQQML
DMwzEzMBl+aBqAA5CmuXXQj84hOnYCXk1STJQ63FBzJgPjEOminr51wDZfuzoOWW
/P7x4m5OnCs8eq1jZr6IErdeO4FsGuuB3nfe241+zOqJ/Ul/cWn/KC4eW3sfsjCM
mnoWc58nICIRO/MNZkowOe8bbomy3E52U3JUK1GDr53bWHltivn+zGhJI24k2H/O
PA7zQMr5g4HwFpx7RmQdGgZH7hdxNbP8LezTPAnBc+C0qhPJAEDpggtP/70/nOCk
3xFLVOH71soeMNYc9jgCW9M7hmAwHCqf1kEBU5IHYkurbebCYdEzkXKUkzk67ZlR
EdCH75qIfJpeq29G8DrcmVH9Z/t13JLuErR5ifg9EAi11WIcn0cGF/DsQ2d23aPM
WQtPvccl4TU23ed4GYmsZ/YoeAZ06UBf5xeaPMhvKv2pqU3QhGwu49o2VtrhDcty
W+sPZrsBseKuAzkvf0DeYxzHYL8JoPsr9+C7h0dRpnEFsOSdWk32tja9mTp1/JRo
K2kTX2GjvRs5kUFpBznGWZSdsn5NNkmmpA/r3nqTTGzg2OMu8HWfuZkpRUbsqyTu
s88vzo7FIksbAh0v3G6rYw6GSRsk9Pij5a800X3Xqkktimi78u2OFiHhIqrAJzHn
Q5tJ59iLJvIlfGPBDiTwbNlYdD9EzpHMwW9TAhxq28QDVC2ShDGAiLJst4dBRsP1
BqffEYGUl6Pm8ViC8Dgn8S5qIKtGX9zs6KiEZi1lVpCKs2RGQI0/IB50tl8Vxfhb
sjOJepUt6EeOgQK3Xiu3QFt8lkyJbHXiBDVj7XMQ/RpTf8n3VZlaho0OGvhS6Pxj
xkfpNTIkBYdjpGUNn3vpU7T7T54bsnlQbzgUG4xChsiP3eXsPRKMpmKiHdGctA/c
9TiALCjOIheX/D21KZHVTsokWfQ9ujXb9OD7dP8QPpA6Bp83T8HqPphPEXfB/zzt
NwW6OZ4bQd68q21bgUXxT2qhvGufccNTfEQHLK+hgXgESi711ZUiLJn3ctdR+8FU
hNsVZCi7f3Hjz9znUdbjPs17M3W/VZDmXlW7FqQudTB8c+aW8jA+Ifqh3e8df8vZ
SLKzFbsHOCEy2VcMxS/4fcI9TIs4DzYGORkWStv4CgQHMjEiwIdQUvOLkHHq8WHR
j7IqyUzVlzoPVzW0gUhYff1hFfAPDnirjqZNjNyksf5cy1ifWzokk++Tns4d8MU/
jwKIqnImM+BITl7HjKnA8ODv235ezmwQe+GaoBfTgUL067kntsfHP6C+VOIs+oWS
981MLBbwWKExf8SpeYj1aS57aALfVhKGSJHmEFCMJiUHp0LMO1Sba6Ai9holv90/
OJ0mdzJeCKwoeo9NxHytw61N2y2T18kZlXy+gkk6AqNZQ4ou1Y6ltmbJIWcTEoZn
YNdHBoNBO+7+349u8bG3GzK5t04QRLP4aTd5M2Vd3Ns5j0PGNrlfoDnteKhAucj+
SraRtCD0buu1bTbcQ/zwVWljP2BLe0eR4vB78RH5fuyIvI2/h+EmK5z+YqwI+5ni
XBq532HUmCJpz5ncyUkpYnREAFWqYhDjO05QnguYJD4v85S/Ee6AOHZqilKSWK+R
E6EkL4/k/1t0NRNnAmUY7VYASLms+MkOgh8aOAVR1mMP/cmJdLuQor+4IA7mF73O
nbxdx0G8gRjBcxGnDUAI1EU6/4hd4KnyZ6gmyANblX9r2xVm1fvTV9M7uX/wfEy1
FmxB+F/da8zno/1kOlvVIwrBpk6HS09yd98egE4JL//Y5w/m3sMuV+kviQKBG4Gs
XZ2RatYeevl0qBGnDf23ngYX4FLyIEfNqcM2bMz3MIdjwKReiu3F8nqcs1KeFNOI
7LKrmai5vuLYKD0fLOIjdImvlK1ugHTm090PGz9ro/9lCgNRUdhMevWyY85SbaCo
WiFT+I/G7lkFAiK0b7azbaECs198r/q3J8gn+tfiTFeFKxyRVDOf5rGOwZygZe+a
heus8DZcDRaUZ4zW9ndR2JK6HwtlfFxnxvFfQ2C3H/huI9s2yXbDXh/IS+ScPTzi
GC7xM4b+gtu90uDkS1QO+IJQ9KU93KiLYk000UuGEELL2WT3KMvV1kzQpOA8NFz3
uTUJLAwC7GON3RBR2jZEraTEY/hF4N9jKhtGIJnn8XaQ4NRp98OOnAQu7Z+FKpLY
5SD1ZnzcYy2Qfa2cM1qkjIdqQEtt4E8oVpAB32YjBdRqWlaJspEW3NAecI0dfWho
eQMI6008xMpi5ZW3MqR8jx4ye8tPSaoeU6fL8JGBBWKmjX4QotSHuwA5YfPlKtui
pvqWFpGrNMwKysPjJ39D+MxFr81aMUKKXmCqneUOntCLzxI4417WXymWRLUh8+3z
ab+fQZqMPjisklS6UXzwhHzrhIf357vz87wHfztqINh/c6LMb91TYM3BkZaQVyww
hMTxhzSbTI+mpYtryAWqjwdYhlqPPD5oXag+gKcfyDr9nYzYsokCdf9OfiAec85T
oc1v1lyE9VjPHMMwF41z+wh60kzC+T6BvLTGaXaEmm+fEdIYt6V+F9ayTi7ugtAn
gwCNdjBA/RLoe0Lr8MDq739xOnqg6dSojVFwX59E4rysK3+NmgiJbl/R1vRlIuA/
cM+3ye1cHeJBPmaEL5F3FU5aACeXFxf1FWzPifYoO+L47c7jxJ3smclIc5omhLh5
ZTQX3ZF2ongYCmoK24Inr8Wlj4E6ZKPPdzyj1MpzVRJg/AG8YXSv5qfBG3rrcPl+
5dBkCNYzg1qrDr7yUL9Z1pDjumq5Pcsrm3p18ohOVbFKsoZHu6KPdQDB3oyj7glK
mgH47dVFFDOuN6+lJkmIrRmydokr0yOz2Gf0S9/gJGWD5WhDp6SOnqYFmgysRHAS
WA/9IDOuuDGiEFtDeL0VXhEzwjy9pPNGriXQaht78vYcNUx54okiQCMT0UQAe+nO
ioGnL8vVNTOQkk22zgdDvohvNAUwgI9bN1yUZP63lgrQ9VbkqBLzWfmkCtsMz0Gi
EmR4s0omq43FgWQa7GKRkRIjsgZj/G0CiJjiQINxe4x283x04jbpPJKz87HC36oT
DcuM0FRrraCJ8P/Z2lwt9vOSm7P+YsmLJh/cHReD7pBeNkjdHg9Kh7bp4ZWibhzm
KqxYQJDXkKG4sJJOoAeWr2lDfk927T/+u51+mRlLi9x15+FW7DXhRkRbwjKNdSjG
vUtRdY45XCKg889AUsIoHo8h/QE7vmxt2cYYbSKWxdXUEOYURM1vLQxW+x3Mn0nF
vJTO03boXtlMCGrXV86Lc7vzGs2/uzuHIrJmA47+2c0kJPP0CvsfAT45CLJVYJAK
JUJHHqkv3xjUwpasAQiAvD6g1d+vzVELit6n3Ox2lMsCFljNjZgdfH2on7wjqoPo
z0rbEMffwJYVtzFGfzo6FgFniaNAfdUW73X0jJgxHtvKs0v7H95A5DfpBD4Pq62b
P6UFrWD2d2vgdE3o9w7u9OlnDQepcbqHDUZaTH0ddXwsixSAe8vTbe4Lq31xYVFd
lSJUDcqgeyRdQk+zSKmwD4G8G3ZEi8BXbLOb620c5tboXyOTWaN+gMLZJGRykgGJ
wd/lWBxsFvpXugcgZuKRmyc8LXXZJeJ6ITeS2Pde0M4plNNZXq8qVJUd/Qa8ould
A+hU0qpCPYW42zkvERcxttPuOj2bJTjqQsgKol0Ik/1XoTD0JtoSFh4cW/paXEez
F+cNKIdX1Shnh9ok3ZYFyhELlji9u4HqPYv8GFWUcRbXFA5C6ahNHadWvQrmpln2
Z2cAofsEevdGGgDr9hZQGOaJ9s7UKYWCOzvA2Cav/XXr1AvHveOChSzkCpoOpCw2
ir6TpMHmbMTV6ZycqCotGZ187uK3LHJ3TSDjzkERtepnHeTSYlaPdktLfm143Mkv
lpePMS2SmmKKGmAze8A/RTd6B8IeDppKSo0IhzJwY5ATzu8Xn2m37BkdbfYSxGso
PnfW6yJcIP2UbVdRghi/vD+Bmf5rz4tuqGhOl4e/+L+QSi59tkMT6l3RJTLeWHKp
Vw1+D9lNVyfkZX/8d1J9kkhoioFqWcOX5xi7W7gzywqU/4RHUgv/3w0asaoIQlWs
L1hPNuTgeTBQ35tjjH65i1/kIvXzp+9T2CqzwLbxlIwspT6YqceCAwnbM/oVT1pF
3DMK93oTTQ4Qc2CIhcmgy8SIsL2PNutmItYexZJiHSjrTwgpkXbxAJDrNgfKXKN2
WlJ5236YPJ4naJGzJiPKLvqHiMZUwGl/RMS5YX6MR70xoRq0c8cFq32/Bz547AYC
ak90FaP+1EbZkubxVMtKgPXVZTankpi+CN3gJz31DdRZ6rN2owulBzMppWprP3Un
MNj6QUnLJW3YEygEWnRWfZmfHF5TAS8uJpaxFqcP3VIquWo5tz/fVx0fYVinwjgb
dPE5jxjAmG0YPz0gjkW6LlyeAIcZEAbzmJ6AJXlcPi/+0xNzyIVQRO9jIPxCGZtF
pIeVM6maRsyDaocZgv1NHWxUzxfuJQbPpFiTNeKyA49ofJbsBN92/dVJ/FtzB/Ow
1c2J1PJef1Sah3IKcFL+Dc2klxeST01Tvx49J4pFpXh3bf76hJnuo9ucui49wH+T
tCUO0lqAOluDwOcmMGnWpZZxsu3MFQJzmxFTecXWB1QQjA3eFdBhrS4HX0bJwipH
Hw4rvtSFgRTU2kCt2pfUx53ZGhIg+7UIbc+wkqaVJ2Vdi/BOlth07liTQ/eLJuSc
uhmKYzi7ZyYjNiLaP4WlS8Bu4DgGjEIZjaPh125YPEdWlpbR4ViqGmPpsjUWNSpU
WHy4LJE1au23oIrY1u4csH2HRpx4yX60oLP5Oa4bYtD2NXODfb0XqGF2+CKdWpqL
mukY08QYRmOecz6aJnp4AV4oE0jlY2Y9iQWkzozIpNbAHS1b6E0KL0XZ6hkU1AJ1
QA03IzsNpdqwVoPhuTez6arr0P3XB4c138Y70sm9q7d2gpYhpD7wa3T+GUgGqqax
Q+ucRQQnwi8aVnXGlbcm257vNiMHvQ+jk/7g10vl93Oc22T8W1b7FIqbwVKqO81q
8pKTHyUqiMRdToZiFMEabQlQFfP0Lscbn40ReEl5l/IC19uZu10/Lsk9j/KWgAmj
mREaaJlGY5EcT3W+/arxp5QAGe0fBovxI3CeFG4tGwpG2DSUq4qOoy2aMp9/iq9C
MmFGTL3m6oqusYVpZFXn0HFTJAi8+3GO8oN/meEN4MBO79VCC8yZg/0oqW8xVHLk
eguZ/Gvp4BmWHvzJ4n9zCPvwId7sw3vIz4mqYrt1wdMRlINsmr8kBeYanFhjm7EO
36MFuLKfikpnfPrpiTTlZDYi2AZScKFVM5IplvPKmHuKj6uFN6WpB/xMImDGFDJ8
XRTJpxhdR3VZu7iEx18ufg3GoCpUECLuw4+4XCSOHzCdb1Xi8LfCmHfS4QqREpjN
EJtj090OGVjoAXkeShHi04uzM8nt2mdb9ILAeYzTI2HQ4c9NGB43wOU6OkegYK+w
fIZrNbxkHS1LG8GQWLvJpZB3SMh6eRBDDe38g4Z7hVrxsxiuIlxD85P0rSGTrc9k
CcOoeHNIS92GI97mJ8L9gPOMa4T5ak6cM1Wf7kL/QZU44FtqUuPo9ELwLXO1UvYr
YAwO4jibcc/A5NKQ1zmrbjTY0hTEKhwtsptjrusS1khEEx7FsyculMul50YYnACY
jhZjJLRcMCr0Jy72Zg6OGChwTQxBVKvrp4JiHaZA8ng2VNc0jvep9WK5jxFOqmH7
7P28MS3o1QLzav+sGvAtAsUB5TiV3YwQDHKTtNyuk53Bd2iVkz3IOS8Ahp3Ufhvg
d1ZwP21fRqS1KF4cnRshTxNVaygidi2jHGwIHp1EA9orP5MerJVxOIpWk8Uqqt0E
plrRUpFAlIhhJ9wlihSBn+4FjZIzm0JmnGQfr/nfsvfXju85KNTI4yGFQWbIBfxB
0X8k5tvWok5wj7tiDHIforSZh+B0d1Scz2yLqF7YWx9FkThiGEffkInWv1s75/TE
32EsCIr4ySwKBChMjQpb96r2VkFt83oHHUUerxK3pd1+28qbgI6E7IhH7dxcGWY0
WOoAIKQn0oetEvefkdTE4M3i5uXxiOTJxnwfPTWLE/swWI24fLxK4FVrHgaYD9/J
IxvlEXloykW9ikjNPIxOvmldFmg/WyXXiG4KmdD0a/TjFZ7WOh68u5Zz1/y8X8if
BehNEXAROHQ6cjDK9v759S6UP4eyqy8lMbmEXOSAMn0qVJL/pG2Qx+dV9bFDLlgV
mZ17OCwXJh08bnzKuE0hGpgkTo+FJLk9o/p7Nd4m4Zcv+yqaV+NtkwVxpEd1HH+v
ACHwzvxLWLcJ7c28sAILt58D9hO87+aRHgk9eOxQjAXE35AC7IIhuo6JYp+AZuN5
Fh3PMREDfmlCgOwgSnSdEs5MeegDgLbF0B8xdXxw3pEyjCkauLBPW6ZWdSfgYaff
dH0t3hbLD+R7erZtYza9tL1/qBv9Dz6FidXFzERqqJR8DRI+HGblH+t1L/IiSbjn
bek42YvKlqRt7GMkMz1W8QOVsVAfiaDgTdEOy0g+khI71XQr7lBYCsaSUpFb53cc
9LQ5PgTOj9wgAYMkHHGGTBqtYjQAXFQ1l9RZOofU8L87+BVxQe8ufaNZoqAscXa6
bTR1d3nlp+D2Gp1plGw6mZr/+/BVHGVNWy9Wx/ovoXezFdgCcpLkVpLqmp4Wpz3q
e0vSZPUjDMlGTihZXz3st9NYieI6r1lqEloyNHsatvv2QMgaVqJltcbUOPlL4frl
kK9Tia5ZGHu+o3EmUtrdJ51dH3iWTLC/ZX7oEzvRg13lqYqnhH9zJfG+/p5cf0I/
LGI0ylljSqgOYbh50FvPSv/8BtkWBSzeY0KRH5YAh5nZSdL1bjlDKEGcQ3oyginO
s0+Gue26AzzYoa+hqR1fA/+Mr8uYwi8Byyo+E4rjaCquDjSGBfC5Za5BHoNlNcvG
bnBBRKfhv0g3UmIGAqVPsrWYs1JAhRKhX0NCHscyCP7CH7f/umj9K9Mb2IPbG6sl
a4vDBF1NpYYll5eZc45PY1MWE6DQsa9DQ9dgmWToVuPPc0NFHokH1cyrr96VXulX
mZf3UWaTQnJdTrmwePZTZxP1qF04JlgEg6njUzoIIIsXatnwNhc5nF5FtKM4AB6s
nJbcIoe1nwHlaj/LUUkkSubjicG/D3GKwR6JRqD7ZYWyXxA7j6ZbZwRQnKPpFsgE
ieirnF/Oa/OfbPrn0lZoxRTwtp0oZidoyaPVyReiCY3Zo9KJzG0KZGVRNti9HWP+
H3iOSA3Xd8KPyn19OyKWELgStn+VKSqxiwObiSWvTICZyh0ORhCA+CoEHJ7KuaVg
kNwee50cDVjeutTHLGMNoW6mILnqkyS+JRF4vWLWDw72wTlcCNhv18l+60X8awpT
CTbyKaP3F2Vb3mcmG3zmR5MuibgQhH5jCRX5pSwhwTDAD1Iq+8IfuumXo14T4pdy
WPESzKXI0v7EarwZj4VTlHqWmiXwe+HNuqEtuMw+Dts4Rdued2mD5JG9voj2SIBG
iaE0bDK3dmM7IYY4nWEib8PlBLJahcyxE6Mwd1Lcalt65HET7n6id7LZvI3rfrDD
1OcqsLoMGnE5NR0KKqeO3FQO21pwY0ITMM/rAOG9hGNo74dURlXcUzqrZrwTknLG
EzBBWmR9x96w+n4uemrdQoodabDMnl16yvSeZDu4gLoM13Zy8ov6AuAYBUQblIF8
61jWyT/bsseryyyl/iOXBRKyKCYX+493HO8zAtUCVJXIQLM7ECsRLbhZz05BAe2a
Y4VtgDEE33/+JEuIm0R9j0ppT8yTI+fvGiCzhX/cICTSeLs3vfxIpaL3omOHYhUW
a55qqN7EBWihpku7yMQSCKsWiX431FW/+9eyynXnDQDT7jHKVIKeg6+F2n9SKs3r
JOOEJyk76BLjrIuWYS79SP/ftxMUvUekyPBBD3R+Z6GAkI8bDLJK0Sze6R5G4WN0
KwzfAIijwlipE9xfzN6cATsFA+ahVd7HxSX5zPWjtfPxakO9YDWDMYAXeUG9X7ob
AQ2kg9mc+2J40FkZcY0TE+WWw2lyZlHcUK3x6NM9N+YOb29xh0pKRPx+6qHadwlh
inU+gvodQumn6s4lQNxtbHxKtgK1+GUbZsdHPKWOvfedqil1f1YxL7lTk8lNKq6n
iBFf9S+ZsS+DG1qPitNh9Gwk1MmxBEL0UrFUpPKxBUL65VaFGaQdN+aOO9UIC9pS
KwTb/f4+L3VPJHXZE7XBe4IDZLaiNAWiuxotPljQmBfeipZJZIh7djg4gT9U6e8g
/ASxieNWIUkzSr9Y0p32J5jjWQFaTsz5Tbsin1NlXepmtkmdHcrZ0OFGOos2XckT
PPrC026jaCL56gl61R36h9SbUmiLGSbFPVOlMwss18XHtYFNHD7wTWOSV9uqyRml
FjZBnyE253XT6dv1KKl1IyYOtG7fp8QVMjt8UOFPJ8oGFRZ1/ClO/sqmXjRw5h8j
W82BqQWaFKPEurGRreU7IAbDr0X+cEtoh45Luug/wgJl8xABeinFot1CpNhEmRAz
xGagg9tEQtIK1B4mE9RkrZuTd0n5me/r63opIkDCh3SNVD+Vv47vijjr3zzvXfGu
c3gircvZA5QThkD15aFLLor7CQd1UxDpS8QGTPU1gQP4MuuoCBlYykiCtjZOJS4m
0AZ6teAr0yoAu9kHr2RnD/FHyQA+QjKpz8L4zhxkvlVY7GANkbVRqNMPoSjTyvRd
2dcJE83LHPV/UMHZqYf9sFpJQC3bbIBCdt+c2w0UKHRXZoNIfdzYT0a+YB2IwDge
h75R67E6guh2cClf2eOw/F+ZuYny3J+0eUyG6YTbv+l+vXMPCS+3LmZbiwUSy5+r
kWbvaG+J/ddSdOAD1qMSJMZF8+l1BVDzOGTfBXW0OUO4KDaxgOSL0RZXznHvYa4B
2ABPQ8Z47VQCsp3/m5a3FE1z4UzICSCZQZ9lmbOWG9RwDU0KG3nUCW/TZ8AEafzb
m8uycbvBXlwBy/LXTdEmRY2IuqAHtBxZzv9rPSZHVxiD9FGy2f4Gddq4CiXQl7IG
gaE6awJqUgRzyUQQgKKdIsAbWFA/xpnA0PiyhIXpINoyDIa5MMMz0tyrlr4irrJo
AXID5TQ39OxRxv4gqhMlo2X3TaDlwKfsGdZk8k6xCBHCqZKLDubOkpTWsTSTwWL+
THjy2VZCuGgDh8YYUHng6qcwefY7k0RNMZeCrwiDNJn58Xt/1iSnSZWgTigj0DV0
17YBcPuWOxHWadsdGU37nOJNeWls9cF5x+204Yk0tfKuah8e4p0M5vGUQi+waFXs
wuva7BZRPwpD20fIAlIT5hO694Al6J7IK2uKuwg/sMyVNQ5boS47sS49n5DCHSdx
uk52R/Oz9dA05jqMOz2uwj+9+rj2ewi+YOj2QIFpqLuwLjGUyB416ZTlZtDPlMeQ
ZbTmLo2lXj4SJTKiswQpkyqPT6QGqwy080sLYIy+nr6BrHY8Z8xL/qYvawjDzfyD
xSMzcwS3CR10Q0iE5U5wL2lLng4BHMBVwNBdZCgELUGRfni4le2AAFhAKZkH03yy
TQ/3JSCsfmoiEnwsXoV4dI2z6pRwREVxtAVZeNVbkPMlAUDXTbw25deHAn5g5bkv
11sdweNZFiTsfGpUR0C/xvhJqRzqQ3Gtw1mXg39RNsIcEFjiIoWAVIewnjDpTZNX
YCshaS2h6dAvmE1Ie7KUNQo9cglWuJBMLaOzWUeTwHw0g1LI4TQ05G0BR3cS7FWT
ZbqqmhhDGJpvVd+pp8uKdRI558gca+jiIg3hFPwYNmVK4juWSqTH42LJtWq+lDlo
qJxtGWDuvtCpQJe0JdbPWT+jYYi62YXHWTLnt2UxL/PRAht9Up/+7lFLl5uHZtmw
xV+1cfStbDctnt2/VlHijQrc/xl8LFrcYKwK2oswT/z3pOF3uqYU2xjAZR2Jfey8
YZdGB4JKAQf0d12/Xs8mLD5c82Rsx+dE8G0hIeN1JilIoRNjN3uHNfTGaKsMQ+DE
tXjqDj6nzGkVpGFaDdK8tsVUzgGYXYW2U6NNxFh3OBKPGehzzW3e+HOF0xbzcJFs
quW9iDvH7ARKZONf7lnPnHbsv+qOaIlzW8GLvnJ/ezuyneVLr9iv8oXfzir5jTVk
he5r/0qX1VM8G9TP249AHu/pu/7TYjC/1CSiH2k/ilBxAhaI1S8+9MWU6aJ/Nx2N
fbsnLjv0thPT5HThQCv9DwdWFpQEVl4aXG8aUWDBaYOjVn1jtQbBczKJAd8sl++j
QV7YAw8HU5VTIxAnGhJsvvttKIBdGcpJop43B2uyb7jp8/EwXte4TovO13VAmueW
3fofMd/StC6YwnESquAGeBE0opr7CBY0+m5T7Cf9VmAe2A/jRRddGsMRd34CD0OO
ha1wkQD/Vjkx6WIdErMtM63UHiS+fjTbDsT760TzMowXVn1jTzXJHzlynw6JoOsI
oi5fApbSWVu/j0WiIP9ADRIAzHe4r0xGETORBSHs74+mZDk2et3ygF0lixJ15Vp0
fADLiNq1wnpoPklAkOn8b5IEn8pFe9UdLTynqvDAaeYZNSWa98lJb7QOIy68Q+WS
foOI90jDH2stOB3i9YCxBcOD7uUiOUlLPZ2Oz3EcCZ819lozo+1u3Rs5bBrBqYE/
JcaTSs1mX5/MY1WLV2l2Aa235BdsIvCW41KLdZ6TYoFozWgWADANc9lvQL8Jgv9f
q9ovSN2LP3KHOOW6h7cOtEuCxTKeAYH3jSRcLLyYpUVLPtgI8+ddSTm7p4m/ahP0
d600rXpENbTJR5kLzwi51JFrhG8hzI06m+yg6zLDOmfn1W7rN8ZaSJ9AX+2r91jG
H/T8qruiaK7MAgfW1yI0cH+byCMbvppLi/wKZj0Sr8aCCgoaiVmUEZFuKU2uLbFo
4LA3QQUs76KBK6SSK3BUfs+W14HGqkMoio+npeXsfv3E32yC1g46O0Thj0DsWndV
yq17jydLLhtaLQdB17guHwED9fiZ0KpXbUCpj5cbnEuubj7K1BBIHmJS4xbWP6jY
FkkcqS/28yBqarj3rE4Riads6D/coUfFTymRLIVvTYut5lD188frqOI72aU1uh8U
8G7Al+aHE5aTcpvMOC6E2U+i+4/I5M/I2Svf1GMGank3ADv7KR6MDI2JWvXG7WRO
kgOfWIeZ79OeRQljNrfB9eiAngeRqaR1zgz1c/uBYRPxWvt3gumSAVKpyM3f1Xf5
7+4BdMuvw5kDpEFtjYWeGhwLjyvKC9FaRILAhKc3u64bArRoOXZ1udmmHTehvZY1
NCm4ZwQegCymMbMAEBFAiflGy321KTdxANm3pkzP1g9/jt/kaPvnNEq2eCRry+5o
RHqDBcLPibnbgXaHzZh3DAaT3eqJ0OKtO7L8R/wUA9Oj/8pXHQMAiKnN7dlYkDkQ
Msfot6nmTVqD3cMUNftWW59ELQQpFgdKs7w8IET4nzaFlVp9RUf1GAu9KJD8LZqj
4VAJc8r4mWxp+odXPoAmMPyqN1ccknEOGfCsxZyn85/4M8ViEIM1rN6p9GFJy7/+
OgvO5oT5TA5kfFmM8QjVzuPBVZCRn1+5QVplmEXPRZ+XjxBhKudfA0zSNByiNIbu
/VhTt5WTWE32+6O/9TkoL3fzXYbmM5VqiaBFN1IAlfm8UOF5wLwWJz/zmecp93Wd
D8d3j2nmDCqfGC9BCpPgvewJyVoV2TwwYZH1yrKIC/N4uBcbxTbcaa6sMhtFwZzP
26r68UDmDEhbGxnCFGdzeGSwnUiwRuLx9OuSVvOpnrMNr3ceOpBvvDPDxwSWw5oi
Dxca/cnqFBqyKmYPf7NTSDBff+3Xc0KOT4KAbhOjQ4nQPcVJCk/jDUqSUn9AoKir
kFPODSHt7/+4aDbEntM3QO39Xo+FImjjqAvulq/T9MSaAvy84n/01rnxqAIPYXoO
XMifrYG2hNd8EdY7JSsuqmkCDlGex49C2jIdnIHajJFus9k0l4hWuqmRvPg2NXZn
YgyDEJ+Ljyk2ijzgGk0fShcfRhOuhWh3aJWyKDm1clrwPC+mfjXQwB+j+hrNaDqT
sm7OfHWadctNXAPYc1x00qIdrt6GC0t+wDxQaVElHkq4HDSo2kpOQHu8I4NP2F+N
mzv3Wg761aNtpY24Lnx9+T8oJkM0psMVIKnjBVgYkU4tkPlUHxvBnsisGgAuj/TB
HJ2+yvKkHDehQanfx1bQPSWWtA+sTdemQ1CJSmbUJL+fOB3NVKd5Ra/wK52k1peu
M1J5lL+kl4rXRXtcRtrDFqe6wJoxhI5wjffBCgM51j8ouV/XFvR6jpHuYXyPeMH5
MX+OTaMmrXSNz2+yLDAs7tx3oi1ngBYf1ALZXdYFFoE+kaLEVC3qrtdXjA/E2VZu
+bwalsL9W7lkrtI7uj1lFX/1ksUfeT6JQhCfztpSKMWlVR6lMxv/EFAI+7rx4/4O
u2Umzt5CsDVmidJqvt0p6jiehZBJUeNrnLXDfHwo4Ff94d6MhY2ARCedOWk3ObKi
6S2I/sEiXL6qqF91RQ0vrp7wpB67mqmp5bXeFHaP5dATWiHh8+CEfKG1f/vThlyj
QkU85ZKnby8lHSAbP85JJiVeUIE6ck4VnoUAV3nDr9g8uG1iXBZeX6F4PMj8FzU8
zupn8+o+7dpysOOu7kKjLFfV7miwud+xlT2LuYC/mPElrdLEH9qtlHUsfEIcH4it
EGJGzVjAa96IWewpZPH2Jlzo+q5JXBvUO0qwWdlqMqPWKPq1rzSJhVNCIadLCS7A
XMgLq+98sLNm7DZrasLIPb/20U6vFpBTVJOzvLNE4dFMnaproswk5e2d2ltGSQsj
aAanfF09xHX/xq3fAkdVmEJQt28jIwwiObRcSaIFIFo9eDl9G64s2yicvOSWKJGX
4PLzaIY+/r6HDhi9AZPktwj+jnLaTdh+VmX3hojhP0Jzf69659NFP9rQBaHKsg3p
awtxpzt2eM+2k4f/YdHjFk4cI0UTrvY8Ko0jfr1FoPIYKd1qVXXGfp4HGZz/cmwB
1QLEFXOOb17a/0fUsY4CVvLcmw9p0Hv1g0my9x0iFmtU8b53CDT7LRjE9md3VPYL
E1DXs8p3RB4nR/mqJTDISZJAOr5DIJ6Qh5DGcr3sKO8+4P+LAcVMAoKqnaTAiRXM
XtI2IVWSgG9vtvMdxLt5UagRfhhj6oJAmkn2AQ0V36dpF/coUQX2rx5PzdQBxgU0
z6w7L61GMvi1mGkDKnJmGd2nOsUrcD3a38GaggBovFOAkyXvaGYfnxs1rHlCAb6Y
soKtubFK58/2dR+beb0CKo6Vc6e8mPCCr8LWRlEqaXpR5+SpNO67/WxiZxf3syUa
YkYfrxfIZYY5CDyKjy6JNBFU0i4BXy49iVCwjxKG0bIjlplzl3+fCF1o8ROijYz6
TKCpLB5r1c2pffsPAwSRHEQcjG6XMAvKx/FoTHlWuZVYOwk2ai/xnPDL7RD65LMO
hJOLIlCNVJZU+KiV9P1IU8J83Ex/4dbzINOpxLQluKivIlUHBMFL3wvWKIFfK3za
xlsC1VkaTyhuf9qcKsDy4tGCOb7J8OAK797oIQ9Re64IS2GlDiSWKnjPyYVzGjI3
Z696a/EF2k+ZqeqUvUbnYK1dnhYWYZdPA2t4l9BDJNIynw1o7O2OyUJl/+N5vsQd
rtjLb/JryH7K6/PL6e1YtyHhENHLMmfb7gmjcW9qgoloq7AK4Rp0kq9q2/zY5TPv
ZMvhgG9YXdkU6Bsf19mBBkAzV3SvB3FxWPpsK7HU58z96WMivTdjhv1zoNsa3Qau
rI4RzV9I9awEBzfWMIeyNhJzQh5EgdSobArhLIKfBfjysjMEM2Bsur4Mejy6c2DP
9GYHkHraYT7dYbkC9oRiB+m9+uknQSLewQI+xseIl+0tN+X2tRj6lqINts8LUxxU
6ni1KINBANc5qGOkjWNmdDB8Cm/n+M64g3B8NSr0u/T1gs6tJk8Hk6g4JCMVKQ71
yRhkIwR+9BGyUI1tuhgKdln3DcmskDzEXDHy0fZo8a6mOnZ6Z6J9nDMk+6BmzDIE
REuCtOTPphQDtCcQsdV00zechZAPxwE8M2U60duNRKjGYBNSIYPLIa6BnUFDHZVc
U1u9NmjOykpZpXSoqwS088QTpMLbfxmUzjTl9NnsCvlHJoQOmjbSICNbloIwhJOR
ToLYhLma8jQRifTAeLa+bkFGRn8qsDX02d50s0L0PW/jpvZSrVwvyfV/tsnqJcPo
J+nSxw04jjgNjdl+u7oIVsr8IB4Zn7mtyn9AC+wPkVUoHus6KrBtmIn+MrPFGRfz
BOWT7YunPugWAWeBvRhOkIgjMQoTYmlZH3KuESjZAkWQ3dIIQK5zxrk2XqCwZWRa
IPeW+tLzV2Pgx1HGLmaDpq2KydVRQBJ4EUCJ7k/S+IRgmoBkhoXyDqlkfBsh2qgb
h8wzgdmj4jwu7nwVTSudHPKKCAFIqGcB5ui8b7Sy0pJ9zwv009ka1oZ60qyilhQ0
blaS13jOMEfH/AcULu+ylpC35p0CRfSOg6UEgA87WdwdAF3EK6DDoeG4FVIu6jPE
dVaIA/5X1bZWh3meBdtfj68OWPKJSMdQvmqywtQGlBoLYj6/br4gc50P90oxvRcv
yuKgk/gEEGgzhYBGGjvdpMykaXclXpOe0kx1C/PQTUyiPKT6xdXx7CmssuXbb+iG
CcE7wJbbiqqBxo+ad3GZKg+t/JYT4i/ign26Re4wv6lxICMoOIhuwb1HG+ZSDVZF
jk+vqGdML0cclvAk8JSDEfD5kwXX2KyIMBWTLw39nPzyV1td0p1X/OBwJTy0SieQ
jbg9vtuqstKsbn0C/Udhfva/kuVEHzFdu/4L6Pt+VD92AbqU4t7X1Byp0xbnTqAF
nRCJnO03jh/vst/yfD+6ZX6ORX0SRnVpI5vErhZZG8TkceNnB+x+fitw6KXxuY9P
v0CShCfF2bW2r+mEC0reYIzhSKN62ISulcWUchlDR8mZZiBhuYYcj7mRGGhTCidO
MX7GbKH5olVzooOONmJZvkJI4jfA3Zl0+mf00kycUWekA9pad3GNllkkYIYixHIR
Cyo2hlpbT0N8ivHb17i3Gjl1jJSeF1P08lxadQSt4LBXAFIeocJkYVYE1DPCkILh
YfJxUnj4dl8ONEAW9c8ZF4tUEPNxN/OftNR5IyZ75o/Y+KfYBuarSybVXIwvrJ50
BJ9l26W1r+ByCLTvkDdX1r35Uo9COJOyuqzmMTU5nm8XCa6+GBW58QKNEYCAcKYR
SMIscwYM7SjVGpqC+etZO0tFstW+Tzkwk8kjBJLyVYdsO5M3SrncQoalwmaPQkNp
pRggwo2f2bj7vuGt7GV84C9QK/iAuVF2C/TJkmFrjKZndo3wft1RkrLeHITAh4C7
lLcI0yqLBWwxOl5O/S55gU0Si+O3N55K4t51WQtb1rJY1iUlD9/8/FGNGTLKwekf
FVwOtpsDftdz6ke2I9J6fYQFSOeHcLK0wvfJ8sk9mKgQsdAENOfS7eYTA7w+18ky
vbh6rsHmkKiD6jjXm2UkVqLmoVnSzVDuXPTvI51z9d8C6SJJJN24M4+AkDlqRaSI
PDeiNA04GL74F3hmmbBrrBLbizi4E002t0WVWz132ZxrH6kAO8irqnk0DrlU22Vm
K2iX6i8ZCFPEjNRMKkPjbCsiMw8gUcKU5+9XU3++gSc70SXzC99ef4Ks1s6o5IQH
/+U98yKIUNMPJnBPcGYPO30QXmTpCofQ0AQ5lhkCQOfhVaXBCdVZ6dPJd3ZTPjeZ
H/wHnvrhLqvQpWTRv0/T0GpdjGWFGA6YFL5lF+BEyAbvo9l13qhMSrzci40wiABm
QISgsQk3loB9z0+fqqGYX7v3f8Ob2KlSwSK7MTJ4b48vFYm5xbHUiOA0DsYtLDNx
55vOTU+AwrgGcxCadjurYCVidnOE6f5WPTPLFYCPrsImRo3ia9H4Ek2HI67xc6T0
q3/r0tomwWNwA6Y5Za3hu5CPdBR30bnBpuLusdqmzFsys4SCxFArcVjFhDGW3FIu
E7TGKVfvT8HBm448Hih/H+VmdB0nmu9bbRxDKRbIGgHlI4iGrh67IQUjSwDjTibN
gR+mU348Fcwk1uyzK1aX5zvTNnMROw4yBO2OWPaax/GMr7DUvijTZFhjE2RUJ4YT
tTBupkbFU1yCKFzcwWBxST9c6gTI9YTxnZAMLi3n3bXMay3/SnHi1l2ksRrDVshJ
mQGXhp3LIcnLOH9wjgeO2lD7tE4wrVLlxrDCSBavyTFLrZeDHexfmmwEVOjSus5j
vkGM9ZYNm4ug9D+FdwqPrE3bVB1Tltky1K7dz5zfoWBaMipubXxacfhKQ2oADmXg
sWCm3smtQuWdcul5dCo+KGkC8ufaVqzl7avGdeBm/LWW3TcwfFfzy2I1IShSnlXL
GHIJn4x7CEgyCA55eFRoZDHYBf5m3YfqQZyMgXEclkuA2v1tgMOPgeDsnhzYAKSW
J2b17vU0bl31T6Mgk4RVmpoh6ho619qy/MZ2kGa02FZ8VSGi9Arrl76GWzYsW+Hw
pFCqBYtw6iWR+ZmiZpDbtLYbqZWBlSCSJcxjlqCSYN5RO/DwzCtgUsQWwnHdeGWn
/4bgdM8g4DdChzR5XEiHMwhgSo7/vWNO7hFRgxz0vgrK73TNmWlQnI+KWsDhnjjp
aPiqBroUA0RuAGlzTjZn5wWvQy/D9HjjoNUWSs/g84f2Sku/KsPWe/e5AD//FtGP
XwBueDvcyHlzK+jkiH49B/BFH987R3qV79MgzXbz0HmpmkL0iyysRuZKX+BJWeGl
hWJbWvIywsBgpFZxpXYzKjMcctdSy+vlTGgNTWd4wAl1laU5yy7Z3eEWJ9oKs0EE
CSmV1hcbNVNm+BoPf7WaPHQ17FD/w7j2nwcrDEMNiFiqNB1daEFgS4VBo6gyaNgO
kXjC9Gx++hl1UeL412sJdMwcE9g4blsjIbDiwnmTREBNeZHhXNu+9uYQ9k0+RrFQ
lZ755yBiy/v+V5sxu2N+IZkafQgM4X/yNbk85IOSI84u4sHQrC9cbnGWnh3WKcWx
DhE37X2itOqXebMXm0JNoSxF70vEtRfL2+UduBDAWgPxMfOxC+8EK24LArOUC0sL
n4NAZmjLB1wG1bDbx60qftZloUSWBK0F20IefpRkaBGY+BThK6lo7ApKwFR4Pa4s
4tIyn6afG+ga3Hdh4iKw2LgBebHXT1v+mC+15WrK1K2tTinRs7gi7BobuHjCYEtM
K4lGhReQJv0XgMPDlt+fnTThjAv/3hOfO+AFMhXrnmgpDsC7AM2rignX2EA0otbW
g2j5Nu72aIdwiOFHMXn6SoX+576VoWdzXATbxulKacKvn8YaFOrzi8j8GTJKy5yX
l2LKXlXUmchf00VDlWyDlNn+Wgg2l2tjpHbBrifFX7sRRI664zkHaYI14ubMrLEP
nnroMKBgG8QJ6yJudh0akkchKs74nlazGIeZ0PGqJuEwSnGytTDCpHzpZstA2eEa
S+MPVvjHeRkHRx+Pu6yVaUH9BtnrwF+MzxEUqC7Pkw3okSwc2n4e/uo+QfSEoKLR
fBcuvAgb182fieSw9lB36/WNgParidRtJm2LNnqQ6zTD58Tno6g2CSNNiIyrWirD
hf/z6nBRnGPlBQl7AZwPIfRDPhOUxCNEEakainCEHo8wr/Q5k0DUT4X+Zd01QBHd
r9aIAOyoyCMqo+acA/hOiD4IApEj1tLpyjb8Sl2qFo9hkxyubeu33JBiIf1AmSVe
kLx8vWvLCFRhG2sgCUfeodnMSNKFdP7BokqLZGiJnXVpKmUQtdA5zQSqG4WsDcHC
/Lkz8yNlflpglkEL8MuzT5Cl39/j748c3ueMJMWBlj7Gs7xeE4SWOdI+taTlClSy
VGU4G9NDzWVngcg9fmC20JpGLkIQTQ6JoSbVWEfT6VB3zJRHpZT42IEJVZEn+v8U
K0arskXpwKO9beuHS8aOTmCq5SaejPLbVakCAPUWqCfh7YFgbP2KyNlydieuHGLk
aJ7EVKg9duxqlV9dxU6XS0sKVE6A1UofFLSKJ1RxEKNOeYzcc2SkLkI6G2Yby+tr
ftlykfYesJak62qCAIgMI9db0Bz7K6cE3JoSIoIaMoFKNZdpUlngjYLZZHa7xY4A
vIbORG4kdpZqWU3ZdaL8NGYuBFYmW4oJeKY2irG313DuBzRDFQuzh0VwCoZSWV03
Qs370g2eD8RzSH/JXHqDNEUVk5mvnjAZmATnI24dwWkQCOnBqyXNO73YcwChngVT
WdSpOVfVoH7mCcMNxlYs7yu/eYzpkdNucUTNtC9kFA+E07Lsx4Qp18p+sCvZeZv6
q8i2xDX312/f5GXTKyO7pU0Nv6LO0iw0NgPbDZomOwBz7lIHs8Dglb1W/x9PE1sA
eEQ7ELLFimBPJeldpdXBYJx6+6OmowOL610ced8tGDkUeO2KMlf7YV6MGbItVJBG
sYlXhflcBelT9l7HLeGqr85iJI560oBLYQqdvdG3OOrBY1RWgQOrvffCUDXmdBhL
3BGqzf8pQ3JRm1pw/rb+nuE0B/ICAPzrp5s4E4dXwxbNGEcBL+nrEJlksg9LEjeL
lcGTYGwp5/7+E7XRIFdVVr22AaW8e2XfrLfedlPdKnDPDStCB8cv5bCv+KfkD5Np
5az7j8yVbiGdmqN9PAnk1UPU0fL+tAsaqBCp5sWFqW/grmS9/UdI7zTyfujdqGgN
GO5qDktll8GpAdIaN7W8bh83sSjhJEmkOinKxiyzuWRbQnUEpynJOcNIeJ+J2VuX
DQdlCgouMTVcC6kp5zNTYvNxQmO2jxtMso1kxWOEPBoRKGj1vHpyCN35cLvKxo9C
vcbIf6vopiq5QIpYVK4Hl2/Tv5M4RWE4hu5LqH0Eq3Ts60+vNogJOFgkkz/Yz8kY
i8rcsQj5pIV9kNvkXlE5kfD/w1M5PjkJhWqp0MoSfCVcrYRe5wF9OIeoI7QeXK1U
Joht+MedS1WPBwcu2ColnaD3RwHl5YYjaEw3/o91iXIhB/wWbhGtiaKbWsGXKW9/
4sx6AmeP+Dak6EvAk183x5R6ffoExzNWQqChEab0ZDfNqQymwlE4NYiNpb+vKHGQ
MjeoiGUW2UpBnGGtzNFieQgaKm1I/ebIU2dgusKZHTbnfKvfijeUts16G3Jzbbno
NhtnFpEm5tJo1+YR9nxRLXehQ/tQyTLqgKmTULGOInyKEL5qceXwOlgDIZreXTIk
7uLKXwJOfmEahZ/QzI9H4BDN1byeP29cTXCG40/A1Az+c+gSA3QMy+PW/oOwNURK
QK/ZJ5IyoI0ZCOtocVCt0DnAFhc7K0LPNy2hGgATNf472M/RrXpw2V5iiwAorWcK
FvDCC3+6Oa+R0QAjFwPnEO5PA3OcJgyr6IoDzEqraXcK8OY4C/qAnya/cFEwvFKt
ZgSwBGbT1zbq99CFKEK/bigEsbqSDiJEq63xb6VcccHS2u1UadhP4TPiHWIQEcDq
cVT0DumFU79Sb/rzw3z4OLGJy4dpazAxohonG46sUI6UU0EzyynkijL9vm+RBTKE
MLsmOIkO5gk0rJePi8a8e882Wd+owZFp6hGRDjY0aISD1n7Q4WQ3pC3zPy6Hx2ji
VuuB8Ouy++dLS/xNzQb3bHLDPrZFwTF/UsjPai5IpyQKKKnAPCWNVUbC8k7VNW8/
65e4JgAYYG2edlCFSn0v2VzOfJVKXCh90hZnR6u9GrHNrz0TDbxLY3un0rn5b9V6
RNzr5YbovWy1HUvSILgV1r656GY5TFFxNjc8FaIOgJNntNsWd6hKLs7X9DeGnceD
D55+qlAnFyp9InKS+xUdqJeQYGoIkoqFcrc2aRsTfh5yH5y7gSk/P298NQq3br1N
P43lWQKpnqa+2FrIjqSdThE3iWLc3z7cpdtAhLhn9bM0laba8FYFSecLELT81GUy
0ve0jjuoHLnMXnoaBl1fsr5208C0rCBwGy5BlZ+uwl2nQwhr9JV+Cu6dZZRAKLld
Xn5kDEFMyi3uvvQ1CRalODWlmuOYrpHp+CybCJziRzs/7oreDCGiOOWjAMALjanJ
YzmB62pQVP89lPbwNGJqmef2e9oTDbheWUg4RT1JVc6UO/5RhpTL8hqfBbKH2Lt9
mznmuoKaE9NHKXqHEtVMoQE2fZmlIwDCms4xuAMsJU1mnuoRNEnuKbKqetMyG9BY
Qgm5oNef8DOrtQBA7FAvnqtY0kK9hVWj6irkmxdxhID2KKz/v556ymmQwD+kN/zY
J124kt6bwKQLuIXB3DRJz0QcAgE0/UEKlbsN7RPguTFVBvebhxX26zT+/L30ANoN
qk1WgU+4bzLw2dg4fYvneMrKrgqaiPt08WDbjwwpfMvJRthHlYgazgFQKv8ffMlL
mQdv1Lf3Yy0iurPYC5deXlbZ6onxruELZvEIoXb9NGfVHZqlmYW3U28Dgbvk0AyV
9E/D0PBfTAgd0q2jTWeu8bx9iTqHih0FAreDLUkIMki3T06UMhQOoe/TbUkUqcgw
Z76BOSAFQUT6XOoXZnaTL/hahxQ43cL4ogaa6jPWWvI+1oLwzykr/hYLFYxu1x5i
kRiUl+Ool3mS0XQkC+Wh+AIWGbiheOB5OEJ+ytFhmZz72eOxTi/VklM9MYzOgkzT
eEXGb+Sxg+VPuTTHGxT1I/p6uNJ2lsea67FxAjyHqLz5gV8X2hTNx6/EoiBQ1uO+
BUlt3A/dhSjkzXigcKGULNN/XgACj+V6kGFoQtQfUBkt3PbeyiffUo6yP+hsoZEY
1bF0IHw6GWAIy7e7wrrVFN7nTlfwuwlu+JATpZDE2rpvYP2Ts46KWoXZvOJY1D01
vtQPLXUYBMJ6OtoI5emexRIMgjYrydSd97AOF1z0ijPW4AMtCZP+MhCNm2ZISxLm
cfVCrJ0zrWMtxd3vL4vo5rOn4Q5vR2RTZr87xo7H1rvkJIV9++YL5pROWf0Yq5kr
EArcpelcNRyiKZvpTRKeH+X3BvbuQUFsoyBCJxSALtO/uss9Kid8D9r9G6fagDsU
L+4eMPHfHgzTcezTrQ/Q7YoakSFRXmz/DIOGBm3cKG/v2OxoBxaTuK/mGjBXV6OO
ughDg0d2U3dni9VURqJa50i443j2PDg4N4ds1eEH1STJzBAs+uOcE1lyzFha9qY1
Ff344HdsDxEb4jbVVYwx3szP/iLNp8bgTGNS+PNJjTzKXwdjR9odR/bfi53CIdx7
KunDYdIRjsisGjuBPV3jX0QteYjDLHQbdOyYdZGMx8yuYqynJOmkDwPNnBRATh1S
AU1tGIRrykQc2fJYTECgnibPnIVd1cvT/bnGVbq126tcX1nwYpsEv/Z3oT8OJ4Ry
5EBju1L+lDv+SjCihq25oqvYXM5txgR7cUmb7Cdvsz9adLcnymFcyPT/jLhrxx5X
eTYHII3UFyqyUB1Miw5LI06ZlDBKLIbANYQxfqWgnTFtWES5Nz5ydTv5Jli8yYiQ
ATQmqZ4eZuaNIexhlZSvAwigiLKzgjoQvcztZ6HwBxdWiQqD5Q9RN68MnWZ33SFf
czuUBConKPT9kenvs3ESwmG9wT52mmV58qW8JYWqPtrpi40AEUlDlKKmmu2+xwgx
diojnkWKgwJFndO6uu2OA+yw8xyi8Icz89Kqva8ToI5QfR7a3APWUQHjpaJ+d+OQ
9IWdnZ2KIY9Ukrtwx09W8LlOZ61/PQOixHG1Oi6q+v5z2pX65gAOSZEYQ+qANpuS
zI2542opwiBnFgFRuD8gx1wnIphA0dXAx1Z3BeXVaVz+lStwCGk4PxjbVwq17Gx2
r3gEobvU2vw7ozYAHcX9mzf6mdH4aGjvyDe+JbLaCSwb/KOhK03ns3anw6+xQaJ2
CsSHXYaGAXcn1hLgj8bRxBgxP+wAryXKeqynXUnqnuB8fVsbRPYNZaFMWx1MfXYv
teLV4x7E8N7qINNiB/d65CRJB/WZFp1mLT/MH89psjhtHgXsT8+ncpLE/YVm8iO8
KOJ4Mqd1+sAnsviyD3jToQPiD3w71xWVrNjQQ1ZuI/wqP3bI9VqvE8yht/KHQTPv
HwGmeKr4FwLKYn0GU4Rslz/JM33UnoHS+FutkFGsWpar7WZRljQWPkjWSOUBlQ01
Y+E50yvZmTT+162pURKUP5r20uczJL1WKcAKlK1Ko8ogW2r7sS8QJg09mGQq4rud
peRI8rnONclDwNO8udKcTLIeuuhzuifvtdd9gTPRw3BHOJ3qYTkpufAYaYtYqryC
90XjkEWHWIm068Q1cMrXi+bV8IifpTaNjLyAJ3ZZH9zJHAnRSjEfcN962jVrRtV8
1A+mk0JkRtowaaQV1HNJXAChNY0Y04hXRwoTKX7ncKScF2CJIJkXrvjS2P/D19cJ
eAWDxjHSAChIwD1ygxfXYz+JCsr8MqdBTdeqC2cGjWpWS3p421CcoNwGGBvNKZHC
9ynhfzGCXjv5BoinHJFc6tg4QUg0rpnn3uTfimoN06TGVAhUjCWCaaO6G93ILu0f
rmJSSEfYSFhlOq3tGmRBurWTgwhIMBiwJq29ssnAvgeJqbMdOqcD0Y/uwv5Ihu7i
eYbDrCmqpgKjD54NYUUIVxUIfs1vWisixrq8EtvfYZhWS9kcZrWQfcXG86dILlrK
s0Ow3zpOdFiSFK+7oy1jiVVmQiBLDqxwWjPMyR1U2YSJLoxBW6TCTG7HfGBbARQL
WpeKmlZWy3H+oQidSTQkK6+yEUeZDHR95vySt+Hxl8fjfBHx8ba0hbstn2vCaELg
GGW4ghIeTQrbiXUbLli9VVTseF3IadyE/XcfP6Pxcg1LZ/whh+d7IEH+poO92rXZ
hnGVbvrnlrB4zAtEpDLTRmDxpJDrKEDrQKz74lWZYFTUTZUd4wgJk/GFyVNHMEAt
Ro2e10JCR2wnerZYBaLVcTkBvyQVhQBzgfEosULt8KfsFKxu3IcJAfnSN12cu93K
nfhsnb3q4n0/pVrc8/hgMw3GZp93OVOVaZlSaXz8S+KmU8PsRcngbNMS+fexwDoL
ecko8MifzcPwAgfLCAVXXHJ5wBNFbUe2TBoQAlJYJNxqpTQeMqT4Ymj/5f+Sr19H
ShPa8AIbDnVy5wtTBQdyjB6BqRLWQvJkzK+1A3bmwTK5SoMsRhWunooJlkCJNBVU
x9J9a2c8yexEr50rQZr8v5BjdrPhvG9iGPHEWFBMAXKhz1Hgeyrc1oYLCY0/zEO/
UYp2cK1bmd7NS2+qS4dQQjt9h1HIy11lon1USdJ44YsllFatoG2X9iZKwS3rv8Zp
fETsv26e7rG6LmctIPbMOa8ALBzx1qbSg9T2OOmu3hUaGr+PBUn2Nbi7JCNVx2Pj
8d4vN91wdIvou+TE0f4dH4RZOpFAbq6wcgSwrlzOW4XK8uyP/aP2DYklcrDjkxmg
aLeuHadeLl8s2dATwvQ/8mCLh2px0bLfioN6GCn2w1oO6a9j/nleW7iDTv7D7UP8
Ohi4zOOze1UFip0xWXOgv3LbCV6/hVwQ4itoPzQAGoAo4BHANUh5XKgPdKg6U8B6
BSnjfUQDDCow9Q4PoXO3JC8Bq99JbrcKWIIomQJlSWyPQcg61lqnr1w221gwFSaY
I2NFpJoPBNpHKJGAKVR3rc638obAGTRU4mZSTTtwUPSpc4GMX6LyFMPP6dKZDw/t
fYBuks7Ke5aF152wiYTxQtIeCWEt7RP/Yd7g8jo/h2Dow1jNKjZade+1HKAGa8/Q
iVykgN7/7k176IEYXoMFOzVf3iWXtjcWOCI2DOa9NcvAuxd1fY5Cy7z8BnxkjW4E
5pWwgKB/IUo3WDhqUk9jUVpwNqG0OyVdPySVdhwVH7YWz7AJd6VjM+reeEvRLeQT
15/AcOoPWqQl9qiJp6Acos6BVklrQ6ZaQ7uVCutApXTax9E2sGUiJKDSUvsHoRkj
bEimecr74RKTgm+HqZOS4VZItvrI5U9e4Uh7UsiAxfjNjhbe5GRlJL6R7IVVFJFn
rRMiDLHk4UpB512HiMr9Tg74Ew0RjUlL/i9ngMRVBiYJjJisaquyczHM05kcdWKT
SxLFjPwWCvTQE8jHENlQXcDTayFA7tQ/QguU6oZHSVR/k5WAmJDbxgmBvpWKVEwu
9UoX+mk9Hg+0P/Y3LBSZHTMVpTMvLNkWBQUUaHrx9llv7lJqO0A2fbgh1ZecMPjR
Fy4/WFrgedd31sVNpES5txlzN6kRqoNNBzWc0YkJNq2Y/MWZBB4IpEny8Pt5oyn0
JVOw3vPJ9oM4tBozzYEJ33ZtgjR6EH/HUK5jd9fMBn2TI2X7GDFHyRZJs0pSzPkV
IyAUl9hgvux5evR610Hy5fwlT2n8eiP7cMssVyZG+fCa/sNJlfD7M91WM8C8Tctj
eYrea1g0yoUj/H8ORbdsQ9V+qzZzI7mq9gFkmirFBE8LgSDMJMG56OvMRRPDfJsi
RHvoH7LGK4mYeV8zOA8vI5vsk7l6knrCcC+2Qk2027pHv5I3eHuHLZayD+JVCTb7
F2rXw/8dmRHRr7eG0H6mMwMo9BJoACH2hRdecA5ITn21n+N7bS9BnpD9xhskQ6Et
LCX96wU2Ocu8MXuYgX4KBkTuqQM9I4iwrLTDqAG2ikvxMn+vlEtd5z/rzC8KgkLT
128IlcriVp8QmWBtGemPJYiYg5DaocnHTN1ji63Q6ptVu5mjhbyY7JF92/+S80BZ
eODqaVGnLEUriO9s26jYwdFLJ64lH5CUSprASv5VYWLb0djaMh3I5pLyoZX9vI+O
pIHhmhPVm1CyFoBKXfHZcEx3EgDzNdhIIl3+4rxmWLt2Gv8eCuHr+s5dStmnWrFo
ql9ESQXkMn3HHOwHX/YBJCs3m0b5NoXX65ncSp2m/iFYZPy+iGzeW6s93fLttZyA
5y8vF+KkUQdwO5RvmqNKNQHH+AIspySJzbXoJHypvD/ENgINw9cVu2e8POGB4Wqr
FK92KwT8L5SRwDBU0XCF4uf2HloGNpv+VDV4e1jE/QlXGlf1EQbYI6q7lZ8NFDZv
Sxc061uRojSuYFttN567Qt2J3zPc56Hyus28sJY1GhAJEGj5fTZdwQUsYk14fh7q
+ShV4RgrrVh1nCw5VIzytKkPMqVaYQAIHCltaa7ebjvpQf2EPUna1T062Qd5qgNj
1zAxKxNlAGY5Rg6b+GrG1nsPM+BB9J4t3L3QvTZcynW1zIcVKK091AJSSsZShrYW
6SuZ2nvxxiZuTCUzjJucSgjgOtDqPCVhOSD6ME8QX/jwiDsXfC3cvEDX7LHbg/8T
0FDjLTkOMh1ZgW28ObNrDsAc8VHKSewEO9rcwKT7Z4P+ftYUwRDffRUYoR13cliF
MOXZ+vJAvS628mJv5DS2kyoByuesWZdCdGnxDYzL8ZqQvYT1tJK4nrhkMCMQp3SE
G2ICScKd87jBRwTqKhZTu6YxVQz6CXOW+VkxzM2KZCdZ9J4jPwTrDxene5oAkyXz
C9yAIMcRHi+U2m98CfdVevYw7tDXu9bKWeJGS3Px8YNPexW36sGmT91pP1o35A+d
JgPlqUSZIkyfUqjDo4CxRfzXnMfpSOX3YGwC1IO+6zKgauAweVb0ChJglG1iK4en
t7P38rv5es/vW2BiHs1L6Rw3svqmaythqV18BtYahBfIvTVAGA42QlwT0p8RzaS7
qv2R98uc7tJb6kzEkvGSvV5kY+WGxKyZiSphhDELsZdfluidYbcbYb3mVBchrI+Z
RGK66b8fZr6/Np7k2wlJM2Pm4Eoe9d1O803DOPjnfp+A1Z3s3rgsOS5PZpRglhaF
ZzMYQuFYKpwH4z9thHD4Sp8C0CdK9IXQ9VTzk3mrCvoerA11TbrFgbHhaimmXaDx
ybkK7MoahObnBcE3KdSSyvjLzI1AVXJDStqfM4Od0yReSp5okmZrDzT0atrQV3RY
GKpHZitofqgW6nQeO/d2jFEHaPzmaII6Q95d+goH6Ikd6O+z+9txrImKR1VRbaHc
p7UGm4aVFriLHipaTl/yi4ctrL8MHfhIZAFVvvuNw6dsyi22pYHhypdFNa2MwBgo
KoU8Hvq3XXVFMJJwymKx3zSeSjAaviNaO0OOGrOxO5SvLFX03EL2XHdNwhacyG+y
lZXoVxcLNgkGymQ7+UtD+VMJJQ257ssLRMUFI3X0Cb30rZKRfCCAAFVcvIL86e95
MY09Qs6o3Ffebfol53f8VSyOVJKL3VbSNIHXBs1NoocmSmACZE8iBsxktXCRBUb2
d/6cGIIETkkksuXGnwx/oXfImmNsA+h7mUsuoe50Yra4PhzpSViHN6HA1xmYMNl0
D/9jBm/jTfrbtNc2u12KMoRlOGpU/p80qF0TzFmtOcPzxNwlUKjblLNl8St7Ibra
ydu4nG87QKlHgWPa8K0BE6KObelflvlLxfr+DEkg4J+M+yURZRlprJ30FT00CkwB
x9TyTly3iNWGFlQVaN48Z2L9OGm58+VqDjWXB9RyO0a8B+VJVY5AtP4rYtLz2l7U
Y/WOcvGZjDGIcWfxF1tLG2IufmaUCI4q8rEo8pTRrwaXAHA55rXT8ur+HqGPR9Eu
AT6m5ysws0gymmPSZobib41XyVoXXBs40WEMxokgu1auOSjyd6DlWTnPCVj27zZd
k3B3EOWUOPSQk/Fo24c9lJx/BxfFo7l850Xl8cOw6QmsYN4O1u8tp3g7VpMytmo5
FcqQAHa0nyGROGjRl3gyttB3T0isGR4/CeDjiw8uCZpDU5YVWzwh2QcK50aWCG46
crsT30LJ2mAUQsWz6vj5UjBlP+duXMjdcCHreGD+JpM0QBgrG+qPcmiMA2zhgcNn
cSKbUXdev5oZif0Veej5XuGYdA6BX2n88vWtDtHpn0s5aF4xJ8Hcce0nK8ViWRYn
lF9shMq7q2+CfWlfXZN3ZvGC9q/YxSxZKhc00ZlInr/BOLeQe7I1TF/BT9FBWriA
Aio5o8Wi9PkG/Lc0Ej8LzkrzsVRJZHIh9Rq+KisQHq38HdiKNyK4XnFunc71ZZmK
AOfRu5BuuLdWB7BYMYv6em/5ADXQBRYvTEL3Y+IBZ/6fcExhmdA1lUQZq/2lnwpN
SJsdBkRIf2RYETg7qsqInYOsWdkM8HJlNc0qEGA6W7MneSpjw108i0aoNnJkjO7L
+RwIb3h285P0l73j82e+dMbgmAS4Cx1gvSvTsLLiVpicEuoBtzLQ3/eRGcxLKoE+
zf1IrbPVznlZOacnEJaOzDkV46fJnnNC1mKPGIuylTHGMw90BVPhMI4QWX+BWp4+
6zaOR/C7iYXaw7QwpROUpFF5bnISL6x0nfj6An1naI3PCYbnDdgNC4Fbr8KMm1Ki
4nMKnZVJZ6yDr/av59Kk61G9++lxXaXIpPTu4z7fvkO2WIW7kd2guqLLVZqZq+JF
PZByUhrrlyv9Fd1u3JCCK996FylkRb3BY7hiUWrqNaUtIv9o758wvipX7VxR6lO0
1Ri8Ay+uckbbyrWzpCBGnO/TOp5Nsni1r8zjcEsZT5nfSIrUivSuaC7L6TQU7sZS
MiFAG1AwtKIYwn8ZsY+acdbYk1DSdKqxTmjPmZq16G2o7TGlYzZS0CZyhpW2NaD0
2GgHp6CNjCBRK5Vu9oiRmuXGZI2ooIG++J7q1yX3HYfPZsQYg+cymtoTW9lSPRfj
ZAsXGLhPYouxEUNez9jn1BlgFbS4TxmSNede9Q744mOLLTMSaa+kxlJfSPbFCA7p
ihyLppxzve/FvzmdNorB35huvdUBtVzsEByRfdzvDj7S6X/lZUpT1L1/ov5ImBQ1
qXs9oUUNuEf+7WCOBcJmSc/HvvBQY6p0v9hizSjv38MFB588XiHVWz6r/qlBTNbr
3hbQ1dbxSWjFxjo9Pi8F/Xeo9dxs34Qq5bdbpp5qEO7DzzhK1Twtsg5Gm3zD1z3w
2EtGW8hWssgIoJhKHu/sm44zyBdx9Ls0f9DTPDkyDI0AbaUt7X7MoVJkWnXMa3sD
iWsAshVGgOo9+4mJQxn/iAEso5nhGt1BDDHgv6L5A/Lug6NN8nwuP5H0drau9qly
rUqF19ZkAArJmLzeSg3QQwJxLYNpJA8ICJTNCYYmkPByOcTSAvh59RtSo9VREO3A
f4BEmPec7CZmmmT2ovNAD/TXBfqcwmFf/XrF42L8tDW1CzQnHr3zTZNjGSl24Dlw
3CicdfCvkw9A6IIXSCF6zM7H47cLLiMTKKSRxYHw/K0E+b5HXuKjSmcfr7qGPil/
MpqLKyJjoNNTRXMvsst17QFzb7yD10dk32qhhjdWK31KGsFsoOgTShJyr4S7MjJe
Kl4dRblX1D/7N0orhjXF946AwWij97MWPcPhrFt/mlr5O9NwduWwsUnGz/64ajt8
G3pv/5Yu0MttgfThsep4a/7blWxuaeJCaIrOI9sROn5tmgtkpxSpmz5DeqaeC8mz
pIwe/3dFBr9A0CYr3hJWFeg0G2kwcEckxLmW4susVR/oL7ET6yxmrvs5gKEQLgxx
F8+u8+XlLUfqcRXA6bDsxrnsFlvU81AsWpPaPsYcC8WAgM+5apRkE6uSS0pqhZJC
BlUM7MfEmUJ0GlIMGGwA/dcAlyEVl0zivOrleYAgo+yQU9dfpDbAGE1MUQEZXEo/
FC01LZGD1nRZ/GiECerh+JY3BRabeHorZQ9qk9jB9sxSN6wSygSydqX9oKRUYgFj
Ax+2XXpZP9lV0hidBsG9bGPwToLCOsmff91++dw2n6wMwGatN1tRngWxbkWPNx+1
CfcwJVa/YkmEt5J7SApq0TvbmscUzx8EekXJnK69WETki8bNAGDsccVS6/aBZAOm
5wZ5VEjESEePZ053hoWoR1ZOwpb9GrKicAc9oomwKv1/v4C+oHtf4WDMs+9a1hXk
nTZQmv0cNlU1rfkFyA2gBJSBkv2yueU2wtL8E/SiW+6k0lFnUGn4WdNLWSL5oAi5
6GB+Qkb4HgXAbylA15BRpzxuOgvLfj9spJ1+SogYl/KUm71RpxdE2lJQNPgEhB27
mX/7GVaWqxMKmuY5axJCDDJgorx1f6PWEaeUjoGIT81z91G3VYc1qy2MJbwvwgp6
12Wi/HSZAXmE3gIrny5/iIknt1L/jGDeYEqjeXYVVMbfc2EBJqCUidKG7Mx1imIj
1j6hsYHcCpp4dHwchmzK4mCbVZHoKKX55I5sBmptntMEyFYNBwKLQBX3GAW/ntL1
zYQrfJ40ljKrWavQfaeQR5jhLX3WyHX/h4v/if3Iy9x3osgKIfXvqJXPh2gKVACy
nnxxXP10sCgemqvRwkj6xLQHRgzCC7hXTUaaKqw5Qt+lRaE2qoLcAbmPvDp2pbmI
fPQUIiMLWMXFjJJ5FaQfevy7E+Lo64rlBemnd4Ub2vreXMTIhdoqUJYzuNEOt3jO
50jeoD3/sIa8YNoTXt/ZETA7a1DNG60slkL0hEpxYetH6vJ7SYwsoeTFrEw085Su
2bL1G32iJHyBamFnX6JItXXswWpUUUDyE314KgBx5Fc148zqgm8uE4v+30YYS/Qc
fhVCKFM8wRdO/qz/Tr+/aFd3K2k4H6Y/6TndJKIx2eqM0ctND3Q8/ClJq0XjLzV1
4IQkgPXglznEI0QPmOsVxBYg8NiPN2zLf+vC53+kWRzZmyU7+FnKnn9Atkt5LthF
a+MkW06NLB0YMrbUqqw6kwl1dYXT7id+qWfOllnLZ/ab3/W9M8aYHAh8xOtoE6tW
AtXiEbRNbfK5dWlMM9MOernkekvCVx7Faa5WGb2QCY0540Iknvo25Hje/2+iXdDP
mbQWZrKUoF3KPpJhQEdS8ZWn1K1xK7qpaOdAl1zp1uqo+ygpg4PBi4e+7CtS7R+l
jJGgIg6P5yChZE3AeDzPs/2OSYbOvqWVXjrvvp6N1CevG9IbCak3XxOGXmcJ4QsE
XUANjbCdisAHqow5o0OnlSgulOZ/P01LrvC8lHbrG2uLL/vUNCKxA6WFe/yrjJyj
SVL5ziGjxjBcWJjCg51LmW3fXBO1qnXdXc0qcV+jZRlHCUMiZIY4mJU1CbSPOX3b
3DHbsGSm++ZhFk/cfnrr9gVsggAQswA5zIuwOr4uMLNmYlnoWuVFuh5Ahmkr/Wjq
YfBMnHaJ3vXbrPnJtjxSI9nDDqqalDgOJzsqLiYArPPaFP9hXiEkLKVvUn5mfZN5
x7DaHlsDgvxaGxRJYA7DhOB7yMweaFobe7ig1ymyo/+cXkWuSduXXkHCsShAfHlW
rtldWFtEz1Q7/9W7i/rL+MyWL5XJ3gzHeD5oE4CW8m3lMbm042+2q3YrRqpTNKts
G39zGDAuw9Kva/u0sodNkHNJGcc5U2IEZbd6AdEhKWavfcc9Lk7M2097EaFq87Bs
gIZsPoPQDclw81XhXXQhws9pxmVFrxxtHs29SzjNZm7wA/n6Rwy1F4ZsZe8ovrPE
f6b+mdYRCEsMciqyeqvmerb2bUQR4v6EkWHs/+jkc6LuvtJpeMBmFcwZkV96JSLo
W8x70EGvwFgtokhKLJLtN/POsJbvIEpXXiBzURcM7KRrhivvLBTvzIkMtBpTHafl
iV09mZ9PqlsfzHmV6MUu9IFdqwhL8y0VkeJ3yYrhIXse+433qsP2WDFmdu+tNDcS
k/DXbKEES95P8yjyqHpuVTARKHrN0fuIMbOXUChnBquVFvuo6gIjYlWCAcBm6dJe
0GqfR3vQTLEyK+jYfZlWwzcXEiZ1bBrrIrzeuR/JaMKkcofXNWC6TgdR8wmtaROI
cdvRknrYieMPtbLE5Bi58GPAcO2fDbSzGDXL/RgIK1mdn/I9zsRn86o71gDfrs3o
fK1iz69dfagqk29iARfEWgQs2vUFNY33uR5Z88FiqFnBOLVU6L8KRcn3pFo6/9Bx
UMg1unInxHrs+TOHhEoJSObwbZB8osxO6bJkveMcLmoKtwrZGvky0S1KJc4mh3ra
Lyq8LhEiaFfM5Uao6NIPYHc59D29zIyTxbYd9ZVV5LbfGIOL8fsRWz1nf2vLSz25
L1PqCcY3O96VPRbMEOHIiLaExbDNUunyac72tZ5IQbHFNliuAHSBJFNEA21Q6wjZ
I79MqAuGaqQhpfPlcFYmifM0qswNsM2RGFOl8YQGybdv9XfJeU6AvZ7TOM4F2UvH
Y81eF9l7/pXv3Hebj+epTvru2zAYJjrysON9Mx06bvfuHtWPpEF+b7BQmpBNYDmo
Sdo700HrEcze+nB8mSTi4cwuF8fN7DzFmWq3TV+kuYhLmLI9y6etf3795FrqPCKf
ZHvYJD0C/sKeotMT3AQtHh3KPNeS8Ujs/wxzTJ/eep43isiJPin3zRZ6A6BsNBp6
oY+uoqjSQf++ZjFfNUNkZ4/wVhp0t3Om/EcBQMfFyoad9gzCQ8wkv0UrcyYjfSgA
RYHszL+c90XLDE0dZIbmCLhXkwJ2ClfrdKwhQZHRvkoaC7nPcCyZUbTc6VT6EUbs
+w4bDDguLvM5oPbJoSpXUMoSWxd9Lv0jze3N3ZmSeaLU2F2vx39dR8cpSGKJv0Mh
nrMiKtylvF2CFalRNAQ8cuRCNo1kaODnHXXr9cdIHw0/MgJ6A1dOX+hQ0RBPZqL/
Tzs24OSvN6ZhShIMydKKVaxo+yUtOw1QBEm4dC578mOauJYlkpv/pY+Wxab9fPSD
koCyvBbzyWGd8RsWumf0kNoo7ajtMWvceJRKXj2wSleSSwBafJfo1TaoEi9dLWWb
pelk1QZ5ubCIizVmeIGWD9JipnXQhIBlonTMsV14o0qSsJGiF/ahus68brAUgBJX
O3mbgS45R4ekRnlqMxaBss3sGj5fS1lRByoJeupLCm3uSGMGozWlr+jBKpStYck2
RzJgol1TO/cY+lzfeHvLN5wFqOCuIvdDcSy81ulcWF2rAB/7hwfS77Pqjofy/Y/1
WCMtOITdDePM5W7HjkxWx2A32DW5Ok3VmYSS5D8H1aNoVMlnGYREjriFTcGbVmGq
98D/gxcXtYQnD5z4rjOErobw9/kMsn1hTLRgBtUAsjw1Vj0jh8FjVj8f6JGAuzbs
bRRGzmgwVw/xPmDwbiarp4OHi9LFAdPx5L06KbermWA7PkJAIarCWCA5ealiQeer
nDmdtTw6EIEUW6w8lFVovVVMoDimsX8yfB59vcwYYoVsbSFYmmKFVaq8cf4R48Hy
38xX7iWuPztdiIPvUdL71YJL//XGqn8SYIj8IAOTGdDluHLsMWeAZ5eieTMC1/hd
OxLNl5Dw13h89LfAwQ/HKNg/CdRRvJ0EHIhIxyHYHmKeOQblqpwWdURduvrIcpoX
dIb8U2qh4KifLp7iG/cS4VLWQCT23lOg5MgLWS614IaJzqcbhI7hyuZs95VyOIKp
9UJY4w7oT3cmTlZU0qmCGqzof91zaig2iP6a21DL5zMC6QBOukt/H7vlpC35vblA
3FlUXVlON2l+I/8bbVn7KI8AtuiL9D+zrSGnkoMmzIymxwq7TQha0XR7VKdzu+aQ
7pN8Mrqt8gOkNzjw8IRfqQG8VnmyuLf7I6XsbZWpXZTM/FyEgt2P/IgP3B1sNxSk
KUrx+4A+MZLBY7ADkyYoa+T+l5Z8prc/JExKXkWxtdqjL4xOVmDdh5AZt2I+rG4W
XhMnp+b2bTaFLgd3YIhMM86JrIw0A/Yw4LSl3qUr2ecudneltTfoZ7dznkxYvbOC
TMwDOx949qzAtQIChlj9j7uPOY4+53p5uOS5AevLv3V2d3WxQlCygajHlY5G4GYP
kMppyMfqe2UGJWE1Tqq0fLPYbjOMEmWf+ZW1t3HfXh4zv+i+hxCkP6FsKtj9uuUr
pppMJHxLaJwYYf3MHQk669/UjkaPfCbDv//ZhqrAm3jmpeecF3uwp9nv8osE8g8f
VrUNui4FF+ApQaPGtwCxab3PbarIgQqWfL3GD1ReD+ojogvzV9l0DWr3mcxMfEyD
mpIpP4EZxGpw87BX/p4XukRQD/ioDo9MIVMMHKD2R+RCaFn+revYjMAw81W1Yat2
q8A8ZTobBgD8H1fksxxhnMVnc6WQsAlHSHpHmP4jPSXY0a3x+6rmZaZgF1x39G7/
QMkte9yLNrmATg8S0oqBv6GrWBud+eLygptX6GH3Rv6WKGKlnkkh12awcD7tVUeR
ksX88i19P02aegA2R314Oy45lV38kT+zyhBZvu6jHFNLmQxpo9xjX+qFskPvRQUX
9+w+l7B0P64RE1zdOwtDGOQN8E3zrr4abpeJQM7SFjKM2rhJ5+cF/ASPaRi0qPl6
xYfkZBX2r2CJ3aMZ8a4vVjzv2PEHd54MIE24/pKj70YB2Re7Jz/WlcEai0ZwJBNo
v9y4I+8noIxxyO9MrI5MCVrFbwqlqPR+O2yOxtnZ7rPqqflXEoAxDpcYg7SZT7b2
8h2ruzmsLYSzekS98vWjWzjeUaNt+Wjq4HMznT7ifp4lOyVgDFqD8xARQ8YVgp3G
pAXRi7ucRGSsGyCY8jRxcxJwd9qvwWLDAPTkq5Ts1I8rBvxbUF9kBh7Gk1vqJEtw
HxZWp0UO6PT7cRkkUwH6gMfoXZ+W2wURmRp/784Nhki3fgDBsfwELpEnaLKYw3l/
XWB+fr+UkNlhP6WFnCdqnUzODCK6u0J5waAXnPqaQr2+gXadRGHd+wpPjR86+XTK
1otvxyakQoR5bbW5OL9t+xC9Xy68GuzpyEHkE6jtVGtCu2/kht+9ZPw+dXVkjZV/
47/7LtH/OhbEkv3gDyDZwgd0hdstHS02K4fWDjbVSozTpC4wUlX7UU0i5OvkladD
fD0zojXuae5mGCD5mYUr6+tgL8pd/jyVLJF3R5W5a2UijkeYHT14aUvNoEo50Xeu
n9usBv0jUPPIH/byxDE69lJAvqoFLj2K5Jl8MzFrh2talrENO9RdPqZ1nhfMGzQU
zeyZlMrADnbgGRatE4odFImwqD8EL40klqBeJ2Uf4lE4FT3P9LkkMUGTsmAcN4p3
lAnt7byiLnbTXj5kvzKk5leVcToswIkby47VqwrCrSX3qDoPezqK9SxLA7Wi1LNh
MGtYAu5UM3kO3Pd5w8Nwl2btHQCnCpJSmZ4e1n8iEPE/c0ugTisFlVPXej7UwSk+
qa1p6tZ1d5njCuS2TetIWzZ8lXDTbIFshFEABOuSf/Sp31u+648R546aezZHlWbA
H9su+Z7RrKOrA6L7DVX5HzZwBav3OrCqdJMo+ZODz/dfh7d+qHJYR7MNnDInXFV6
lYPvDpDqEyqXzUsDPhunpVFap1Jw6OEkkFK0pqYYQxKkOkEpztmGkBQFM79qHJUn
4e4rcx3L9Drej2kj+elGhhUC8fVpNXWi6yOPb83Q+cBfA2Bhedtd/rueVgEiEHwO
YkwK3+1KKd3OAXx6ee4owrKcGf3ZC9eC/SbDBuyNPwB6bRNcEfXE3Am1nm4I6aXe
H7LIAU81eT75MDwJma/QyCKRX9inZ4U24qeC2tNCG6ey9MODtPUnIq8JtVB7nUvs
3C6pdOCI6/nIKpbPK9Qv82c2e7WXdpc1HYmAxVQgHkUn2GL60uGKoFaoeZkfkWyF
JxPbEnbXtsJYXZR0oDf9dXQhBG4u3Iu03JJQylu9Fr1MbumcQchDEgme7Y0IPPrM
sBOdb97H+A1s3a34pjfgKzlW5DxGmtiYIjjqQicle4Y4OkqHKP1RrlLvmmQPhawu
mxj75bkzrweQjthhXu3Jt3V/CnCyefaTg+dPVpmfcy5/nEoAgIZT2D5xdO9W1y16
tOwNUTOOF6xt7jJEfbtyu8HfaZeDEs7BnzfuQZVssYiPNdB9v+JsuU7ustpfLsMY
+SyTmqjWY+soXYJjdBZf8lkGXmbDO8igzRPu6+uMrkJg2p8y0xA/r6tg0CbcH17b
OcPbL9ZkiBpxP/t7u4PS2zqlbdfxaaa84B1OTK7SHTD1AVWyN4BEyvANvRTPZm3e
4eg5Ivwn/sTdQ+I62chAxCjv4FTU1KSYpRWa3oKH5fz/+JjlFKriaDJcETnLwOIM
sDGqFAy0XBJeHEg1x4iqdIFiATWpTfyz7eZaNM5428Gm3yeCV1kOXm6gYU1MbH5C
tRUviNKKvSWLMl8LRH+kK3lamG31QHT6rXNfIwZxUWFUCox+7kc/fxkxkQiF3Npc
WPA43ndtMSw5ZrgJLcUzYkeeOAGDmYEmZohFN/wDte8nBoVQAPZkD64TmYpBZgya
vk9gn+ex+UJvVVsn0ZsDELjc06bgrrnENmi+v84oNFLhgsM9rKA6nQPLR38+3dsW
PoJN/AzQjWCErR7r4DAFaTGheMROS97Ylt+vv9idMpHZLRTZNGky7oF7apPlaCC8
LMCiERPj3vWo0IyJTS2OT6MZRv7jaZIniSpREl7+qipCXuQZ2hP5ED5DVEMuSrYm
Jc1Sm7RuJAscXaz8qynBAHefKnPYpLu/8cQU/l8S89pSt0DjdIXvsM1Z9B/IYekT
YoUA5+4diprLFxiBBnRnKy1qvO1CLVpuIcy1T93SstgcWd+wGDBMq8EkRUKIS6ZT
UflGM/PUCTX9E9TkIqjV/Yt4XaA7zs4bY3Oikx1q/9L9vsPgmAc/LjBgIIRXt5hX
mS7MRBIw/f7utYi+5GWyQBd52NDTYT5G6NdODtE721B2oqyZUmMqayQIjY+ux5G7
NFCAx9aGQnCcnE/pQcBl6MrWmBvkErIdo/JKJa4XthjsxlErEyOVPFGWGfBGd9A2
ZGbjwVShFKB9GMPK+Oajb7z3VRAY5PPooUCjj2nEjPCjnO4rNrb+hbBexRElFGXY
wt0oCv5gLdop5JlCQRGm6jJuduCMWoDVgq8QTVjrD9iybCxltm2oVLcRpMgG+z0s
dIk9tGEkKtqhL+gPv8PB2xCSPUztEtBuTPU0kcCqnAEuTs9F0gIIKLZzkGdZGGd7
XR4W/ln0m+CCnkTZ7ATQwRBoqlN0x0xWXdEKeG3NkAo4i+Cw74I7lqaHZNxGmQBx
HgVRpPFIP5VXMGArw7VU8RWQ/ELDVPDHxJAcwSLXZ0uj9CnYQIbWMFzdFXb88d1G
8fHoggO2WxLx0CKfK8r5jdGVtNT93CCrlj2ysoN4uxjPCv4Sfi/7I96kHXDdJhQo
hn5kw+zAEUa2gc9BPBzJK4knYOwhUMJt4gxUjSPpQKQ+osydz7TLJO/Sr6RYHZWZ
lO8OoiNva8+mVWGsejabYjH3qsTWgl5fxSApZlC3O0/CrhTqK79IuNJtQHwQ7CML
AVToIKPeO14AIfC9a5u2ZrfbWOw+iZldmsJ1QLL0awHMOEtYKc5no3LF2glu4V1K
/aqpeIyZ8o30vwU6qJGmNjY21ZIeqEwtvTpuhFeopYmHE+9Q4BnyJCs9TueuDFKn
VU4rXS32bsuZNfdhfgRiqqJwJskdv73wGTeoQHp+Cwkx1PT42LYpHzSUDPtEHto1
63qJquPTif0hHDstdNH5dypTm5xXmevbTH/me84inxuCpoaAIzXsvpsBVvYy5L0n
Z/YTouRYxAHXxYo019Jyc9pGdIPXlvn1X5k3fwSaTCq7jKzOtttkMfDorzDhEa0h
QyihfscDmdoxwu57Kp3ysGV5YXnTtdjpRAhCUdoffCqQ00zHmjRWIIjnCvMVtKh7
+3tSJPGR2pWMOEHpyVgbjkiy53LbVuf4DnU0bIEda8y4nSfcXSpFK48H1qPoTc+w
3t1KBRRWLAJsUaSbH5nThcK7vYeBhIk9oyBl6anU699YkWW/QsQ9PW2YwL6KhlT1
OMdlL19MninvtJsRDzeorZSMwgJXrXlL3tjAhNp8Z9Bbm2afLIo7q/7APgVA7yfA
Eh9H7yqooEBOnKdE3ukusFvEFiRQIVclq48e5wMCzcc+Bl4g2AVsD/w6NObB6RFE
zJ3HGPuc+xOT9sTTfWe5FJLw5FrZyuwxBjDa7yDHv1pumN4oX7f78XpLrAejFmBt
5/hMlaEMgREnPFX7GGxwc8j9GiVb9162njS8KFzFecjYe/p6mnTeW/qOXg9ywHI8
WvvnF+ulmRXNU/S5R45/jdYqgTATXsCX2h8m8KED2nKXpx2JBKPJwDv66zPIWpO0
DLUzci4EnaerRRsDPOV5W4Y5rjkZtluNRP8w3aeS28VwWXkU+qyb+vcdkrdGp4A2
1zG58whlkBEjRvTOVCxFv6RVmolX2l0JzmUBKQq1X+KxtR6+PyUBFXYWiI7kQxnr
uDHOCIXhMiwTSK8RAp2PIhvgPSnsAXiqfPxVeiEJseSlAekjLl58O/AqIyZn2Vwq
REDvzrXdOuQ3UELt4lO/yIA60l09zq5cVXWglf8yzXewhQZRK6QK3t8E4E91tvUJ
U8EMbGeeV73nW4ZH2eBFp/tFCBXua2nmf7IJtSeZ6lV1Ff8fO/+A/QdNodEPfc7B
jiWHaABZMe5kbmtLJnRc+VpbLcSN87wXNteo1yknVHwTTARo52CQepoc2S2xoPyk
pc/fWdo+gW0gayBwoqGB53mCMTHgQXZ4BaQ70B8JJHnduDFfhi980wKsCXXv8FZG
JiKKvFSKVy0iXdgS4jxjxntWLpY/GaYoEIn/HmTAtybzAPbbYE6G+whNwzvRjasm
dheTQ6CmpS7vSJbiQrIaxzJzvV9Wfi99rZHaCdmdTY1SEoreZhyamc4Wcg3AcL7r
PPHdu/WnRvleTo/mIYEs9WkU1WvnT5FEHvbDP5WcxHhu6xOMr4gkyf0SkC/RIcfk
A70bSxpS7L4aQDAyDhqr53PkEgWHxrQNu3iIUCReeWedG8ll4PvsmIfbM6KnpjNZ
l8dPyVUhl6H1zc6jvecBcrL8x4Zz6FgQzGFQtXdbn9ElISNEwx4E5qhgHIR66K+i
f4rot1Ds3rNo1zx+lzB+OrpyAqVJW1qW2b0V3/1SDXgsSb+1Tpw5yg0ZavEygMPh
oRgDvKaK95JryIw6SXlgYwAPz2dZfKvrjOtc+m4bQ44bZQnzUmjzTgTozBGjZXY+
UWGjxoxQAZknvXwlnNYf3nEjLUuwQnpZUZx9PfKyWpAf88+ek4rafgu8WM7KtC4A
ne8G7bgTT3FtplIhPXLsuA29lHEHHbjhdYIfXm6rLH+rnVgJLc09u9xDDMVbaB6k
WNAVSJafLMZgtjnUwZXbRufQxMvOqhLL+DhKGuwKetR7utfISwmBb+j9FX81C7zz
c8iVp5a/tc1vE1GliCHYcrXO5Wle762fsCxRHh6qajQssmW1rPiOlsDlmGSi4ynq
zoULcq53x382kwvIE4R2KuMHGjdrFUSeeWJFOAcECoL6PMdNSmplzzrtHEJy77tL
sc/HA3INP7nzKnj07udrn6qbkpuVMq7V7gUD7Rp+DKtdFPGIoMqlh6w/X0oOB8oc
mzfaxC6sgteIoGV2f6we7tAytkbDzwnnBky+nRurStgNRzqISqiuqoBEgoAHzBFd
o/m+O7SbgYG5F83pMswpH+XmZBT8zsiuYvX0Ai2SeItE3ac05C7zlEmSdfpjqQSy
d+OSpNjqIGr9e9FkMPeIOlI5PKqzRSSiA48Wkn3A9FF2rLH9RAMrhEV668rqj6oL
GFto/p50FwFO+bihaaeWtfYX15sZjX1uYV6l0MhtKrJrtzVuWmoIL4wf4TbJ0hW5
KHL5Yj+KtY9P0RO2tFoQuhaQfdf+uhj9LC0xGpE8c0atqA1ul6Rkm25ynX1tlFT4
ezgR9aM8o5mQ3LxzMx6hNdZVegy5ATKmdKH0dK2+k3Y/P7B670MqbCtOlvQoY0Qp
Ox05X6Kr4TfhuqjM1QfUyrrA9Xq+1x9i8J88yl7p2E2tIvj+oou25VCr+Kxyl8bv
Sudr67Zwq+Rzdp91N//EaNVufllb2UnHyGndCSDgAPvWsmqHGKsoCLfx8s/n87ix
OHvEsshWiELyxG8DuCN9sLP1kFRjLHgmxAydIG62OfL4Es7yltxTZuf9Cahr59bv
WtYiJdDpeOfeEuXBwAsP6MTtZ7uR6X0zMvFE+bqWvElRbWIp1XlEtrOmRJ4eT2iQ
c/Tj7J9HPGxJhC17VIRQ8bSR8HbDZCf0ujlMObUIYPLxA7lbjDM/sF+5mk1OBEVe
FWCn48c0jWJsfUBWOQ0F3EsZriHb4iWaikhkzMZ/vTOhGWdtRcxm/B60qxs5fVai
nJ88oY+KIacTwiVDIZ1898d587VhphuFviUEFDNANZw/VO5UDazQfj0ChUNwyyaM
JrPtTdTaS+y9130O5HOqDSftUBUFzJEKaRFpy3AAFavL0ZMsYdDfcUXZ5t5Ybk7Y
sJhtgq9ktKij6WI+/ZW+IWLXBXGUwPvc6x1sMK4ICEvGWHkxivPZ1Zq9suAdwK/E
q7EJPL9H6Gk3lgC4Ke8xfHpsTZq9wh96l8c7MgsRqxpDsWNKGhJkFIRG/7cYYXvF
ZUDv/GU5Y62yvLpnj7tR9baRV7RPQXDwIgFGLQoK7YhiywIoaEWayI3pIAzb837Y
WYjnXpoNW285xQgmPaVqm6BDtPQLEPTnsstS6RTacem6Kjg1Cj8xfi2U7/iqmgiC
c7rrJXyOwvwS4hsFd7Ipxey5seFDNDAQAQof0NxDnvoIHau4sZ1gpj30WcbpEJBl
cOliIC0kRUp3l8+UqI/ZFA0DLkVUhtp5GCVfuDGSh5TAAOeulOUJxuyvawLbxCPp
PqgmPUbjHqFFSpxKQyfBlZCrcsm9rwAQIqroWJEkXORqbLIsUBT0o10T2aUonV9X
KMsXbiIB2vk84mB8zpDwNvrhImZe5I2baAp9TJsAOz+wsXiNIObtx+T5Psa0jWQj
BiLH/BV5ulP2ouHZnVt+rNNVRyBkEqjykQCB7Q9k64J3KyYaroKsp9j9DvR0p5ub
/Q6ldCtYrGG5Ct4qgge8Qv1egqmGCKAwbSh82X5MC4NnOaz3YLNxjqkZUdSTCIwL
CVyNOY9lvauUEZZQqlvqBvkGhFRbq+IkTuYmRoR75LI/ti3laJklOw8xMNSCMP4B
ytzrzCN7CWpvRMkm7HTFG1RNtrgnvW+CZvtE/anIAgFSn8dge43Bwrp2P4vDmMjv
iM+tX03wCKKeF25NOHVyVu0TB0j942w7GOYCE4PNSBfLHSJ1Fiy6ifO0txi6CrQm
i1SBu/D7Onc5hpD5RFN/mNs3nWSJumnwkG6H5OsU9TeB3zTmOApkBt4hykWN4aJS
znPMEVJP6Q5esftSxMLy1LWz8icSkXphQ25fEZ68grEq3F2qgTeY0hy/iyM7KfhH
NLqWrtvXXwh6G65KfWUo6YqOYraoE2hE25SWQY4yodm60fLom69jYoqX0ivTcVVf
u8pCamgPWiRrkf4Q/jFbB4pufhktlqzUWDpauJB282R0XXK25RCpTdi/lFH86rU8
lAd1K6STdtmybNVH3QHCel6elKhSOl+XEYcOkI1PHtkadPk79o9EpTPdGvhkwUbb
mxPp1UJ8dccRuxoLiFLsJQBXI5rlcICzO65NrBk+Nk+HodtopXzgERQb5KxNy1Tz
fXsJtyPkBtsSK+k86/ER3WwA9j1uwhc1R0BpGwFNyqpcTSD1foZQGqTE0gecnkfw
estg8BmzD/6lKiin8Ntwk6JpdYAVbFct/9qPGCJEUn/yMlVhAfnP5tFm5/QZPP1S
b/e0GVO6248Rbfr8LamYSIXsxo6t6oKB/PZNJ0lUA//JeoaykxNhXFZ3wOylVqWO
W2zbImYZbsuPWwJcKSnJJesKofn9QOhV1UPfzmuUTCx8fX+I4iLQzvr7BS09utJF
6PQitMo/hSiEJ+T7fr0JbwV1IbDPjAsa2yIzZrOBkbMrETt+VK9G2+LgSrTavhPV
duJyIhO2ZZ7//DL+Jrc0Fa1EQA6L+dw1UAGEoT47KjIJoaLt4Xir8W26uvDLLqY8
/HUlkr+vnf2IBNKuReJIhcfPqKVP+p+Q1EagKJXMz61DH39r++vB4cOOirk2ojfU
IQ9E52QXtEupgXMKifeyNpFFa1Sd86LIRd8LUkq7ec6BytAjl0noya9PAGKkb7jS
kRd07NdHzo1ZVgIijjEqNtIhkzXpLc4HnZFTwdDPOnM5+HHBTRJg1NzU4CggsYaA
UA7CAz0iefxBOUdPQ6cqAOaoQ8UKTtphO6Ub6V+jUGrTrn6l+ORwJKftUG4Er8Jp
w0f6krBm3ZqTqeDBFj3xG/O11rECwPGUI/OEimGKUagKmFu3i13R+yQwj2Kw3i+M
7vcHXzoaOfhDoDsRZ0BlgS1sr1h9LjYkokCEPd0P+QCrWMaa+siYdACM2opSzp+6
poOFdfwrccdKbG+qw/5N76BA2PYvvKkqD/ezWJbKRMimwAFSxOm5c8zgca5dxzcL
hldXI6XYiJEQB6I0n35iXFOVms/2d6G0wRVXFO0jAlct+899fcfLFNUrRxD0DAU/
7DlLqsvFBFP6NgUa20VbuQsry9ju7NGWBNxRQYDvUmQvAqXeYla1hYR45/eB7U/i
8CVqqYH+mWEWBUJeI+J1sKPEPN1GkTJT2s2fMn4DRUsZNGG+ddhvHQyTCxIKldvF
ZywdlfMI5P9wuNtRTSMF4FW16SUz3uLDLERTl932XmOfjV9JEDdKfQVGLohjc+MS
dCy+Ejz3t5cq1nApBh4hfh7tH9o3KLSM6D5ujgzcNacV+UBIAGYH27gf+3QXwiKz
EnPCG04uDSeYHajBaetf7mRlJSXH8stwLImNlinLCqdEqhMO+f7lWE452mKjgdzS
VB670MztZmZvbV2n0A+nvp9W5qXKrSQllf133joctohXJa598MbeaN3neUZklTGX
SMki+KMVojtsSCYWk0Xudq2tgF2qQzawpHzSfu82m1KbWuTQzeGkBOD18+gSFYVM
82ghTFyCFLSuCFRfe0rwHzz5TrUtf1eOU2v03Pk+xqbPhIucDb07CwFjQNai4ocT
t5bh72dZzUaH1VTWwpweRv34xndQe9dS+jxojpsVbVmbisr1cgVtJ0XBTJyfbXr8
O8kzVqedCBYXYf8FhfgDTzYR9HqGvAJX6EN7tsM/0KxiVKPQeNEN6MgKaoVbGIzd
9jTEQlUflOc5+J8aYA9vCffBUPy2GghiCe/liuFs1swDAewJBm9+aK93LP33LtBq
cAatrGBic2+rXDhCXceHJgKLy8eyOgvnan1UGbxDx39j+5t5GAePx4QA3gdOQL7t
JD/G3dvD8wYTl9i28+RPxsM3l+KQ7EzA70GjrAhdkuLYlgnTR/0kxVXwjrDyF4IQ
bazXPMygWwDFvPSDx3Y4phmQFu+e3MQEDEeNE3z5PxOpYAeMAW7W0JKBVYQy7UEl
IgtdF0vq8291PQMShJCEnfZl2EHVNxioldIMmAKPH1YRSXmiPvOOK9PThkbgDgwJ
B+/bXcB72Qia/r7HOdKxLIOl2UGEXdko2Xs2Ca3jAdE1usuHnb78pZ07TClH3LR6
H8Ey4rIw2Et6Jdn/sKp5vZXEqZpVWs2R1VGy7u47pf/x4DeWQROFO/Ka6c8UDQsw
KG3ZohpaAqun/t6Mjdo8ReNVrDdOPrdJF7zs/xTseC+p9fs1qhBqtwrcrLHbPXW9
F13sdKOMAnJnvQVwGZqt3Dxg9PYAlPUlao1dy0f41Q5yTRq6zwRhAoXTZgDAk/DY
HeUCUfunKbXoIg8Mq81mxyPduPFAxxM0GkayLeL89tJ/c/Q1x7VsZwg2xT9QkDug
ZDMiCiiRBc2LWVqxh+cuBVo1j0w4pZIs9BSiP+VElRntndpC45xnp7LKqqqCm/VL
P8W0CXqogjJR+TbbuDTbxAAHq/WKC7QAtZj8GTp0O4k/nSICit7su46UQgU4L/bG
Ncz79HvUm95F/VxyKwc8Jetbh3i6DogWjMJ23S3rr6j6TmYmb0QG8Jz11zoPuBTq
xF8dmHQHYxUMHcq+tOzg9sS9UVDPmhdFtpDDUX772Y65FmmHsNcLeGU46F48GADA
wniTSbl133p+Nv66+LIRtmNjSC8ZzTaIflElownttxWuXuRg87ChKDoy7YfdRVpa
3WI9PHkTaB6F0nVwv+CCxqZqyzMOaKIIJGQR1t9SUnvEawchTkOzUovUXWpaVpOE
Tv1t6uBwC/9Y50BBA0icgjIuDe6WjAwnLQXdpZnKpiIYa0+Sle7LXGbonhY6qiZ4
A2DIy+gPGgqTFdW6fsG3afT3gcezjzlodBX4pQ/tWuay/YWVG+b3DEV6PA3hMz7M
gmJW1QKbXpT4YdGoKhC1z82yLPWYtYkhxJA8zL9qJcGcVD2vG/VgR2Devxc5iUG5
QFEOqVMLH5I2IPwHP1QpVulFRlKx2WO92sXQGwsRVXtRUnYzXyqcUS3obQ0r0u7W
hk3Oe+5H9JsbYTwO3LgJOExWhYx0dBSHVCqyiB5c/BSthXAiQQ5UOdroqYF9oP2K
a4uHkMULU2ToueZTvji2W9UV8rQn7zsileR78/2Z/WHy8rgjK7ebyDWhA7P6nWvi
BTy4l8QmpiFYmSd+U4SeR3dFD9F3TJt4l1oUaZqPMlLKoHhjZG7RJwrC4i5+QMB/
qm9PcoW55bTd7DEoNyczhqieoQSDUOwOVwMdu+vcCwZJhoT8oqnUp4Kw6/imU1NE
XPPhPmhMjZoTjO2CU7lBxuPTmy19b6CDAMcI5mm05mv/JWNNb4p4mTFjn7CXWRDK
nGYyIiLFp6cgVsmG2CXoyqP/YspaJo94HTOgZWivGNflwresoFbHrBJmO0sjEYRb
ltAAtFAOtCoarkscteyxNhQp43PTR7P8vBa72rAQsuhSu11Ec7SEAZLyft8opvMd
Y8mJtvbmp0aAS6K1OCazfwQOJB9CUVcF5rvrgm7NpSXJKxxITsJx10hmdNxXUrbJ
907lrb1rZffufHyI0mz23YOCuIYI7aibpYwc+2IVnDsbYsY/x5xvxXWP6f4b893/
B8GyXj0OIz/0cP2d1W7RruqRBtHio5r4Nwwi/Ham9qYRYBxliAZbG0qmU8FZVElk
TjjZuiXAn0Ltuob92FqClm1a5alo+g8MYZ+5exUwOhd82Yvm77edU50vaw/Une8k
KzH2WSVjXZufMX04Zues71fhuZOyPqnbrxeuA+zBuPvHFZdaSjH5bm42UXUF8e7I
Z3xg+IJpjQlILl4BGkzd2AD7FudHfasjlbp8XT2F49OtWqqJLQ6p1Hbzy+OCBWjh
tIo3A9M41ohfWc+A0UKmlepFxSMN1PuFL15MhDTt7DC5GCSGHfmZQ6XQS4dLAmuk
ZC+jTBRnxShz13u9Ti7OOuSkfIBFYkSIAcnUwNJx/iaCPdJnKiF0+zKTVE1huCka
O2YKf9HJWrjPUqpyziS+QmkD2xoPS8bgsyShmmIUSWJzsBAy16EyXihmMx0H81ww
+th6UGyr2aS3gcf4qeSBcebBNlQjIzwPnm0qxpacKbOf7xUQigv+jed9e285xyEo
qPrrcc+P3Q6dcCnHhbqgNcXhPvGRfq3WWnOQbEdhm2GXtLjx2zBR+hCGcph1fKqk
cPrvfg3vv9Yq/XSVz7Nxo/QTQASu8mpAvJNdm207T2t/IXym+Mluq5i6woFXXlRb
fOITb7oCCUSl2dyWct6wiIaiZCYH5UTCz98o7DGt96EM/8SBtOERcRU0YaWjp789
nZykyFanUIuAU8xnZRnuhaK4XI7zhGv1Oh3yCRVmmy7RtFRbHS8NGTgm9odLAPFE
xQAwMpeyRrlKIHCm0pIKKljD2OBdyYtiIvxgOE3gzxg6dvKeY6yEyQ42QuDQdkLp
vlOL1DdNhRO6yPpOnp/v8vde5DZCAXudJQSvKW/cfcK25KtDDG5dEed5pM2p/Ttf
k1rvRpw6YlMPj55YBojB5K2cw8ikz8sEA7mLX753+uaLqF4Nbr2FpYyaetVBUBYP
HsOBbwcmqbIem7Y307adj8G4slOIlbF2SHq9je4qsHJWYSWj3CBB34xp1ATcTUxw
2bFobljHTfMoY6l/Gx/auEvBENPbGg7SpyB7ZVTHxKdNfW/Llb9T2tvJwzd2vEfY
vawMH59nLk+qWsWNCaH7XMFF8tsBa0iUTk0bTAX1cOgoJ+6iddR5clM5ZsVEaCiC
jnxVXfJ3dWgjeA4VVA3VH29o8vZeRhNxM7DhFFU/1d8rl2r5TQyWSTzejwPJSPWd
GY1/7zECvx0dzGO9GDCLvuTH5QGCWFSWgWQ98Ew1OzjY1XSbr7bdHly0/LdELvzV
kxpcNdWrcmKP0yDx1rX23sJHBzZaNFZ0abU1LuMSDIBnH2dAAHpVVyVlQ/UUtRnT
p4B7i6WbhoS+2Ll3D2MPkoubAq7FEcUYS61pSGNf3/+GzL0oRHMkQrGKP90g4Yog
+dPOS1kubWjD6A/SCAAI9uws+Zu2Pya9OrPS7KdCf3geDiz34LNtiduCR/h4yk2Z
pHWZxgO5ckcK9k96LX8IXQwj3VTBSFUJpmBUTl3uvHAerqvS98z0F/dd1Gijn0M9
cL1TF0TR1VLgmiXGFp9BK0MGPq1sOdtcZIWMoBCnRRisOAfuk3Mn+T4nFHC/7cGb
/FH4pZdpnLYRLM7hnEr+S4nk+c2vXi5+4KiomHvIqm9ObCTiEqgMgFG+cSX5DOFd
q/AAc+NA7vZnMK7EkCFJjwMJAFvnmwp+P+k3y9rxoj0boJY2fdrcr5PK52WhFSrY
KeYBEJQnt5quMC04QPSZXSsngmyxbgqpta2STUtqJlIqr/WYnpqwLLMK2cFnH1aM
qSP4U5s9hb3f2g/YGyUyt7kG6QcPVjUr+o2o+RSL97BzVA+lArPdhPdiD+KsSxSU
RIbNLJju5c228gXUyu3nJgtPTOg60Aiy525Bd9avYQ9KVoDuCg2Q7qpFmbtjaHqB
87vlP1CcSWkiZyeKJpdpgH71JfjBfh1sbstghHqEC64ilsnZ0145gdTbxooBF/8/
SRmPi9MZ4oVO1LAiN0a/GL230zrbgZFjqjFkRYSImcfqF8dxLvFDw9rFVBNxETT4
5BZSFqIGssHibh3Im3n1eA4emKs8KpzTkiLOH/zgP2Va+ALxYSmh4ntvMxYbtMSu
Ct1QpsIDFPgRg3jd9xdLvUNCV1Gqpl4VNkIwYGxNVekRgOuMIt8GGjPDJZcMmm2E
QDJK3aEBHQeczZ2FrbewWB+Xqi0LEWKH8evTmnX17UbCOnEPxp/MFzcyXs+nzPDy
FzEHxg0TEhyLRNi/97kJMJmQdHizAjO1sK95zuk+9gpJecI1hhpoylQg7EBK1jAg
9nY2reWUOo0YdJ2H9tmv2PFfMeH+h3xyWrHP7gkb0SX1uQTyy6X8wYULYkIFJKq+
pynmp5s/VGA9ecSwukWY+V/iN7jfHqojxsNMA7qggqtFwVGTteA1kxTcw+awX6JT
uc331WksTacZm8+y4STrAmIBPvzhSN0s3Bf1EusM3gf0UwuQrs8lgGZnuHJrDxXl
hHRj4GZkVcoL4XyF8d1TtxjuLR3I51ygkGzU2qbq+wBfZjaESTaxmzNd/1ISOnF7
EbS8FGR5Qb0ac+1kULpkVJPAQcKzlk97bZU+12m0zrGdxxP5/GVSVoD8sVX/d68Z
b0UcaYdbAI5P8s2w03Ls+VUHoG32pI5E251djuoOFgrTY36PGS+wdR3b+IH6NHYU
ItqpkpilrizUYS7OtDVQbya5+fK/S+8HEu34TQxCZYI6fFxBVGbhKUe1T9rTo0oK
OGXsj6vS4Wvh5/wYn6viPcQo/JgCj9b77GSTe3w3geRqZmKSopxVDld2WKdgbzT6
/TnnxN5Mjtc+SNSzLTzLcb0XABjUgwaMKiZe/YXhMAwPCkVsrbW8B4KkRu/AegBJ
oF0LHbDQ0LAJq5G1N6HREzm7gvs0rtCdG3KO/Y4+mVkfR0qSG2o9nEn2TGPYx1MO
sYLkl4yVsnIiHRp3AfIOQ7qFy2Icrf94T1okWQhBINzIc+x4jqCdI8qKu67MuvfO
N+5zvHVZl2YnhbHpq1ONzsF6ODW7gfYkETI1jH5HtswgawvyK4dIV/0ealrGY7iv
Mxj2VqbfyooAWCMiZq2pufo1TF0oLIEk8JihMAMi2qXKTefsEiGA2HhWhE+vBzkL
AyPlqc/5vGUHHYd51Rj+dLizC5wapXYhBdqy/wXtZHN9ZxEpaS80KfdZElDoovdJ
R1woifFjI0Vc3nQwWW6n5ullIgciAjO8fcPjFssgLATlpFOihtt3FDjo0XiyfbhQ
r4r6ACzWW7e39OX1nlUFRuj7b9zc5OLDPkfSFQIKTpSqG5qVRidr4Ui2iAUcPAPP
D5qRoczIWAiqa6klmNae0HC53rMo5k/wz+k6/4vOEPF5iOZmoaf0LsUZjUCa5id8
PRniLBiF6kRPiQVYEd7lRYmZN1Wcz04gO17HIiGnKF/QNn63N381h+MZUn1K0+zW
+tnZwHPvzI2j/akWNXTGW7hqgDt7O8EbZ/Pm4NWoiH5yL6KScvpeq5CubA+E94Vk
sLNoIPki5J1mOkAwP9A/aQvRXOPDlXaBRwxX0P2EjnG91AeoVq/yWHVizRhFH+9v
6o5IbUL8ObaJSbMgmDDOj4juKDwxRe0LSAMaX7CvbOFrchZB26UiLBjyMwRiSfU+
GKKUd/elV5c4E2NbWvbCsvaSl9B+x6+DcyJbtOnbiuDKlK8R/RXZy8sawmvB2Zpl
dlvNvQtEqH3amOGHQaYBT2uf8nOYCb5qFx8UZjLgIPGJDgwqBLtJTbwmLp7tcz1b
SI2LY0A5FQWCqsb8WyckdQr+pJNHLn1cX+svBg42YpSTle7jwrBrWRTeDWJu2NYM
+OlpYzPb1OXxpxm28PV1S4bzbp6hF1AuiAF11P0rWXhMF46rm3Vjk3Rnwj1E6zA1
5HTqm7767kIuBfJ1xn1nHPPMp7gE0vnYx4Jhkbm+eOKJQQ0Kbhfx2Fpf4WAZtX5b
4N4iGckq1OJOKqB+h4B06tYcmiOjf9pliKyVY1IS9ZUNyTMFMEhxG5OuFjDuq7kj
mDIj1L/WmzohZ1Op7N6nRKP+PI9zKAQurpnYHtMA9K+VUqdxRVhjP1jivdnRmDA+
3Yj7qOrjxVZZ8PVGyL4x4qGCzULe+StJL/a7mI4wEEXKeE32r4F6HE97rZSMGSr+
ijuF4i74T/FzhpqF8pC8TzmzXGA4ysDCo5pVNVP4eLSOIv7QkqwTSG8p9V69GSAp
OeayV2ZFoYzeF+SCIQSNAqYCwxVoBUtyJZeaoVG25aAFrwiePauutU602mV7zQB8
q5EHSi3nQ+SsB+seEnUFtrVbD8CnmY3IMn6ZIrOkwxPuE6nKbYseJBY8In1DwyWB
OZwIqzEabEASm77sJ2NNC4MYtphuBccKribGl4Ot2ZSn14QNNOSlHoj1paQgnl+C
COoWg45fJRFHc7bIcjSlTXiGmGA4w/qbo96iuDz0hV3E4H2iKLs77mByBegOfLtf
q/1nBVWENar1CGdF3eMawLwHRWDLO65j0JM4bqLIyc9ktPnPSrchzBjPe8+EtJE6
6S3eQ3if+HAcZuYSn8pxqkRxdrG67K/tm5X2u/AlSBlbBriyjaBbX3x2GqeQUQhx
4shfrZQMqky7P8Ayaw7jaVFoYiyMcu0d4x7/aZgiCSLFZVQC/UGUAonHKecC0vhY
w3RCfuhnFVdKKrbsYLyJzdFga0hIMdRKGM3EjOhjQdixL4zSNwcK5x09wdhcbI2p
E54jjiaCZDPPhdcV9pPgFrUim7F39R77ru+hLGANjg2mC98acRqP/KdeKT42bkme
s5n66NR7ptmI92tc51Qlc7M+ygRPiug108y64pENgshlUrTcX0THITsNmHQLdGeY
rdtquvJ3vnYdeAs0te9lWQGmyCBjaL/y/j56VdJfzPHEkH6WAoqJ2M4wNLqjTsTb
nqQKqFAqO1WznV65pPnXHxxsa0+Aml0ZotrncDgZyXCqNq+SRlUH/6qL8Q0uSccd
HoH1UkX8UyExJlmXrm2UlLlWONdhvRFBI4+bkM5TeOVfDABqeyHHEl5LIxlIGeEw
m0p2Ufc9C4aGEJ0+coyyC15M2EzRFy6jz0TIyaXNrO9ffRWCylOwQjCoII3I+2NL
foIal0pR+Jx/6KM/BvvTwno+wIc89ZXCUEHzVg4TyICBlPbauRXavVbMc8ZbRwDI
QA+TO0lIMqPIunHjdF0Dnq5oH/TDhiSmA5aWmPX6aqNCKHFMVlD7DVQ5vNk/c+mn
Z0Vy+wA5lKRUn3b4NFNVMDuiRPzvIvPgJsqPD4NdLIvrP2CKAvM62gdBeroNwkFo
a07R7PuE+r5lZzdYv9ZRmhT4OGVHskfVfLFwRHE5B0l3kDyXvLLiLvNmTGTOQN1L
vM/Ky05/tAr7uwAhRS+vId9S76Hera/aDWvvCvJsY9tvZty6YHTWz9VF9L64ZyOm
FwbsK51rSX+4X5kjJwzvwG7d5xRHw6SttHVt5cc11uf/losCsSC8tg/AR4E8bo1P
mdiVQw6EYk+6xnTBSsHBR9U2fWH/NcWaSUQhQByWbHs+qNhWEqqqQrCXE3hROvoV
2X/dHADGrk9AIX045OEqLOOcurd8I1CyRwlJmLqEm93Z27q55ykVJYJT7fkI226m
on3wg+AOmMSmuizgYBq3el/zJat88pSnTeS4s2RavU7O8+8tq8Ymrd0cA6hUEr1Y
z08CPnvjCFIlTYQalwqeOiZB/2/VKjROxZeHqdbG618y1n0neaDYmiYqmSszji9m
Vkhm/bpXBwIZ/Dba0XwBQh1yguVgq8T7q/Acyr3hFq2quVZLjoCvHS8Xnx4iMEO6
js6AyVRBZwWwgNe7yqU+voD/wrGZLaclsMe4PzSU0hjsMkNPkOF3c8dq33FK3dPR
v27+IxBdLFTRFo9nOlWGwv3cOmWaNdhqeHIzejjOtCwf0CnHhQcctZb9Yk5hIM1b
ZtVBqK3MSeLBXbMGNfws+MpxLz4IJQ+EYV4IXI/v14IpfNDwjBa5DmzT7Cl2nfxv
zYwZ9zhMKz63QjGpmxKRI+JUwrA1lVHzUFOr6iUG6SPdIJvXxt1FcmFJ5t0jG5c7
oMiHXKVJIYGULozPRj/sueJyErvBcua85IIygZW/3n6F/9wKGGR4JV4asm1ewgK8
7HrwQMyLnGLZCTcG640m1mmJJ2VosusItivDl9GyKw9gqqCSj7Va7Z8D/OTtfxdd
nD2QtC4GXlTHbnlSjA9k39tc0Ttlhq4jYN2nUC3teIUnVaUB0QWGqweguu4xujFi
dTCmHzrOxnFkhu7OhDty8qQ78xz3Q8Vr2YjVOq6HrlRuwMb9lCGML1btOdQk2Acp
wVT3zRa7rqM4hvEwjrOKS/n2Mbx8wMRZoBq4LHEkLEnurIAUaANhFlSlON01AmFk
Tzc5MVslObMdfryWS0MOhNr+CDsiCQyJlXOvodA4PCOWnSt0vDvXDgoJuB6Lmj6l
HJvTVO5iyVpEsCZRnaIe+cgMpqd1rTBu+g9+dqiJ5qMxvR2dAnaW5Wy7a2hkHCqK
Sk5N1PtoJTanAiY8bkqnRq+zcDkGGe0S1Mgpi0aTveNnySwoKrtypAck/1HqnuV4
pyC4yAHHqSPircIr2XorCBfn36sBskD6SVeDhQvOGqAAXvX5k6tDKHjQRq1q1d0h
DhtY6VYs+P1QXWUenUvbRp6g50jmrd9Qq4c+8lHkuCMd3jGnf1k11Ebrs/FEGhSo
JaZHIjA4OBhVbthE9RTd1e081HUwqf2BEhQuQOwsNfmLDaaieYU+3vfAR80fDd5w
salN8XGCGVSwy3hT599649+Tv9KXhuLKdLo9R+kayWcKr5ryBKoyBq82pCjHZvvc
BaBlSwzXk//LvqHPrnYncXXVW+52qbVFw3fLtsfId6oO4Xhc4pmxkvdb7PvLsXRN
6qW/JlgAHH584sGivEnNFu2JxXiTzbH0kh22cUA7xD/UmzVGhYaWGlAkiiZmA5eQ
T5b50bv1vx3BBgfpWtPBs43kPRqSjIhCglmofyLZh2tfkSbxiiNdgj45KEYCD+Xc
pYMgLnoJhqYvsy10U1PaMxmXkkrjgLONzel1rENGTtOW54+SPPC5cCPNcbKudMSz
HXjc+0+1B25KZp9HhTUXGpMY/NcTFuHET02WlicdYf4Wwz8p6vwevIqq+x/kRJOO
fHtf/oRdHALUKQzgRNdr8d7MIjPclkW2ovF0cxLz8Cep/VOxw3XuY/Oax80VoB8v
MBn7GACvRRkFyL192tasevEhI2i6nUSzSdbngUZxUR4uj5pPuzJnjz0iebGJu97S
C3GNxMQ6etC4zByrWAALxsIv1UalmOFYa0Dr07BxVelB0BQslQwQEq00FYi/aoMu
VY1CxwfsjeOQvivR/j3JXnxMhLgQjnNq/+wq3ZvPgVW75T0dU5FAJMlz6lt3lozX
bSMGN1uNrMIPnQQMf77QGUlbITUVDsfAJIMWKcFccDKOy9GqlPpRV6YFkpwxPc7m
kkkn6IrNDBTBgXfkhzNtWjseW9Fd9fzrByJtCamEXTWv399KDiJyRD5cjOqW4u5S
Tz7alhq0SFkCOUN2RNID2/6/gZeAGfAOiy0qnozrVpq+XyzSmHYliPfRk2qNW0by
IL8pGrgfKH03EiDHzM78/xObT2Ofwrah7un2byzM/MRrmSp9ak7pFoqYtVmovOek
2K9puUoswqp22UNxTAdBBFqYO5cn8rwHTQV039mNap+Quq4YFeIS7vVLwloFNn63
Ph1gbt1o2pnvHpwryx149JTVJhFdWSktbtva/9ugYLFFgqT7J+8bcoPG+Krp/uAQ
MRVC5Z3Kc15wYuZiCoSp6FdbXoOItv+iyLC6Ya+VJOg91/jM+/53Le8x2urltdrB
6rsJcAoEU+bN5DdZeqZXuKgSJ9/tzNsRMaxlAsAFwRPl417syEa+AxYVMpF3LrlF
lwaV4saNKMyJTSfp03gb7XPSSky4vQJA1koJ/uvaAEP6HWQwNyPYmKRI+/YpaWb/
csRv0lWGLuAs29r5QpEub/hMUqUD7s5wtKFoB5nHJ7EXw1oKFBvsDyC1dlGe4ZW6
tTghk0z/gd1BeRfg1lOkjV2SceN1qcuNq/J3Ulom6paWSZ0NLxuWB5eYWcayQSsz
lal+xSQJfjqa5dr7jgS9DzR2XPp8OEK9GM44LleFl/UVqD7DChgM6Lxm7cSKC4AL
8EsP1DdFeNbHrf0g3RV5lzs08qdOn8PJW6CiuhVRzkWGl8P78NMReJn/JkqjvDlW
R0qK19C+LfRqKAKD7uKRanJ/XI54H3cyI1/GWVqv7drgD6g/SglDJcpHrnn2FxKH
k5IinWa1xUZ/kebVarZaw+zzFYGJE2/SVhgVfsCmR27L/Qg2yq4vEOnJIweu5gO5
uts4HlxUUVJqZ4uoZXXc4uqrDnxHTjdjbrIymdylJYY6VD9XHeg/25kx8dCtvXJr
KUElZXyqkmK2PpbAZhq9zsBgBz+pxvePIMOxGiTtzXwe9MFNEl6b36l5jeh96scd
uiIun30o/jATi4seQKxBQvMKcRnMgsZ64RMGQZ14jcM9bNUQexg4iqDPATsRjVOz
GBv1DfZfspge2LCkPiVs00kTRK/+NB/rLr11Yu5vaL6K1rEXr9Ko+tbYRt7PSYKr
qDm+QsJzMHQGFH5eiLLE6dvs7aOJz544jDc9IjqPjAvVSd/oJalSI9EwwbbgqxI+
zcdETthX4MyRepk6eZ1SPV0KF7Gw+03EWFXLLr3CaoLItZ02Sp/vYx29zm7mYsVR
bXMJqqIPU8vQcylzNBxsgvgDBs9qkJgJMPEXe7V5qmKxriGZKxTSF5ujgchut0NA
v1qEz/U/k2p1cWxqrQ9LIoVFKN8xu9pT5XIHEardMOiCBz1JRNH2UY0R2I5EGI1r
0sP45iBGm1xqTi9Z6H+3lWeBDfPxabjOgmHfnJMmKke1jYIQuRb95eeLyv0oY9Xe
rXRqqiLT0zpTE17+gVXHGpdAJdekTg0JLfEZgeX0bBLNIrVkLvvQJmVHKDQPFnmT
ZYOwwcVL0fOCDCymRICDjyOAe1Dk2XS0g7CEc0tMsaoSITN/5krOzauGnhoN9ngc
s6VkeEdCqb1WI1ZBMiyvrvzYXlHg0kby3dh5koF9A3ocGkBKgYgE5+nKNWVemBWa
xJiPTd/3Tu1mkwhE1o6OB51fOUsA0Wa15BlhEGwdG7n8lyBqXpKUJbJA2FzObPly
AVxdE0Q8S5cVz3eleacQQb40jdCRsPL7vjd3LJlwqIZhsKPq14hxbqmzORjnokuC
0ffb1Eq9Vu9uLFL0LEasfdyPv4wpBZwLFt5Kc1O3Tmzy4tejIVuVhJ4bas1RQPUD
07b4k3aWwXtXOBjVms5hjl3RKsrAuDF4v53XUl/mLUPHVtt3RGpFtOJF5UhDzQZ8
m8c8MR3nX4tYa2ulywWLcTN6jJCxOEEZbLxlzUEOzKiXAJ7qFQ6feAcrRvsKqxS6
UiNDt0zIbFzdIiDOkUQGCd92JhqgJs6/+d1449SGxZefE6wnXMRhmf8nxgdd9uFm
pg5Zuc5+jXiieUYKaXvQ//aMfXJ3LllhAxXoHz3JiQ3MXvn1qlbNi1Y+LDC7Ak4W
QpmwNNMxdGuHd15Lhx92/QaVtl+6IDGpYbc91P7WY4WD4m4qry+6txxu6XWilKXl
Fixkug3wBDMO5X61fyHfYDAp3c6lHtnsLy59jeBwPhjjpBRAUD30iuYP2schFixq
HzuQFZI6JUnOSePELrYS6nwP8vNLxh3zN+mCTtTRflBgFbcdYNbfm/t/d9qt4aKO
rWy+ps1uX3FR3vQFVxHiaCcPjBIZXA8JRv8XXcALxto75ExGTsq25lNmL58deQSA
1Sopth45BEIsZXbv0kAxDlaziMAsOgXWoEYLnyIYc/T/yeZ0rKJiAHUi9jDZqxzN
mniz3ZhDydFjJgG5+rJS6AF2mdHkQRzvRGZv6saSFLQqX/NsOozJiySn9FTgSsJj
9WPaPh4FQ5ajGPHmHwvmIDTEfhGJ75zoPmjhWMvs/Yxxj0Y+pJ6h3UtzHDzL5m8r
4s74kZBBJGF9SL7Htxf0RddIjt18zkISEMjgyCKWHstnMnisDrxZBWzqskPzfkEV
QSMQ4PL47d2kHjwyzUsQx6XJ7iwvmf94CHUyvVUcb5YbB5XmZiH9N+vXIYyT2Oy+
zZt2Zd9FSP5kxn4qWtwpCUjwFKpb8ajjdP+krBFGEmDyvHPXLMria97hrELv51to
OChIsCjPDS1q6yXcMR/huuLHNXdz6CDRRKckcsd6IpXiaQ77PoE7XcTgYIgIgsjk
/Sxd5aGfae5GmDe9gGUC3EgIXVEvbhcTk0RB8387QXGLNrSP02oLU0gD1QYpEoZn
6RDpQmyk5G/pLC8f827eANuLJIeN7vSvDTjcqYqYTaGgkoeaKORJl9g81e24A9Ey
nGaeEnCvb0kT1gLH7LCaoAMhNsqo2OHdo1N+XLA+qWqdl2viO0wLnbODZSvcKii1
tou3kxAh6qbiWqJBepZ29mMHH2Py/z22GoKc6wSc38VI9FPUpDqK27D+5PL1EZ72
bY4CCJ2BIz0AZu9xhH9gPJ0CkPbZrtn/8WMmCHwWGImfXCTqtcwPy2XtnxfFoRk9
oFsDjmkkrKfNggdPH2gBkdA63oc4JPc1JXaNe7ZxSVt9DD7Ayv5DZWrN9fdA2eus
vHXj8CKrLftdm8nb/yGkdgicjffV6g/d28S5wDBuC60yI1Jcyahbqnk3h/lO+oEE
RInEmDhSY2k3vKYIFSDA5ZpToOHV0npZ73ssSOX2NOZBKmhtx5nJ+HzTl7hs2Pij
Nl7kjiCFqYTc5jsxRjX+WBpL4Eksm8hxjLG6qScw7HNA9nQeTPHieBxAmqHF17vL
FyLPHsqvBlMcQoEQmO/PEJOJInySi5orB9QPfmTCDHUj43a/sHUzr2d1A/u3pENs
46JmD2IhEzVEW5/GibvAby6KAKIcGfHBqhwX17kaMwHD/eIVpDB1L8YKpbA3zENo
nuKnmvSMPnwNISE+pi3qCJ71Nl2NiyXO9ri5TiiDZs8wX7Sqw2ch/PuUJd4pgIqN
Y8gw6Utea/3jHYbq5CEy8bq5ZPfn0bF8lbNQ5enCmdbanBzlp8jxHV2ix3JzIBjA
Lf0SMcYZvdAfoUM+WqKdK2/AEaXuvTZcpanRiTm0x0bxJ8CuErFgb0M8SzBKTd9n
Di5mQsi+gqhvYWr5o/jYtgmNCGZT3Sc5o3sOMVP8CSJCe9krqPxBqKbSsSznGgCH
SFvqTc5YmWsEpXekR03EVg5D4ZAOMia5lGKRp8iyEpgiYifhc14wgGtVEbqQfsTt
6E3aJQTobpNADAcLt81O9Ckciqk/6id8Xms4Z43NqW0dhAwN17bmh3rfRlWSXZWW
W4Lzehn7ciiBDSl3Kdr11/CGtf7yAaf6O/Rtaxsl+vhEIDCrxk9WngVD6LIF9hzQ
A8vnFp0UafcKTpJsHOYKHPGVlsmruuJm1QLc+VZeoq+gmurjgdSGcW80gfRoWooh
jGqXG8JVsFP5jkgQky7ZzpzimsExLSkEUqXr4gw7rwch0u/veF/TG5zUGQpagFkV
iaFhotlNzWbvubs6jZp1rLYl6IrWcT+Dd2h8+qkd5PXXyYXwmtrhHoCeDW766kTI
a3Q33SEFSqTv/wIhS1eVurkEUKgpmwBcdFMz+dZVqa6xpAE2UCMH8vIeELDiLGts
QEfDObmb/3STLfjDM/NVCHeTFjxysqad8oh9GVaSvocPn5/6oZv+pjDAXhCD0w0V
BJfxZgFCHJDskqVhhtCM9M0//3sp9jrb7WdICg4TLVhHpd70IleNKpIVq7o4s1Em
sZmx7WA1saoLgQhuINwYDgkW1HqkrD8R4lKgsv2UV3c4xcGb/sUuwcDrCliJkMvv
ftqMA+byn4Y5VhJbbcNkFjcoGl7cBDS4URGa/Z+/xm4SbTY9OFE/uOlT4KH0SCjG
dd45N14VtwJgfZkjhpFVoj5o/tKZx/k4PLGUHSVzc4PqPha1t2WJPL241VpX4e0D
V2fLxrRMLolvbo+7nTI5Q+6v6kDqGPiAe3PJfHAlH38JbD8As4npzcurZZVs7BTX
yYzvdWhWYSqDP87HTpdyFAKFYPS46VT9XO8yCWUBP20Xgn2HiwAMqCDEwzvd3egP
UpRvIk1p3Sh6mpwXmnZffUi16Bzl8HGo1w3AyrSOrJGJ8afqOxI3i9b5F8UFC0ly
M9Frnutio2O61U33KBQ+9AC0By81wLP5tA/qKmnLcYa2ACZrRIEIgeu5S1eiXmvo
Uhw/bpAwXcR1vuNNO1JnNcIWUOA3Jwa4zBlC5mE+GrH0fF0Nb3ZbL/Jtdr+O6rmP
Ep6N4Dc4ywBJXCy3BwSUfA/PCM5r4wQERsD1bE3jtIUgO2Q/O1Qosx34+kVu7CXt
P3UAUT0Awj9pM16zB+2AtQqNSDGeKfMA26XTRfX5zP4L3/8mmvJaymyuv7HRxgSk
kBJIs9oQXrEXv4ieMPdQQWvCT7H32F+aB5C+jVUmCbBvobVDFEF/xmlxDDd611Pp
CrvHcIII90s3YkU9VyE3Y6L1xmOTX+3aia0VfAuQgKjPOTDjj+EL+VfgsKBlL/Qj
FnskN2/zlOWnc8JmlB7F6QEP1F8OEOCEK+oaEhyE1gHg9Qh+ksrFY2u216S2QnyU
jsbspIIqc1/G4rJKqZg5yqotZfbHIClJCSSSAYjwF8yQfNtF4VccxKk0HoLw5adX
VtX6nAs+A32BKWwi/dZOtAiJx8TA0rMV1lhEpY5OJdMTsU8a8/vdXBQMn7RWvOA9
PsZ5Ey+1gCPWKKawMRlonuYwi4Lj2DTFG1BdXMdIz9Z3sMNnAoWXLrh6VtiVoBui
82asAIS7sd3Cs4cjT8F8VDo/v85aNWgMdTM4BdNKrDVVoJrU97N0U+yHgrLxdyke
BwFgusP8RFX53dzoIy6VDcVQLiRsBYO76ZtvKJNCQ/0SogxX8ldgbGXPAmStHtVP
hSWfLqCCYWAgFEbLZqKWV6qmMjfkDO19o8QZ2guaq68T354vIz3w9eo5igfr5srI
lt8hemNUtYCXu6V7GIJ8QmybLGuNChYZiqEJ+Ga0Lg7Xwki+LC+1gKOZaDFgauZ5
aZVxUiry7KpLZI7TuCq0I8ZyX7bZJL+5nlhIwgxDTKCizwSjiWxDzOHieeSccy8Q
G0Hy448+bNbXl+cS2NmNQA7rfI/Fg/HFwjdBSVONViIj13eEUbu+8em8OeWNRUHk
mYwr02ST2azgeJvJ0OmOAMD2naMJ+PY5GY6EzlyDFKeOLTY8fzyw5uvWJihcHK3w
LdNn4oQSs95inuJ5Umum4UHeFIxFb/iovFhsE/YSZJwKZxmNTvlc/iNHmdAW8HLu
AQ8P6ngZ6UmqCIMdvdLxshKGI7IqPLtBMWQXaOT7fOI21gRuJ07mNBjNjcYbHRnU
tsuScfX0S8SpBgnxhjpl4/W0sXMCXheIXK6EtEEynSLZlamPVUinXEokPNiymGsS
RUY646Tgz+QKOpxXwndnH2PmhaY8TqbAoJi5Vuuu5mwOyUa+SG+YfCdR25Eob6dX
IkkshNlxWL2K0XQnOhySivvFfU/Wj+AyBKhzFhXhc2K/3jSdA3RMKZP5IhrDbUF7
qe2dl5eJ1MmRBwe68vi3PDqZbJevkovQ1oilO/dHd/fFLeRhxx+CTq/ivP1NL7+u
7ynJ6LFotxoXnXzIrsR7CaexcixRjrTRCHiwIxHCGRFwELiNMMisLGuuPDy+dHbn
lmhusilL3TbqeKpzRKXIkibZePpiygeKjSu3pgxvA4njPfdM0RI1Wu6yrnzvCkyy
i8b/nXfVji8+Sj/NnGr2xDeZPeQ2omWcw0fOxHWeJ36hnU9yQo52bQIBkdP506Kz
MpduoqHJded85+VC3aVDkNWWBS82IMmEz5feB0P+LLjVkfOsMTX5utXNl5PLe8CK
83ZKI1SfAg3qh80FPKhESRwfi4EoeepLJ01OD9+SPP30GYixxb3KcGGSlX4O+mX9
ogLB2hd2+HHh2xqTQBFbUm6KrD48GA5jEQ+fQwPT+dwqWmzZoY/+eXVJ3VDGAgUw
ZZ9x24FJHwHesQySKLskcIg9hEAo0QJF2ynGCYzMGcCC+8/fHJMvYxsQQ+GzMxdk
gPTc5RSks14V5IhQlnQdYfQTpsmJhzuaavud/3qNPbW3daNMuH/G/pmhq+a2WBzO
p+jwOPG1DJUNiVpXkstAzd33H4a99IbmNsu69aQ2d4YBYni79LSBmnj5EoITI9Rc
GdyJ3XRV1185mUHmlmj2H4imjkP18iGbv8CJhE79yGmMcyUHPsKlmbuwGQkuZsBr
vCypsOhoBcZlUxPPXL/Kf3mqaF7hH1egEW0kERhY8aB6ES6+/+FVFyjfkWLJ61V6
y51spcDAmuDadI/PfDXcmhuRk/GaBxUu0XfDLsm+Ihdog938pBuURQnwjdAd1+Yq
+FTgku3GiaiROWWO3/SWMURYyd70n8jkVVAjBX4KcawRtp2L9y1vyfE+GsF9AAv8
7QcjgVkuFHyuPqEsyHbdsCbpu1w2EgTboxHDkcLI35HxeKyucHBCCu1MzDhJlzlx
5lzwh2Vc6WCngSMcm3WIyLc3Ejyb/m8Cvj8LJvK9b9c50Lpa+FlfFR7hnw00B7Xa
Tu6ARsJkGFq4v8EVRMIoS0glXzUMEJSsPSdK8fs9kQ+kA+yzcVg0GZFBI4W1ERhS
8gOAvTNW5iA0l3C6bYTUERDeM9OfKSgYNFhC66Sv64wt+vjDK7Y7hwmXJa9mrBTo
Pj6Olr+EOS1QXdY/Z8dNTvM4/Tru7PhS+UPqKli9EmuIAfF8k6rocMmAgu65kONY
cUvlXxng0C45rgbyo0yzUdZYJrPa+kr3R50pcHOsLJ9WcFdDwjMpI2OlkGr5pkD9
C+U9qDaKUZaNAUA71CHX2Fu/BW9gJQr9kjhYlHIAvoTLt99kWU0DfrVMQBpJ81V6
hKCGvzV5syAsR2u+yC7O4yBPO4UYDfbUp/2itwafAp2o1o1oXZAc9RqktsxhX3M4
M67OxRzrJQ91qOVWghkFE1/EF5HInlNLSEWKr/QkWcsNaHKHZ2ey9TMMc9XsNWq7
XVOcI679d0QwdHmIOHy2Zt4zPqn0adVkhyDWPi5qW7i+3K55IOimvQ3uR2crswS9
wFXIGdJX2xCCwsw0K40vBoYK1v3Hn/IadXvRX6rhJgAYo60mkDC7pbJabDjpCOuS
ywqZZ0T/lm9mQcOvbvrteK0Dal61WILJuAjdDoX0Wk3OQAr4NgYOtyE7PXNUOpCQ
H/OEZB/mXbormI84DHw4GCQWzOlkrya4Qn1P3hkfwiGOb3XqmZKVkYhWrmaQ6uHb
msbDskbYTUi8GEOrXI/H8FfqbrAX9Ch5n95qhCFF1ZbiuSL6XwPiP+ahVJixPTuv
/AeqNRBFotnmZfNzr53aHxjOtlqB9XzmmtRbcuwnleaoo1talw/Io3yefP308nyQ
j7DNGAxWhd3+jr8HCEYWCuftdooj3ydvzInPGAWUFJZBCvlY5ApO5NQRdqittCkY
CjBTUCDGBXSlpclfMVvIQMp3QVEv1TXgDa3Wl0HDrz3VJZgDWE8SUiNBKmDTMvsg
nYv0pqm7GbnTnI8tMLB5Fhj5265Km7lhbyDXcG/OU5LtOAt+OUj0GkOy9+vF1C5i
6Cht8v4hkfKjguLwPF/586nOdI0jbrilwhocbvvvAGVSL9HUYlG7Tmwtvd/Y+OaD
SVEBEQo+2W0uI2n4cn0qiXEGAFvXx15qeYn6c062uj/Iv0EdrDc/Etf2APwMiyMh
L+Zaz2VPsGNwvctZA0PCUfN28+/pylKgugrx+xYc/wg8UTwl2zxFB0g749PmclQe
KGa4xJ2OT9Hy9aTawAc3D0CfbYawPTxXeWdymBbPzDkcYw+HmfvKm4lZevnUHvt7
VnKp6Xq4PvKLGCgUfgapZ93SNBDHkeKEy4UPf6EWRZ0WyfZcjw/28aAh7iL1yVVH
V8g7CnfnwMtFiFSVhvzfFEBKqcRo5ht4wPjgG/rDKSqxfwR/bunXeijbkwLXl/22
Ts7nq0pwDn8sWxnkhvPhsNdTVezqTEJmUZ6NTJ5UV2QQvivm6O8/yKQuN4KNq341
S6PJJ8Ubiuw4WFi3YJPrNjcJ069e7wg3Us6dYumR0HjEcG/lfCRoQ8xAfv+dGLtA
cM5WIxTYAf29tB3uQkUY8+be7CgyMhHiw/6Gxmdr/9JGGX0SQlROV4wkMC3lUkBr
fCHy1PCaCoSLYFzdecKlUHOKbLa7T3jNgTdSR/urWfWxmijRY/LFUOzecDOlif+9
pZzat9gtp9OPqYL7bMjdwYCSaZuL4qf2njGRLqzB19kPDayTBxF9ozddaC+P5P9/
c0aPCu3ePwyF6TsrtGF2WPnixTcpYCE1/rQZYKdnRwDZo6+Na2FWnqlN4LI6HaeT
V8yLtG0I/TLUw8ndBBPWvtl+QfhWTiUKowGPUmItozLoHPUKYp1xLVD3MvGXCp28
mFdgH3JBdB6i3GiJSDymdmmKl6gt8/hH3ofkgAeU+w6JuI8Rtm3Ch46vh3thhfFf
T+ak1Fy1sd2VFl/3w+TzElcXf4SrjYjBa2GNcwQtk/1Zp7j5qUUGS8sYkrmsPmJt
6rRmrsTgr5wy3bycV6xAg0B7IYI/rC9N9/JowKj4bN0FJeceMFGFmFEQ96J13e3J
FaojL+F3HOLuCPGzjDQD5Z5Y0tXEOOnz0pAbYEx1/Iy6lMUII+K9DgFw785cy2al
OZZN1TXZPwjnBetKOKl7oSnTcrLg3T7XU4kV4hYYFhAqSsrk2M+RGj011W+wIkXT
kIPxUOerNPQvqOGFPXjH0IdJv2sQFqCkvUaiPrbhfTn3gqNW7cWZ0EbqIfQXSldi
x9uOxlLYBCCKcI63RjuRD46vnNz6VzF93DRE3detccGHLNzWvqKrcwGH7cNyk8VI
6ZEeQ3EV/A8J1T4p3ZxYY9n9h4AxOQp/fFSVuhltRgCyA0joYq9XHB5daKtgdmtP
k4/1RqqYov7GwLFsKRYX+iveCU9vxIkyGqGjptPFtiDnikFWUugMSaApWdfPZsgr
ymr6YJQiGiqRgRUKn8Pk5a8V84+zqpX81zRhzV341LGxHW4JGvrD5/OiQI2hudY+
7g6+eicjAnxU6vqYINNwybX2IyVzJHf7k+rs39p2inUdpmRxcJwRCRKDkoSlHtom
SCQOfpC+r05LSmXtJ0+qGHLoLoAyfLUqGz0n5aBfSexZW/mES0pgSbL22QI07W8A
06EJBJLQ8M6RHFWMcKwO/rnC+ztm9wcIG84gmXkWXLv0wxWDSEVYRHiyZe2zRNDc
S1HDvGbqSpJ8+p8lgmoryQaBlhx6GgR3BtsAC3LPBTGDagOHWk0DMeZn/L4JbITD
qUrveFWEMgzk02MxFzegKX+bfNXm2gP9BxWu065s/oU2pKSxo18u5Dr3FQiiPFJi
SHUwlWZJt3fBSVNGw92zpz1K75EUV9HyF2X+MaaHbsEIDFfTuI/v+pC6gMcwLjCV
rbnVSuycVsga6IdOWAu3fd8ifP4SSZ8md7i3iXTDgUjV8CzIzjoRLNbdePlCtvvG
pdXg9cYyYPpxuT+ZXlGN1/2M0QyJJWXIZNMF1e5ZL7bZO09bz5MAYSbVKx1EvWjD
6OjOTBksB3PUVcUivW40lpP1ttwqajG6tm9wvioBFPGi29CyGie/9oKjiaxiIVdK
bx6DmTqScDElHb5gzhLsWpiZIw3yx7u6ne6ljEPwD2tqmzrdCL6ODT8/Ffuo6Dv2
2kPhnvFx3bzWs9Ylzn8Q5mC0rybjZ7kcQoKixryOnzpTEt3d5ACLK8rQOm6alZCx
Q98EhxMOyUR38cBtXMAXUo5KwwuH6jFzLdZ6XOOW5FwrXu633SwtTSxIrZVEW7IK
OmUI8qKg1yBGSddl2IBwQTPddhVhFs8VRAvlY8hvOlq/l1xV0++IZfKR6H3U4i5U
/8P2+5rfvov2y4uGdpvrQiiPU7yUXnnO+ue1WUwbzN+C5YVp7JD1+E5bJOghWfPg
WREgCRLv/aPEbtDwf7iKSBo+SNv+OLfHp5QYCievpDNA/as/8/jd5s1++woAGqd6
393DTIAxQqlaiPrHE7Pcg3/zVkOm655tU9lL0O8QM3bbh7Sf2x/yydicjkl7f2pn
LmFNOmxNDP57Qa3S0oUAatAsFsqv0zFMNtVwCgCSjetkV8gJIZCN3hzXdz8h1OQ2
N8nl7l3AM/IaDv0U23n4MAYeA4A3z+5Oq3kAaFuPOyiLvxLYTJGocg2x0HaIisuL
ijAJwPwW0pdWm5W8xkt79YQZFQy/nX6sGC+Wao6GIx1aYkWMJXNd1+5I6WahcuFf
lBuG5iS8l8HisU8l4g2xu4bL/zcF87dJTaFzzNEsusabSrckg3L162vVl4/cKYrp
BDd4Vk0AFzfjugPKKjQChi7PawrZWDVRIpreBPzKBwcmpr/Ak75PWAII2aULqH+1
NwIuO9eyLjmmuDuOaJZ+vlXGCbmNvqEKqzw9+c+1uoUDTs460y3g7rMO8Ie6WyTz
5m/4EezSeJcTotQ9jVRGIKqq5dLPpRid4InphRHXbnnRJY7gISs6vwvuk6b9jQ2t
IuLidYGljU350eXkBr0XUqeYA/NnLjlWw17KHKNZm91grDH11a544mKR6QvgU2QU
lOfP2It/N2ov+yzO78Wl2Ut77I0gXMw+ubF4QqidPWXLVq3JHNR7CJRfUC4Jn3FQ
2CSCaHONeaIcaECkPtYxVK5tGEyZY+g6t89uQ20hgnPRO1xbcEhOzweWPrbSbtXQ
8ioYYjMoMrFwUFL4Z8nae59rl3vfg2UcecADn8p3hpK9vz1izV+Gyarm6sx3+fro
JLfdRe/WFvJOEGfFCF4EI9lslX5Txa96dMI02Sy+dNE4u6muJMPooPD57pzHcBdE
DbV0aKrfat0wuPl3lWOcHX9HqrrA5u13PdIDFfhE89RHX0UjBFR92UL/ZYNTT/cF
ldVO6HZOiqi60gwXx0wTRdZ2cm3Hdn6Y9osF904W5pyDNK6uM4UskzVaT/tE8tq8
SI4KS6hpxWSdc8JwurgRqYCPsxzaRMoA9cxDtTnnNbvHPsbP2WQuZC9lSBZsr/GA
aSSGo7GqYp5syRAl6weyumFGwGruCQm/vX/BQZ4ct2hSOiPiKU4zXkkQlkh/Ilii
2dlCQxDGeLoETW5hJF1TCIkE0XzXPY+F1bK86JmlC/csrZhonEeDr4d0KgDkafr8
4CI4JqvMPgJaIpkROnWZbS3QIc+qFUL6e6H7fe3lUTCEJQ8TCcNdAMF1DH6Iu0Pu
On06MB8PE24wlROBuxJjKDV86mtjgvs5CQnFuAviC+nTuc4QGAMM4MJv4skgI63Z
yeB15AHi1+jPEmH320ec7/ARMDCNZPz4DCGBL1o1are4MsD00QJRzJnIuvH7gvx5
mYwNXgIvLnj98nhzlFPISUqJ8zFaFpHdGVNP4KEYXyMfYRw6f2UvcvZXx4+Qp7mg
RMfHjb/sKRFoDQZ8ZW/3HnfFNH/yM+kEchKTKADgHyxygCpZoghtUO3Wnut4cwKs
IW1OOnXxn1Hrc6yzJVXe0NRWW/vEwqqv/Vy/JG/MiM5+RDIyZnkeWhVb8WcR321r
lkf/vOecEaDaaA4SdsBdt664EcdBG/hPHUbfv0tt02DZliWub7KTZEdcdG5G4UW5
AUQzpFeQNFO8XP9zVpff2/CAmpbC+ScY5OA0DfcQG3XidfD2l5BbyiexTkzwXCWU
kRpyFTcpN/AsF4/VjcKw+xBNYNw7sSfXalH/h1b8wrcjhR2ycanbrRxhRdb30oAi
17rBwFelT+oIhAyZZdeKRqDMMpGHYJhY/R6tE/E9D5O6eJpXQIdzlXBDT2+ng48Q
QoQz/9zfYRxEMHec5BTwYLbjEAqjtjUDm+FDU1C1039mN6KYgMkoGPmwwVWhHKuk
rmpqci+OPL7xxT0K+kq3hxupIGNmHQaG1vM02SApI3az6Lb6nM1AS8rfQup0tj3i
ESP8KetX5WYsBUAfv97rLBsymWF+klKvQYq4EuDhnK5iUPY97lrPpz2l3vLDLufF
cb6VSnx2bD2sUICpUzKKiCq3gKu7M/nwauSm+jEi/uMZluU8tlZ+OxDlnJKvAtYZ
u7yqz7x5HIA0vzYLx+jsrXzd0SCke8rDJAoiMH1fNUXqWqS9oFfGM0Z/MTtTd80S
NBem0fliQWy2fTmHM50D4kgJlFFc6+oRckj9cQ5gfDSZo7EOOQk6xN1JXlKXXEGP
0tRXAFNX2WqNctL/xJlPZJOWVjuSanrhUogwH6U9Y8Q4TdXymZZNrJzUhLMGtZUF
hIoC9vhQU7YSXFuvZSgkQBviU0j6Z0dO9vvt5Qn5vG0XYh9DeFIGyZDoJhz5kHYV
eDOFaqyeJYpcu51ff2pScQGlG2Uo8rjFPatJ/cfigmRXVR1/IkuSZbrZcLhd9pKw
LUVrMfxiiTZLHVg33OKsdJukkjcBd6P4ULGfUIRcHunfZfyCand1SMZqzMZoq1Jz
YCK4PWGD2t5UjIn2beMbVI0ZsCRVeroIcJarM7h/fquhy8aRjJLD7DHtS53VD4Ph
XfVkLikT1beHc5SIzD6AegIUyaClpL9aGVpK029IvoG6ZdL59R3LP7Y7beu7wiyl
xoFbTDW+wPcFYgCiLcYOFWbQYyUGIxztprArrdSWUNJULo1LOWLmXzj7tBxCPXUT
nl7H2CrCpguENbmbfmkDQZgHw8DvOYXaiJdQYD9FyDFCISVBBExcNAyQuC8tQVK4
3KRG9KT3xhjSJ16C7IzTLmLzasT2O1Q4R1avLGs5QoCTB8/m2Nc7whfn1g3szNrl
qWz2iRctGMktv0JBhRYYyAZa5IGgcg7236vPsI9+24akCogXV6ypvvrqWh8jWDwc
/owCkeXRfahXKpQtTysWpP0IqdrqkiJqU5JK6JgiKvzSYydLRKYTrqD0PY8jCEm+
Lq00C78LUpxIxpR1lOEpqfP411Qt7J6XyA3GAxodIcWEB80pjM/Kr3AdGRVZ0HAK
3x2JNtWf/IobzgRZ89l+Z0IN1w13CdKrWyDckhdOBqn+TuzFgMMmXvFs/TNcErc9
B1YOIEn5s/G1vxbp+VK8T+rRTRP/y6JHxRbvFluPOf82H40rroMxVxE3vhgMv1Lt
hkLo/+/lud516wpORfe5Sr2TjbI7Ad3oV5sE28mjLdnopRuU66x5DBkqhfdWnyAI
Xo3t0xE9g8Hu7yffoFphA/uDBIGGimX4yml2QE9SsvXYobg9PbheyZJe5ukh1TRC
V12FUkRG5ACkHnPMWV3mbv21uBumYwuHlPrq4qVM8vNGmuQosGlX1AE1qCrLr+dc
n9pWckaX3jKYWyHJQSo9CYNTukFznvWZ7SFTzRwTNR6YR3igfdYdmSLX8KrE4o4K
iQ7xQtXk+DW79WUamuvi2jU3hbjCMtA95P6yd1ZcmZn2QwM2wexaGEOqyw11qj7n
VV2zKNJOC4+gms7ucL2oqKxzh28Ui+BkEMG5qBxodS+ftec4hbjT0zP9rokbndKw
gTBl4B5avBnP3ayCkgXzYS0zxC0ZqGk0G8pGhmUL0W/zihyt7CbKfJ+2On3lWVxO
jOJmkO+UDfw9Z1bfKWvPy2lO0XEBCkizLtQERQ7tz/9LOsRSJK/YGVk/cj8l8El5
TpH3uhCIqL9e/s1sAK90/twwu/Cv+ZNXTUZtsi6osgYquOLo4mEvrc6F///G2vb0
68PIKnE1mc8GOW3Mf3AYYg6Dtz5fEWAOE0mlNXU77L/VPASpD3UXB9HgcHWfVvu8
5+6FQ36RWXZtMIfgj0bBC5Pt+dexA9D9M5eAiGcUUr7xqmDP7wsemBS9r/gjHBzM
+OrLi9mbsBDTNuX4UpbYqsi0qKPmLXylbtb+nvVS/uE5oPkMBQyvRkTP7c6oLcV4
+oFlXcT9BCyMNexfNWR6gq7p4TYhjqyROiLyyoONTv+j+ehQV2me7ua/WF5PZ4q0
qPCJ1jRJzAJPbn3FEwG7/3n6olu/jNaaqsQpXi4mt247uDYb3YPx3on4zYyj5cAe
rRaYTCn8uh3PV/CCjM/h5MJCnHri6eAa9BiOiEDFFQ485D4SN46meUYI1aCarPxv
oNK5mF7RoBxFYJikR/1Qm6HDB713/FIq4O+2uimXvDieSfLoXZLvvyROmTzyTqrD
uu0NOGNu2m2sQNwakLIrFINY79XE8+lid0SDHQOUjil5s9TuIQtRX8sgv7n14TAg
RRLnP0f8PtVOHAx397zJt2kJmAZHdrdbs1wBqKZQPDLDAfmKBRVXBP0CzXuybuzY
nn3kDetyWJtgHfzCMuI/2fRdoTIq0HReQnnSmB1PKzJ/ouYUasUFs6+VrShqiAps
iZJtHUIcFFVE33qQqTydIYd5WtZ2lby1k34LKFmFUEyS8IWQF9/4+Lx54p3+X1E5
Qf6GMY2m8iqwujV3DWMoCjVVLXCnC6LHLhM43BwYiWZgsMHZ1mpvrgq34ZJd/fMv
Icwj1w7ehVhNyYqXb0pvkX5i522HErr2BHV+K9XOmJRdfjE0N8U6CtNh4HunVpLZ
DRNx1F++JUo3Jxlz3S3Ogcd9Z6pbiJUDD7ue8csFcWbdhRGWWXLzEBgtrsdj4uJ4
eIZ4zjMm0bbWW8O3vlTkGrUIRdWS6Inbm7RtsoFrYUmD1h/N6jksB+GpvAX95C0M
TRymCi0rqK5nKJ6yhryBPoFV9RXv5+lYH89tkwLOuE7kdeAsyaVEAa7XX4A/+0pA
3/FAyZpMhdtMOPZ2yTv5JsYGl/36L5JYYGh31u4TqxvQaR+Gmmwxcl/os66UAQB/
gRXIIyqD7TeGkGSnsmr5iHlAXtY2/mfqSOJCcaRCS9H3dkNjJA0/o6B/wB+jvgun
IIEsjHrcTHalL+lYH9aH/R6SxDOjlNbFFrreb8aswNw9fMRlyKCg8dFO0tc/x+pq
I3lXQT/Hyt6lfz4COpE/1pk8rHzIlshLzi0VeOru+vV6MzUBHb8IeWPUENoIfqyV
jq5lJHlD5UeEbxuYfx8DypvNvKSHs8qlhKUjFZMhMXoi2wVAVKsHw9rPZAGLJmpK
xa1J6ALvcfhhGENjMHwLp1vah1du0NuvM2rZuAkNc84o7F4/HiqUEO2wu1YOG3qk
o8ldJ4h4ibcQNGVx4qQLz4XCRO9G0kq3fJCH7kRE3ui7hpHGW84Tkr4adimDPjUG
X17Uo6L9uE5pHiSTGei1xBpttczynGEPFWWbjxbfkyzh/SGtnKTk/cFV5HgHfDxh
NZAoaKkr8+lnaojmnpQtvw2nSySzja0iZUQeA3w0QKAWcDxiZMSLVRg3tvj3GWFV
4TnycYRmiOB2ouW4J7GqVWLfonaUGdTKSAXPkpKPHa1M+o82QOG6vqhgsBaXeh7X
dp2v5cxG9trYd2XXVQvA3mAub6MjX9UzFtZbAyOor4I4dyTefIZIqCCeb2kmAh09
u4YcLxEsK8CZ2vQ7Z2bSw5ewwu3gdoUk/1NKa0pU2D1Ih2HVzKwMmqtxlvfIaA2Y
64nziIL7M6G3O6WDB5h6zIgQSug1canT558bdVzEYqaAt1BsiqLR5KSqB2Fk0One
kGjpsVOLfJv2Qk13SbmfOuN3u8+D0x97J0Rg17rFDgbHojDQaLG2YTerJPoMTt2K
CTQY/oh/g5PDRmNMcYPX8I/NKhMY5K6QgdB6HLhGQKuuRi6kuZjn17jLUEOIUpa3
m5i1oqTKQq1HFSA93m23bbA0wYDto1BNiFU7dkJQYtxYQVcDQvR7PS/ZEK9rNN1K
AGhE8mXJq2tH/NJC3qd6FrFOSwCboIvO8M3ZlILgk4UCBHdyYGv1oE3dubeHLVxd
MwyoL6mETTbz7frBCNyewdvAA+M+zVOaHiySu/GxLf+GVIhPeelU9/+Crfl04+sX
hO5E5doWbIVkH2zM6KSYkocWc5fzq7qntueprJ9mw8HZ/sslVPsPN0qw37bMPiUR
OX/yY+aaFokxBeZsZLN19rsRPMqKscyEiR4kfoOqxxkrAV4A7+GUc9jI/ihIJI8X
MqJAY2t5dshyfuhc8cuJLUDQrw8K+OO+ZHBow56zW+kEKIrApRPFbGd1Q7X0L772
GydElQ4virZPPsqDwz1XTf+O8IdNYBVjtIQwncWGa8Be91fQdpdGVawYMQ2AClBK
ttA8MasgH4KNP6ElHYWJ4o+u9/NwDizsiqSXwXbLRxYsDB/EX81bP7UuGpm7p/sA
Qi7+rv4ZQR9zOupMVonTZ4M9NQHzX5e8YcIHg0B14TVJt9EvhcWn/3Z2yExy4Bh9
S2YYSV1szVxwseOxSFflYSsYHxwoiVQBOimDAojj5MX1ptwuxrd8BlSm+5C4/KMY
8GWvpOo98bD0rx10aS4xd9c9p2F2/OKeZB3mRCpBnFysklKtCVTYHJmubREvGF6W
LnjjbBSilWsATXDSz+wTrB/bYzZ2WyBdCVc7C2ErF0uh9WBZQ1rHvSbTnu0DwElB
lk9Jkq7s28XVbcSziaohgHnrr4TL50o73ecIjnFBZjq/P9mYAgcHEes53faDGaK4
zz8q/hrSfPvvJ3Oys4g0M46U6NulTa6pEc4wtwDFcksYI1Y05kz8LCs+LlL244Ox
KZO71HzU+8kb1+k1D9LuGlvnRRpU0H/tRFLP+nDpiY/XYmt8vhZE2QpunWSNUmhP
vgTTgGihO1V9TtEWh4w40hIESDYOVJ9RHX7KzBLalZunxdzSjtjUWLEQyzflxgDv
LhyJ8wwsMf+COLshairFERR2QAVNVnufeO29yXGQEpa6z97TszJ4Y4m4l7NWpUay
aqgdaKGPVdnrhdB5oRXkXzds3kWaeoVQ6pkSOaYyVeoiuzlVi+gqPtO1bNOEYIJm
jIIXese6tKh7j8C69RKouBR9SR/XNLIYULhqkMQT0wlHNsy7y2eWKAEQ2QsOTeld
GCJpjqNpFDMm4qjQErK7jhlXGbDAd9uacfkHrn/djml8dAdkHMxgU2hKOUbmuwTk
yL2B6d3jaVcS83r3f3jJkFjdZ+/i5ZA8KbcERQSwPCOtuEKFj5D9J+jupSUT1hp6
MeaPxayzYXf6y6XWvSAx74rNfGKpB+lYCw/uRbwuDAFtXEpeFlMEXNleSU9LDXNS
2mBdNnwJw1LfqIIdeuWnnY1H/rZ6/aTfPDVwU4Go3EGD849hpZbrjCGUdPmBmos1
lUZ/mbV1w8pOuzWO2dTNZazampbyhwE6SymlBE6uxW7ioulS+25EVqOAqzKn7cZx
imj805ANktJYSpa5JHYd5pYz7EJ+rYYkUB5Ni/sagTZFbgMzVspGxGkCJv7tXk+i
AVaKD7IFI+XchnNBQUZU7ICu02dQPpMJLtiFgK2okF+WgxLT+Ec9pXZr/n4BFt+0
mTp8PdtnMrzjwTi/NLsXW3JXODomOAhbwyXPPcHRbxfJQInRXktd4KF6SREZnKaJ
f1OL553d+qDMVMgMCJQRdOMk2GWfaUfTKo9u9eGT3eSIHt4SMLyt8reqSsMWQ+o5
t09zvRnAsDglJHQYq49NrZcSEVuiKXH4Z+PvrUsTapdEKm4rT/n71RNm2tCLvEP6
thhy6HsuikcxDu3hHNL4UPh8ykMWkMbnqXEzWzoH695FjmRfQhm8R72T+DQYxBoM
A28vCe9semu5y9zYIu8qYLwP1dBVsJaE7pQjFPFEISi8iGo6htlmU/rkMkx5ZowT
FdqtqhixzrrhHA2tlYCZcTEW/yFbH0qn531rfxzhkBjPb3mT7X3wouvMT41LRsYX
djjBHglJhy6dxzTVLI+eQL1VBnI1ACwJPmxmoBN/50QQCet+1TKXlpRos4m1Ruf3
HUq3zA7Dt2KamRVl0oFDzjEBlUulMyLM4XJNM+LFWlEorzKvciJ41lVVfgghacRb
S0ObeSkwngjwvKZ9R9cpALfWjU95zQJG+Q3kyLD1f+8FTCss9CangL6u16feH45v
9YZuKwPAeas+yKWad/Zgatip0tNQq2eYNWeVRRfrMqdJ0ilxRj39L2UKGWk697U1
IO4kw04QygRtt4KsBR3QcDhttzWD+xxEY73oYHwUOtvxllFh8sCoNdcwZtmkeufx
fOcxjv4FWl5YogByIgZIWPU5MloyNXfPP1O0aWGwESPgl/4QKUhhjQ1TJMU4liPi
o+IuwkAN9Myx6mlJpixMRW9kjwbOIaKxHIJxPOFQtrezdd0p38wXQh8rr8tXiC7G
vJz1zJfmknZ2pBfSz9wAH3fg3jlJGnUkbKI6jsQjQuUIc76aXo72iyfJnQWg5N4c
WOedNgSh0Rfvn4vVFEmFB9xZlYwoyiogMZxJ/h4G1OxQlj48TFTlcIEf5wPwM8F6
9U/G7IgsRYb/F6Bi5RbK8wojKf7J7E0P+s6E3hosZjAHnFADu8qp8+x7kctH2C4c
K3+iA6HueU7HX6OritVyHNtHPn1PiZNkScYawYPI59mGjyG5ae6lqEArcRwyYxSB
hYoKj1vJJ69Lofm1Owtz9M2O65YdS1PkGpOtppMdUZ3Nraco3NoFXkXsOGYmcg51
SscSwShbCmn4JanXXE2h/2uVpPrviIsPoDZvCwcU5wVttwACIr6gIIHwrqoIeMtd
j5mt1Qcr0nydK+s1iWiDergmxbm40NMJKgGQcgQlZpZYGeHQ/zKXYoI3M4FEWbc4
4jRHZiC2Gd9+2C9hGfEHCjGSSBh8hPx1vj1RAdEnwa2gWODTG8BfsxerlyGKyPbT
3BZTiG8ut+LBdyFW4nNkzaR00DvDVCwaUQBYhiVfI4B+qIl+RdcF0tSShw7XrVsb
TxT89uaw745AhBPiD2B6ZQ3iJJfu9Tr/bkqbsUm2jqOk4hMWdrVE+MPFrqKv32po
YLPfpvp5YoGQpgRgzz7qXFoYo6iP7Sbfymn7ZswXERoMuLpXI1lkXVrmzU2dnW7h
8inIHb5d6Z2maNENQft0H6/RtItktV62XLgZvoXCVRD1u6kNV608DEkMykZwh2DF
ChogxnBEhcr3ir0tutdEVS8aA7G1lgS+qOM5Jp0Te5jpEy9LNys6TiLW6j/IHw7z
vlbu8WtN5IDlVvtJK9WUKJuB0dR+sNIMyo3uVLWfC+Qtav6cvvredW91FMSQFNw7
xdruujrKbmEyBzOBURv1hbc1EEehesmFPEUxd863uRUCVt3wpekhzl+j+/7YVNBQ
feP1aWPvIXExPIyjaXvJ1OmXwqwim2Hgva8DjW0n+uDID+TxBVFcnpgAQ39v4yDy
FOMeGxgTshrNQPnaPeiFWCQCt2wBt3IzIxffpyqROHkeKQH+4bI8atks1Fvd6/Sf
D/FfRRBSCALIANZKTbGpY+L/Akp0jw+mNh+era+e0bVnNMWiquDUwjzmt8gnwiMP
n+gbepIL+99kXF9dCDXqHCLGxgl5ukZ7ANSV0mvR7ww8hzE5WTc1D4PoxOcUvX8m
oygAJ/Ov6gMsoRw29BxMRYmAtNGQnJdmBuEnY1XIL68SYUV75nyrh0pqSgJZvsd6
PMknftcL2UhgweGzERs3M/o7JJGDWtzbdHn890VfeTlAsF8Q55btsRatBKee9XYQ
ix9bzUBGmZ1XoSwHhG01uAlKJxHKqmmMOmd52kNS80QjPxHpv16y4a9ymLbiy7Zq
wPAup/DNV3CaGEwSI+z7IiQq7ybj1zGa29fVn1k1Lkn25P7kzoyLmobnbPna0Cmp
lTRIVAlrFdlCHyxmxB/LXXH6l07aF4wV8QOhhbrWLY+RKayot/9mGpu9ITF9Lzs7
O/HRPVpB/bIcDDue9wOjqlgDAt/dmsW8OpOWduprGfOtzPBbehMHnfC9Y914kNNl
I+yo+ayT6hh15fjs2fp5P0S+IY//98exr5OD9/QpFvPRytOJck70HQZ3gl/rMiBm
ViNwa4ZLjPHDCO5CqSOIbUPGrQUyIJyYNSSfXXOc292SWlZCDq3/suOfcvTK3eU0
hWPP53FnGtMnZ6avsK7jqp1i6Ms4iF788HlUxBivCKdleSXMkBBM8xPPQILjBEWr
Bz6hYDtPWs97MQ0aSEiJltPnYc5VXjfsQtN4zLhfDhAWzaiJV6xYyBAfKtnqUj/o
wfFcG5j8ijaSvY/AblLV3qZfdiKUsE9T7NamDi419nPzBp4/AWdqvtWQS8YXQTv1
+tObz+/wBeujc/t+hBcI16N8/AqGYBCHUrC/MqJDvER0egJH7zSZVdKGBhPtoGH2
THhdtoAROqddyf3W/Sb87dDG34jvozzLtvxk3MmBw5FJCq0q5FK39pugZBPp4REv
Y45n09w/mS11Wolr975P44G556pzKB0K45QB0VcG+YNCYQHmfG6n6Q9hm3MhAX8c
oyPfvshNS1k0LGEsyH9f+iGCxFzk5mpGrkG+UtunUIJxCVYfQcCWMOsyUR/+m/2R
UfwLXIhXxrcyi6ootgx/iLv50wRrb/iPtIqQ9qmAU1t7dLl0s5xJrRFMGeHaUZdo
aMHEtCindenCSRxDYrT3U5VgsNdUl3n8fuFsATZVdnFCRfv4ndT1mTSMu2pWBY4Q
tcqrP0WRugEhGG/dm4U4ai+fCjzMT1ufoFH9N1/fnv6LuvX7F8ecnBHRqdFVSsKo
1ETe610jDcajmxDdtkdEexy+k5L7eRBHExBsxN77O6ihwnw97Kf5nf35B5p0zlo2
AGQghY+SD74TUTVRXgoP9PIzh19kQFWfSsILMxiCL1guoTDFHcURkn7ZbJzHJqvf
2WUSOC70we38TVFts7U9VM/Oq88IkkC7Y/qTnkRHB/a+MvH1rxjMLovSq+Jaw2HB
vuPF+INr3HoKX9MQpW1aiOii4tQ/9+Fbt32NjZVghAGGRXL+HbFUsj2m36YbfbCF
L0LhSw6eu7Z2iIb/BxDxPGuEOHG0RyEKecZsYKDqvMUp6eoligk/T5ODRUNxTo8h
zphzEZ59gJ/CJ5iQqQdxGh3U9rtV+uiN3It43FpL5R+QOz9RZUqIH/2DxXkwMiTS
PDluq+mGWIYgciyT4H2cNbfHqhK2LW4MfSLVzIpqNg47E5CguCKgq4PaIR1K+HlB
3DOknUQy5EYIr7yd8FXCTdRyzqoMdnEMOzDov+SeFKM5soEab/kryR68WdFkWic5
GBVjWuCrJMMoYgCdwt55WRw+jIU4sL+H1xvezkDt5EizjOwJ1wEHJGsJFgnTXKHU
gZPuDRhUeibBmHmYhq2CwhyGTn18jO3mLo9mXV3u4jfPhWdfea5lMGXEcTbaQn0d
XMgyQp/GISzcnnDSiub6xH9F/y0vdSkiOL2ckwqTVQS63TN5wcD/KiYP4Cr7QvXw
Rd9HEmIwjkwl7z5FDLKkUS4C1TBjAr4Cw/nVwVW3pYZq8gzVNN/0Vtl2YqAzMDyY
Tn1Ed/SmUM03Kf7hxZE3Ya8Jlvv0QAAsbmtvj/tEaoxxhSwWNBlqaPyJT2dBBC5a
5Z7ASaLmNczceCEmR7iw/hmHN48juY44ShdqrzL83GZ+SfnhbJIg7ZirbvLDtu9P
+JglakMg9jnhvRoXWidR9kUpRn0AoLpOYC8P+sYfJW4VKxvBcJqWHc0Q4xcshE8H
NtGjWozjge0OzUDv/oG2+EwlXg7jYsV0Q41ceSHQpnbVgsAgqFNDJLoQCAgS0jId
bWl5lErqnBdRZNCtG5WHe+hICW2Q7ExhehO8HqhKQu8QvTXAM5JpMM6eVyMfeMNA
30quAb0QtjV7AMG9XQ3/0t5ibopLHAFpEJpRnU3FYyJQOjbkEP4q94jwllrcyLYT
Anl3Ka04g+3GJjfAMqZHLeoGRUgZS65lFBD64GooFYNcx7SwjK94JII3skAZIBTi
+EUS3zGG7jNMD+cP/4pXMJgimoeJrRMF8frLXJlH5kVrrMZG/i6QXA7V/leqyIOo
1qWwm5Jvvq6YZNepjv2Q6Fk7VESzWvi+wmOP0aAqxZYshNO0WP0fARFs3FGX7ahD
jEQ7YH/Yxx934vYw5/n6IirJ3cLoR2tme6OpsLd+DVoqPNxTC3k/ki/+jAZNegRW
QjZkhBJAFljvddWmaiRJFVxkQBWjI2qkRYtr2He1wFhNk68HGOIg4Dd9sdpBunF0
fgs6K0quKxzii8tEM2BO+FGmtRBGBFwVgKgS3pdRUMSMNHKbl52PPHOt2w7+7exz
AoER8AJENLu+MwAVd7h9NZDvRu+a+IHjXFNu4p27rg0s9fAWUWxRlDzu7OgBOtBD
O6CxpbgpIVq01n2KcMUxakY08fGjffOxwEIGkQR9MstWxypvQOM8afIsKdEAXmiR
HC7vkwBfgq8aOi1FaY+GcIpbYL8Kl+YKBvD3C/Rq2F001Bw29X/fhfw3VsaYYnRf
erv0XcA1k7guQ+Snz6hm7kGbVpDkbQK4bDv7x8kPxLbiIvOWboLJoLCbYTgwSFJJ
ddCetvgZwbEEBnml5S0cN/cJSrZZnbHDttDc/VSDCuKn+ESRbBucDZFU+DfFB7uu
0lNahh+6dto3mu8Q9AnKMthxbHTV0I308VTh5qWUFElbphdij+QayzhGeu98bm5R
g8NG2X3PwOgI+I8zr77hPDOijtTzMWB22S3Om6AQM7kY5iv4fDVF7Lnmu7Ke/WHU
xQG5wmxO+dUju3JcEB0unhWlPogkiBQCmR6NzINMwpfAfv7wIzgEDSBUDE8jfuKL
2ibgAC72COvGe38uAz0rhJ7TyGSriwyOKKVLF3PmdErzf3gt8vts8SHySkV6vZPO
bkev7r/Ntjms7/QOwlKXtnWxhXax0WcMqt9v+1recbrlFoZy4jSkUfD02bssACBD
E8WAUHYK0FaapB8vmZvxw6vS+044G865x+9yBroTq3cgkbNbn47KY5gqOADrfzUh
4pPcly4jt86RC/ag04jRmbOY55RbvmTaV1Phk9f/IU1uGZTvB8+DtplnfNBppvEC
+iHTcp714qStBSGdsCyP+zP+TbtNM6OfLjgcERPrpjBPNdFDpfRmCR8ePGQdZkPm
C9QioYtVIAxzIKxd5jI05ZQcczIKCdj9ECR6P8bQ+AgMxyTMknh4eKemdY97DPin
ogumRvI9ssKKLVjdYhGXSFLvAcGy9aUHHxkLxTd0pdKQKGAv55oOO7A+nHbzDyDU
yM0nHUIOf81tmt4PvqmxcVXIPYrdDQOClQ8NV9F0oM1N+RM4CdQY0jXKEnJA8OE8
adCNUk5q3/MH+l/lDpQQe78ZA/uja50wUjDzqMNTfzfQzZdLEC59H1qrDMlDAnPd
gkm4zf4N/jdDzU+kIKdeqqxIaUvHvNJz3GT/lshqfp8tNpdqWRiSirW1q3dJXWnK
zVLnJim3OX2FsWB/+LZGalc/olOU56tcBLvD429lNd99td51BwRZXwRzd1ZJ0uyN
YUZDNTuGBrela1iOlwCc/WL9SNB5L7JaZreKsFYwDyt4ckQLKfqlmrwvU5iuyqtU
56y6feinzm+n+QdzHZ0WKOBgBaXSsZ5rCc1uqiaz/5iwRLfl1db94ootUjGg7qP2
2HpGS8PLe0q4mmv+Us84YYEVcDhd6uNI+WK3EzkFLhPpjHoJ43uFxeEv2eoFCo4Y
RCCi+o10VvKl4HoIgP8mNE50SCav2pzb/OMHwBPTRuDKVfBb5URKiulxWdem6FFm
kN/XhsSyjOV0eIy7GG3doUHmjyn4iWfZ8cb8r7nMnWUcg/Jnpbkh0DPo890LKOe0
mR+vUyDuE9HDSrdVbAtw9AzQNq4RpaBvQDZKL0LdkwiQQ08MNnYHimwXirNzO8sP
fIS1kYWfyihDYgGbOYf2WyNt4huwn9IAyjpviSZLCkGCF59dhLcTCGAiZEqyCOLN
NFJFbLZzdlYA+wSYjPVXnvd7HzuA7WOG4OGh+N5uipgmVDCYb8LoESZkHU25MdhU
XMFGlh34mio7YGjQDKJEXNOQGZ6u24ZyMMyRhFgPDDjoZojLMt2yIPIr5O66MMN+
WOyL+73wXFZLjmAUMl6GWkON2x6sKsMFyvvg3ezECxzMmgl5RV+KVlhto8apc0M0
4XKZlZBsy2je2SFgm2GwgFP+NJlQT2pOhsV/d5mYJBEFnGnx3AjrpYyQ5tDQNTAS
+3VVjEvLdgZDBS3DW/ia7PyTkQ8OtImf8DTAaaoNsv5IirG+Bkd5ggkmYMbupqNy
5HpWK9QP+ckzDLtfcbAPS03BUWMrOdNMt6L7lnd8ZFxYF5hmKT9tBurt4Cwo0Qc8
27f2vfvaZfXwDKyoVrIG+5HcKPrbQxlJsmyP6HSvwX3bENNdAeotAKRW+gqOTO+q
ZfdZbLU8oz8ZUMYnbNNCQSFqDT4qfwVzugYImtnn6E9nxnBtP9olBsDt88XptIEu
zs4GKvoMvyzWUw9BHBDFITZGMexWPz08RqRtQSSUb4Gco+yF7wtxLuEAZ9RnUaOY
WN7t3BLrtsuRfSXBIn8o5zmgkQ3mwDSjIx1Q/fwE54aKTpMIqkD9C+asCZO8bRmW
diLzeji/BAoVnXjaftHRTzFHioZt/o6WaFghu1/3S5FdsBt1FCSMLQCvvq5vkLgT
U5OGozNECnsXUFbZwRUzPRcCoFwEM66o77oYdK6hLwKcQETpe/Z8X8TGxu9/hIwW
U0XmPxw9+Av6dQJYxXKl6sSom7ORgOqHrcop/KhH8cWYExXAl9BRuXTqpB6Xzhve
nSUy8dm5/L8sEuAi95TZSKEh3ggZWAVkUcqnN0Bj0c8zbK2ZRZcmJZ527JWOl5TC
ycLBJjVE0svEoVGrM9ZzN7FxFJ08zaZwsmPsrsHXMRk8ZtRzf1DklahXdUPfrNIR
YUFYTRVBP8XG6wDwArWthzh5j/XrImCHeZ3VetUQr2lk1dDC5mVdGpdLlnMmxDKu
zYCS9B1e4i8CT46uTfU455wVZzlaeXIDs2NLdFE3m7vGwkEDMdQH1X/HoqWvml35
Xf5QdBl3RL3BdxixATyYKeMIeiJJmBl4jhcHvmwMc8OIwNm1z5QyPS1beG5Lh4u0
qbEY/K6pnpQ6eHflCppwlCPGfH8+I3FmRkDo2oiPerW6/EKRi0QpHruC0YBpOshO
f3R5t3Geo4y4D792wgLrNiqxVLCAujpc5pY3+m+huzZsWsaQrrZpa9k0S8YPSpd8
EpIfQBnGFxMqX8eMgmLSq2q8H1DGM2MX5D6qVTKNl0+UlYfRIvr2jmIhUfF7fhyg
H7VWyzHft+SB+zQkpkd8upPn9RCpkdYhS3m89Gylf8PQqkn5KbEjf4qXr8XJDjq+
2cgeyVRzDx+dZ0EQUVsNpgTqRUKaOGoN/g3lWYxsdRs+JzPfsSJXq+pQS/YZeoC2
g1tMpB7LpuxsRNoxNsWr4pAIWH9kiJ7IQvyzi+c7mbyv9XsPBXxar2RRO7qNmv6M
S/5VF6II+gXDX9npTdDC6Cps6fit5BHROW9B/2/Q+GZ8RLWorwwkMAut9ZEWo29s
Gv9SRO3Ql2GbJPA+IMPMQKNCW/esi8bXicBx2yBj2lThs9tcNUUBES2F2agLtqQI
Ank7UkOtUhewG+o1ij/tFUZCv4WdHlkqLATbAAhv6hZTyQm7MtAmhHrX500QXvmG
vwj2Lqvz6AGuhLoHKjdXSDKO7QNfXrVVpxPIkDYXbzVu/qDyOUuX8tn/kuYDWulA
un4aCpUxymE3Dtoa7eYLox7apMk855NC1qOOeMc7wo7ROr5jF+tTVBuiFda7YiSV
jk59aRdfWNKyHdUV2LMUeCnHXhqT2LgVxTNgYdjULoi0BPx3SSIdk4nMDVbDLDyS
X/G8GOJIZHZp1nnUcSUeCHdKWkNk7z4mJwi4uUdAvGJ2C5ZJUtPVXXnpjN7HwoMM
ftH/9cS0jMB4gmp/u0cU55O4wTGWcSE2/P0oVLLnY6FaaZOXDILvoc36MYK8irbk
94XLBwk7O3YkUw6DeBKJmu1HX6I1fgWHNEl+G2QKShk3xD5HzfSoi+mV3uxjGICz
ozksia1GjLZfuDw6Suf2RWqlwIzQWOctjh566kKmC7Fb/QqS/yRv/K7qUObDMrIi
opfMP6kIvi6FvKvhvG7Tu6n2hbg8i6CSdky1B9EHp8qdh762L2ICOFVI4s7YVGQX
BSdOp2mrp85PBuT1iF8+tmQBK8kDDs1OlWAi2txv4XWCh+3jqlmrx709q1fZee/6
IZ7W+2d4oVviyf0ECecWkfCxLh4zUmSJ0cDfemsgXFxHZ82+H9UXsADIJGNhRXAN
LHXf0NKpEsbxIBNCa2n+3fFLeE6+yQ6TKbnASQZt63uZGKZY9NsL5KN72wPuV/JV
iwxP1KK2Ui+i/eJTNN4i5IBVh655FYSycyxVSMBYfndHak69/UfM57ifVnHhrPYA
hUjv6QjqoALu4xglzXlfqqsLWKLwSvcP+QapQggztFLsirq+sR6/RN6KucTb/pC2
DvVLjdF9wR+HdpSRrLpp/7TJGTXG8UU/Ez7LaaQlWG8w9bjdY1Ynpe7YxQo8XYjZ
jLG3X7IP4zB9LB3i5Y+d1VhBYt3LxSzJXM004KL9bAdCCsto0+KdP/yBWw4n9XOP
AJL4R0VinZq76EP07bte3m6rtb6zGNwcpIWEispe5aE8MEkpBB9FMlwXns6EEjCd
/f9kXVLd/CxFue/e7qxuFIXV/6Ppnmd+BycMsk28bGi7V2PYyqn/TmKbpV9t7qsl
Ip+XcKNSOAMeees0sNO65z+NFSDZc9lzEtqTBxxClQ4r8WBtefC/5rwjSutY0DXp
UelGEie4Ugm3MxVEQzKeWUbw9R8oTxKLrJ7CO9rGG/c4JCtT5TTjhpmX4G0BbY3r
T8xqOGccOxPUIHLG8k/pQrDNncV+J0G39s1Ey8f8oD2UHeaNsUOiFZAeUe2Lbw+L
RXGF8xe/xvq8F149PhwYBcK41gfpz2y0Qpy85QvqRGWko2pdaDPpsZh69uf8IF6n
ufrupsa47t5JiOIkjKb9y2ipX+0F8/YTXV9YvFdcXJ7EkNpf90yBqiqkr8b6aOOY
gidp+yi8wO5ll2lM62QU1+O0LJwgFSuIt995Y7Zd2GA2zpolREqGqvP6E6NFWMzD
yhQNGgbJuYbH2slPyENjN9npNOv1uv4rIZfeRelIWv/Hd/tNFB0gpg5OjfpAYOQ4
eMmdBQghxs+uOvtbg6Y2YToOLU0QiOYkcPxIMeM9IsBBovC4FqB8nh1mg+GHw0Me
EP9e9aOEUA5RzXZ9clv8UAs0BeuRXKiI3bX7grOY3WJcpakgAaoDeOzXHHLruuOy
R/7QLtrP3vYdcoXilbgOJhaW/q9mBTFsYP+0Gj7kFZ5WJIFiS/fnBmf1yLzQyQaa
VN1h1XZhHa/pRqMomGjx/gnXehiny1uvZ6ZZhDUQVN1jrFcpbjjeELc9fEYVupL6
RRN5AaY2Jnid4eCECuAmrbgEsPTxIOVFZZzqz6AfxHpPL12u75GfcjuqNuwXQVSb
UUF//OklIXbJbstvSGpogIK2WCEfyQwxd+I68SimTqguuBscVC8EhNl7heE9hN6n
5z1EuoySPeQvTrD9eoxBPmiggCUT7Zx++8UBm0d4I1CluqmlNnuS9FXYZ1hl0R4A
+oPTRATL9wfcLibloxaGJMP/m2Nug3EElSzLMv/Pr0XTQS0wie5aUaGIpMrZUYZO
Fd7cyT3nEidpZzmNb/08924RpMjCcjKi+pSxVjVhvOedUWUYKXWGyng10PZUyBy/
DBSHQq+FgexbtZXJhU1RvBcc5Bei/xO7SUtCQIiBafwQK8yKqCLiqFsyS15XoibJ
daDwoWkrj2zpHhnpyPaPYpKUZtd+CzKcsTLtSC3JxyUNxF8fA6XOnMU7dnwUhMif
zZmSXx1XGFsE9arreGmrjv9z1JfVUxgXsr8HGyoXI4278eWK+txw9WGyIe0HiON6
jMCfx960b3CYS7kzZngD1xuTiiCT1ncD01pajlAvoFKMBXAqRE2WOhvHvYokiIrG
VPxWCkJhbpP57Xpxy0j/by5nyrFdp62q9ACAUgb4E4phckPSJzXXZKdrbGXMyZVH
gM9U5mTdS+d33S2GWsSUQ9wuPuCdudssiwkgfSI9trNokA2tzZNRPduL81jk0IlF
iDRdAbiwXsPz1P/pHLQO5doclDrmjHx7uLCOQ06cTH8nzC0L7YR9FelpFBAbZvpn
rE8LLr1IUKFubJ30EWLVfud1ueTcqcPswzNmyPb6flwfAzKkFKRF0GKHUeOIeefW
sdrBAEtAPfY4Zwsr6s7EZQO5B1P0IcUKrc+uTFjo9gYMZN+N6f3tech5dJwMMjYl
8HtlxxhcCVaaAv8L9Zd0TWQd+kBKj5AafilwKj9QGxVk76DXyFtpA38fanR1McgS
DMRju9DM7V21neK6nNqQP6ZduMOlcRRzsztKdldm8pPeqKxTNCeP1KofLenvkxU/
if6Ru0K5y3VxkSy2Ef18FXJSFinP5xAgp3FYLgxW2Dh7WMVjeso9y/Qa5TDxBFYK
P7gxGf2dnkdXxvXoViXBYOhDgO44lei42jutBHxMC7sBmB2LsXzOdbisdHL6Idq0
hUyERbcN2xy9CjXeBp9jA6MeRdJNrn2X3k813ts5+kDGrdrfMGsbzetM79yqN427
V1X/MrOhGIKjEgsZffdrVuBcNIGRI5QdtniQkFkHSzyib/6nAecx77z5AmbWqIO/
xX7HNqvzucV+1vjtkql63N3mJo2dIP2Q8WDhqFwD4rWlhx7Y/2KMgMxDtI0TOQIC
fyAM5qvoqzoGtiZ+WZ9lou1J4PD7rbJ5TrplY2ydy4zGYu02yYlC6At6xUDD86Hz
bdX96pPpctdEXKuEF2R2vAQWHRiDQvwh+p+bVBRy2XXsNZWexVmACJHDT3ByegaG
oLc6UuBEr1p+DoaG3713yS7PsmLS1R7f2M2VEkDYBpp/19xUGQUgc41Dn5HfjfZ6
Bai25+rdoWTGL0iWPFA+g7g0T47ROp+nAAKXVOVlgTgN+9jVANMNuROGLoW1/9+Q
c+OAChF0GovI5SzQvOo/pAIoKMioY1rxjjUmDaska0TmUckBTm4dZ811ty3EwFcB
AYLdmr22MzOubKPr4rOFKozI3ww1QbE20Cmwy2OwdF9teuFySdnTgbDuhYRi5fIF
skn0FK01wXCixv44F0GZBqbaREZ1VeRl5s5s/E7JwXPW118CPbbc2H+rgCHSOf1e
waD0rICP4vLywLVkc0UibUGg8xfDZ3Jk1dCamZ26ovkhjAWgcUMjRFVLLdDIYL3w
1YZhps+EwfuAhudsBx6qUsHuQsYkYj+B6jU5PQNdiQHe+Ki9hKKNCtWTYc5H3h3a
ApynD1fw8rR1+UV1Py9eTRuElLWxzzqAI+4wl8vFBmfZkmt+5Z3Jkl9dSXt8Vzxe
OPgTL0mb4uSf7KUzxNDjWF1fISR9gW/PRXEXKdW3/cIv8k7Nv9PIoTtjxZXEdb2U
ocqPwx+/RdFj3M0iJf/WvYCKkbGmFM1JbRcKCO1SGDrxqougYHIdJljH5f7yEoi7
LYWKQfaz64YXJkPXd+AgLfU9TNZ4ZnnciaN8fCak2vwGt/c8fh8hzRVwg+g76O7j
rPj8TOfISHi+HOqBFOgH5BLqWQm4Ay2pfWjOtMe4AtTee4dyNsMgLERf6Tov4YQJ
ic1Pvh7bWiI4G6PLGPSesBueqQovSV0XeWrW9Me1tVijyncNbx5ZXNeZsIpLNX0A
cRxN6cnLgEvyJJc2+ltthqN3Pyh9uMOhbRGHJZcr/ywkUl1670lzdvsGWSA0eQhf
7i8/rr01VOTJw2Aw8WBByifvETGWNCHf3/n21Q03LxsDrKyYarbNe/wEkBgV34/w
UmMde/I2rfDx38dPv3n5Ux6zcZzD/LbNrGXjM0P6cvtaHf3IOtcVBeHbEiIs9804
qVecZODqBnpgaTW1uhf8WxcLd9fsfr5v1W1oH45QLrYcQ7DAuby52+6IEipmi7EG
N59LKJ07EkjBJ6zf/yu/BmBYHElIfvKCbveb94w5k+Yp4OOdhqw04TkQD+4V9skg
jHM8OXRkIx4q65G9d+DeKk3Ar1hErxZy5Sc7ujHuna11PO+efGqY4Mawc/+zIGk5
zrcscaZ3AEHtotaspyoGOVAEHgbwuF6+utKThUJWpJ6cMP1OAt5UTi427aFLxCkD
GtHtEn0QDsNlBF3vMBHUecc42pHUnlMxoFLBboo290dV7F2UfWQH9VrMZlpPw2gs
sZ5xX86xyHptWjcX2a9Lh+lrO3/BS8QxsaScXLGe5Um8NDmDzYX6AXAeBXYNPUlD
spvWBnkp6YtAmj8bBG1ERbZRhrTB1G2FYkAnllWQ9n/4+BaIu3RJG57mgJznM9H2
0lHOMKdSb/neh3Ou7gkqNLxnS0VZAvreBws/+JHsjzP8XxEpYhLmuPLNsbpAWKM9
vRSG/PRyBttSbxw03qFYb/SauaUNfmR11FPTEwofLcAW756/UZ3w+9bnSo5JBqEP
jiUcdSn5fbK5OKAIzD2Kw1kdhC3I4FPJrPlCH4BxmR3QgY181f+c9D2INOQAN4xl
TR8wt2HN5XZ0cKzt33s7rk/K9TDlUnE/nZbd0NCL24O8+RUOFPJSlSXo/aAfCt9v
0XFo7ilIBoZ3zy8w443t9PnNxWxVYbd4zxTwTzm+z/0oYwUD+sq2vjwZdyfRdY7g
5fa2KWwbo7bX5ub/CynJQqoWiR02dH/nKLe0BXq5j1ZMcoEvBJwc+R//ADahoxx/
IGk/V8pT8w6Of4SyGid+cW5081nNI/IP1ZpKMSAT1tKlFhpVY8Snrvz4OPPCdgkN
RsbzlqHmcBXZ8dfyN5xIFDPyJJO64c5WUpl2+Eez5ZaS85v8Tiimi+ctcXbccC3G
2/Y7zUN5Sq7imKXJ/BalfN2Bai6K0RHHhqOiN40G0ysc3V5ePsKg8+8+KSXJIzIn
+3TEefvNaIDTCsvN97yh+xb2HVdcqmMqlTVmcPVraxA+Gvqlv0biD+H6bmg1VCta
2QeqIrCP2rWluGh+TObrsP4Vs62xftscl/hXmn3EMRGHNpo3VLIjeCK891Lr5+kY
1PLHgoUnKe47zU3nBXweGjWkRwXHAopYgOwroNzfz9y3/QSBndPzpwEyYbe0roaK
5lI0+dJ24PXGAmu9Arf5LrMNbmtnyqHBT31tOiIu0nze4T+rwtDgPwGbTpl052yV
UXpzsLj94jIhKTQ4kl58g5TZV/ygc7P4iCo6WknRZ4QboRDAtFwz+ZtAc7LHMV14
2P2l/EsOtpStum9KKlb8DEGKwX4tqHU71mxjLskem+kFxhWUASdUhKfhFYq3VqJO
CCPuKEkJpgmK8M5MGyyL/LwvLrx6HNEBbmmHKf8JtATXiV5GfDDtQKMVbrBZFV3p
MqQP26leL/h+vwwl0dEQen/0uOjPR2UvsNpr9ZRoz7NTYYQb+F8Ub34oOaKZ8fVs
AJNrR367zl4SjVcidG8ZGAF2Qkj89s0BQLo+pUW7vVrOqiZk2iFdS4z/OnFwJkxT
fvKYIaoOsLihDUagsG210tGD4MK2fHfQUgJJSedSy7v+5kJZXJ/jkB8DjbydygoL
7Mq8Ct+RfCkM3rpkJGoFmMQTEoKX+emfxTbaggDHpkkeiD7RoglHO7pjGBW0zC78
69r46pkO0cqKnLvMOaJEWMgQ3fmdIv/LsMZ/ZAquY5XSMCj9uJXR8A4PmQSIrlhp
ICb+C7MwU7rlcjj9g3XqfbZ0yDD5p+rjfTiOlijZhAxabV2sZmnyZixM+1oxw+lY
74KL2aQjUWJ4Icwmi5xh5/4gDQG/RSHz+2JIQRhzYu7EnKxTaU3E0y0bvWmHMpjp
gf8KyIK1uDhCB1vuIxoc5y9kyUTWBXgNn80LnjGmAIHOiYqwFBitqHhnJR0SzvK7
VkxAPWeYu7WfQQtJEnTUdJjOW72xOxfE9mF2vXbkx0HzbcjCEnB/CLfqA9qDLeIU
+RbVMefmgG+Vcb0McRFTMMvzwtGnO4fAypPIJKUfBWAcS55PJz8eFKwYwiUvlIoI
9YS/kwXmjdcb79OPM7d59PzXSGKATQxWSfOP3YKOPSwd13d2kQojPPPBc4QGj8BD
rbyplyfJu0DBcamar3kVg9AKBBbrSWDT2P0FjX0KM747e5of/0OFfHJDhiyKimRb
ErAYQ9vQKGkxCqqQ3BTvuGWc3A5ceznzUObFYVB3sG0Z0885D20wLkSfVhR9IJT6
oFp3WoKVXHxNl7jwy36N3qDYi853JIKnL4QeZYc2HKE3Oenf/O+J3u4g96Y/o36+
uMs5uheNLOCLooQHc3pS71MD3M4a90kxE5yc8PyiIrhlbk5iUll+gSe/jgMgaq4D
cIlfBtcqiQfOwt+BJzkkisUD7Yo2enmBtDQ6adSezEeMbABWvlAGqAsJwZn/4C7q
vaWK3TnYFsNAXqxytK/ln71bx888zEBCxyWA3DI78v/RquF2rF9mEWFnGGJZnT5r
rR83aLYYug0sJPmOzf7lZV3inmzI+ftRwdg1uyGe4oRKW2yZxF5/N0uemi6PlQp5
Cx3JuuJVfe7gwf8pZ3GJIHydoDJPbEgTsQ32VBPQ4dh9/6X+BWSik0jqnv8Qztgf
5hdbPhKKgXeKllZCwdldc/QOruhKUd9KiiSDcAHlkSO4ejPuCnSdUnxviGc1yzMR
fp+DzCB0usU6sQyAKzWOiddFL+QrGQ7nOZd2M6atJp0OyHazL9MRTAWvzvku9Xh8
JXCMTfgW9J9bzaDmcOD8kiTbYcC2SClBzCwi+FzaM8AO+s2pAMvbgOgP0TMUvWE2
RnCxuWgDaBaKciWYDbabVM/6nexJVSO8+Tl4kUofrT3Pe5rwua6czVKMoPeMGupA
Gwx60Qbfp9402teDYnjQyR1jX8gh4radcVvwXvED1kPrtYU5WQmaTNwwg+D+fqWs
64uVIcd55PilSI5z9MuR8RPs5reIlIS/qUPFd5ED1r02rzBEAVHBQjm3aCd2vcP6
2sr90GYmcvJaF9HVSLobQlGRHA8/blGvaPll/8ZljGfPwXv92iLXsdXGSBCEPZyx
2x7pYz7qJH6+PsXVV7U3+Qyc79lUHo8pt9YGspYoA5qi8aQ8tfAxzn0uJKyZbabx
RrxZIHz2nPyOpczVfzWZGrDw8bRLhz8UxHi/YHStYsBSzjd3yHsoy2QX8tQM8oJx
/qq6xuaXErksvDjYb6g33B6Co8xd9y3Q6POHEQkDZ2orIysJbFdh/IxG7HNTg3uz
1hdYgLIAKCfmceSeKVbWwiyX/84MIER8/sLw1UmWoqTlMJeLc4UTUCA3Q4/Z4agC
Wa2J9c9zr15gimYY2cF4eRhbPymQ+Y/Pt4fp2qyCsShezo21JFDq8hlkvHAc3DNi
s8mpHQ0cil4+rcUOuQVo3s1tfeh9MiFzzIByHnGNi6VkbJFy7mQa4Uvu63OsXxUn
FknkUVgxR1quxd52L+3cv8NYX+DIr30N4N/M/cdRxnTZZKDFOs1WLHkzN3sIAtcY
djrAkVOo7fWIPFRbjsWr8IEXYy4JzLvRs3/cipogw0GxpZZxh4eHLJzh3UXc5kB4
3YF0VFJX7om/py74WatCYelhI6uRawHDQaoRwQmYMzqwAOn8ZMxVFHDciMe7I2Yk
IdWtf3TRsanqfgxUkCscKMsqBXF42E5GpfYIHZBJCUVYHB1pVbomGsAK+6iEfhFB
n/rhYzJXw/70TNRq7WWeHxx9O6pZUM8wGqBvdy4sQRb/oeqXNSzjyvqcMYVeMBpe
olT+DW/Ruc/e1Bff8BsKlaTv2Xsrs9y8lMg8lliTi+enbz9NxAniDrYSRrZuj6Bi
EWrCpoRAP2+97GYPQ75CHKIfN1tOCCeQfwpPEKZVgsZOA7zGNV2INtRMNRKXktLW
WAQJDvf0D1VcCuIIYKXggRiaS2wEE7p9FKqrYA3sPZGIm0HXwaV7m052ADKQkiTP
8DNWkCVhybO0nRio8baTFtMLs9iOKhWPz9vEr6Ui/UBrOuOnSMz+x9G1ngwQ+yZf
Sn1E0gMt7l8QRJPwwNZL3upJeTMvjyE/nHGEHyKn6FHeU5eVBeYPCowr+amJiQXY
mOk4A+TrwJUgsZZp/12XLYnRA/eQ3/tLtO1ei1gIEf7Gp8G/f8QF2HOqmamaurc5
RaCrWEfpQ7XkP58+moakIB1fU0LiWXXl6ejfva7jMYVBJ8PqRHLlr9Ejc34xMLLF
AtsYvGWhxv6muDcqtf3A0vlRKFZQMutXUo5HZ9JnR8hoKJuONGDycLYEevt6SfQZ
eYFjvvcRSPDrMNp3TBkwvA40joa7RAP4hrlQy+QKSM4zN9qy2Ffv/28gLT6AxOFX
zZOSKm9eZ49wD+1AuAb/ud2WK+BwyYTInI+8SCoMffK9aBXk13x0jkjbqEgk7PQu
KHSiVTJs3VPcd1cSPya9unSR8eJ8jTvpzXU/bduTcp8kLBVBccZxcVUXE7etTgzr
mrEG+02oN/ozsnxviHdJiL83MKz4Ps5qiTEd55xm5NCcRoWKvL153xXDi48nnijt
CzFnzPUP02Al9fTMlvAmVSSRwIVCH2c/NqdOpzl4Ff42mZHOGl1ESo69n//pWxbz
sf/1oF4I+iM5SRbpEY6v6kJH/fyz0RqAUARI9V9vxqB2PXIvszBi0a3yVk+kYkPf
Ns9xl8nphVfhB1invWQBAD46ybiqueXcxyqkfsi7+unIhWyOlXWk/8q8gpBDlr2r
dQ/XEtkRmU++uQS35xO6sitqUUyO8eC/sfwDNKUJRSi974hCqtNL6IFYCUiHiKEJ
uzlBwXTGVYeyCLkd1vNv9HN+bllVw7Nh2zecNCvb5fW54z17FEOUpC5rm1klY50O
8a7ZJ1ZU7OWyRFiCGDmPX5fOkrC7EZFDjigUNEi4BuNz1kcVCM6+3Tz0i2pokNfG
TsmO9r3xaALuFrTR9P8o5+U74CDw+eOkPBsZxVzLvlCt3T6RoxNYiOsX62x/GvFI
XQXhF4gNj3tTW2pMwTa3XOHWmYEyrAMDKnU4l5RubJdbAcE2lKlQPU0uiZn5owFO
5Xoxc/LAjKKsRHfpW0JCIdEuhZLH+RVvtFh0iZJMeH45PpmuMQ8m8nJdfTlsSbGy
QXzk/D1mBY4Lc8cltMz5clq6sNWlzrHA9opzINvHaIouBEH3m2NPboA1/UamGBsf
TgeF+rEbnJKXM4G9bRJRGURFpxstyA4M9C3tg64sdBViCah49GAcTaXI4VP57DT7
aD7pffeNFbcctWS7lntBZ8fT6EbHREaSKh2D3S0mYjuFFFkFq0N2qRoNpMoq+VT3
itcd+pE1k7fsFOGHA7vyxeT8GGB04hTTaDDWzqP6B18qwhZ78Tke+/32VGjQMgW9
5+b4eh+agkZ6a2lWmLewiQe4gBGL54KRIxeBhFz/YtakbC8pzjGDc0dL6pI9qVUw
ZdbSWbybmy4RNqYU/ehs2eQRQhHMv2O9gJ/8KVT7A0yjtFFCV/gdJHN10Oz0Nb31
2K7Vb6BlG5K1yxzGqGBci7FLFWdAySYM7Y4HSZ+6kx/iuPzpKeVrey3kgFxS1Vsv
KP5Obsayc5dFCodrju+FVhO45LfcJTheNOoSNb7bXOI49Wo7QQ8Pjy6TimjRh6ai
Hm9WuhEpJ4+NUzHToB3iTXNvzcK/hsxm+WGFwUOuO3EYwmjbNEJy3pwZzl9VPdKI
kvGisaoR7i0XWU+/wpRIz+LBdMQIVe96UMZA0SgPZeNbD0aCgV0HrtnwuOxwZtfj
ymmIMZx54DgsSacDCO8gpo+FJHzckv7tQLm+OSsnw8A6RBWy+QkbIGikKqsW3cWV
stskzyOIN2osAwBhvv0/+vJ/g+OzBbLonl9B8E5oW8ChNzGLx3Rq7KyCNtPxwI1B
L5b3nBdXZlOcaZQp+mfde11pB2g7l/0h/J7BW0GeohEWCKUJtI6k98QrTww0KecP
Z+3GUHVxacIhw9sseDMQ9eVGn/v3YM5dLk/vNERqTVQmM55mZJ1/KJn3zyjHyK5v
nGRXFqgiD3tUDKsSeAMzKmBBurZ0+nvxamZwYuFfqhNxv8lvJc1kj+T+3tjiYLWt
HCvQgrDuV1hWly3o2QJmFnk3mBysi50yleuoaX8SvSSQcG88jd2XJ6Z/lgQqFH9C
NS3t8aWEvxgr3uyD6gqQYNLf6sCC6y9Q/aZYJnubUMh/zta5mCe2fHZpGk8yjHDn
Eihup5OzsMiFoB5/WPfLVvz7ekei6F5VWIoIM5Mz9IiO7uBH3hgakd6N9A8W2RIf
sRasHk55if0vng5iRNlxDZ6kBMvEyW+V3hs5H8v7GRjHHyqp9Dzpg7fEfN5u8xbC
Sb5zuE1+hPK40EP/nNUoMxOQm8tmWIPRAVaSYm3AQqBQh0/1te7vA5pIvNfsnJAd
q8JgnIpvhQ7isneuynVzZYH5qTswDrksdaBOLZjpgybO1CYiyc3qaBK0ZsPal06r
Td8Axxny5jZAX0O5zAM7ejJ0rYA/n2v4WgbKug+/htVWvlDek/YvQ/lJvX9p5Km3
1Pd6t7PK8QNvDCfcDTpilx+cMvJuG58rFpkjjiUe7MSGUF3eEGsXYoU8NVWDwv0R
9uJ3oy6h6HX8DNu26S841Qy+FLTYYKzrLvQ90CXybEGWPOiji3r3WLXuSFh6dCsJ
2OpRjlDQddHGeC/rxu+OTleiL4nmQOTcDJ32hlcwaMz7iE7eDI1jkXiKy1Fl+Q22
IsDneCWIEx4vStJF/y8InB5/i5Z/RQB4EE5ipXv6KNcDd8s6Zk4oF4W+p85Ctp2j
7IAAoQaGRCV/UL/Wm5udp6mL1iEVwOiyu/kyHPy5tbXZkK5hZJYoTjpTIA5YRzlZ
icNOsM3gFyzY/8CppN9dqcA2rvpxFSVi0GUiEQ5RReU+Ot+k3QUEQacRS3+T+8L4
vZ+Cq7XmIeSHvIulVSVElB1pbyenWy0s3WztvXwknmPnysvedEGYHBdnCDWs/PTA
V31BlhrHarLyytkQFL1VI+3LVmhSawQ2qhgwpIxFDd6ix1b+s/mo5p7LP6l5HENW
WkwA/ujO66i9a7zswjqoZMIXCYTEJT3WHxQHAvrVQd7keHkzIoZf7t8h21kGadto
hrH+SFoHMl2ZBJHGnhprTa0nWcVa/7+rx5OK7+ZHZzI2aOXZ5/uAtBdsipEb+lbY
pW6lgh2cbYK56Y1215NqnpXaIL92+D0sAvNjtYT6/ZcF59V/r7XTaqDFRns3rzOQ
tNtUrKSHUZtyUaItyxTrddK+BM+a4L+OKhsd8vhysIOnDvFkkCzkeQsjzp2zhq6J
gP628LsDT3MslRFYmlpPuAoS9/8IlzAK9kHcCYeFL9vQIpXpI4oAHu6KOS3kkKBC
u7G+A6DKmGQrM7wK8L40T1HtA0oKyfZMjeMQhbsw7bHXpuCFDugvFeHigubHPcdM
1x3KEgc9hYhK/yH0JbgufCXqT5HXdC6m+hUZg6thi0fFenjOQtv+fvg1HdwhLtFo
5LfVTVqami8/FLIANV01SVyVDJxCRs3EAG+lVAw1q/O55fBXUcYSQNb5ydszog6r
NfR5s2BvmvRuxXKnuvmfTE+4XF4TWU+n6PuycvFPqtK4gfR9mie15prIKau+7i3U
d7NUsACleMw5WWk7DPa8IPQRG6amEGv04DH04T8YTxvrWRGBshfFBBMDyiPq4goX
OggiNHXK3fU2roAa7zTL81knkcauR0EnmerR5O66Epz8rwNuXXGhjt2L+yJ2gIbj
UIZsU4SvhmF2eoag33p8GaVnjANYmrMiLg41UKjd8G8tfhX6cfoAIjvh6CmS3/nd
Zky5YSUtA8xvzjupE1eHpwHfdfDNFxyYt/kPQdU7lTRQppvVhm+JgAHkXQgHQPnA
mJIVx5/BgJLoRnHeKYA/KStx8n3bLbC7KETo6ZFOqk0woAi9YPr+n6mZr9+iCkog
+NK1VWPxsKSuXnu/ysgyjxVGRyHuX1dWWYp99YD4lHlsKAF5fwQ2Pd/1PRBoWxcz
bterTybQ7orRhHPZQVEsVyQlUgDf3te7AkJxEuSBJVXKi+0rMjSISkQbFnfhqfjc
2MK1aVPi0fs6CysFlsRFnNWK5eokiL0cWwG9it062AYGveQ9ISKjW0kIaKM7ADRB
6ZkudgxBpRIsOH5kddGffSsSbUMIKh0D5qpx8Yy6gsPq10CM+LS4BM3La4osw2gv
XiaAUGEmR4N9tR17ZhcvsKZJ1KVq3AOJODVfAHwmSUGHhh0k69Vk4kLa3aTIDpOR
EpfqOo2bYMHhN/+vmJ1nfXOymFZdPBEAvMJjOA78k9gSxNj9NEZ8Wm7nSyFSYoJF
PdmjCX8IkpQTL26394y7qJy8N93hSbdS7qutqScao1THQ1wIwgcuFsKQd8r6Nx+8
AdpQ4FmCIKkU5qV6nATslbXEdRnY8g44o1Rhb/Qr8RnMMR8Rw2qczH8gFzkFtK0M
/M9EO4EuQscoB12rHuxRdn6R6AsrlmTTxMws6DWCSRuVgoyqEAvdY+2KeJTuWfvR
l1XnCN6UA1vv5rg1mCWzId2VLQEPhZjNxNqw9Xpu4YlbBWeETXhJoMJJ/Nv+Ox6t
yQ18jRw0Il71WcadCRRT3LRqIYEbcB3oJGAfj1P9V36xreJTmA/8b4H+X0LeXU2K
vFci9UqQE1wOJgvI24Bk6As1gyPwwtAvwd1nE26vN7fdU917eJCrwjMJ4c8zdq9Y
ZwApKIc0q3g0QvrPFlnUUWTJBUJrhsYTleiPP399X0JIv3M/IGjDBji2Paz5xjOP
KuNfNHK/tiynIyInDvvPJlljJftQHLBjIcQ1+k//vnV5ML3raJ5OYN8K3AK4Nh4Q
U1aOnKy+aAJH7o7I02pKpUyHwwBxHWzZ9z3Kop/B3C92rhcKW4B53nMF+UiIdbeC
sKgk13oie7VyvJOcbcZJXQVJHfrnyxIztqDG6BHEQGeJtVI23/S89vrTqLOCAht1
wPkl5mxPaFZifJwvp4RsWzLUhZFXmDu3YiausarqyvnXoPn8RRHmae9e3yeY3LVJ
k9cJ79ItzxXdKhB+/uIaYbEsbEbRQ1Rlv40eSYivga6PSR5k+XdVlmbS0b9H11q5
yORcdf0H3+XBtBCXgxMgjVpdYwrbfcy85DWD3XCIPhXKQy589mRaw8RDS1U6dQS1
GzFfDFK9dbDqT47VLTY6TkiIOuqUg1fAYB3hApx1V5Z6wNX+qCsc38yFoBkdEoxB
0I/kr0D7Wnfmm1YKVl4uYn336OHOyP5Hg4Nrjfdcg3Iq6DIxpgZc2++wOsGZC/4s
+fDpZT71K0R4ESMOBJi69a4RlXC5+7keK0p4bg7jj1jtnJmcZ59e1iuR9nCg6R9N
s637Y1teTbaFpHNwQLTahBYkOtT+rFPhmntEzG1UbPSiYgzFMiQk2lYi/7dS2GV4
1PEgcTGQgmGV/v4jp0RWbvMtSpRGHI4/dr5s0hCaqQ+IQ9FyJ23lU6XUuUoGFvy/
D8MBSMpKaCiIapJNE/xPINoxzZNXCWxbCnWDNZZRflot5L50/cw3UOm9hVJvGNfw
IrpC/+I7f6V71svcxNrqqgm2HAjqxrPJOzCYUzLzzs2AX1pD2qQkOB+q5/OsnBUQ
e3drYzG71tkLFTtK99MA+DCnzSiDDbJKZ4bvwYh4lYR7fGyOIrf86gQjFIPLwDXk
gMVnFyMfJzMnEqjMeDJ0xCx2rs3TKkOwBCnnmK3ErNJ68usnB+hawnxrM2++1PBC
L0804vRLi+11TLLfiOBJvt2m7yjX9X6j0V4fczsvFpWxv2sEJdfynUWURFrqMKll
GNu1Bo7U68U00PPCxXDz+aY/nlx7MkUliG16Rc2AUji4yRLHjt7J7ZltQXD8TNqY
0iKhXAIF3Sx0zmV2YW6J3EOUv0H/f6QfadBSlI8Yg0RiUVpukQ4VThuUeQlMsQdU
FkKO0w2ImbU4nMoHrexFBy1GqzxBzCmvrI7ubkY3cxRazRJEShe3TF4hai61rRup
mVASLC8Y3z3TJzllYXq6HlDN8wgIelMf8PjQm9CXbL5GQGw9G4k52kb2QD4WlH9S
B5NRod9thS5Hfg1PxFw/cWkOBYs+li9kaz6KvOIuoGH3S/ujMiStxca7/lz6xaOk
Z2AaP8Ui1DOvdmgtP7OSPsaaNfBZgC4AZA2U8dK1boLHJgcb/7LRzadUWfGXv0Ut
iuWoQkhFGnkkGnEP1eLBPumXxCUxkchMmKDmwUoqV4yB067B4k9f8nI/fIpBA9L7
NHIiwLhkod0o4rZ7sAaNIiYNdGEGcKqRWJ0d2/d+2DKs2r/s+dZcQNrBnvUZaYQt
YZXvK9DopDN+RYsjJoMq7HK5hUeAEnqys/KXfBzXsPwpEazpEuzmRQ+CF/i2RqzN
4Neg3qrz8vNqC5W2GQJGGrimpI/GxmPepxfxzNB5z4F+C6RxGlRIULKRDgjWDv/z
GxNSOmeddLWlCKbF1RnGibLns+1pUbHn3eAtReWWowXbZ5TQX4ds8DFzedZ7ifn6
8Ssg5FmB7T0eqWqgtCCy7n+dAXNCWH4Es5EGUpuHKlgU+UzwPJNytt7NvQszbgm/
Uum8KAuBx3JNwTzMphBE8QnEXgJfLFwWxKjNKwAV1Sbq5u72NBNekBihJJMe2bwl
jQBrca2ArFVIx9wgvovKyK+G87G2phrfo/Q/Bkdrvrlm5XtIFNeC1LqA2O4F/Lqg
PC0cxF9EL3aE7Le/tn9QXBJ5Z17idUlAoA3fDjP2zhzsxe0CoX5HVbm6DCoDQBBe
Tsit2xdRFE65jSSJDo7DfbYbdaozQULF9qABKraQFKM3tbBd/1lplthG6B89Plv0
4wAUQbn2JLJUffPS2l9KGaBv/NIUJpPS1SfowuAXnpXV9UdzcDXN+4r4jM+TRMZx
G42M4sxbQvhFre8r+914e7CG63f+3HsaawAb3NR9oDN02uc7fY6Q6nlYsA4XMy1q
7FkRKczDMkrSzT3ewopZ8nwOOuXl5AkCJPlnvq6y+vB+d+DZZMPzt+fY6lhLZF0h
zqbJqzKzZy+Zf5lno03KVr4lN/rS3/28JKiWYOW5WTnA8K0hg2TdY4g44n0Lxdki
YC4QgW4285j2oAbe3PFeayhQjegU0kdwIXTV7pcomwCW1/pRWB39t4gf676Bt1zM
hSXqmxI7hIApSz3uuFUZAF3cmvDweuJASor9nl/eOTiHIQsrxx/TieyoXLXpHFHw
1yPEmiDb8YBF3bHEVAU1pLwrQyCcI0HmowMVnmjInM5WesHlqbcTE2GKOB8vupPq
oFDcByLGCpTN2142XmqrsfQ0fjR/Sdv10AthY8zL+ZdcFoO1E1kV7piWLoOuz6U3
ozpTWu+N/0mukIa+xSHs/nQQACG1otpSMQL8BYKWdlj20kBNG/zCCvV4CrIxtL4n
Ky+jZhl/oSfXpEjVq1AYHhfFY0pFJgHxfGsKk1f5KkzQ0J/Lm4EygxcUtgaRIulE
neFD84uKZKGcIZsbOTpgbYU78TWz3W2JSPBrq4JoeNGjDFksx2aMtxXcoYVTRRbD
C8uEe2VyYd+MeDb9jacP/eJ+WMXijLOkDysG2D770EQnZMKtJp1A2WEAt2I0sNOf
LAux2PRiMYJKUpvFn0wQlFJGa2fj1HCkcJ087esAgPEj/rrqca0izrPqauVnXrlR
bBToLHeDJPGMpvXb+7xZCRqeGrnsznm+MkwB0qCqgcmQaDKLE2tWYb/0KUD0g96J
Yuvcf8NgRrxvINST5Tel3L+db0ne0oOGspAlBxDY7WsPiNu8ZYxEWSSTH7F6+XOx
T1m82THrvCyko5iUlohpenpwk2t4oNkTRko9Uvv7lWHKrmVcKlXUaHMKTK40Xjp0
/t40fuOaGoQ9G7LSc1eaYv3C/YPYBCCjnFrMi1YGYPng0MFRszPEQ2wA2+j97Yr6
9HBbMnxWkQp7+rLi1ngHqbVJhplE710jQUnWw+7l+9QbZ5kFpoCPVkgvSeigKRM5
tDV18SCamoE/ThKiag9mnIUn/ts4sIFv/IoGpzwILOuE36n3e33dMrSV6QpzOStY
YGW3ih8dPNfD36y7s+fh5eiRU00brnXi24+tf7b+WsOnbkpbeJuKuNs2TQNv1vSu
mJCc/3gPc+85+NNTMqkJBxN6PLqJQeMjUb3VHIQ2vIPAomkR2RrkrT2ZClbrWZUr
i0dCFRdFsTRHTkxqERPGFbgGayIXL5Rmrg5QiT+38UDAroi/jWTNLfb1dfFGt+yn
G581g3XSE510fXNaWZpBiRErFkclL4ay661/JSL+PvQxjEbUZVrF8KGlNB8umKMO
yTl8FEZv0TJzq9Pr4VN/cVvUewXBL17Kdppba9bAeyrpkCUc6iAJm17842HiyI51
AQcs3hW3wIZOmmSAY8aq/3+q6e2pTxg1kfCs6m2iTFDt4ooSaj4bQwB9ey4VwXAH
WQTAtDXJQnTLOAsMNSGX6jvBfbOEOL1a7JaCZqvpO5OVjperDfzGYa92yJiFazw0
6QqNYSMGJlif2Z5LqL3O+yO/qVP3jS358g0VbFAq5pIXQoXBWXymOtH1ea/o6ChH
B+4NFEqyqbAHlzvY9AKYf169E6KRTP+yv2gZp1pkC97TEZ3/OgrZ3iiofLHxCI45
KJt7Yk3rMxinY5fMLBvHizfsia4eCsNTmsqAbpzSuehC+fzSTgsaRg2za1YYPYim
Do6EDjKwnCyD4ZK1Jet8Jkjf3Borq9Ggwz11YHJWEtM0qo2m7A0TvWA2GZuhdEKA
F5Y3MFFSobfgDqwYkJD9AUr2VHecy5d0nR3omdnzGxzBQ07XFWBQTKZPy0GrS3Lp
zv7++sp/m4N7Uxrhklp65uspKc1sx889SE7HJi/oLJCftO4y9MfVtyofDAlNJ1Hx
XneDB0HCA2EBpy8ELjnX09GIG9kzkeiOPG8dk59Kkp1kiqWpyjKaG4chTr8nnN7g
CewKoZ2w3Kr4USDH4r1eSPXNWYLrbRvuD848sl0+u5yvPqxzqTj62plr4M/CzETf
eMXW8+VyqWky/RuOGubK3fJ2hSDuJyTrYU/wJ4fNz50xSz4K3P2ps/GJOMiRbgzv
TniU7s3YouxTA58kviWQZ2tz19eWyeumQRXbno6QfK3cuqGEkWB71T3WQrvaT3Mz
rBSGg3o7RJ0mtfPAtKX1Drb0J5LyJhxS1exuJpKhEWO9VDhSo3ccJz4rL5j8kUhW
q3cUtg4nEe+Cj0dgOOS7QZfLELziEj3k1IfiPGQ2wwi+sVVYLwlE/FmpA0VqgbEj
ar++pP/T1yIlv66afaRrvONL9UPA9sT+ycEoidZn7MuC+Nk4fkUDYvLbpqSofU5X
kD22cWLPhewr+R29eCB8eJ9fuqx6DtC6px0bfddzoBcT/LMBpXohMjfpkeVHRS50
LP5895CQoKerpe3sHNguKur3kjvowmY1uMz69bYJa9jeGk+LgsWgxB482uFrsqmT
aoaKtAYth0iG9ECh8MVS761ZgUf9ipZ2AHUkts3k7zy9IYEv4NYwXPR4MD4oiLgC
4S4qpaa2KgjAk6vbj/+67X75Vspljp7gbby7OQw13w31fg+Llf+Uftiwf0FTbwy3
L/JB2o3c2iLB65J0gMFFvfON2jAqVotyKhyKA+WdRQ3dVTdBhGE+3EvkHIlvBZUl
PaxBKdtfZXFKL01rNdmrWbOeH+lDeO2ZvvNBquU8FRgr1+jA6NGYo5S9jM378/l/
ZQrR0LlcxMDWBwMgM1WjgovOTBDszYpDyLgKNyfoLuIaDepk+7tY6geHZKr37SYv
x67r4z+m7NdaqMcaTn8Rr2yuSD4GOxphfdVFYaWr9k7uR1auJVQ0Q1/cJNs1hCx7
HHQJgBLnvc1yK7b7hlaHOlrdAIN63dZUXNCTLa9ZqcDhCeuuZtMZ2VTnggy9tK9l
zyaMdFpimQFhT4MbfbY32c2atl28M1vYwfofSJ1Pj4AIqz087BKkxzmwc2Eq52C6
7WThxXGlfrRvpB5jVAzRt9ZTMIXr1vhXb2NuGSJh/io6GA2hcHsTf+Xl1N8YCuVR
7upnofm8ZGV1Qfjxk8UqPlwqSNoqC0EzW6lDhHAYZ2DZwTIPkT42PNDXGx70Ssmb
t5ITI1giCk6zjhMkcvYoph067go1GYXOqrRPGRGFNNJyNY0sWHieJIRZv5/Wc9C8
DTtoPyb5yriVibbxxpeuEB72sHXlZ5R9H5JJzFlZ73ymvEsk1ZGUXxaXw18ER4kO
SYo12m8nnb0MBi/PU4mZYlCryDdBpxE7XpeHLQBwJo22GDiefqbI3CWHvJCG2Ewt
Yxnsj5FYMITNmEq7aSXM+krAvfwUaKrFECiBNVXyz7726oHxLcbEtgVZncfJ9Lzd
m+7cNPkxEhiXsgiAGGLFMiGp4B3b9+bLc9cKdgVD72T9d3uROnRKsDOG2SjkMprd
Bopyoo7SIgWPFLPw0ufnOIbkg2y87h+9aP4sg7ha5mIlP5GFi51Rck1nS/ckeNO5
yzpa9jFNei81vLhvxgmmhjUAlquo8hL4vs5wT+DJOozEYBKJDb2RzjCkpL/BmttC
3jT2qj/xKQTNqnp1JVqQz1s07Hd6d+9OxyhRo9PNpdNdHE70DvQ6FKX9qR2KyQ3A
V2x0ew8MadPay8FoOpEll3DX4qS9uEEg/TWEu1FrofPnnPU5N627oGCkDZdMutEb
UCn5NimASNqIu8zSGO5xnRlLdGC64VpnB1LRJSpG7qDeCDHQbDMj0MDHC/BYsCbz
MjLHGpkj1VfAJGciO5rPtbXV3Lk/Sjwe4EXl5pw7RUupuP+clhap2OJ/1pG7Ra3R
j3nzZMW0aF1vyG76jfUFV5/hG08tA9ZyX/ZBVU43SRYaQ4+AfFQ9hI/XVCf9jW7j
ERI7alUdtNtyup3v62RlDJOWvpl9xlhQfm0Azu5AF2VkyOWMOxpFXAkrLJgSWTYD
67sJUFsTz2eksXrdCaEPX2CYvJ1XfWTbzwbOoFwOfsWgnYrC/Sjees9GURfJdGlc
/+aYdS8jV1P5K0HtqOawG+RAcPp5b9pZNn1IOsJ6/h5EIqgUXuBVyL3saaMYeWV3
GY9xS0gUQvAcXL0ODOOfyftXjrld8G6ePeOBXRtI5F/Yi6+Jv3TFTEPXylDLDYN9
ugDyBqxbfjWfeQ6sQmYjjwFExk+pHPBdwwaaXYBxi7vYGlE1aMgqlx7AQM6v9m8z
NZnELThGfvetOJS9tP9nW3wgIJDHrC4vmccDzCcKBzersGsV3wqOqD881Nfah8PK
B9tizT1YrDTuhXcFN4uBCBDAtVQ1gCV5L2RTSCmm07UfOCTina988ky3qX1UDo41
jdWwVl3Ml5+2Els2/x3/CP7VIz7apqXEse7EgQYGNJqbDcAl3ruMifzOVtC0Syc0
h1wwAtJj+FnyItwgPF47DRq8sfeZqXmx8cfNCmqeA6DGKS4YosPZ4NstJpCZwx4+
yYmwzdn8TCUYoOCMzupnwzZEs382EcAa79WSTMxA8xx7Q11OgcAfcJmoyaRgp1Ba
3A38FalRY4Q6qzl7eHAfqAa+JUndExW6ZJlaoyX4yyhiXCaGtcLT6lHnODc9gTye
xjjLqAjvgYdIMEBpp/SkqCFkb6mXBkPHcZ7Urmn1xnDPU7PTPcXAmUUTteDmu/RC
w/XJpvaHAgIzaaX5r42Neku3VpkvgcAUwiu6h8aAWX2SZVRGaZxrOVguqN1uj3Kl
5kzL/ot/5U5q0eEYo5NmWYxFQJx9S/FQ/tJMTswDbwXl4bIRBJlejPE1SiwUwifX
xSirCqs5etlQoDrfO7q7LnvmUA9DLG4UCVLEMV6Acw5QKWMWqKKetdQFDdvx1AyT
xXH+Z1xGcexJdQ2hjLoLbWV16Mw1uCsnHe7frld5YeNVse7I8AVCoLJvimp0BM/r
Kjnb06UQViHIX4ydwU8ojNXeuEQvO5uisQQtiE6yDoaEntvLb0FFUXv5Dz7XlGuX
rxMoG3wP3UesGZTKIKCJVuPjJctSV0RalgJZ6uksSW9Ca5YfA572Puog6DbD7luz
Ymypc2LDcdS0a/e7ZvvGPc+pl6bbrllqglItQXizFU4sn52Id8WMd6Tx9jd7y6jG
NlAWaUNGMlprhPfQNq8xvBJ5AKguJ89OYXhr79NmZHvAg3DP75LjnKN/Iu8STGt8
9zz5RMBeaampMIAd2raTysiMxbfMt6s3d82QfyJqdhA8a1/kveRU6zeu5hgdQON9
+6ArRflFXM4jiSK0wZTUZlZLK/oypzgE/WXjdS/DDO6fQWp1BnOYU3qIrnNEtwtK
e3lBRTw5UMgrbEviKKwLsqGNu/ymlEkZVvszNAYSmsG20l6l2DXzN19uMT7tZP67
0DUl74Ec/LwK9sHgb+37kjuklglJwNfAWTjCPsUHP/Y+IoQPODsw/+Zlq4mcVPl+
MS58pH1HKyMJqXqxM5BIqxVFF1/FWmdmP9mI9IuNNXcYeLtiiZGt18bdaOEgSRV/
GkdSSZwq+BGNP3O9gS8mmKcqeLZSD3hgLxAPUVNQj7D1SY8zWu1gTD4GbLJzwoj8
VDUguaqjoskkHRSeojjdD64KVWBkgPzLJsHJ39oP48nnr9v7RGw+k0W+hY/JpZg5
wTlW36cZlHR5I8s3JR+CyK04v68TKlz77Fy4Kn9jjBkPxWD10M2IsgceeQOfwv9z
fygNDF3SVgLCwR+S7sGXYhacRLP1rXjoPRy36kXZDUBzuy/vYmMdxIopiYuKaXyU
dVpwGwUk30VN+3D2smdNZDiXUUpk/QWmDwmA2lmm1SdGhS2fyslOAgGrdBPauDzy
u+D7cEJTG9lP+JR/Ebe/O9+7l7p4V4FUWCgCYNuZu9rmL+HI/Q7B/BUzWyiMfpeT
Ae91YkASM1bSadgufSbZBPJUC85OrqVL+MFy7UNfuBnWwNM72paTHA165Kds6wUp
TMGJdifbB/PXgROlL2iTCDXg8MVfHpCOX9sZGahnnJ59hMFHldPBZ2L//VYpJemr
5/pHJJ+UBXQqpsbST648OLK9SxjQBtYvXzk3ZyRLnC0COlO8WcI7tQsMRDf0P7NA
WuPdBy+yuVGaYF7A0FrNF/ldG5zL3Vjx/D4vPOrCNpPpr8rgCqTvO6V8RfOtzA2R
Qdygsoihuiv5UCFbAB1NQt2FK0N2M5yBMxkc7lFhQVfdgqJizcszwhk4Fg7SW9mF
f1ujye6uSf2kBbxKRNII6xhbEKpFFkZBvLamFiNWREHLKGWYbib125DtdjC48PbE
0S/VIBEVm7KtOt5AqmXw+0hVA4ZSqjzPWDdqBOnEg4c/ZHzuIajsUs+MNZa/r2if
wsAw50pzSD1hc9nLAAeYGGPc25yV2iXB/CHm3HToQfY9F9jq26m0GcwUndCvS5xE
++6tPpT/CX0Fu05q+kir0Cp+oFfUdXcxEC0NhBrh3XbR87+8WFblIrrNCOc+oOhT
fkBPYTNZtOLJjA0qM8R31E0BuD21i6gRRi176WsNankVJfuYjTpf/iZzjzDlqyoD
q7vPW7mWil8lXk0Q9QL0E2ji+iiTAFO3jHHLwhNVj1GpR6/pcEZ1y6lbqDA/5Skp
ifje3YTfRWppUkxFoATDMSxqmslaEWc6ALycTQj/eo532i2bglsUkoHnRCrz2mLP
EEAeUWcPnu6kZOHp333NIjjZPtLZgLnbmMLFt3jgODOyBmDDFhbrHUbc4iIB71tx
2k95vjzoY8SahaflXSfHpUJNbjFQMQtrtTcMGpvpd7z8fwvAEeP/CWDBR5P2g654
OefftEOgdgeYhxnBxn4+QASc3NF3W+w/dc+vzJZbYSJRrUbboIA/33KA6XkOKNQf
+A/F1HnRBJwfIYjCAcCZ+hJN2r9EmoBnrgI3gFE0reyQS1h9q7hilVGaUJLGtcnn
GmzUliwMb6gjKSW+NqGjOCeTwk7G1cLFAm0M7lBkR2JscZ5YLpZfQ+S2jn5uGEwh
N8ip2kdAim1HJEck2s4fjjaD/tgjGu1w3Wwu9Gs+ezRXQal2eEKWQMS6jxW5OtWJ
TVFBxbbPTdN57eEEy3GnYsu+Tr5rpIsMG52cv7nFTOPi6Lfad10opCmtKAQluBBZ
o/3PGNjPzG9nAi/zEJsrcjwtzVFjZQc84J3uHw8sI98dfnyT/eYNNlnJxjLjkvRY
J7GUgaLzXothZXuYaZZF40siUvRRd352HK0NA+iSF7OEqRfTJNsLz96GCKHRkGQV
39tt/jTuv00mZinnbQr2VO9XzAyAKDXPLps36XsZb9jpgND52BpSJOy1GH2WKCuR
NpCSziO3QuFz1Lw1COHplx2oXFzy1b6OQywSd/+C7Ns+MGBx+NPBoCecM3+ykd04
dzIaK46EM5cYf97uhII61/qvfqlco7ii+uD4c8pgx+UQO6WSNYyF1ZBHiABsbi4h
fOZECIamCvvwXJ4YeE5De6+8eevOuKMBkE+iv4LwY5/tlg8dTYn/r4xoORaDrDDr
htHbeM1fqBtVK8XIJuEKG3Iby75BfxDwuyPR+/IAGK2pCnNb/ugHAVN4LsreM++c
9q/QjWtLEiCaQCvsZAKOyW3NDfV91dMKX7/k+xkSiEuusXz1iTL7055kmKtfDbnu
7xuZMeq++vwigJHzS8DfsnviCg7xUmQh7D1UM6U8MWMWEvA/KZPGuGrBj9391mbI
mS3nzqpiFUwOB6ObDTumaztjqxkGTi0mPWER51sroJjkv9vd6CeorX8oXsNC7YfN
vXjMXQVOncs0IyiHZx3yO4AJjpXrbNdDJH5Ps9Bom5vajbeF8wy9OUL5AL1c9VYI
V9nWslnQughALR+lDvhje5617yA4JupJPSD8UBe8vIcCzwdtQK6gR4PHiqq04E2o
XTe3TRvpJPMFKpxKjutEJuPnQJaxUhpHAam6zYRGFU9fnSutCrsFe/1+OZvVBxKg
D/4B+FooFxZsb2sA9ngVyIoM0C5ndGh1dTlt6aYRrxuip4jJCd1VyQFgELW0RnEs
zWo7HF+uuHX1INKHo++TABsdiX0X8kORuDXutVFG/VV1jyVy/E50SZk394RQDA3J
h1QqFQARBIArGYM7NQvySvJZTySNfsqReEY7p+fwPYzrllqHukoFFwXkJwEQ7jyK
yu43tJcMnP3piy8pYLv6reEWRPE84F/lppOFDNehm6DTQlTD9pcD7lzB7HE8ikBl
69OyIjpb33QaLd+AcF/9DshhnLjfwSq7mXzb8IjgFNuxbxN+5iuq91P9u+arg6ur
Z1yRO43Izjcf93Mxi1ZaQbltF65drou3imqWmlNmtj24G09m9Axc0XOvg0CFaSEo
BPpcTJzyxv2Ni5ZNH0H5a6PNn+zjWufm3MPBSBH4ao5lo/gPm4jm4fr+qBiNfc1V
e88TOgn9EQcLhcFVYESmoKS0ywXVmMj/qxv+q7K8NLNHCkNf4EEk8rApC7tBMBv+
mGUnuXSlFlDno6ZVpnbvMmH5B2kAY6BOSlnc9nLePmFzoUhqZ7X8eTvrq00IOPSJ
aiED+y5Py0fD4na2cGrNT2CJsHV81SA9qMvQCw8pW2zgey765/HKAj4QNfXnzL9J
6YmSosB3z7y1mCZuanp7yQTUEF+eO16frN9WyPkA9GeKdqStVLrTVJVA/ExVFzT9
oGIQC8j2ZA2pXeeyt2cqWF0QUCZWkAQX6nT417XehPMBf4kVGPWfKd2KCSlTJGUc
qCJw+h5xsYmpjdYyh771fggvn+wLkJlBzs9BSaCkz7S7MmQk7WReW+pvcK1txlNn
fJtClwNtZ0FMdNmGLK3sNzyFVuDUDkRKZ0RhK5WfwRM7PG7yoXIFZrOCI0QauAw3
89hfOX23hLYIbFRaoMTR5OsIy11ctoopebH8BhjnpUoKxBZLo7cRXCeg4pYQiIJ+
D2Y53yDNEsuBJf+t4R5JBHUIz/58pY/4o6wIPYL6zgUBH517PQIQOGcS5lW9LV8z
NO9nQ0hED3OfX07ghfS8B8nv13PmlylPIZkKSS7G0T72G2RoQc7vbj3OLow9DUmy
1GyNqKzbY9WAZlSPB2Ek/WN1ac+FsLA5BhZSvIqsVbnpDrZxohKXLszvXPHyjG4l
z87CWHPUyMrs6uirRqv8jQZ1F/sOrb44NLPI6nxA470GDmemut48EMb71fuKG/Oj
/J2QUS5o/sUZ7XvWHeg4epfWOhPWC7kQe/lGYQLD+a2gqpAVGOg92Lew8cqkNNXV
TjByijPf0Q4hRriU8VSMUFVTbrRfwsEwQEw2K/aEF1QZ06ysrwvCSA46QHzLzMC2
zn+vEGBK9CzoeMh1+fJ3O7Bq3YDshYp21TXAR+6g+uLAwJkebCWvVxAHrpjlMsXq
QPiWERdbs9trA6ZOKwTnsm6YLFCXbE25ZYd+lYJ0Hb66nHNyX+y6G7AiqJ0eSas6
vYeDI9DCAa3nPDZQEiBhsGu4qozAgg+mGZofFHDYcNaWYnvCuGeObIS3pVFCmUGr
Cv3DQ29YoOoW+Hr6DTTz060sPwjGc7XEQQ5tkMSOKWKgwrkAGlrpB4C/9HyTpJE/
SJCzz+BMKNurPjS1AIamIhurMpN6isf/WL1qWXUFY9j2OpxFjoowld+USGEyLdnI
vKm7Cg3B6Fjtlu1PAaxd4cb+43Bhd/vSkjJ25ncPAzRprtbrz/24EOFv3bqaIyYM
GFfl6ktdy0ONxIyMXE3pEOlNi9r2oPYdUmeCZKn3OJoH/H7wFA17yXpF5+7evUoq
tqusefabaJ/JqORapYO4vw8YUyxMfzGUTXFrfiGTAUMAbT1Hy+Et5bi/A6GTyaa1
xRXALzO8gUSH7gqHFiZMgxCmGoNOUYv9ez94MU54zR/OlQ3OGtpoBRZspv0C7zUu
362p84wWgJMXb9xgVVIMnDGb58zYedDtrmbfN17y4veZXc5Wi4D+49rAQ7eXDIFS
TOMSsrrXIFWSSopsE6o/zqGnbL5iavfM7nWREmDmGY6eEhauQl6XeGW1VzX59qwP
c8rJTkNGv7v1/GxGAA1p9y0nqX5zGWP+1KiIN3jusW5DQeK7jkUei2lhAW4oewxf
lCWKziWO35m1rPOfkMjypdygjBxffN0pLxP/VBGOTl7IHW79vM/6lpJlm+anX4FD
khKQVi99sYisHUULDmbkgy1cX3DvkL7mcCkU3doe/5hhomO5+hzvwgbT0ozgq7rt
m6++8fbmVMiMCp5qVAuvU4GHFD9QnK6lhZsp9YnP2rXLMCk8l+uRlVxXOnY7n11Z
qXE+kd/Z1Iufi/iHmHstYt9UoD1zIC3atOO2TENUMRNs2FzP3DmEMNrQodW72J8O
38GKdgzz2JZhwwhzqZ+ezOQea4L1WPrf1ezHduoUYr5BaF87nxk+QjqCG/iW5DJO
6eCQdF8N2QiwuxYdobL2CFoYeHEvunJdMnLzPp230vOzcDe587sS1w590nTZeadK
wUsNyhu1KZmLcdnfgMDY3GFV5y7KPFUSqjNuQeqmqgk2TIEoZakfXB2MwZJtIh9P
sGd+nLlLpgJVIvSgNnfRvNPc6LuLmujYbEByLwWIQhA908AKpCtOGnLcsOs47AS/
tL7T68SUt8ajdXtuV8o8CUXGeKkGWPTtNSSO0xDufgCgAfjbI+CnoNCd8n+OPTf2
cDU3OZc0zTWJIqpaI2KfZK6LORxURf98caryH5RrX7pRfeIxd1KsyVrMmu7T1nRj
ncF9YrFHak8GxCV2tOdbDNWEL89qNoqFubH/awPFp9NNQ9W//WlQK9J6LoHZRGuQ
Ulxy7tUk6QhuB1/hETDx14z/TzXNBy3yKT/gM0P+Ujw1xYQQtUJuOqlcQsIj+ell
FDKzloB3xod8KElptKuMtdsqT4WxwBxNoehiBp6hB2XrXTuqtjtsTMpn06WrhMgx
qMaltWroT/NTqV4PJsCcX18nmR+dAcL5+fcgJgI0mTn4SSGOF3Ak2wV6PBJ8rW4R
CcKL2zrWuBFqmMUEN5ByqHw+Nzta9VPLhQJfysHmXdtNm7RFh2BAMnHmEneIioPr
6ATgEgM5vOKk2BJqiEkdIJY3w4hyg6LdK7G4w6DdeoPsziVR5YD2Rmq8ym7+jxAc
sUQa9GjcChaUzvVpA2Tu2SVo08iKcuYcgqS8JfDzm/VGZWMoJir8jikgtoqEWcjr
rKpm0tmFyaNohZUpgUrtJcdfSC/ZGgNxXXJxqyKJ84T5O3L2XUq9BadcYaygcenX
4gba8tQ23njo3OkzXm3lAgyrOlK+4z3RZJW2Ls1sIjzXMmLogU8kJuIJhB3+EJsp
Yko4hvGGdtjCJFVb5RcoAm8DnkYo3C+3GTAfrh5E2DYDUnVj2Wv733qF7Iq0dNJn
f4b9vgbHqF4FN/S/qucUBf6Pvxi5GAdpNjFtF5uxOp29l4uZRWppdTrzg7iKAWys
yiPHHfiNXgSzzzDCC9/XXXhGO1u4dsbx6p9m1fTTSiOedkms7LDIhGEf18NB7wnI
20KZr20N3UIyOPS0KB/9cIBKctUBdARERLASk8RaGDsVZyRXGMOqLskzaMC0sFZ2
gqtNsm/eUWiBt3CCljDlmRFo9DjYGZGbCynVEclT2s54Z1juoMKJJjERFigakojc
QcoV/b1qkeC1vx6sRzbSkXJ8aOfyXPyto9FbAyKCKqJbXaI6GvZHTvs+tz2lM8+e
7+GCpS17g+mHrBrQGRciN2iPfFuB01Klycc86xztVVqqI/eu0635KqX5360n+alX
sdyRFUCl5aK/2yLrIzJo/cHiZpnCqyfMFahKhT0qUsbJ9TFrNktllFkKEo+XH9Xs
CKIRAOTB6G+vSY89vACH2LX8hKKTk7BsMcJkDF6F4N+m+Ef+kkLPQihzR1BJa2MM
kDTYSrKBAnUS6cqLjXCiUSUEn05fib/sF4O+DB/Ynjzo8ffK683RsjI6O4yGXVnu
lzcwY+U7wyResAtg5qetzbQj1+WmBvV2lUV2kxZS6yO3njT6r0scglZIvN3+ObUa
wYcsewtzGzgfLTk8nXKFYbHGJSsDOhKc5RiqPpaqRwRPq0jG6NZ8amIkjQJw3VUa
wk2Xe30n7zWxyQHmxgP6l19PuOvGvad5BML5ERQOr8LnDDEHNz8bfqyuePUCqJmk
5n3iSPEByGeYcyj3sZHoFWs3yUeR4+85nEcxcng8MlSJL0EIUVcTnv+/fe/ia4n0
MEiBBciNJuQUiEOlpy5JFnWmvIM/L6OxwdomUsGggGlqlXyfzRYEiGvZ0C/4WPPE
13j4JCK06OEDit0owfM+iqUX0VZOSHnFSu/uzYalEB2w3bOQ7ywAqteGot9zsqSi
Tpa1ZaDa+ok+WrK+IHKWb5Z60fe990MQfz6nbbk1Azo5VPUZVkIS0oilPq6OLGeF
0Po4qcwBtQRPFGiK/PQBdc2YAOxQStJqGeDge+r7gy1qekcttdFSdZfdQoLSDPfG
MdWAhFl/St+BKgZIAkUgh8KvpeTV6+S1GpdCoC9iju2etiOj21wJgabT8uPQ4ooO
QW6Tjd/ksegIwl9B8VThY4pGjn2IHness1WryHqzvlJBPtdTjTnlDuSpguw39hN2
0WGGYmbOevX9EEj00zrHOsh154xVCUduMcDrUbJoTCtk0at0/mw+htj4RBnwPTvG
mqdSd+kAbun4khLmOnTb3pi/3U3rbol/PqWbr0M109uXv7xV1wVr8fQXi1d1Xyi8
ikFiYR2E+bCgfororVX502EnrR04Lyw2t7oo10uk/TV+Nmzp7bCb7JeBQHOmSxGw
Zp1PTkSnTYU7EF71v7ljGIyxIy0wMqX+r4OBVP6OQmObwTcSYZfLXYJVPzwNliQa
YYNeCpIGnACo5c63ozjZco6DPL1cZOWVERThf2KGr5I+RhXG2ALrtfMOfZCSTJHh
xho1+SoRMx2qVJWdtfHMLDFCmL3RrvpC+RryXEmkAeo07k6hMSY3C04katHvpcCI
dmXEhvH1PI5LRZyXb0IVGrtQ8xoaDoqVkov+ac4Q4dUvdnBXsiJd1IZxQ06y/B79
EZafhkzg+7ytk8EB/40rY6z1p61i8+DsTfw00UZejzwgdy4BxPCjsnQEmpwmOb9b
1Z1ozQKJSxzA9TTLAqimAc5FqL/FfIL9HOkRRi75zVxlgEZzckjIamL8RrMIH3RD
uAYG15KL6fKJ2FVzdp7Gi2a/m/c7jv+MjQtKqC7ugJmtqRyyQCti4FXqyNsiLPCJ
Myt3vNuk1uVav+aZ+6F0FPoNyEtfLhOrqqRL5xDW+k664zdk58gIh0KaZraI6BOh
P+55zFWJLS9HEuiR4ejtDzrLAtyhi+br7BYCmUVxwtZLML/ilr6bjt+xFY9ykw/C
pQx72uQV58xueKLTsTp8x9uBW8mBzptOXhxhjfYw+DvSdlMLyVPjaebOdMEAGSqK
wE/R5SFrWqDWOaOPXN7z8X9NV19sgFnC+k9bpG0Cx+v3/BG6PZ6ypKf6oP8v0chM
ofm7hJI9Od7dU9zAVGnMBZOrUtTHobRhbj70H5YV5+jZRWCRWk+AQTqkxLHG+TPb
Y6qd2qlfJ8nnWPzmzogeO0HM7wj3970rsO6bu7eqgoP/a4RYGLCM7KOIlqsN1Zlj
kOr6vroNvC0QJpv87MwVSoj2mIYKlrxVBuTdpuvwtZyIYJd7gIEXC5w9Slppjvdf
LZNZM+NeWad9Emws3PGKR7ZTVb3PypS/VGuDVS9muIUJAOXFPFEJyzrWN2LnpISQ
v8zEIGCdB4x5yRGUroqMOgCL+pRahURTbjVxVN3+Wy5087UiLAa6qJvCPo4dDrVd
f/r4c+QjNEHeggjgYumLib5UkSJ7ucNZTbM5D44GIsdiTJAaiKRsUD/VF23ZBnNW
Yx2fnNsoh+/ebO2swJp02YVVQ93JGn5acV/EgSiOC4DFXkT5sGK4qxK+j+hCeUpE
KZepxvsHmCrYlC2oqGunzQ+rRSBfVF/o7bhVl9lIPQX3hB2q7niNGWH1yesG2iaE
NPL4+aDZQhIKjieZEUii5JLR+yxnTMJCyXT0K2IB3FOR0W4i8wsNLL3XbNqmdZCS
Kaw4Vx7re74evL3uf09kFNYmSyghV+P+cZcWQ4/Cem95pJU6IyGE0GZwImcGfBCr
w0PwOzni0dVLi/Ek+zujQ5g4IVTvR6aVpFjrlduxDwCGgS/FZodWqlxTX0O4peIa
O5ZPCb+l25knQ6azehHh1zcI1kwJTI3sFbjruXy1HKTITHy2EDXmFI5vSYCFXbkk
EMhX7VjKVyXc9JvoLck1O7nz6XEBNenRL0dtohSkXtUoJbEXgDrZlliCnyd5bIMy
tl/ilJ2HJ/tkaBG7YBv1ZHAVrDfVO86923dumRzzF7ekvc5BGjUNTdTcXgnA4cV6
o5XBOvuzTwE5hN2avXh42Bb2hJMVryHFATSivRuxSmNoT+g+LmBApi0BUmV4OS72
6ovUZv/dEhAiN/DWGPszzYx2KN75rqTHjIaTjqRd6MGjEBPgJhMZu8fVJrnUn6RP
nYVTVVLjH4dSFGm2JS9hatc19uEOGee2qJecMC455VUoSY8GgXHEPeQgQobWJQQC
62ScqCsoKk0ROpE6Rn6ybkCY4i9yexrbgtOvBrbvuS/z2GJZAgqESfZm5NH+XYFO
D9sJoPysLg3KCOaKMyRjyFK2dqamc2CHcU9DpSpe+q4tdVJcMyTCr1kyHQKrN4ER
hSkFu7Mhx25L7eE4umcfnY4gOJN6EaYGYS4vZGAB0puOKSG3h3HwIx6wLQFxSsIc
07NrfETVh3qBGCrSD97sCvDBSSgkpyo8d61U//iiaDz7z759XG5UskaogvbEz+W6
8yxqczMQ7enpd9Yb8yOQMcDCyFScKg50jiz8yhIUtIqxxQuMRh+00DvB4aLmr964
2S8Mcf9IMBWYQQs0gLLzoUu4NJd9w68ALiqYAj40faEghvpRFMfeZbOMe0dOfqzG
C/xJqS4MPsgdQ+qc4W6sH4UPG1uAwig7Y1P7I8KR5gn996ZWumpeiIl6Qkf0yq/j
P99yJCJKIltrW9JtPTznw+Id/WY7yA0R0zuJkxuTz4NQlFKUmD1eDnmcEaYk0JcW
pOBMUQ3OArezEhAZslcYfgCe0Hop9fwfAY5Ha0mvV3ao2dfJl/Xb7HLzGnpnRgmm
oy0lQvM0+PtOw1Nd9jXJTziehN6705HkEhxSjYGIFzMR8aDH3Ga3WBuWapIClmjK
uwe4VFsasO2rIwDsThfgLs3rfvNLlFPlatq/9LVzGsf+Egk98KxO5H26C4Ustm/O
jPsMSSaBfJXJPWNswpSV6H2Iia16HJHrYn4r5Tu5+3UiAts0RkVLFR9MdKrxm5xr
sCft/9ni5IW/o65eTDeAVVN6DnPoM/uUeEkUjgzxeAyy3N0C00SdDqrWdPvnUYQL
YHWfhTbwDx4J5JQyfBD5XXgkq9d3zkgGKQo2Wi8wdD86uU6NhIiLEm5GI0vG2/lb
wPjtUFqwRCizh4v8eaAuIc+Pnncfqa4UVLRQMOuc6kXNzVwkgMZkZ9Ow5y/IL4yj
BoVBVdry6NimqZOlJ1a6QqmUxHzw7GJyH7R6AcsXMf3U+RyLRw/oxz7s0uDQQ+wP
oKsVjvNXHU0W9tyyCdIeCQWdaRAEAkyDGlj/EISBjASaYGe7JoSu/EfVWraVTE0E
ILrWIY/eswx7AaWut9OriKyY9mznnJ0wlpzkN9QiUnGLTdRzYl0jUExNKg0RFrZs
qxGhq/pw9UaJRxY8/l/uNceks9jqrazactPed6YejJmMPh9rnwaQEQEMYoG3XdMD
fSbBp5skiQnNoR3tuHQiwsvrKxzCB00ntg7j/EyupvM7Bn/QlQxIkuCanwnNys//
+gqMuRpWj7Pwv5HgYJ1YN1C4mEDu+07E3TXdyW+cWV+6IkxMNesYPJlWUa3QiLPd
zdh06r5rWVW6Fqkkhuy5rBefpvoWjxvHK3jBW7ZwRSOUOic6tHWeuvydaHn6OI4q
B/plERLEfwIitVytHlNn+/d4+5v674DDKIZGjllrY2z3idEzwMsaycPXQJ7v8OpH
hWdtuZ1EaP5+qBWOTWw21SepGeGLrBMce+mTWAizJVHego9pIeexArsTuuwJD77e
IAqfSlJtBGhBHPoGofvvhHiufZlFO0tAVkHdSNL/VNRckK6adMjWs/Rds3Arcn8z
9enb3xkYTC3XJRkRuJ4kIO1cDLMY8oEWYfWmWHShyigertEBN6C399161gntMmAo
3k3FcwcBfuodbCup1XM+8AWc3sI2fFSXqsMHl5/LGWiQFTp0gRs85ZpH7bg6nzm1
njhJGss749W0wy0WxRp86x+mmETW6k0QsAbVD/9gmWNtw8Uq72ifOPpxEUhqvDTc
GKTB6sPbM5nKiGAF2k41lkmC7+aZfL/dVLH3L/n4N/gFMGMPmBjdenpNoZ91F5Sn
TmUDJUU19L7f4avsa3PsMlwSHnhY9WF0krdquT0x3UFod9tFo4u+wzZOvf/mN4zN
l8q3kjPmEwSKdtAlw8+ecluVE9oDfDHzs6b51DghmxW1GcrqfOr4R6aduDO5SPVv
7eQl3zwtZvjCnJ/DwU1N7TqmsYgKWSFTtkgvNsaT/Yghz+BeX53Rle62p+NQtsSS
oW/zGiP1qneWNYK85K53SuGr/aZa2teOWzAm3U9s8texh1+Raw4NijfTAIrastmw
FDDXghIaVB3CE4/KWRrFmiZStw//c36pMZx1mQHikZMVYGCK9b/Jf3P/uez9Qjum
CiItEvk3f3RY0HQyC/weXJq8OUVcFXL/iJwqxXK+X9oDbp0jaFCeoI8ioWSpvshq
MdVaD9zruVI0dtRMqm1BvC4IYPDXAGWKFNXtdNo08Le5+Qp8nz56Eys0eJ6uo6xe
vXOWjOkMpB5kC2v2xooBr0VYboscXirU3T1wxz5NUBuhgd3vYP9ktUtfmRqAiSET
CUZwe5oWBX5CuKdZd77aRDgEHP7FcYckbK/bcuKQfsfyVI/rfwq/KmUQ/T6Maasn
cCaDoEwiIWjLVrJK1DXZsAU1M5GdDlJdCPV11PFl3DMpatkJ96cDjNa0azGb5BeH
eCAUJL2G+Y31IeFYfm7dXSDKr78VQPz+c3y/0BanilwzU4xslnm95sddCQA+DBvH
Q7gwz6slvq2zdzPJ2cxONhtPajSDLt9UFiIK+5x69QB/g1s9/upswWL5qO4r7l8+
yCKsdX8ERXxRMyqfGV8Np7V0ahiyEaAgnPJn95bMyVYkePfFIIWvkv/8PXmJgNIk
8RNbI6JwLrSdjY7srFI2EBxxElyRjUbUbcZq14Nb2Qz6Yw0FZaskWvxX2OyNT7F5
8hwx8aIV4N0S6slXHiOWYNVvejjm7Udlf+uBOR16F/Lz3O9wUyeFgSKvyeeVp44Z
q4mgcPO5mlhqK6fgOGTFA4UaHoAWKISIjS+ZCt+OcPym2fuBudQt2ypoq4G3id5Z
2VLmEVCm76SuaNK7UcTmpmXCV+hNS3mPR9D5IwE53CFsP53MjuoGbhPeCnJNta8Q
k2hVLh/dlu/nQrt80O31U6bdEs4Ry2EOosaekz+sHAJFEIxnzifI3PRQQQoSMf2W
wtVN15SmZWVcff93PIJ2lu6EtL5oWm6PdAM+Y+yYIXl5MFOg1AN2UM1JYHmqwkBw
5lHZgq/Rbg8ZSqgXXxSY/LsFMXm7VTc9FtKgutrH4Grsl02NUUP0OitVnZ7aiHEo
EZFHwrFl1V0Wt5Q16u7df4W++EXs8+FOIcpwmyhNH4j/xssqz+O5flfMl6wr1ETC
0L3a32UQbkSODx52sBoCvuP5+PwsPgBPo7JosCFYwBFHGRob/jgvlcwouOQSZO1j
ygf7aZDDb1+9BZ9vt0ipDouGzNAHNwDGIe5L+m6YJ1fxkjcdITCy0KXVpmor4Gt0
9/HBSJMCwic2glU12RAu2//UMIjWwmfvEd78Htxm73s2hsWixz8RzsAcs2nt0WKP
v0sqsCRXLZtKL3MvvKHbKLa3g39hDwuuOvdhiiDWQkPTZW+9H6SKbvos0nLZUHwF
lJYJqVC6ME0zW3/ERuWf29d6ep2KQ0JmxZNooler2IyK80AjaSDX3gwZ0vqpPDCM
hcMHFei0vTDkDN8a+uOr2ncd0TfRov6cxteETSOJhKAucSF03AyYFoEA7AfimjoF
ZuC0b+KLApW2ENq5UjGodhDbNAV/vaEhZzsHPh/JSFVu+JP01o3ySitg4s//egtk
5i9bARpDWpLy41xZB7Fjv7GwaRuEc4h1Q1izZFkp/8Gx5QN48jdeVJFJNMwsXhx9
lU/wYy8hPAVHabO+YXHdAgRf9OlcZtMfTBIJskqe2bPdVaBZ5PmCtqCJL21InrU/
SIP5p2/v6UsthnHDvNYynKzPbCKnbRHTwgyUBKJYGCXGO3hnrIFxVOuoT97YWAKk
6nkKSo+Bn6ZVrsk6zI28L3Mj0TT2gt5AbH4hLpkIcr4ITQnKLIxWxClhuCgV51ET
a09GVbSQcWFcK0K5pTVEiFZEuhrhbu65Qt411jecwTevDPJUkS7ShaS90kat6s/5
gqh4NZRJOjKF4sfdEyHvO8904VaRkW4ZzZC+sQ5Ro8Q4Je/85LgCP8kLYxB2wXsm
KNPwrxtmY4oLyd4ysKXu2wFoUZqqTnu8ZnGDCrlGNdS0hWvIKRHXjdufNIks0dyO
cISNN8Qnx1owLDOhNIoj4aLTExFQuS1CicFCx0oXAPJzMOvDHTo1eWhYvsgnRngr
jK7rGygeztaaC6DSq4ewcKz8IH33H3wpbTwLexObWt1jhway1Bdalc0xnNky+0vl
Qmr5LE7/LhnYpGlTVEyhDkisFyoBk8uIDk9KsQ+xRSikStEmuvv0u5NZIpcFLbvE
l1uixy10Y8/fBZI802Dufgmj7okuFH7+rqlKk86FgX+2p7/Uabid9UtMdWgVhJju
KUSFZ3avOZV7qMszwl7iqdthxuf1NRU1oEq8v7EAmltmKjG/ohNHaZAQ8m2Fl6be
+YkOdzH1qE7ZIyHQiAE4XW6+7j9WElXGVN0Ec0eV3CTPCzct8wst0aihFWweIh+E
tUht46DxbO38R719q4P7NGSiyQ6TwuXxi9nF0hk1sfC9MWch1mgeYkCFL37KwhUD
RCaZPSTLEwFTTbfhuCZW5+K9Ima6xsNQR9o0yNN29XSrlLM+aPU+kbvgJ/ArcZdq
RJJXevHgCnpN2pEz0a1tigUqG6nSNeZAYMN/cnT9GoYaNbuC9i90ergaj/gPb5GU
DZwlkL3kSSt2v6gRhPbZjnvobqfA/nBFzWBm6TfUIJJe9W6hfPPH1zIFqiIAgCg7
P/XH/l9l8jePst/YqVTpZvjoNNboKJmenZbfP4pnyc9qf3e/rKyvwITlYEVv61wZ
SSXfIC0kio07qTVB2PSvJ17OsJ6haXHm5epEepKRQFqaII5XzNSyG/nEwkxZx8us
qtFd+/NVMUVil21HzZmLbd2hZCyER2i/11quXY36eSkJopJEyzdJNK3cwolThkZV
2+jtieTjCJR/2jH1ISksDq3+lGrUEOserXsn0ixGm3iXUV/xiKcoNJG/jGPPl7nj
dV2ZUEJrsDyEwdtBAmdOW5fjDV8VsExctKD6CgkYbo6uSLOqSCr41nnri0iBU193
ktdPGEOhgf6VXkDoVGHZNF54IWEOlxRYoCBsvnhCCkR2eOuiK48FC7rjjJiUtSf+
CPdsYiy/VSx87Gc5FH0yPb9YGPAntsZbQ4yjFGufEhch5fquoqin2/CI3VD2g/mp
rK8UrvHgCGuTjhU8KaDlLklBO+nrYbWTl9eIDCVSH+xWkfhtXwqtw6i0/l0z2Aop
kwtkq3cHK0I3TPN4klJVWfoF23ShnuvEhZd4FrcLKM1NTaoJj1kqHxLoLH93GN2X
Ks6gPARGvApNvx6vQ4x3YI9jJGaOCGY9Gdd27WmyhWMLC8uK+wsLZSVZ9A5qZ5pq
+j/bHVJ1jtvJ0BeVRUQg318sbbMZp4qbm6jBw2Z+jHJ9tjK7ollrCwmcHUSR8nkD
cvRRVmizp+wUCNaJg4766DhznOvra/h0FXSlhE6xJM7ST5wnq/De5uMydvYKmurU
kp4rpPjrQiZGVtzSu3ItShOImb+0QYPDbxuGQq/FzCMgoN4uaicF+awGQw3EjVOo
NBE7n2I0kA6qohpXO38eNBx2QkAYfit+j5YdMuQE49pLI7JnJk0WQ+y1A0PHsYlh
4EZ/l0xlB8lrOkQ4+j/pQKFABwB4HUd5+RSk3tbXFDntb2NwcjBaqTKbWWUsf9uV
UfyeQZWnNtwx3htCw8g63VQ0UB/IdX8I0X+ecHlvohM3Egg6GbU0kcyrl4HIx+m6
WEnkbLv+tV08ZGxnp6YR0GiW1CuxbrVpV4Og8L/UsFumbbvKJIPdOSjOdDi+Vs76
WTcyVgz63gppW8Fhm0pknOycdkaj6xG7uDOa4fn0i62y1fpxXrREN+EQM9GmxGRs
AYF42EFU3LAtrtEjhdCiwjKqqYOdNvcyR1wiGOgP3MyjLQYPqGKbSGdT7Hj4XNvr
FzFmatURcHVd3B2WnegUMNi6ASYHPD3sRKRcGt4FrFCJkT6D7JPaWC4Qy8AXW2Xd
+gG+/1srrxvEwN5miTuP3flIpMqK2glbysPu/HkbE30aaaF4epSlg8RQRp3HBe3Y
uQRIKIjNnFU5o4sXZXpLfhIZ1L5MeBU3IFjYJQt/Ssaccgcivr4Bhm1kkIqyPgVu
T9MInNFikrju4pXLj8b8dfJD6do4x/Yv1ZhK38hKaM+75j1RSjCCM3HpDR8lz0cY
9lJ6/tC0d0GGfOnt5jLk+yWA2CyKeNomiv43HTeq33AzOjOosKaoGd4unHxZB76F
/JrDQ4k6cHG0GhKk/6Pf4/k60829ifkL+xUNKQC3MK5WcaVeEnqHX49x8lIc9sgq
mjUqLhC0QsQJeYt3h2cuqwKOX0ylN7PGMvbzRtI24uyM+8AzNvaSr+6LimBZYALS
mq3L9NPOQmpH5ekonfZ6XkCs5eI0u1fYWxUDLyqmPWmLaOR3A+8fqHqpRSvSrZlE
seHV6CMWzrA44n0jgF/NP111bdhD5y7rBgLSkkVDpjo9yklTPk8m2oG4kn13+GfV
4e8U+S1wjTv6rmedzNjHuelX3YCVXgnpurRu3tIvYHxOESx7pT+2oh55F5tUzzhy
4zavjSu+lRA5YLqZmmkQBXoq1ISK7TtDk+/00Pn23s2XX8oTDovOP+yTSYZMZhgl
ugDv7omVjZq2fxfUj4W/gk1ePmgk7RRV8fK2QPmRyYji5YMzs3bjYWTMw6IrhWT/
taQN3He67VqB+hxgq9xOaN7T7CHx1c/BOjGOM9whjJJz1G0998LCyiv4L6bU2OtC
iXrxf3FFmwQq0P6zkjChz3Q28AQT2Sk52TIL9MvLUbt6uUoqZbbtf6iw2sZppURX
O0byaureer1NZc0kLxWvFlyYDZbAzTiZlh3AAKE2iNM9jb06f/I2enN55qWJ54v6
q+U6nJvaCb+wGHzRwwwbwAbY4ySppzuB998F7C4ZYd/o7frDkoo+xCOpZTrGlAkG
qQviBPSmVIe/OCxhRvZvKsNZFKOQ1TGgLp+W2Hq6cdxT3k26Zqu7+zes/ijXnZmY
lAPP1ZLNNu8DxjsVASxqxIgK5SdnGcZs/SnhNHF+VkmLw1C2zRaILvUe3Q+H41k2
nYrp1FYuXRRCNyk3PBzi/eh1pTYAP3U3+aP08vDrV0nc8zcOFdjH+1yC9MC2qtv9
7e7vPMiUfRZlzsf2NxHKzfHS7ygyVJbF5H8v5rXbC7yB2VOcizEYqfxsF376JYPA
QvLJNK2xRvd+41M9Kld2CwASdmFXS+21Euj12kEfQscrt3GzS008dMX4zpoOcb1i
TeRBn7OQNa1uXiSJ7DmeMPbAd4/aIJ7yiYoa8RdRxZjT1Ho+yLHsCmxZGeOcHSzw
vLZJ0d8NsDqH73+Sz2jUTZjM30F20Qb9RJ7mIxFC36EEedEW4IP6UuVBbK4oCSG6
7CbfijcSW7jC0KhzPaa/kqCYEtjVlkw4p5Ud8GUfkXoOK97NRk3QO19gx2lx4yAL
sHPZ30zlIFz7dlr+1byqUu4kTh7S6cP8brgm9v1QN1fPNunrg3Rh/Bk1/gx6ozzu
Lw4PH6W75m4aV95tPEvFDU4ccx8VS/+rxHJO0YtcDRGCA3n0MRIXsBPzENxVozHA
VH80Xn9+5yXq7lo+Qgmkw7NRODN6riPs3M4vStw/gPSzm5fMRRg9piE/Y9Wbk4uS
2R9AbOIFDqwD8e4UF1bROf4ChfqizAHRaUqUuYFIzsF4CPveooVJsu2OLZnZggZ/
mw1kCS6UqIPijK0obnAdo5vS/VmJhfa6oV8Xl/S1W7nO8Ib0Lri76JPiqy1V2eNA
tPKsEF/ATIfRbTSm36fEHVITQAXMmdGlby/brg9oOYxmPPUupK3VC56e7kc+uO2t
iXGPnmcPy5HuxHcA2FA+JFXUxUbWyJ/UA8C3BbVB1PKpCUwrt3b2FTy+Tdn9XCSI
4j5lMzvwTkNfKOt38fS8ikK9RtTWOP8ll2urkkW5Ki9JqwAGmmToyMeBjQ2BWzBh
/Lf2GmxRk3X+DJruQ57+Qvh1Cn54llMuAuYVDkIVcUBWmpgOU8KT4uj/lTdrDE/M
sNrDe6BlasHrRSEiZgryv8Nz4R3EPeBMD27T9Gsls3MOclya9k+xXJ47dNW+jWt4
tYzrRQp96Rs+RyXUec846TqfldlUrvWfp3kUEvHXMVh332S5KCLmTQIi6tDoGhOc
kjbK7js/xLHbzUmmH06WcD81J9Tmwoy2y/h8Z+cPKXTFP6ccI2AGb6ZcSByMuwIO
VWqoq6HMfogyXJmydcEYqtEUzonhcZYcHnFz8M8YD63Byv4YseV0PkI46GhZh6rX
YIOcU/AV/cmARcZeuaTeK3puQ/vuKpQ+xz2tAGjaGwLZuBBHw0ITN7TXCA8b79s1
9/1RsqjpDpNDdUrdkaFL6Vhs4NvHC5kJEJZvb/148Wa3SQEm1oNyfVLtv/F7QJr1
ghotoq+xLhciKfuBwv+LnBILcxOSuZQokd8ZuvBC/CQUBIHcHfPovMex6YNinoni
OLK2YVM/HUAmXRLKo5vyh2hUFH8ri/aCavR7IVZ/x/spbLT6nQTKmnAf6yUtlmO2
r/isUw+glFIIj9ooOxohws9HLh8/+rxRkm5vUvEwd7ybvyRd/hSJj74SI92GXVIa
M4QvrV6CAZTsOjzbrlTxj1NwSuCrbmb7cju8g27t6jFGM+4TQOCUCBwzKVBQpb6P
83Mum7HAld3gMNKz+JNKnTHSEt/orxj5Av9fxffGj8HVEH6zK/F/r1Y5Qp0bVkSx
hiOt4oSX0nkXA2p/IzmXDe23n8d8FHQKWbMO9PwbfkbTkVVHGggxAYgRX3svOq4K
ZmzLcFT5LJBPggpOAZKKiRvvCiYRuX1QDQfK7A+41QPF6e+Iab+o6kiaLPDo2643
P6FiCeEQCMl/9orpmal1Iw3ziRkVaJPADtSeXgfdl6+g06kwPf9fisSiu0am6zyI
MF97hWH4q8VxV0e+bIkgdsRS9G4oFoqeG8OyjSfRjRwS/6fzzbOVybR/UhfWnMH9
XdBT17tEuYw4frCMU1l+dxJmDO3BzAmbGEzEhSw0HSwtCdomyUrlSwm47Zv+k7Xf
ivTl/WatIXabgeD0dBk2nvYA5NCPmQk6ILy0xsNhf5L+0SC5vZZE8F57WhouL1Ep
QRS9/UnM0XhlGOVX7MpBmiGC4ktdJ/vSs9GZjenDVxaKmTI0Lk426+UCkYb09R0m
cE8w2NDpjurfnP57scL5iKLFKW8kSawXT+SPYtdhS8ZKL8tii1VRB+HpHsD+pw9M
KLVm4ii6LomPLJ1SX+C3cAv8NV6o2x/6nLGAF46Ds4sMQDxiCPrrVh9cOwCMBp/0
wA2MfSDoBh2bAyRnBXPLN4axRTS/iKIlhwzwAGCnFcrGOc210R9Q/xwhLA15Mxt4
hF0dxDOsQMR5wJ2dtWuBbk0AToxcdgz9pAKhucyCdNZ0D7Z0J3zPmJrmn++ihY6X
8MsqPZ1UUXAiXbyGUWrtrTRh+cx+GRuYHZb4gWKstURUGBgkwtLuiCo7JPNppEM8
DUTIGAt84wbpP+rwh+ZvS7d/+zcK9J9SF3ySRe9Tj+0EF8omH9grSruUCiyJBIkM
15pC13kiMLisysOGbWRAQqh/R0v40UkJqfRYRxgJGjw5QlBBBWzoZ2WcDoZPbzjr
q1eadMMeOaGQF3EMyl/SzBzy5juDxrcQNPsJbbg9z2ISgyByt2wADX1V5UhKJkps
ODwzmuqi6sxXI2nVNZT96rDajnMZCumgsI9s1a0BgNdpvrgEWZB4CZ4XWWk/qe9t
2rw6JwWr3zRKaRBdOEuzucHb/qS1NGYdo4UA119G+zfw3LmQuBjR8xpLsF1MGAy7
lmQArIUFGmglKTt6WVNsno1PboFsu9VLHs0tD1gSWs9dHoj2hvsgz5aBOyiIU8Vq
BdkUY68nxs7tAr59q4kRKlSwGaJknOWdWZ2OhAPeij+EhsYXGQUkcpkgh0nvc97q
/uDNsv8/eRioJQ4Hn3g2k17PcRUm9NRV1MPYPhOtnOXUJzf2AktTqh0XLNbei6IP
/RfrhltPE3oRRNBBfVreZagiMxNkE93ab6e/4RtIiR4BPZDhZIjNx9FklacLBazE
J1h+hKDJ45faIP/s9wBIqXhubfQ9u7M0gG2p+Y0HyLvNe4thsLCwAEKuRqYC3R9w
eAbD85NLTU3AY+AP4IgiKs6PEAjLZMMYKZUQqYrvJI522mKDjRQJ1wIR5wBDoPfe
5bdK08lxi5NpGue9BuFLfNdWMM6b8jW5AQ7i+wfZUYLihYOKcy9n0/xlqVNZYcKO
vswNUryd2/W474AnsAB0O3gMrj4xjj3fnFF8p7+FeNmfDO/bQ9KBANOn/dZi7mTK
W5KGCWiiDjKg9hSOKKh8ABR0z2PppoEnJBgfqetoKqeRufYImDdHrIAacTjxaMZH
FBjKXBoig2fbYJXrzZ1IgmzoDvhpayl8FR5vVTvKzVxkUpno+hZKV9n/9qHaSkQT
iimzdLm2qNoyH6cgjTQ5ngW3e/QUCw8/uoDBuC5faKOS63U9qtGH8y975FwgEvZ+
ZQA2fa84FwIft+u/v+DsXB/k2oIlwAw5DOYCD8c6XCJhzXjns3sspkzr+ftnW37Q
VHBOx5drswfGVzAIWL6Hk3K6gecqJO/SgtzceK64kCLBOpcZ9LXSmxaNCYqkpcae
XwdUr49FCphck71uRaE/ZdPlBYMpn7Q+qt35ylzooWqGrSE+VJDINRPXZ+RKIp3W
gbAubfn41DQCOnrxr9aynFk/ZfBf5XkmmLhVJBArHsjptU8lcRlHeaKkDrL+liq3
9p+1IOT793rioV1B/R9BzrYThriqIrL26Yuz4FbQyqslZu3B3IAmPX29witG+WZO
zKtSu40N6Oq17dtpkK3srd8Qju/MN/i5CvMFNHj8/UtnnbQ16cYIsyIz4tkHkK+k
MU3wMJ5DGgsrjWVx89YbsvqHuKDB8XKaTZZv7n0UcT4Om3VhImvy9ohvE8SVWRLK
dWJ7pTCiQIRUShTVFSbazOY98DvPGqiiRV42RKf0OI3QT6aiEcMjeVdvAIfhIcsi
HJXEzeft6VqzCWLxR73BxwuYJR/mbDW2lxF/Yo06/iYl+a+SZG+SkasgQgZNonIz
PDLnH76DXgAc0ucxp4IdeHr51P/73svBf2j5X18zRP4oUQb5wrXcsR6Fd58+vgNR
6hqpbq8EMe6HGo8TjjzhLjjs5e5r4LE7OvVCqK37KWRZUnGv8GYm6egvZkfBHWut
yKSmMktCNFJKTnNZlkPdkefdIDlUpLnY37sTuzkh78mrt3U1oTbgET2DJLLk/tBH
Jy9QQdyutpsO7rhw1oV5D2GvjtWXe/CSuw1s3R4ms6lWzTpWKevvfKlOYkyqV78Z
9P62s1PNo3GS5hFdLea07oqtoN2cFu5RKSmmjAWtBYrWcK9rwpdTySPtMpA3lCEl
YUbSWjhmlsEnu6K5dXFY3xWzN3+O1bd5O6CTnLF9+rvKNuT9XAt6STtwl2sQqD41
H2DwH9qrchxB4Vkr2RVtNfBuFtabB+UzZvo7Vyd4C0ptd3glxTrOkMv8jkZgQYPb
tnuMELVtc6IelAhqcGEMorjP33i/rexWKSCq3MOJAlyfnjcr7b6ol1F30BBDxnhJ
zDup8lmy29VhmrCeKKTiza0BQA8GxSueM9VNJ7A04OCcvW0Ivo3zdG1h0vKZxlfe
5mK9Dba1E0wbcdH5af0hrLPVQvtKSwi6D8EauLUNWwoI6eEqinrAO78ldsrbVs/o
i81DBlDeveI4oEw1OJHTNQjLfm63CxncFqUFekn2moGFSQXKH0PC6S7PLeSzi5E7
wOUShze43XCYK+1nO3xaq+t6HuaBal4gudVvtH+4eFf1Ym4G9P61nBIZLet0C+mS
opJDuq+fdm3ZIkhRj+HyU3w6MGCrHKZZnRswrTlK+H54rg6+eo5H0LcRH12IG8bv
WpIimhKFWX/fFDgTgutcuWN92sZnwnTOmNfH1uM3SE69tgR9aycqBr/a10o4HVOs
dCxAXBlu4UUYX7jf8y5Ne6x81LCafIK1t04LNjEOL7Ze9JnqLsS8pHBoVZ+hBmdY
EPNiXtSumxi9dcwQmUZwFJfg3BGzXVGxiPbPp7ZuX2FR3EVZRrgPmMB9e1VgOaQ+
on+EN8QgeBmqx85iHgdqRtxl9FKaSfNYdcgoK7H6PoICsrDFv+GcYjOZRkhVrbLm
e8GW0P5fdrjOY9RqEeOErkZmClRYSPsUhE9zl4gw7fBQsimDNTdRHKlf2e8Lzt8E
Uow116Fc5NBN0baM8TkpOIcPwv4/804Q+8RmqNWALLa0jeqVrMaxnIz6TeAc6b2P
Co8cs7eI+e8xf/5C+NroBnHZmHUaB3f2umyNw8+ALOE3ksbBYS0YeHEPgwCvVRU1
kD+dyCdeYQVtQf5lsUE33FVciavvW77ldW1cmzZWDxRBbzglorjrM6QYbZZCDHeJ
HNnadSI4BN83hfG6v3nLZDryc+u/jQeMO4s2vsCL5I/o+Wzaan+OuQ5nXJMBuSDS
0jIGd8WvM2pUkq/EeqjvsFhyiGJiX3pSc8IPEfS0iNRJyqid83mgig4dKIDoE7Wn
M0yRefOg6JMGshllplVX5YGBT9JISfhfq8hHJexX6PLq0dsZHpyZ2VlIvJxFzMG/
B2Zjf55K6vESz5DCvkF7edMp/nr7x2roXtKdtfUYc+OxBOSsqZdVV78eVjVg+2XE
gFISDPGvPbRRCdkDCluJE+jvvgimBQhyPKIVKz4WPQHOSkDri9USXF5SxSePaCbv
mD/aAvUgo6mVIhGigK8wt8+4KMrY4YGdV8SkHYBu5Gkb8yJsn4q9e6kIWFXEgZfb
0aJOvChBL7nOeW59z+R16meoOd0IFooraskX3zyfwnFHEZoLcRqlkr1Kwg3LMJcM
P7DZu2EbQCwaD952P7Eby+9BL6znaFTyT4xKp0gJVwoqUoAtimGhihOsCfuppDdB
6zWMxgFpTlApwenpk7KWu+/StgcJ6saZIQBlEiRBa07xG7ifsk/NTMNE4k2DyCpP
J0Ds/POAIbnQ0ua6EqI2qq6CbAHKNwDnUDCyBABaRh1uP4xcDhKvRpjnUm+PG3SP
EleaHAsK9xblRbFdf84La5EihNlaO3KkwilBgXqWCBJiZHPjgw82hkCgDwlQmBDT
xz1zNQ5bzqFB7FntujU9R0fz8HfvrpdsFXvLtaAz8NIXF2CriDDbKK2sjBBXNyGP
mmaajTLkRk6bPbRpn0CGcYLBCMM/i461xIsuIR7YsPN75T3wXzK5ALOgiXmWQ5qg
uaSBgAQryZFGa2Qn/rR5NoMWgQ1ek/YN9SJSBv6GdzWG9vlsfxnHh9M8cpocMmtU
XuJAkfAdL3R8jU5lzHA5pjBDP63xXbKkahfOqlvMyEUgdAD4E5vQtWvpHRogcrqm
bqUeRI+14REAPefZEBR3RXerkrJQCSzXXYtaSOO26b/HqTDlkciEgzW7XNso6DVf
2r3rACyI1NGFH1XF297aLfdhb08Dm9Z/j0sb0WyNxAfVDovD3FJ24/kXv8ltBHxv
dp69GgZ71aO3atrYNW4ULCN1I7k1+gHfmvDsU1cz0GhLbJANaq5C8rIStwp/KlfF
43vXe8v89q4zexhlEYmi+RYTo56f5sbyKLh7o2iFdP9pi40G5xuKjWUGAD9qHm3x
W9VbnkRqVCLmpggeDX5i6MGAYptisABrZFkXUhj//TOIhy/AcC6wdmBynPw28Qp8
uWIRDDstGYkwIKLxWzjq5hXybn2LehdKb8JdAHIMBgz//9FT4qQ2KusMFr8puqrZ
gtkxCt8NNOcNbpAxTcQl1TNsA8vbgUkG3/TCyy5/jhA2O4SCryaEYn6cUKzqBJbh
f4lgjt6oG+LifFqtSOuhOZunfD4W0KfJS195sq/HIyEpVnTVcY+yZN6lbd26nuPA
D6DqUwDycyBtxew2EbbQY8O3oVq3z4CyAwmcee3+K45XTTSoHb7KPgF+qel/Otw+
zJ7fj2X0m7BpkNArA6c7JAglsyteke9pDfzg7bRNK/BOxPpRgnymzDHwPJnwI1j6
BGs2Fv6rXHf5ENdqNw7OR7v6SXgq/W816QNLWDbQEftCHGL7/7go/TCyLY5gbg3x
hqm5JisULDlWvfgRL4r7D4gYENb4ujiI6d9qs/kGEu4t5NFTPQy+KYE9W69x256g
9KK95vyPRd50ftbiLz7AlCAokwJR0mq31VqzGE79RD/Waf+UVgOHFS5Vj5e42NpE
o3FOgxAEPgeBXJjLPnV5xJD9j9RrCpRQjTXKDciCfCqX2vZCHowfWoQBoDxvd+o1
yq8iUGeyc2iF3QrXBWxo881zD0FAP6XYYwO8lOYHuQ7FE7icNT9nvC0V+ZYfgrxZ
9ENmW/I0dN6CAJ1I8Ywg0RQhyIGEMdMuxwG+/NgOVK9uKv8aKDy1fX7bkxzQJMJe
OVj7n5HvCUzrPvqJc694oZk2jpBP3Kal/pTv55SqQ9hdIblpSpO2d3SJUPqWz3zl
kndm0GtSytgNVdC4wyWr1pw+floHYiVwjsXyzOIOdlZ1yeZxFdCFgakm42XiB3Da
ivK93nBXdvTgTIfytwfd8Ogvfe1HDSBOlHmJ3qYDA57A+Dxkudimutl+vgGyMiyK
42DsMKfMwexiGsT1MnXuRWLwt4U9Zq24EIgi2W76AMi4wBAE+ZC2derBrlevPWN5
E5EKvcoHzShi7a0b24OjapJARQRVfNkZSkdnE9eim2utspnb6UMxk+dhIgE9OArz
8VusyA7c5/Wx+XirHReiNz36GbcYlJgeFLU3Q1u7uTizMJgZhwCjGnPuyckmVT+x
yRmoa2eivkkHkRrx5FEwCe0UOwXGwunYlOU4StNsVvAjsHEsFYXtAG1wRSU0Lo/K
yTDqCLafxeNDnt50j3kDb8KLNsNoaXX6NqEx3x4ktGfs77DzxJd66nJPpMT6ucsa
hw6FMvEfBkb33noibUIkRhRbvvMyTYiy5ni3HpNmEcGoo++JOkic3jpWB5Dc3zTq
EVhy1as0OCx52vcf/DvroTBAc5fIqJM1fnLoROOx1fev7LSpmLS/Ft/vwnfJ80xL
OkUvkGtYQNI1sbA72GTyfAEZXf6V7p679bCJ/jMfTzCNHsCajXRfRSGJqND0j0U8
vL0IejCEgVZq2lSu+9cZPEt60J0U34eWwAjbV75ewVpCzYw1+Mfrh6gFiOB5mwDL
eStr9ZcAXJTqmkE8O5JvTFc1UpcyyXHWKCkyEUf4u53R8gZLzXROngqTDLy/6Rbo
By1QWal1rDq9YSk36V3IvXFI/Tuqc+bDUgkcwWVF1DOs5os/9V5y0EbYZQaZBoZq
0ZSVdihTlysMwxXaX5GaMJMKQizGWdLOju2r5n3AOKP9Vs3a3WlJ4FhAdKEfDgz3
xISlOzrxkiv3QucirzsMqwFuU8j5/R6hjJIs8eqxiHk0zbo3e6UUxHXAnFs4/bJI
sHMV7tv8WbZuJqdGNXvKSuOZEcQVBR6sRQ2f54mvN8s064EdsSK7/JpdYJ3VPtIb
JW9shdrJgiFkFPAITrrhZIC/jbrm9qIzc8x5CXcXiftxaUkuhTT6UBhL3Fr9cnvt
KgJ96Vjt5z9n0n86NUEOZdgxLu2RwP+S/abQU0Af61K/y+Qi9SwkI3ldE/er1pvG
9RpaJ0wpOjH92oykfLApqeOuMsr/Ep0ofS7LRuEqKCdeNVl1WKySwMTi+7Mm7bPJ
N2TCoBwsgF9ZCcUlnfRWXG5XhTByl/YYx8Abgf+NzYiDaipYnCZZNTBLEbrk+QaH
/1mR5cB0c9Az4Mz9D0K+CUw/7TuF3ziJ1yqoNJ2CtgjCV3lnSEaneXVOzYuhzyC/
XCu4uMrZnBAkPeP3V18jffOYsLjqaKh+5Z8+QeRsO9XdJT8H73y5pCkMohC0iRlC
Z7HC1gzODZMPeWq34vUL/nIoEmEwofOOi5109H+EkpMuJvQI0kazhUrCnz+PFyJ2
foFc4R0xiVLwyGE7gcTWA+joahntsXZZpTqS6zEUrbxScREoaXX/+SdC5ubSysbh
H/qOv9Ccj9UE9821+dkYyYDQU8l0lAxNz0IcS0tNh9hDaPVvTLZ1mizKqW04DpyI
dTcA1p87iMEVdhyOC++tkq54GI3m1FO5ldIisgvN8tTNDZUHs8dF92nireulYnKp
JJqAr1f+8ra78TX5DmHgj70Rb2NIhEvPPOae710afAKNvr9W39MQDPthWnuLmsBC
4QQuPzQ3QKJy/kDHDbuNXlHVOinRntHlNywT+E/yvdwo8e6ba+wmwhIQufSOUXJ4
rqMebB7XfeFoCh9x0UrHlYKvS0+Dj6C1DNAyucuelLj9lBLRzg9yO9ow0UZahAVb
Mntj1j2O7GEO2wUILsAYpEax6Fb9JDI2PeDArWt5fEW/on/Bdx2EjTAoHEkqNyNh
o/gY6WD9ga77Lk+oHVVeYwytiMOtd1BwpfVYLea/zG6kz1Afd0R9NdRTRBnoNmjH
DvXbFwWj+JCokzWzvWqXFUPfS01AEsRcKdI6Xgu8PqJjTw+6W5bihQKIIBffsUb5
PMhjuoHFXm2dQgQ6LjbUSr38fERHzYYzgJR9WAHUi0O0N2L+SjPk4xgUK2a4I/l3
WzExRyGTqF6hgSmkorKJcEqHV9XRSAAFQnvZNTqTSJBBXucrJik7iNCjpKc6rRhd
Vcwknm02XhU0WymwmYV8bv/NOa44YnhQeCIPvqSOdQE3wodiyDL6WLVeMS3xC76P
SBfrBynULEZDuIZy9zV2yemgwjpPN6k7GDwaRJy2nrTcVsiB/+icz0cuEdO07WL9
AxBhahKfo3Tk6gj+GumSijUUR8uFXhtp0qCBOVQ/MX2KtgILjXqx+5wq/1SESN1y
74TMsnPmBCo96uzQNZwuUzKSW7qBMA3OlyYbbniXspiIZezivty/xI5GWOsna8Wj
bYMTUdxMuJk62fXqu/ht5qYAz5VpzlaaFClSmjCkPzNCa9WBy8AgwdtGzRBEL2hM
+CpgqFUipIDKwURpfcF38ECODTgs0eFhpFWy24m3ID2zAxbT+pOwy+th+KjsREra
9veqyTz48qrCjxQDWJX+2C1F+c5/vSGl/p+FnnlPQrIUrcsWoK/VjksLqfcd+uC2
3M98ZQn9TqDVDmKWA8UvUjrQjmSbdZZtDqfniL2i+/wlIUbh8lZYfUKvwJUwY2lp
l7cG0Fje9YYU5FLBpirclAlm66URZMLMdez+QOK5WhC4KQe5MYM5nkg27sPE01La
FSCNtb9nakpappBHieBwCVHaRei79Asc9HPGjpgnrawgDYHzRRtQhHJxYrXO0JPp
hTMAMmWen2RylpqFLImcAXsNFPrLanhxVhk6y33a2HHtgR+x7+BFGgXDQP2l4zel
FiyEyrmjtm+5Y4AIXPiqw7m4FRy8FEYVD39AxvMfqQ7KnUpOGhaRpFwIVukkcr1p
we3tg6lmQp2KduXnsZb1Ok8DvJ1dcr1zGPN8bKjo0DhdUG5LnDERVtAN7+ytt5Tf
vZT5jH7R/kYyJMdaELr3+R7qIIhKcPI4Ab1rZTwWTHakChchEw8/EMekGizBVaaq
JuTMjk5cbWehFlEuESrgBxLtQFCd5ldqEvPIHwonb8n2Q6r6+sRTMSpmvDHZ9hVK
xOWYrLKE9DKWmfltTa6ihtaooE3aeH1LF/kRZd0hNVMdtpfxwLBTJP4N6ah+/9yo
HekLM49Q52faTOxDrBlhz3NNY6mtVIl+BrDSKD05cITV+jtfINBc1phtb3x9zNvU
JDaTRg+k0IXKhBbFph+liWz3htUu4VDTk3RfkCfsjl2NBW0YanGkXBbRrIO9cIS8
eFTLUN+PwwzGKakDL4x4NNZ/CwyxjIYqyEXy/BoD6/C/aVx33Y+wQa1u0WgIcR9G
zrXZnzIjpcpGwh3f/7TnnmA1WryERAV3Y159Rve1DpTJjrtY9P0SWv/+cUYhLaRd
BAuNRPAaRfkGdIjKCavzvIiqx/HbQoYoWjmrGCjhKoFG2wincZx2BT7aR005pljr
+/9CbxJMPtZj90OFI6AwqtzJemeySS868JVZuGH2FMg2z2N9z0OdiLQ/w92uIy0P
ANQGEbckYrkM/T14cejt5dp5IZLDIR5a1dyFSR+PUAJDyZK9GPos9mjb2rvl18Vv
gQ+nNlzIvgdDAkIApt8QT6UGPs786/39NJ3QryWcXyxxcjUe5NfQ6Jn4TFCAcCtB
oSwuNr4arLNGTK1D1OtMiaLYf5ILFJinxaMJCyfV0mkzkQtBxUZGre1rSV4geJIg
BWinrBu7Pqf8a1naxm6sHxla2l6T05qurfa08A0Bu0cOut56PklB+QjDV04lbk81
y9VbxJB7l+ulHQFi53CrFsEOzlZNENrigFYhoLjgs9jJnKLJHmmtbUpCrQeoz6Mc
FkumHJsatjbk6kCaIXy4mrZjLYItTVHSNksFnPBHpts4zS8IeOJjcBANyk4jh+mw
JcL3zmP1/QttRMOOVL/sp9lhgbLLeq8OEGxTYEVOglwbYmw2TUcwMkJ4wbH7NBmG
l9by9Z2d1qlZbG7mqsg8B5c3Fk7lM5lHOX7ONhRQnIJEXAZv0qpMlqKEED6c0xQo
EnPOXybvrYeQzJDSgjzAbLz5Lal1xC+fdIxXTUyq9PwU+iL0JjFSp3fA3fAucW/s
t3DGGvmcjD9euA3qBDOJF7bio0wyq6eu14you0j16R6Qlxy2uFP5zV+TGuXBh2GG
CKNT58Ar//+FT3TdYiGTks8U+85kkp3xFaf5/4EGN9ChUBV6hAeE0hmOiSC7RuX7
ygqd9Zf4RPECgFyOK/vEdAx12kGXpBCm3PH8XGdrTqFfngSoOOrr2u6hdotE8IV2
6Y70+6zq4NQR6vQHPe5VBeLiDl/gq8pfQqsC7uulqrTnFJY7mwpIpptlG0yj+6UI
tpEVEVjIHbE7av90S/cyVIrzI09i+yMZlruh6lB6L42Lm+xf1D45LbWfaQ0aNtMy
qyD2oFoA4FClUEpAXJRzFn62Rif9Q/U1sYklMHNP8Tb+3i9mGDHobt6aoI+zKnlt
djpXYH/6l9nInAho1w03p/oGDqlSbCmbV9i/SjlrVOCydbFEz16EYy/BzUyzAaIE
YYLxtlbr6d1VOQciT4ghw4Seb+DnbwXUfcYWIPbIxR0BMPLhTXnHS+3TwM/hYZKh
09c4hxE82FMskvisJidt2YbcgEYWSQ3y7kHow4wECsBVkuqSIgWXaU+XmnqvnndY
CtvfPBUgdacchFwpVsB91fNbXxQVW6hJUERQYBOcGNzExtF9M/DJc4MvN66si/V7
JCJsMw/CYhIus08ygDuRCtTj842r1kgOSifYUFW9BAFEljIKUupowbGjJrgYMEoT
WjmRAm08iFeQdWMMJDZUTvyughmRLRAs+1TL57FgMc0KCYx+ieYUJEV4RIixCu0f
S4pCq0/KwLFNOKg5f8Ptmi6dCunIrVSboFwjweD5k+4Bj1+plc2Ox+Z+5lBkiyrV
Gnx3/JbnrQRKwalluhsID/lkULWYFWafMTmiiApJW7iH0DfgLpOf0nCkyfwbh5hK
CZk1Ebdxf5WGdGnXTZjBCZABAGm9ILEEOxkJm9m8YxstFF880BjuYfrtUBdvsoCz
wtIQJEHeD6+PLOyZRhnV/Jv4ASLSTY7Gc7rIeZiUbbI15KzgdZ3PGgq7eYZ9rwWj
3T2JnOj70682TxANXjuQoWXIqUc8nwCB+QOeQCCHeUnddPTpBAbPuemOkNDdbKSM
1WpbnxOyVbtaGVSx53XNOQELv1CuWY377UAdKxEER79jP6hBdItXlBdl/K70uaDT
Z8VRco76WhXaxqOLlFgSa3BTTJFTOylx5VOzsrUH3phgEzuzzIrnPX9xuLP1eZzz
icHeT/yOJrI4oMuh9ut2gQzYplwpuCP7LHfOmUVg8PA4fHTsJGazhgW15v0eGWO4
uxeib2aqneurcUkH5KXA2vSJREXvweveE1c5yzqwwAoItorFYkzzEioBkqM1yxWK
2dlTCOcqTOlCa9LeWTDN4FPoCuKu4Pdw4vaYLrCd5/mnOzueCvODumoJ8We0JeJh
i5t6ALNJLnt+DfvExusyC+8+YNG0bYU9ODeu63PvysSdMTTRsX+IODVmK2yeWCH1
S1GEWOqxypZMrDVCDfzgkptKuwfgBmYT6i9pOlJXgKIQOdDSZG00J+Qn5en8kvMr
tUVnwxzKRwgO7K9Tt6LJH0J/bI7dCCgCJ4F9SapobVJ8pdSN/OZWmj1mRiNP/ZRS
RnB4Q1/TAOtUXMGi0yK1xpR11xFUKrgwPQL8dp1csn1Rt+6SAV9zpNrJLua2hL8d
1rOeyFSckPQTKzrin5ulqVm5vktrIhAVvCQOsbNzfd1LXXwlUHmh7U68Xx3v/Y6I
y152QZBdgCJOrLfwXhlMSaFiZCB/jmB9gImnVeGspusZpHsztvorYPe8XKLKPkw1
etvjO+802J8F3DXzRWLpJH6iYsIvXawcqlKk8Wt7J+S8cLSbdzsIfWgQUS3T7aqi
10Jahql9+EcAa55C3+Tr91XE4DjI6jghaSb41avMMbFSCu/taQIpiNUAl0wOloIK
VJzJD4e2m/BIRx1zla7UUDKSS6IxZMUsOUrwN3DID3+7E/5/crCMuH8m6ikV2qfd
P9GBD3zvQoR0SwluPYI0hO/+Rvd7JU4ei3BoPhST4SgjmIpgFJqLMioc3um9QoGL
wO0+FKSKy6xDg3nWAwEzCydoRX/8SWwehXKkb5tC1UkB/ak5P0EQXOde7YgJCzwC
FN11cAywRiuf6m2G/6MX+duZx37GTOJwK6RcliRCFFPoOVbuOqjwQUlKGmCDbup6
VxdaoORn8iTEEnm/B2j9is0dPRKhdddKdAI0sKdHTUMGfGM5mrHB86N5nm7ocgxi
YOzUIWajWoz9jXHMOlp8GvTsMLQOyWhTfYq9tH3oxkL9hidu98f6mkneA6PrEIfs
FPrwl94b4Y18UOhb96RL8R7FE8G0SAJRYrViJdbnM3LkYmuEL1CPLrBex6OJpvRu
WuOOELMaLn+dwBTDDrHLPTdF4e7nWzZgDBXiXYRrQ7F6mPcI5vN9aNOayp2pHIM0
+zZEcqLYM1mEqcVqvvt8zQWf5kXcp1QRHO2sZqu8mFxE3us+W58jBR+I0GgrmZ4w
C/oR4xo/PBjjeSI6KiS868OJahb7gnk9ckbPwuXat8ZuAtFqixEXqsBUZl0YRphl
76swddfhLOpwSa/i8eyKsevgf+BPr0GSNYlq/oMV/tZYmFyuMriTEEM2Y0o1ic8f
Jw6NlmiMPqfcaHddUqofOoeV11bnhBqc6aKMnfrB/HaL339rS/JirSzw3ivhB1tQ
7LMSGLpcXF9Nu5Qbc9VM7Lo8VhO261jRb7/143anRBOhwc0aWaqvVeuvOGnwS0tA
/rKlNo+3NRPW3h5QCrxdO5d7kFjPBbH50onvesF9rYzpCOIkF9RzHK5fZL15Cyr6
1Rk7ooUMdJvNWcsAsaN4R+Mx3B7IOW8sFlLxllVCdyS6XS4LJ1PNdW7YpTrc4Qrm
XPVrwa+KNEjCZBoomsfqZxYdy6Ol4mpnM5DKRk9Mj9BE1vF8vk5SdOIpvJiZZhyg
olIfa5ItMARZss/36064sBSI1UcHT8KI+LSDYTowmlPVQxJNKCUI4CCcFEsN7fIQ
C6dC1EX0/ofKZfVtEnZZBE9EE0LjUunNx8ml8VSni+HvXKdu91oLnwYP99J3gEAM
AGB8aO3H+MGWlInG3JEUoK5mBHtWmORP3Eiyle/3D4x/Uk4UVwTJLUgy/MR+uTxe
QSTQd94yfIUUW2BtGyFJuPBpW11A8ybeL0s74tHLDTXP1zRofxsbxYqp+CgV9lxE
6uNmeyZndlbBbrjDycohRVZ6sC5yWUTHdavaUMJYGK1saLz4whszyMOquw57Yuxc
zGwKREcct4gZHFo64IWGAMOX1rplmnGXSPTAaFRolryf4xu0yoAc/K8WkRJ1RyRJ
G8l0R41cVvey69/SCXHzeA/9QNQraO6n6RsRjzzYp1BXs5n/gusuJGQny1YeydDe
zygF3nCHsEQWAe1P8JldY4cuEVn1/G1QqbkxkKI+Kpebv2G8QyFEMjrLQ02h+EN1
FZKdzGCW9T8E8pIFYV38PoVouN51+j9yLVaT8E8h5+p3ysTWSkcWAVx8Y1+HQlOb
jPlEtG6wFgIMVOonBH/D6atkPntXl0Bf2PT9v7UkkkymIoewiJgGbfOFxfc3caOr
74yWhxKFeQXXg2LTQNFoAYiQCBHYcWdi/cPNd5pT3A74Hbp1IIsIeJ5sOzMgovJx
butMj/YoTPcmJNol71ig3C/60fqmNjnkQfil1LZcd0H1d0MkHQ8gMXYbzjLbt1+Z
ozjpPmU988+IilnzvDmfdOK6x0gqPpXmY36CYc5nDAiYWeNdNaxXtwbKxhomiiW6
a54pYw/zzJpyMOOZZmbBVa+yk2ywItbS9Eo70IgYAZMz8lxHoTHvHd6QXveiIELH
6EE/y4/3nMwSC5JPAhOjaCeRsAdqb9LxS2GhZMynwX/EhoIbODu6dMid1tJ7yWAr
ivE3Dg5U2GNu7ucS2PldIly8dusnNJ3iA4kavWrqvseac4lIGPYycwC406Sqgywo
GHsHhKZdqEcnFoUoNsFuKu0mMSHnT+EAhOp9BDypJ8DolcxRriNI8e+bzJup9Sox
oUnGN6XIhqguyT4pr50xoXf6Dau06yjnYUDUOsU/EmYfp+BxbiJ1X4h0JiYgcNTi
YpDOLr5cM4L7KZty27f2L2mGmLIPMQF7jwRPJVoY3rIHYwfmXgTXlOC3tKaz8WqI
n1CSNl4NaiHOxutYrs0891KWez9wEBC2xFx/iqilbekjkJXHTtK2mgerTtkz7hBC
ooJtuOYa6qm4Uld3xd7hqh3d9M2EE/1B6DpqsroUypIyx2tUx+7S/9rg/ubalzny
0rlcFVTyCJE4BbyilJcddNFi/1qNbMO1CYgfkAEmLAGZpcLcZMR5atjMvvDKBxgm
PLCiP9waeweBphgKWRoyEdq44HrlUI+sC+D6xag4WasrKE/1Koh5gXFOkF4+p/ot
hkavF9wXhPeMM3VfPNImTEZty/EqegIQY6DvU42k6S5JRJEiso27c5aLnlJLQMgF
ni49a26CwdjmlyonxeGqJku6Ftq3Cd0ozYxy7MLhV4r8Wv6m/ilCuVX9ycBzFWQb
MjXwflyCJMDKpMBkdKHYfrPBbMVXZ0aBUhMKa0y0IQVmYtkHWxM6AF3WJmk1fF0X
s2FH/j7AExoC6uyo2IlpnMqEco4HJv/95XDx1XLaVFj595kVwL2ONdSZBqcRPB39
bd18y1Pin78GuR+JLSgqYdKkrd/9px4Uj74wOfSw4mri5VS0l7uPsfOytGEn9+Mt
nQmCzTnubIewlgWqlHIEGxYWKV9PvFhaxHEfvdvJQyve/DoE3ccPe7P5V+hm5rr8
ObhpuGdAYt1kRVB963LyAKFT5kEtP0TRPvsKZLWCi/EIOUgSh9NUt+91rek9nX8B
ASw5jiMiSGExu6UGAvKcI1wFMCbbV7I0wXfZLJbHrgedFoTVUJyTHUsZtLqLBOyR
CUbz4A4wpJ40Rv+9v20DrUqlzgc/jPdVmc/3yhjO/0M2+xjsH/W+U3hxhHIe5auh
dLHNSaF8yisOQr8Kh2dBIsHsqPAvPHonodD6068FAC/l29tRZDNliPUfjN4mziFU
RQYoz0bth9W22mwTTky00KGzoBuIq1qZHVBSDVeHV0ABntjhUQ1g5Rro+ig25Vve
2zKNxpA0yh2rMFzMTRG4jPRotBs/3lHhi0MMk9tF/kAOtnLVlXB1KHnkXea0V6cs
qNwXUWuyxctQxYkTRV3Xh5+rVBQtMnKPp3T30YVo2seswytUAEbQ3pKaWzeZ1SE+
TuSHFYGrGaKKc/yQTZyY+CINm83nORnasZznQq2U5hUNJDmZh+PHbKt1V2zEsyiM
WEbnNAGvM26qsiZd4RVfwdb+VPTxkeq8fsZL/oQs759sE3GHHQkJH/ubQpZ4LX8s
PRAJ/zPYwLIl0wXzzdnmkNu//u+prNfnosuUy6klaBuC+n6HTsqeRAxmCWmIKS92
KdtTzy2qhWYYZnFGDUlpxETN0VS9LRUlLjzvwvV1waMbenOEQ15ND2PRZnk1TL2J
jEaftkCxgVaBY0xXZwNzmOtXzh0kcj11WLBFLTc62QrPjZ4+p5o0foHsYvJdqXfc
p4O3QDsHImHKUU9eLrc7qCH2622E8T66n/oleUD4cjT8rcUJ6zBLxgruTWs377v9
37sVYoU/HqTo+pnoKKZm3zv0L/nMlxJ1rGvPnK+iQUW1A3Nzw0QO1Np7gIBZ670V
G9vfANckTXPsEW197+jsgxY+i4M7eaGlOy9HmvdLQEwTvvfhSvvOvvBaqCV8VPyT
L8/oReRhTtugHm+u7PoIv/uZIOrqIlFBBdDnhDcYPqFg1HVMR3Y4c5emQ87kx2Ua
Y1NQDke3JEcNekQ55+HwAQXdsE7PfXEWGd3fIwM/IqmG7Hw9pPeL1osSCFnmeHVL
zeiuCh5hu/eZ4S7zoc2bzkq2Zljzzl7dCt0CCQRQS7YxQY5/U4nxJNa5dSUgfrf2
OClOH6kg34pSTnzLltCz954aX61hCUVRc1mWFTKcDW/neevqmvxe/iGYR3mWZK2K
T9D4JGhGHXQsMVHgMyOwdbeFSXlEFHj4QYboKMXENJ1F6mmfvfspicCvBiVbjQvT
pTTvoWLoQIATPCgKdEeEowpZgCN5zubr5b0TuIuM4ganoOSyqqH0QeYAt1hZ2o6d
AdySWpR8tbU6+2W44uWjS74oNtUxlO37NhTjXAzRHOls5B/7KarmrZ+U4mdbPsJg
EjX5MBR9vTL/205PxSAit+Yvq+CPUCMiYed9/2AXxYc/02M0PH76mhMDjiomHo7M
NV6+LmuXND/slDL+4BfDWXliqicvMgIcCgWFozt7IcbmpLLOXwKtdPYBHqhaJV+H
lr4wDOIg3WH3p721lKr45bR6eI+Ao8tNpKlUmtKQmo1Cw3OIem3B3fYwoF4U7ukU
4rg36e/6MeItn4oij/8dvIjTIk7q05wT+T+tOjNQ+En6XMZ3v4a21cZl/+3gwCMb
RZiOksMSkyg4EJk05rlEgL2GPkm1W/DMd8GSvQQsZ43NEyUzLrrH8eZlkvXdJgcF
atTv6DAHsP6dZlwc3mM6Yk31ojbjVRS7LhJbRxoNAQohGrOj9Fxyt2j70LDaaJcj
ReLSxms0F5nXuoO/fyu4Un+MwwsUioJh5C+pr+Pvk5OXn/QS/EfeGJNMRE32GQmb
cyDB5fAus4B6F3es4IGQVbXfyfeDV1T5OmnLK3K2voD0PKAeP2gnSA/LC4mtyOxT
eeCL+Y4MYvFEwfA5Q0mHYPdfZfWzoQ/XqYEJCEEW560oLWfQ93dFhh1jw4Ma4pKY
n8Fojz+E2oqZkUpTR4cdh22kt3FkDFZt9lng4RtYWyicoJiRHG5hOIiV3virdaw8
qQbSPPMsh7wSqJxME7g/TaUhOYlu8+2HjPId6ilbtmpkboygFqBbyQWkxOuS8VSE
WHF+qujbZZyrozm9iZjx+eZrPKzj78WsZxeHbQQFIcBrIbgep0JBv56Skxprd2f9
Wix0inexrQZKU4YyJXNerccoKq5+NfnnxN/3+LOiyBfnn1qKLiTYKtcUNP/FD0Ai
X7DhuQPbcErQEWSKVPAJNJg2hRrXRfy5fYO2Y6orxtURzLgBWyOuWv9n5BV0duPr
QuUWFG5rYQdEaIg16TcTp4HBOlKbiVQ5JTiHkEWabN9qTGDvUQgYt6mg5zpXcJPd
8juUPFWxLpNHxrBBG3yQuBhyerlVFEjo2Dt02CmfBT5SNDukL8A9HQ+0xa1JHCTu
/NPjCRkbqzQl4w8LRJ5VMzrc6TDY8IppESpOZJ67rBnP/YYMWNcFe/hAeU7+iF6d
hRySGsTqYijrqMTm3qexdVZ2AuzmW68GBhmptQt83HaEJJ9GVJecEbMFlVCtfQ4k
7u8tuTFrbDLrD7+EIFetylDDzEvS/Dln268PPNISH48efkjebwY/4qVCW3psAwgN
G64ZJIUGpup9Ck/2II8IqXxtf4LmTQl2YZYwuNtA3WATzpIdgzShs+aYm3y2bWtz
luyxhEYD5JtYlFmShiJier/TbqInYfXO3ziG8/GdqBMRAdjnTHhVv9wG2vInr8Rq
JBsZa4dB4E/rTdeiglEw4r86pdrQNjl+mV4n0mb/3zvtpW+gJj+QhYK6/TpkWPFH
pBeBkeTWjKDXYAykrUHZh6bouPEh/v2HyAgMr2022zek0TqHWZsSfykWYJy5SDqh
NnA15In1hBNYeCFZZGz9eVzAPL4SNdDFOE+TctGmW6KXQgLhYfWlN4OKNKSIR+u2
98d0B/j96870SmFvmvcv66lXaYrF+rVvc9AXsX3egJWiWMvURUl01Cet+n5fSWv9
EITKXXvmFsji4f1RmCpnoV0rndkhX3D5bK9C58+SGlaRZ47qRB0Vp+swLRYBubuU
BKv65868wUbCWBopePFblEDXnmDcz/W2fOw91OWNRjdXfdG5ueiVOa19zHUiIiKy
hfa0kda18e76MCZONKZLn5teYfbWA0Xy0SFCmUG2Yj60iR81dQ6ryzMRZkOhpvWe
rxfVif40sZrCK3qL2SWDjsov63tgN592S0dPvnc95BQZobPqDBZh2AAgpHAopnOr
EfyAUVzokcBjKLovcuF8DoGIhyhIXSIFThFJfZRHfkSCbXn5Z4WdogVKvsUfG96O
V9ZUEo5h2EdKVGWPgwH9wVtFs8xi9fjfj4VRG+NMPDILNP9WivCMbd2Gf8qnv/AM
aDmVDvCRLZMGjQlgw+6uy2Kkz1Kto4wmZll6cBwpInt2qN4XDTdyfWbW88nBRwok
xvKX1W+MZZsXj/1jarDnzxQVQRFJITvJHMZkBoH/lKKjgL6QEfckvWD+f0DK+PYu
tTgE5iLR6heFrWwgHn5zdbkPrJ/XhTexczF1CXt0RzwE2oOKTTP51rG79iOqE+iq
f7A3H2x3toVGKa95SpYCe1HCQ3CCEidKyvAuFB6hSdnhxqDQHOn4OlgCIbYkTdo1
GNSNgsJNrQXusj9OTQJsPFlydMWGbcltccEPpY6dxVEjxobiYxfLKtwRurrjmrkq
E6FCnMcD+8WsF54ix2y8K/NCXCVMrmoY/XypAnC9DaiHw8ziyAhNbeKFl4EfiOik
nUPupK239hdF7qED0QVtW5pVIKe+6Z1SbEIqswigaCoPHr2PyVdP48MNWCAITdLd
dViIlIBqWwsSMr/6x8KdqpNEaIfF45zgq6argePrZRb7JXuDHTvsmYiAcRktKxas
3dEgB/A+hECl2FlrOJmEATlFClk+bt/5fJXd4/0zXeVC9kkN2A+QqDZf7o6lfahD
3SHc4hexcnJdCzPEyWFgRJeOK/SrBDxJqxut6U1cBfi8vMsOGlc+BbLHwmhK1DGb
lvSkdYQc8zgauNJ8A91edM4jroE7X4QZlk4TlRD0+fmfiDFrQL1IKgj8NNZUdFuK
JKXVWD+gjWC1AWsL1idmqP4FwY6qYCjhlLG17BsK1ehUVuXLgoHyz9t0tGMbWdIL
AUcKxsY2evr6Q7COTnycbJb7QGWaQZ943NO+RVYc+cauIA1iZCskrGBJAztFNb4X
vJbQt/sJoINmiAFJoiRJys4VqA/1vtFXcvxLH/eNbqZ7sYJry8Hpx4ajY7tyIbm6
3+GshcgSib3dNodpx4SxYr/ypjuwWIvEzlos2JmGvwhVfgFSLvBzNblZUPnbrnuw
b40EAq71DPTCIbysNmlMzG74J6FlutnYtOHIKaIUwbrta2GLvmGra+hb2ZDhXOvV
TkDOXm+/UXfzHYwou0jz53b9jeXQd2zAXg0M8B61JQucCa36doQW55sSeguQlq8V
P4wvZfNQIFeZM57TuJsXjBuP02WoZMyOFbzrl8zmw45r1o2YoTS5Z5QMq75jj0Oz
aEYxUSPCyEUTYtzgCixVzLJmzHbIORI484W4AWqudqo+v0Sw3NyRKQOMRjwmIwe/
gefmBIzzUwaXuUYd/ER0+SW9MHVZVSzCVU93Jx5nJlUh/9WoZGT9Ldxlc+nvHb7y
LxEjYgsfrGfEWUUbWIDmst6xABInrm8+n4unNkNHBFfX6lA8uArmeNHu4Hc8HkZ0
p5b89uOT2JiWq83kFkvUs6Ope8vR+nMahO9CDFwpvRRfUEOiH9kgNkBVEPAeHb3h
hTFYTPxh/E2pPkRpmLzFoDdQpuHqp9iiUvofZA48pGQInc8+PLbO6Dzd24wVz6Kw
r9C8W1JphalkQHAg1KC/V0T8mC8q2FsKOZQu9MEPUXnqZTepWZA1WfsmaabQa9V0
xdCwDnF1Z9G73Esj3XdK8dBzYsg/Osk815ro0eQ/bM4irvc4t03rA7EuYL/wi1ik
wlKyOd6zMZrNXvVLSTi5o7TleuaCvWcRtrCJ9AEpPqyNOJfyEprExXS02FXVvUSw
QUQ2toY7vkPLTgpMseJCUGBRQBBK9OaVcvzzjNFl36L/U5rDcplPMtBQvPqFKDGW
0m5pC5MISObvDMRHCEc2z3PZ/5SBt4ZVd1wI/wkr8ZqqeRqWJENF/4FsqWauJUzq
QJHspb2WVrpx6MS5d69rnZBORN4ydtLFXz9QbyeSjd36tLzd+FZW4urd+ncy014f
ARiDYDQEqvd0TDtmCu07HJVI2k/6lJYYom1w3IDRhbK8pmDz27iorgz7rqQygxWn
DLH28DkGj2HyM+iehgkH+W0Zv0YU0gMnk58eOZAqOcLUpGBPSb8mC/rrA5Iqk9We
EjcHLW49uC2HXUlcLxVLlzx/cZdYQEi7vBPjvTSyvZk6N4xMngYFQXOmAgbVoT5j
8k22ZMH2tWA2LApSMmoA+3K08td4OxlsKpPnW8aY15UjvX1ET8AgsXR0C7c2Kr+2
3QbVf6YLiZEJvq2Ka8hkop1yTlZVeLE11qJJywGiMfS1ibiur3QFjVFNpG0JVk5/
t1i8pYjXQu8kjuanw2ey5aK+/qYLNdlRjHN2BxjRIFbskoWJT+uTKjkPjgfgrR36
uMObMMHAuq3E0yrQzDcXaapty0VVZDr0eHtDyPVoFXUrRzZXkYL1ASs6pvmgvIU5
Kr/rInmQK+sedZjnIJu/g1wReYKVSYIpAaq8Q5d21UcPWwRGX/+dByitegK7OOOw
ix13Hq2BZFws89hemSFJOljqwRv0m5baqkSYvOvJgJFnz646L8ed+NRB5Wyn50y0
29T9+i/Zhp+bkcxxbuEpx8yV8MD0gMMRN3dGqq61VmFwda2m2nCVLvTLJtcECeFQ
aMODUvvu61OQKSjbcqT1ntqRBy464vkEMQVqli84cd84XfUSEhMYY9N4P1RoUdCv
2xnPxfSC/9wpjKNRhzwmiUux+zRkh9SPARri95OYRN4tXNLt6SOI/PuRSQbjRSOz
nD8Td3k7iBlcw2QUAtXXUUSKpFkHAd9Olu5AKLdjRnfyo29BNPepLMbH7PRoyM6F
DaarRrBghVf22Bi8rPPom4a49Lh2ERFJlK/BWG+3KsD5tPyKw61vzjcUuWETMvAx
QVUl/FBXoZGl++88Nk3d8n27GmkF/OS0Vrb4Pa7HvUN62oKP9hI2LL0FiKd2t5pi
5aoXrMDdqe98VdET3xn6gkeR0/SH5khe1W4XPLWTNOlCI/B1z9SMdbAjw0UfgP1o
0iPcE3p6cEcq2TQRnCe+1aWpKtNdqF2eh7F0OTESEYLMF/fdsFPDOqhJwzp9sGq2
IoqgTqxkkvPpsGJ0tONvqPxPYrtI9z6oHVHpPES1Vgop6A4GL38F8/nhYkzyD6yt
P4xUOxGrsv0rYBSi+Ggzyuj0LW1OgrhYVCo7vKhftg0B634YbQfFx4skN9M46lOn
2HL4YEBmIWykGk6qQmKVnmAi8gXFV8dDmVX0x/KU1NTR9OY092QyaFvAuKJPVXr/
xpWJ1E4j4tQXu8t7WLCeVuiGmafzfmvOs90KAN0jSMjK5V82PSTjeprXPrX5MY1G
j3OHnXigI2gWouOYYispyQwSnA/UhGyudMQS3xV7RkISPEV+wKRcFaUXfHamat8Z
SB8KvDNs0JwkuQ7aOGPLHpOn9d6e3Yocie6Qpd4zxh48BGFTtPJ01dU1D/s5DPTD
wuImi776dFAhN7hkvOB4FFkvUy46P16WSClEXWiGJdNEuMQlPt2xczivCydAEiFS
QBmA+OgxPZwDD5XJbEmohN3+3YlZwGIzlpmpTueVhEjAum3kq6x46fwyrIjfVtSx
zE9uAk8POIIsUft+7jtidL/gbomOZS/c4KCB/KDOeRzl26UrOLKw+UAujEU9BB7R
CiILXtcs4FLABa0RCAZSvGIA7M9sKbkj9soSZRwf9AcJEgXqGVWenbECMShNmneE
41k8kPwtRgso1ANpB5CF8xj/+ClA4LA/o0zAQFf1/sQE9QA2mEoo90cqRkJjmUgO
bAqTXjH+7aR+N7bA33eNNs1eUrLLBsflx14QmdgH0JkP11o7jKW18RI850bJ/LBg
uNW7gx3jCaKaJDfputpjeoefGHUj4EXDF+f7fUdQcacbd8pj0Ok7xpR+WS7LsUBD
ERt0OhA23BzHwVdT9mNq3Y68EiC8IB8qmwtFkuJcH+h+n3d71cRfu1olhOlt2X6x
f60FQZNrqW3OBkmL88eV+vDQ7B+OHH0XB6P5efn7c4VYqFTXc42yLEMzpQVSxjBl
LhZqSCke5bw2LS5vxcQAOtq8whD08DHJB8DLmQOnMI92ONsaOSdQ1cIDoeCkAaQr
PMTDeyIdwPGK8BB5kivj360o/vFxyOVrTsIEu8wH0A8QPkndN4nPNcQEJEOykSFA
SQ+VDOzMxkqlPVv2dZlv6xTtEL9d2MYe8icFKY7Wp8fo6mqqUe1gwk07oAMUjhe3
bOrP0XTVyDaAv59eaWECOWspZyMvGovFZGP/iSHpzEJzjCJ/jEuQ8cDstxcHM1VA
RQV1ZDUntfC8cz2YbeikB+FRdlCDUlMxCp+OeoVSL/7CWaqqVDfAp9YT9PjjD5bU
kw0JeIfIgvHy8eZVN3mw/ShDC5L6XSBQQcVodjLrHQgoFBgS999PnGayiyke+amY
rXRyeCiy18AQkqyinisGTAjC8sdENyguCtGDiOK7zA7aubWOwM3ywaJ0Su+9jQbm
U79xcuOnkI5k+v2edPwwhIZe/EaUB7optlLg/vOyjHIoPek+gi8z3Q9iX2QX4aRG
7wTtrT+cYzfQS1Ni7Uwbu+6AUPK20ASRZICOMAS78ZbDAAYw1Lfj7KnxxagzA8wA
P/Ik9OfWx0mOrEa5wALhmi6W0Jgl/KfWvavsfejKb4QjAl+Se3r5WmZSj5sJXO4e
STIcrTRa11RC38McpC7QNkssHrWPHZvfgJRFOE0txPbFCRqqf4GeKPMj8SKuuYtl
LC8h6kJYw2WFWAlJ+pRAqL/tPRqcwYpIaoNN73ONOxKJBBQK7ISPOrq/36BTRT2W
CrVXT8MYfDCPE07OPv3Ks5G5c6zhAIuj5aF+H4mUOgu9zB306yOafvfwTrPbQhrs
/wzR9xYzc5jlNd5W/zC36rMBB+6wZjVSgVitq73Vnc5dFyju+yZYg1Uhf0vX61pa
w17149O+bsMOgNTLXg1BoZXMiCoxdPRKWdFb11WFYKtxvcRufIwNmBB5neSMmTvN
TPUjaP3pTc0GSiRyKvqFadrRxYr/u3ECzHvOzv8R8g6UAI1O4kKkaStEuSp32BdY
1XyNQHVkxymC/Y0fjinEQOLFf4aAMQDRo0IHzndOJh8G7fOb1xJEofiienKFQ6ik
dSgGTB550RYhH1NGL9prjJE6vpXxCNp/jV+Anh9Os9cEe+qTOkfTQZqW2t715NtD
eRaoOzEsVPAD94q/trJTfk95KeaJe0UjilsY7XnOn+88WUz1v+JDtFj+FIXHt9M0
6xKxRlrAJs8GeKACDJ+M6ygDBfIM5aMU9yOgacw+J0sf9qbIxOOoqywsJy9rBJG/
NNU40Yl93/FufB/m38ojr03Pp1b0pnitZM5coKsiUyn4zEEur9TbzuJ0bWdN8cxO
Lw1V9QRqaWH/JwBmHHD3+0w+AdOUW2wKMkxz8hqjeIcf9G02hadvjTqR2h7kI4G8
UeaS+Xd7mndDLbUsSoCs6h8nInfpKaxuBo67OypxEfD/AVsFDyK1Kc6M/IdSZYXu
0GjKTXNPt8PCe0JVg6OtxeWxXQl1ma2rCXyX10O6ULSNpuKDxg+ryCHLEqP1BPzl
0xSan4hyKp5gVzgzcmJlnPNnatIpplJfWOJ0JsJF5MxWd+LbFRRtY4t8vMB6xa8N
i/EUW0ygoNiMOBToid9L3ss0Z8I03bndj4ZpojeMLEuDL7RSCLWMcG4ok1YmwjCw
SqJsyWGYdbZbV5aQf38Q30OIgfwi5ZbziAhfDk/64SzoSuqwnOiaph3T6fxTPlb4
5892CKu2b4BFnef8NScTE9XHoTG84ueJBqMi29M2RxZJtR4ns1jEeNITyHbLYHUc
Wf1hN66n/VD4MziRq/g5GXSXo1dkbVJ0tkKSAg1ANtlf7wC56hYpdRH0bftzL91d
glUyliAB777yw1Ibk4oNz9Tr12WJ20uzPZfdcqDgvqJsHAkaNhxWuldUgdbMjQaw
p5dBQWxQ4Y8QJVAVh/It8s22eOepxVN8d5ZhxVk51wehdwTAn5kHPWefxloH5Wi7
+7/45iGun67nYkYR7plROk6CJLD/4is0S5tZFZSEO/bdhTfoLiQ0RyCnT1YAINN2
s1A+7SejM80tnc7Lgtd5jfMsKRY3EeKwZuJUouP56iuUVo/tMFxD13d88H+Vp+gA
/9tPTg+hTpCWPCC2lbd851pdQNx8uG1dN4eneWS9SqvE3uE5v7BkOpyAJTuX6lUC
ZMTmQcXVq03udaCvsZFxKQERK2zoTDCCf+fJOztqVlpFoUDZ9ln6/KX4EVjizg2v
omn6VHxvBiPybrmM2AXlhPHLluwUhKLH3DYZJcAM4Liz6AwS9mueApZcYPAFu3Wc
jQ3Z0vY6fxv8EqF0s0jyFNhnV7eiOi7ZgqE/57PAQBSxT/wF6NjNtCi/vENhfXZb
ALOqYPPJg7PrRNwBLzpeOYHqY1xXCV67ucIC4rV50pl30PeIJuhSNkwiAfpoviIf
/PRAaGG8HEEyuqrwQu8YIDFQwd+sthQiYPJiZgIhyv1yiEaJgID6A0UW3Ent5o1O
wlG6uv3SDyV8abD4W8GZvWPAgHNCDb5FRg0dlsxkB8nLUcPfCGZxee0ohK7hT/7S
9wzKSELgyjod3jrft5cUsiLASkDiCKSH8avLIvG3lNqK5Fhv+jDy/Ze5Nfb4glUE
gwpA4Re1gpaFv1cfZDzbToIa3cQ4PSAB1q2KHhJNiKMjoSMjK+/kk/sTH5lcDX0i
ecGHHrWqsDnVvsJ7HqSU9wT/EpnmSuFXLGRTwOkzQ6VvjAA8igBajYgE3efy3Wbp
hM1e5mkC+YLA8MJtgRtwDvr4dJponr/iEfQUaWD2TeYkqiB+2aKelL1/ppIFguyU
JNIHCXX6+KQZTLPZSURLxb8S8CUZKr81lwod526rfCJCgCPS5CyKZhr5AM1v+uJp
BsWTvdYyrjdYHltNHhI7sxmaJ/LVIX+03aN43p/bA0nvEq77zJYmy3API/Fyz2E0
aEcKNzi8fTVCGdOF2yI/iqDUE5Vfo2U7WBIvTckphDtKctFH83M9JrUFnFW8i7vq
uAeC72Nf1cdpFrenrCb7XiF2k14kKn7dq+i1VvVb08JJhS5bt7EY49gKhry6Vojj
bp2QUYvuRAxKZtCdY26qHE97o9YOnhMOiUf3y/jSbGQAXH+ToYa9DPADwx1t/5+0
Eq59UElsaHokPYlbnGfiNbAI8y49Jnicf3N+97hoVUogWIgFM4wMO5GNM6+viNkb
3QkOcgRhOyI/lYOe+3OlXQwHkQvVrfXsrRqZrkeAaCGA6nd7qD1/KXHnU05ISI7L
KhFp+tV83GLyTOMsaixBjnu+gM4B9OwUVKLnQpLkc1MC9zZA9yY4hUG58WelbbAA
huF+vy0bvJYR5B16x4yykEImSglPrUjJoS6rhFRKQssRPTLwNcb40XKg3hZAQAUt
ke7mHBGzoLGxIWfHSg0ZrEHFDDI7k3xsyelWFvtw5hJmgTGOCBli3qHpZnAryWtE
aIC3xtR/NHd9Ukug7mnZfIqPyLqikCtH+mMaqNBTTc5nodLBXwUkR8kpr01J3fU2
v7cD5TXhwMOkIEvJQuT7WW/6YbvtzRSwqkQfyq9beyG5gSMGiKtd2A0+oQhPQu2P
KJd4ivHHBP1fR1qXtBx0TieJs/SfQZhvYp0Hlc70ZlbLySY36lc/yLvk5Z7TJjOP
ikP0IsqsmhpeB0xhPVm0w+VoF2g5xvtQq0cbipLBArznq9LyTUcvP7P+wAuRXl1F
OyMl9kzl20wufiIhlH7bMs2OdTt6TUr94S233P1OF0tBtWjN39WrpYDPlTNJKwvF
J+1Cakkaw1GxtBge4w8QaE3H8p5CHWvbHTqQjFJBDCPCPy8QcCD81XD4Hr7Wojyo
z559tYNIzuqD3yVQuEXF1jvjVdYGoY/oDV4l/hYLpnQOKp/MZrS6iPwgCPQvzc7+
rv+BAypWObpOw9ogJfCP2p168BPk5mmReRajOnbfnbDvKw96AvEtLuFc4MzOXnlt
DLZLMOLn//6RlpI6+SHGXc3ANtpEMphujSGZ3Jd4oBVUcZ1sPDySr6grh8wHgK83
Ju6ruIZyKH7yviOoyIIHg4oX0t6Zkxp3piTFpt+oNqeQLaKB+GOtdquI3DGJm65Y
zeHRqOmsnm0kUv3UHuJfWY3xbC+S5yrGN5SGFl3Veno+UQwnHn6X6ZU6FUvk30y8
HjIV6+3XagSSXJZEeXolvGACc5W0tQCCzTKUSLA1a9Cy7h9CQe9uN6jmMSdvpRCC
pFT6A5KCHV2opUOKipchQOR4Bndd4nuU7MHizkIS1ycoVSjyPhpcU+hWy1tkY/Gs
YSCIEomCIKdLIpvfDIy1CXLqApBkrTRmoNZ4ZorEEn31lM2ec72HTAHMLO287p3C
JViXF6bC6eDpabB0OY95BvUcQBCBoXpyscwvZb/dRhFKXuaACfLTDjutp+sZqNMH
aedYj9ZpWz1bXB9oca+4tnnzVHSQ+R9s1a9u0MKD4BdFedvy4676rWW9gvC/vCxr
kPs+VNoENyycyfMz6v4JIxQjizE0WVowAjIJp5hI8DKdCi/C8ciXVWjAlmXGWhRH
1ZtyFQXHVKHv+jFeHEhO2oZhfLAIi4xOAyphvO0C5PxyD6ByNyyzneMij8pBxLi4
MZ2f88UEfk+QcaIS/AzUhxrfTeYsoGTDStI8siSPuCoMSqVCZeGRJ0CQ/OyUGP8B
4HN+d53RR9h4Yv4cruylA3BLIMIRsYJwxsfNXXb/blouQCjjSrLRDOdNYQLg4EnH
J+eR0BuYgqEDIQfBTyWfljAfLixlTao7JKpWtlz8r0figjIRvWFxQ1A4n68cva+F
ueD/Je8Q1mbSoHdwNH2BoatcMj6C0Ch1Bp67+75PKeSQcaJy2U3cGej8l7T1oBSI
zYCaefrgBaU9UtRVmbfzLjqycJBOpaV6gBzodnQ2Ixf+9sjwSthfMveV162F93Oi
89Jym4cxKlOA//dHPUdovukGfpRzlzBk8xHNh1v08fewc2V17ktjm+aeEK69vMOR
ObiIdDxzJomjQE7ZFxWkb+pdpto5MJxdTOQjQEh1V/dVbCchKOLMCzRu15mmnldc
l+nSoqXVMjauWfPopWuRvSXPnOOnIvSkQhQl23XsEG/WNRVFUOuqsOzngpBwd+JT
9BJrMMxYOEk0mpV0B3lsvtTBpqXFdnd2BIjHLTR1dQHw2XkREIHCOseB6Mjn6tc5
QiY2bkMNoIstqm2UTuTNPqeB7aPyX2DbLCrbSdhVHgRmrJ2vh2mLPOnNHFmW+pFW
EJrqi9yuU1tMTs5gZL5ppkwn2dIUbloJwAJRfCgDEw1Bqeza4G6MkHi7zscpJdzZ
Ge0o2UUIeDXu1sWxb5lt6LlQeGVJjDPJ1qNYpESG717bBZx7tlIGR863J8QLR0/c
wnD0lmGho3E+25NQK69fNFd1C3A0KWlhntzLHvofBm62M/XRv/geGyZjGoRtodH0
lvIPAyIX61rHSpxNiMxEz02BA2BIKqdRaQAM6uUIONLYa0RIAKrkPB/WMc1+DLrj
xvk/xLJBiByd7AZQRYO3B93LukmNv31ig8w5mUBCjPFbakMNhp2AEw0/chYRvp2i
PeYHsQkD1U+h+yrnkXvKrLxi4s82XWdCXgsQrGPdGiIE1CaYYKMIxH4Wep2cIkwe
oh0Y3733OUyhWJHLpxdnbdVhbfI/uvpLh1ZfJMQaP08FVydtHBVCyBMn0722dJUt
n531WQm31F9xmcdcDuqzfYweW8kQuOY96BO3Y25pw5wmdxucrqrbuiQ5KcKnedVZ
fCiIPr0XhTUFDS+G71wpPquSWZe3Cov72/umIaReALliVpV/xYP1jhtMiVDmxkmg
YVqnKKdrfTSfsHZV2JfDiK1N5k3W9F2HUK7ts+aw6PyqHx4G6eNN6hFxzDTFJU74
pVSepmXPkXbkq018q/00PvXKpnv4kAxAixXIDsr15NvV6OqkZNwNv8mhlTavsJe8
70glWd/Cpri9C4lzBggRPTiyOHxHpW7k1Cp10wvehYrnVVP3EjtRYhANvXtwzgHC
a11tnECTk1a/UPBv3o2z/22/Y9QqXvnhQD8i64XmF/k5PlKG549Z8/VzCdjw5ylS
PKIVfhEQCSmxT7fiqVgTqFAtRdaivBPi9xkikbQkWAikY4erTCdtDmvXPi68MLDe
H374iiDhYlwVq3+3+760lVdExppLOISAamXVf0mectJowR04lpWcnyLcdofMjFDA
4RNjS1hRIORhvnhuSpa/A/9Nw1W37fxLnSWQAjs97ct8yyb+bD5WYIeWF+9vhHta
YM60o70Jk4BV/0K10/ImzcsutMhnZ1eOGoJhP8CXFrmmCu4MnYV7I2++0NEuCqZA
LsHH839OErIe/jmhbfxNjw3aGPf8AEbjACKIr3lBu8gc4tJjEhIiD+Jf7o26rauN
ENHCyZFqLJJG+RMtzKUtsAqIxsvroh8zvN7Mg4jbhOn4YoVRkZzwpmrAdI4p6VnV
xzbW4F3cotby00yEUv6fqyh/rx0bEMdTdNrASWnFhxYJQDcYuWFPYLMTKJaM/6yd
hD8HDv+rKCbxnCxIFMJ0zkTJ8CQVB2wRArfUKfLf/lr1ZRwMpynZwKiDYQQGVPMe
Na4x11guFyqKod7Xun2/tZjfn+O1xKmpgliyD3iWRH2PlbmD6EZbY7qupnrVey6k
2kuwHYWz59q5pMYlyNAOYfXpKQ0nnn2lh+9P4XijQL6hrcIlFgzz701lXHUXqhyj
X70tdRi9RZwZdhJVko+KbtbSTIoPpF8OGroxKDSYhu4o9TikGskDpr0jhlQLxcb0
/Xljrq9Wssi7ZZKXUYssc5S/+gCu5Eu08O3J2VscCDQm5UTfAlMtFWdkbSLEg4mk
AmPeXvLOM6zuwxo+Z5lOi+SUQFR7Kk5FQVM2b0ezp5VOo109ggDOwe/zgBP/H8ky
nZf6LJoxXXaWOUklU2GFifzDAOF2ONJKl6kUuGMYCT8TzcT6Kw1zvxgGMyQ4rM8R
Ddz7oxm0kEn8/LcCDeLspXCbNoXEpWvhRji4jXzIBJkEhC5X/n53RxdubMWa4FlM
+evvEFWvdEiWkrOFf5mF+MCh+W7SIj2DVDWwS71Ko67Rr4UugRmS3uG8aKhiBWWK
8M8evmAq0y90mkZVfrPOp87uEcq0jsjtVTREcu7ZHXrSDhmzbCr8wtP8DrYoulvE
wMvR/rq4nphYoTR9Lx4kPkYJA9Pj74lQo64SQonh6as/hlTCUTlVnGJRsnn8WHeT
gms2/NwRjaaT3Xs6VHi6W9QRuBNybYnYuOj6m8bJuh44raRONTJGlv9q997KDynr
nMjIyM7yWRrODu8pxB3Bhxs3/kjjy5isnICRJQdUoRICd5stBWPQ9/KN4/71L+8W
7oD7ZKpOGodXtqcRpkjnZFOr2szGVKQ0wyoh7umro345xyHGS2bKzE2F0y75FRYH
`protect END_PROTECTED
