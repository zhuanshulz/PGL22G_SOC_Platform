`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pyTFcwyTqA2TW7d6lzAL5FjWXrN9AD3tnlFv+JsvBq84SEuc+9qF+TEAPs0BV4UF
5yH91PoGmEdZRj1rGpUxDoHxrpl41z5nZwMcdHvwcKCUrCMF3n2Sm7gvpgzQ+IC0
JhOZt2F++hcV7HkCYLt9mXbpJ+480C5ZIAE5kf1fxt1/z62tkOSi9FYBwXsMEVee
SOJrhVFa+xqDasl8ZT4ozRA3QAsG94MH8oCOJtaAZsPGeKNyIoUg4uYPdzDXahrv
DcE6WJeGRavFUjAVKSpwjMhh9MaDn+p5AIjqhAtLRHMx8/1S9y/0x5mEKSKZYPus
qIjMmHisgtDouYitBc7y/cJrM4bKKd5L9+V1Ru3NKu/5mijRFuVYwmw/7V5yn27/
1NE0Od/4u+gucJA8iOLlSg==
`protect END_PROTECTED
