`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9dWjIiZ1y6sxwC+rwPjfStAB5rc4NOaEsZoHrNsBcifDUu8H80S8TAwNKNpe5G3V
TR7oXGV6AREMApQuZ1l/LQjLPpWA/jdRkqgMhPdEGUSXXUkaIHg/S6gJTVp6pvYU
oTFNMVG6kbw8HWp/Uq0tr/a68tahuJCYKbA8lqDBdh3oAYIQxx2WacXBG4KUa1zv
/4jYs7fdpGAU/M670VdYjHSKfjf2IBns3YikTQjjcIK3IAH+d9tT38gO9XPg2BH/
AlkoENo1jdMNbe8IOUCHxRQu+l3JruMX0dI88uyExKuwPExQos9Mh6x9nVICxg7m
sjC98UvD/XQ8DCab9GOY6JOUlS96WFOdpwHpnj/QgyWlC8mU5174tJ89FmzQmTzF
tKedby6g1Jwo2AljEApOSDFaJ+IXi9bQ27FkscygbmfJPMViXPOWmVyMONTXa3Z4
`protect END_PROTECTED
