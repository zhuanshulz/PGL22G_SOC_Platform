`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JBYp3rjQV55+NY1b1NjVxQv8OgNysUYbCwWJ5O0CWB/WNuxNA0zTwaEt5Mwt6g3K
gy7N8ujZHdW5M3EV2kS27+uqz5M1D4s2knnvY1mC22fAYJyPJ6sAxANPIDJC7hgg
akODfl82TZ6+il9d5CKO6lJlDQzoW0ekFexC26CFQUW8HyOuGeBt253oXM+Zcq7D
jDEFC4SnzUvZprko9kIIZ+AC0Kwy+6gQOTBUZgO256ExiIq0SEoJKKU+ax/z7XKD
LmsDP0Uw9T026c1sqaBVs7ItkHGZ5i7weMSEnYUDMU5Bvt0n5MHHURzPp45F10Qs
Lje0/zU+arsqy6WP3W1ncuw9ltl6pmxmDIcYH1njM3yYPEM7Fr2TVl3vaqtS+z/f
35uHuuXv6MFZn62MPfoji17XjMAIQgEOiG361X0G4dBGwkY3pKec8UHknW+SGzc2
ksjB86/jhXtZPFXARAygWnjB2VFd9pPnb77F9EMRdKH6mnnraQo3iJ4Z3CL+4C05
ui970yW0lWerDMiw11FnYlIeaGTw/fsGgXsnr/ryVUsJugzg4athYyrkAclR8Ux3
0iN1otzXyy0XEfDQCVSC2/dvLYHB1jGtI582e0i4ROJArt9LKNfGnSG3pMj2StEd
bDeWBMBmNlVpUxp2o3JEN0p5SYTdbqS8EQwErpHXgcGYLcWWIvdG7++4KdL3RGcG
6RRw8cxW2nVIcZTlKm0mfhWr89efVYCdcMkNudSkbJZ6uoUxZ3kit6n3c6Fqmwf3
ot3mTpJzX83CIYVlknVoxu4WTFHimbh6/fBED1bSvSzs2env8S1slL7X5R2PaNBA
zUTJBUq+kJs6NfIuocTMleVmADISir33fKiI/oNBABZargS1kV4cHHrBhRC6Zofe
UlWm5nG9djvbgueHJvH19mCSyewZQ/KURRnKQ6C/s/ZyrEaQFY0WxaJ92gPbd9Hh
3bPJsvRq67UN7+yJIY+Rc8MLYb3RdbsXhJa9jnUSqAbd682czFOoBwSJ64R1zIy7
ejGfhuI02d2avdiVfkGyeDD96NNTyRx/+qHVWpYtap4t0nW0XCklyW1KZWgp5ZUk
uibBE/+gSnV37T1Cj7EKDLddDtyM1lk7R0SXVE5q/2YdBFl7hOIZbDKgPIqdzXVc
72FHGmrfINweuV9ZpwY95pDTKja6FK5nmPqwgDRL3ytZFa08LBVNGKT/FFYzpcKs
kHOL1oUsvTre0mQx8hU7wyI4vczn0+aBBbm9qCmNNs46PkDtzchSesa5KxohI+N4
HkjcsVqRh6xHtuVAKVWTQqCelVdPu6EyoUtdu0yEb6kgezeoa168+VWMh+Ci7IcX
IOnmPwuS0is7s3XrOddvoQ==
`protect END_PROTECTED
