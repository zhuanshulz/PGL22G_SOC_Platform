`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1CNz+9d0a985BGwHMpmuvUpgAsDhhmI9S7lDwIgG1YinF5c0I87sc5G2+1mQqfIJ
/QYhzcgadAM8JrnUDWBbLYmPDJgrXbamVrv+UhTISb6jeQK5bJvoc3NZEN+okXh+
axR0oqcrDmomYYlXl10KrGXVHOvYEpQcEqoUnIxDoaeha3NoCxw1gn9S9megkKYp
/Iawf14Ksvzc/7BjSbFfvXMhkKe/pMhLOztpQYxd0ACLpvZoJJjykEW5+s7eh/In
vxeiZAtCB8lLni5jzg15lz+PVCxiuxv/rLckBt8e9hVDMU8x6Y7EU1QRs34cURH7
qc510So/zgipJo+424IO69f66kHVyK9akKQWI1vGmjpRi/b/6Hmtapoy8Xvqt8n0
/NNLoGOYUj1IvYjpVc5vSLsfxdSsKsslo+U5g1S/qf4CCOV0DIJ9yUKONMIUMNTc
6TqGmu/iJGizzcHyXDxv+9ET6Z6FWIJpQJHKoiuFA6w=
`protect END_PROTECTED
