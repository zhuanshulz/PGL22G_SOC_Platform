`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8TZNdr4pylUgQvGOql+MpPyfkVI5GEEMs906czGlDFsn1levvN3au3efeTwrRaV
88kXOr+jItNjx+ZvWcAwsi64HvXG7IA0VyjghEXMGJT7ZptQKBCjARcErrhar7pm
owhj7UU889B6VaM2J1xi3EPYOYKX7834ml7KLIp2NtFn31LmCU5OH1oJ9gkoyZM/
uck7Ss0Ih8yL/9qDlompU2GwVr4gstQjH0YpjIrzev5fsthmIM3YtwaqLFKJIZxj
n60iBT9kHp0KKuTezyHGEuV+zHICinm9kyk1rzqm6DhZflzvR6V3hJ6nWDREma1p
D+1EUiCQL/RKdJ1ElQW6M/FQCihSE4neubnrThz0ytYLrzfsh1Ht8dnXYMr7eAVK
11Eux9R8nyhdZHvqszbWwsmZBErIVqr//iMzkVdGMZyZJOnxJ0raYqU5HI7TLDpI
p0X+U+wubDGi7otS6adQRkr1XrOZui9GkUU5enF4n2e4ldLIa0UuVNv9Ke9OzK0H
eGtEmJFsokb0/3YdkgzJQdN7AJ7vIDU/csCfHmbGZz6ZitTYmz/7HGlUSrgwmbNX
ODxumN6Izy2qfyIC5v/4nw==
`protect END_PROTECTED
