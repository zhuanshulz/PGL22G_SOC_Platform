`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QU8gTJpFgvtWQbTB4Z3KaaOhmX+HG6GdRVWlK3lnZYOmmM6r1+ce4lZ9DoFuYZFl
g6aNAGLD0Jm/6BFyxwOatgcmmmcQ45fyWVRkl+wcu7b63+T+u9y7fUy52bS+A/94
kb+OpJdhtWq3mJr+rzu8dgjU0NV5D1A+Ly858s4WDngkbD9lPA7BSyDd6kWvPvyF
2NXrCx4dkBn2Nov9zdAVCfoqIzqK9PbuXPvtpcA85vXEnfYvo8+iIRZZA5/glvP6
yyy5B/7hUv9fcW87x1jImSeZit++aifn2w/0LnHoRdAkaPgNvH/dqEFCoSZmggcJ
0VTe8ILcq6d4AxJU+xV4Uw==
`protect END_PROTECTED
