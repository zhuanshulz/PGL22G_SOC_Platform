`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lth+WMRvwqqNtFRosm/ruOYzV09HXz2P8s7IolTiTLog1w6we/O2LJTEg0mLKGVt
MeFyQhjjT4QYSsqEG5MRwDK1DwOlVmlsppwdSr1+iHa/8yWxwdrq1QAVT7tAQCne
wlkn6f2DjsG25+NGX5x05fAzZQZV8COQngkHMITiGkplI0mK9BoJ4BIpZRhWKukN
5WR16OXAvK0MgAbkpWThRjblFkIXi3pKFtpeSnZx7UMqzHs8pAjgK3ANJcb+HSV4
Gd7Z+MhAfzbNaBVPGAsNfCh54uVHz4F9IVnSr071jZzjUcd5hdoAp9shSlVe52i5
uV9PJBtSk00oaRwHWaMvZLsWZmYxqx6b34Q5EiuAy1fpXcYtectr3QU3vBD4N4QI
cZ2lUOUWJUZ+/7xehH0MdQEH8wr0uYw76zxkeFz5XxR/DXyuGr6b9d37Yg7VOa7j
TF4wtY9XU9irDUz99ZGlee2PIdakRpselvAkwq6X/C+gf5hY2qqwHDisRfAF/mIT
x1/7BR8rKBi0zsbH438+EgMs51Trztp0ClOW8dUyhrcmUZyKAWOUt2iJ3ygYAWWS
OhKibyMhIBhhKMvppeDH5QtEs9Pbdls9eXKicqf4uCXgYqsHhvVGm/MH/bV0NFVF
J0IjSIDELdGx3yCbjijSq34/V8hx+42gUE6LBkjKOYZnCtH2Q0IKEDbTm7wGScPO
8JR3H+dG94GDQUytIX+CouLe1UGuBA2gTxx+I40LqOHJg848vka/MwxIW8eeei3o
BbPZqS6gHmi7bCoeET+S0xQYc476hzftmmCnyJspJtm4vw4QeLw/G8oyXSP6bv6U
D6mhFwIHYkYaDnw7Inws5aC38J8T/vdXC+CkuhNj7EVhi7Rf45u5Fd+jkhsf05si
AChtHXptCYO+37OAA+5zjnvZko82BTif5BRC9BnEyDpYJ3NQa/Jla0JNYJ03o0Vu
vg+bYZ7XmPZ/i/MqXLkKRtE4v5nLprSUlzwn/t0k+At0fPqrMiKdPDOgqKAGVgRF
MO2N/hLUeGT+p+OaDpUnsVLtntg7cHq3sBkq4agoIK4qQnxkUyK5S1i0j5WQ8YNC
XwzfVLOkRhtGk/WGG9DCVpvvqOxg3HCcOjPqRyrXRCqcmkb4gTU8cbfACF65/7Cg
nxU+M2XVxM+4HRVfXsO+iO0iByTKfH6GUAJHt7YpvYdfwcXQz3tWiR5+h/VUjTnx
XPs6mn7Rx8w7sTHwJhOXoQ4cDJb9AIpUx4PmdpVHDBiXuL71uQCFl+AclqVHZ3CT
7m1YQpD3X9NkL6AvVRSs2mVmFiMFYqetCaUxh8c77Hw3dK207fjhd+oP7t/srlqP
137HOnETyiG9p6bROa5jPAEHYnTi4prIRdZkU3pYT0aVyd+IalURTnP6/x9ww34p
/Ts7PiEI1NGL+Ynq70I78gwssiC/Q8LMEbX+RHJO2tvMXf5+CAkn+MfzJmjrpCoh
O4+33KJxxSG6foKhjzkYjFMcHCu3f9z57YSYFCsIChi3PYK30nWN8wvblg/A7C4n
25rjbSWco1k3xkqD+hTwZXGCF94nrdw+hnUMUknSuYHOgMqlDIXOk/XtVyYvaAPl
udNyortGR+XmRKD1ItH2s5PD5R+O62fgPLTtvnrhVOhvg24c8f1UzEgoENspOgpf
MkZRBmdMbigVjmoL2iMq+7kWBqMQfZXJ7qmlxzaJ5UHHlAOHTalsgtvnxpwZJ614
piVAjgGHiZ9MKt/RQFih8MmJGWPio4mq+yAlt56vxP2N1MUnZiFlhrfIJAsq6Q8P
uRcRW2f+D2yMJj/6M2A6oJmiOf/BeHNV/BeOeD++SmoHAcoQ2DeeD0Fo4X//iRHS
eT9WG0FT/Uui2DAl9s2hvWChp1rjZx4RwcG5Xx5ifAI7jXN0sjD8WWOzCpmHKNhH
StqHHYw/QY73XBQsS6rsLvRGHTRwe/XDrlwvwDYFcS9eXbEk8WAwDrSZvUlRNXwr
qPCbr9/dr0CBf/Nqzy/4kDIg0nkFuGz1elUp03vRvdH7wGPr6+lFd0ogT9Q2koj5
EcaNVLZTfamlwlDzEXu3RQPoBBXuoB2QIDZ192Mzz89rTfU5zKWu+T1NoLsdF06A
2dRxirn5wtlrSGg3yz6rA2dk55gS7RV9PqvQCWTpsQlLNKCkSgw98ZJNrzOdzGDh
QC1Fl3XYGm1l4WAGSsdboo3+y3tqPORL40znmpF9rC9O5Mo8+DDKHYo4DsA1poVL
qo8fAGUCYQjWuuhGW1O88h+rjpxpYjndNiQJSZ2VBiEDGHrZkYW2TaB/caY/BkcH
30hH0AeguY7JWuIOrsR+XxEs6GcLaB/oK87uzxZRkOVS2bjzCGDj7vpSjTWoTLuR
gihOGpCTDS1VVogrIpbIkDMVzdtg66SzdbHTQPy1kpHwZ0RRMGMMQq9bYWvysQKZ
dCXOidLr4XTCbH8EQp8S+VhTqiCVg+57LWqzvER4fWCEhIrg1LEIGa5naKID2P8B
HCONH4ko6nUgiu2yXD7sedmMoDSt6QVtRWPgaBm27Ar6w5/57VINTA1Fy8XpU83u
0sEmQBYTjxztXka75vR8rBnMbV+7cqfSSRXu+W45CnESDCadHc/2iVTcI1KseeZH
qojtk9vBKnAbtvVRaSQJYs2HusmKuuOucF43OD0QtL2cdLyECgjuo2XmFPWfJfBk
J/07Qz5jujyId+NULNhELPBSd+LXL3VgM213WiDom06LjVWxUooKSYRl3SGiBGIS
QUgTIaW+Su2ut3A09UeJqRAnRUt9S0XeIywqJPTh0hH5VRXSwZ4Q3daK3xzTNa0y
AZeS+iTTme9rZdqQIMvhkF+r2sful9vA+5ljS26RqX6JgvTrNVHttTsbLPlGS8Jv
P+8nylrcyFReMa6BRknu7r9kBB/PeKJ64PfG9El1dEZ3k18OonMtvBtf0S3wNOEG
2LDOnW5gheJAB2KD91CA07ule7UGobnGzu/Bbn/YD9nARd3UoboicxGNSJ4fWqlF
R3xExOUQ/u9qt5CuT6tkSUxnud14XURaJ7ABYU5WLwFzlDQ9Jb9l2dCUZbnUWjam
9mRy+MixZbdEPNcJWJWhQUCTpciItXLXbr2C39krpsbmp0AlqOy32Cbm3JGjm53o
m+ru28HUGv3J51Bms2se37t9RzvQtVQFrmvvu7G3Su0/u2UED2EdXqoUub6cJjY+
Hh8cZSahu7B9iMOhCTQ+Dd4yVO2qtYHXL3po9eUnlFBSLckQ7++fOp+W7WqifV4I
of0a5BN00qpgI4rpFmlFyqvTLL9b2gQfWViYXWYn2Vs0RCwUmo8TWovqsignBeI3
Co+WI6ML5LmuUUSh2qVXkqMJG2K1IZ6LqePYAuaHFEAaCM5iaCH8L1SWniXQ3xcs
vIYKH43fr7NgUhOmkaHthvle4uHfqcFKAYlrwwHCfeoDk5PoyuZOp2RnBI+ZiV+D
AZNuUFIfL+Cpep9IX5bqq0wKdsUfnWe4tkuq98OHs7mMXd2UQ2HyRieLhVy7h7Wr
wfz5/wwuzcE8dHVuWH6zjCuzMr0YnGoi9vmM4WlmMTR/Q2HNc3xhTQXCwsuQtqP5
Ip4xUro+CyFnX6/2Tz2ST3rAtDNm9joAEwo0SZ18K9Sqzlqet7iYdDpn/qxJR/NO
gmPRPVf2tloGGmTkb41E8ny0U31FRaVw/acRYXeJZLpx0ITBXj6ZV/k2BlgVCyJ8
Cci6CdWZI6qtdR8Eu+71iPnGApUS8lOUVj1pExViCEgo4SyvqO7yxl313e2fvgfG
sJQcHhJyzkC2PmXwvkyNwwSHYmRlW4ZPdoTUq3GvPZf2muykPmxnAzwIEGBbZGas
8x/FthN/E4d12UtmI1VgXk0mHyP3WBih6NQsy59ZkW4XOgsQTMcamrYc7/ez+Rvq
QBwe4KKnWhHShDe3sL5Sew==
`protect END_PROTECTED
