`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gj4b4JJfOLMQy+J2lZBPGmOMyCFAQrUUDpnfTuA11MuVppm/J7EPrbZMquPrBfjY
qBWNeday+NO1enHEsqE7CFf3M3PQIrITx+48P1keumzPEk5eLKMP6H4Tqa6LuVuK
d7g4bhiFG7L+FxlmN/pSqIJA1wdIuYcGt9Ll0KmODNmVdIo2z5YPS6zhFBC55Fu4
KIbKe3FZOU1wT9CXDDcTbV4Xt0F6GegqrwXEmvnZ+LOp/JXdLePzBiJXICjiy9FE
+dEsagFwUj5DRpVBlHSAXjMti1cSmRqQIAXPHoD92ZwzZUFFVpatgMExeMitZR4e
eekPjhnJasth3yOXrfGfLqY1MnOSYqpS51FbP5rkJjeuNZeqJLETgEf//ICrQ3Pz
+c1V4032XwD6gPMZ0X75S7Xu15cNdEW+vVnIbOL8YrYb8CvdYGfN/19DCKj2EH8T
0vFGgbk4DwbOslZrwTBZbTB1XFLoO5N9uM7JEmO+vxil2TccJgkVoeHP2eHBw04R
wvi9DyToN4sDt9LMboAPz9hI7iqB3Upr5QfvknppFHKdvPyXcicwjUbuPWJnjHN9
VHt9gPQNi9d3FyDOh6Oi4I0CbSFFnSmrhapSNoD3F42uwSmgOi7C0XIpRQy+x4N+
Zwq3t+bI6ItejxYITmF9yXKhvUGrIvcX7h189qz7Wljsd0xcHfz/Ydro1L7oUqZ1
BefKBOWUN4PF0b7ZRAXb0JGCOSthW2yid6hR+8V+3iZEFL4bLoaRB4xJyaW/qkAr
QeNN4fJfF7cql/WzhVR/9HtIXXUGTHT82GjWTD/W054=
`protect END_PROTECTED
