`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bu+FY7KEye0g/ePelkcO26GkAU0tNhVyb6zk8ncdZ84GY5iClkhGbntyFSR5mpE6
jUEAMi/LErZLBXBe/6Lh333+vUp5XFQQEt+dHWBRm7tSRt0Pr/f9for9QOg7KO8d
bG73JEWSbSaGeFIB6HNGeK5wNhCc2zk72T2t71p2aYWewEfViSNz/VKqbGZvWrHL
7j6Lzlx8AmwJPYYmbNQfFjjNGHBMYZCOfbMmOzuBssdjm+8tLvP84dc2UH0TCsLV
8cgbwyak/48mt/mDyvdxJtfviB9ck0bEIdUSbOpzrMucUC50vZwr98ehZf5o+qLK
XlPrunM+/dOyuDgwFC973Br8aQ0tBgVzHV9UAL4Kw7bNChafT7szCjwkxlx2VDE9
N+Oir4ixyNNpUqd49RLijMozraaCRd230pf/C6wrHFZ9gEKCMW4zcnKPEAW1+N85
T4nZDmasblPbumfSRXUTGK0jSdPt/yIoOadWGRkpBbckMYtNSfjnqC5Y3HF7AjGa
HrncNohr4147BCjFSElLc+xFeAQaQwJJSrIRwY3oKCV+036sNHtliG7YPbBGbESp
G7mhQVXbGmTW/Lo5mHX/qKV9xFce2d5h92JQrcpw+Dk6o+UJYos+fkkaa71YMnoC
`protect END_PROTECTED
