`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zZUxSXy63CcNTNI+hkQLpUJ7Uriitjpr7010FQwR2kthMRNqZCt3LDFh7nuT5DXJ
IQCPfvGaLc8Y44epuV1BkXgJzFg/KcZ+rlGCPWsPbiSIlRrXd/h+tQGaT9/UFWQW
DhaApIP0dzewAVLGUvt/JJsYWhT+k7kp7fFl541110NTxX+GGYaSy95BIUoem2y2
nwglBjzHgI0g/UnijkFLWDuydYVL8K+bcROMvdQtxBYfB0fesd/tdSiAlmuI3eaR
VUU2PnSzWfZ6LfzadHf70lLgrkZBkv0hwOoA3kxYUMFNLzUTZPZiRktkWazGgzui
4dOQ/7Kxv5ayzBNZYFrfHglU5/1xA7kR0FgDMCYOZtwCacP20Tm/d1q15nFq/5Zu
Wa+weWPD7qs0/14Q4dEtz09SAqgHNqp009C+GuKfq9UmFkG75xUhp/kcipEifYsH
IROJcBXbmHPTcoK98buWsGVgYasNgWQpE/k1ue/qz0XOjSpEtJdAfoTvCW4DSRYy
mc6MUEJhDFJo7VKvTaaFhbstTkbY59u0it3OXyBj5XU8CY1FhwUpfvqlRUSsJMGW
R99L35S/l++BgNLwPT1hguP4YAYA+MG5F5ExiTyock7v5HGdpDuaY1aLsxQLjyVz
dENN1TeablNtAIuumYYuNFk4Y9Lv8ZNz8KlzbQwkr+KIVVzYv+QjAZ5dJ+W4hM3Q
fwCRPyyyF1Z0Cbeh/5oEirIxbuMSe9RpjAatgwlRa6g2B7HlnaSS/ElWvTEHb6o6
Qm1OCn17LQF7qfWU0iKK39kujtrfA/bfv4WfymgQ+nJ2Lo34jk9/P5L9sqeDvwfd
6K0m1q6YKW95+MLlZwzU7+a9SPW/BH739O7cOW0pm+PQVoqNxcgZ50W8V8VsK64/
OsaSp0H0Ev73nxcCV+trlHb3C8AMJ93h/W6CI8nQ06sUKXmQpdbV5PQnhGV+hs1K
n8usdVC4vvHrD0g1w3YowkgTXHu8RLE16ApOy5XOcQ+ChYGDaSgGxWZxmIq9MfCJ
qJlAn7UxRu9Ief1I4ItjlRg1/2XseA6GAw/4ajRShJFFGjl/Z0bkOeTZtHOmzK+q
JIUh2Q31XWDOyRahm/uMW8U2pqGonHhSEbnb0dsukKpL/u8HCuigBpWLYvbbIi5p
ltVTXIneyfeBLGJLOb2kf7HFYlulyMNk7XwRjY/xhtfoch9eyppnege2ltGnpaXR
c0kraDAdYnaCPfQjxAHRUpp4ppaczO0I1JZWr68qjWZ1vGTn2Lu02tojdV01UOJJ
IoO7jcrt0gINzvnxJgX4dw==
`protect END_PROTECTED
