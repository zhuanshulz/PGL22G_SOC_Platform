`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T33HZdXrqQGPnh0PjlNU4i/NCmFdePkQ8w0OTWPa9aKPUSgWBiNVMoboUTJsFdkX
ItNy2lNgYztQWPnJ7kEt5tgy0MecXGVTzVnuLzzcA0FHD9LZFkZ6S2Cn5e0sxhKm
DO1RaqE8GJFD4wPqQuSb1pu+WP7QyipykF/2lalipFyhc9qEKR0x+X3zCMMr0/k3
aym1blT535lymIHXzOfTIBPuwC1FGUjzEEeANcHpYqM3WRDwA9zJtHx4VrOYsIvc
kddsK7tCwv1f5WVLWcFFBJksD/f7BUg13V+J64utsp/lr83sjS33OdRB4g8W69ym
P2lvodvp+QGGoYG73Z5Eq6YV1I301cfU3ThJn03vywPoolTvTofwIWQJiT62HURL
omHeS2ABr93lCs4SYLZtLJHC6Y9KtVnN/3FpVYscvFfuKhto7qYm2lj+NuNn2Za9
FBudql+vebcFJlC4CBIbbhT55cpugwNbw4d/eMnZgf15+0T5Fau1tCeMgZPvbZ3N
4P/NIy9D+UqnlgLpxEzHQ6/NMBcuqh8T/TGj0uyZtCDVJajhc0QrVpBW/FhI+4EB
ZLYweI6hN3U7AYOZQdQklnPKt0BRdKO2GkASEgu4u2c1u99NNxXvIYO66ZdNdia5
bYQlfjmnD8m6eoekV1NqaXTKEMHAizFWh0fcLgHnW2Gr7SnN8CcKnwhm1RLF1SCI
ThLAiOId+1nyQbMRc86/vWk3RpRn8yAy5F1j2XslkUD4mxXmK5WTxXlBMiyz4eQg
YQWiYSKVxUdfuzfjlyyduG9NPegohw2vZjP5rEAVtBBQbPmtkGE93j4I0xeMI1lh
BBIwqs1jYTm3mIT+all1WPB/kIqN7mlym2NHpCm72EXkBIqiG95QFjkVX6jwpsrX
APwrTwcAIDG61BRN5gdmdq9EQVMhIlLlB+nbbi6I/Oe3Vu1mzE2vaYr57dREQPFE
Cu3e2hOnS+JRshHYmggQntfWTiFrpoSEe7iFs/Y5tOdYK6zf2AyuYusg/84ExKPs
0c/E/RP1XP333oP8F6hQ4GBdnw+Jmyp2IXoIL2mUVMPgwsqh66AD6qdEpF9tCVYz
ohs3FqaH/kgPI1vVqkKpC85pjrTWjjYpY9MHw11NV/oLUagVD/l0DYDeGkk00G48
qgeqZe/y8CeI4F9qxHN/BRP7NL5XNgHWAdpZpaSCslRSYIHhRhF6WL762e8MEY3m
isFuaUy+4j7b9k3fc2xXUvi+01cykwu10EDAZdZijM+ULJfqLtqwH3viBG37XmgX
NvuZVpqKJkxTdNMRX21Bf7TtXIhd7WhqNWssM+kiESVwG507mz+Lu9bcRdw2xMYU
zoT3SSvMD2UvAqhMv70HrXJHhvEZ9BX9pr1B6j2g9h17gIdJoKG5473R7/t63IBZ
2JXSiUDmqFtRNQ8BWPbbUSyQwb+wYGaMsVd3mrk2DtJ45AMJWX2f+QgkAS6T/pv7
zXmdh3aoGkDNWShJYePLcEb5vRtCLaAcXQHRK6gkNHTMcKZ4ozrzAuboQwSTJErt
YIlFT1cxEjIRzPvA9q2/8ytNkhJfwNvm7/2QCUJ2Ftdz76/Kc8WTplZ+a5nBqqu4
rRuGs5gQy0mFz/US5oYK0f2+KGF+jfjevbwBjOKZQJoKckHLfBCYjta31yAuxgsh
W0WH0m2Xcz/NnaBlVcphQt8ur/01KpfUGUtdJ0HJJifJ9y+bchMepz0N8RI4i53A
s9yU2jzWBmX9mKj4j3knVnS8qKKAEV8g93N3crZStpqUYNdfUw9MxLftpcIVz/SE
CPyZkKllEy6vnp2QSZA/0Aw/Ii4t4Nfld2Q5ILiLG+NqsMdlTeBtqbKdrH3TnAvm
3YWCt6Q8YNTzRXQwi0iz+XJ/sX+Hu+ubwwERsaOayPXk1ZDexe7sgkOdnaPYJJND
2q5vXF/mwtNUMQAiYosGLnlAfxRaFLeYF6g7Dz8oj4p1FXNh3ZTCld+Hnw1wdStg
YQPfy0NdYJKTuy1QSLsjZTmzaqlMyUdqzuXlVlkLSqVhc+4YaksPhR38tjYLltki
BioKxjr65Fd/no1UUO9erj1KZ0LCO9zelbqgxjsuaCVURrzdAK6OgsNbkRpfEL3r
jWwSH0p+CGHKq62f0NTIhNuLyBwUPpFkVTiTf29k5A0hXY9TYLmDkzCyiW8Hr7zu
fYMJozz0fw0DnCq7AHzQkmv2V6gt7QSxWuX0sx+MAP2juOsGqY+GFwLE1XwQfIfo
9QuK7b/AQ2llaC8uphmV/Jl+KT63cak4IfcOUOFxvFHwBXbBImpVfksBdXaok49w
GXWH3qLH6395U+U81SNV1mXg+UpQvcDAnDJPK68+mcAg/m9mqIYSXqPBedtpi2nY
Z6RIMcqT+8qw4oPlQuemjraAXMQIIBPx9D0I9XNFXx3rbOSE7JtpL+7ndqa1TI/j
DNyZ2v2beXbsQW9/hjFDI9pWWjFWkrUq86B/pi2TNBMEKnNk0SAS6xRGkzcdUB3e
0Dpq/DRR2WDIfZuWBCv/4fWv8bHrQN0bKjEKHF7oVgS8WFz8Hnt4xveOy+7+XwUl
MLwp5R3rGLFC55NXw42XkuwrZfjK/r6oT08ZwWQWxgxQeQHDmjYqnUFFPEIJwvUi
jLSTFiAtlLM/soe4aInrxot00+dM/uDZjMQWVQgW0/x1PoyR8t5TpNdJlgohlj5j
5Cn+uxx+U2Zr8CL4CVqUTPdoB7cFaW9tZ8M3kVzLmiuGfKrR12neDM1gSjscnZQx
ubNze/DRSYyiVU99b9BcCNzLJnZSeLTLB1GsdycvR3qYOZTcnj7oCYJkfTlwjw11
`protect END_PROTECTED
