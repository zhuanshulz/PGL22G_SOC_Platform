`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DM2/C/myQZch+kjfMVtnA5qRw3bCdC3NwG4xFfNVmTXqdrb/TTpbvUz/v/Nrdzjw
SJjkAwob3ymr4jSfHDcQzfRcsjF/urQ9y/DvgHUd14ugVQbMXgZVUYRekCFF2vmU
V1B1GvtO04OMHrW0ZcR4zw0LmsqtbaYN8ik9BVCmOgA8qT34xZThw68jwiipOq9y
ZJLPvr3290sTwyyXEXvVzMjz+/S9TqZat3Gg8C/pJQI18N+fakklH/LjYeuJAjnR
/j5yJvbP7G2w0zgFcJNJ9jea9sLYltrOUXU4QM0BS0WRBQg2yGTpqNRfOb6Tfc73
7zO0vWgqycnzSWZZ/4xHUnzcIDlzwBHVIGsdQkLflxXjhKyuPXbzdU+VtcguYRi6
IFytPYYRalaUBQ31qfuwvEjDkC5RK4VcQezDnqtUVknu8R8l5+IeUFF9Zn4O7NIU
+TiI1Ci1GnwTInh2r9wkK+qLCRN3RGJxixUGTTwNGFRAHHsjBlpWMa39dErqvcoj
xy9IZqdMDqvgYl8YrRw83fDmmIkvBgTGR7x12hUU9gVZatsZgE/aS/QAEJQ2E6Tg
K3R99c8D1kFWJy8BsoTYE0AG4aYtbSDxaRkymxRN/7spXm4EyuNmQCUoJcZlC5+8
V7aof62FoPVRx0DKHI8ULHH0TCowfc9zLdmIhxd2395o86cGbKNHwUw2yYOwYlG+
W535YABtveMyjAAIXdmi+CN23xDPUZ+4eDv8eOpGbzyTDg8jyii8npXddUtQS+u6
w2Wg/H0yDD8WWzTIezGgaOQ5z7igk3XbxBMxQk2XLMhy3+5fQw1QLspd5mooWuK1
CVfXU46Ac83fl75JbcSjrKSRVBkCSeGTQvLUTXNhKLAhaEUlhB9DLkz67s/0UHTb
BZg3XmKYV9Ixj/YnK6AfqmRzKjb9wjFzTrWOtJj0fgRHpzMWtdKBrJ2LxKwY5FwU
OkVrD+3mOLQ2SfC7sYn6+iiMo0o1Di+pdJITl/aZ0+LNoKLQ6YMuvTxd4e9FY0C6
T4ocNSAPTpmfSiHYtNUK5M8dLK5fvsnOUf1ovrSgqaAycfJzcj1G0+MhtXqScI/9
cwoWWt4Dv+AgOb0e22rxh6uB9n3zeQCpAQHAuzOvARVf9PcmZoPyf+QLwY6y9M6o
Ul+qPjH/Pkz1PdFtMU7mBXcjOuNQMpnAV3re9dstq4oDmQ7UluXKPebR7sdu2cYr
9lnxqL4Dtq3ZvEPVUqMstmvig1BvJW2aivZABAJVmQV1tWjraOAv9nhn4h3HxLeg
wpOma7vY+4kdYbOqYgwZGfyvOecAZ3173ph8xt/Ll0O5G83zcsPdTYld6f+tMi7w
MQD4LxJBCjYt/JJjddWGPAMc1K9ohFaQpLPwJLJP9pLbIhQObZ3Tkfo9ZmKmdDNA
cFoH8LCf1utpUsLAlEWRWyeYIGXDs9pavBzJdPhYxp+fPeT5PX5Cvd88q/gSxKXy
Ke2gL2RAxiv+asXye4lNOQh4sRT1Bl4TazZql8wYWcgzsqsRHX/QbyLbA0WL6PPz
T6E6VvtDlTkPZO0K9lnqTgFW+hfUoSyoD6gpFseLdOGi4Lc/QafFqLQ8JsgO+GgK
+Cg1xlVROmfZpYPFBPuwcZNbxrauRSOxzLzaKAVVU93SjNPKqh1axXS/HcQu3sNl
n9FVVqutegSgLfCGwIH0euTD5VztqQ0iC7e8nq+SEJsxx//f4/PqfoLk9X/cpCqK
u1Ut17wtsHkm8A2dI0LPM6RMyfzzPSGBGz/85BXtd3OflaPocOzGoaTTA0QD+9V7
sxsLlMUZizRPVtgIHiJDvi5tQPqAAESTqsre2kyuvOKw9ANtm37kR0d9RcKSBzqH
HueaQj3Zyxypogg4bLN6qLtaR1iGXzM/I8+InScd37sey7MlkFlF8jCw/IJANg8X
yv9zqmYx93Y6Jy9dSnYSQw5ze8V+SfqxZC7ghDpBfBJOLUyiQ9HCvfXCyulHfDJi
+kXCw9+ahHWYJSXGq8QoGFRiZUVjED8pBXU45+H9j3qAIi2wDmF9Ow30Zx5J8t+D
mPUD6JmEl9lflSsbdVotnO09Q4FiQALK7TjtXmDURvw0nx2vwOyKl+cHlvW4E3eV
vhS0Uk3IsUtLZZU5rQ7GKCly27AM0HTSpWS+OVwJQhB3O2m9V2ru/HHlYI+4+UU3
C81CuBlAlL+/A+JCdf5oi0w5jZFNcCBChGt/Hj9oQvjxVrqm19MF3m3i4ZbfQ+2r
wGOxcqms9F1Sb4Ropy2ffcd1MaVSZtgeg6j+JMrCUnP6G5fRpEZIBGdkhhsMglAK
+2gTjNVxqV5+M8PaYqZeoCCkK1AsIF6f695s193PlUxYLZoNrSl6FLzWdVESpBQj
LRR6yYpErvFAA+M2HkqjEUFwwcgck+Lrz3XJAcT1Yg/SyQjjKqqvFaccq/PSQMt4
Uhnt8Z4OBb7Tm+NtkZqFz17/TyOT2MH2PIojqYAuDEg20yg5Qz8rhrjcCUjJKdmK
MsRRAD11PGlp28GbIWrRef4S88tOamL+MBofsRr/EzRPn+Se331yD3u6N2QfIsbF
eNSWMUoZTIGKbcvpSQi3JwgIgLXaMccWRjBbso5gksh12aTcgpUdhPNkbgd++tN3
kvlAuz8VXYRzeszWQveIFjMytM15h7EgU8dIIGY0Gtp8cttKwlm7WTEfrknMxhzV
2KifT9MucdXixNk1i8gDByNTYs81BU9qKSB4c0tWCb6HseMd8UKbx/kmicZTKGq9
ipEO9pQF6uDMqQtRLmbGqpyHThEmlH8oym07t5c/VT5kAJj8LqMCF2MvnqR2qH3g
vStcGtTsmEpknGfQnnXIAtJnjUg/rsQbyqsUITgbmGETx/2JlxqIvr6e2rjj9MYi
qOX4e4tP/cgG+qaVJYcV5VFHS84D36JPm7csWmvwKxmFKpCNsGlHLlMEk/XWZhjA
0ZaItvNP8Z9X2ZySamFnPBtJ2NOFZAsuQIojy03oCwiUH8YNQy5JTPYEwMBGcCuh
UCO4nhmRm/xZHJoZclWc0aurjBPnMroyxU0Cihg6hlOq7EJNILPKN4+U2mJGl+f/
X7KuzgAb1nn0nlFB6ZAVwXvxee9JmzxNV9s7QxNk/KaaHzQ2WQ0AXhrHSzVJwu4l
7tqg5dvGz5mAHpp5UnUaXA9ydKZ3a8ja7tBoObC54PZjw9a5VyjeAfjvv+Ptd9t/
evi0WXvMJcRa40Ff5+VZ5biTYlXYfklCYkljtDVRXMmWTqxeI23hvyOCSKiAOWj9
HiHT/egQdselloJDPse4Yw+i4+ob1Tq/LpWHDUyKiww97uMIAoQdkidb87w3ptFl
deZ0G60bxq52doLg0rdnsX5BT84nH9iWaj6pUsp+PV2T7CqkA9PkEJZRkkl5EjWg
LOuA0/I3YUdRSmqSwR1xbw==
`protect END_PROTECTED
