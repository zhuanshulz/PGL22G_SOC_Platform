`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OaAEM6WDkWvCwA4v2xCUZ9gXhuq7+lierwgadd4sFyQ7sQD9FiLurSPHHTe8TsF
B72EwImb/XHYQ2wioabB/3G2ikPv0Z9SfvflZmYUech6kdoPubRUhntd4rIiG5T0
srdDQk7n3J5z3yyKQveWsRlaoLreE/kQT/z7lJc6aREWN3IEpYvtktxz8dKN7TzF
4738ELCGolBpYXfwR095N1VPZel4/QswegsaEc6kQznCwNxtYKxGiVgo4ZaUVO0Z
I+Po4JjtYUaXb7u3XpxCbfczlY97u0T2IRMcIx2rBoS0oSNAZrlpNgfWcbw8HaIt
ymsXW6jKf5LdxJzca6ETtsw0QoXVVaz4c5gnjEiWcZwD4nOUOEz9cI3HPFvRjc5v
vGG7/tfqN3lYFE5Upopo2z4oSF6YJ1wYQ+oWqWBQxqjcrOOVxrcRoReXfi5Mz/Ls
g18c0AhX1530N9drkBRALNYprgaHku3EPiOrZGeb9vx4jVzvFGWD3lqbiXY+N0Qp
/s1bP/bgRZil+JpxKdSjh+xHkP2ee9F0ueCd2cNen1oWvR3qzlSVho8m4xORhV0u
9yaURoJwvY5YvCE+hJDyP+B5Laq1Uk6j5TAu6s+8aEsdhDLXWZY9f9iiBpCHT/s1
mIGjERFVgUgcMYAWgfpCy2X5OlZGKTXCfrekIKNrQsPoM1iviMxtxpmIkn6q9oV1
hCNtoLqkbKDRGJxX3XvpKV5g2yWY7MmcjNMom6Efc07cmetOHFNiftvqC5mj9yrw
4WUjMXtVQw047fo4HUv50qA5HoSxJg+tcEgPKdlSD4A4gQIBXI2q8LdXJ0fPWieT
9lez/pgtBLwzKxIrnhoziUEBJ75Vnr+gSjAFjP8SKF/xZkdUUwUcSw4GzUy5O5JG
toKPBae97rtgPv5Tgjh34EdWa3/UQ9i7QHhPyerC+RlXeX5/k6nwJqCBZ8yFktwg
SoLiZvnaskO4hziAJEHvd/aaw2vCgrc4WedBngX81gOBlof5JsslKXCnpmQisJOh
Owq4GW+Q9oLjz1kHw/lNYgaFDgfzKJ2Z3TeGO9f0+iYs4Jp28TzLasd2h0OsucgX
e23YJKAGktCSEib1c5x1NnM5NPv60++9tlZXj9Hgc5u5gHT+sZXmvnvZ8PF66yYx
ut6bSPRhWVOSkBSICernlLyf/+H9kfoyMrEwzzhI98n8jVKYCNCYqwJiZmKM1BNG
cKr3VDKITX9Q7Vi92sLf0nATgfkH3DSU/Y7AvTd2WWvkG10unptQf8Ih78GzQL2o
XN/d2TzWSKlLh7VYDgmCvEMN66qfVt9m4CU90wruePglWTAxjzK4AqJdWKpieuCi
Mt9YFZCVLW84b56l4L2qlMrbOrmPhsyOEdhKkAubClngMHFt2NIHFzrG8GclIa/x
WpxUcD9MplHAxKGnR2cbulXzrc1MHeyYC0d5vcXRTMS3/Vjfzo1oEMTyy4eSdmm4
o1j6sV8YP27nhbPmHy9aC5mkjTl+9uAbEW51l/jKKsXqp4wk90bpm8Y85DZP+Di3
PCqnhe2wTYtK7dXEdXgSep8ey19p/EVSZbRt1gir1w1ELqWmt/OHc/qfaHLtwV1v
pGcu7EwU70u/Olyp0OsYUORDOyrdzt1+qG8iyviz8ERu2MzB/5bIYQexc15PqUKp
55fDDjbWxeeKHGJaLWwawdNuPxaNKNWPRt+D2gddbYyXQUZR/hwNDgw5xm6lfPFZ
PHYaM8ktXhGcIVvyVbvXwa3oyChcHOYfJJMF0pAmswGw+6VH7bUtfIIxFKXqe1q8
tU4XF2y2OFmO/+X6pscUzumQFIOcVi71MG9sdS3P1c4GfdL7pCWSbhxFvEa3BkMX
q9oaVHcNJefDrHykjtJsOG/dU12ykqChiWPqmpwlTr7unK6ijTjlYfLIHC/ZQir6
0PkuVbsKAGKCSAhiIxAoJZy+TspEQ3FD/NQLupGO7O++kKUtccWEITVJSzMLJZSQ
5kYFSG1MxCtoOyJOEWyJCzAL95fVMtphRHZgt17l6H9XzUHEUEORulQlcwL7AcMZ
JkChoqAGuAY7KU7GZQle39VOZnplwFNXVnrcUWrp7T17PC0Prpt/VWJCr69aV1ZA
gWmbafCe9ymmj/Wd/+Ot665h2DGhziHS52pNEkn2W9fdHWQyAmBjej97zOxl2QFS
tjnxWyqlIjT1LdcHJ2jEPJgmQ1gSL9xWf35w1pA2vOSpE0yi+hPCBFoBPFlFkswG
asRdPQlNOQLFRLcflxEq+yC2QJOrsSzUpln0/TpXVjpEbNa8hOSJ4aWj8kJQ8Cb9
eeVgdETTn7K1HOCwiAUdIv4yTjSNzACnTwqiXxTkJ4/hWNfjjazugZb+oELcptuz
jk2kuawUcb0GtWHmw7Kd+E6wHo++K+MeJDKN1a9+aiVYawpOpOqTkrJNukiyJiJO
80jPOg2LyyF/XpUP57SXTGYwzwVA9vth91/0iGux4mumjHmKyHHakR1SRVfP7C0R
0Bo+5aiO5VIV4cyqWhl9YMgb4IbYOP4Ep6XtYWh9L5oen0J4tOVkfN5URGEGhfWf
MC0fHOfJ7P+XU74I2oX4XOTVulbvx7W1M0FiZZTLNUT6V7tUn3hulxFNna6MAbSv
CHv4w6+SaTlTo+ufEKkUWkJDv+WE6uY39bDhKaNPQeqZP9fgas3876nGUaOTgylG
U7ODWhX2GTO8TETBggXfo+c9dXwUgHp7Ur0g4ukYK1U5Frt6qCaIaetbdgBC8TFP
9WWvlIC9z0LNpMCsP22xH+FnanuJLbkPcT+PJPcwUElaDblImKJzt/oC+KG6XZts
gpiqGAWBY4yiWb7lgF6pF1AEGyTuQNNjS96l72r6s1cCfnG34MSMURUwbtufJPA9
oXRLSmQXcCFRx5Hqvjv3pMbb9HxMUs0/57Rd0G2IHc0K83be3zyAtE79jU6P0Ndp
arEA8Y/EFBLqnpf5FzKzokueOvaAuZcdbSYClg4t75HpiYjQW5Xl/01rpCD+NpXy
LJ/5RljO3XdKUqnyxGnPvUzVGB4R0crXUJqL30kAFn7BS32FPGyRz6E8Km3KSyFr
L4EwLQAmwo1IYog3ORqGDtVjYusSx3o8KoUI3lxxREmM0ItJYaqJUhMM0FACEexX
qC+IpAss2NDAL+w5jL22Nm5ZhUtFQ86+yc48+aUbgLjFgrEfJmpK+87rPkTsZ7a3
Q8XVhU8uTgecagAHpCXTspwgLdB/TTRg/3vTIQvME3qsiOLNNffsw+WktiK+Mr2J
KgmrBdGzY2OQ6nYqHCUA+YW0vfEO4yQZBzM0xLAEiCaluAyRnsDTmAyHH8VirO8N
sC5duBZWmS2GOVsBrsnHjaiH1Cs8bbOMswe2WXgfEfDumvio+5yxH82KZKlvSuy4
k6niA8w9rVhS+Cx8FzXJBvjA6to8Dm1Bj/UFArVxBFA=
`protect END_PROTECTED
