`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cw+vO9fkgg1hKbH4TLg05dFdMxYGDOLwS3eMXHotlMUFVtT7gif673leLFifsevZ
h8xSTM8ztgBS4ZN0WLkMcvurwNfU5B0+whggjRaJloB7qq2K3Pn9KpKv8yikDUrV
JkLVdT6g0DQWbXVBu8iv1a9+dDEj6PhShFeCuOGWH4CwBa6X2XBaPaaUYgFZzuNa
ZfrVTr59z70M4YnU3ibrZNp9pSP6iWbDhD57hrOH+qYjjMLVGDliHppN9DpU+XQg
U9Uv7X4igKcyr0miz1KVMEb+UftSwCG0EGa6eMdWO26Mh75aXEzljs1VxyW+BUrz
LzpFivnV30lTUZ8Wle1CxSxAqHt/SKMonsFKHQDkg9hPkPVTPI/5Br20D6fbkXJE
spucgYZjVg6ZHrkc3FBZg2RrJ5aGnBM2IMxTWi4WOww=
`protect END_PROTECTED
