`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQQipCy82yXDLoNDFbjOl1QGmqUm5xUXQ9oJPpr+/emmV0QR9Iu8dU8fra6rTde/
A9At0I5E6a85DxYS1iWCko32B9PKIPQ6uB8pUUGYICWqW1OFdl0ayGyAEIFgmh8h
tNoElJn7D0CD0p3YRpKFe29kxGVvjEaxBf9xqQ50+VyILGSuairHsbTW0Ky2Jxx7
WSFJr0kUHe/DY2OOy50cuM1KnmKbWkSHngXCjoNnq7fohKZEmx/wouNgzi/Kuhai
v9eKWfjOW4ZFJB3LdYBqBxT88EPzHQ9q9SShgtjZHOchU+mhrX+y52sxmIwZg26H
AgQooQA4a1JETE+j4KvhBBD73FbNxUDapZCHjnyqj2enLLaI7NDx7q80QG8LkKFR
BYg1mqLc6WVX6M23f4I6iFErOP2hztW+PU3yCGtO9u1UNXAhHRIeU6BCgwBb5UmG
C/qgW3H9Q2oz168GLKHA0zsjmq6btl7m5LMS6r33GHjJTnf4qSCugAPwNvyZbuVD
neBABM8PrTdXtaHzA05h8lXzCIJ2NGzrA7z4h5WgWhj9q5960s9eI7HtB8YYEUhX
kup9KpfpL7t641wWOgbASA==
`protect END_PROTECTED
