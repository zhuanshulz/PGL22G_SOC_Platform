`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DNH1g0iXqYco7wXqpWeomnH0koRlp3lYNYEaR8134qoWTT0Tmx26pUW4XX6YvdKw
R/Ec/WpURuoBMFRCGAwbotgpkWoWOvh/RDLi69OmVE1C/v0oqrskGLMj+Ds+dsAy
rzk+4FubVa85SE+4f5Kb/fYMxofNRK2Qm6DQjBmR+UPChOi52svVqfFCLh3zerHa
J02yWFycvrQw1B3Qou9xUxggYX44kxJ2B/h7b2fzagbenlG3r7gEWD8nadYu8yEe
9hOfnXtlltp1ZVMYg8Qc0Fn7tnQ2Lq2fS/H9mNV7HA0blfHvKtuHTURIsPnY5we8
QT3O3+H+nn2v4BfR/ZQ5l41qGkm5GJrcwldmPCV7m/7tyXu2/E4wKO3fmG4Fow7C
3gzNs04mlvZwwgiQury3HmYXxEPl6hvn0fmpliOGCGlfUKGzcK/bAvoU0wnc8j1b
/xZzPjTxaCm0c6ojp2z4reKVTh9/JfI2FqqzZmbRh1jl3FeDeJn4DP1KLeS0+gVg
E+BhPbsCOJ8deuzPuO+Y+Rqu5jwYHKSzZ+kNV1qt+y/2vhIT4LwxZO3bT+6hB4Hg
OXIhA5DfYkaaGVmLL24zF9Bxz9jEW9ax0M6Nai98Pc9bOE3OinFeJfyA+56lpCqM
hPUd4P9SiQ41gsFXJeXTQ81GNfuS3mlPgrRdPCoTMmF5WSJtzfUTztQndn3ahHvC
ZiS6tIDqCJqApHKELs5Q+UqThN74IGCb3CWTIUMzeOOQVpxjLcoN6rrHLoRbff3u
zLlZT0NZB0/Qm4MV1RZQ40W3S0uFneCFfAkTbp/GOAmzoZsRSHsbWkwJav6a7O9o
cDgKzUb/1uETNpZy4/og9pV5A3otlaGaVxcjsCKLyTZzYxE3ceUqKvvkRJcWE6rZ
bLbCdTCUuJIuMrhUEnWhtENHr6NIf1qc2VJc8qJT+Dl1xMcCYs+OZ55MF4QYxwYq
MDm8IWcEDW3k3LzaFkOrCqe5gGhyFrj98rvyQzW7yUkTepqbEFi6j4BQmPDstyAi
Nr9iRR9lBhRnLaOxo9rxRgi4+32qe3fwu1ItDnoPRv8bvuOgVJYcNP8AN/dW6Cnq
TvKpskDzI1r+xBEWOAzKOBMPXHyTqrMcDiMgzsOW87d39zlczlr5BEdWhOHQMEBW
OjSQao+iREL96mPnMefnoRUk7M8OM+q8skRgZ3+TnVqBryo46uO6MiTxI96O1Rp5
LP5NFZ9zhr3mvQtruN9sZIDkhHGmS2R8KkRQh560VXY8xGPGPl3wP7Qhrwl//3Cz
m+ySxVz8o3tky8PUkEdTqZ/vcl8Sk8jhwjA4h65OjPyEhv9OWxzxH/KfsDz024ID
MfcmDYE9lbYtCIRDpcnBAIE60S9u2AahF+PS3e4kpQjMuXz7VXsPpkd9uLKgtehY
SnwkC4YlJrFoQJc+1AkKAD2oUV7kIDm60xTPCawGxnC4x23mKIopCGT0/9Uogmz3
E/s53QgaviMvSUlcvmxZJ6FQk8v4rMo311OIu2YL7m1pBkZ+hYxeVDEx3JT9DwXs
vuC6bQCNk5P/tD5q9Rx+iZPsJYKAOj/tJTQuoicQW3SkArw4Iixb2HAotEMrEH4H
fufuLz9DVH7kGH6r8RpoMHd6o1aZvGi1WOBT7GiVTJVmmDhXhS4TBI79sNj4qwVS
+k49hjV8TSwbA7g8Y1kBMS3apW2P2f817CTDGZ3aZJgltGeWNtT8njlwPq2K7E4h
IMlSaqvk1AK/5cF+/KwrmLKCU+h8Zlo+6OzBp/b8N1Z3KVYJresZPCFOKueZnsRV
H/p3/c1v7iUTkDCrCwI2K8TWbr3ULJJjcZsOUQAAaLwoAEcO8RctkolhU4eYnttc
ojSfRrTaTr2sJ85KnaBDVbFLuf86krp+6bAt2pl781jGaLhRX1xdIBST4tF23dci
6U3zOJzICLo0dD3pd2cRZ0nYk0uwFU8Rhjf2OK7r6rTW03CMmFYrztDEPtnLZ0gu
0MK8QK6RihMfTVXeeL2ynvyE+GbI5sWDlxQIo4B6SDBgzd21R2kQ727R0y5+mqNK
0RGM7ch/HFiNCRUUwF7SQypPWaza+gl11IcaDUId7Gj9RZoH9cGG4cOx2l0K8cFs
clQk3AGsFfdbcRqKz+SnuHuA5wo/XIIQ1ox7IrRKCMB5MrjKcL/WgfmXIBkuIvG9
TsJcQrFy+VkiKUhE52ajKPqwSqUz4GYaHXkjT4VklpFc53TnZseLWevFaEMl7PFk
6O8re/sijCaVg6fQtHfhYHCXA32wVgp0rTdBMvTMDE2PiwNujHCBRDxd+vOLPeKv
gK/W+nPKv6V6ME+avi5yGumkV89O60ZtOAEu9Ku5ploMQzKc1Z0AzwdH9vkMOa31
5Mz9N4b7uIApruvGeHqq5MIZy+r3dG6Z8TiX5t1lgwc01w0m2BNGmlapUmJ/Bjkb
d/Ifmor6BFL1F55Sm9XHRzateKSbQeoxyr8NTbl/EC5UAxBhIP2FJ5U/0vGiLjm1
x0QEM+L0BbxfMZc9/cIM2asV+A0OcZOyGW5XrGD3chh+p057YVHYfdt1Lhm7i4aH
8tTQpOJl0BLUafGTA+0t8lPpnO8MAM+4ve6gYckHIf2S5RNAc2pZI5NBWwN9Dv5/
o6UaBYweUWFszai3GunkwfAvpP4RN7iFJspkAvaqZoD2FH3Q5NU/JnBeIYczRgXA
yb4ODYw0DeCQ2NU53uxdHKEALBIZC2gxCj2XrXdsu27alvuckcUJ+uMsnMEdybOX
4c1PuGKYHCM7Cl4ojD8JoQm8lJ+R90sDcpGEZh6fHoOAbjHbmYoQKNmL/xRZ46y2
A8/E/kylBAKGrgQWgxdXKrYbIRjz8ViNJAX620O/8IkXcbx3KKCqwXzbkPffF2yc
geheoSm+YEKAALeMXudjE0cQbov0GLMdYTnPNBA6XaApkoRpGFUJwOu9pief1P9l
Ll+5GKlSHJYjW9h60b0lkoVHORCQdqWxugW8YUH70YZQfluqCxTwWR5YRvi+5C33
WGu/RiQoC271DjxhWNvSeeJS3BnWJhxJ5teP6o0xGa1yil06HR/ZOnueX2LfiTKt
z9FrM2Jyi7sjCV4ntpgRv1UlhuvaqqsMfQ89mX7HLqIHhwnQbRBx+gPrkOq8dKEW
zwIv4qyXjdeXfEdd2vYvpUUmK3eYV8mdMNe6QYNdTS3cbGMhl0RCgFY6nOcdo+QE
3/KCQZdGZ9qIzw3/2yJeojnfeN6jIrHJgDQU4FQpgMb5NN7jEheBvXcsAxGmsXyw
K9eltlOe9YT+HPmMK/Gg9llX8uwMdZjGyI2n7TryseQQfqWFXt2HPvLaNtHYfZTH
bMvA7UYIyYngGx36u0NXRgDMf4Nn3FA0FiGpUu5Bdozrhjj1+MZnMQu0IOEDge8G
uhaQ9pcwIP3bGiiuI9KOOE2mBx2BcvCVwAgs6jV0eRz+ckxqt48QhInaX8K8ih8f
zlpSj8s3a8ch32WWM6W063Fa1gQORIRmwWiOK9GqcHkrK5Uh2gz74beb/Rkc3hI/
PmheceV/wWCfMJY4eyrw/7v5yyXgS5ekBhCLyhV+U7/xuaTfuca93kH881n3dsCo
enug/gmpoEMQEBvbqWLhQU2/L0lHfJumEmsaI8p8qQPRZOjDBv8JV4V3v/VNnT7h
G/ktjyChfy8t3H8mCcsAhrFfr0IkLpZwxsQT8fw7zQjYTQWTs8SHuEl9PZCQ9cFQ
VqSBFuX5pTuIwBEKeKnXmL/Bl2nW9u8GYHAnVdddIUfE5/ZgBb0xRE7Cp9n1khvA
PXTWimZ8z7F6o+jbde9DC+kbOjhBgmOTQZfiuF9vt3MrgMo0rSIdn91sNW3F4Jit
We9kGg1GOOkiwOVPxYzugzXgxETs0/FkKFoKT+YnyavETdQdGgZk7Nky8AH+43Qw
cHg8WSrxCG3yg4E2NwVI1Wj+8pPvClZIEcPydcOKs8MScCct6nbDVWek9Ufmr7xS
P+Kt7+HIf1BOZ1kKR4Wia3Gq3DddjdDXsWdAlplBXMKZKRc+3drgp789I2jKwyKd
OGJ44gPJ5Bswjk0bb/RMOSDMpBLaWZ+2NQHZAJv5Mb54kKHQGf6SY5596ZFhxvx/
0DO6jqp4AINfLrMvwy/I8+n78sHY6R5hgAwbqSNjF/lAj2HO8Mrr8oLAAUetWPbC
heDj2+e0u4QgJReoDSAigIiSojOYJFwLRXWfPs0A9lytkf4zmRvZXmye08KhsMSF
wX5NaY9RwhLqQWREKk2Ef+MZcpY67VEG9MdryVI/Cy2BTWSGBmsEI45mNiWtcExH
HvMse4+Xylqszuz3mJIVCsrm2nTjA19rfasIbUbPFEIqbuLsInbQMqz1dpfQixUn
+olzYVLLTXe/m4YbeElHE3sLs9r2yh1u1DYn9Sr1nWGUSGfM0StfFSWqDVCgO/Nb
t0tfZnISniyR64PjAd9veTf6xvuF6ituwOtZUr6oBCQ/yrjOWpMtyULrybyal1oM
OX5ZNU2uw8KgTLncJy4urDV5QJXiY486xQ/3DOFzXwiJuBaNaPMyOPwFCMU1atgV
9hLmoj8OBXhMJ7mqZxcCu4OowNwEXdp71QQhAgyqEwM6WldDeKOr2veAdBgyAl4L
2xC4RHEw+gBhQ7IaV17Wt3MRMWEUn5GoOoAI2QSay8kvE0J2OaafHw+GfywlhtVu
lbeAhrthm6748gzfGqNI1WxySrcbmyojozFbJZdR6MyTk1MQqdhSgxr5iGc1YHcd
9D7AKhuKhnFUOtun3IsAAE8tKBrG6eCIhppn+fFMZMEP5hLOEJNTEcZXyaXQb3sg
eq9eqVNyMy0jfFGGLVHcKMo1+q5yS2/wk7PLIWLzQEW/Co71X+md4aUVYVKYn/F+
L+6DZEWA1ztjug9k7Xh4uDPQqiZgdV1C0OgLmAbyfnHncD7/52N3eScy4JJqE/fr
lNvJ9d7TgyJN79zHm90/xvVF5m0/d48Q9v5JDRWJ2ML0khPKxYk36iqp74IJzzRx
xaGU1EBhavo/RP14gXQIO2eGwS65Cic4ViLRa0X2hrwIODIWyJl0lNRQdDpXU6jK
`protect END_PROTECTED
