`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8F3eGkJA6pMb+meO+GySPVgPFm11wy7arBqg+um//SJyZ0SQhFW2af4/FKsRRFvP
XL6d/7IIUW8rAPvEWoCbZ769DauvhQn6AQ2jcMI5hmwdiWv7DtoJ31bEqECAATwx
+FKmB+lFy8JDGWTJ0ktXQrGYeejasExO66SFZRj7uuCnfyWpZxoQP2aeNpoqqq6+
QL8fh5VTfs/kfJLIiqZcbuXtHfRWCpvXZ3GYENp+ZIXUFfo83VsRt+eEPfVupFft
CK++iNSn/4Do41Znxx6yjSbf0H6VRtAlZaPna/QNX+baBRSWDZRHsJwccZWbU1Bb
2e4jR6oN1MkJX/ezCdm+zuWpOXxRaO7q3GnOFekvNVDm3SkfYasOTXwRK1lTpYGz
nShX1NZN2WYPFmYCBIzA7hHG88PCbKqu/1w8Zdakrayi/hM3EN7bU12bnXTdAljI
RC9sphPHTx3xB7r4GASLIGNXnzWfJALS2QInC4qM6hRSC9ly2EOIiu1ta4tFcFTP
pOmU1nOYgX05Uq8gl48jcuq9nH5QhNfEWMVurL2hN3RnHFm0kbBWmdknRY6rk8+a
/Sb7XRKL/4aSk6KqMIGffjQ3dLvsDFA0qcbX7xKfLChNcLGUnjn3OvPz/Hu7jGYt
XDP0nmZi4243K1ZkTJiaNKb0r/G29du/Vkg8wNv5WE/bIIhHR6dXx6kbH5JQ27hR
oTTv6ztlcpfzsFXpwuscZZBFwc+JOkheqBfItk1u+uFNGix8hHV1CpDGUXu2bFqv
GTJXbzjw+G/LjzLBEVatEKeq7CewgEuNxuUZtv7M8zAYfpCN4EtC4cjpEp9bE/V9
sj4gJQB+IzXZ1kQ7Gz85itjJPHSDnGgmL85zqOwn7cFREnLgIrNjJtJ6sudCmF5o
i1V07t5RLvYiPn8neX+ybyl0rR17XU/Wui1BLbF9hUYVoweHYk1umtPXVArH6/+n
BWrFWrfHcHaDwLN6KqQYnL8K1u/gE0V7aMPcuzdMLI70vyNKxOsyV0nXv+rHBh01
Be6dA3snOOC1xV7YlRk1HwUi6wIE0wkbGHDWn+qgSgDp/9fq8RJ/S0zeT697gZqk
x3ZVXQSfq66KpSyN86HqeE7KUKEYq4qd59BuWl6CLSti4WlxRMWGa7PDxJFPtaUs
UsKpQoPgg+aHJsj+eWbp4km3ab9n8D3s9LmFTSzJUNmmki8bRxt9b7w6KvDBWh9Z
DRqTlGrNLEeSp5bGDVRm1vfJBHsGVSChIRICMG1Pi3gn8XOna+ppbBHLRl9K73nC
do2cwwjxUzhP87wkP5mWOv9IIsSh2xSmQWIfMqMUF74/w3GGExmPMqcWuzpnde0+
wE6aoa9Mi90yNhLcrDO1iBZbCjUbjH5mFNN80I9ipfuk3wRE7QWX1xCrc3fvwBNz
L9o5n8hPWqzEgnUneV3hfW/wdZqc3+X9pvAZRWXzVdSLccyHNLFnR68Hd/RdWwIu
FHW2eJ/17joKFU+qgNzZ8He6PijUb8UYNxZC1Y7/gaYmx23ZSz7SA0phwMWfjTUF
ZarlKqgYebNW2tVAwU4g7SUJaxS/UJixmJotCa9CjzgcROIfrbiR8EpzkWS9slju
40abd7VWjEq4ztJW/GDjZvFx67nEnkHT+WA/Tp0M8FTA0dX57K9WCzAUDbAU+xDT
hTz1Emh0q8cQYBDW45TrG87IMCnCONbdkixC/AbgkC1x9Ud1BEcyqrEOLl7QInsg
fGJzz5ex6yEilBtPNlS91vvyS7v5dXJEbcFlQd/XKzbV2cw3iElAwRCEqudcoAco
M15/UhNNEveC5z/lM4vusv0aVrq2gNxgx4bA7qIoU3inhIn+JQ6VfcXhAQWH//J/
QKl5vd1OkJHa7I61fzsefCuGlfT79tcnPvs9Y0mhb7tC+cdY6wcLEcb+n3TEZ9fg
bjgv4sK1V9NozjH5kXIOT1VL37G5TyQGCSqEUTpB8Jbiluvw21gfVtt2Dfjp9O4N
mhPzsLD3qUwmRA7NxWi8pQyfa6TeNiSLxwq7yyErzHs9sRfnkB5J6B6yTi0M96dO
DJVwIZrbmhxjRky4JJnomn0Egc9+Qd5mt3ggtHGVnI4oYkBc4vQ64aMmNobcDSEG
eMz0oweFYi0pHV+hb7XSW6m02R6SAMyIqhF8sAsjSmZuh8VGMu03EN8AFRW0TURz
qzWmfM2yEap441lNZRxhnmm2wY4cARsjm51ptSLbE1ANJoW4SmjRbTdShCFabqIs
k5AmiS8aIrFgapoZm6rqVn9owJUbHIepgHy6F2y79y6yOJP3fTIz7qEt/a52latL
0DOSBvJbRTqbv1y/ANPersPkjjO6h7mP5gNRSuOnNYJLHZzz833cIdoJr2jsFfq0
qNrosVtTBl5COvwKDa6tSqV0lEAQdNTDK09PNUMnMXrx+totBcLwn/zRkKiIazwR
dgeSF6I0EyfNJZmblzTrsDdfr36Wv/dwkYoQr8WpQ4x7IrND+RjOkO4F87naJUXh
SxzuRESVIIw/DWk2Her2nOCk6EFVLB83O64rmk2kFKgMI+sPI4rjpWfI2dgQFIOl
GaMR8z3ISJnloW16Nd56JsK5pB9IWoDSfUV8NOun/3pZp1F3h3JrZWrPqaZV0Yzn
v8YGlhiCkHWx+7hOQ1/ttiQqsLld5u256VKWsO3BO97vJ01Zzsd7xUcAsVQE1aGw
xQob6x1chv98VuckCK+bH51IxPzI4UZN2L4NgzCD/nQvS/2J4uotPkOOiLfpNABK
SzllijIWrNDVs+DfuFgLLSqPRIPg7IK0V/BKeDC+zbHqENGJSmwPk0qcU8t/tHH2
fx54HCSFZekfoh1NM4dHTsTn5YKXl5+sL79PgWDIwzfwFgQ8nuiyWJHT6VhSH1rQ
bQtQBh/FfY8Iq4LDpufkLdu7hzefc76wobKoCcwFYfw=
`protect END_PROTECTED
