`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F52zCZy1PoG8DPin8SP/cg/tKCEUs9zX3134BVXhK+GFAvPmeRR7MCnUgwfpQkqR
ZRtaVkbDtKlXVjZwVREYEjQqrZK4M7re6Z19lwwMvdqqaguTGAemCQwTOPQOq8ei
fpjVEP+x7h3T3B/1JziUuICBHHOYd+o9Wph9yom57QBEllk2kcOG74yW+5DV2h6T
IjqO+EQHugtD7v+5YBT7XkiN39f4bHW0P5SN2XNY/FPmFkb0SNhXArnJHbkw5tYs
EhM0xWPyxkvx7ODCXHVPL/Ou3pvwAgKaEAjTg7GwRiNV6C6TTiykm64Ke68I8Rdx
AMakJjpwJVjKIRyUvUgr6A3uBHHE2LQkrTxb7+W4m0lnp8D5+1iRflb/4NKgL05i
WVjbsFHw54GrKLuCFujxyXa+KwoC22iQ9HA5PTrSQ/esSeoTqiMSiC5TygZxM1KC
LcHkkHwyy1AHXGYbDr/f6soAFZjjQnIo4+O/yTlVsRvCPikzyxTvN1Ch5WFIcwq+
aK92C22xdi83rNk0oa1Pj8FzNG4SqVPSUYjMkwwW9hrT15FAq8aeZTsh+A+sCgVU
wAVfjhqzekFoEzQMqWH1Xi/5HtYCFZSQo/HPysdhzj7hU9YborCNU+hbNOPasgeb
iArX04pN1KzrCIM0xd9hsxnyYSvQBl7cMMo+pefvZYc28h7Nt8+lSbEEqDC7qAzT
KudDLTM768uu/VgsZVtBxlrsJRHW6N/yzjYKJqCP/KxIPE9/xO59ty2OfYcvkUQ5
bVFpPhsuBdLPXoTwSked+eDZj522W+FmP9fgVyTZmhqyRYo8mIsrD4BHri/kdBeF
8IJWP/C8J8FjNqFoeCBCUeV4l84GAFmGM5dIg06yrCnNBts65sa30DJzG4aqbTGS
5oQqh99TCUH4GS9OuXUkEZIiM2bShpWLZXGwsx0NvHk/Od2FvQRSGdn8/LjWGbp9
x5Bp8MxmxFLknzqJjFNgV4bHx+xJU8JeVYQkmnty3nOHVlJXcUTeGGKbma+mehOh
2f3tJmGslqj6BPa1xH0Na2dHpSm9J2rOSSBqc+3ZTPzfHzegeyWZaRuZ/5CROsoP
oZbO2SRF+Hd7JfYY1BHeC09zb45tIaAOVG+M2PbRwjnSMwd5AH5oMFQGHKuqpOwx
396sr3aUMK9Ut1dvgLkz7150wPh3/ztUcIHrKVGd5qUO82fvyU8miIWMns/NxM9Q
KnBR4h0EBiY46KduYkMu7eyBqhcFObTJLP+LdS0inyPm0raujjnSJnKI5E/hyQyv
UFIZuhIXseAaIHS+pmNr4uuBHBjHgFtXrmVT/jWM4gn1Ba3fZfDtmwiubz6OV7Ur
wrDm1JKPMMemIoZbbrwAESHuY68qWoJYczzyCnzDXdFIjPCPe76DxkjGCGq+oXi6
XLUrNcrjv/oRb2Ns7rJel5Mc5AwWfM8R9a6ohMIMpwhs8Dh6pKmaGUnxQAaRe1fF
xn3JSc/NONBdvm5F9Rysfn0lhmiHea1gpFm154ivGn9CaSNWlp1mghcALWeQdWCU
8WrsG4HgXuaHhnyphFL7iKUCKb9C/vcijIgvB+VA/A3zjweSCKscle4K7FKED9CC
82NgH5B4dVFzPjBUbB4/cUjJtsBnIHjynxHtsEC9r1dtsS3qVjqTr4lw6zg5oEDv
Xlme4AIXQoaK8PeB+G/9rLi0eJ0j7TEW4Id0Ir3qRT5jL1rr89pbcBFTICBAWL+a
9yPAw7tEm0qnGp/mWeORRtj3RGgJKw5T83qFjRqGp1XqclsQwtyz01E4frDbt1K8
WLnSHE1azeAGcnlh49NCGT3Lgmr8Hr/W1bYJkhPLqABfleylUPjKqGNLXslPYRVn
8yvB0DDp2Ytqv0pRSaC2RmnnOKhDInfFdXC96V9nDz85af768Rh/Q2rF0PXfj4i6
ura47WL7qxTCoEq+5/6nu1TXizynO32hHEE+qZzZBcHKQXXooTQ2uz+/xxuEz6l0
EJWPN878IMgSRNuBHOh+O2w+wJYJyNoD3iHAmSbQoXczHLL2l6FWf9pjh84rnxQE
yf7IVfw7QzDHKbA4Stt4tqHR/pN0eBfjMCPIm4K+aeLtKSF53F3S1QFxBaZr/QB2
JJlF21LjgO/NS6dbLjjiUbJp6+fNn18r8OhhcRrSzrf1u+JbJQ3GybjZkz0u5X3Q
Y+r1Yl1AM3a8ohB5f7wAOg/HclrixHeAsVZ7RvHECOfWwKKExCrc2ao0ZEdYbwlm
ROS5i4MyfKQHRWM0YGMvbf1tN67v2BpGE9bq/RmK+LO6RtKKywL+awsekOUI+DrP
kNzfamhSL7VfHL+GTPU8KJn+5M03ltnVhf2Vr3ds7bVjkQphRAGyh318qiedD8Q6
e2qQQUzUaPNZAQmgHqBtx5U7szzsre91QooSX7pgd6Jubg45IRLzW2BCeJmb0rHz
i92nhW2B/wwjDI7aOxZfRJuTq6nJddVSnjsff5bIRJYcFD0DRsZESeuWipciAR/y
F0YIO7+/IGOPpysfKd/pAZeR4zI6ubKRhh7N1QWNjkoSVWXVLikarEfLJYM9queG
HRFVWBU9ZVgTyGZYI6AcQuNR6UL7mr7ZByI+rzXuGVsQzxVijMMYwjrDGEgcjUDP
41aD2FnqMfKv7Kv/GIRGRRdm9ccdh3YAQGwQv4hEsaGIv4EVQwC6KgKERCEBOjNm
nLOhRpKbeJ2yaA8n59RevPX1IXsrwccAFrijOU1488hgeeoTKWktVd1L9psL3aYf
elPB6SIkXegU95UhGUaiXy9TYmjHWFGeZ3e2tRmbUEc8OK9PemiBKKY4jqnNpASZ
1SQlAamyLagk99L6ojNKQKXd6uzFrhXSV6BRQQLVVfkf+E3Vm9RVT9y5MT6zQgXw
AsvtC5X+FjlGi2p8EPnNhs1yJVCkR7UaCuZiXa1AE/A65zNWNTQWJdrzCiedNIzw
Z79ygt5k0kaEDzF/abu4UGTamRFXcZ6R+/X7aldhbg3AI8EuPM/o1O5BGSfb9aTT
NbKLw9rgYHXlCGwRhnSjJD3TzOwVF4Uw+TaHwdKqcb3P9DRJInx2metdcnTIvLW/
ZbneanVuRGsdiaWC3Z7XKCzRhuL/kOy6pYgko4ixYEiNeWMzEpGyfMmWeM1fJsSq
SsjXOypZIbI/SbU6AQcGks5Bw4rk6t2PzTJxEJeaHwpK24az3JpoSJ1FxRLU/wQx
S1mTNE1rs+d/XKZWjZ7rKdHEOG4pvcPpQ3KcjOn3spT85Tcu9QvioVr8sgTdBGPo
PFiWdob9kWzrG5UOHUWz2W07qpf51Khuvi3ez9wwPwKlFhJFPadeTT9uZDzYrK4j
S8Cxw9K7a9FAxspE44dRg2aZViEaC+SpNPVQsk46u7Vf7z8sabXmPkkgOhD9D27y
vDcqJqUEQKqWnhF/AUMFvnVXpJZCqXQqfWTqMp/9BIB5sh+U0vPtP/3MPGeeyuUu
Hb0zPv06fAH8sHnx22cMaHbqybHwE9s4sgWoNAETSMtX2IOot/wewpbmXuEg6k1j
lQ6oiBUEpNW/cPv5QyGxucYrAxU96QtQckDW+aPejJ3JSnsrccomjQukZ2KA95Aa
+hgfwMZOnBx/dJyefo1yKMusaBGrO8+sg49TR+Jf79Ggob8xvyAixbZo4sdub7hR
4ghqVQcIYkbWlSz6Cm9HYvO799DngPA1C7j4NOnCgVRQeH9BwsIuqpOHRHUadm0F
k0DWj2i8BwlJOh7knU02htCnJ7tN9RH6gbPGVSMlp5xXYCXJQo+Daz5McVUMpsyG
finipJ5b5GIPeBvG9iE0aR13kq9gg4rv7jj+fCHPLXFelV2VYzMuSAbLRjPCs4Ec
mpAiVbH06ND1J8XoKAS/0LofGABOTIam9oKwPm7qOizXhevCR+vewgC2TEDb+bxl
gdc+1QMt1Fg+XreCDl5Np/DO6dYkxhdruJBzMqAjrx2soUdxYLd88zh+pfzl7t7v
CAtFl8aHOVMhealCsg6nHCgTPS1qhLw8AOhr/NibQyEmqj/bmKCh7p0ynRuOw1tX
PdXFt8PuFtkMpcLzi/1yU1GouiKmDJTbG/IeEaOti2T/yMJfmSyxD/wywHRU97Al
ySV/RvhgrLw8AdKAszeCiTyI6xMwzUzahx51YXEzMSS8epQguS4DZlwNhp5Yr2Th
FrMwVfLofI0no04S8xudg575pVqBiHge1oWqY+QOylLvqs8ky6ojPQa3uI+GoIwu
yrH7xDjezDqr0eImqr6z0vcfKkNdcaung10vxUIl9/jg0EbKOCD0d4220jSn1Pmz
IBVMwAhu1BTfaSvWTAi2zdE8WxeAiLPmVnK8Uy6Jwv3IhaIIR5xIhYunNmwkMRg1
2dMT4V+uSrbyu02P1Ym5Y13WX894j2A47BTSo2RiKpB3e80rlFXEnrPNjyNFSm+V
BFpYynTK+XJI1siPtyHz6FoiYlbYY5s3Rgye2zeJmuQo430xy14w0J506ABrnz8L
2HSr/QxQbUZFxU3RLWGWYXEiKJuCSBgneXEazb91ex2+PbSfNVKGEDIVTcxY9QyU
wtWKiyU+TaO1xweN4WozaDBdCUhyVLLtfH8/F31E5wL3OOO2nokUn/3i+rscUt0+
x2a7Ma01AABiBekyU1cRUUuQHR793u8HX/y2uplR1Ov+s7YrfRg40RR0YYzIdPuZ
dhhmGJhwm4WIOe8nYNQjA/qgAHgdsgE+yTno15dw4bz8kFVIXqaBCbWIyBmKqBii
aaOSOPQhl5/QMtvobkb1emjmMfHcE6XY3CydtkU++KqahF4dNmeMbraSQOawQZZW
yUVeCRGPFTVuyNlRAvQsMWlgOpvQvrKjl0FTBevLtMZbcqJf5rdekWpa2VS6oGHE
vmtrftbuWLaW4E8htlSMYF2eDcQdIKJqaJQreh7y49StdhWHyWH8Kg4F2IpkeB+p
MrA00DAnrqU7zR/6LO/IdgaQufnTr18+Azpk6klrmJln0Ww3IgQdb9xfbXn1pAOm
lGTF9Ngtr3WE3IQJssvS1tEIHeGhDC4PHMUG+DGR2QnJgMZAubTeDYPPxS+dkVsz
4UJ6BqX6qn+PU2uDKq18ZCMRRnvScyzhH/jZ3mn16bqJTT9oPaOZAErw3SaRpzwm
FSJTtwSHQXYi4w2euL6nF3mW5n3rCR/ludoFbG7s0h1GSyriQgi9blJ0WBtvOphT
ESGzWjRQXKNylkfhUTkQCFtPi7uI9eYCUXJsPyurxhGh0fTkvsgQrkVAD/uimfJQ
dnLdgrXW4QfETXbEd/6Mf3MxDjTyO9f5krMVFco5gCAClZ4bTglS3Mnyyw8W7EGR
eZIfx9H4ewUDoQ7o79onl1/7ZJrZXJJ9gIbGt257zg9xmpceA6+xAeO0M8K1WvXb
pSxSgv+EVM2+g9n1541BVSH/QGewrHkcjjkrhUkCJQ34uPAchPCb/2ByXXYe/Q5l
AZlD0/Zd2cCkiS6o2M7UV2qv9KZLMq19v/Hcr50EkbcCccQ++fZFjIEXA4pP4utF
1ya3r3U2bEwuViFYhlujRW5GAspIyVD/3ZIiBsiKZe2LxE7XKmRBBGkZ9hqtqsDz
dJa7cMGVLDY1CbArjgplTcaZZTT+C4WSX682HE4JA2XKjF9fnYj7JuNyc2aURti1
mSR+zdiK00goLBqRN7vA9XxphuU5MKe9k6VBhutCp5LyOnFHxLpcpGl1cPFda080
O0ahyElhdH+9HcnSAHBiyPhWZvtfnoNNW+Ch/3gEWUkSIaa1+R7ciXSwKB2CDkvJ
wxpS9wZRBdh5GLliZVbPWS4MrE9ko3TEtz6p+p2NCpPwb9As6mV32EaNHpCs5xe4
RAVVf7x+ccIUpwDsEw30avkQF7Mi2z9S6hjHooeskU0eOzKzyFHTotRCY3SOI/bq
AYQ46vHMmtJV+aMen2S5/MWfPCv8JJK2NCsr5IEfkvQqgv5TI9fQDXsyqKVGDQQ6
C497Js/q1IQBZFosxK/Nq6weKGj5aBrU6GBAUYIYfO7ETnhThSIlHitVbkdBwLfk
LKUhCZ33Tb06V3ULq2rM+JgAwTVU75mUszWXmlmrUL/lRPvLYYINRMVFdgWdx58V
yfrUtaSXwGEnP9UV+eTLH3Q+llGOHq/mD13qoqBFYN/PGbmjz0DvzDvQFpLJFaH8
xHnFbn+p+143444kUED/ZNFkKav1B2V7g2wIShegPrv4eBiGwkBYCO02cGLsds3Y
B7rjg3jSL4rGmvsjjru4v2xlhftUGPdbiGocZxqdUjSB3Un3Gb2kleNGMXrbTkye
pEtJcNWXlmqOJqotpao/S8p8ziJZsMUH07xtSqZmu60e161b491GtZmODcdqKg5l
r2y9FUjWcnkMpbRlJAxZaea6WyRcWba0FAyCRUDUbnJihDi+kl5dgpeFcLw1lysM
UTwXxwR2DMXhySQPjyOltM955cXggRVt+GKV3DS2D5DB9Ds+rysL9oMLaeAZGU33
Tcs99JrRid7/RrIgOCNGya4pZncUhQjwcNPM1mxefe7fSn5qErA87CLS0Vmva+nI
8BvZlOBVRkoVoHH0O9dA1A0WeKlmYORqUkkNFyuBaIm6tYLIbBYXhdlXQquKhLki
e8HYWDAc2U8bT24sF2VrNn5GK9fMQ7BFIyooHzhWF32/0vYVyYi1nGwbK4VPLgl8
Nv5pmjRFhcZHOUg8a9XPNU/PVSjPWkb+e+xLvS7zLOyvEzEazYPtMQWsFL4Xp2Qv
jLykmugAg+hcL4Sc8+v9lAhA+MY+eSSICPYA7KjdDbjerUERwQE/2fDIJji3DkrO
zjIRzQHVmxFBrIf93+zb/GzS3CSUNT0uWihNlT/E6RJB0dQVTqUjTkcLnIavQ+ze
GA6U7MIzSWask0LCOAQ8DuuFP62qmVEuSlC00SRE0S040mUwSdiTk79a5NVxUs2T
n0DNxQwi80qhEiGw2h9wCFA1wZpWZVlcEK0Bvf4dM0wkk2Ggdx0hZYVPi6E8wzol
ohoK/yAf59hTWszuUgPL5zarQGnwna/aDjbOiPrvdSQO6XYnJ+7pU2RxC4pggXCu
Sqz4wMyre6m2DEHh751xJj2RE4HfqmQ5ZtDDNElkna0sGWfcmrodmzhjdpYgUdz8
Mymb/hhpCV/W2Yx9pH5Trc08o4guRQPviGSuy6PI/XJC/rkquBQbETqQVgFiP1Pr
yxy9+hY6/Gk/KnyrxkWFgBYTbETmCpflQfJMZO5k7DW1GAvZkkojUk69fgWttsCx
EfnBEdBZwZbtB9cLainGZK7xyCXEiPwz1qZw1jpQCUW6c9AKz6uRbOBqY+1PkJ3B
soRB/QXTUwyW/0h5miXqDGndejdZ5nePj8HScki9R9/lCgbwBkcap9yH4ycO+7J/
MgJv611wVa3i+bT2sFg+y80x7vC0xNmHFePSBN8zX4/+gfMBgh9Y39m4rd9o8p52
ZkX1m7hMpE5wSRUjTYdhZg1p9dhRgydQV/clkOaXzTGMMTLaNmAwk6SvlgQbd1j0
vU4IH7oJa32ib/SoLqW/1HvxEdy8szYmW+DhI2ErC26G/Joub0vBCwWOZvKLrIe8
E7peUWoxlGD0P8FMh4/PbQ==
`protect END_PROTECTED
