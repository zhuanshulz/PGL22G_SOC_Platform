`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f+jSL8jxRZqIw5H6mbQgMEbJIHKk2ZdnbR83TTu6IdbMtfQt/iZwtPVLUHKUkqkp
5ehGKuHgGA+/cpXr3Ra6+5GNfzv11LaAHkDT6BeoyiYD0Qhk4Qw6pWJxuLNK7abH
gBmDAqxWT+CHIF6OjW4DWWdTQxHy/vgklqvSTKjkcCkT4f8Y3h87o3cIzRZOkdsQ
a6yCuTpmABIhQILdND4hyf2Ta/BGDv2Z4CMgyd/u6zxWIjAdX/aBMQQG/0/saRlr
OjNlXHLb44QxuzBxLWiAmZZFgUXULO5/Q51cDLZ1fnZIotQnrm48bLrhg8BbGkye
NLNJ2SJUnMg98VhQW+3m6t/InyHkSAs3GDhqgpfPQqqgLKBqCpBwqgCl7VCAHIR+
4jf28zvXeUgRFWDShg56kHmNRUZ76FMhkbu7RPcVIgL71cf6FukUK9x4HrhB8OWe
KneNYXCdiuHI9VtmDUaIlWgCNi/IKUPYXs/y7wlvMU2aF2NZ/Fw+iG7v/RpluBLk
00WBkkw6vOOaiiqYrLvP69+9j2L6NxhOZs6r8nk1DdmLUG0rWZ461PqGHJywQujh
u70ci8kNU0TSrwE1ChtzFf5cxsb3QMcbs7sBPtL2aVtTSwQb9f04QCiymUj6EG+r
hW72+V/LqpL1YwmhD7bGq+niQj7KOZwOn3+Q3A+MGOCGjMBRHsXUz/880W4twtAd
0pawqVw7EYwj1Dd2f/wCfraNM8HR7MEri8GNtfbq0oWFHdNt1ljmmEi3TP82jIc6
NdDuiMcIhgDHrNnKIBHjNaZseWpcj2JZ6f4i6R97hMmulVzRomUDZvRvjLYLbwsq
PLS7ZB5xzATToXmnr6qHoRmSIssaJpmYGTteGHLKTkYMRXrMTJUdSpRnY2NZPr8o
90CeRlpTgszDPCHBY4XNA3v6hPC726+DJt5FC/k5cjl0cwY+pZ+cRG8DcyHkX5gV
M4miJqbtFNI6LRDHVmweGYOHxYwsgUpjxvSl7Uw71JI1D2EmZPgEeKT214EGndk+
BGqVVZHprMlDcel0j8AvC2sC/L8ME+GaHEaF++dPbCiGUJBLjVMJH5QQXKywMaSe
dZo7WpcBrYrN0y/nLaJ/zlD2a+ptTg4VhlJv8xbHZNPc96Oy0X98h7FxK5JBqQ4X
9HZlPryJAJIHsbJRGXQOQvowYaLXW+pkvczscZZHKBwPiek0DRnoWFCtLaYiSCZ0
oadt1BMmpcVNhEnPtQTvNvyppPPDW4kML/nVkSb3ouwC8553A9BHGxqEZli8f6M7
P1C6QD+hVqIxCn8oLwCb+/L3zcfZWdiFfQWn6oXBcqA2DHqfSkF1aO5nYdLK/BJ8
XnTI+pkYVFrw2VuZ2lsZ3QfH7pbaNCqAaP5SljJ73Cz2r2sijEIl0M0OfviHe8a8
ljVAecQUVERKSxijkTofq7WBWHAm0qVDFaLkn9YVolfhjYxoSVPf20CoXoqHi52t
aeYrZ7xwR5QGkTYXBvusN34U4DxBVH3YaTyewad6WuD0k4JuITUYDwmCC9bVTqW3
HcPmAuy6QUvYk3Mopp4OgyCfHuliQbvlzHA4H4pUwpTdNeWAnLmcxjRenC3aHsz1
y1UzSHwPiF6q1oRFKzsxr1Cmocgq1IwUPr0Mwuat/raUdh0GWMJX1EzBSYA+EuVS
sGsJwIvuOAI0O+7X0D3ZOe3UfLxoAV1u/sId9nGJZM3uexhD/nBeLqAS5fTI/YYH
mcVn1c+idB1nCQhz9LGFTycyO3QgOYBuIIevmxLEl22CEHFTUtrKW+7QHcRy1Wvp
ccrmS/odIuVC0fdmnndS58aBlXZS2M9zXdA69/KxT9ec9pubp8St9mES/vGJ84+Z
uL0I58IZCMzFpB4MnZc9N084dLBA1l9UzcpRuUng7+V+kHr0znSU99bMmuevcSum
9Itn8oyRaZJdqVrG+e4Rao3EDI3j3Ltwn/ZkJqF+gaUWryPyj5qv+NhXJscHlgAb
g3dZaSCYXiZ6FOCKl5Z2Ua+mC3uGvGgZLBQpOz99sbNPnasLt1/j/Vf1vaQdprq/
lIjsPBLMqc446kgLRLzh9GaVmJ767SH0cA793m1rZvETVfY50eHd0aXACy2lSH7u
lavdHOkgqGhbsQCGXCXrTKC0NFPYNftBN4Xw0GEnj9zur4ZERvwp1diMcNyFKYk9
Gn4iXUqPv56U1VZa9tiVmuratT2C16GYsUypUaeLumm07k0NHhrB94yjw/af375D
WfKXm5ZVbRYbKdY4cZVlu8DNwMMlIwErMwo7jVhGyiLd8I5XxaszvAtV1+cuoKuk
c4RiCddUN6hfzPfIpiWl1AscE4tDITdacUKZ4gnXE6Q4Gi1NJMii97ryMXtarrEW
HKoQEva2nBZBwk/I/deTYO+PUwSiFykdzMqkmSYE9V0lTm2cftcOOpPkE1xETQPg
CCTOMg1xfUknIxz8ZeLe5ncCLurLyIZpN/UCG9kndPb5rAOjl8aGVU8ACmBCDIcM
C5qyzloBz3QRimtkE/L0gWLr3aD0FKZ1uvZ9k1+cjaclVYjEUcRu1ZkVamQY1yyp
3X99AaI1iBqFojTIHLzRV5cq+EEdjNeZkZ7KJbuchqm1sOxdUJRbHmBczNezhrm6
Be4cAwSi0Xf78eMzKyuSC58t2mGOqhGx+ZKtCwKTv9LLgJaBANrTaR/ihsZ5ZxqB
+WgQz19xHVTkBEF+Z4qBmy2lsjyV9yeUr158SD7vQ7S/aQ8g7hE/8I+wc2ELFSeG
FTyNXmGN7jawqPdos3beJ3xUpVbuqyuRE1LbjteC7cORyo4zG4fbBeC5XpW8MuvD
bV6fJI6pcRs2tY7waocNQfnIph3aFkgMZ3lP3wMWpLiIrhttjTEWfl3Dv9YkjaHX
8Lx5/TvvoUYKU7G95mJGU6TS0UJjuAv1dM8EoYa/4TuwB3nIpdHBdfm+WG8zAgo2
UH0of/nGZQN7OwpoSBbjaA+sJHBL3Hp0VPqs9tHOkjCy5wIOh3hMHeJRVJpOUgju
FwUf4TzFI7iiPxNiuE8agQskvnOsfC3QaVa714RQJ/vD0AWFOUXZmLKqoYZSEJKY
DZa0Qqcfm1DerwL4uB6H3BaqXFtdS9EpHKow71dYM/9uK0v85HoKPRHi9QlEnwjM
g1RrIUlZqqP6egYyiw0E3P6/vPApM54DCvQ0LIKPuuieMxt8HOL/42pp6gX1YG7C
goCKV3GNgNJrRl2WIgYvtz7BJf4+aHwtASlsHDuu8TIF8+OnlCbGadRNjRVQve+v
`protect END_PROTECTED
