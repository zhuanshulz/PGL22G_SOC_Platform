`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1A64SJlEtDQCXwdvaMq0ylDArKGrVUKQTIMvpCK8tT7O+ugHf6GAyhHbUJKzISL2
HP4YXnSFBrGPIjqL1rOX8oWPny2pk+KQ9r+0bvwT8XT7JG1U69EkBdcx50nAKwmm
EGV5LzFokf4Vrt+Tg8HCmRf/lHvQkMbX6VVgFOmA1uf/Vq7Thbop9Y7xyAZFrCws
7NqvRZoj7jaI8rpSEzfkQKG0gVAm1J8ntjKxmyvehW21BjGdm5ZkERMTRSG87JM1
oOIEcTxNebVNUSnJtxeUVgOzEmm1O4vaPfVHBT9KY1jsaWpzhTNWZ+j6PoV3FK3p
mW3+JVer1KwvrxcdVokfjpP7FLiK54GAaLtAZFc3m4EsSFZRYHoG0bf/qE1oOJWe
/cg3n72d0OOhHHvRJJQeFSBC86MsHZY1kHe08HLi0hxN6y+E7SEsvCqCKqRCj0sV
/eP5OsWuOONWKfS6IaT/C9AGkMMFkQnnI2twAMPcN+NjCHPDm0w8Hv1ACKOD90r0
4tcUT4lxbup9UZ7AJlL5wii+7beu1nUCS8qu4jGIOkEks0PMF4JKphBW6i7WPjg9
lrrL0yuA6DpKcoXzhEgmUAsSEOlOx8JciXOSPkOLwG5NZVn4Vie6ySV2bM05TyBF
C8ds0HJ+0CGHG62lH8LHBw84TmBz/3UpGpSi6CnKRcXIbsEhnxPG2HmTDKSBP0GA
eyYN0L2elq8OVvx0qAgVZZn6R3SD9F+kFA/5QP1Otkfwx9mWmjyOJLPapaonudhV
nvXlYnQl1vG8HmPK9hc2CKUzX2gTITMcz1OI06sQOCYH25bJWMFHUYhxagOHr9HU
3GT2XRn/n6cxuBZYbZLkbJr4tHKew3FM5H3sSkK/46GhPCFrO/P+/GAyz19fHHzB
OPEmZLyXSofwDle/5A+dkgnC1MiD/dugFTtE2fr4dY7tMjC33JDHF6NJ8o26oPro
svDLAaMAxTcAXTpOmRgowdI50uLmww4blhauOW8aw74tMuwLNLs+0Ns6DU5xJPkT
WD5pk+qChZCQsuGb1zS0vSThbj6++6dVu412tKgUd4wXpDSg/Hk+WjhgyCYUg9rP
qZhQ7xaE7o5YC1YMw6jutcP9ivKOs1xhNeUfBEPZLGxM8cJ8Xov6buXrG2FHVvBy
dpjTS8mefKkdxB8dhld8TnOFPUKfTNvDXUx0+1Di7ZPwBMUl0+zETb71yvD7VoH6
nx8LH6y+jIr2arbZfB78tJ5F3ZAcZt5uAg3WSYrNaqyaRQ3efZxxkzuq/Gh+WrNp
CdB84uF6s3sj2HkrkxjhP2rdsOxdqBFoyAzIdBY3qiGwlSOWh7OowvrMm0Mya95M
7GSKG7f6etEyrF6JRDuIeY9tsn43Vcdg7Oc2zDmb7C+J5JTgsZpjwW0zh+VCEtjH
lGu5BCA0PgYixmlQtJ3dSV8NYB115eRHe+yrjGfNpn9Tv51Piqh+FSMORNogcIV6
lrbe8Vm+chlVujqORc3KF456jWPAjjtil+7PonNWm1HTr2eIHCETZXir84N+iUuz
pRYXMPOE0YV7uoll5OCT2Ez2gxC664iOj3LZESiZnIi1UULbcWKJA7+tmT1S7Bau
Dkd7ukz0JD4UF5hQng3OGlOk6MKWhvh+kZ1pHTEAI7jb8VAR9dtQ282m2xdsLwHb
hwURgsXeP9Q7reZhlrwnajzUIRJjNYq8L8m6AmcJQQMFaSdm9OMZXalot13wl7vi
GPrccvyJ3S3miFLcrUOv2UJljwZs8XmIy72FX1I2Dul8aP+ue3tLmwT5LnuRnuG8
/yISdfILplhhMrkawxWNTbzTGHWRvpYd9CaVJfQlnPtlsbqnBnTMN1Ht2nRcGGpP
qEZjX4vQpi6pDRb0qDg8HJg7CUsOPdroIBsF26jtZLIutW55pmue7GjFUYmBJoOB
uSo8JE1nr1XepKELBbqh+o+HVb/F7fvaxMWTLn8RQJvCu0AAlWHvuuUqVsmvfy+/
XLZuuCKBfPIJmPXhQOXFXOZH8l392/TaJlwTDCURaMI3K6j7vbAtAR+VzQ9Duvde
JD37otH2ihhS4o69Esc9chEk6eSSNXSF3onBDXfyu7JzoSnbCOTLwGzczk4Zk9dz
xZHB/wisyMLZ+m3W94RfYSGvNPA31fuCpOVZPl0kxDeUP2e1uxt5y462+NFgs5gs
nRlLZTOp5I+Wplog+srE4Ugcf8RILkJY2SUkdodewDXIG5AoBg0Bt+xVLcfzvOwZ
vCrLYkQIXC2LM2I7g+tVo/GO5GVd2LqO49HUmSU3kUxg5JzmGvS/wSBXJzD5Yfel
HPKddzqWImXUWtihVD31PoJEncJS2x9Ykhk6wliRm/xayuI8lEXTrqzpDO2J+TSg
PWI7e9ok9rEabnNR1DwA6uui0P/3N0xwKoKWhVSKhs09g4S88VFZtCZGzZrHB5++
mQQ6HqGsd1NkzFV1Eu6scnRLlzHGBdplQ/lSn1+HgYrsr/UY1BpuA8APADpUvSuM
DTjZnKVDIxICrKzy/IhLwt80uY7KzdK/e5mbxTK2BbE=
`protect END_PROTECTED
