`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXsNtQ1wJKCjv+qqCfAjFimuPBDXgV9d/2rgFQraIBPAyeI2FoTxq/gk9EtwKw5F
FM2pg3Ij/XOaJi0naWfq7GkeqJ7sSE3dkRiludxJxVngrtwvc1K3u5IofuCHiDDz
5YLnL9syp/Ju52/4SxvktJ/fGs3RFZvRRrsewMvzcMo62/icOC/HeyTAjWRiU4zn
wMyAV7Dl8ME9dIAtYYqXEbXS7RoQZcBp4dEq6+r2g64o3pU/S7scZ6N/Zr5mjsMG
QrBAy/163NRwxSQ44aInrJCal6+UPJKCMFW8ME9VC+mfY33KN9HvNWrO3o5mUREM
3guvvBYEAxHltqcwfyj8X22ecfqUbpXdnVs1SY0XpAB53l5aOlSnhUKbzcfunDou
vw7QdzCrtNmGFIyYNiJbdGVUO+phPrlDHBymcQ979pzeC7MV8gSRz+5GM0jOc80H
Lu+gQ1i1zy6MuyMG8DpZzc5WLc/1y2qjE2CAa5CSi4dIUQS2nyO20v63QMa7Rxna
hq/jtrA9u45WQUjEiaxfu08dREkSh+J0Z5LAz2/+5oUE6MRf3LGJk85g/h17bw1T
Uv1qBWIaWk2kURXQ689CS+qsqElHB3i2uu3fPxrBxNzvqAMU5K9jyqn5TguYuENF
5kDjg3jcBNaPBfF7LqiM6T0L9+DYpVGIcqdS0a3cOjzYtYr/C/ByX7p6+CEzE/mz
b+fzGVR4BQ53fFP35e1O7/H8829fTU1QJf31r5B6LDOS9Gv6IAOsUBoDsGdIU3jC
OioV2iQWkPf/Nt6r/4a4QCdvcdJRQ/Lb2Hl7lHlQuZIb1Tu+2p91RaEwHAjm1r+n
JXTeSsbyZ2R2bmA6av9Y8vUVViMNQoIFfYM7sRc45o1oBfXD8I6jgOx2qQk7S+3s
Q2TZAtJGkqrNFg+MY6WYSr661hkoimprXfCWfVqttxco2o0CH2uj6CwvhaHvgrRu
eGK5/BGpc3Q3nljnIm/nvDiX4Yt+M7ngfyqoCDs/O8OaiiE9ablanxWPLKfI2wxO
EtgETPZgROrkC2I5obWF+8xcH0G46FF8xENDaoCqlq6qNLVV5fhDLUuQzK7D619Y
m3rI/Oe7IiqYcgc1qcHCqcPlpf4C9oTDau1bqYsKul/seD/+rjL3VTmNFY6dzHdL
RWZ0xX6Kp9ml0H+RRUnCu9OJnI63Cs356KhUhfk1V0Djq/nKO57+hbEYw7NTwEob
5/CR+3r7z4KwvIH1UYskfO8UYFaOE6PaFGUM+YTdnXF5wPjKH2FXWHd8R5bgPYwh
M8Tu0ITi80n7zT/v/skRcA==
`protect END_PROTECTED
