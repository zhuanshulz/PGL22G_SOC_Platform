`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B0gM3wgh7M91LrLlSNXlPq5+lGzT1anvAme8gERzZZSaAAds/AnB8G81dLCwvMz7
7Jwu/dy+JHv/KJ2tYPU1o+pBR3/y5cBbDvNcaoa9Cb1tkeHcjYQgHIrVOildxoe0
Y0i/SbAukRjdoUGB3K5upD5uWy/NjBEhf4TW5zClGOmo7IoBYDeFcb3TA3fL0mrq
7LcTL1IoGfgmERJNap/oa3O328Y7VfbNPRU0KXstlFyx5x+g7QNb+0DZe09krLdR
i0tBfXlRpnBTKORffLjelcdw4hwpiYUDUQUHZZmi0+lHtIE0WzID+LmZwef3apKj
Dnwgn62GfRBt9uzFk86crw==
`protect END_PROTECTED
