`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cK1PRG1D4f4rx3o8BmbSviFxzLPQbGMjGMZ2hSw0qnjjBiVe/yx/HkfHAWjENGXH
kSSGOHsGjvYXXESpn7djwO6a+D0DXUijDBe3o41n3l3nIVOFS05R9KG7F6HoniIG
48HQREj8nujMVYwA/zt9T+2B3390jkqyz/26YBsMMyPeOYCxIt3gIuGQv5WIQmQ6
04AmJHI4btHd1BzUGdYic8TfFwKaPTrWc8+a76bc9QKAHLXvjx4k7PSOJnQhKlIr
nb2gOluKDNSq3zZUn7jFRIie6PvE+8jVPYhzW/MMO42NumYapoSYsX3M2wRrvFg0
e7Ou6bF/wl1Dnx1Z7iIMc5Is2+69s7+AxbFO4+FqpZQ7HMxv8mVF6BSTpQWiXjdE
mWTOHTWk2ZDIDzJnumUXA2/vVhF9iSmnw9Yt9E9LRrpxtkzcMfnShgAMUA5I3T6I
1C6WZ2ueOZc5vP75pFZsWDiKQWRo6GuSgCYOFCihlIB7dgy+AeM+aRupj1zy+v+u
CI+HDP0sSxgAkPFLFH5i0aa71vUmMqLBIdQ2PXeohArG+0tOL4/Ig2KFeysP8QEs
kJPUzgkevpQA3NAsv1gB4q4uyCps6C2KKfmp7H8xHD2yVBCzry4b1UT+yE9DxO/a
4tq0uNuYsFhUr0rc3e1f2Qn5nluj1YYRmObLbI8tJ8joc9BjIw+uXSU7VIe5mRmX
tQQ6VaoqgszuqwQZFYtbCRPsyXSVs2QS+WeRZzHP+bbgoZmDbgwUjXcGmOOGpkQo
NS6quSqV7m2OC5zmgPwQ/ecsSNoZti2pSTNzuj3EyvvXoVC9Qm7/816m/93pOM2+
VG61gm2PG9ofG2/ZRFWznajlYxuhQLKpCvTDD+vquzqCYj2rWI/8mJkT03L1JPsq
sr7/6mZm8cdRF9vOV+o4uNmx10IcEGpfVwDb5NhmHz6avnIwMnXTwdPUhOD7ayNj
rVkwQzVEooh90HFG563J5wUGF3g8Ng6oF7EnUdUbfTXKMwubplzsu1ETkV1WoXYW
muhJdeEjub/wLBSmYvbVrZCsMtSBQyAp4BCJf1zaVwO1j8HpZjd3dbuVep+1/JQO
+t3XJ3RZjNlAyyJmoh0eZ7/LAjvrdExvfAKqxvwUOsM0xCalXA35EqOWI2SZnrRZ
8wMSM/KiJ4eUn00Cg+zI6PunAzjWeoCFrlQh7+n07Eony5q3QyqTqcTIjo6wxbtL
Vy4wJi28vBDGRfS5NB+R5hF/HKdJXW3b6HSFEwvKlnIoXPoT8mb7TtnIV6/Zalox
aFQbfyCQWm99vrIpu/4JUMYOGXh/xWfNGkKLbxXblybwh07+DLaaX5dnxMwf4ZIC
BM0Ihon/ofyf7DBKySF54F3kQwrCA6R17bjPtvSlRvjj8vtc+TrZYpx/AlbqKrmN
vkIjadFwIl0p/poif2soztDABfGt0vStjKGRcltv0JmkZnsjtcuxVVoAZ7MPbauk
uYvOcWX0U8g/SMBjX7eUVZizpsBxK9Eb+YCGu1msSlzbBEH73AT/RTd0rARWLyLs
uMYyJctEco3nnM3KuP/+FejPvSTvLnrVzBo9J65s/180U2O/EzlwYV6cH3YBcz8k
nC0VWF/bDFgj8xWkq9s79YETBVdpfhrgnGHH0y7IuFAG/+s3aK4CmI1Dg8C6vYEC
BveL5ar6GyhsbrKwiOIv4mEBJLy5/6hHNd8PJmVlQXguzIvphPKZNPlo5dpk4T2V
MHy5if68anayCV5TKYWsgWRRXBh+eydHjhUUeOb79buIkWjhBWnNDp7f4Wh4qWzz
8muD5HaRcvgZUWXHBES1+MCbktQDElJ1U9JblYFjR8nzoBcGWa0qLmwj3tlIvZnQ
4+2MflCN4WRQyHZpRxbeyN8AFDrIFomAIySa7MbiNjMUu8hfD7e0+s9wfoaHaxys
+nicNDytHWC1mwR8Ro05il9ukbj+O+UW3nzL5QTiunW+Byo1zVhENHhSd279xvxS
7UEfH22FXQi9Pxz/T20rBXiz6LYPqBuKpaQ5/K8pcQUO1ZNQiGWT/AGwjOY8FRRi
XJbxEcGzHwiqtYeN5+YJPeLmjFszQ+Sds3usIysYxvXOeJYDd8hR0fxlVzOz43sR
AWlviQVdzuGYb71t53xfr3odWeDaJFU2WgzmWN0W+aTjqIrmBoP/HpaL2mG5RgWW
bB2KWa9jzxl0sMpVmky90xSTBwWE8qHNW6FtCdpQZcXaaZpUDUhr+GVcoLfzQukK
OUgqkCCjsMoZFeklgUmAk3osp/qsXSSOZnIxqzzoaqIntLRr45pVp34v5mybqv0A
eqN6wTiqbE9CS7YTEJNp2tlzgcft/s7ag0b7EqXQgX9k+bKO4TO+Tt6XRdJCchHj
6mzZAAuqzFcP3kPY4hbeBOwRVGW6x8HRD33kFrXNhZt3VmJFUDG6Hjipjw+GR2h/
7aYZU5mQ0BJdi2KHdo+BmPc7jUUXEwSWgysdUV+Q8KIx6sRtrVc/pzdkcBXBT2bU
3BioNiNTHvu9IpvzQpo4Td6SO9KIcD9E0cnBHPhLHOrMBRTBTTCFZlqeowG2+sX/
8EWux2+MwmJLDcQDW4mMEM1tTbzRhg5FLTXNfvj/iwqOzsS6RjHMcO4uoxhX2Xs5
FHVU8VjogNK1wgW02qE6f+NrBzVqcFaNigrtpUaRmUo72u5L3xibpcEgzOiRv4nU
t4B9TabnsBAbzW4DwDO2X+ijB5rGzm8yvFAgh9MmAUVipSjZI1JFDQjQx+u1PqXg
ijSe5R0HridKZUptkj3u8QjmZkLxwX9XGBywBM3U5kLIFfUFLxhyFzEA+bxOkJRR
rNF+DuHpvhrbG59SRlEMfosWsfUolHLfZIUCMJracbt0srWOaWXx5+W7JfGygkVB
EhJ6wuQ39b8xQcPah0NSLXawo2o1d5Zxdy8wiVuwxyVGSut6VvmHV5QDDCzmFnwr
+QJbU9PwuENBC3SFBR2lmxviJi4owqGv2irQB0gts3R025KdrMiSG3AbSW8/kW9R
7S4+sh7TEoELP81GOXQUPMwekTqnW1j1Ulx+MOSTn6cePKKqG2tyel2IYxjhW7iK
vymbZfa2cq1KY8+KhNj43eQ0zBHsRgKJeA6Q6qdTWVwZUPIFXyHVen8Tpf2VhQyQ
kjbrJiCvMZ5UHFc5nSXfHP53Lee3bvQEW0JlzZUqbily7lpSjj0n2JRIcU4ef+D0
dW1srR9bUDkzDpa4K9VEvCVv97r5BVXCnjgBrD5K8P2+wSx7D9dNffuuqR2ePx3N
3oDf/8V6sycnVVCdALcrXwH3Bpa7oXyYVu3AjTu7NbJCVr6904JrguklnsIs56sb
AOo3tFpQ83vXJ9CQpxp/BubF/GLb+mc0hiUyscIsVAoxha2ene61UtrLGfOOwdtD
rK+H0NrPg2PoD6sTuvRR1TFaZB+z/laUSKgW6Sg4AZbTtt2B83yxDt0J8Gn6JWbI
35ixQcD0ehu9JBFe+R8EthJ/FqRcKBWprLfJvDMHSgDqyaQge5X1ljoh+A3f28up
YvQPA4fBJeWaj294v5mBkLjM0ubXEKmHVOUHwVSXubFlnfsozD/wonLrwdBoID2X
SYGXZKPJ0ayrMeJhpka7V6U3vnPGcCpxkUFKxEFmvFN/8XWtGfRSWMb5bpoO4bgC
92ITnYctjHpq/EWuGpzbiwtRIMKYvrl6L8UB6NIRAPvklyrDg0FFnCgrODbtYrjB
MW4tUyz+9MBMLFTZ/d1ZrtpnLerUb5G2d9QIqHPSo6atc+r6hBrFRMCCYOBNmAa6
kD9rLHtPyEaKmkT5BQrgceDXacm3lHPWUloXMFToL25VjWJIEFwNSQah9HnGgt0I
n+/HRt5BdLq9UwTeb3ocbIU9dkgSdpxjvxfuQrMwZt81QxVeaHrTXY+lIgc8jtyP
gqrWqv7luZRjYeq5gDRcUbkqLX3CeKhe4Q9UMSnppt7Op5PDhV7u2ulj7KoyT0mY
2/XE9w7+Z8SsYoq/NsSzhnTxQyuID721WwMB4nj7wqWhycnpDTI9xT2mhwkPIE9i
ZPI7Yux5tYSJ0oIHtGMTeLoSZZ7j9PrzBcuI9438N5pNqWYPtgNVYjn0LWllOCVG
X3L+QOnDAeUuiHQpHjNErgirm/zfGiu1n7pVSQK2D9BDJED89wZM/jnK4IuhLZDm
u2dC3YW71FunvSOx8duQN7W7zgi0GXq8JNsCWhEoGM0xHFmogLPDAntsp5dXzg6W
22PnckGz0s71DPqDlKzuyQOn+cSaIRxt5Im9HSQTr57lDYktF9eTrnb/RpCHSyxP
/luPgghw/ybk9OCUF11oFf0DNCbT6FRwXs+0OKRrdKSpTtU5Vlzke5vsSEplCOoe
YQ6oI2Nsvvkr645KjJAWscr7q3nXNwimsrLc0Yqq2kUVDA2+bzxZIp1MlsBdtTec
DgHO/BlMvaAFkDMsLHw+2QomEGwJMDz5hrrTcGZ8rzsPScQTZDcnTpIZKEUFhn64
bC8rZCc00dvo5yAfIVfGIW9Vj1Q+gPPUiGiglfYbkJEFA8ABJcTAD+cSh7liTec4
cyETwTdulUNdjfWfe9mDkyu7VJP8/4SpiuyG6wlScLlntMeFkyOpsmAA2UJFI3vN
6wnWpZ5IuL1w7TzcV1kg8b1oFMNNjjnUTg59Mn5e26wkfpDdaTCRT2Js5WpWnDqe
2FcuuG4p+ztm6mRwknmgj7gs+W0xwR62LZxzoWdoLiOcozWUwnlPRf35xPGeAv1H
`protect END_PROTECTED
