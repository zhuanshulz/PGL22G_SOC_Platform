`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0UdioH6R5AuXc9bjKFKJhXZ/I5pFtSB7FYx7YF3lImhu+95ZiaEeS0fj0FZ5A76w
JpD5dNikmu+FlUGgEcWctNVEHAhm+PB+wtnJz2Xbm71ayMZ4vcDF1L6BvjLwgvCh
4rV5qhhKLTGM1+3R7kxmNeCCyDdaBABZpzALoClZEquCXv2QFd8RFIkhDkTx1KbC
abth/rdiZHhlFDkCIZbH+Y5vyzJO0kuYTGumVcKWQDGnlYu+ENUdjmtzUi9KZ/9n
NdOmEyIpJLv4+MUcb8ls7X5ecmGtN6O0patToTCRIKtuvCQcv9Tehm4elOHEKwU2
64L0M1+6WOT1mbYkkdm3cmPDG6sMAKw5+GlLiQA8aPy9FafoFBHTQWmF9lE+MwRp
6xeIvtpkiNypED3JcHg4yzGaR85KxR3tWM/KATrsGmvgjGoZZ4zQlvSr5l8o2XMG
WTVNoRv3yo8uHsijnR2/JRO1SbOiNUII8BwGXWsff+lQ6pOqDWr1sALmkUIq5d5O
9C9vWSOfSjOi4jl3fT+wSyPi+4ci4UZAQuRk0h/2Zj50XiJ7BfXvataIslhw2zi9
YfuopwtQMTvESR/N1poEAnkgzqY1gf5yFA0G7pR0Tj6jqOHQYbwj7aMoZWmlOaJK
v0rpQSmXan9XBS5WhF73LOztoTpARisEbGSJMKZJv6MaSQwIVFWsBZeCDFGKkKgG
qcuhHpqnsb9YY/1x9l4qsXYbE254RYcSJT9tK/QMoNzS6v3CtzIpButTIIFHoAve
BghPN+iT4GhLRJjPgyTqrlFNLukPLBP4csylYb+SAV7bR2+erw/GvdB9aIUKvgJT
1Ge7HFX4LppQXAely3FsFVz9ghqxweEsXazh7v6vDi5yihw3g23z1pylcqiFl6XG
nq+MoY44XnLomba5zAQyjm3JDKU6nOMgOwxwsrSV3KaxKBLUwvKxxloONosLVg7e
whgNt3yZX+MXa96hv9Dc8+ziFS2Lh+gMVXBih3UTdEyX+qUU7TntMmPyHakvxJ1e
Dbdxp3WsQiRbF9sI0/385wbLB41VbBA6jn3GV9rRX6bxOC7wGncpXLiqUMfJHrLM
ydFqsTFJFJUgYHy+jt2vVA7JUcwPl3oo1IWFzoP7weYJqHYOS9AV7fbvd8yF2y3B
Y1z7HL/bkZBmCI8nnFwFsaYLtL2f5qmhSlFJTj8j5HJ00xR9f9Ft8axutYYBzt4V
1HFIXo5R0Jnrxmkf71GtlUwjXbdgGoaW2NanIsrS16kdgqddxtdXOaQksus7Cxxb
Q0eVE5SQ2+/U6r3GnakVWbcIEIaduN041O3zjVPf84JqdtqOO6Fc2oxfo2Z7UtvK
eoklWmJn1h1CS1ppKlHa4Et+M5xKVGM8XMH2BZ03wj38qHXFd+pNFUaZeoOA6BqH
Z+Hu8efaFp4PPa+Hsd3XlAIsnOP6h3YyqYZk7TFmAdgCXlNmLeQXCB8mHamAN8QY
nmYA5kNkl9G3S0fMk9vGcIiEPZWSa4Z/d8CE5sj2QJV3dzYwXzyLqo0J/shIU8NO
eGjcxT4rR+HKejMB+ugOjXFe7XbJL8XAROkPeY9mNZKujxbjafkD0EC8GDqqvtuC
iBuKXCsU/7diNBdUQGlQ3eV848sZANun5PLOZB/anCVXHsAGDx4k8IO6pU5rxNtd
bANZcGoXOhtHZM1/CvY4JuzuQ0dblae5+pud76Ybm8MpCcr8xtYqnitH629lwuVC
SsOSVwY/KTFoYRtZ1v7eJvkOS22pKkcKAddWw9huDlkif5Ai3BZu1HMNk7mmW1TS
CvG52fIDCm9eTSEE4PDyDGWSTTCBETqnL4zkP9+JNKVffGylZ+eFg6hni++plbyQ
fBoCUSD6q1Xiy/VgOZr3BewFC4tt6Kel7+zcL6ly7KWmhPaVPqvQfxpT6BOUv8BP
BSo9WcU6WHhm2rBBP5E47cbczH9GAIp2l/iRKNbY+PyHGfzJ1s3qOxq6h0Y+P1NR
L3DsqOusNDhklJBvtykeXCCqtidrTY2elJigx3uxqPUzkjoTOmInhU1lTH47BkHf
X28E3rMChZtz1IX1rJ51dtE/VaDNxGSY5KVQZAYaIQmKGoqUBpg2rdwMXyfBGk/G
Y9+uuBPow5/5vDxE3XHDFe9nFy15jD5uYOgMOO3pYS7Yrkeu+K/1jv1dpbJkF92A
kI/s+wsDr9RSVFtGxPLDHbQugfec188+eZ9G+ZFWay/sdPYgBvkMan9Dq0OvvZL9
WyBX2jGEKcxUB/dlUPz4devWgAr9ITN0p5dnBZLnaA2ysorNf9IqokHd0h35aR+x
WCKz6d9gVRb0leBVG2fKCq9M6sMx+7fdYOEGRhqPQzyWA5vqLiUR2iZkTFj0K+ET
M2JI7c9mjD+KxWjB9rsAk3KQfSQPEqUG2oGXCi0eY9k0RF/Z1bfgESPjH7bd54LF
cSfDDH/gFvvH1NG8HnYxmaQkfzjysVlBuu/YDXN7Dx6XkMlqtK5ul7yeBb3wd2dg
To/PjU5dO0x5gOE2w69nOkkC/zvYbI0QHdse+hYXTRETnBl1qqjaCah9j7ktZLKt
VQmUDVf5s22tFS8HQtU9OoW+OGrf8xsIbCZPtVIBXoTU5xRPVtMQJpiqV/EZHVz7
vbCBshXVyE2xls1sJFIwSQ3Mhq3/Q+hEWQ90IkHjzksgzMtYX37sJkT6mhtKSRZ6
WaLQScshRlGSvnSi9g0EgYJv2Uxc7OuVLF6MF/oenwYIZi9/FDHLBjEBk/Qi5EYu
vJvyAHlYBOeAy5md3HWOHF/+4xCv9IT+CVccI9LeEONCziWSjPfYS9zITCTvnmxa
2rOsf9r1CBGbRzm46f4f70H0drhQpAzyT29AlqOd2AI+v+7nRKJCRB5aeuAjTFF2
BducX55trPzZy7CDjmDHejdmmj94FIzlU7GvgrFUiXGewhMuvVoxW5+I9Cgh9cZY
xVCkPYMVfEwBE7xVt5T62mzeCabVPrB9l2kMr9V3oPlQ/Oo8d4fc8yEDumAjPN5R
+vxPqS5sDui2kwuHkS+K9sPEXRtLoGfwxt5FfhOUJ0+j4XKJyA9crAbLF18b/K6k
YT64ut2mebFersabDBxlJtSwja+CCvzhyMzsBfsWV5n1c2VZ2CObioQpTrgr0HhE
Sac2CicHth/1I8iEvm7kqlvSjo5yVyHQd2UCg/yTFdFWm3R0loa8Q9cCygMuQMeW
xUjQYNmfzxxC6mwSzGUwAPqEfTL1JC8jMaPVKbw27kHF+fmBPyWkbSr//aAez41K
RdS7fPGCUK5RRL8Sgudkxv6oZjxPMMQqD7HZxLTs8845H+FbsZmrh7cNhjTNMG1X
IAsS5inJrADud6iTAiyzuvNzPE9RHD96kTp/wyRQ5NDZCbmbmKbtS41VGqSPTUIC
tEqrp0BT8wBmW1cwgIvayK3j4u3sjY28ZbspGbsLOypgTrkdrVFCAvSVpuwEmUAB
qsHuzkZdHyn2vb/Uw4ru3vww9Zos1i0Efieyrjoq6SBLZqw67qdMpYBtxZyufFXZ
4KvS/yQmVuBcg+8Vyxx3r8WIOGhidNqJb3KYhdVOuf8=
`protect END_PROTECTED
