`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pibEit7hcDAC70NcNxPH44tYUr7ZM81D23fQDJPV3mSzHRfT7kzFxcv2vBJXvELg
9pAU5ePOVictQEj3GZrWIzF3lbd4htyG1335uxa6ODaw9pCK2LCOixv6Zuup3ADk
1g1GwW9qGRuqfgszcWKzTnclXiyDNvX8Yv8/qy8nf2n3W0I3dHEvOnyeutIHl5/m
UO/rskIWKC0mUrJRhRDn/dITaJTbhILYs6g+DYyOCmvPlEipcxN/w24FN7vB13fo
7YwJFpVpXUctfXhL7lbgpeYpKFvtk8D+qp4It9cH1PAe7+njjs+K7mo294gXBz7B
bi3De3fuRTA6vJ5dtDJmKdGkxut/ERogni2aHTL+M7FTNeRt8sVqVTHyuEOMOC8a
4M2Hn0bmvrHIoSEVRRgA59TXCeGgR3t6PxwqLElT/Z1tcWJSvaTqMwU7LHPCUXWZ
KPRZ5UKCPtWRt/6VX94UJJfJHdPrDXdz9iJokEapnZ/zNvQOQV9D58MPkt3VHmgV
RENR6uaortOdFcDU6DTRTXUpAosbWO8ypDOmOXy8ImLkVijtnjM+BesAGyS3r6Y3
asdho8BD0ohYyEGF/LfOBNrPJBAi/Omg78UJgxR8/PdzDJnLCqfEcF0Olqeu7+cr
v0pDtoVM6/zIivNhATBTP/FXlVPyC8uOeeJM6y7U9t+loqWXjyj7+rR5ugLiRcDW
DcSdhnyy09cyySS5wYpxXBVpqVWPgwzbzUrI6GEYVYxzeIsG5QXkmpSiWFfMDXKn
Zr+4pamOVXm81hRvKzv3cUgFrvdOEGbXSIDUOH3lPMwwta+Mv1R20xYryS9Tp2wQ
`protect END_PROTECTED
