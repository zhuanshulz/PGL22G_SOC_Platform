`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
clRETSonfYcMSrjGAcEzI52fcsc6QH0i9ap2CVGzVCyGDCGZPhkSusDKMO+9ci/3
sx+flP5Lg61ViD97XdyXCwX5I3hQg5hTI9jAxfmMWOJkWBLfCRRnzu1+edkPQ7kc
1IpI6YACHamAKaHuIap+s9dWuo9yBO9p5Wx/rsrYewEfZt5uc34Pi/0bUHooIaqv
TJ0OqZnd3zZvqhQTJTjOWC5aRurQ5QTalR7yKqXQPLMCcwYxynCGQTm9rIv8rr07
fpNWrYOABA0gVgqd1yXSlgjdlWRqxiBWGPgEEn1+jK9WIPesg8h3ppEWXnq+0Ind
rxmAqJ7usAT471UL8QotlXXiyFBpOuM8ukQ7rPIC6Vo=
`protect END_PROTECTED
