`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8R7PNqW+ryitMJKEWK0Gus40ytQQvAawtyVs25nsW5eTEhUbGFzg4ayCGwawuNF
eQoFWtrbJObqcp31WESFeqtL0LvzbSADyDijZxmxWPVZUiFYEtECzlOuEHKAV1lF
SFQxfkaHPn/XDXaqOC4bdFlJ7z+uXbI/5c9Ui+fVCs6bxnl1PEetbRtLlhJiubVT
yVpF39bW6mhTXIrVVLSn6+qKqaRR+dPCA+0qB+5MWgr74/JiIHzB39ZhAeNZikpy
hKMbrghExoiY9EKq9UdSZGOw4VEZT3Hy/LsbSEqAkic0jmNAQjj2fJwzDqJrisYk
YdzpCtRKQy2sBPmj5OMC7aEq8WEiQ5Pi3pEBrNmE2T2JwcyPU+5wK9njRvOxUXNj
5+cvJHatVoIfUS0XrS0G8yYGSbkrf2CDRWZACd7LxPd6xXZRiO7asPs8V4roNeAo
4p/b4h9wZePVOa4mkVyRDHsWnKZalrjQubvyE5MtuYZTCeygxjKn2FgVhL9KxkPI
9xZ7MT/OfeIL38dGVTD+wC/QfVXMayL7UfqedF/KcEnEuX1ppHudeBhjOM1cgSDy
xqxbBz88BeVuzZIjAlJWFMVmBu/dQIzPRbYT+QTX4F4dXbtOplwvAB4LHF21bTb3
vuDEsosAyvX7H3Sm/zDZGbN3GFqqMEobXfb0jEnp8Rt89e86pYq5aJBEjGiv+Crz
XNrR4cGtGJBe6AeIWIcNLkMJzZBfOzAOqjC6iO7b7FFWUafEeABpdHsqnQx0dsyf
2IJ6yziPd4sWk7Cpc0TBFA==
`protect END_PROTECTED
