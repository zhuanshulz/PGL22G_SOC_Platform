`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWAxORhnE9J5yOxzF9U338iSUvoz4/3xBcY26C8nYuFdf+Azs2G+seX/j+43EDUm
BQXg+946pZZVKF5rxEB1lbxJ/D28DjVCIVQE/TO7yZIK2lLJBvZ27BpjsEZs8xH/
Pon6ofCKWldspDoTdcJomVAL2yCC+OMqnr5yeMK0ewOd5+6P2FAAP9LcmyQFiR0F
gaM2thn2E1LZGQ9A8cDad2/6oxP2dtodeBzOIpgtJPsYpRkhuHJRxOIX+sul5u+4
78a99u2u3XmTd/qZzdtqtgUiUk4tnw6Gcluw1UX2uIIsV/XJCXqaLNCwESprAeEm
p2avst6Y6QuWIIc95tEuC7+Jlkcunl6Oi0oH1LJwU1dOEFhS9+9yl+ncLLRjexQy
Gt7J3DumQNAXUWTzUt/hlq1dhFg5F5ZH83E7D+qfY1F9ljpnYqxSS/lErY5Vq86T
TYc2P+9NEzb2VSznIBKJEyrYt4LsBm9tJBdfTC1nI2nxmLB+hHnvIDSvGTmQN4uc
7nIYmCYNi1DuoZyP5NBZ+wzGRwUq+e2QGOjZ9vrnQtjyIqYLeqZFPtaZX/VsYOfB
/35AlMSyYGXndwuFjwqMlQRoNFWC9osy3/qgbK9azHUW+0QzociPbf0VC3DQD75z
3fl15VsFaTQEUCjvVojt2O2NXYmZHzMzvX0KVV8Jnq+EfTnnJhYQXh49IG1XTPjC
5FpU4hvFWlsG6g4hsMDTd1eWIqBd4scRb07LDtrRHCmhlJj4KfX+cFGNRk6X53u/
9W24qiLgH1Ok3x4Tg2PedOe9eJwJH0FFQ9KvshwUMq71oiE/oe2q1dyoJZ8GAu2S
Ub5ZUh6RYRpvMvEUYNF6tD+96JMKBJo1LSkqAmXHsNxv6E++XgBCmm2OdRjqxj+s
e8B0jdWnOEgNKWl/Hq6YTjOyyPPYS/Q5k/rkBkHLQKGmR/5hV3wkIWBHbpe00Tyh
FSBZaii3IBWr3InzUL90orqWR16L4GxXz9NZpuYvo5pmXhTZAmbiFiOOa82pIS+L
QOSfpCI8yKh4qiH/UCowyQr5vT0udZkNJjOYHbVfsicSdhB1ZFLrsVJzCAte7Xr3
QtDkmjst6FAta8nwTu98/+uD7OLOskLBjpuQL0Wl6opo0RJ71tQTWkhLs3baxVAK
4rAeoplsK0xfrdSy87dwZa5Z6WLzyvqhMst7AVu6H1VkQEz5PNxSl1wCmo7Pya9k
bvDvrjn7jGW2INo9LAo/G1yho2ZOCe7zMcrnRSYkRLKu/YNg5x4FNgIxmnwIsshP
zLR+NEw1wE10hVf8HdrmTIH2CRR/H4GKENGNX8dH88TlUbFHqJ2DpzEh4QC24zKG
pNDbCGoPOuSVwMX0OSMjqalVfJ6vjX/j3Ot59B6byoXkftP3OJJeyOO0Gz4M6kbA
rtfrpv6Jszb0Qhj13MfdFQLv0gC87xTwN4Rf+1QizVO+eOJhzy7d5Gr4c6lbFqmh
h/hZFLW+8TKxYtXBQQAMflU7ZHdd+Jcvl5QWrUH6UtqqKQt35uNk4Zk826FL9kQo
EEgm+jKEIMpEgrdeFk9Vhh02NHSeTXsVA5cgc9qs3lhNr6AwTsiPxkQS4M8mmBcZ
CCZtvHzyMfuytOuUdtnN7e54MRVkV4PQ0yL98y7g2ZKo9HouSOMteZW1hueKk/fx
N4//2eNC6B048YD+UKwHFhFJrjVen4B+R/eOk1TLqh6EqakRqF2tKAEVrodlm3bq
KjUMNXeSATYSKnNOxLFOzh1qtPalUyQBP/7YDx/9QRl7vMUnYI9i+FMFxsYUyGms
4xR7+G6Dpsnm0IV1kxia7aRfLNjXMe/PcKpiDhPM417sJBiRx9rmTWGoqFMOu1FF
oreH1qEbPTn16rrzso5fluxv/xDWQCPlIQIiObH5tlZFdd8qiD02aDO2LeJvOP4N
PKEY6YY1QSw9WBNQ3fEWAYWu3+o9q0LO6GdZloIrpTS+nLrvOsKTE2xlxPbbFnQF
HzXwCIZZcHNl0NgBbbc3DW0XckZe8YzBgeHpfMoMAN+25SUt9eYbiCzWyjEClSBM
HOklsTOy0jgSQN51hlpyoEO4AcUHZtoP2xBqxEqtWcpVqrXGbgH+fx4GhzDFGsrD
3lkrrDmoiGXKxFPG9ooerCYM6vrzUug3muveZcsK8YNIiLKVAvuVpqAR1JEROiz4
N4a2Lwnkl/4/E+PUX+aPy12kHj5K9V2JpSjXVesBA0lCY0ruVvcFe2prFuaXODOE
Smz9E4kts7nt9PUatQ2WFfFLtrb4bhf2dmazTpAHQYwW8mwCzgOi0ykm2l3z8K9g
UlmDqpOuvclB3pewiF0tl2xM/+8xHUg1rRq8EsYietPwnTRX2iYkpE3YuEsVNrM8
xK5DLtxA/gxBuzQilKuE6aO3dkfig+D9DptU4tmnsg50S/yJkhsvr+pxxbG52Sip
xb9yLhmXnO54Y/fls805XouANtgjaXT67MizGshSmrc/YeBlYsUTOEitEVrOz0O2
XuIGM3/UXZDodM924t0cZCtzcXgv6Poo8P3DPmjMRQ2spdI7xLNvLSOzUOYqsj7e
YdKS1ToxVr2Wz7XJVdHZ4jzZUtaXpWoxwijs5KjKPIdRjWJ2DEoUMBhUrbeMZHw0
/vtJ1eYYF/Mr9O9M2XxgDxw2HDlLBwCjRYm5VHAW0/4fDAAGkqBEkHj0VIjbyHHw
ICpUwWqpllJEfPD23R8NH7fPlJho3ETnIem/oPgyobkmf5jGOxSqRL6J6st2cBrZ
Q44Pwt96Y8+R71MoSrPa4q/bPxVj0evsfkifgOTDlIXPEoZNztF5jJ2EEY9w85ac
/ngDvHPHN1r1dUY+9xfs1Q==
`protect END_PROTECTED
