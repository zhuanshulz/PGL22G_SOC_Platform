`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufSeP10sWkaKgh9h+T8hr8X5lUOZZhDDgumiSJbzfPGh6ebd4e5j/MKkVA6Ja+uv
SQVp4nQRZV448Po/Ja0aBLTcuJm1mFoDrCfUcb8adc7Jta+1Jll+ltuP56zGXho1
YTR6/UUvn5QeIdY3G1dh6EZJUjVgRoe7Dfn6Pe7QISyuJ3zS16Jw0QhgZzSBFcMr
zWbkSVWmvACrGIlOlZ1LLf990inrHJr6yuxev1udXyr+Qwe7bva8Xq1KpsXfx0HY
EEK0HCQvu3U9cyoWfNp1zML1TpOU0rWfxSqYrj7n/u8DlMIUI3dfj96YY725NqTT
zCL6IbJQiJtdH9XlMJaAerT7FZgyCX87x7FX2SVsYjpB/l4J1MK0P06ECyyLYcGO
iH20ATbm3MFcJ9k19Op3NvWgEKN74pUMVlUMxctTXkz1+w74XhjTODPF2/U0wH5A
`protect END_PROTECTED
