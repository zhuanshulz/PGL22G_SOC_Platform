`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7412BS3cGIcWstp3WTSdaDDxU155FPsr9GMzKRB0wjsdDgEzRQOx/MbSi8+ZLVqr
vXr2ROwKOmkoL5jw72ZvO74OrVVyc0qXpxvpPc05nOb3QdF/u/s3QIgZ0kB8obKZ
Cz9EpVBHx8uDNBNX4hF3Fdfo0GAJ/BroKntIofLGWc/c1NJUTPytT0b+qVSEGhg1
1FXsr64DRqrPZTHXkxdRa+AoLo4D2OwNoQKeQMXRZbjBBJYnCiVNlwQGA1X2+Z24
CH7NTw7JMzkHTChAwd7uyuuvHGlytrmbu6Vj61zfdQkxzFNVNqKmaNm930HG9lnN
IoS7q/dMzQGZMlawBWW75QB2Rl5elAF/pFjJQ0kUqNjZplWeuL8snNIPQ5Zqtv5/
XWZ6C76ZLX/e4YecY/TClw85vdywoVo+WfxhV834qZA0kQhcDP98tvzCrnaWbdp1
waLxYOZjnzyV1UXjYlGzPbxbBfHJMRgcJhUTThA1QTgiE2aqOZmYkJYDnGyYinFH
XYiqpfmr38upy9jhKi5dV7YONGSpmA35ZInipyzr4HR8MoxF5Et0SO8v4jka3W1u
bH58WKZqTK3JBqmlxWayuA==
`protect END_PROTECTED
