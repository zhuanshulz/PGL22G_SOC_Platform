`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jiSEv/s1khaFgeV0lEvuwU+jkWPfRkUrC3Dt6suFRlG1rFurnL/AcivXiB7VRWro
9X7fWcr8x3osF/y7wXU9EqivhCaoe/8XzFKD/KTDk3cHsohe4qb8eex17wT02D8O
+vL0izMbiC2dez0X9Ar/jdQMbY4Sn+CmF9nIYA4QmmN65RuynXQ2BCMf7KP2IVvQ
34D5tFTHTbh7UpgVpwlhFnzt7C7XYz3Iq0IPAU+0a0yF/euALJZ1jD7Ra+7LUhyo
XNHIvOZadOaPK3ynffem1E90a4NRCCKJLcNRnq1pDM41a4bl2gZ+aoiU2OIPMn76
W++6CXxndjISgv2bCm7jLuibnaQb7eT4/kuyQJzksaQ0zJvGCIf6ymfNi3SOJCdU
A0fW/cR1Ql1mRZrEvZ6rZh7O3OzqBz6qersJqbSpXc2cDlcaiEfEU+FWsg8GCVYc
4LDE9cFVJSHN18jkQB1XbexOkHosxFImUAXNbsbwMMjabRGmYXoFd57O1JB0zhkz
0h6nSDN/Nh750/Ya/t0enSE0ZDdCrYPFI5EwkKye6qTRNwn20EVJJ2R8n3DYiEe8
oO8xyAMBZslFSuQ4TBW2U2bVqbCGdoqdPrdcgiWJ/JRQndig7D9jW6lEVf8cUemw
Xpz2nG43HVs7jEW5TsL6VOIBmgmHUd9bcjh2t/czHDOhKcTtb01CWVDJzk88UL59
zir9g2KvUt9lpqCykIvG1RK1rQaAQWDvMI0DpFzegbrS45W3AypH4+SkOrQfGORF
6eAOLYDp/sGPTXDWti6MOl98jzuE/1r7PL16f6+vV1C3gvxHwO0WJo+QrEvSsZa6
I9upbkauA1dMJATklAEYx64maUKq9pxMMATlo+F0D/+K82yDMAHAcowq+/J1lqzX
vWipMwCCQOX7S3+vqB5TLxJIy+zq8pDHigQHw0wxPiqCSR0nBBnyhxyocvoKNZMk
/XIh6Ch23qh2OeS586Ac+sU80sCgk8OKpno2MGHtJ0NxnRHYN2GjvHLokmO3SUoc
wdAkkFPbN6bgULL+B6yTINF+UWgS9Ox2v3HmEKd0V8Z9WTm6MVfsonuIyToYIIub
5Vs5/LPHPQEmbEUO/m3flKpoCcKYn09NFuxBtKeun8+sYFDuYRwcOjP4MAKmgvh8
SmbXo0GIF2c/p/WliG2o2ipDdTmTf2PAKA+TQeTif7jF7wgfIktSEQT+LcZeczqu
V/oHOV8rU4N0zW3ftKUt1wJS85UZrmYGkA6djO6BiAB0mu6HpHKDc1L5sGi/jyba
l49f0DYB+XzLayEEmp4K/Wign8OAaZcw1asIYju1WqCg1go5bAt98Tcb2b7VMAEp
9XwAOfzeV2oNMp/vq6v/BM0gs0O2852TUpU6c+GD1kYfk4IithoK1Iz5gg1BfWbZ
aitqhk1C4JTef40YKZLc2blm9I1NLOZTCkP/vyTERyoRn+fHKPfYPAJzi5V1rQdZ
+fQv+C3NrB7mhSud2HJ6dolsLQO3NTVfehEtDj6pxfG02Uu36CL7aBdw6cV/3peT
X2yzBdE12KPq4Gw01fnv5aj4folAaqKE2tlhM8+X9aDOIb2ACbdw/H+OgR6qNdu4
UD5Vqy5wtZL//h3keC/qEidoZReqxt4GBsmbWN416NC2dELR0DDLXVJcz9aiYB82
u3OeIRYke2SCbOnYIG2QQ/LOcvWGOZ0LuP7veE7dqDPRkWLgI5l4M0S3bM1ADCbG
fXSOgAtYu1qBHV48ZUqo/z2R5dId40rnXXMXHj55XJPsd4JpBtTWEavOyGm+pgn5
kMr+ZusM+sglkIcSXiLBkFfofXjRqWMcl3uugA5U961nJ3AGvUAq82yHxfm+bW8b
MiJ/2/yMSGO6TLaDGUKi/KJfL/zIhPGn5xlrdAkr0vbxD3z44y/rj7EdcxQq+Koi
4JVd8U2RUwa9/CRGT7dvaOFYXZcBxlPlfzbYLvRoxST+ZpROeXwYwdZM/A3/2T2P
Isd2KRA7EWAdjHOR4DLF2g==
`protect END_PROTECTED
