`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KawZURpc1p9S7GlC5FXW/TKH+40qrXFpTwCBqVXZHWxetDlpevHuNgnEl7eoQgku
sTkzSOdCXONKwnoH5bu0nvw8FehCocBBIiAiKQoLylMzmd5A/l56SqN7EhS0aXdU
txxG3jDsMeWFIWksG5FgiPdh2R1W3Qiey17A7ILBxKxD7A6tn7SSihxte/CaHkyi
rNIuueB4SH1LT4Jl5kTKGRFRQPxluz124ni2u8jBTn68S+WL9hyNjqis1TZEbSWZ
xhUQ4MerdGUo2NV/4zbS8VHST5y60H6PaePiTSUGNG1VBd3RNVSN+zTeKvPOeZWz
zDUlgZ4Ny4oNkybA/AwuPzmAfLx2LVo27Av4Xq9eOR89VT2HyOZr+45jOhGK4ux/
YYhUUQMS8Lzyyc4bhplxooG0I8oJd2XURT5K2WJBUPE3JJ0kVIgRXYbZdLP+0TPE
6f0f4MJtRMmUSUGKwq7FXSuYe3fZDG5ozsKwdGHcBxgPgm+v3o7c3I1pnEfJPpiy
UquTwLOooywputEBICfnRwut38rdU/zU7ak6QTWlnIj6J+puFfjyrHzagyagrvd7
6RN0+YVpYF3ttIXZs7MQbREnJse9P3KrUnVpdkbLVkrTInnhUr3fTo+yupHiQqkx
zk4r+3Pt9+ZJjwNL9Puydx+kWnxD5BqWvvra9oXLXUO/K06FfecmOY6+cKsWPxz8
L24O7TASOk6a7/e+s3fwDsfQ7mkkbw39Sk20Y/z/WnWe/q+/nMTOVvw9NvLFfolj
xuBFI79FHn1YCou+VlV+D/A2bVRWzqv7jzPl9ATletilFSUIcqEO4QLUlliM/vSD
nR9Cg0LtKq1jldcul6czWwFTxkxP1EwFajr+v/eXgwjV5stXe/+fZVhvm1yWl30d
ANtmyHq/M4IsQw4B1B/P4Qf8zhHHRTIwPEBbJLKTDBunMBGusRDMcIgpcieOPc0p
byRx9fZ5c3W1yzUTJqKtwq4c0cplbdiFTYhxbhVBZE2vqd4+soJCoC3NS7pKz1sL
78aOrZuA+JH/WVa+B58UVzrw8Id+Jsfsq1XuaiJd1LatY2uzI4KATJh8zH+Gr4tf
f+q15HBM44Jqg1nQ7DFWIX9HIE7OSEfXbuvmUR1osMh8MJ2UVfxvB2bjIKwDbMpA
tEQ3xDcuNvLOI5Wbr7Y1iAdiIpE+nCnmVzeL6Df1DFt8Y7aNmEGV/5Wf1OzddKEV
7gFnrc0GSBV9vR4MH5pCeqs30bwJStn+jVw9seiQLyB8do+unmN1vPVfoeNQDlhS
u+5thRQU47fzPFnNSGX4ZLQp/zEzbxsVPO0XE5lDb5Gy/u6GLo35klV9WwvOSXUA
sc2t4Wuq+yslF8oqT8UyxnvTj8Z1lGhIkZLhqwHYRB9saSXdJnjhrcdAViakVmue
db9Cu1nFS5q60/fm65Tm2cqpV6DT5XQxMSjOS2vAEj2BGT995aOO1ZzkBkMZH3wo
5+FxYAotu+ZKWxdFs0IijlaYbpGf6/a+nczPKQy3x5FVpIInJPou356dlRLdEoOo
hZ2eMPxr693oa9mx+nIetjQVMPIM+HvyEePYu69WlSY=
`protect END_PROTECTED
