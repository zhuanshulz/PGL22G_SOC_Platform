`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRfwe5x6/C5OH27Nia2//LIrFblLE73xU6N7/K2aLSArDSiEYSvaa7wsX6Q6rnp8
92cPxx45gjzM9TmUm10/bfGZ+usOWi3edWKDtfyvMAov+bBQ+03tPaJDfgAuYnMv
mx7fkLhzbOB4ADI/4HKZIdDSZdwg9SY0I+11C0UGDaT/GqJz3vaKzpFVmYoV2sGm
Dw5aZWD01SHkgFPKv9PM/j0gj6XijVT2STXT2PApqYtQkcHA0GE/IhJSMSM9mt36
4cTFVyM9HEfmRfnWl6lakgETKIF0SN2eYNeHvOjiRY3TBo7nv9kx5cYu2/2tN9va
oOhgrFgTsWxt3x+ONwwoPT1Ttb0POZ6+8rsVJWXKv/5h4fwRyMCYhjTBIERyEjWv
F6G7xIm79u2AOGvuCnVmx7IZC7QF8ciJf3s9VncbvBp8N8Q8Unkf8Q3b0pLd+Mqm
jPQ6amsR9AFyTAiHO5zcAytN0S5BgQ4W5eNwnfwDRQDC4X9fSe81/IEda1Jr2T7E
EoA0E4WJJJyNCMLDSUORAuwwzl6uaMPn7dhKIQbaM9fU6nAQSeyzvzVY/V3l2DEB
6796rC0thywfI24RtmwUzHvYM8SOWf77cgEo04q62YYe0PKP+16dMQzKUAFLfUcN
dVtDuT3CfzM6fRyghSvDMvYOqfBz2ovZAP7zfceXvxy7FiIyFyFKABKcvauKJoVK
kSTiCvKHC5zRjm21qHb5vc0KqDA/gpqTEJ8ol0M99k8FRCd/2FA3Lq/KT7uu7EVL
Zdt/Tn30AV4fY2kBPwD7FTGc90egjFsI9wTXIJgU1ipMlRK4XUtuEgzkIOvrJ2IP
XJS1SAswgsY0mESF1XHsB9IvJDI59eQ9jhKI1YZR6Ui5e1+dBYRcHc4emB5QwFnf
qSCLjsQgF0QTyoHjd/FGTYNJXwhGiuFbvGaJaFACnINgUi8wnwy9sWemVWEMUMaE
ZYgLTbuyXDStvljYI3vwmuLkWiUsnuSh28bu32kR2a9y6jIssaoDw/2dyk5Sg9Se
WKtO0doiyrdnR2P3BUIX31cG63uXAcntZA9tSnZBH03Y+Pw/agxrVaryvJvz8IBr
dAjiwNivDMhLv4mfibUvdg==
`protect END_PROTECTED
