`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QspdQ0QJIeIewvKGlrsAtLry5mEdR5TChA1NFcnl3BHCOwWaMiGc2/2tfBO9T0r
lgcxaV3J6FM1pLsIzDi70AecbyvRxXU8jD603hsFOse1wi65FxF2FANdB+8hOALQ
19EdaaV+y1YhRKq5f6kSRZY+VllHhkb+C7EU9U/zuF3wrC8S6lXdUU5g09wJNVGq
o5G8WF1DYu680D5Ko1iO3Xutvc0Odk8umly/PPc524ZRLfZkOQBJjluh86AFTYIP
9vuWypfSlYKuHzmBqi0E80yfSbh1hJg0idZwjby2NN6JoR0FuI20G5GnA8XsfQiU
3aH+xKETBX3fvefRn7dNESJ/LXy6zcnuHe1sMHg/IKInyLNo04bOjiyrcKgZQYVy
Pg2/80z6yknXxwlNm2sae0Uc9Xfh9dGItqdhG2Zfbv3j5RXXH9HOosrK6f4XuAYO
ZaKO4CP7TnBgogEQn2+VG52fzxocGB+DWqAJpBEYiK5kz2XXEYMIolh4pL/38k49
rqg+KCaVh+RTgDGxZw2Sed6lMgm4CJrElJZyWn0i4gYy00HhWi8ET1XTSVv3vAzj
xJoBTRWWlbcgD5ZZUZDLhHm/57K9vtelOkycB/5aYZ5NIqAbI7pNBhXug3f8pp3i
+ch15plfggbTlN9Mt/5buCyBYlrTIWXZ7RpJsh2DG+DSsbJ0GLeXKX/pJ13dFa6F
SEaWdt2oqu24ZORlgRiaaluQif1d0LifrBQQM+1FjDj8R2otR276GYSCY8CcTxeY
NqLV2h4r67NDXedPuJXMJreKMJA/HAGYlY9d9zwibXNrT9khF09qJQ+HbN6g4J2K
VBe3a4jWsvw+OjYp61pEW0TAchR3BKW6PxMD3TE5fpm82Nyf2zRQJwJXuQZGYpu9
2Ye9Xd50H229D9ojTgjA2/UbU3FBaIomUuKkMW0Cuwg6e1iAZGqzPQLH8iLAYc3R
QhP2N96wowvv7yhI+3TYDpVhehhs5fNDn3gy80y/vDyD/tClqcsMGoajwovEHJlL
ca9AB/N4b8QCoaLaljM2k79mFo2oOQpZBJXC7HlBM4XhGBBgAfc9yPZj+HPmel1b
F3LbQdId8uF7UKf9FHbwP0SeA7YzI7V5XGHvvGFrCSmBWLBpnnjYaZ4uq9C2ATRu
R2tIFz72WS6S8cCOMO0/Sy8v2BUZxJCkbJ/+jOrBiNEioaPREzbEkw6w+H44A1oM
7StCqt4d0QKldwHDKp/j7yNmq2dG0U4tZ7ZQFLPwAO4=
`protect END_PROTECTED
