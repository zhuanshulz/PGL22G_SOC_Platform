`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJbTPFFTZtrFy15r3056ib8YZlqn75W7IPLBdEByQesY96aBMME7AZW4yR/LAPQU
zj4Si2cOXn06lbaO/HJG4eZ+LmZ88xmiMOSMzDW8VzQ0waBN+zHZpuHGtR9prH0o
fR4/5hWgu46MnnPncAWWQnTkI9TycQ02oe36UOzp1AsnNCT6k4pvzHoGkqQiHkdK
QU5HjfZqshYMORYWn+iQxpoozo/n2HmfRHPBMT8wWlk6rDQjhjKoP+GY12KNstwa
h53zQ5IT88xRGoY0C2Uv3N8x0U9sjvQowTmsRYv0jnZk7zXS8nmT0a8L7H0kQQ4S
OSscs5HgmLQzV4dsYzzxrq6pDDSxr2RLSt/ScGQxvv1+DDE9aQLbbfujQcYbXk4q
8HG0fjZmyvAzLlwlAqQGpqaosGu6pbMl/qsy9YeR7KYuq2t+5FFv4DBgo2fDmpY1
v5itbkpt3ReUKy8RaKFk4ycqTBQaZvKbt6OY4AvqF7ffW95imSLTycGIXONvii5a
FKxyZUiAwmJ7y+liFXhOwZil+GQ4At4e+O4cJ7t9rRSfdIi8MRbe8aDdrPVnXlM2
4VRdCPEh7Vbw3Z1mpALy7cFzN295JyOfxNueflaNQU/Q8ojkoQ7oF9cQ5+tVV6Fh
w3Q3OS3W0yWAhS6YUYDPzRbrz/a8HF8Xv+p4GyUcY29YaIWvDEbZqimm4iPRVfPN
G3x53hkqxfx4TrW+ynA7kTl414f7pv29rDDdMp8y99nGFQaWNARNRMSnKt0wgrGX
igtQdUVdVRy3VAVSqeBeO9z0/tNNp622IAF5ht890ppLUnp0OkAEszLllG3wjCDC
vb+7VffNeMRZ06PWRk9bzUkscBm/3g+nYETf/28xXbq+IPLrLivy0L+bbSYnO8Qe
WD1e5OZlfMZnFnEXbVdu/DhwYFeaGCN5dOfWzkx/ErsKfUk+hswo+K2i08mYf/eJ
eMtAaMxIX2WAB9untrBNwmhmIg9i+Jv/1nVr4qQc2Jp2WSFRzWBpMV7qGczm0SxV
SrgKYADl7wVm58K+4PnU5E/VNAdS2C3wkeIk1h9vhgw=
`protect END_PROTECTED
