`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QM1anQj4Nw6fjQ3elLnZ8K4inroGKUaM+QczsOA4RoU7BuU2Z+Nu2kyPh5+1UykX
LXkVOIOgXWk76JK5cMTEB+N4SrquvvO6QHyAcNTHno3mtlJfM1USNnE5s3nXkhrr
nqOw7LifeYjdZ8iG6SWBPKbemm3RuoWJa7Wzlxkxvdo3lV/2gulNAB7quWwwk/Oc
Od6BcOi3zSdr9fDjOFn59XhBcgEGFp3Az/PFSRBf7l0R0YcPmJHgUr9m+INzRhpX
u9l53ch7efdCrI0ixENYG46WV6sNSED4y7VQ6uLSwLfAcUr/PntWJTPT8MJoZTJh
QrkPd2qSiWT4/AG9i52vyjNWY43XaRNck+QuBLTKRxPoFOX0tewmS6RK5QdIiyh5
XnHnfUsc+Qmgbh7Y9uJ6T7HRaCvZiCBqcFn/ZUnCG9ox7MmD/8rZzCRVEsHsH5EU
aygX7QOVTHGqU3wjXelmdunowhwrsz8D5bVUXSsce6Kilwt8mWMFt3vGWHX6vpSi
UJeEsHPITgRqTx7U+0ZezzItwch37uBy20WJWJpDRB9MsZ+t3imVXDOVlbYrvD+q
ZuJ3v2kdVkuymdG5QWf5FLx5X1PnceEa9R3F68SzFRVyuN9KHsbos43fHa0Go9BP
W2Dvg6t8IHEYORQhuaYMF7Rr5nDnzYCWBWfPEgzPX9ysEZ8VYy1W7odQS4M611Y1
y0PV4HKnZxPFQE3bLkMEYtXvRgAAXSckLSOsp1bfvh8S5IQOIL5+VA2JY3+Wv/4T
M4TkHa8cjjX90DvZp9a+Y1oJSyFL2S9aZSApkTRy2JN9dsvD206Q4I4mnba3+SC/
2Frk+0IkYlYN1bbEpNswEQ==
`protect END_PROTECTED
