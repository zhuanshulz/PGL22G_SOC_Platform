`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjxKnfSigmNpmyQcVJsPE65TX/MS8GV0ho5a814wqV+13PNQ2Ppd+KZyCSM1kSpI
GNBsQBym3gA6uiLNZajyk3U4X2FaX327Xbg+aV28FrJETlGx/IZkLQzO/iCFDBYa
TLPuFPgXQ5EOEtscwEfD69b0R1/cIIDcu+XrPM8FDoswxZkM1KQxKZKGc3XMI5+s
yMlxRRuVjC5eSLBb2s9zl3A6t6MHlpN9yYsRKXHwTxemQ1Aq5810G5CCN/jHRfXX
1icaOmZI12YiHWsdCbeqjkRb6s6AsNKQ8F+LWp1Rw/QJzCXjUdN7cNhluKbCcdPh
E06yQqhD/9jmw2GZguion/Mp7RzQw/mKQI0MAkIhRtIpYInKwLSoE+93dTFizwBV
DtHx468egTOFwcPUeKXXLxp+KOrPxxn/lPPNKH/UPWUfsidL8ijcuLP6DX/+FfLB
ms8gqlM5teatmEO2ySj4g2NpRdhipeGpAZAm67OzqUkcN67d96YCicf9TBdfOcbK
fPPOCCofjTrXBb+tiV0x9qGHJANU/c3pQe/Dg/5C/fA9WppbTp8Yqjwlb5ObQh5f
362vbcJQOBdP28BB6w8yaddcgZgs/PW23c87JLWsUma2VKGocgm4pSJ2Hz+b/v7W
9XrPoLVt+CbyZJz/e3hUAsXHf8Qo3YkJBa/Wt54ToOUhxYccU/jwLupIzlNz4r4I
Lor1tSf8QDmgQX+y/r49Oh2Box7AoSKWJd2dCPn7XIgyUJwGYWpTilASOZeYvlDj
EAH0kKVYddhP2n7iyHry6plivLT9hjBoZcz8YuRyrwux1AKF/ImdvkRTL6PoSQAY
qGkCMnl6VX/lt2IxC22JX+zq6B33EvMOMov3m+mdh1C3Sw9Y2pyaejsALHHP9Sc5
Csg6OoTx/ZmNrWHKu9xBnOi2pnvr6GyiJXpdc7PUxqz9yys5zaR77VlnL8hBOB9c
c4WaKch49dKZj7VlNNTjribFlYofFV+LJy1G++f3OiXjaBhgoYqR/uJyA7lf1VNR
zljrnje+8QjAZQ6a+sNNpThgPEJwpjWzTSP7AV2PpY+0jyqQSDir+PpdRarXFbEa
U7hke4RYB4OiyUYeWuuAhnGP1bCjkf+hEveD2o1QJ4x+55kr8tA1SEz8RVp6CoNe
xerRyP1/1yVBUOo5T5BvU/qm0nTMahxM2eA/eMBfhwjDDRfjByrtNLJUcCUo+XGz
+gASiwXBGkE1yPweOpEEOGt36rjGXre7CwTLUOAqsi8=
`protect END_PROTECTED
