`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixKnEAOiFMtOVgYa2tNR/9f87hog8V5MgvFQ5VtVyekz28xpt+IStr4tnkfWTWnn
OnuZqea1I7QGb7kR79RhLqWsAk8srcwz4gjwN1k+2aIVU2CUnrkNKCUnsd7toX6j
IS/6oK7mNXZXASj1lmPfbxO6P+NQZx3qBthuvQ3gZKgd0D8mKd41diENUB73rP3m
l2bZrZ/yU8IsN48KvPrl2zJzi9vkb5HkFuZiwTe0BLk3x8apswihgqbVhjxLM3JC
i641mPXL7vOICEL4wepVKFUVUqB3ZSpi7MczSgOHRRfluJT4xj4zcT4MreVXnRWh
vKvz92Dum+wy2+ytpeCsnDw/fx9uN5b5XnBmUVobn5AzplqY3XNyzCnsgmSqGyZD
YVtj1cZy+7l6F3HmD1rNAX4UZZA/WrfZmu+rSw6FPyyeIzLa2Me29s2uZRNA6OLM
kSNnOicujufeqKh2qJZOkuogl0MYTPxyQWIVJVqKxahmPwwAxk3/0XJWYVTR3JQB
yRUsuy8u7RiBA27xHfb2CcbZA5T42g8DJe684Vby0U78JzncgYNSnhxxmxlYWqrL
4T6d6YxWgK7DOWMONknAfE9h2hb2riVugqD8baflNtdsO6x3LPKtlpAB8cMmk3Al
4B3Jn2fpd1/bKT6DiGVpTw==
`protect END_PROTECTED
