`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r3ih8aJOx1d+U6OuUcEGzOlH69FbszT6af9j0hEasGT4n9AijNv+SuHpP7k6oPil
iYH7Q774nCdL8v4H5G4o8A4IkP40tl9DTX2z0ZrMkbXXSh29MFU1macmBhA/1Uvv
DHtiT+Y6Kf5679/nyuLCLMHUAoQ9V4mEDziN27dRcubdEAdETXFlLLu32lTLsbZg
MCFOuDPddEkRb4RuKWZrGzS+r2Esg9AbvNcKLiJ/viDqwzFDdWJwGeG2vLI7hWCT
JcO7SmaPI+WcQcDUQ1L8s3kg187OQLJh6Y5Itv/ObtSMxNvUdkNHs5gg/e6Qo0R/
Z96bowbAy8c06ghXo2h02rMRG2bP9RMOsnnOI3kjfuobkf2PWv1fDmEtyc0e+mYS
ceC+DtvQ8rXAipzMLT/cdw==
`protect END_PROTECTED
