`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggAMGBAYFVbIjGLEhjv9sd1EbBvFYKlsKUelyqtsGhK5iGIQFyTi0s11Y0T6HZSa
shJaD0JzTepiAcoiw5U3jTn/nm6fI7vfcNfH9d7/fOXufgMfwngjHNavc8mXIwsK
DBlBvAk9Fb4IoH97r5XyQ0G6kYb6lwyqo2C6iwYU4Y/3BG/HnPcZKyWMloSWLQg4
cSMu0ZOvKvVblyqrYiw/g8q+qnQifszczDY+rytS3724JtKGBVbhje7Moff+6Q/l
aG82LBczVn/UV5ttVZceiA==
`protect END_PROTECTED
