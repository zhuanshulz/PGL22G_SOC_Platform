`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXIlTrXja9GIoamnT3qNPfplv2cvaHcbkR5y/aya8/LON5Yxre3POUx8fIuhtS3e
O3Hs424so6jkTjYn5DkeKDSQObGkSc/Mxm9uY020sVjbXKbSytR5FUJQPoZjDeal
EOB97TkJLvIdNkLnUwcuT/BtiRU9so9SHo6CUYkUqPh5cIH70ZloO2xVyy8pQ9ue
deDo74oC1fO1NLq+lXOW+oYD4jXvAY8FoLOCTMj9GZBPh6xbPmykAK9EDTA3fdTh
AogX3JZ84OE0aIxQOAHHBDZnJokMB5RFirYWfObeVj9+UIIDNg7xRvV1ykEIM0jz
g9vMTIJHhUN2PXZx8VRWNY4gMksJDaD5LEyGd+KJOc1/Ruk3WHs8UdNFhmRkqd2G
MlYQ0aS+B3nt4he9jS913YFm0onwy915k6wqgA2QYY8A5Heww7mOOLzi0WMFpme/
wJ+UtNJtTorNNQ7P1uO98elXgXeuDSBFvte88buWfUQwugJ48a8mL2A92+nFTxof
L++quWcci7hc+igsW2I9i8D6Ge3G3fupP7gNqtxb3Wg13apsrUB7Fou6mF5eJpXh
IWACiGJlvePJjy9vMKqBILNdCP0pXjMgO8cIRZvSAC6xrJUWuPb+k8dq3pGZGvMz
r2onJCt55vj1wNiD6c7NRORB48sIKu+yuFp1Mv5LQWRZNyC/5cVkP4xwvJgsrIGN
FL4KSCWHBmnS1DYbxmTn+nNNWfe10jgpA7hXW1Cyt/Aanjx0kcT7QfSpLkjbSeGZ
3RvmEA3KRp6kZnM5YRrgPsWzvUrKFhuQiUtEyz9dTz1W62IkKhkBo4Z2WnADQfQU
R0OfftTWBSuM1RP+A1BSbtSh0qm9MSk+AAlmw2QzAsoGR25PhPWDK8kN0qUgVwwm
ZlshDYs47Aq25NL5XwVI4yBSMtaIg3Lx6wh76Cy9RzubFLINPWHeYNawUUssZO14
V9J3VBM5xGJ4FnA7ERR8SuB5T9IzIutux5zv4Rbqi3+EhXXEAhbs/PW57c5fCzCE
tLLatEtAE0uBc8EDtHx58VBj08ZdYsf9xOYwtADufK3O00jC62nu/R/8U4W1+tP/
OlRg6lLYGjUYnBougZPnRzrxBsEIf0HXUUvAsHsqcdz9xh2805Ep/BW+sFi0W77k
8GoydMOnnpVwv/oBAQz767u1R1NqMrK85KZQ9c8aRSSd70ysqkaqXUbNTS2ZPAgR
Np5wfVSRxMU3FLr5t23b6TJm05Quj7yZAvpVFEnDnuy8/NlUKIJ+cvSw2oVBgzfW
HrZ9M+E1ptpQ33X5FJoxGyIwxv6M49vPcPz93LvOV3HOh67MiHRHn/+GAZCCm8u6
KGMxDC2Sxw1sUE08U4eMuhMBNR11Sb6NKzshXOgmt8UrV9nLZtoIaeyEeK89L621
yJpVv4Jz3L9XBU7y/Q1lZn/13Me6OAjuYD43ED+FvxlfeBIBnWQVmfM1jii8B2R6
0zx3i2atkJxgN2XJmm54Kp+Yu8Z6zHqpeG8/zm0rfMWUkMJOoA5aCjbqJB69wV2J
SWJ43wuPsdRslbaOia8O8kx7xd16qeRp0to+I8F+sMqJCbObNsM1YEcurineCa8n
JbhFzxcmpfPqo5tH5/yk++/NkR7AaYHGCBvqY8l+lrUHLWeA9g8a6RCOVesjBihG
xA0RFL2UilW6lOiogxkY36ay48A0XhuDeMhZgz3kPb9jS0KJr+P58yuhDqR0AxBd
EVqz+X+GhrENAS9C8c5P4BTxlP7U79x7ZAaRj1LLw/vQjwNmjNAy3UnGcHtDO+Ee
AM+LvgZ/TwrB9Rv5S2Z8DML4SB8WH/LLohtZ3VFz8vQtZTjhAT3gVVjrRKBQovVr
DB7cf/45OvAPOZUUfgjpz2OtRFoR8gpj9pV+GXQgpFC6xLK0lCAlC46M5qgbu/x2
4DU1/4y6bFlKK0fzlkvcd0xFcNQz62Hm6aX94+1OrzJGGSCOnwu5wUBEGTETtz6v
2B2kV5I47frlTWoyT62SJ7DQvL9glTKFs0pEg1MydIZdyAUv2S+7tHZo/dWv/XGt
pezUtghSCGe0N1JvQhF0tWqlyYEMiyj86V8eUS6qdCN7B4zZyMyTAymUAN1VS3oc
EautPykZ302OrOQOd44F+uRS7r1wAFc1PIA72kIROFI1KwIqHMqoDiiZJHa3pe0p
r2L3EKdc07HKa6aFiwbrNutROzXIlPudTGl5vy89/jgat/GdEIZG4Lf1ZPFdVZP1
3xAQTsGm77snMYAiVo6xQTtPhTlro9Klrw1nYuRgleuEM19mHMVWZDz7yaewwMOF
6ZxZ2ibiH941G1E08NoPQrHmkon/AU7RDniRleleeoKz5qK+gZOeNEP19y+5vfaf
hguvCklRwQRifJlodzDNzKxXHgNTRBPIJ84yzQODnMkwlxy7boKtawIj0vXPuMyX
ATbyPRglhEGY4Y2w3zqMzEMxs4rMzcbZrOpyxmlcy50TZc5cBT2ttwPQ9PDjlIY1
2q/pnRkmPSNY2L8ofKaWwNdHpwwldcIFbG38VV/zDeZt8MGt+cJKyAo7cFxqXUuI
N/njP+GCzhPBxfRFuRBMZqBd95o1eZjg4dawJNJBAVferuANtLkKodK/IINJRrXm
ty+tSZpI5zrxywIhIH1vMCTT+N8DSx8t0Vfs94G5S/x+hOKkADgFelMjUoB3bx7M
+abp4oIbKcjyQReb+oEt/kMxJqbQCg7y1sNK/0UY+uAuEAvE/niEWRG1cz4Rf0fl
4lwHsyxIPeAY2sPNMlQInu7aJyxNcLxXPK2E/0AqDmZD+egSOqEVdH4JdXBaK7yR
owi0kRNddDVAgpuR+LPCLySxB0XgAanzilPUyQoo3QTWO8VGRqkj3R/3BW3LrEtK
5zZLyPggt7xLJz9tksPub02oO+H1Zwl4Eyf90be4koboZwiDQuZJEDlCEA9g1goL
ORHld0DFqdbRedl1FBBSaC4Md9kxej21dgI5J4TFkJzx/cHViuYwmnkOo/frOogO
BYZMRPaVCkWxTu/NGa68Ia14DR2VNf62hnqbCVMp4DcDKzTEvmBlgqBhEjkXLGv0
nV/ng+0KFVkjrpxtCYnfnWvuzW6NbPeDS2s0l5YhZwmQOCg6A7TrmgfMTMH6wfxl
mvSKPWudjADZQQd0zGbEUwZWU8WFuOHg7OY4mcOO7b+paXBcJ3T0KSL48jBR/yKm
qg5q9A/AZ/69+T9sy3OzPZlGhM4IMjgQ1zrv6HpS8swkhRA+D1CD8pR326Ztg47f
S01vCHs2inhfpkD3qylQsy6nrMf4Xp8ooQ+X8r3yT5gyvIP0uRXq+DRoPc+D7+gv
WQ/6D7aAvYMLtFrlv48zFf3ZD+32WnQ4uL5Cq/H3Dsztr4wQJ3V5FfNIQs81pKbV
3KN7aviLvE9YF3UAx+4o80B2lSmQxK9drtX/bUXbTYLWJpAWj4/zVXpvC1uHB2I9
7wsl2UYRCZEPJsyBzuUFSxWNp0Ehiz73zDZludsPh9yo5AySFNy2sBTg1lkgJ3G+
HqbPsdhYJmdkLAgdhhnzai+JgcjnOXqibstnDw7W2jA637hdiqIs+oQupFjR+Acw
pNW9hWUBpvT1YplucHitADJkvXXhuy/hxHQkramMtOi8idenIB8HrcGD+hlPTQj2
oJrrVrNRuGM5Z85hFho82ykXKTHWr3K7P27OUTwWDjhO0CrXlqjlLwj5pQPdf0Ll
STppaD5iiDZzTgM2svCQ7ZFZX5t6GDXthyQ2vBJWy4AiezhvHhSzVxotgxb4B+MU
5pvXsP4qtJVtbrvmPAaZx/DrEluALcyJc7Jzi6z7LV/rUcASZVftvMuOqQWKmYgy
dZOZTqf2SyR+Jiyz4h3s4CGHdGcPrdzWJYUmh1B+P35/pbzxfJYqhV9jdZUDyJdt
dbKT01TYqcoJ3B6SXOMc9aJMO8GaWx9mmmT+JS6N6hgGxgHt74bjS+5BF2M2Acfj
6Z8Jq6VssZNR8gQ1J5yRIN3T4uSnwF9JkiecOZLjOlAW9mQmXxAF0wK61KTStb0z
MPEWEiZZN55RWtUXcVFKUVtKId+98HY4ZmsHxvd/jeGVDR+GlLaisZ4aCNdY9oHb
FAA3U3sGjplaVwiOgWxiRF/xHPl78WfeMH87KTbhJhSDks6LJ45QZaM6U5ud/Qj2
ncxdMyVBGsldRxQQGWT+OodG3BsZ/ybz4P5xxVGEbeKx68BlP9Jcqcr5wQLZRrWi
I77PywJGJ3usg4KPXFJWciWFO2ek3zPyfPm26toU9Ol8myxiY8Do+fjSeDf2DFiO
q+xur6br9BvBoznhj7Js20nW6cyJMvLVDnSvcKDL8/V737QFXmElO6U8ECAEqfwK
9Dm3YkSYI4jAkFw7sRnPMzyTeIPSfYdGKe883qnTnUHxf+wYbOOc8L5PVYVxebXj
`protect END_PROTECTED
