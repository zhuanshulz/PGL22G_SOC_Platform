`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8W9zWWRhgNSjzSisOJwZC8uAYk57B402eJfcuqqoCxXg5LRXmBWV0/R5xWnBFP2m
d3i7wTCNkuRO71AVyvIWBT0xHMmAukFq92e+ocBZnDUBYFSNYGUcy+LOQrPXAzAj
RRPlceHPZJG3gBzrpdZHM0cmd9QTabjombmvL1D5GOmUamnsKOB+MVvFYRAB6+eB
BrlMnyhGnknycILMknOX2TCrO1MJ7/QeiAEoKuK99kWPqWtZa8XcWssaSrxwsTpE
ULneVQn5v9Et/ZGfR2h1NdUPkeyVi/fdQhmgdnT1ypAT9ksT1emALlILrnjK6OKI
+ip6k2FuuqM5g+TNib7MTwSRk40mitdcOHjzmXoqot6YsPLw/jjYILpuQoW59r+6
xibPmCUC5couzafAEkJF619bMcibxoKr+Z6t+IVTzeDrF+QRB60SJDkXwcFC+rM+
su3zGFHl1NyoohZfMJtdziZ5Yv9HYQGJyCNcmmemkxevSx3wCSesZlt/nmWGHjRU
IzmR1oDgzcJ1lWCwRzJZ7GuZiu+DyU0SsQXDB8a64oLEssHjX+Skul+Mg1fy1yJR
UGjJBXK8qrFcg3HoC0HAIg==
`protect END_PROTECTED
