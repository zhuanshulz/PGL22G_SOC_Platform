`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OJJPPLrsQZKOJTb3La2wrXg2aNbo70l2AmFwiDjTrJFMxy8111tafo4c552Gtrdt
u8bfZNr20NyESXoN9nlOYs8uDjiO7gpK+orXYQot7yHMnB5d4HakQSn7C/Q6UDlw
7PJS3DSj2EvjY/vRNpVgaE4UNoor64uGNx/bte/4Dyoiycc/Y1J1+i0WRspDZ4F4
4/gfyWAgKCI16mrpnYiJ+G2g1RVg1EhsyXHWSn3aQ87cUNRWkN4OZVpFjS1eYmzO
xt72v/wxKEAFuW5GeA8LXGVuF+LQFIkw6m8KWrSn+Z+rryHFaQ2EvVDLtkjsNSiH
086p5LXBG2SfLtlOofoicLzRZ/RoYz6O8M8KOf64pZ+xyPnRd4yaft9z6ZSe3b2Z
yEaSjmSavZ/o2HLx0QnL4ctpIkK6kfU3leRnTfXfZpeY2qmLGOr63cOtOT6JfM4U
9L11hLj9k9IKGFUfSF4JIWNpJPHJjqGO6V6U3duUXtjfpp83OnKNeyKbcOQAFYNy
o/MpI1PrVgJCF74E0brK6bfeud1P71eLPg6NUpLJnfvOHAyo5RTsNllIIThPudqp
Is+Ko5iKZbSpejHTSBMNHgoTHFBsveZz8gKj1Gqk4w1LiNA2PbmWe3czSy9lt7Fm
`protect END_PROTECTED
