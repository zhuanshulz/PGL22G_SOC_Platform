`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqUClfPCoKtEyd1kYaGfdq3mOHQkAjI8yRMpudunZ3i4TSM2YRQo4p26y948nZ0K
BE+5qIYiaemLbi7eetCD1eq7uSR8fWOx25SLeAKJV2I9i7wrv/Zp2TgUaXbhb6rV
RY2yTXlbUx/uWUN9ZJ52fQmQg4xRCje6iWuOY1nN54gd9hUKi4nTonR/l2rIhYiY
a+HQ+tHgXjoJe9Bo2bQ2OkknDmA1rNHKA2SjVBZjBwiTH6pszd6itvn1UKdEJKqJ
+BjbzSKqimO9JUXoT/NzqEnKffQUaLC4NZDDm/ekEkuDE+yoMaf2JzsTwddElI5D
JMyZxO6KSUR9qwpfXpQzCXOcqexzaM1Uq05VAgb6KKYYcSDmMgLXuloWQImNhSWw
XRGib2atogIIblU5nf0XTnEvrzNSpkZZfwTAs/Z5iVWX9Nctr1sdFCBIxd23E9A0
lCMzIBXRrCIHUEtqR0vpne41Ogzpuq1BiAGCMrLyAInnrbUVZMlfvZQXhSpNUoSv
gX8wEYMFOBddr68ojOAWrdmT6HFQKryEWLHHol+P8eY9PEf0IwNy60pWgFrXCh9P
eSGVQm8JkqB/PTydSNS8a8T7azOCdnT+TwZeZkec6WbLPFn7XYOm47w4Hxs2Uo0Q
MzipwUaSrCt00+u2X/0gsX/qVCfICAGglE8WqSeapDZUWgpyiB9XGccviOEixLa5
hFMgGUOIQYmVYzDVk7ymaL7gUXvq65mF1cjjgopMlxunJ1knX7FPAQ9JnLj4OlWS
FINWULQpyQrWdWWbOfU+TMiQvsHpLVlqdaKfcrCLq3tXMP0Ubh3/Mi8IW4yWttlz
iZ+HgsHDs8kO6cGBHEwVm7cz6cB+mfJVpIiF+zDcglmqqe8QDk3mX3WPcbHD4OSB
hxGX2ucn2NQYuw0cegyC4xfZHN+1b9Y7bT7BlSem6L+ejBi53vDRhAwBRvkeD4VF
cZ3M/C9CTenqf+y2HxiI1Z7ExSDa+hze+eNQ7txljvVcBf2Sh8VX3+TMO6ZpV5rQ
cou/JacDMcguwTrcQ4S+sw40chIXrsyRiwW8CmTI8zIV29YdiPwUEqS3grx2brA2
Xgd8LfNdYDlDfprk4qqxfIGv2Fd8bOB9EM6IJqWnyM6SO1jpNLXdFrk5S/zeQMcg
++Nf3iuVjSVa9w8PuNoJuN51ThWorH0p5pd4ts1sgZvVGcW4CywZr9CJ3fZ/+NA9
FjgdzRr0PM8HwW0ru97QtoukXgQ2/fWyDP3FsmVGTvjKEWEYN4YxDSi+1oAkGnVO
ExqVFiuVnvxxX2ojAtnn+vZ2oQEUk1kZfRPUdu74/dUMssIiE12/iwJAKZyf2hSm
yZa48s0OUOW56biBoaKRqGMbHGYcbsC5BVknBB1mUDqvufj5A7FeqgnVOWESY9RX
Z3dEDPAIbSSzdUKdGupCUU5/rGmAsvYCcK4nkx/VFWx8noEZRfFqNNKuGHHTdwDV
8a57WeS6Q30I2FXtff6YxkDnuyB5j9qemsVeFVuAZGFmbqCvpWXhYtB1d/3UtyVC
fP1SA0b63TR6h8o7LtkSq/eBmZqwsq8EV55LDevFL9XFfSKIj3CRfrzQQDxTcREt
nxAUXm3dgRou0g1t8q6dsz04N0v9nI/i6CVnfp1wGtGD1m+y3jQZYSza3dUYFnIR
DdJe3oPauJmxm3wzp613KYNDjSlLVI43s9FFO5rVrqOQAOZOUGquXphz7vV+ItrU
ZaOWkK9yU2i6+S2l3LpuIFayJ8A4fzXiPHn22gSX2UH/ij+0bOKb0x8kvFBDeeSt
MuHQlbm4Pnn94miVvcjp6sM64hpzqGzgfiN7C58uPrKVji1+DXc5hi1OCEzceKpq
cNbH9D4h3cSzeXgHMeSpXJqSa45Lr6HGg7oKNEPbP4lLh+2rdCnBBVSB4k2qE/gM
Fet+rm+VhyHhbldZQ2liT6mx73wqio1sBeyiuIClgc4ITTBybI0Su8NehDvk2qkf
d7ECt6i54y+QDEh0G8bSwoNEFWOnspPg7aA+VLCYSYx/9xysAlFhhv5AgsfQ33FQ
BkZfixezC8YiRjvJlrzdhVH4Sa+ecPfqQYsqx9QSEI9XR4qUG30NwlRYfF99roOW
Q5WzxL8/G5sTb7lCJXB4UyySPeZCrmmBEj3leY2oSekBwTS2/XzYSF7DdsG92Mv+
Y95a2pOEzMUlsx8j3K8odQzKr5zo1FzMuUjGZDQQZ+nfNwLqZTcx/mskqACcQz11
8bU9a6DHYQ8tViWjPa/UbtrXOY1Rc7bBun5K9Mgdq3ie60nOHMEzotWIbUheWK24
e3ILrgqrG5oZeJ7U1PtqhOlYIyctWTmfolsXiLNOkY341rLFsYcKLPwsOgtMAOOX
A5nEWagJs3LdcCbjmOkLe7BB+fd49Mj+4J9+ejo9RDpQ0jXhrOLQdvOU01xCSyMN
w+x2Ma2+cT6U0xl4WE8VkyDQbriUv3CbzW1BiagDpVQG9kJ6tOZ+0ITa+yjPYgqE
Hoxw4OBA0gdcJnsJcgYCnrTGR1+ie9E7FF6mZLKj6xzTFN53SEXiLRpGIPag/WsF
1QOatPujGGksP1dsXOAJstEjKVSLvyAq7BJ0VwjuLIMbMTCvoHta/x0tcjnswfqI
alYx00sKHa2rD92zaExmdsJscaTj1VXukWKuG3JND+zYs917Xzo+8lAbm3MuBkjF
JYmUanJIKASaWQvqUahXTUpUlsXdfu5jOsXX5hUQ5B9cC5GvgiV3/fINIrMocHT4
5NDnPHNRmp4e4fWFujy7Qax8M4gyrTrpPjG/fg2NnqtOJXqqQwKBrK+DD+4Rar0X
0V70V9i4VtanNMia/t3IF09ITNfwIt2EJSuM+BzERqCKt5YO57z6oDMXDCMfqFbC
IwDT3TZN0DcOw/FQBbUs1MHAAhrQBaK1lvm+nNUeX9LIDdggJ+S1zmWf4mcBLL+f
uIq/C0O/yOJLQL44BFRsUY65xT54CMIhxu4Ou1gUeREwwNz1A0yZMMmBgJIQJW4y
2BMtcXy0QIBSLriGOcUU7JaTIQCI6sLG5YjWh8jHOKBN2RWpDsKCQZHyo67iF6dm
6rnT0zY17wTkiCMpe2VRgV2gDAVNjVke4dUGQwJAYdobxntJ7TxedKk57rR/tRga
oON5AWycoOJBVGX9cq6v8va7NcniDPYyOApesSR/FCGgoRBAYcknBg8N0vxaFKMh
VUF8b5xrvzqPI02th1iRkjFbcc9IdzWQgPB+9UF/Rgzvmn3zZQryBvyKfrjCls1R
A3VmYZWsPlIqX6o2XafIDrG/tgCr+CpltiGSM1ict0gV4lCd9JEfFaQrAHT/o4+A
kJGybJkOQ/i5EfErLIvYNNrYGVGEUp3Y5azDpRINWE3jKxH9lmqGghcMIsbDMQX0
okcyYdxpDuzmz2563Lb0T2XUleEP0387xBeejvOUTnfrjkFPo+JVWWh+5M9VEIKm
RtzH4aYQllc7Q4Wz1UJbrk5n6vwGK1hE0jmwYqF5ppDop/ax+5qDc4x3sBEnngM8
q3xWEQoBFXK/8HByi0TgdmDiyxKDyS9v8lJyrUs1vY50aQUjHP3diH77FFs5NMVx
esSQqRyofpqwUoV3r3aDdEwz6Mo4RqTAa5FK77hLOyUwrDPvseW2ZoemO+JFmb7L
8a11Rcq3IbOLJ9sk4Kh7PwewVtfswEccbTKXXK0blxw2J8w8WdxAdLskWw+/GzfE
0OKNW4kt/6bbvbBCmwOpjzyj6qHjbnMuUWjgm2UGazDXrnRSqe2rPTxhEWd37TA5
wGjADXSLgqu98GB2F/sP2xS/ph7jJJ19lrP2wMwEtIZ7yn+Ww3BnU/5PutgRnG0+
Ct4FS5D+mejbzIVRLxgojz4L20TEuc/idsub5WSPbOAZxdGilYD7lqPUGl8ZjzWF
keaDSQuTMzCEd/8sWKGQ3DdP07XgPyqQFe41JUer2v5CD4OlLWBr9R5yRTh556mD
Grnce7y0Km/VW6sow/oYaOWyeqgUFIfonamog9SdPy4Ulis4Z0JsmWApycaqX9OF
9aiO0Y5WwyGw/5OtRBRWpVHA9ZLf3C/+EP+RpyHuEA9ipM47eGpTVmCM8AJpSubI
jJxfKWr/OrNgt07bblEi20PbAc3Sfysd+C/o8wMGv91HFPEJ0y8TxnihFqDzFnzi
jgiYKx+ZonIZfX0IyynEY0p94kJXJPv+UlX00IKSlZ7SaObWJRIYovKCxoY2jbaX
JgFGwu2L72d+TT1cVUVc4MevQz5VDC/wG8Cu/1Oim8auia6uf9rdf1dS8tH2aDPj
zB5VoPS7ZrWnGxo7kESM4E1VDms4TOaAZXW+Aa2ST7KHW7vbV6m30KHCS6VBnpDB
4zt9ChaCoyJJhFzXMTxABf1Xtn4hKZiBNTuE8YideQ7aY7DPMO7jW3v28jGJfAEZ
++ozrXwvZ99ule3JrDQfuu+a1q0/z+21TUSjGwxA8KfOJfVgvbpq5yceYgd9Tk79
etP8QaBLOPVJlbOKd2CsBwk+WB/xvN/dds/8Sb4vORMYaNK9k6NYobgD4fFRrwKV
xD/UxpcBXGrO1dpclUWSldtUDyU78kQXyZ+XZFPtOzPJyruDWOMke6CynMvcQO2h
q7yoVxXvm1lok4+4Fo0m9oXqbNnjXGcIj6yGy7zv+tQdrFgtkoi9vHQTt9SZJmmM
KpbxqMfOvGVGVavLStPc5uPfwvUa2I1dFg9TiSpF41JcqrB1JRimfLtdBYoPxVQu
EtNntTNNutSd/fV6lsuUDOIg2lxyV3j3XatI87J1c1Zj7teReTazBPjl5d43kE0C
kswbL6exa+btrE/qrd1tHI4Fu2KsFLxJ2YqynOs8gRpBTCpA04reZ/uQ4nBlqAVe
QKeS+NnKA1KeqUH4BED4ZgY7weny9w6R4kT8FTq9dFqnfPM3rGux/BgBsx72MN9y
L+UZ1fEwj9NKOORsqEAb+E5YOs6s/7wT0FUvmXvmPqNjbwjTL7wShT2yc65viAws
hqZeGPpyoMCwtaL9/Y2miqS1mqCUvTybmGIXnFvgflM+90v9Vm/d/oHrkJjUpe7V
viNZafd8DuJ/vDHoobDvZSBF3XHb9znioVV8Y1g++i2QWlhMn3fO61HCMBgtHx3X
R75CC8fFOWFalElOvcczwQB974KIU5VQA81zw/wgkU1lr354b4rvZc0Z6ADcqGwZ
aeOh81A1UlCJpNR5vgT55VvCmSqdPFSSmo/RtE27xh6yCHQvXa9H9Op0lKzHtExF
dn6lOHjuNhWcIeVCe2tbpSl1tUz9W/cJjfkUfV5Z8l2cEzr2Hv5iaygH6HCiu70l
YJ08YtdhWDOgEw9vFsqBRofXU7zN2389+IXqovo6noMQwoGiCWIreFkHUpOHSx5x
DvfyCkiKX1M3mGUvWB6bnuLfrCAH2xUatAY8cUj/O8A/CGOcvVx37yARqQZ+U2dw
tHXzCP3OLJ3ph/P4qkC80OOI+truq3YtslP3yG96oc5Hf5vyXhD9mFhUxsFUUbxl
aPCYQFwVsvCAx7pR7q0SLCiCpHl+dmckdC+gOyJN4FwidFh3FdOQ9tT4i8ixOoWI
FVLvQtZxLvE5anK/jRZ+ua9k8m4Ojp7xYZIA24nDQZlPobtkVCZU1RDqQRVWd8bQ
hlJ+G9bVL/MzrFAChibSoGOgkRZ/3eZLk2go9Vw042/aY41aOzdB5DV+QXBO7rpX
Uh9mnEiOxy9HaoC5Za/iwqXRXMnzb2e5/Cr0V9vwmpXZAwFG4/xox68N6ocbMAqX
GSpho+3F0o/88A/ey0SPPz3UpNKOGAHPmMrA5QtIItRaseRIYGALb7kqA5gCg38T
jgOuVw7IVAicyEddlgdHYdWFib1Z7y6g2BaqzIGB05PQ5T9+6VAQvg1qE6kPq1+8
gyCxpWKEJKPeQsdplkk2mwcpLrdv+ymDEWB+GRIYPDU/oLtTT9HHnAAyRrtDs2Fz
ju0I2tfZ1IUHEfUbZvqV5Epp6X1V8kSIe7PxM1mrBw137xG0h+LWO6MUcM9voDej
1Cho5E1F9FDUvvf9bJulbH4dWFhe94OQnZ/RYNQk25dCbgk9V/+nLGuL5M2v87VJ
FBgFFypob4xK3Heqf/LCPwa1MxH2FPuZ/0DCEL2zwmlikjylMpeOrlL8XolXp9xR
lZt0+qKQJwVGM38A9oGqOu38PC8wsWBtl4gdmobHWt4v7X08nydKfO2LYO5zMM0l
2YdoPvkNFJmqJRqjb9Qh9GjZQ2mWB9hvz75H6BPqpzTkO3kAydTxMGfnhO+cGN6+
WEvmawUGy+OkLyeJlenooWtaScplBNI6IuKjRNlTcHKakdb8E7t0NXsdBvU6HMHA
X6ptMUkaRJR42FRirKQ2GkfOnGKFaWIdgMvK494Z8CA018NGjzh7GVEmcK5PwUyf
xTLVh5Xv+QRCpvoMzYR4NzGTMDOMLcfx8PJNWmtMw9zBUZodWIYzwlgO4tD1kMUO
r90FrPRyXd6kc/H8gUo/jOlSH+0/TyiUp0P3RNCirwyTF4WbVW6yi2LQuLKdhmvx
sCKCX//KFa0R5XjhnAPbQpXuoUjmH9oRCFdbaWwCsEJ/UhGLVb9Cf98TM7euL6Wp
gZS/uyPoYCAuRDgFIasQul1MQll5Y6/0L0jP/PiQpkfO1QzeHC2YDcVPFZCR6/z7
xlGaSOfTJ3FmPxRp2ru1lcrw3q+U+Yu5YEXGJqLXhE/y3LSz2drF7EHuS9vLVBXw
XqIP/Kh15Az70LDxRzeVrKuRmy3GjR0lotRxGdzsJbRj/JDAdSh/+Vnkxv+6Ty7S
SI+sM0jfWqpR6BPcyGo4VhW6njPw7uemj0w14N7uIsUXipWQLAUme5BQY9mWl3DV
LH6KQiPqEqMppWqJXDirhg2JAJMjjEzFgqT9aVy9PzmDGeANSh4YDlSdXJW/7aN7
SU1s0RRZXU+qFVb8bI9+PjsMuGsO8MFw0wRcaBWsf8D3xMcv+qgTRV3UV9RQxPyW
TCHcR6Q9FD107mjw1LeSvkCQ5WYPNlasz4WQ4fXtL8xMnZ0aO9t+geck6/bxBx0f
LS+ufRmIc33vRuB95Gdfs8CQqXMRl11dvi+Zjga1ySM1rxJUSE3F2xsUhsQAFZPj
aOR1u2zCzP/kMWmP/s7dTI/HChmF9twne92fR+Cwy/Flvif0zBS+6AluIFFSpaxr
eIAVVO+1lndkRsbiNqDd/rWbBqCK8KvpA7kXbLR9XtR36zT2hTQXxjK4KBbJIqaK
FmQhQqSezK9sIWak6oCXU2cEqmIiW+RIY9urQd7s2GIi36hWHtxYCxjOKhbmblqq
v94VnZ+xqicyzFmWdDd23BBq2KhJzZE8VGFZdUW9mTDweoEDocHVVSJ+++7hGw4r
+SNl14GjTtq5Udye8sbHtYGSDhQKyM7s9SzghQJqLdMWDfqSi8444KZv1kXywqUX
c3iw38dcEjfXT72TD64TcQEBKmDiX+SeudMasfePmux3oxR8GIcOXCHZ5C5VmuWH
hZJ96zrT0tE+Vn2MVsdjJe74WkP0CJG152axAFWK77ltXsDMWbyhTTGvz35Uz507
VQGEWGOc1TFH1v1JTzrVEmRoVPxU856BE4LmJV+AvFmddYl8NAm7mvbsITreUcdC
Irob2mU6hEvDuW/3pwcSrWxUKgNt1lC4nlZf7qbaVZFgtsS7c+oHCrcwXTf4sF98
P4GmcAfHfGPt+guevHIy52gS8b4v8c89mIXyFtI2irhodQY5r9tW7ya6aMuoFZPi
cQZakTurB5wdKtA/+hMaXg==
`protect END_PROTECTED
