`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tud1t+GZZ7V40cr0ZvFE+MmZ4lpzZlDoeoCTq2yGf0tb230xCUklkDsfOGlu6I1a
TZQ45LCpUNw8wI5h2r7Rnaqd5/5GJXeDTfVUoWyhHxzdlejzuZsnmGqLM286LupH
vdYc0dxMZVHxZ/bHcZKL7O6LsHNRkABx0NGJm1PNAeEM1Wd/h6AinLn5ymf8/WHS
RyY+UW7L886bcNbYKUoA3vJQP11TRp6sM7Cc1O4pgUH1Vd1+IOOHtfkb4ZQyxTEB
1PxxUabs6992rfcdjUN5WxjweyP7eBSUGMxYGTL+jii9vJ03Vc388sKhTJFnEzqv
8/z5BbWG1EaPYfaHcBEjZlIPInqEtKetwh9rlraGkvFHhoQLCCrVvLL8JhWaxnul
P/4xNMZZOD0FIVQEgBprO9cQuBXAeBrZD5rhRzJvXG/W/pYVQg8VIRPEw8MN1ye5
LNSJ++HtFxzw3j/sSKTIyv76koa6WQILIGOiqKR4+Pti/hIxQ+BLi6b4ZYQPaxBt
23x9hp4/BvCyl6XvFEMhavxUxelGfZnLXUfMFhy90IkOqrdd9ioysf3/6HSX9RcV
LmNbWwmS5suFTkGdZskZI/f1AFTX7daIx+n6W6dwCLTbKHIIrDsx9aDK/1r3iU15
bzyeDvsPuplBKtDg7c7FVyFx8IWFCKiFmHFZ71trTBJw0N/7BJbY6ccFSfdNidNJ
Y6V5Qz8waAvB/fa3maPcnddg6zZ2XcdzRxFT2U6MynfmauIGkL58qrkqD+j79RJZ
ezfpr5xwnsoTDtbpr/9kbBmAFvGdEVquw8EmkXXLLWr5Tm+unRr++ZKvw44CXPx+
LYACt2JGqoxB6yRJDXbkTuFSfFzsBusof1mh/KNuT/5sPs1IxXztALx8rgW6K10V
UBO4yJDBSLergJ5jai5Ev0AnHT+v2Zv3kPCGn+ZP3sv3QwfLp1G3LNsrjWIk1Rgo
ayqvJRv16KB0/EcL8yUEINuPYqurSINNWkjNUHLNOosoZNJJD1iATO9cfOgzuiWy
06TpTTe5WLmndlDBRNH1NsjTMt5lg83zTeyXJFDlIm6nfpwsTGbQCMuWdWcbzymx
U17tIfrJGPX8rKkf9xylZTVVkyFzUGPS44ayunczAomKCwzMREE2Z7JyhO6lKufr
miCoksyDMySreBMkmTlaCdppGKZgn0FGqaHUSzwe4g9rUscndWy4VaAC5O5nKJn0
utS9nWgzyqTeV5T+Fd1wZpoy6WAH70mJWZVcjnv2qxrsL1uGMWn8jIb+QhuJkC1Q
zXJ4M3ChZeiTHfZjYgmILbqcQaKWJIhabmgG7vVaWdp7QnCy1+yMxjO60VAEso9J
pruBY41pNr+L+vDWd+e9eQZwIxCCqGSjoVjYN4U10FL8WV63GKKV1kGFVcFNvSFd
xv15eZg/3er8bYTpiLxT1BD0JgS9dUzPdiD8AuvaCBcslu8fMTOiqvICR4YGIK3a
wMHokUcon+F2mgmleyQy1/Db79JlDb3pIIA06mq4H0NZ6proV5/PlQ2ag73I6mLD
/QPEbg3XTuq9+IS35uDh/zajG+JVr988ggmLT7h3b8LiqAgV02fbNTPg9Cwb/pXH
3nsZ+DcP8485wZEpAQ+bWmTkWG5PX3btH2+lcibCSDJv6/WE4bnsyGrUGshpkmzn
/lNV2P7BpSRQL16y5CtLBXB8UBzKH/qkEkof1hwoRPAMnKR6AclmEHm3FbOuq+hS
LUuH7mBfhJSWHKJ5MMag0wPT3Do88VpXjcdjB6paEA+mTIWDY0B1yqErQ0P4XN5q
7c4McQwZ9x569BCZnQsBBP8nqWObfE9zFCKHrYzDxKJlvsj0jVdcZYfn/aHznyeM
yJyDlFcnCFVAfCBCvC+zW3/f7TWQP1igJUHBlRui3y+vqMCDHvnCrHj2YXZkhF7l
OzkPFUp5Vaa8aZdDVuUnfpIzA2si7d7PUzWwqJDhyv90PZsDfYvT3pzply0CqzZT
xSr7JljsGSADBNk3kXbCY/JtsLbAplociwJhvGVBg+/wohJAMODfj54CR39IiklW
k1TwrCUbb73YZGpwY5Fwa8YrteRlHGD/v2R2sCmbj4MWn8tF/YKH0GR/XtUNnl1n
1o02UAN/Mjmq4aMxjFhevw/K20ZvEuE9XU3iATC++8ZrmFwt9or80c5fh0PeH2v8
lxeyvSAArkzji/3WQLeEwiruRV/nx7GRz02oAVuBsQFl3f9mjYctISgiwjbAl2Ho
F8sMPXLdj0FadIbRPJNRbHh2rAcunp1kO83BdP2LDVIFvw/nNRTQ0gPL+7hSchTz
LTZyGqMRp3l3yH6LsUspD2s5pifDWmY8UZq/oANo9JNyHfgQ23Imcf53U6HThq82
f3mwwN23OB/NtyRdn7e5tSy8iLBEcWe5747DSjXrR1zKZCA4KrSABhi6YzIeoXYj
y5DWuLrr1z1GkZJrEQnsbDsNrHdO1kSNgqG+c59HEMrklWn1j5r7wquKiDJTGe9d
9nAxeuZUZPUYZAaecSEyXdkqy5KS0uvP5fGcrVo/uTj6IUXEeG9s8oQJKtrRRlL4
WUEyub8TCkM7JpE1HkjTMtJ5rreRzy4HU8qMhntia3VZR5c1XlUFFcXLKKmvWmNO
mxug5XnyTmX2AaJHd3PVaj1c6dw8JMAj5nRSSj2HwvmJRoeN2XqPDTJQYUoNgCdw
8tK6QggrEN/Wg8apNqZEXtoNj+WmQ69on+P05x392iONEWMMJW3+hOKWDbAdkDfr
LtoO9VCroLBOhSfu/1ZNQgY/Q8sSZ8kokmop17hjrFXUIUS6ZGbfn1yTX9g4vt5T
1bIUs/Ttjj9xpKxbI9QehtNHBV9mUqeV4mzIljudtlI3+0Mc4yLP9KistYtshcgA
44Uo9oP1K/AjcU9HUNH7fpwAp7lNw9awHCsPeHxOP/jHHo0prEfv4UAtCRxT1cor
mV8t4Ps5SEQ0xOXUgAldH4/sVk1HQ/jRL1NXpNSt2WHYTrE5P821GUiIWD/LQ+Mg
+9suCrmT6ZwwUYEmOq0AayWDO3L5bZU/h0IJnKNjnVhk7J3RMOyZ6UF1nLiVV5mx
Na3LaB4H1C0IxNSaIcxwMb97n48VygqajRePkF6mLL99eOVn4nSQrcg1OFscXY3N
N9srO4IJF0XIeR03xs1v97A6wrviiFEAxyOM+iq+7E5eTO52Epj/E0F8cJpCKr32
bLQx+qizvV3sV06MySYbq1cytHanfKqZC0LAx6179ZMEYs6aSK7Jlv5iNa531X5q
`protect END_PROTECTED
