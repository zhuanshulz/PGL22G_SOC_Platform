`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qHTbJVfdXbYXxdZatks8vvJqEXkY2LTUZ29IQ6uK7L+7vkLx+NOtX3CA/KoOykvo
TkOMwpDKeak+TmYyYusakTSrgyrKWKK8QJwZsFRX3aNrg4p9J4K/xa6HYgKAmSZ7
BVq7wifVBKdnnCHhXgaXMTTjPYIa+REqb4d4Z/vTIEqXaWCostwElylVaIGQw3mC
uoUBxQlxISJRU8wm7bOqT1ZamKI+VUeYCG0Q8sHe275dPFhDrKlkwAQdFK9XFzjN
bjn0zXsN4m8ol41h/DQmLQ==
`protect END_PROTECTED
