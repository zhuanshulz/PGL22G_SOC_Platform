`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5C4e56PsUKr95VuW1CzUAKsBmnLAlqgbC9yyT3nvfzHnTVfPdimC8Gnpv5tzTeq
imr68BIZxlLPpi9RLHoMIOdAbrgUrm/JVt9RGJlF1+L3KjdHpyknt+v1F9OoKe+N
HdUsHzxDM2HvuShA1Nn+scm2COkjJyWKfJ3JS33gQYND92/+gHoBLUvflOD7KEom
dvqOlQjDBTMRzz1SXS3SvvA0YG/7sk+jr5YtKW99ob0Or5eJLl3PUvqxYXyQS+SS
xyVVjAnjPhRlL67r8vtTIh5Wj+zngY5Tfk5+EJv/BOu6vxBjIi8zrkPL+70qwIyI
dLPAMDHaiUIremU2x28ywUxbAaRWfeZEd6EEs7734UMqOzF5aXIzCI5gRcsMHGl/
6wL9iSKzmmzOsH51Vs1qEIfumn0BH3ptNtOkjqa7LfcG1jRtwWHS2Vo6OXPpzHW5
AN4a4RgaFMocymrYwBaKeOOxelVvLbfUYIvpmiKH60Yx1EiuuP32eMndEJ8APC+Y
hVNdJcmK5aTsaSnRUDSnJkk27Q0QKULx7j+pMdSQJNr9Oe5HSDRxbiUMmQsslN0b
lccdP/CU8a7yJE1Gp/GXYSCJ7eR2pqkKz1dGyN3TwZiq5T5tcijDHPfBmDYngPbu
Rl9lpyrBj/Xx1wJEdNi2K7ByRntGjYrkQPqF5Ovgp31kSGEINNTaQEp8/Jia4oed
VA3v+pPhDHRUi/dc+jypppJLMLQraMGzT83pagxgGwpWuhA5wjYBD/QigCzdr+a6
FvEYnd4H5QL9kazfztH6xM945FQ4T9LnmEpeGNarugsGo9yGv1s3uxry3/D6o1F0
Lzsm4R5EIBeieYu7xVh8X4khEFPf3JD1osk8IyoYF+QzjuGfesbbU3BEc1+ArHwS
t6SFPPAJgOVeOtWsr/Ik9ywGxmRBPKbV0BVRboWItSPty9EBdcSLOeyEA1qTm91V
25WZxIMlL2WMMj85qiZygXnHbJEyKVdZmHsNg/2BWAlrn8DKJC/tUlRrN8zwWo54
f969QYqjXFL4EDtCpVd5lCRMD25ntHDLyj3X2SnI8uFbPZgEMTUMbx2fhtzBOG9N
DT03ZDz/1n3j152XH2WLomW+13qlpO+n3hdYKXqzd0X7GTwhmeLLKioIFLrsdrQy
f1MmoaxOf2fipbGvjEejD6286rXqAqfL5MBHPQOM+1FitveLaMNlXO12bFbPm/Xt
bl5seTVzTzsc+nwP002lqiqaPyl89WYKTB0p5J5QjJIGwfkNQ3KamjbPWd9SVDUE
N7rLOiDFoSgRkydCLWcIMylQPLWrwmNdxK9fUphcR1jvuWc28ch82slvNWfM+aWJ
`protect END_PROTECTED
