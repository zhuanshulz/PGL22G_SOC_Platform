`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v+4e5LJknetgw+3Nphlw7c+/VupkUEOcBSrrEKK/HTa+BG1W2xfQpliPt6Dv+V0o
mAP5jsD+UswOEogn/YWsWtK4wClcsv49ah3UlmA63b977THVBy6zGVwrpBeJMAfO
D5K3KZG+cknDGdMYvBBmr6EJTC8Zq0fcLkYjYJRhcfjX1EjOLqnsmbc6NUVCmdzi
5XcdAfSmjcUYz6VaS42HbidB5P9HY0HExFUrPonh7EVU1yUsDkQ7dw/lBD4+1KBY
eMFI5GOKjWd0nkNKGX1CR1M/SNFE3g2u2UNtFdztOtt3wHifB5+Y14A7L9SQjNHn
GfwJaulwM2p/yag45JCtri8Xj3YiNfKSIv/ZymtFmVsa5JDllo+ydxX2xDDlg258
sUUTk3wsClfZG1/r3zK2IbrYQ1RXr919UyQI6YiJDOzqm/5ANS+KXpAfyMr0Uw4Z
clGI+WQwYbHeB5GoZVnwoOORu/2q/awX380kcx9Wqi1l4rB2IWdHYVoO3tjvKorg
SdzoHCkLtwPYRe3Fpr1/vnHgohctsYOWr0Og9mE682kXLxwMqAPJBxthaCvcJqdx
R4H7iZ7vEk3NBrxly5wR/xy8/dE8Mzp0Z95Y5gm8qqf6qyQNKffVk8tuuIYhbRRF
xbYjoo+SUex5ikmU8pbD7rYltzrEVvnsZr8gh6bMM4E2YuMxbBx8gmP60+5wF6K6
QIE33klr5TXkT0Gi9fZWYVLPu2n8frYtPcWFdQPcuWiusTwq4wnjkdDqD+LoocGg
w8brFDn6oOM0luSm8fgdIKd1lVukYDfk1C1lMDV+pNd4KsifCgPb2guJAMO8VjyG
dWtY6YSeSvoEw9cAYp94PsiktFhy95v9gMvvDdUfuoCQXLERVhIZoOxMxIx9ryqT
J4VylI366jGKVlQF3EktGIkcKtV4gC3XfpMz+B7v0kyXK1doFpJKT6aTOtreyb5U
JFGQs1TJHGVD93ZcrNIuXOABCPtbjlkxlqULkOsm3eYYTau0FHV24K+lF90w422t
8ErzwO4hFZRIrhvjewSm7Gxi3EkuGDWcyMRJQSHu5PLxMHtzyqMzyxtBH3z7wrEL
MUzfGATLKyyugeddGT7VC/XymzHY/TWAHshC4GHPaIfNMhl2GVKC9krP2rrcnI86
MpbGbKLlriaXW+knpR1HSZBatetlnN5i5AqAjv8siwTAo05HHho/An7aniK+Nk2Z
4NjMGpoYVGLSzCMl1YsU0k/Afv3thIpQ+nAnYpOwrRpBVAbzKmLHokQB+MeQ+4ib
7x/fJLtaxqYcJOWm5tZv39GH8FWELSQOYhER/6ooUkUH/rnMRw8AzgmiqFDY7NH4
f4oI8WcauX6MT0Ap588PqxE+3+XdsEl/9MsaNBNETN5+L0haowRKVvegrMiTZXc+
e+EApaK4Fs+CMIHPazl+6B2V5eR5wvaQjp7H/hBsNk/eYIx0LJwIT/7kQpWMdae1
IdBtC3Oi7dZJVZX8C6G4OXg4tEEcINOvrF5qhMZjRgjXwd8Z5yQdM0PxIsY836oH
gaq96/RY1yxKBDwgqUyA8Z4Lj4f1Ln4M56bzGzTKPM1kNxvfBbkb1y7Gxyp4zfd7
aYdEBN5fvVoduG3H/OXdyippNyk32d6dGPQNCAEG/GnQIA76b/bkr8V6CX6Ju/Sb
KUJEWoSNhTSQ0G32XnfGpUKspvoTx+nifCrb0XBU7vZpVRPZyDCp812BQNzEZTz9
g3w3ADsoZAdxy4baK9hCvfJh446fwwXSzwp1LYJLIC/3Iwnp93LxqI/Thz64Y94w
ky0mNndzacDsrqJrLeRozNb6omvKD8Cpa4ncsNEuBsJlXTKgEUuTLD8hl4EvhGTV
iGpW2jQywu9POpxtO8ekfCByc+PJGQalBdeUMgktpv1lanou2wiWm5uCfuaOXBAQ
VqWrfRLTppvFWzs3pUk6KiiEicqgg27+/r6Zxz8/gRBLiF+ESYaLRcKlmOBqzomK
K2CVDvr2746wEn1V8E3S572zgD/Vm+u0mBzYd5zMRzge4/GD7NHkqdHYy7W6Gtq5
me6x1FPv/z1QQFBwAy+9WaOwY/6WWmAu4z3x+KGsw61yr0LOLUP11cHQTBDj8bgH
oE6LdPNF2zpVqNBXX7dGPyvyRc0bjXaahRavaGL6zeKQNlBI+ZeQnCU8D2f8X/Em
574GenjKIa/niiO1lan73DLFrbDDx0qdiPUBoFLaCVI86PDmVJNA116udst4ev+W
Jl28EKZq/xALO557Cuu7FAMN31AnxN3xdWpgYFplwFlMWlaI8UgYxFddaNgosTek
f/tZFBMCmflsAGMxO5YrS1QTp9Uhh+AODlNiOds9npUmcsK9nW7erOePW1jFHwSs
V3JU+gD9b6o/Gx77JW3gax0uvw0VakSgiaRr/NA7I72g2vRwpnG9RyHx4VnLzMYi
fW+peA5h3BT1mn+kLy4Q3k48p2g08twgJws6kYEO9aRFQ/iIM+ap6Zhk5ko9epFd
NI4COWeAd2UmiYFKx6ETCXXNFVUWE/lpF5Vi5eJXZjiHufPHuYv3F83BY8kZUKd4
tJSjxTALnd28iWMzo+Grs5pei0GoCMYeS8S9DgQ3asHxZdELbQC549/Yn/aFjC2P
TdiNIelHsGVR8+vb1B/BjMEQyTBVlKsg5ilnMEU/eXQsO9e49RE2YFFIz9+dzVGw
oeigIqUv03inlWe6QBmkj8pjOcZrR9A6v6NRyvHYboCW00zrlg4zJLn74cYBmG7+
RVIpAimnZwrKEHiq7iXFMpGK/1guGipJxYmZKHlOSnWBQvuHLy3kGVX4ezZVhbpw
afqODc1zmiF2nOd6KoA8GEFT/FKhS0ADMdVmqLbEHdzdzfKkLsTgMbACTftzVuax
xR6fFQJwQYakmNxlU8OtfIAVRKNJgF67UuuBD8lCpjmU2ve7SK3jgYQCUwUukew8
QAGXfdKUL6b7P9BzhkRr8i7R8LF+8FZ+E0Q12LBWvOpDyYBsOFOzrOS6iAAQr8BM
5yvFsQmy3byyFyjrNm6Uy1BkeVO3S/Y+wAqwMi9viLCvfDwEZV+uEB7xGJSnMI6b
c2KO4e8zrbdzZnKkioiNU49zpKY9ZsUXTH0nxAtmDmW8spyD0XG45MpWWyn+z9Bz
NuE0hP9I1Yaf1/LWa11plqGfKqBy6pDzWUWO4O10oeQ64YwNb1qhkErYFr6925b3
NEQMpX+HvX6oh34Qn/kiRzIc2HkAtY2nmKXvFj/BjaRG13818Yl9BiMyJhVwbbpC
WRq7ePi3kSSo31W1qJOgiI7mIfhtq4Vfp8finbpZT5ee+7ChOPVpH8p8XJQEV9tS
Qcys8ybl2SMvUWyZ3/iQvzI5ukYOvN9maFT8nCPpqO0WC7eIhwSf9cDRAPzFH6LB
2uHkfdfeWrCh8H4ZDiLrCgVRJZIECImlOVd3SxVqqBMkqK3NHy9n8kkLF6ANspVv
v09fkJ6jDlt4DOshaK7tbvHhvLP3VKBZAlVGhp0cMO6UcX41aUAdVxHRILQey73N
PdcQ40vuimTs+P/HKK/n4YqVK8JK0fXyAIPYAShFwVZOPzu+hGunjl69g/DknUAr
6kgXmQFqjlUgbTw3njLwtGSzUkJ2rUgffqPvWdWz3+g537w/CNd5O+8sN1Y4LtjZ
pYRoadyo65Sjn3rmtFzGkdanNuLGq26l3o/HzlHKSrGF1lTX4P35xuThk0J59pmW
6ZpdWm14pP2jS7yZ2dkzmmI5oZ+Erq2c09aHllPrtA+CwaRBpY/IQg9BY+29ox/m
b+OFICx4tSjBDn6wZgt0qSn2CfSsVPJFXwGvUfAWNjX/dQPcoW3PSSL2x7YJX0U6
mQc7OrQkEWPN2oOzLiS+m8d5HCRpN5+ZK+sY5MPWw0PELhXQN5J1e/e8GLom7pIa
NslA/x5lyCuu7B0/FbaUwD2ZsyMVNoK53M6pTnRQUUJ3GzhMYh9JBlxmoMrJYkos
ogpanoxbNnQXQj6A9Emt4IAGzqKvHG/ul1Mh9/Nq+VAIv9JQFmNISmUju1rXp0d1
bXo9RfAMidemYaHQ1AqPjyEhHT9eUqtu+/ByxgC5SolOSLaqSj10M+tkSLpVGCmf
4iHXuebve2dAwTPHq95UhXhEEE4ofjGC+XypW7SbQb3jWPOelzH34y5yezk1ZxOn
LjGE3yl0C1AWr5zGJmW83AE0jVy81i8Fm85gFelmevDpzxM6uHYyJR1EUTtiIUQQ
ML3QAoSy9GVmkZHBk47Tyh/T6sT4Xe7uOaSEiqCa40KMfMxGWOzwwtS/RvkoiHP6
Hd/v20TtNwQMRR7yivEcjhHNAKzMULBfAbGPoDj6MpasA7JqZmW7bNF6dKF6p1yp
Ljf/RrTeGK0jmMqGY6+UoyEHzhsZvW9jhLneicRkbggcd5nTNfwKRpFJ80FJNADW
0it7JuMLhPGg+Chop9xxiv71mvVj94sOfFlm9/fEJ9NUlOSsCT52COjq88B5BsSw
qukMQDxO0zxUfOV8knSOaPya/PEUwRlaOjGVOyq209sdOXPH2OzBWBniE2AZEuhg
hMtSJCVrEnx3w1ciasV0XcIyu4UQaeY+pJbca46yWG58XajMzNQjmWZA/+xNqPkx
xNtmYMqhPDwv70MqWjjPakYuVF2j/A0+0rv9ThAvppxLHqNivChkMofIbdSL87cy
kPsHXfPpiPFBgSK+Ra36XtVl6JMu5s9fKnMPxYZPewfvVVGFP+OTvk01e2l9BDYC
hD3Lh2Dgyd5ZStJH0rSC1MCFVgOitcGDivPmoMhdvntFwMeoOYxD0zRJI1CbEO7O
SqHBOJVOuXNglw+eB61YrC//txjQBX0cAA9ekEebkdUPsJxQhhQcL82YtAr2KVR9
hRfpBWNU0dgyBkWvS4eElYe9NvgMl16Otdr1LiZzO9gM3k+sxp7gk/bn36YNvGUV
765+y6hu2vcb8zNW12Xsy8wyXFBefQwF4kIAJ/Bo/4WdA5DJIvNme9nf92lXtJOt
zU02NovkRRWmzkGq5TmgMzZ3jWYdgRd4qW/gOHPEs1has6L1W2yvIRULWPLtWYFK
V5PPAO7w6K4yvNe1MGBjHAdlT8FbRDNc6qgDj217UB4v8WHz2+/rOzmMEAVHqjgR
eefrLrxO5n/qyL7EdvkELk0idIs4s7xPFH1GqEeeBMKWULQIirPLBKPBtU/XUtB0
/JadbWjyHLNUzN1hOZydPXFm9oJvwmHIDCvYvm7LBSFQoawSyfCPHnVgtIrN7jqj
Oj22lGiWedWALUlj/RLLxPHHpb5Iay20O7OU8GD6HBM62wM4j70OaG4pLS5G4N/1
7/E1mFC5M2i21peWS9GjDc02ZxJRV3pnnsHYU/qP/7Cnq94U8UXgoz4UqTle7Gym
u5QKKc2CauumNgORtm3JuED+OtJ8GARpCPougMhGULhh3d8RYNoQ7xg3v5YvGc6N
4Jy5Lub0I69JDnS2jNPJkg==
`protect END_PROTECTED
