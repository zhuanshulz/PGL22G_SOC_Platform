`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
goOwAucfoC7pVnxHlC1YhOP+5lltZT67b/VvSriaiZHOWZO3i4y4bXyvZ9yMLkJB
LnDJtQumlMm7aafLqhcH0sjJE5a/0TvCUmIMc2M4kM14mJU3pKiuXsz/3VdCPhe2
UBLR2bFkeCHNK6HRGgFPc9LQgt6DtzaCqfYjQBeotDRnFgUv2w7IhVWWRqROB8aQ
7s3niehmC34EROinuQcup2Jcdj+XNP9l8FXrmyr1NvFgCzGXUs5mwga1aVTTbZcK
`protect END_PROTECTED
