`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjSdPGmt7vGa9UtUMizeWoM6ZCPNYym5EEIW1Ziby+A5vA1fJc54fBb++F4RFHve
OxE0upWCZg5QHNLr/HF/oTBcBg0Yg1hoUeqeme/nsM55a7QaMlUaM/5ohDHmNpBA
cpm0O/N2o0w+Sc9lVOsGleamUrfFErIQjAy3ov3pYS95eMlihmWDcJfOce9KgKoQ
Gedpi3Qz7uJzGqkaW7gwFr3vmIfzXKj8dkLKHBi1qy7rv1mOBzuM7Tp4SNvmUlhv
rB+UQQr57neADIi2Bu8oN0GwWZ+hnYZ3Hp9dTQEO24ESaoapgVY7u+LjgGbFODKE
1t2sXXgXoqrOCxz/ugKqjlLq2UBt8+XhHNbfc0MuiYn2Lj9222GfXnMEBN2nxk32
X4rF3FjX6Jg754/EgWLCAqHkfKjEZL6FUzBfcAgSWppDLY70+cWAEIvaZEwTTLhd
R8QDCGAv+By5/H2dhOMz9UoimZPgZR6/RiYZxarfBx/noHKfVXLBTOF5EBojXIx6
o8E1KnKXypPEzi8pSEzGnUbtRG+hRLAB+TBbDQHkfWiYiiEycRvJO704H/GkMpR9
CyndhBNJMLdX+RIYhNNkPHLDw8IVe0+YVLW7LB6PYL/qe1PegAKE0AKYgtGtQ7kP
6B12HQtxbRCE0a8+rGvIMktYbYsVa80rHv6w9uFhdFjUuvrfHjDaKqFFjuV6Aps8
UdxLGAUcvsVBvXDs+WtwIjeRNNd5K+d1e7Vc/NzP6lWQYbvTNOP1OZfiBb/8kruj
2YDRV//hFw8gIyMM1s/KhtdYf5ClMBTclZnS1gz56wo=
`protect END_PROTECTED
