`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KH4qqJoPyga3Wk5FQaaalgpP4WvdLeaNQ26rk2WI3sZLc7KkCIall1LCeQ4MHYMS
hGvBb38KDJCg7aahNfHg8E/Wm0Y009op9JCbqN34hnkjm/1oVX2GReh/yntq5kDV
rZ6BomCeg8Or4kwfII1lkO8GnsI4GYRoMV1N0hsGL3JKcWTCUvFLKZ5JueSyNslN
Iw3WmCuXKVuDFqM0M98/HRM+qt08XMAYLF3VaMQ8r6yRaycEQhLqQhh0xkhRHrMM
Dp/KY1xQ3f2Ys6xjEec83q4rIFof8iEWZTaSOYNzcGbx4xZTu0cD5jMQ8iLVv4zo
vnedPm4HdLlEquYQcUL0U5owoglqw6zUn1ns24vuboq5ZHuM2ylPAXKWj2Z3gboq
5KXJfm3RpLZtJNWheWfRu+Z+uAGNDHXcpkA9r4f0VUTwfhc4u8xkeZ5Ga1OcjolI
qBOqIpnl81P9LFuRAfvMy9uEWZvq+l/vbypGmkZuhH6EtS9nZaiNKI8fbyTnasQg
5r0+dBVhU6BreJem5SyBKFeFp1yBgvqMkWLWBkmNSvH+DzSIxk1F1doOu7ZghPLA
enlgJklX2mGCaZ45VO40tCNfIIJpeFeT8y/n5qPUtcPYY6I+kMOiyU1H+pTqgUH1
xc7g5CdhK0KEmzfjos6tLVC/uFUgYFkcChsGDKSl0kQSYIftu+JPAGV9Gu5HYTER
dxPmQqHlgTvgIcTCvMEBZO948PPqOXZLV4bZFMfm4BmJvyv0JNjiZ2G4zfRoHrEH
l4NjXgQHtx98D9OMytZNOxQyFxQeD0W7Fk61RNZ8a11c77o+1+sVTwIEHu9LKzwH
4QJCyvDVSEyT6tXfZ9UnXkX2n+2O76eLQBH58dtaoezyfq6wOdqC5W33yklIChGl
nB6XK476j/rAAW+NiCsjwzfO/uYYKz/3iXgRrB9elhWRpy3FyvJUzU7Me6RQjHDq
aSwCk5DbKceR5Ue0VP34KHnD2+5J860mNPyLgMOd0tjwOG8b8CeGoz9of2K0BEkX
eMkMQSTGFAqVIk3mkwX/uu4lsv5qecGSDU75jGnsLOrqjpP3q8h89hmarUUgPu2A
CjNKLd7wKFe2dR8BDI1XQGQ7ctiiWVIO8n5VH+nqr1L6eLVvTlZR9bT3Ys/GHK6p
wkty/aWXIvcdpvwpJ3ff36FFS4WPBHhXp3as3NwSif29KnwYBhW3Abey5GmFA85I
I4990oKgZj4XiGkYUm/Ibqc8ltuZ93L5oAH9kRnVxlbNO96qKQXjqMTjFccH34hC
j5cj8/Cs0p5meRjYphHVr+b3c9vBRhVqktHA9LPr8ubS+/j2a3939YB3BrPSPoUQ
pvgyVmyDajFMUkuI9YkCFq8eEOcGIwRubAqdH+p4M8U4nkHEwe8LhqesuQJYoheX
uachQz6projPKsENGOhQIWGPvzkPujoAr0chnUpNrYUeV7KVDQUGjVgOusKg28p2
gb0gNDT4VW/Izhh0t5/DsB7vNpimMzfHhC/K+pOkB72cYeoy9Ixv8G+vqTiKxyEE
sTRU/62C19ePutfQwu17Qzi2Ibut6j6TLFAWzInMRFBpINvRapAz020j2uB6PcwD
MWXzxKIf5Su50tgZgyn1ImvcRGBFtyPNRvlyhZh6trIpcgyz2xYSmxoA8U9FzZZB
9svy/IgKTKYfIL+M2r9T8oRdYvQ5Y666alvbhAEAdswhTT7SJI4tTpzQGoXM6i/E
OkRLTC7aOZx2fmQ8u6xI7LgW6sFCnOUpRmsJr8eTPYu5DpTU5xzqKdIWWGIAEmQT
rBJsAWfXQ/mW5gTBdt5KXwvZXNnuEOkRgpB3UYgrhrtRmt7cYBC1LhTZRZb+kv7p
5I5uz62gZWQDh++gUVi/5MzZOBI3XtFnQxV45fPCquUrl/ufnvLFvpgGCSrQ+BeB
EzPEFcqudaVH7JhKJlYIT04QBwBAXRDze2RpMIOw0VCmtXk8E5/0tdF6sEAP/Gew
ygBBkjCC7EraFn+6428rLMuB3H4mMhhVhmvalFLKmUO/2zXpIFfR9sRaUQmi+Meo
ZifjHdgwfra97ID8fEPbW0uJ3pkp91o1pBQHdG188ytQZe5/BqYUZc8LmsV4ayr6
uJSI5GX9HIm2eEh4/f4nx4xFqy5RBTPgD7KjnK5YhpqbhDcRxCBljrzBcI4/05UP
+FDAb0jFqw540DfDWBRGxbFmf6nKE+HBAgk6Zm+ylqIUmIrbNTn5nVqx9LIyDpUB
MBgjjOei1FAsWd3xJDYJqoZN7F8Yw02SBC1XcO1qLL8636lstjERg/t+C77f9OUL
6E6Vn2OOFc7cmRsh1ZQqskxSHJmIzsrFQ4pm44TOeY3W5O2CxE7HiNtSP/XErDUj
pMOGdp0sQt+2X8s5ILsjKBC1zD3qG/2ktKNrH9K/OdBt+jr3LuZHV45Hb0hymYOK
vgSH/HTtPWJ5vTXxEeLl0HxVIaLtkyZycwxLmz2V0sw2MVPxKLlqkpZtj3RNhEj9
cnVl1H/GHRxk1jRiSVuKGsdiqDqOtd3TSDV5f00NAGo8AAjRjQ7rh2UCtMvEtZj9
mTQh8rPOH896P66pIgD8BWZrd3Tzqlj9rrBqYIZy/e0M0t0Nkk41AzaQqAkOi3g+
1dYr12LfhdPyVI408X9CoA1StH+uyGTqhaQkt0Y9kGkfRCRs5Fdh4ypoqBIClbtR
RSsBU6+wFeUIEYmN09buer54w/8PO9Ua9Fe+qIgEJCptj4t6HWHD8HwzDrdQLMbt
sW9HR9ViE5jPPauCoH2fbhDKw8A7nVQ/3/qjABkBgCXXmlaDVap1eJnRr+aaQCaJ
tOm2xfWGY0oaWypTeaJXj6FU7dQX1l9lnwIbMzfRGQx6EeoEct75mhFgazdbwus1
4G5Ro19laM54nNnDBoKOS4xpN3vsq46A2n9C0+xAm6/hXYGdc6eZ6614iMbGNDwf
L+thGwVGcSxJbapryWTnTtGu/lp+4x7D2i84zsY469IzOwyt1fpVjEGvr2v7umQT
1IP9QnTF38d1fMzDhPkOajx49o85koc+ariwsxM/wLamD1gev3HP/ONcql1jSltP
2BQP+XX99uTOZFMDcO7XATbx2wsAqQubjyBdmIDDzXhDqtDvzP9eZPoOeYWqssJp
I4ExC+jdsl95pQc9sN4weVXKbCdoTUhpdaAjrvrrvkhPCsQH9xIno81m8XMNergU
0ZJtfIEGmDN3Il9tx12aG5ouAajN5Gm3eddmmTmI5NFSxJF/ZpDYmN7sQ9klnyN/
JCirKo+1Ww0nrZ5jXJS2L79Y5ljgt+i7yGgif6ZvizDdJAjY2AMbRgLoS4iWWxZp
8kCIB3dcipnZFkPGDqWR+HzvQZ6a1bm1GmS0IrejzaE1p6QCvh0LMwqlRZ3/kYI/
PvYXrBiJj1jPdvcyyCfsR4vqsNedc39/CLxqxkgUI+6npqAj5IKKYHEio1f+CL5P
ZmqY7JmyU3wRCpkUnwmzh2h8WwhiUYt5qAJMX0wDLN2moZ4ReUfThNatnRmvyGEC
MVqN8nf2X1npW8w672caG/7EJb6Z0k4Bq+ujpcTJ09T+LMDikSpk8yQ1rKq6QS97
OboOESc2X8Y9589yUvgYy3tL455zA6IIF9pC8tW8oR/uWkH9z48fTV8PvTLCZ9tl
pBGdU5JbgcFlQtO7fB1tkmoBPUbLi7MuMokj9AR7NubtE95Mnv0Kslx999kVL9Tj
QpoN/SPcwo2ZQkOd5bnkf1Ngj2kT74Lisy4HF+O2laSjMI0Xb4PQt5ieSxvWjXji
OsQJ5ISL2PSBZ04YdMUWPhjT1LA3XdGGxqhWaa7x7rusf9cJZXEASi+djvFCE4rI
0s4HqdMXpL8TlL59M/7BQ3EJBZOyfa54boC0I+3GH7C3kSec9V9E6r9ScfDeEIql
qEMLwad1fyFOHR9m6eGiCaceZ9YvGn0HDkTE/OxMkttUYuvyKRavYozSUg/z3/hE
5SwNeUZO21wNYhM7nKJVUcX3ESYJEl+wFljeZt20nUdGIIDlUdOjJnPI+Lc922/8
VDHVx7Q+zfJpfR5Rss4JosVj11OEVjrZRxZU9SLS98I7JsqwfHGyU4p1ZqmZp/U/
TjT7bSOaxQMVCto37uWMA5hisoC0/DRDAMi1PdUF7TMRbHr/e+/2fDIlIqYEp35s
JWFF5CynFXnO8Hj6HU0ZgSzdHHPXci7DcqJtO35HNf7OT2XL6IgpUyOtQ8WSj2LK
XzwGbOoW8jNF8Ue12afmCpsXCz0ZDWrXEXolMbvBNMt11o4kVoKRYAE0/bCbyk+V
wfa1GhWDV1QSABfkc7811LOVlVGcC6HMhg9H75W15dkDhQUhgH+hjj83c7six98j
yckoV0jfkqW6Qvh1WwLVNIUj2S/gi91tghgR106Gw8X8UT+H95LSZrD4+WAROxlN
5H7JLpJ6rv1Kyl4OVddsyXG9prVlP0qSTBJnZ5YOS1Mkh7S59Foqz92jWw4jnLPI
yaHPbBz67HTokfTTEUTkLCmtOzlP2bSltJunWZBx4j5jKcfSMsysdUVyqz+E9hJi
wPKEz/eh1TXI8Rj71m6raR2npKJ9lIsjE2CeAxyK3ehEVVi3I/+/0mjGJ8qRAETi
iGAEkixXCgI2Zfha6CnfNklLYh20WtZaulnNxpd8KH3Zj2m7Za+V3rubcOznjztY
4lf4rn0mKEIN5Bi1Xg+gKqTHsg9mszZxHvO6CHAyPkSEXufSfL8iAH9kFeD2xhtg
dkwxSgwGndZE4maB8jJOsGckTV18ZK2jqHXMUZ8bt4wK+z/S0eG8aRrcqYNCFzSV
l76fdpncvGStmvWnlMbQvgajj3spYhi5Ni64xxCq6X89r4JnmC1c0CEYmM28ZgHh
2CjhOJKLmVQtlvOJKXuUhuma5gDBDgLunGicGEpVMYRZJk1PfqD7wNtvz6ojgK+k
jchW6K4aTS9XaSPOq1yFdWxK1Vufk3ltN5VaVwt5rUADInjmJQ2JOTnXneCGIvlS
ZTSOmjDK5tu3PG0xCZT7yFJD648YUmR0Tm3/hv1FAIfSTfG8I/1WRUPQeAqSdeXU
ufMZrVU6Hzoz9zc1Hh1l1nef0fyrZ2Z6SQ+gp6QSPNeNP0d2OfIFmCQm2ELXINwj
2jkbGG3WMZ2pgz+PDKUjwhMq4Q3z+frWGJYWHeVxp6/XlSB5Qivn1sp+3kAH/kho
zqZ0pjv5QXVIlZSsWYHu6GUzQow8lKET7PKZrcL02VhQbUsgdG3ifoWGz2suH81r
IWqSCqnblZms2LA8xfTVmZVxHSaFKj9L8iwuK9KUCaQV3+PkebBeHDH6J9rpOw9w
iRIHeZXEmKZquiiIZ8zKSjh923mHMF+sb76a/OVz296mgy6xJDw+ydfOYYx/0QGP
yntlE3aQvRag+Dh8RfWWBkyKwh3sWez8Kl2xYbm8WIIsgnAafOmCPj7Kd/n57FrG
AX82+Lm/yG7OpCWZMZHiaPCEiFK+l4ridUbiXCUpiH1r223KDqgU1uC73zhBZQj6
CXna79EmzzQaWochDUt1N+j1O7Qytb+N7bZOJ8SLRXzKu+ouXakC5WGpKvAXJgMu
f1tBIrOLzaax5rHPb/zZKBA8ecPa00KNAJNQ5fXihQmlxo8PYFYMt+kYdDMAVK18
/RFNUT4UCWTOV1kwQycmcDKz+lpJWZ/6slwctOCPGcoi8aJ9fJRsuHfYwLd2iBcM
bMSG06pXRvnTfU5AB7yrHqNk3fjgc6efz9nsvUq0YKjS0wCIVnjS7x+Jh8sYVaXF
VBnqkfB1LOExrXdIS363ZgxxqcUdqvYMz0/EjnJuBDvKwmcHsIPD3Iol5YK4rLbF
qjELYQA7E2K3a19a7Uv/yR6z0UQBQixILkh2XqNUMGGs0Nda6GkhJz+LFjyfv3L3
npkljBWrNVFoi6ISU0rXlqmI78P+T2T05b7O/OD0zxC3yndA5mAWlAAYTmjaJlYe
Lq9OtZubLLZ5bmNirKnrpMFhztd3OKFWkZiBEiCv2E6UnNPxxySV8S+cRCJX05dM
K8DIIydUZZz0xh0ddxq+jpkDm+izu8Zfa6zt9liazEbpCu65wrKz0jJ4e4ziP7Cr
MCNyrfM0AHJaYqZZZ9zvBIcEBQ2xB/OThUcGDNf9woeZkofl4cAjZYOpZBxOFhfn
x9c50svru+Mf3FYcDgB5+gaUalRfwK3vPYzEjsvnooctJRNVFZoXWBnkEE0fWF2w
XsITy18pqrXbiOn8KlAdC+H1PLoenOMoW1VPPrPJYJYQxbl6635YbO1vCngw3LEK
KEENUSshVGnlxra20IgI0JV3ZunYCbwHB5nP/lzrnGPinpAPLH0EJ5JKHj9IAeRl
t1tDY2dUIPtKj6UO04L/vdPyZIDagUhjcxXh9MZBGEWMqxm5F8m/47b6FN66lSOD
4ckNUBz2y7YlhXbLVzZmj49D3kBzIgkPl7wOidY9O2xqCicUdHGtfgGO8HT38HLz
xetsRA7uZeOeiwWPdXSSqCFS4zklkhVvRXSh2WhyNjJKE3TTb6UZKjGv6CRw21ZL
MXWUZMNtVf7PM5f2OvFRZGVkXV+3r3JpValzEARADxsaVcPNrhMQbvE+UMaJIh/o
fhi+HqQEM8MrNeUdIF/hgEa6yF1s0UwFEAjsnN3PTqE0LBCs7Rm19RnfYh8bATRy
CCC2pQCauW0U3K4Eur1bPCxZcUgsqfR2nDSAg20NG3SZSw+z85NOEEpIc+3dRizb
T5Gj4Ey95ebk4D1f5Oq0fg8AOQiGvQtomoffc/VoqslIaDaptMmm4jhGFJIJZmBN
PcIMrBXR/WRlWkncDseEZSug0aS0+Jo/ETy4G5P6ffxN79YW6E9ZT2/8FmARj72m
zYc0PjokL80gCTdB7PhzGkDX+Zv4HWtH/0bEC65P1II4VE/eijbbEzuG3xrQu8t+
Zmq0vytshEquEEdmh2uE1mE3C6kAaN6HCqtBC746YHzpXCEI/JE+MC9+SNAJKx9g
0NmIpFTX1ILyeopjV9cYBfNNdI1AkUM+9df2PXz4NQ9TfjkEwI9p33h8hRCMnHo4
1en26nvqJ972s4diKZE31XyE+UuwB0QYbLOzA282kFipbvTtov7Vob3MbNy0y0/U
R6D2k3bbdBxIvKCv/pd2ciwp0MhvWWM45lJU9UokmS2NUKLg2ORE2HQSFD2NMaUY
7Kpb4mpEJTXHrSfGgpMwEzKzNdB/61QjZfYZaugoirZPZSZz+QWIfB+UKJrqPHwd
frdECQUZuHoXFdYZrp1o5Wd4w7TcEAxChi/2purWSPmIxYy/NC15EfDl6CzySomx
M/fu0o9yntDNaOuTkzve/MSfxJ0Ow2aNS+KD3RQtm9Bi2Sf6250R8nMCgZF5Juog
5pEYsner/popoOHPdmdGC8b38dsJkcgRRjrrweiOF1v+0KnLYaHWduPTMW0c+FZL
FVIKM8Whgi/vQT5l7szoQIVPOahGmAPp2Xox2CWa7inr1gURqhYdh/F3Cf4mf5Ng
xbWRpULXz73F0pPvN9N1+QQ7Kf7UzbHoYLBBUdduolzmJxfWzw7a4K5xvvD7amdu
+TWJQY/5+4HXW4OeEKEIvD9bHW0Iv0kqF/Mhy8Lx40Uf5PHnuENl1AyEUm3SAEwQ
ktxPnQX5YV3Jn3Z2QqvPYnoraVhUI3c+vIiegUdSEVYcNPx1uJ5hxb0UWZKZn/Pl
fvBty0slN8afpvqPxksWCJIor7CP8rQ3I4ZwDbFVN7Bh217VSQyh+OK+F0ReFNpr
kynVkNBfsK20gMqNUZ6P4E7se8K6hnSN3DP8Dbbwd0tVpVDQv6u99jM7E2Uv1ri9
/ARB8G4+HkC/9FgLCEPZGqnDe+ZJt0Yrcu1cVIS+Km0EQvc0zXM5lSGrRIDQ1wxs
p0kosx2PPuA3IIgEG5ZN5H2Ym0O7fZ8wJdDJJC3aYHIB5QDiAY3k+0zNTTPDSST+
bwrBmSjVl3fXkOlSnNIuWMstGswCSijc0gy8LuAJTwyyJp17KZ914eCs+uDjTRA7
55ciHFxWp3XtfGmTsTb7T7WgU43Ld/RsQy3aSaxBjzXAuu6HITt/0jNrmPWTx+2v
LMeKHDQPVocENL6Z/63NljVyhf9qsI8gmzPHKDLYro5cGB7jaYM2DIYMAQa6Cr4K
fPrUWBQVCKojW9n1glf1TR2qKh1GTtvkYNaLbVtQRz63JvnPK1CUaAApcO9zPNA9
W2tg0hwdFSq/G30NaaIDMKyb+aYC9f1R4Dgbm+08s6BwatKmLxzOBCI55BhmxM4J
WXnvDu150FVoBfiQsEzMR3HtGafnv9+gwrg7ZYdYsuUT6twaFb5xk52YPrJ/NN5G
wI9UeIYLe6O7ddjgatfZHB2GRm8IC4NGVzLoUO3i+G4WwfPQaF1Ka/mEzjWHz5A4
qgqA9HueRle/PQQGqEB9hkbnp80tACvK6yjZMXX3K3GqMimvEsE92+4YTKxzuPOO
64uyt+jwtmV8Xe+BG97cAi0WhqEIAVVnKFpT726jNOYmo4cb5RBTgDG0mJYIRAPr
+wqMPVsq0G2x7hdTri2jIWTATM4E62lr1zwhsr9PSxi5mINZ1mo7vdY0tYBlhQFd
NV+PfF8AOxInlaPTYKC75UeH5BSC+uwBxX8jFiJnKyjao1Isv6hrwpUpFOYfyz97
HUzL7KuIud0Piwrdx67Gr/X5WlrdJivNxfvsJtz4odehKPJtxZxyI9twpBzoJ6C8
lB20wZ2DrCm6+Pc4ruL4ei+YBOHia1bE1Vxr7yyUuzIVzwm0oLaFgh7rr8oolNwQ
1H7UvfVARstRwANuXgeEcN/MIZaDJN8Oqii/VZ3l+WI6yGpW1rbjOPqfZbQfWkS8
s6tUuVwYDkS3hMb0PQdM+SIRDOXHIO3ZUxoio5gJkMESW/D/hVBvF8kkSZ93Y5hS
TJXI/cj3ayRRQuD2o/l4WAGtMg2dVQf4ScR8phtLiPTR2p275upidYmK+fCPvhql
kcif7kk57u/SOrF5qhIJnpMQEDauP2KqN7cIcqqj37XH7M8NDA5Tj4smhGJeo+MS
Ve4RH62A6v+zaJVVRXbLdvfAT/tgMFanP8LigMsLvvzTwKS0KXDRBx15ye2iDPoI
7xTbXkqt7LurSXPmVH3+6CPwNXMWUJD1qZxNprs9407zwAEGKgVnst61hVSSDjC4
Ft/FPpDwgaXq6B6HOTabyF9xsN6/Oq3k90uXaJohHzKkv9OpIKHXz2jLAySOSmkg
xAxHSNj3V0ydqt00jRClY0mAK/ECj73vOua1uE7+yuz4w2epaZh9LmZ/3eEEZh1X
8rIU5pxmvL/CUJZMoiTPsHucKb/CdpSWoSWM5ptR+hOn0lHzaNq3EO5C6Ukjs9PX
AY8aOCoCRpl+S8bHkIlOlT09zUURhsuVIuHpXu5DYAYth2wItQiF0/RR6riD4If5
1jDEtCiBE8w/bzXSF1rUBpRGc4uCxXkueCEMnbC1lV2yElehm4jEUqL0cogFiLIu
o472Hy2duyOgKhnQcznysamH+zsV3EdBcWTur++6XH5QTmcQMTMpqxmjoh91EINs
OYCo6HTMhBGjXuXINH/502o92stPZnad+G6bUFKuL6M9EcNJFD3oM8ZYHj3FwG94
zxWhAD5+dGv3BUPYYEG46Rg8ZO6s0q3u8jVp6c1DTje/eDwkPm4ZRh1Fgn6ZHf+m
QI84n/TD8T0RNrahadg7mDlDSJ83enn8InBx25stNtq6ausRaSRbkrPf0QdXcQVp
9iPRDEc3lmieRkXIl8Jo3QPBtGJGs819w+KsAWCu3j+vSmK9p2qAYHlMQ0TEpNG4
U/q9vuQJQxNKnUEJyWWxpLlIX61yuRm+OlU6wjNGlO2Dg02b5mtAqsHi3mCMtx1b
Sk/ETL+lt6rrf2o9qssPMBkBvkfy9tW2W5/Oo5BlvO+x7qwPnNO6gGGlJGKKFXjX
amhKggTnt3f9O3RCbnia0hLj32IsuMSi7AvaSa67D50e+ipb7DoiTTMSDNTD7uqH
zpDaHtJs7sZQ2DnqESzw4G3hSznicTxU/jh34/Oox6YA5BqdsSBzgt+hlsUcx9iX
k32fUDYZ3hVGcDfMgcb2OjKqEHLNFj7NKJ2kZB3uLdztdgUrfx1brRIxtp8ZzN/e
aqE/d7xZ+EPicAsAL80Uijx6sG2nNlLotn/HCsrNMb/ejJ/+GN2VRss6mAeu4J4N
JRECPpp+fzLIQ3pdRXzTzDBGoRNBcCBGxlvxI1Gkg84mOvYg6lK1l9cQopVZp3an
6nUlD7psChKYzFZg406Dk6h6yQAFnnCY797C6Z6ZkFLKi9ThCVBlCzzGSh44UbS0
TCOv3a7ACrAaBg4U59p9Dphf9BeoZrQBTKsCkokBW4p3ThiU0vqLEGc1R40P7pSc
3NsDJXAiq0gYzdtQVIxxPIvlnMa1hj398spzj9kKAeGr3sY+ZWNBWVmg8v5Hk/f+
GUNUwdRW1Qr7csw9oY65Rt5nyCHITXjEdd7tprTGviBZuFcOiAEWjd7aPpa4orLt
mJT51D7atnXVby5tWAPTFQFF3MCXCSiSUwQnkx+l6kT5OONRBBzm2MKT1ZYmldP6
J4SuKYptt7s0C3UYJHpmn9Fqi8HrMypUFnxI/L2id+yPBFkY89gPxokMGTWiy1/P
LFD+GkicOMtMBByFIlDJiNkZP92kfgOwrNdA4QYXBGVKCdma1KgBjIBUJRnOhxoq
ppdswcaoDWUflDKFgzhMXn7blEwgBzYT6Zr6Ktf/sLAKpyYiJqwEOPwilKsAl3r+
e+ea2CsO8hSCHsxteaqNwonfMeYr10q764dp6lApYfgeKhI22kJt0xudjioAN+bv
CgBpTk8SRqIwhSIt4wP3qqipUcQDxK9HS7l2BtSreGaW55XlhCdEsmBg1RTzItF4
ZulTRLhljBN7cQj10hMd/1H26rFw2SwQOvj7gK6VWrsG2MQQvkbvW3KUUNSECJix
YHjrRNKHQEV5BPVIs/6pPEKr1MuSOhr5DRhpbevJrM8WI+KfddvcqlJnOsMjlqbW
tSC5EAvJFgKes8tqkIS+haFx8pBr9t4Ro86jMwfshPuEy4lBGOiWxe0o4yoUEujI
Ru3t00dkCnRONO0WfdpPUXj5w2CIDQqJOvoWqfm+5R8+jm6IVXglXTtbAvcrw60M
2Vjgf1wXTXgZtY/Hbe2qtGIZUuL4NNYvyRpZf4r0zjv85NTlJ90NkAgPMKlgzzN8
MWJEY/DaUCLnVIyfp8M+X/L4OjkTwI4q8XKGGCMyV8iOvwyZw/nSt8vZYiK6JR+8
ZO1I+0Ece2kIvUCiVnecnyg40UMCsqkdSenUnlHcx6YrEtSvhgQJmt1R6QUHpcQI
yHUgw4BucAk8+yQ4CKIna2D/iGF2FAZbG8n68XELhTO2oPo5enDJqrj+8GslIRkC
OiX3T453VwYFEJ6bExAEXK+c7gtJxNm1MncRdG3EdORm4GcXlJLbRu5DU3sqqjHZ
A+9CS4LffYWQeRQ+7RRV5D59nJ00y9CY0C6+6UM0kMtp/8Qn1f9al843f0DmM8SU
mqUfXQmbckCdrrntPSuo+9mO/7VVXGrXGu+vHEifu0lMllfvtt4zQ9oWlCfCflT3
Gx0Tztj1ptE9ohRLxo5nPmomS2jpGm8CSBZhJq/pzJSYI2aCO9CjO0gnIUzZuFCn
j47CJveSfaCZ1QmY+KYgAcCk6+dR+NlURdY3pdkN44VqSnLU4Fye6ccFhWIz8CIQ
5yyjW/QjZhmER8NpIcwes1N5vD9d14XYBHPA9YFAu2DPhUyBqFIoNfNOx1bFujlB
tALtySjtXXYH76mqph5JqSCBTMQqEdRFZAhM2UFNIq961RMrdYsxc7pm3HOinfJj
Hyd3qxLUx7DAmooZtu6RfU4yUMixKXigcWK2XnsFuMSZVW2+N2AjhADFQfkrpSSU
EK9Yen0YqrR1OTzF4EeeZEcQTxIvzd5WpzuniwFEdIzMCKghYSODvQB4MuWoGNl8
5UIt6sERwTD8EXaWiRL1GxZe3yzH346dB4j9HYkgbCne9vYz+Z/y76K+vBMx78c1
ehvBqbW6RFJO+8v1wTN3f5lEiVrIuLl/2AOilQoL25gE+CaUBw0qdFO4eB4wCm63
/G7mByjOuCSxrDGegNLWurh3NIuXIBFWPszXmmsyu6IM/eQ/TyourXb/P9VU3rmT
BRYNGxdVZSjuemo6dCEE/PapHbrfuas8DKMc3RBprp55OUetxqQ9Y1acZmjzPtZt
sg4QCVJ/rp+PGx7RskojANvSINzmY1tlFUJT5743uwsR2F4vVddDabaJHvnMEH6h
IbM2Kg6o1D6FYqZz9Hzgsk+PPbJADqLP0JGe60/zcpyyPx9ZI7iO1/0HbsONdr8Z
eC7LxWLS9H1c9lYg1lWRiucCeoXB0rD/xjc1FPtvvu8UyWxnzm4ixVloSIZZGS09
LJiY5No1iJUcjkItPIfm2DaG8kRxUIF05rpbq2cnxCx+82+3pJnCEKwyQfQVTfMP
X+pgwWW64aUoRgjLQQhw7xxyBPXCr1OUF/oXjjOj4JHazubUAdoxKDy+ZtiCPYkH
myfdy77vXZ+iLULhUqf/34P4AvB3HdXkeYWLVC3p0lClnGOE+KpOB9iYilvQpw7r
sJwubQs8/vG4v3CMT7o3rFvA20qLc1kPkHsDT8sAeKg+nYUUarATSHe5RlGeB0/j
CeIzqE9UVkMW2K3d48sIMkaIqEBVi+WcxGZsGQ6tYC27hSP/qt1+pDHsrkXwwg8s
GYbI0r2THzNOpqyDdz/A9rB7/Ei96KXk9c9k7PIyIjSJdcftpzNaBdPkHZxTp1ht
e4hQUibzUVxcws2x/nTwRkItfTrxawo24l3Zwnkp9PnkFNgjiz7142ekihCqKBZM
wE+FYTVp46O9Eb1axCFHLPGbZ0Ab7smJ5RHj4+3xNwBPSlFwwiykDTzasx4V3su8
8A2XBvOPAVI+mkdSjFvdOW+OLfCa3dinoxcx4d4PmoFoEQxrRzWCAHBrA2Tvit6G
0G+g6oTBfm5s3myA6Jr7/+vO7VLg6KOumJqvNW+El1Lygu15nzkDNQvuweogM6kV
K6DsUftlGSgjBJjEmQ7mn55UQ1B1pC91reaEGjrUDJ8ezzcaQFdIOj6olAS/VwaG
VR8RFy+dVGYPTPexESIQezmAnr9+snL27Efp33ADSjDfVfOstcDoNgFFrpX6ucUI
Us9mSH1BS9i6sjJNzkqnwdS0YA/u5HD08KVFUYc+jzpZOgF8yarZrEayULb260Jo
U1KcvDoxB1e89TYIIu4dQlB8bKWtI1GTNpV7BukYo0f6mTIiksTZbqeAhvF1XpQT
MjHQ+T0kCirwPnWab43+tWZq8ecMIHfFePQfB0DSDuLSbKE8b792zGn9WgrHZsr5
F8iN0mrL43mTuq+WvTdVbPPUuieJv+8Jqg8gpg1CFwHRQvJS/1+WtDIPVwKQeUAN
LmSSPSgFWFjRe4L0Y554nIhMOsWd6XsEZXQilYz5A46vv5C4N6XP2XKJvg2KebB2
68jrJLEmcrRLamQbBQdhWDvCQvPY1nBuR2A8EBfNLVaiDoJBdKMwaCmrb4B6Vp27
TC6DUaqBlTMjmqw2vbYmFkpPbU/0/Rcb0wJwtogvRFck4wecRTR2RBxtdYHav5vt
oE8mXXQ7Ve/sZ4XRhkWPIpNkY4cpDuYrCGSedcYBCM4wgB1TD9Ql7iXpHqTCzFN3
itXLaE6QcIcx/WCLOkmRoHrEN6odD/oL4P0rTRoK20LiHTtjwIhK3MAeY+u9hycX
5ePoAwSN0bJ1BVsamV9P2KI4V2EcBQN16JQveblvGV8c5w9rs6EVavYY89LHm+5+
q7NKq1SEPagXJnK8YZZ5HiniOVKJJpTz5lfoYChxeSJn7jkYFxZUKASntlIkgeKH
zMYIMBNmFzCcYhuWBlybNNr4GSZ+7eN1bY6mOLlQACktqBGFQbMqUprIPQOng4y+
Q6snADCtGM9/6h1M9nJX6n9Iw7H0vb4ftnHPfa7S9Sy41I1+XcCOsaEN5DwlpU/7
b087KyhZivv4TcQyAPg5Y9hHXkdi6mcqnfHkkBAzBglvW9BstrpeAJqn4TDamLK0
va1QRB07GR+o3e86wnE1nBJmn54sFsdnLGLcMQ5mpQk5DxeEr4zFKbDvcus6I/Xw
xZbuUmBquKLBALSI0tkzW1BQXCm8o9G8r4h9Eyn7rVn64PO/E5Ex8kSFS/yEmqUb
gfgJ3qGkr70OwHghS7kVlbinMIb08t2ziQY4DjYWK0FiUnDFHWsZPm952PSsEujo
pYJy59IkuYdQnsQvXK0YXJXnMgwmiLCbYmvNFN3tklAZv8v+qfBuQDVROb1Yc8ZG
rBrCfdFxK3D8paiyMarJJ9t1+fVkv7fYrhFmy/5jRVKIG1JvYf6jWO6h2HCZUhvG
8+qLQGk0RXj27TYJhic0Tc5FSthHwubeSSOtIvmb5eJpp31BhWUw0tN2Mob1yKHV
sALNfY67gR6TYYPi4jRNZk3ibW7RQx2m650e3fG/Hp1HlmlAQ1kUKQ0Dvcj1myMj
zdHnMu2W7fEsRkUXWP/LxhYXbG7hwtCfy6v1ZvvArASZqABZyBLBOHzJY448GeI4
bbn89WA9TO4jr7d6gYSVE0KN6jHOppZpa4SaWAt1fm5XHy5j+y/5kBMzA4pkpbK9
mJKCY8pPEy6EzvzQAintMkoZentxEqlH0aUNk3TBVgq6KNLwQxT+NidOaq5vAkiu
XarrBGTJksp1/PcOgPbrdf7wTjCj2tb7BYTHfW1OVppQoRDMHv9ufQ1j64R7XLTx
BBwxvxaluOJmDKxCnMOkXx3Vb+9AhQrd1Umy7F1Gxr3zgfibcf2ujuGQv2+nEPfc
wPURvgME9RZDhnB1dlc7odhRSdteICExUle9znn25kteyWNphGqekHt8+JrwhW1t
lQ/EJG8DXYjb7SsyfdqiLSJ70Zqo578cYFK80pQjEb5sP02odHKt8+AtQqKNDdHQ
sUUdFQAX5NmlJpvrCxfsl7EGiYmhatqH7LpvABDVnsH0LnbH1KQAuwSfYaH0QjsY
US5nTEPvoC8ARP11FDbgF+DLpeBGQaGw6D230CZruHZicb42RjhFpnsovFxi11TM
QFtH7dOx0EiNfICgKILJsAXaysLyoVqAH08/INTqrKZ0jot8hAFEko6GFjMOBo6y
O+yjgXdLUy9RaI/uHdHm7mYAHAib78eLT7fbt3vIOyeGABs6gcKXEDEak2hsDI3Q
Yv8MwxKMPYsang7jdYnw7QW3YjPRGjY0Yl6f3x1RYceCH1Uub36AajJa6PH9YzFT
3O5Qwo1IUms2p7i+PQ8+U5V6RoIgml8wpxCxerZXeH1jhqrUuzZ+cDvpOLdRWe0y
qDr3sWbeDs/RrHb6a8YVDo7DjBmKvJ5VRLXGTlkjF3UC9QLldPqTu0fsIOChi8B6
DiESATBevBgvJ3Y8/GXo9dbx85ApzVC2iBGfmb6A2NlPkLQ+BKe+sOoR4PMOf/t4
blWOOhVDSyDxG+HkOLcF6zWcXwr/lpflgeljkvmRUvdIYz+1hqqUSjmDBVljQTiK
qPIF1U1Vp5sSshvab0AH6uF0lCUrx8vM+VpSKyrLlfdSHv7PEvRA3R6LNj02qblH
Af/LPc+ACZGvZtdD5RcOG7u0dUagGX0+IwWbzT+CrJTFSeSipQAOTj6y4PsVa4qU
9k1DcYPUvCQhJZchxV0apdKlJxdL7HOGn0tPwyE5MM5iaz+lVxMThj30d/vXYckm
wXIA0UpIaG3OJQFJrDNcYMHLo38f77jrxS1o2NQ/PvkL9KxRj2g3g7KDtj7m1P+g
DhjwYzWOZpvi3mw8oepoargGbypO4l7lruN/5RgVWe5szwkwVQigfxBrZuMhDMo7
+qZu/MRxAWawK6KCBRNz14BCZmADLIhX5Qfoc6bbWIFVFk9cJ+g0chMf1joJqS7W
+xzjJoKCmWHYGmBQxvH1zUomQCKm1mvBvEFDB4jdb4ZSVVoa3GoMoJX+74UN5dSe
mqHZ55lL4BI1XM/C3cnU4r3FlMWjE7rxuGuxK5UimcYxDrXcmRcwN8qxvildHLSj
mPCJ9MlkKCNb3yQaHiScH+rq9P1YUPOpN035DeFSgXDfN6J0NvOv0UEi0Cj2V0ca
Q9nqXsLAvSsXwx/uJXKxQdGwqG0ajrU6eVDM9Zd2MFctrjA1316L88JQ17jUoy+s
0X7vcOTeEA45BfNs/PDRaU3eNCcubL4rXRuJ6TBqS+Ney1Wgdi2NtbJpmmv/uj3y
+cLjA4KE9w2aZmqJ7k+mrNGbwFNHLEpt3Tos8oyFb6RzpdZwq7pDfu72iwL9JHb1
MfFVi993C/HMmR5fd9D/kG9sIeK/VEq5Af85D7gyL9Lk4X9z+k6z5AVf9ZE9klNS
Z3zsXdw2VxMqNHFF8u9E/I2Pn1VJsaHpXjIViooYux03dq9LPfxT42F/CTFL3jD7
+Go55wTebHO+Da9qfJFssL4KVprBDc071sCDoKWtZYQyIpGu/kZ25cqndjgXL0ED
MDZdQV8+S4AmPWr3uM5udIhJ8yBUVGrCf5SuPWBivkyehGLt3MpCu/IppD2lXvXH
9DKnjYLGBSvvJ/UUOS+bnlm0AW9DVJeVZT8zA4qeZM2SyyoGeYhkjoM4hkfhEmQb
yIHVVnBSY3k/D5FInc01REAJP0kJf1u0ZFikgL1F5/3zlRgNIT7SMyuUG2uYoeCS
g2Otwlyxs+skWCwmZqR1KPb5sblOw538xoT7FpZDx1CnUe/bapNBX6yPwdXbDxoA
5NnHjyubtoCq4xc2sImkPoT1xDzvzrMGQ8ywtKf0VcIOc3O+BFP4l53h4Ed8j811
sCYLYowWgdNJ8aPXegE79wyFglaRK1YhIL5XSQ3DD7A+hecIe1iWvzJW8BXO/S25
gLAgmOQlXSLGk9tAC93sh7z6zE6qgm+a7vEcfvzLOV5MlHcTHAI55gzTAOJR6Fse
wE9whX+dwZE590c30FlPayCYpQcGbHcLgyWAu8/M9zNEbWNhI7eU8m8uOKBOYy0i
jYgfBFgYwA88/wSY16sMu7DPI6PVzMgTm4E1Tk3W4702TWxYR7g9mDz8NeMjtbY4
Q00Ej+FgEsPuTtUlCozVwlZaw4onq9WDejhFKx9v5GMVfkgVDYePJhrh2wwGEPxR
Cc8tmUvEFZpgQcKr1cdvyg==
`protect END_PROTECTED
