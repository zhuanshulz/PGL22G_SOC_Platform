`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8w013nSpblhJ3XzSmcGCnELmqG39mwi2qkaYPqM2tlUDRZ1qFy6W18rRLX7HfRZf
f0HrV5gJL5p4ERpRMmSgweSVGIEDyYm9glM8wOHWLQcFILhvkVgHDaI7ZvoyPyfO
DYRzou4+Xqv7jFyjh5Gj+vuqAr1biQcsAXB6tTy4F7zA5wAytb5zVcaHPs5qLLEQ
bxWCSHFKDunK9y41wYShtOvCrIDCe+kQMYDJubbE6ulrAg2TrwdFGHX+5ABbQ0zg
EPvWsnyFIOgOH4OP1QQD2uwVyr3M5nJe6aqHrZk+AqHndZnAlWnZLPdiCAysAh9v
wK/75NBc3UxtbRQh8ZDKu0ot5YpMeCOrXncTTOwdamHN+hBxSu6wfwlROSUeC3ZV
M1etVuUGOLhfg2nRhVtC9bBlWrHwp3Z7twdQUO85vBoBOfiUHhtZ5kKXFus1i1+J
2G+r+RZUgONnkN4acoTIqQehuxI+p/0QWuNzjag4Plhym0Ne2Hg1PDcpFzAUBlCa
7m4s/rXJmgD2pHe73OKMVFhlOVQyw7BxIpdrP/oD/g5QqiCeJHU/f6jqGRs/QEWR
MXu8Fzx/iE+nToHnAo37UEFzjE6E+GJ3WfCORJjwYVnCDKZL/fLEDAQpZF7DLBbp
Tb+s6UK8KUq2al/aMQ3Gah3cmJYKpkkOdXAmEz7kH2fmuNgVYu3x02sRcfKayYh0
`protect END_PROTECTED
