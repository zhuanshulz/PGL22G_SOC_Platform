`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ExrDaK6xL/RRPwvKKZ7H5M6sOMvsCWze6aFSrDG+Edft6wW/EWALEvDf6OdrneA5
7foCEW4a9gXWo1sxOv3OXGnb7GwzOZtSeX2pGpx9UPJyb+xaxEWCJGr0RA4coyw1
9OApngoeICFRJaESSCcQEUqgikPJFukY3Eq4ZBBDg6odH1+7A9sG9sE4tSFO9LJ/
XyiIbXU8orwUuvnQoD0q8YcQ2+bTDX9+SRSo6R/Nbwv3115lx3/HL5nX2RRTunYg
lYXrnPiyQj01FJQ/zTYiyoJv16w4WWl+RcBZwRJy3U68JsGnWDhwRHf7U/oum/VL
WoQAUgjQZXxbn+9QsxTR18GPRJyoLaQe+7phBJJmj/nYTdWoZPKp/rIpy6CA6yuu
eOFHOvp5IiULOrEO8WYGkSDUPF3hM2lfRsV156nm29MR4MuSp/lBngbZ+5PcY2Wk
iT+PiVhxdOO5cw1nj6cQ9Ycd03l1nL6dLtXcrCOq8GY5gTEEPfbKESxMkCh3RuNc
aWyBoPWtwbqtHibEXYvRyjO0W72l7fXI377TN5xqGX7xDlOAsiGQ/KOFmm0LJ5KR
tDgLKyBHQao4hTHpQsYrvqR6L3fJoaSBAEIjgK8W/MxrQPqYFC/8P6XnS+XEWwI7
mxOmUvfTuDdAdHmkMD0YyYWEqKY1BmT0bGc/FgYE++koyPtsxG7vXN44GQ5LWnXr
lh8f1bOd2/MvwzwHYCBRvaEBHEjQPy02ghpOaW18WKUiT4cTSAMbuvvGrhX79P7p
8pcc5YZ0Zf0Ec85HhtvTJzTJVh7YIBQqV/Oul3cYrV1IlBiz766m5LLbWifR5eB1
pUG6Rg3RFSxYaLWUGbL3bKxbXp73BKkJmFbk6TC7bYAZT2CX4QwLEwSKP8c/7bZC
tjc6rwTkRYM4Atp9xFQDKL6EApMehPYv5bNG/Jlvkkyh2oCCB+Xfm4w0EWxa+oYq
gg+aq5S7rKWnYjZLbmmxnviv/ypyV06TqZj0/0qgT668vrkJc1u6P7OkfdRoIUkc
4PU4savokd4AeREOUYRRO7W9/Vlv0Qw6dz96Aidx5pWKsg2zLvl+QVyFWKzbATkI
jKbO/9AOA+fT+ABOYQhAaUKj+bDsc4CsQ5OQIL6+n0M0IXwKJ0YyBPp9hJPTMfoj
nNnZmnwJ6AHqOUinc+hSL2V8nxw7wX1mkEq/0GmRs8yWVtLEgmLN6rxvnIKlcwZP
eYvQxDgGa71qLBsqTvZ+W1/d5j6fchzrmwRFmktCK2emvU/H5wfYYH92XxGebxM5
bfppWwL8TRqg1WtZQy7YOzuDV0g5rlplW8ruiXV3fycUKkv23UBFEVQn1rdvHezj
qe8s3kJsi3efodaDIUJ2G6xZKF8xv9a10aiXJBq8A7FjHYBDdPMTznhxHW8cQj5P
xtO2Cv3V5GRW2WFkYQoLpWvfmBCiuT0bkcRyD8QGC/0jEkGHppWRgLFSc5dB64+2
wF1Qh/u3w+b4YIJ3oROuZQZ/31UsZYZXjQjYLifsMSW3F4+07dBvOjaBubszCfbY
8EsOrhzEoikqlaDanqf+lMIiZlVaJBNiVH6u7HI3MCko1aZ3MEI02KQW1I1dZJMn
ZnzUpPjtHhLtSxBmqynWnfzLrzK743aXgF57xqB4NTJX1XJgomLV2UICqZAoiqQQ
4P/E9EDM4AAnHnsgPKS2MXjO+PZRmIRdLitmD9oayqBS9LSfAIkV8g3xgh7JOs/A
numvHBiyjlI0bxcVIGXnC2KD3vkCjB7I/G+K28k2htwFX4hqnwdYdkPVZ4Ds4WwO
Dte/r8gQEgV0f6bbhzLMIyQblqNJiY9VbBHXqam6x8fmrh/J9G0yxpqNjudyDD7E
Ysgq6N0OayuAyltoMD1JTGOhEuGy7Gqb8oNSzRAiL1nFpLkXQcx7sqxRxKyRhutc
JKpMLvBJZvd9z9AyGHXjQzGyJG+aeKxAc4I/hRZUW6QjDjvO5DGxWLuVcVx84ROB
C/axiAgFXTC7Rf4Nb1838udv8zkAVsKVTxE6M8Mmis/QPhvDqsx+QRGL0pge+OaW
Pxj5FG/GAUgCpdneO1fNLGvZsHY/ErbC05vBwxm4foh+MVes+ABCDrpqW6fz2ShJ
9XM65fuRi4MRWNC3lyFis1+sEWyho45S1pehFOabCtPa17ZZDHoZsK4z8wHEFw1r
XqjMU7pPCGM920yWOt5/b4g0yVj9al4/mBNGpZBKgpmFZah1cO4AQohBijCISpuc
ILubbTMvWAWjsp7LDa0MKQ9zx828Vz01UahKkze9D9QyNSbOyJHl7ENd+Y1ZkUVh
Rta74EMXIuPLrKzvyIN2bKI71mpnMJXhrgYggAk56A8ryc5tOz+VT/slzE4cRp/P
4jCkZEmTQOmoKGN6Alr1BVjfidcu/SUIWMF+qcXDKf6UyrXyjEFhnvcrKAekVEdW
phoe0G9kbIW/zbvkaTXVCgOrU5LUplCg/u8GjBLOS7vn/DbQa7+DgpC+9LkCyPxH
i4VQ3ajZRfeivVebY19gps4yHR4iJaZ8Aertd0sllvM4ddsKLzut+Zl+WWYXp/nI
SQfWgUCIB9wxBNQUP4kMclpBSMq7zqHS0ZzGHGmYCbJ/j0MMOwMhb5xk1Kfyvfp7
fJxrfcD4iYrTsfLzCuobpmeG3zyo5Fn+gxxiEy5Wm+lOJsxbLnNq/nXQV+Tce0Qm
WtFhtQBGXAAhW6JcuaIEj4bfw5n4ZPsJ7ckQD5G2YVpQLp314uxjIVLxRfukpUV9
pp1XmIY0iE/HVccFmMczpeYAjxE1GktErCRI7D3J+Kk5e1BTsNf5c2Dfm151ivpU
0eKqp13M820pNFVyavULFLgtpxaBCPKKokn9C6DICCsj64UuQFRO6KduH8peUcA4
h29IRBNXWW7s3ngX+jJURAcpwvruPrDf3CHlCAGulj5IOqUfWBiraQ7GvIZKo+4/
wpZyEcCASa2RGsklzSgogyJYUJc5Zj+Ozbk367tB4memPXFjNF3bG0VvcQc8qyWn
JSoj3R9M4Z1gt1RPk3HHIbzVv9qaBL5+2HAuNxC1dwLlDCv1LEC10E6OlXgo8m1A
gkwArIro3Os8HDyr43zpFyZ/CxQKGMqUSkcqPsyvkyGLMFcITcENt3/IZzLLOTo7
zz9GzSGZra28oNQ1ShJwp5P7PWsEgdAK69l9bbh8lS1I/T0EAtO4NWqOUQOZ1g1C
C5fJAMFNhd8xyQAM6x0zBp4o+39uZucoDekWkqstEd4WxPK0OZNSNOsMcLYaoZ7D
1UfJyzUmAkHiaRvQw+knYCElgWt/dWqBjJ4dzOEaAbAL3dn+jP6+SFHPnbAvvYrm
hf54waCABoOmnPssv6+TkKQ59BmTAPBH9brjc0C8glIxYeHkXwF17q1aBCj5FPIu
TH2lh1u3Ifc+FWE7Bd+0s5UQ0U4PQRBam4tI0eC4NoAENREvd0C7lb5H5lZJaqgC
Qei3QjUcivafGZoYJBUkRqQPeUfNVO6dbmjnMjyf5S4qXp7t0thxSokb3VV6W8ZM
DtPEbTDGl5UyUYlVxpyn/KO0YAke7flcrk2zpg8T5Jcbx23WI+chG1Bg2y7NIl1H
l3rdHcsWB5UFFjPB2DfLf+yAKibSXZZvzyADzsqiuXaBy/+UJIwdCid61KRcELq6
h8+gnkAm3afWcf72n5y3w+qSf8+C1JlW55czVff9y15vWlEFQph4e0+70Zptejgp
X8Qpq9vM+lFZodU5TWkbLoBIjAnbb1HUkHJBimNJ/5XXO03XogRiZ2RlziZSLLrP
6ctbUxEcutYLTgT7ZMcN7d+7tuLh5K8OhyShx5i8TR4dUV8e4I65TzR4C6smZ+5O
qPukPB53v+FKCDK1HzNgKQmtnUVRnhecRjxSuSLO0zw7ocCNKY6QjkYehp5oiGDo
U/zCv7jpMiAHUt8eUDl7d5Or8Qo3fF9wfXowjHOBU9NHldwTYndZyLeYGjpY3VVw
x80olmcLyPOCmE7PaTNFZUDuMw7onD/iIsb3Do4BYZk9Vyu2fR7OOuJjq137PmvH
B9OYwXv6kT59fyzzhJSBU5OICQdUqzxuF9pYOrCU1PZY0aVfGePQJ4Ae/7JSDNGd
n3JAsQHvBwc9c00EJe5+CoYYdbRbLdaEeyT3wYPvfP0tmgIVxCkBcaOBo3oZY2DD
oIh28sqY0pAVjuFOWXc5vUG4rghwlg7eoQ5eChoafiCvy6nJOdhjXxVBrNWgsgwe
J/cQUQJuyRPRE/P2wHNayeAJgyHXXFbcKqnHLnbVWJaqn9MZTcyKSDZAvHZEUf+4
fBMKwggAs8BB+VsMWRNDEUt4znGjc+Lny6BCLzJoVTRslydDj+b6lS052fFML9v0
Xy0Io3xR4PEy8hkIXsnMboDxeZDAooS5Nm8krpwtPWF5v0dvYIAaOgM+zfLT0hzj
14jZl6WT1xHlEZTTbcZwBH+2B4lhNucI0tPbg1IkoYF3bJ6chSbm5NyCbIP9RlcZ
7R+nLSfmxokR+HQhsvmMNdTME+K9t3XbuxIn7RaJd+DVG8w0raGUqLKHy372sx+F
rriWYxCoNcpFWVe4C9b/SUCdzXeA3gL9UW9Om48DW5U94uwLH6HaGY39+1QGKpjF
YNS2GAq47z8QrcGq+VV5FlhiatnhS11J5FhDfOkyC6m4q8J0GNAwY1JQ0eaD3iRW
w8wvN8S3EWLL71+br2Mx254h95tvuRp/ineFkrAA5ombk71BoagGCQ9vGifW2DL6
NTN9HR9I3nDOmyqr8z0HmJV9M2+xZussmdlETwUo3mbAEUbvirEaWJxvr8epaJAn
txtIClS5rriw0fhKSJV03a8aYuaEGFqjl7kbQhr6Za56Tk7uLUYyrk32KftrhBm8
CViczAx+q0HpkGi1CeCOnpHGgbKngIl5ghn7k4at86IkZyCsdx9113TimzaVjV7L
0PrDTgDZkx3oR7OfsB+Q+XU8KPbv4ETr6qNJALMWzgn2jwsgF5aNfOpdDqa1IHXu
GHm1EDyKpb4GC2k5KrmW3XMDeGHN8wKr3sasrM7GyhWWQdvqbaN4DEUwVZuRlx52
BqPOSGH/Es6eRJTLNdKyO6c91BQ+mGuoqUxELCfqGY3/8TpGPGarQiydKr5St57I
ky1T1VjWdJ5GuG1B5E+FP1qwpvLZBDMqWQ4VqCz1Nzctc7ldAP3ecaTc/GinwlTk
ijXknEY/halUr74/o5z+G+M9fjqQC0a/aH2nbfDV4Qv9/Dl6DEPrddhqXs14Kn1S
pZa1s5PKESDkdqk2dxfKJ2GFmlcNH1d2g5ww9izrrMQ64Yvye+z024XBV3x//fub
GwTWO2obU8wl/rFoAQrggYDSjyRWtwHU21kdxBPvSBZpq5T0XhzUdidr7+M1w6jS
tp0jW2k6ivMLteTXF+R02Copsiso1jOHQtNAIhgZBhbUTMCTwFoT/mEtKfH789/b
N+6xYVQSMqEuD5qr+G/uMsjY5nwe7HcwMZwcTcwKmFgUDUYHhFnb0jOXLkYnDrFD
IrGHIdmpaSfyYoVqMOZZssp44sbLqJDQKJZGQICxilczpXN9Xx3DqMj/OB/U0k6a
LMIPUWzoKPF4Kvbtnn7ovDo7QY7WxpVDvHYeMQID7nk5fZHQypJj61sY2OqEB/Et
Ja+lEeLMWEIG5//T+C3lWORau/gM9UrybQU3EleQmBfuKON/6sUr+E8+cmy/bBle
OXlorFLu5oz20Ext3yXZ1O4GwMBmsVjo+qa9Tcfus90bi7LuPXKHbLyK6RtLUJC2
3kitDiUQU1qpVAqYRkmO0xTjvpb7YsSnVv3BXn4XTwJbQvzY8mp/UhDxRuskyty7
dojKfVifntXq/AxZHUyCxQ+mvC/lIIKbC6uJLqKMrUTgtaUzuLYYHpJADKfth+y+
sAn+x01c/bzmWeSxr+N2AZcuLOGiGNPJuVjFk80uZ/q9JiGUq+3aOiMaz2Vpp0yY
2rmat5+adwbFBhd0TkxXizjr2m58VvvS2QjN9PQZ6F4OnITNa/I9BVMpdxpuKnGX
mqoSniLJTybRUg4r/aQocPXLcXHjtQZWHo8lQ/oaf1c29cwzGEnR0wI5jxMx7YOy
7GbDurGqt9fim89UPLLp8Gugyw+nZzC21QWu8e9qWkL9toUlqLCOYAEMi9rnyEIt
sTIeBKEyC9mhXFU858Iv4ZmcaTbjy/kGXiLMDJJN7C81H1mYN0lmdSLUoN+mSJUQ
0MdgYHdKsXI8y4JJlG8lDeoGYRfu6zhqgTLk4QjZr2q5rWviDqXLLlcdHHWoQDwn
M5YTRqsWE7LpR5Wb1jrZroZHB7Tq5lpqugz1rkB8bKwfcuDykRD+9gmD1SVmY8Nm
XyDX5OddjXEVvneUzfeTZ1q9H+dfKJFOOMHaVN/8RkMsQuW+wIdlFVaYoB/vi2BL
uo/JSWBOwENmV2VpnzkNchjJylgFELCAcG5gwv2LKHtOaRx7z4phds2Lg3ARV0dQ
2W01Ibp4qBlzxB1/LklqILNxMbVCQ/iaSjbfRwYIXGOpqlCHln/T8v2kOfcb3D2r
jgJM+9ph66LJXx5UUipwRHFsPqJGSfqJaStzPKOKVKbR4UpFdAGBqhbwPF15hLAm
OAWNbodSTQtkmJoViLXKFP5E4QVG6VYT/G+emeCgcjw5hX+OpR7zpND0cb/9NMXS
S7ynKtOr7L3bJLocZsGPUZc+Lyyu5iOSd/oJRZHkLC57oKY91aAnA1bwTDSSHSRx
8kRAB/4+kBHY1P6sXUxrhDk6bx0OqVTRakyfxsQTdHmc+/ETpVOrd/QOiTJsQptZ
AOcZ17t+rYPUk2fvKftAqoV7HcbdOb1tpnJNqIPwReeTMWm87DCZOk0Om4RgJVfh
GIYjlB+XBGSOS9KAqa6TW7oSNGFftDi6Y5PyZC6I5T+GQg3PM3zqIVnE8EJ+1Rf0
iNojkIKrzj8NO3BcaTwkgyHXw5ZkaPM8y992dilOsEGM5J8zec8IUwigEbMhcgfK
x5JypTmTJd5s1OU4lcWRJNwv4chEvZ5KsqSvHhyMNt2MiGwJF3JzNCOCqHNARVTz
K5s+cRlGoomkQUdUeDBkDxS6zSguEHfhd1nh4tBXfVwVFUTwWjLGhDhlUeuRXutL
7llyxp0Pb7R7eI77fJgc+I4gE1Bk1rtmU6l5odgYBV3t/ZxUANGs3MroGMPsUagX
vQYlqkrOoDrfttrt4UEfK8yt53Oz/AqTY2yt3zU4JLgxc6BS8rL0rlqo5UfKNm+G
s0gW9QL4/Sy0wyUoVjqNxWMQ3ehstVcRcaY+qPJ5Qz4iGizIVrnRHQqgNb46RJdP
rF8l2Pauhxyz6mquu8lYpGnABdJoFAZuAG/qPfvQBSDF6m29Ud5Cy8jwcpyVs8AG
lsKbiamA2zHYanVHR4xwYmVIzUTzDJm+faQG1LLPiUcqdEvvYYpBRbFLFvDoiKEJ
9I4niHYui/Qt4zJKgxhJ9Bq6/pw9plWcpBxNlXZtlsZkYSO0hWDz0x163t3WVS0M
2b6Jhs8eD6iB2/FruL1vRDmwH9ku/dpbwysyEJavnjP1RLOosYWVRi1BYaY+zBeO
mP/ko6S2wU7j3xhLvL3TPvOVk2ttd/Rp3YO5ognTctePD80mA73A8P57civErHcB
3GOlUW4bzv+A31ItR8cO0x1XkmB8hUNP8GvJU5wzaO6L5dU+XZ9+q9LYMsrOTkS8
IMFF6rGJWVDUFFu72BaiCugIsRq7qVstssmmULmW0kItRaaxurYv4Zw9KV+GmGQd
wjUf/K85R2og/TV01WdX1DktqoDs2iCX9R8cvzhEdnlu131Hmymc6Og50FVzawYI
XkwKQT79wi+mCD3KsqmAsp4BDoRHcy5BzoN+aBHbeXW9fqE25L7K+OljusLudvAe
YEMA1C3pOQwSxGMDqCR/QvJ25B85kVB068eVBoBlQ6uYj9Y2MFniky0gmS1kCtpp
I3Al/7RYf2Z0sJ6fwLvzSXV8orqWEj/0hwi/obiH4Faxtcz6dWLetoBwm6ViRmn3
fF8E1CnSTZpS5tKWf8R38gM929todH6vxT4qEgw3YAReV1+qbfY2Dh1b6sDLJZXd
BUk5cgOa37XnvqtyKdH/j3d0gZQdtqxucz+myKRySZgxJgYOPfD4YKd4fGygccdz
WPJCIKuwJLneGbI1UulTTvBnILLq9Lw2Y4Sk9c1l1gNquUKIxTLRXQm9sqybej+k
5/VlkOWYpR37Q5RXQzDUCGSkAAwd1aH2T0YtkAx3QDuNMKt3uqsIWNnSMi4MU7d6
LMTMUQkPj9GbRNVEhNvz3rz8jFiKSboIh1YT6WZayQgtG2hKe/7Lu+2jrktpVc3Q
4XkkJUliIZn2LeK0W0MmpupdRZRixhjs1vt7/WLv6pA1ldHT4QBXuLKXwIfbbP5v
5dvWwROfdnmZmUqZI2j1pY8KQ3xeiK4+vu1ubfDeEsVeqgnIZvi5Ah6se7WR4ZuV
9sVXp7LrP2pjrJa0DiU85DM1fOE/K51Nsf/6zRIaTnbhqiGQjalOZeNQrSqjKNf4
fw8saX2kMn98Ks5Auk9g7V8na+47k+I0SJ+wD2aZTQ1RUn4vYYUBq5dgwrN58D7i
vl7NdepQauNLYvt64YYt1fdOVFx7w9XDYcNjXQwBsFFd0Os9/QqRbmXtYqi2SXQK
NvSvOfInrCBryQ3r4RXnwrkwa13O76+LHkKrMqvbSS3QoCXbZkIj58Z7nAyGf9L5
dtKBJ9GSMiBjiScWRvmfef5mB7hFWbIxm1ZMQV99G+SZUvdu/uNV05+CtiKRavdJ
HLTw3q7hvvRyj1d+k7K+3P2t8pujO3j3KmwX71PH0JIsAmgWH2QVooVePbFFwTMj
Y62awMUTE+yG0KLDBnKZQ5fXOIewFmqYKcRUMGTfdK+rwghkjpRt38zIInFldV7w
vXjj49Qj4I8B98d1tALrBIv541tTpyjcKKVogfFhLmT/6/k5WL1SDYfGeADNW5Uk
0pyR7RuHPs1EJEjmhMzIDzED5eLvOktUqHx8VJD2XaONcIkYNJI/GI/sf/yyPXNB
cewhJzL35l9sIs95gDPTkYw28iy0q4LJIp9puIjSLRRKBeCVtBBZ2hqEsMttJkCD
A8uUHlS6A+76NYKOcyXF2xuR4r0eobNHnWObB7g4dAfUa2gBOv14rbjWJ2G0kaxi
EfM+A0OvExDwzOBzCJegWqFVJojqJJtWGJclZRmbAt8yS+g/Hori9B8KC8KhIFEE
MSg0F536IIX4CCMRNBKmb8YS4uYInSXotT5jl/KnsmRLYO5McqR20qiImhg+AaZQ
AWBGUFU3dNS5LtGtQGYMAev2egUcDSxSmUeHjOfk/otBr5V/+zf3isXrkvmLmurp
3dlkWV9+rqnpJg1WYNM704vQFOc0PiSrx640fGx/kH/sGQ3BQxDuFB/7F/kqzxu9
U9tDG2H4/gsZm4er1IvJ5Z15o5T60rkgqgwZ/cGdZAOxRkuvqtPbVvn47SANXH7M
DlyyGhR58THU+LzsHOpkJyBfnXFnv1FPMNxWrN1hYoPkhDzbcuXp3tPdxo+5PqFC
dqEt7k3QHTUDvbaFb00+nnLlkpu/3BQEBCagZSoLWh+TXJ8Vs2h9Bqy+D50fUyGZ
E3YPbePD67sxjMbcNfDylbjKTId/zqupCb0AGMc/F6rrnw5xHtR+Ii+pivNleKff
7o+xuU5NWdyYRGFOcBhFIsXNZEnoX+BkOZPhjDNfhDDDC+HuIeAcMnDvRvzVAW5+
teXeZLFRt+xUoVKMYUTDvz3hkMt8KEOMTtYh19Py1dFcqZBMo/CP1yImwq0v9BMw
g9DzdOslOtSDLnLInvVyjlkKwACxNcbnOyVmZQM5z8rdOnnTkg+EI7TUstUmwuln
cBOgMG+sBD5+WOUS7hOxP0+ydPTMafsA7f4k84L2li7NTx8IEc+SzCz1/JtHd5LA
fLhHj7uRDBBIAwJ+itbx6+f1beQpLcxY0ZaC+U8JIhTlXQER1FdvKoTufPUy/3cO
jeVo94dwpOFQHMqCSQg5Wr9961zy+qz0HAoYd1IPO73HnLi9MgFAdY1c7F5/WTkm
xPylg1sBhyWeNrQENGVMsDW61eqwhqPn08tevYLJ2ir6pIPVZYhIplxu69Wut/fB
SCOq0L377ItIF+gdCV7p+kfL7GUEm0b687jixvDFs9xxe3lAz0L/S7pNKPuPwQqb
wa9qMZSklNQx55AC05kwD1BrPHPRsRjq9DfCBVFgrQKz6hEKUERJVbJ8aGFDiy39
rDW0CXV167jYTgQyZjH0flFkM44y5NPeH8cXTuUoqCZbEQF1EZWJ7oMTI3wdLJao
HGLk6VsHIL8hlW+y6/u3MK0TqPCWQRW+MCk8AP3QrOqYxIrRWLOCIyDTqv0Y8JFD
GK+wo0WGD6orF3P84Yg30ST6vI43BUdjV2u8p5uxXbrxsscnKEVrVcX+M5N5chq9
nZt59/fyV0oPH6Hsz0gimqFVxo6tk7cuC1AW6auYKvpU7t92cr+nmkwjO5U4QU/f
OrHAsKz+4PtDrir1j/aMsud8zydmeAYIl5W+2BDnF+/vmy2XMYojstAm4HWSPeLw
bX7h34VRva2syXUANfitI4zoeMteD+SOxvmB/it9YX81EkTMGCE2Mw/1wswycqIF
6sL9MVjxnUeY1jIHgy/206eVEIMfGj9rRo85Ja68G5z7kDtza8QMan1RMlc2ZJSD
scMAK+Qju5NLmeojfWqL+3peUlu9VSGVRSlSLpkHchm0eZmFDFvRzPCcjDSAiKVv
JH6tMq7yyx+on10xGTRFk1P8qgC6fN8FAUT3ap2j5O2zmEE9D5/qI5RJN3+vmIYG
lSjU1aFF77suGnBuw7w8ljpHVN+w5jhsT7Nlqk88IJgQdnzV3DLOxXMTCNeGQZWa
/fYaFwrUzKPJ7A3IJ48R1xDV+lkfkYBApGuJDToMEX3P5UTqR1dOeitKFYatz2MH
e8jM2qhFIuDY9wxQMtKDYx7Zo4Xj0BB9aplR6lePFXXYoU9pulKWMe6yiNNwwmG0
yb1Q/jfxpw8xOumZDgaEDW84T18liRwbpyOxZH9namiKNWLzCHfKnilI9VJ7os2S
kww20PbUleB1vAtN6BB1DgeIPbjhdNzMAuf+qZ6bz5KoLWw9+k4U8FOlvd3oOdqI
EQFsxcVl5H41NKwsxPbCypPx2a4KeJfPmPaqX4veqOR1NPc05VYa65SBM+nD0i7r
x8Kx1xJsj84cKvUT1qrOQgJJiyfHGarpGhTtIjdqikOh6121nQWUgNPRPEjbwixn
z02rsmYK8g7klC2fnMGdhtnuEt2pxR1c6s1/Wdy/2JFWfbhT6tgQ5+Tapqk08M9P
GR8MidChMQ8iOeS6gKUphR/Q7JTFrSuppnUmyH401Loq2GqiLR3DMPDm40vhZtHh
mh9dPuLs9iL5HVJVrXS7wyHmizz4ROOziJsDrxaWrYQMh1oumava8Mphl1r5WPtu
+vJ8OmdMIoa23rilqEOanUEjmkTC3aNA2x2VKOq06RCw6Q7EFO4l+gyvDiawYzDK
lFAbOVBMqLE1wCSAajTVWOoA1mLsGb74YA3T9XE1zpOOFZLT6lv7QZBFULHAk0jX
knuO1BeU8RY2fYi79IYkxTADMO+Eyw+p8PuvR5F6K85Wfsa8dl3NxUoa9FYrzwRt
TovjGdih0JTz8yUKeesphPekfd0PghAvFX8eMAohLq7+d1DCSg4pCDu+0V+vi60k
1u0FjKEHg+VL0gNAwN6qaK3W4CKSyABe9fPv3PK6Bjz3DFpcS/KtsfIqLpgvscBL
H57zBXGZDhHS/nqjMJs1Wu34qcKmc0r/zTkGOf1lRT309fOOw9zRvEJNQ5gvQ4Vk
eZzAVxqWw0rVDwG1nvu+FaBh5hYJisG++iMAV8Vw/ny6sLVNab0NLskqCYRscQPk
gMZbuH7jE/AJs37aA5GBC+9MuA09NmqWR2gT0EXh0S88ERB4s03iOdcUTe4BCzq6
i7b7dv+CY2b2NiZI8NvALMC0YNIKzC5kfojiMbEkC2CNK+AIUSbPCu+ScXoW2gq8
LkPUJ9K5IO7YTqkN9RE3aGPcx0IMgWWpfWpvztoiF2m/AV3IzfwjXmxl4W+urwwG
tZ/fO0tj+Havis1VJHGqr4ddkEI0qex3dZYEh56ch+ASNfe34LBQH4TqQAzxenFv
uaqvoHdFBa4Zd8ByVntb/ZV8ap7fB9VmKZkgbwjyfF7Iu1ZmUkkXxUZZ7y++tGcE
3yjC3Egfu9/QSnhEvlR+UnLS430P/cZhv8jPZBvh07bDrUZ/KPgNwgI1GFZrgaW7
SFhYKHSA5IAizwnUEZ6IwVKdJLHkoFanGKRBWsKRak70l6IQzOSvJ1lGFR17f5po
lCb1WrvWmONKWDyhKZlUF7RoBs/Kt/jNZKEKB6dz/0kFwNAR/uKb4pMpbVO74YOe
OnaYdPSCF/TyRd9VsBKubCRC91ifocPfXdTyydWf/BqkX7iQGsW34UVfP3Yi9fcP
Zp88jQXcKayQigbcnY+JFO6X5Z6YTw3rEFXk1OKVKfL86llfXOLK0MeOgV9aL2Du
nNrgrZfla36JfTIy23LVgjEsayqspRti4EXl3j/TZ4U49dn1QzJTqcbgX6oMeGXb
yyZpKzk520xaBIeY4GRBGnivoIZG1KvX2VSIZwkc4BnGJHJ9FBEkWy+m1n9X7qaU
sVZk/GsMmLDrgo2tI0UDoEh3gJnIC3sLCiazPj6p5acPwlDYVAbRUL4BHA0UOWBq
+iFJfryCAeYmkqbQf+MpM9EOc/jtarVb+f2pudEjK6e/UoSdcRpolQjlzQI727ju
x8NOctzafFkozgTwEdQ6DqxFXCbYQCZUNfXnqhdsemNb4Yq65/7BrnF4tUgrj0mQ
pNo0EKnPyk8jVdkSWNCiqA3HVjs5c8R44q+n/8+epoyK51R0HYRs0OQcRhWxwWeg
XoYqGsB2q7TXt1NRoUxB6XWGioUDPVi7bT8mXNZTafpRDuJ97kgNowuuqdYBsxm7
TMnlA36psMkcAaijYwMLet8Q5vfOrGaQW9kxH5wEYWcf1YFfb0qH0Hp0Lh/OgdLB
DQ68sgpiU3ZKBip8zXBMgoVfmG5kcDsNJT/vv2krAn5IY+ovHrlkAYE0JN7n1SfJ
AtfWpsvVJeVy1W9kA8jvSdC4BTpbaqksyIeXgKw5lNEXMehD5i3LpipLocPHFhn7
YbzpPGfD/WvknF3knevsiWBFcwCjJeoK1BJc2+zIUY9nfsZ9QvgVOtU0TFbveuQN
lS0GrzuKcAqUo4FDlzHELMq4lIqd/kDlEGazLaizrlg4muqpPo25h3+Etj0YD+L9
WtB01XRpUXvOQYLWwW5ilgFkm4S/nLTRCxB6nIdVAJVCaFsbEfP2aqP48rtdZw7m
juHMj5LkjVXlvPXp8W1XRYu7YbE/Pge1XIYq4kmKSlhJU8SdLL3OozGJv0xfncTU
6gGQehZGYcUxWWFSJReEi+HKkpsK57waVO8wD1UNU6GeepyG0C7jr9Ob88XPy055
KEtrmxNYKSQMw4LOaPIvsm7buEgJZMnvcZ+GyjxsRJ/bpgwqAhGm0fwtNZnnMtKN
sFRsRJlLFmncsCzMbKfIw47JTtUt1/sR4w7QIJkIxg7w4NmSIzcqpLrm1VIeubJf
5zs6s4pxapIXYOxH86ixZq4xB7t0MIoIixmLU4STLHPd54T19Rg1C7QP2c2BC9D4
CFuW694y5yoY/G+LOvPnDh+sYcF1EjyBi+FVz+ZqdbE7250SHq+xZVO9l40Y9Dtf
VDaNNnsMh2aB8EZVxEmczLBNDpEE0+v8tzbOtWh3Bg47SvyMU/Nb7NIhcHyW2ETk
ptIupy/w+8LkJ88utXJdY1WqkavWtucB4rdW/SkxeZBYcz2Vq4SeM7nMunr4UQZ5
pos8FN5d0/vT0SjDmM6iweGILMqS28reRsJuYTpESuxCfyBkQuIEyEc5h6ebR5Ts
3L3dR14Y8ZsDcN1/HrriPyYSLK/2dq4oycgE6EOMhck0Rq3V18iaMIudHPNlnng6
+O4j3zK5AoPodGCsblsLE+a8EAc0tO94Hr0q+Lk8vD81vzKa/K9F0VbimjseJUck
MTGVXpuqj0BG1Y945QGbyrWliZB8iu1q4yisjbpfEo07HC6/lgxn2cfS9EdtuCGu
IV2W7bEWN0cFlUC5i5CSaMw2jE7/VK8fT42j/YOb5HPIUjqSENnrp4VLnZtGwoCV
/qdbYKhzGQYM8YHzjeg5yQ==
`protect END_PROTECTED
