`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdQgMNgfcgQ/2T4TMAtqnoGys62QITLIbpBlm7nH6+cGvENAkS1OPjNT60adB9Jq
QzFVU7hAXZ4i5QYZ0N3nzYOZJdwD7f3rR5KX0SWybkEBVKKdgJa1lO3kvW2xcs1F
O6WwI+4TockSxk61s95Ar/kB4PXp4PJ4JwbqcJINb89IQmtFmsN0JKr58VwuQkB1
dFI/ZSMmUXTVgxRUEM9g3S9XKQFB5L+xT7ZfPSHv+ZnHtNy9CjM7UJD7WX1W/FL8
2HbuLX2GeSkroXX3mzfDk9jNtAdEt6ptnSNm0+vSmhJtjUTjgNBssxaS5e1NcLZa
dI2X3JneESOGI8Bj3ujflzZ05gLyAHPbdsiYUKl4AD7rC+5Ykn9209NegnWVKaCc
dtL6UQXuHfLdG5P5jQ/U/gCmiF26q3Tm3YIF6E5ivPS0jYF5rwGNciB9vEOHblJC
V7tYXtbZMHgHuArQfVQqM3DhGTip+mIDwBkp/Umpq3/fDI0hLqwJpyzsBV4FaHWE
BzE+R0dTjSb+Gcnf8KKanfBETdr0H9psG+EJlQINCBazSalZAS91jUrhn3J69f5l
mYz+Z/mwIwjM6wVJ4A62KJ6rPqYIWRbqwWuGf2C3zfwYLO3ET9OWTwpks56dbH1I
8HGxNpm9/sWqLayqTQQLWZmKpH+VzSNnaLK/2XBsxCg=
`protect END_PROTECTED
