`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OdL8kYLXk19DWyunzPZJVHFf9njzlTw+hyu9lET5CGDoBfe1IFDQKHhop9WV3bK
GiR54QY7c8wAfYeVXwLLKl8Jeo6hgGOydKlj+w5O7Ne4+77p6eZ0BJ9vnfCAO/Xj
/DD9r1GX6J4D+H2wEGfEN8+9z3LV9rRrUCLpFejV5bnqLhb1Kc8hxnIyuTErbrNV
kbvodGfFJikbp9ee6+UebO8uZKjAOSuXRvQj6BAcekAY1fGl1UIkUTINO7/NoQsq
DulG6kB/Y8RlZIHMrRh9HmkTdN2Ud9PB0JJjecH4lTXOGlQaIZFnnFJn8DRoCuYr
dqGTNbM3AM7kr3SM40B/d8CkG6h2YzIhum26Mh2DAGCYfufZ5RTSVL5Gv+gaivcf
OtRBcm65E8YSA38ZkqqZMZRQ7I2OiHWqR77m57q7r7Lu2oqiQNYoQ1llBVrJCoR+
hQb7ys345KPnVUs/FBPAqK1a05d4Dsneynj8AJ79r5Xro4dCzrc3Ng5oKlKmytbE
1HA+wkeQG1ka/0RKECv2GHL+NRrO4/x3trVx6y3+H9bIMsv8GIO/kE9MUzjhCTiu
CCM8E6uVhQAowXUjCrzd12/hgl4bBTjxEdmVy6H69P5QH3+qnB7YMBnGmcS2BOjV
5zis5isoFelXmV1L5/PhChhaO+a4Zvg4ahibiTgTRlml/tD4y+6n8w/ms5uWMgYi
cyMrtkZJAY7pfGGEVEKvnVCIze1QrzDrTEqEFM0N1T4//hJVCbB/nTKqDVF+CTrB
xGxvXnVGen3bPWalCYaSdQKU9M3c1wv8SdQnbB6yLzRHwbD8a70FEoPEmlclzLTT
YDf9R0iayE37AKE0tkK0xEzf1fazCDboeWtx3Yf+gfV4LEPb9MpLN3aVKTY4K9pH
eDjXrf8R8N73HOFJyWFBq6Gwc/qAw3vTAbInEOzTu1VBRMhbiyn7bdMb5JmDFbJa
TjULATO2gxN2s3ErGl6A00X2Px5x+u3jHvuLy+kX6AuEcytKwrbon69yGVw5Y4mm
FqSFQdSszf6HnpfH7nGTD24B/12Ddq6g5h7bVhBwwzwMLId0uBKqnCoYyzCrjk4P
35Pjg5KE9tWV6XQme3OtAgoYL7/H7pPTlPxSAjeUFW57vVX1GKZsvLg1HR1WT/RR
Jdll/9/G5WNrHy2KLuKfEfig+kJLm5TDLD1DRCEJ2DnINJXPPPRnpLfevS+7Kt3S
Q2hDE0I/+dttInwgeC2/zEj0DwD1ef3p/V2lHNoyyrh7CQ7BOX+UOrjQviNvndXz
idTbhIBeomJeui/5txIoWPa+FQDt72YZkDlwLm8U7QKTZDFqWEYsiTKg9WY2EKkI
nseh7nUWFkP3GDoNHHHjI6vqWvpw0WlujQbJ79b4iYfAgUe8IGK6bfNkI3Hkhg4W
cpgBiFn4bDMyF+YJdW1bSfZIs+equKlqrEIfg8EgQU/dSriows8Z+fWrMeKe1cee
JHIeM+Ct6Hv7OA6Aa37uQcGWi44a1E3eg3rqhrV+9OiFzb3cC3wTHBpiSOtjTjhv
MnDqrxm2VQLk73RiGvRM/FVUaNOn/gTH7UBPZcAXCSEylfjpJSUkreqdki1JR9f1
wgnAtZ1sujakQXGa6l8OVezQ6zXtbSqfkJ7i7qwfpp3wkHUnCex7zzj0sM/32t1z
`protect END_PROTECTED
