`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bG7oDIaZgHdOnFwFd4ZsI7pRamynGIH8SHk3ZKcKe8GMqt9ha6US5ZI5yuJrWGZ1
TijPJyxjFmJ1i+oStcqq79x/CazsoNIgtOXa/D2ZGLCiu2DXyUbvF9cz4rHcnj7O
wIU+lIkNNRrb6b7s8SQ1Bg1+IejH0D5wBfKsFW5SFEO9OM85r4yzwaOZ0bfOsTdL
QJGR0pbc9EETZ2CHGzqRkUjeNm1Fl23ipPZGiBZcD5+TjDSTumKGyJxIPHQMahYt
rno+09K8aPMA+ToZ9MH0/eUIZ4RB5xSlU1ZPu4ESFOwYKf/nQV7p0bWFCmNC3QXx
EFVBXU6Nms5M92zP/tJ8u8SnCHBz/4wHCaGEomZLF1CYDXmUj5/lLHyrh5UEufQz
pXwlPDbVbaixBFZf4q/y24x37ItBM9QOSS2I/52Z3IVqZGKBm8xtgHFv05za168U
hRWPi4tMX1pA+uxMsFc2hoSU/KiQyYEt3JDjGYiW4taKfMblNK4YkORizTvwQrKQ
NvUXaR3QzPVLJApwW7fV4vSFF60wV4yh3yQzcYsbSPPdlTrzsS+pzUfIxBEwUpQB
Nx1ogeiNK1qUfsm/HMNDeA==
`protect END_PROTECTED
