`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4q68Rb1u82ltqqSAjwiEp0l1cdQ24dQNjewb4/iCnxkZjtk7go1F2DuKCb14xguG
qrBYm1bx51mRKRevRShFasMy8kfQdTn/Z7kFZ//jexfI7vQTwJJjk4tqVgpzs0Fq
9NeyShOtCE5VNmed5cJXdYpinx2bm845PLv3q5eSwPevjrdZYETAskEjsEz3vczb
5cWA4nMJ7wNsjNuUn/pzbFOtk2p3lk0qnrC/Xvuzjmpbx8c5V+4OO+TARGv5hGM4
s3ibQLzrOJ0sDldwwjf/Ettc1G/2ngikYTs8+oAqNPSeUskzbIOgC1tWi/2SSeoH
BfmH26rxk3N3hm7PsqXX+Yyo8fls5hl01PDy3hvKfcXYwMzwcKGtdE8IkPor1IID
N0r2qKtglci8uF13OOreqp6Icxr0sSDChdIS6376jpGi9hjIBg+ANmkWx/9yi+8v
pLSVCfFp0ltH1oDikviSNg+fTpFfukL2SBY0P2jNdiEUA/5kMy+prUCDMpN10NUo
1eZyW6C6fnVuIJad+13+8hR5NFOMZYoS4mPyO+v7Kc3W3jq3Z92lJTgo6Ow5JVSJ
P3a9toCHFuEkcN/yIuTOu+Of5z5hsseJ6XFjmN8QJu2Fab30IuODBpl+Zb111BYK
95IncXVc2eUcJlaB4aIzmGr3aPrbjLIE51QPKwpdipVfDS8bV3rdynEY6dyyTPxU
p3yD9A61jb4ceWIfcBdqwtPNRGzQmzhbtMLPKNrNAOJ8BjjvnBPLqslUsVZHndTV
I4ZZcc2X/W39ZlUZI0bnoeSylKKhOIBhSZmNXHxG+EHg06E6fEZqFSQ7Y5zQGMsI
1F3gralSPcMKKdVdzOGeoKttHs6E9RD/SzDrDlJzmniGqEMaAsqaqUS7gtaxp9l+
r5NwoLeHKmA2QYmhH7joT3f810TpJ5V/rqqm87Bsyc+IKJ7IWtHkIN1f4/piQ+3f
4LUPZqL9s3HjrMg9MtNo7XDWuFfMmcSHJQ9LEEvoM4UE0GLqtCr4gOxbrbr5Kefw
fmh5kofoQT0R3qds0klZTx79ZpIl7NUULvm3fv04u5MnbyZNVjk7rw4uYcSNhvEK
LgqJjc4Lz+r23HMgt+qb1AK38klJ8W6Gfn8yufcTVKx+q/jNnFeTKtP6+DqJPvfo
jqiN9+RDdti9syW44L9tNqfLOnewGmtu4ACtN9iUCuDncjqSEyDqShK4Zj1kEyF+
Vy6sf0FZKQUMXAane9TbYF9onodJNfKhPByyxcntaUfJsdgfyvJ68whT5GzAP9Sp
nkAo37JalvAh1Kp7e4gPoU6Jr3vZl+XHCDD2Oalgk4pB1F9bo8L55iQIuO5wvxaS
IiqB8mr64Bs7FsStLtvgGz0OdM8BfnMi9kNEuuQfft5VAEQlSi8oBcP3coucDYnt
RzNYby1UFoGTzlSt0MDAzg==
`protect END_PROTECTED
