`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5uvNH4TtAAqlqtiRX1aVHdbiJmRTDpJcJgPt16FREl8QSBtHkdjMyqQGXpqg4e+R
iioXlpOxhDRXTxyBRzGBOvO1/Eb68GKENAJwP64r26yJ6B6PnMbsb5BfSk7fn7uz
gSsP2b57Ap5bcG9DKqGNKWy+9yH9cAG+JMUZ9dkw15GsQE+gzBOMefVTqTDHs9lx
2CvRDaWcRNe7Vs45ZPjWd3ltZFJeKsGEWYY1I83Q3keukD/bQAuMd5aZEI+5xsjR
PSdxvUYgUtmTWCEqIVPCEnpS6DkMPbSHseEL0Y6Brn7x8HHKqth+S8V78LLfcW0F
67ENH6CxFl3T0hFG9fGlsroVIKG380aUeSdAE4e2Jj9eZyNQfVgGdRPURroxwB/b
g+OGIBXC85gskrEmaZ+u6fOTrATLGof7Bke6nyTwBTytTAKT+REtH5wjr5vO7ceX
jHm858/d6IsgAYvjDEdRcrL83KRQ4jC7e7zrkRVeWHnJGwXQk0XJs1IOCNxRxIzK
4TO6IpPSuq89cZZImAuGEYHbp3Dn8QxG7JU8dSujhfwSxAeBpyWySDaeqoH/SOrh
AwYVM/Yxio8/MEqQ2nf5npyyboH6oLbdRS0kBSym36dql+uoXnfIZozpJrpbcZwH
x2w+Fxr5zxayl04OrEZqsSfkvuQtocQLAzeIsrJGAyjmjlQ5uscMEYZjsJJy8fzg
eyvSmvDJWcIxIiwVdznzNPtlsySEgfYgyJTV1JWXV5QoPyfrJga8xerZSpnvH7oS
w0h0IKtYxrQKLzP63uDtA/3CbUzD9ZSjpqKisUCTfzncEYQ6u3bvIMfi6fNVVb0u
dbFpMXywWyLcxPzX/LX9UuKTRm1vw6xEqCaJi0dE7LB1ElHMx10HbwAnWlruiijV
aEsGzZmmkVyBCRvGGymeYwsmCBGv3F76DJtT/JZviFD+lPABHAzhYeLiQEPynUIl
FvYqijEddNEZkpPbH0xbjY9wpCZS7HdjgMH5P7Gxg7Zd5ss62+efOFCTFimHONZf
rnxsH8vP6CXqIe9vxKDTbuu+nWAn4G03+8sbcWcFHnqkjMqjq6FykKHrRHSwdBVs
NEiqd8wd3nstc85BFnoL1vmYKnk1mQv1G4h9J8HXlqbrTnV8ZEab5GNb5ZkOIRSF
YXVtzk3RtDe9TPRNPJoNsTGgp3jfZ4TtVUtiFy6xO5Qh+VAkK3mOLQ0jYiEYe8+V
nwxDMov13XQOWIvvC2ghrScsqREgxg0qf9/hFwGsoIn2jL+jT6pSb/dp/rEC8Kgc
cZBJs33/qVtP894gVvCw/UW5a5F5yI4k4G56UcsCPCf7N1RNdZCzIvwOT4QehU3e
ahSS5sPylLNpsgZ/7qvWxiqXNqpfuXFc608fN4GW9A8x+sTTo3TVzKWXuSGrpZeB
ECGcdK6TBdnkNk4H9YCeMmjy1Hx9g4uZY2K/e/EBAuDyaN07u48Qc2fC9i6wY9Ue
vpxhmi1MG8Q+/SOZoqppz0fmPVPwjqJV8ZYUIeIfhj9i0+Ohd/9604aIzzEUQJgR
SnHoSf9XJ+ZP2cV5EKuUrlcvf+tyIIYAmEJa7PmDuR+Twd1Vfik+rwUCyv/XDGOk
eAz1Q5iOz7tDIqtH6VI+paHnodziiOkD3l2n4UO2U8pEx+ZaPpHuxwoxBK/V/wzO
pkDRGcPLgkw+szHqAZ6flQLmvXvjRQ+p/JH7tDKyaDmoVtYt/ujl6gCn502xWZiR
CLa38osGXY72kwfLCo8LKSqpL4arp0PU9pL81LJuxZg1AXDBsh47CIjK8ZYeHZJ3
`protect END_PROTECTED
