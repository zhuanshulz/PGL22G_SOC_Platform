`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SZ213EWp84T4yu2hnKeuBzfhmGhYLCU4rrSw8CCbsfiTM3+bNJLIztI7jNu12gUt
q8S8mTcNnlEZC8xPCgvEJq9nz9cHDdcyC53/0ogFPtXTsf/sphDJjMg8JrXNzIIi
WJPVJIZ+CTLW/vkzEmWEz3fZcqjPe45sjwAsCrH8ItyZZWiGwcMM+US4jxxPDPlv
J9mwHRfXABzw6XBb5b9vuQ/mahjOH4cOIotyjZMw9l5d35L7vqzA1f/EVqVZFuH9
DP2VffwDWKHe5qyjxGIrXivnkv+24DgoD7UaAsDY3BuMRpFlVCX9SjoPvxrgwU+Q
K+SP37Kp5ZlkfJCg0yKrA+6Fymfm9OmKAw6wZuMf3mo=
`protect END_PROTECTED
