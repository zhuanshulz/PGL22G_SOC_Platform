`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAxCk+6EOwPtcn52S2Bi1/dRFEj91cCDRmFkdPyzy/v0Vp48Nq6r3TEnYlYIRqbO
VnvJtudeVjoYm4wAAZ9GvNGYRpPhllx+PfZol0Z+mbYZZyj2Thhw2TSHMrrapnkU
uklY6ykTqlZna4oy62SqMKART5kqPQIWG+SjYCg26h4P0kxBh47WvF/E/7GZdOTF
xjfapTT9ApswdOnnuCTMaoVLQGRKit2dqgqHVAhqKgzX+9JJJtiFzCnj2OIA1HmM
TQ7YWJD1bAyezKTEVGGLExztNzv3+AMbuZVrJpwLjXzVB9TdAOvKKyO/bIU7ZDaQ
vrkQnaC7gwwhA1ZWzWnyDJAEYyUEO94npEb9KyDK2Bg8LzjgN1YMcaDN4xxKxXyU
FV/yGrqO4hKGjEwiKfqmqNzX+OUzww9wQLjxvQ3acgo+ZRLsXTfNhjWhAiYorZbn
4mTPpL+MmEg9qIYDfb9u/1kp8VYKeADS3dU1V3raR4ZFc+G4OUMLpg3tSF/Kcmid
HfN9x9t30dNEikt7EC+NPO5Bob5vGkgopNjAKzL/gT2Kjj2huURo/ImeCqt6GCHs
tGqRL32w385AW3oMiaW3yM+3ACEiF1E6oU0fcuSwAGxnvhSflYioBSieV14pm/qq
7kXbFfk9o217W0rD0L1OAeGn+ioSeAtRazvduZzq9Z1Dd+dx0PL2Y9SkutPlCyvo
YdK/Q6ydbsp2qSRC5nwHBZgXanb9Uq5rOd00OnAKu3KfBqCY7TQ/D0MogC71FHXy
oa1gvCuT65elBXwI0YbOx3Rk8fU3yXhJbBTh8WyKz+0PLJ0/kpPYXzIO/DCc/3/j
3FV54ZL1swZD/Tzs7X0mtlgNS8R9h2eSuz26jUOSzvMJ3ST5pT6NQpTSf0rvvbLc
YCEELOzXiHrAFNo7oNiF2ljjl6DSi088lpLX/jBXSEtmdxXr5dmhYbdUM/sPz835
j34eGmMu/XWzMF1hPrIw6NmzMKoYvDlO5lfunPQ1r6RDV7bkUTVUSc9fpA8yMPEG
UF5U9UfKEwI0EEFzsFIvoWI03uDG040gq6TCjhvgXOb1Tb8hCUOa/+8L1dnMQhMr
kYIN1Q8jM3U3CGfe9CIB73HQ2StXDfCyeB/cZbCjTuVYWENRrDgxGKPUDnCcM5vx
fp8vyOEOeukZrV74JYHbGuGFPPEe6XAbazwMt2LF0wmJwdYstfoPMCUYK1eXyfaF
KniatTa85v6QRZW3B4Z88zLQqBt3XkqoK14/4A7+AngDqT7wWkiPNu04LV0idaJl
9qK8K5MLrUDr5oWeB2wjO2kk8mK2LmevkTZ5V7D4GBE=
`protect END_PROTECTED
