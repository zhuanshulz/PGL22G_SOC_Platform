`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aToG/31i4u3BKH5vzvA9h5qUlCp8788GTDSWXmhz3GDTxqPKoaNN+8mjSBBs2Yn8
EHyJ3xsZm20FmQSuxsC14NQsih7ovY8+1bTBZIMGZyHS9VL9BdMoY9nqxbS6nzwU
LAqY8eCizuhBtl6Xj83lQde4g3w4vjmLJr+UepIgJOAB4s7rmpk1nEO5htMPtSlh
YDTca7JgwEoaEvjqCrRdapgxjLyf6ThcjBsXwjYSpfpmFHz435t/8HmLv//z6TFN
Lw2WRGxZo3bGg+oQWsX0ZOJofZEQxKaLyRtvSvRM/3IvnpuyXmm3t5Z5w5rzfED+
YU72qBir4NnjywzDQoUDAjYLJm+qSc/DlAdCJfFplBkEcnvlZr9mZROxIH8IzTv/
zv0MZUURjVLm3mbp+/+GkSFlLqwDo4x4qfXg+6F9PnvoM3Ers2FKHih3YVCQA6JC
ZTno2xXUdY8D81ouEHly8e8f+I0/N9CEwVGjEwQnuXVMtToRE32vudrAQqLk3xzg
Y9vfF8TeDmPXKWLMn/vkwEsVo+MCt/CINSla+9ApHOc=
`protect END_PROTECTED
