`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOp3qvJWtNoG2TiyxCm9+NgFYJtmCZikIYLe/BnQRYyz5eX/qzTHhj3kZ7DOBjsS
WjGqqFpXW6jOL3pesJDfAhexwxZkkznQEdma5aGFAcR76fe6/YC9G3523Cza6omT
OKYwxjF4YOXEKVM5DKsnWP2+AeBGnCINDtkqOtw3/fB2PI8O0rt8sMm60asR0+ca
JZEh46DWBT3tsW/YkjDdqT3G8reBmBKKgmoKdSPYVBFwJqVn2tXMA62ta+25O8je
siXBPitr0idTYgUu8aYw3lNeN/ud584Yja70eLdFOLCFOZtk8AYrsyvk11xpMFQH
KtQkMNJw1rQvRiS/GpafRqGgVS6bTLi2MQ6LVYhqTmftt5WxqKU3vtdd3rLEL6Qg
r+FcwrHxJ2Qd+qfq/IJN+1ZVnixvhes3Zd/yBybnkS5FnxXkQfgxxoFTbcAmxYxP
lgKRvRT47aVS8hKwaNmiK9XiR043O74s7PCKsz7XXNwpM1oEwST/4Mftb32kZkV1
RnaOF6LbKOKZOEhq5QBfb4FtoR2RJas2TQI1XuR77P2RsX+vIuwinMdYvDDtih7Z
Nbb50Njfk28llX8mmiAvrbVngbuEBVJlXHKQ8EFAKBd+keCAFYdJiRuj9rZcKcB2
pVSd/EtFiyHXlATvPPlDyALyg/ZPZPblzvn7t5Shcir60/JMpXZa5PovwFGOMm8d
RM6Dv+VANoVFCRSrDnvZVilKKfMSYIAieUX0qzei9llLS8wARW90b9SX9m/EafWT
GxrMlMt7/chQXxkDZdr/qXUkbHd5RuE8I7HVgh4+3C/jEgSaTMx5TuGWPlgCMJRi
MtX2typVLYQta3vV7STLaYngufPIuwynnYaRe+Z34QkZpJdYNpjyVwvuy99jHCFM
d5VlzWnxZ8N/RSKoZOLZ7CRj7G66+0tAa0XOI7royUp1j9zG5GJpgX3PJEfoqOLY
UnDS6MsphZ/lLj1cT9UwnJoq50QRfREgp0KITWLYskqdbURziTj4tQdzYkc79LxH
ehEK1QIB0ORsa9awAUi7m0+jPXawfzAAWnt4lbfeGsmljUIggGeZEsYwf4qeTCLq
pdL7a0C6kqvXtSdLxEeAvT74Lpmpagj7UYAAXB07Q4TElWZMcRl9t2LFEDhG5Dns
juaYx55W44d9BQZK9WiMXVSZ8RSEwEeEl89EsPRVTCVc5RXUnL85Vz0JFgIxAXeS
+CtDTAvJBPel2pBGdNLDjN3Vql3QSuPVMsdVYSyNvTB7f2a61cQEdTwiRn97CBHy
QlW0PBtWnMj/Y+5Qy6g88xqSbuwMQVS0bzoEAXYbkmip5l5nP6TFd+duoHxMTy7x
zZcw0PcNjoVafhe6qZPs9d74RarKc/VmvM2kupkHBI9/b833OogNmYkBQUcpiJj9
XVRD0wy2i0ZM4gswgO33Wq6SyhrybO/xe0HBvaQQPNzsyJ0nTzUraHdSIt7NwcW8
pIpQccVD9ShAOoGA8YbzhA8NGni8od2jtNdCFPvMaVWA0cuLrB6DI5vB4jKO4r6/
TIog8RBiVfSom2dt1epXTpV/nPeg5lB4MJ5GUzTh4haLZGLTI47jh4PM0L+Ljs/3
xiK6BCID5nNnsMP6lSwloaXAaozVNrbUlEOK85XqCTAyoLKz1jcFe3EgkbNk3yTJ
RX9QzDdiSq5z814O3iRikQUxSfoflwPV49dYzwAuUiVF/TBNCd9xkfMSeWnTTe6r
1kM5LaBwEJH2bQqZxkm3IR7GsA+SmM8JscEB+7E/7aYhbHxVAFcOENbe8AAgKBJx
EghT+kRPs2vNu28rHq2UX/hbM7Br4pIP0TPIXO5URr0hu3qOFILH0U4uX9+5bgXP
eNz9suvGaaTICW9RydnAEUdGi+uTlwZbqiJ7cKDXL8xdTvmnblg0jFzo1xWmXRy3
juYDKmLXeYK7VRaFNxBFP1njI+zFD9R/dDoPO0MZqOdCLM3FmtMZ4b7PJEbvBmP+
WUsIuMi0YAcRjlGKRAnrdiK/jTTufxpF31tqX+Rw2ruIxlbtD457dmY0UgrlNwMG
oBT78JVr97OMAcIlTYawpOMzVc2TspaXF0xJerfHWFJo7+4ZyzmBG0EUi1G2IhW3
RwZSCWZtzp8fNLz+dwllN4pRg4nzeUKSxGiMi0Lbuy6zRVT/pExxlH737kWSpaUA
4doc6zpW5vTuMoE1ZchkkipHDI7NnL0mVrrHoEiJse6Zyt/ZtlJqbq3ZY1A9OLL9
UQ3Y8g92vqXp7Gl6pGt3XrkrcwNVOLOTD9o7SaIFncwIliNAGlHqt3akApexkKan
lwUQo8N9vGpqr2MBK33Y+fkgYrwpbweRJXu8eMR6FqirjUK57Nl7CKsiZ3DbRKXh
5jdKUF6jjKJJ2LkjFc+WdUuPOTJ2mrIhyH+lw3IWE0817NMHPhxJhEySpLY6WyMG
y7J8MseOwUaT4uxzUf3g+YVwHSpG9IQvklx7evKB7UB0t5nyA3q91JxhjyvF3OY9
YqxLn7xHGQqfrf/zT3ZAJOfe6hRt/HoUYJxzZrqi/tmBFcCOKTndX5tPHjDx4haW
70sXtZNF4Zisy7ZRBZqxqPE2ArOx2A1aQysQwClDwridz1xivphKMyDxfuQS7Wro
HUh3QRSScDfbSXoIq65q+STyARah+VUVtdwXHDflwIH4f8MklUYBuMrV7OhHqiYl
XW0My/ZSy8HcubYhDkeM2OuZwyTsuc58fY8DySKt6bRC4oxj9qP5v3se1fnGAyrr
WD6S+HdLESkIVgguZrmZsk4HMqfY8GBTFL4FJZnQt4xbTjGp0II/bkmK6bX7MUs6
2i7yOiqnCoxtBZ8UvVHFwKIg4sjl6MESUp3LTA84N4nIcVuZ0ZMlgljVx+etR6TD
6WpZ3Zcuc/BR1XhowGIp/+IWyYaB9qkGKA7miQdcKrZELErkIxKYOy3Z/bX5lHap
Ga2918nsqKCHrZveMx9D5d+KB8zH+OIr6vIiAQV/BF53+nick2VBx/Gll9LJFsM0
BvV1yBwcHvSxmZghw4hQtq0J4nzGO2yEXWlBvab5AdngT81HfrB8Sbywbt00cItc
VzA5LpaDsdzdIAVP0I2skrS2Vo9qL/NnbvPOpWI7r1sRx00aW1A2I2UHNPFZdJqc
Db9qM9bvSKFU54DtmTbQEKyIlo4lWXLn3nTDH6ihhrAU7RgzqsM8SoFQ01/0TAu6
CwbqpYNmJi17/2jUMKk8SMUDOP7k3HjxhmAe5AEHMa/bNxhDpBHrPkMokis67xtg
yWlZs3Nti52WXomaK0ZEDt7Th6AAifkVM3MBxgL+b2F1WwyeA4Vz6JNvkVKXPRwY
gZes4fe41Uvqzkv8rSpMyqIvNLKoxngKohQaccXVkczQ9Jfg3g2fiP16ZSJgi+11
BhyS1qkBkql8zbEz/eWyL3DYmDKka1/AYR5z1KghrwGth3pAJ0vNNLb8xFzByX8k
uvwTiURnnXRyqRuAR7YuZhH9vCPd8VMzldC2sFrqS1NZ3SEsZAxvZGtPKWBRCPHQ
EpqFxzw4SPRiIRewKSc1lwNezKgdX7KaMtnCzNxX8XfExcqLHWxG83U09bFtosZl
7zxzDVIWdlAltPh/ub8xN80AhWbEebnXz5J2bcYDMm501Kfa3n20EeJ4MlgNlb4N
Q1eQkOcx2FjxDdkyMO6kjwWSDOkDGot2Wl9TSpAu4QWHNAijHXF/WBELEsSmweJ+
/H+WqEBEl/tsFTlbQcvX7TWUShAZT1JlaTfaOBH58AmYkybtnIdIY32gjqngp7R7
U2ZGt/OufmTr3F5YHFJHc9Zy8zJmNlDT603tF7ZH6Xpj5i3SsMQDbxDKidq2kVei
xT0QDhK7dWLINSALHo51xsULuuP9OW4Gbla4WsO3TqrmTP2RPmL5HUJ5qlcH98+S
ewdmbgV6ba1k+l2GoDIujFh33fIGYWAhae1i4yhPxKQoG1lZN5wkCCyyy5M3dXzA
LCAg1PBkpNgoX/uBvd8tXBf4CXbaMM7AQOL1WeZVwR2dIpLVfwkHBkJnxnv96JVP
ueT4yOBQqtjxuuZYEzr7qq6mWsPYNKE1/39fD7rXqkeWXFhnA9kLEB9tY2Ki0aa6
I1CsqY2WrrccxcT8ifpEnHdSTC7JjouBNEZMogUm1QUQs21TKCW1c/lLhVBMcd0O
gV8joFNfRU4cF9Z9EZ8oHeTFh5U/YBIs7hv8HFRSt3p060dlZhLr5TavKMtjFfgj
CSXW9hKyPCW+oBqZS97Q+BGl+EkEMBdfwlNuydcb52mqGOfmgj0ifIGUHtVVh3z8
HIbFaIlmSKjfl7e+59hrnWN0g7mtNYAfXMCqLpBafQsLGDjPHC5HuNXkf7KkhnSl
ljZWFFXI64p6rZKmYXmzve8/kAs+Rs3eD0O0cerk+cPD7raebHhdqIg0F8wtzDpP
SovJtw+/aIK+6bMq5cZw8Y35inhJwfrKDytYOmWAXWbm7Q1tx3G7RZ0JXr5fvERG
e/HNT5r7coPhKYYVKufK1ZHv6na/U30XX3OYpzKRlBw4ZmFGh9VoGz5Hw7oqkFX9
bi+/SvyCU83tT06LmKPYOJIC9GT8AtC+4PahzKXxeKqQm7L/TaoP8zWy2MryL9cy
cZNSkrklOuezoiS+YI9FJst1XuCI0umIIMKohEV6JKvglfKSPq2pwWDfR8rLPC6o
EqoXxkPvi8THMky8/lNjRoKayyGxg0drUmFaS5Fdd17gwc2C8F+9yHagPQJhDe1Z
d0Q+40rDHjS7CIhT0O+NiHjIM6dzeb6reVsYCDYC3yCnktyZQ99J6KHrePMJ7r8L
Ne93ChwqskAPJZNnvyCnWDkbg7rq0FIQLhqQSOyFkjlh1XMxHslYoDdNkPPy253C
7GWbQ2AKAehKydcS6y5ob7l7OvCSQbHe+V8zZ/wwhcJU0Swo9NMIsu34CsmMzB1I
6TpUpGXY7PGWkoO+NO32ygoERwu3mM0s2XlcIZ+4b4O5dWE6MriyaWileKqbhi4B
3fIsTC6E/8tQvf3wOJ93VP3J7L1KtJofy8iBziXO8eGQK1b5D8yxn4DcJ2rNgpY5
9EV2szbZlh/N0E7Ja4tsIpPIhmR7taTbONb7sQnUl+NBApjb1D5/VkjoVHPcVkH6
ZYh59zoiybuEE1/qDqlm8k06Ze7AFrPBfcogq74MssVDH3rgclyKqJxiRaynnpuJ
Ql8kIdsD+mVD6IpvyG/fl3NL5Crd3MzwptnlVUwzn1kVf9CN+9KYS4DQkHGTOb52
krh7LF1BFvdNUOYJ8zIG0VHVuyng/+ZAwoe0m1mF/bdOfrlSBH8uN6kqsSebgz6k
lKM2a/3dttg4ZufuqzGj3BKQkU8TsrZHcWYzm0qq+YKVjj4GmwQNfwe8qqBcw3M7
UnDXX26DSXTiijKKq6TRPOynK3QzXjzezJYk91w+EqT78UiaEsA1AMapgZnfF16i
ZRHHTl2NocIKgZGRow5gP9JKc0Qa/lO7zhPAS334wFX16myPqJ5fZABOuq5xnyAp
nAoTkciE8xV9ohfmHgJB1aNH1Zm/wD+ZBPIDu0cDvbCBGngHCUoZLXIAOpIsFoa5
7uA/T60IA8wCB87M9Es35fPSdQIudhjn1V8N9ofSGZJcyKrSfKgfyLvq1AGVLEI9
f387mQDHXcXlnIHqQAJwmr/lX0ExdWERk1d1FqLldAQNfDBWfbZTQxpufr+mNQo+
YxxVMVRZWxZ6cu5WYGMMBhJqnFJfsFQ858QnM+oVO4EF+duJQvaQAweeAEpAf9cP
WOjLqFSlHhXuLBzCGXRXaQQHG0H7Jh+GhE/hM30V67+GeU1brOIemnBWjtYXALtu
X4CHt48JlFQ5PeLDbuZzYyE/lt/WTQck8f26vBTUZCmDa79phuO/Lj5W4WuVEci9
7y7Nd+EPzEb7ab9qwbEE6Vwr65vQNzMfMpnKMzlD8YfkJktlEnZh01K3mxQBaSpa
u2amLxocwpGsql9cXxyS7AA6l2wM6gpJPb6hlj84g8rP/8Su5ZUmzg8sAQ4oQrZ1
wYG2G1z15uSIpZdUahzYdkDz8A07jGhz034gO+K3cd9qK1TG/IJX3Pm1wZQibQby
/+rlhn0kwFWBrd8zu5SPkdMbNf/UYmVaIfbyOugJthXF6NB0svIixIUFvVvC3+qw
ZpH57iwXv/v5AHe+ClXwsn5KM55OGNZuvLtoJKVUMffroufHeE6TrIYHb3Xp22lf
q6jzGWJr8rZ+uQ6kcmgsCRdPwLY8H1e5uPhoP7AAVSKRPw/DiPDr0YTtWs152hUf
Ty/LIi8qdIRTgR0O+9JGzykDXNhl3DDOLMtc5WEABNEpA2ZUVpCuwNCJmIyRF1yU
1jX7BvQEKn2oTdQF5fI99zd4WjU/be38+19hEK2Qe7y0E3Vh08ryOFx33Tic+o3d
R00zrCGBXBWw8pOPC5Xwc1Xyk2yK98ABer5XsLyN5jb5wc0TMXgMeNEnMk81ajuj
NVmfL2bngH1qSxxZzy+XGS3YXmc0zQce/SopuFAwMJ6ppF72Xtr8X6MqQpm/PuEo
LInp4ehE7hHVZcOLHO3EyspL1QDupc8LuZd36Xr/uHU2nFOTwOi/IiaxEeTEwYGm
4Q92LHKebtscfUN6WLGbJ7/eIp+rAUJ4jjGFCDkKEZqzVI4SKkqaiCCU8GUxfg89
nbuByCGmw5VCkoVwk0kKgLDrMetV4VlafNu7No+AfgIE0/qBCY+4aTnoUVWX0K9L
zxjjimgcsP8QpWQEtHY10z9KLX77yOdfu4KJFF2ir54rBZPCgESRWE5UhBXFMkDU
KKZO1yLnlammgh7gIGl8JdbD7t8D+EpTkEnRKehWAhNEhl8t2xbxxiSiTVl9vL+8
YxrbUX9cIbPcXCSAj94lx4wnIJqRKDWjCGYhPgxcd9RdpTQvqIXOUfcGkMgfYtZi
nED1q1QtCsaS2YY89unYlYjiM56K0q964oixaCn3gyluJqv0UQlz2ZgYS4YjaAzn
9EL5vQCauEcYwkje3cvsnNDjxeDk2CnRu1HdCZJcSBHkIMujc6+g9mhVfZXz8R6D
4KeDKpt1Ydg0tf6jxs4dHm8fXwFAiWY36g/+6OnfSe6HnCS/kevC4R5P+Vt0Mrvu
DOlnafY6QVBXNhzgeTdGiFaj0fk3Jk5J4qUl6RG7g7KBD5n/dm/J8cHKp/seAkkr
FgDbaWB42c1H23rxEk4a1eC0QyES5Cv0xHoSeRCvk9djdgd14gTIJArsJheYzXN8
YuK6i+hG0JgQjRWi2ZW2aj+n0Pdj5ymFi/y6fnKbVFikKEtXXNPNiW/xKLesfhTc
0ffcKTylWZJPHMPt1nKA731gdY4MO9VdxxQciQE434uHQASGtr/eewJcdj88pLwv
fHjy4Ixxs8YBBivVsyl+0XblhgVQgOLcGcquqpjNBXJVgWLcvO5l1aJtYkd77/+c
jr2FI0+Gh+xoD6l92zhI+5MTYOQgdJcZZLIATFT6wdTrfYzInBxd7vEk9eKjx/Fr
AdtWBTtA4p3f4WHBQkjvEU+kCoKfcXxXM9dgW7KUd1zn3GhWFV2+p71340U6SGcZ
Q2GMbq6skVXeylZ01sYHo+VTBoNSB7PDXGCftYz4xgo8w641Xjss0N5KTmBYGWjG
TgZrB00nUYGYegH0clzT0fcb1crOjSbd6OtJ5raTYxm74Oyv0iSnv2ihBtimiP9P
ThdkXN7q+piAGL5tbMMVWfUG2oyB0WuG748dipOnS03CxHYE1I45f2d1qNi02msy
lRe+rz8gL7O+kda/4r1bEcatQpvQ63iwGn4Nb/Neo1fssLFUhwisXe3g1Poh+d2y
3hksQBIdNDmTGzQpT03GJekBLL9DQDmc5sV0NGFpezzvjarfCUhM6WEhUDnCO0S4
nnK6bVWwbzczH2NZZ59KOrOOWxpj3NU4oz6adSK821To5mpmmYqYx5XBDvWWs75B
hip6pB017x9YDl270NFlZJj64xeSHzQUlyxxiHtydbzzesb0PN6i/OY93YTpfIhX
M5Q0USvCmvEkV3pydQaQF6LXQHebba5io4ExVprqze8/TVoDIkjzqLzaCTw6vvkd
9XbnmCRQykENAWQb5jFPT8dWPkwWtF1FTmof6wnTdGNtzhe6z1sA/u4ViSkGlJJZ
RPnysP496MFM15DK9RvFJUQaeGVbSEladJwIoxIAt7t/4oa4RZc1W1B/Mz/23FSr
ZCuUJ+VRWRt/FWWWkoHsAXSu61yVtry6wbLB0UKzQyX9ufj8cmRk9fk/n8N8jxpr
u6Sjoti9Mq0NhSdXAd8aiQU3b13BJ+81cMDfg//pL7tJjRPb1r8x7LeJ/RgNOcLH
gpewGSJpMpG7kl0TbHeodOZSLceUy2PXjinkIOZF2Ma1cteUQfU0eF5Q0oIDp+Su
HKD0fChFaLfJkt8Gogd3Y/lvbGsvER9HgtYBEcCjKJ6wFwMSmGbfrk0yfEuyYmMp
74HtKJ24ffbEzAChGPYXStgfc8iXKzvUBGoIvFdwoQUZzna2vQZ8cpcdte0Nd0vZ
lV4WBkHwX4zcokNSJXuJ9ImpuOS3AzRyUzblYgQ+L7e/orX7aP8+0JTmSIIsn8KS
jzZy00hQ7hNQhFhKdY1b/8oP5qMDLKbpLbte89WVqra6ehaD/MLiedfXDmcW46Cy
LPMHPrRF/DyOQEzjdu6p749FxrEtYZCrgPxTHRi8YJ6e8tkGeG7xI4v/Bnk4vOKS
L+s5YRRJ1du5cWli6B8n9pOAdayb+Xfk4iQWXK1RJ3PUylEVr+loNeOGNN0Ziil1
p8GM3p3O1hY3hKO+ig/pWkcFY4kJ5k/b9NHJBN56GekuDzQRJOoIgwU1j/we1wf9
cMUWiEyZE8ZkYwBgvh0cfkdJrQKvW7D584IU+6mVHiXZ4lAHnkOiy6Ia41U1OOGG
VJHGqqnyQOGgVWklzEehaqqqYVr6KbOBcQtU433W3cW5KHz+PvcRSqjXSkwGLZrx
At8OMWe9jD0+cg9TUxngs+yp2/nj3LWrBXY7GEP/E3Rk+b8DLM4LVnSRUphfEfjX
uBA4IVuZnOEW+g/lq3tUIS4OMOYjdJA1/mtHcgudRCRcqwUOr26wA3DbH9qQXyR4
wSZWDxjyeD43wIvUUnxKpgH5CX+OIDzwi1oP2VQLiJN2Tsbeg97QPxoz7QnagW3C
aPSUmVO+Uizu8r1nXGfLnxMLjf33hif+G01fumOoOiK1qfoaaJuRYvpJiJG6eeyN
dNIla3hVkVhC0YSK/FkYeW94UiK4ZwXh3IlW6xB9/HJIx9VjJppryX9gUw+gCyYk
It+yPHsZdMZhnkjVBgOalVs8VymUZOVxfFJ3YO14djbbQcK08Po+IuRotv16G+xi
pdUPOH1Kzdz3oz1ohhd2x2LkcKL+rYaN7Em/idgyW15YFD1D9Jcm3Cg3zsZxliIS
42yMP5TegRHNO3DNWLuAPQMg+E1x2swEhBY7v0UMQtpP9ETgFY7AUvbM1hPPwFC5
dzSgU3UpyUOjZpHVPKoatzrLhbsQC8Es2kSTRSODfIfl6zyZLgnJDzBBNXRVuuCm
KsgI3TjAdVSQF0Jfp1YZ+SAIA2z50tXIXsCjrnA8ukWda+QgvXIq4syxub3zT2mX
rqTyla1/4tp/qLf4Dn/cUes3Xeepn3IiET+B/YvRT8BOCjo1ScSVECM0GFzXx7ak
HOuERSGzguan+tw0vsrYBzy8QVKYwr2HXS9op8hIQxWc/0gDZ+Zhv48+jR/chZ2r
PkGOABKI//gGcXJlbs+HDC842yF1hRVQN+VnqWIhpiqQ/ZfpALxhIozlkLBpLk7C
6QDj0K+zv7l4LXF15nWhqZSbx64gdYlHx0YPHHAP1pn23pFC54CP5jKoQK6I4YIG
YWTBsHT+4dHXdGOKUwoaGUcY0jg9VuGB4K3tbbDjc3Ata7BphEpEUQPUkC62AOoW
fY1ZTfMf6czZ02lbVtYKRQTuUgUo0Wr1qsfYgxrbaoV/eL2q+o9v7Sbq2MTMgBR+
+8QqTJC0ek+J3XLW+WcKEMn7eQVmoXr94f+wDEh04ErkZU1SV6immbzLEMNCyD5N
tAeJ4IHw1zl5DnkltF6Fhl+t8I1sfHRDL1dJ1nAxYKe0Ls57b78mSe0w2wmEyHGO
RBzRSIFMG0aB20hVKcoko5wQ+OOAATr1E95cIadbYhv/W3tMWwwj44eipZKN8qWt
G0CPDOdd9jI2Iwt2bDnXPJMedZq30rFbbFgXLtp6YIOMu1eBykMdzN6QAAwvV/Pv
dWaIkOGFR1HelgQrVMAWPyRjkg1sB8tCImyUryFm/JkuQLyeZBTqhsZZCv0CvaBb
7BBw3kP0CXxud2xKVU0/CIE1pfuOXKhZXmV/yhOVnK5dANEa/v71T0onwcHPLwSk
oeFsOt54Wv/eBKNL0C9aE1R5qZG6r2zbK8IVt9n5qd0IL6zpmRkzmi9RJUcZIF36
3s3QMpFfVT3zvLk94xMntK0EYll9zfZ7l2HkC0OdHyD7gFbD8umU6d5X66/LFw+O
XduYk71dt/8Ww7EqPUrpu44JzjsozSUumILsUxAfBfOCFoWREvP3Z/EiVnDgVuIO
CmiLPyK4WnnGtcKzJ+0QjOqwtsX1SXh0M8gjdAZdIAldrVR4SUMR4LPwsOnk50Zv
gQ53vwcKM9tXQgPGBd171xgviOe/fH+6RxtZ753zDi4mOrxjAqkIX3VgBkeHiFKu
vkEUjiGtzufBeZYFwpCYOodBXWDRbg6HjqumFbSv4lHx66NpcQScQN+NZhQt/Wju
sgyJUHJ4fKt0WcXSNVwAY5BZSdo7D0CRrFnvJ+2kUL2iYaq0SESPqxNlkL742FEK
KIg89JtTrFkc4ANz+VZm49NoTm9OwXJ5pBoT8EB+CKWMhqf0e+tXkKeP1Rzr7AIL
aL76R5trKOsb5y+YUDCLS51b19Va+KaJJElznF78SoqEm0XTFPqSCcCM7OPz/3Vd
DjnfYqKpxSRvpYO8CN2PvZSntf4eDMWOumKW0RpP8GgpBvK7MzRWYw352mr/OWEw
YmYEJR4Ca0q9ytdVH0wf9jGfATzwZupjps13fTHXeiL2OHsslCqsBxNytMo8H7iJ
+KpfvrorlDgmhpWDsHYh5M5lyKUD/CeErEiwaXAhnLXOdEKm4Y36LzrQkDa5ad4+
b2NNkBDuB1swrWp0RnO0mCCWEVtQ3s07mDmvMn/QG6ypT/LMANAqaqROE5sQ3Owr
+tsATL5Tc1Cat2f8MXWjVP4AAeTT4M1WU7KtlNy/v2G4pC45sXEtQzw7Aeu1xKQd
v6IRwk3pzftjPsN3DUgfBpgp5FbFu23pc1549HBQ1LUMfBn/ycMg8QWwRPczAiiI
DPkVRVxLOE6au5iAK+quGNBRK3vzBlMKpp6mIr/hjLoSQenqR4D1yeznp4CYYwDW
iUkO8SEf+irjeR6s0BdfU02ZSgpVMOu8Mv7JzgJ3T0/S3BHHKu7HK+3w61JsSdvu
X47X1HBkCj6LODIj5bfhP6ZyZZiPOe30mhn7C4mpP7PL8ZF6j9LI1xOf23Jul55+
S5n0dscxv5MR8/qcXuaQwjagme+wAp7nTAmIR0vRRgMqJWECMQrSJH4v+FJmzX6I
EXJkgmEALdX0olUEOT8ABEurrUe7YeT5uy51F0jfGUP1grnYf5Y7bDmeLY/o3fuR
frhUfRybX0cozGEkYaM0afGsX1iCmqijTweQVWreLtOApV0xKXUyWt0TrerQszd4
8WckaN3OFJXOTM/VLFhF96T7xD7GOYjMOCzIQu3NQCzHQqKpziRr3lGNacNqTYHT
5mR4SP916QCCW67ew+14UrGFQEKbELIA1pJSenzm6uKarsXvVcZQ3KinAKa+0UYs
zqowEApCraS4CLO1VMKJBaEFEYi4HCB74azU5twegonKQ3PKQnAKe8yfDn0qGaes
+gNE2gakXKkfyFZ9u9v2831KDfxUbppH4Ji6wDLwVSjyg08g8ioFxzaBCoXWLaDx
g3Ld8mDD+x2ZG5A7ZuQ6yop2Sjmf4dGRR/Twl0Xx6/Pd6KZlD45L6hHx8I7Onv4D
J8cE0orQstcLbQSM8HDSPMk+2TVIFm65dQBFm8BrZIO417Pb+Afg7haBrhDNAk4k
6Vs8YmubQDyLT0I+lXeOGtYLWrm0wmwTIdsAvWvTuwDFFextMVDVKotwlSrl0k5V
xGRVcWi97UKUQkZJJdbxR9B1c2UfR3042a3NPO/bRPT2ZvFof2DfQd5paM6aM0YF
r1ymnv4UZ4CsmUTk+SrWtBwNHJ3AR6q9I6R4oxwaexAWR2tefWhYqLq/gtTxQdR+
xEjmmvHyNRRM1JpMGKNMT5/1Ms0FjEfRcYVPtX7bvZmAEdB5mYvuZ8A+6VgF+yYj
YQsAh9acbSDW+bMl/9iqCibwN4MP2w8AG7acSYyYpttaNMzmcg8EhfvA3WQUHg69
P0MA1z+5rP/e98OTNz0Kt6C2+JMQGoH/etF5uKxdSOIzcVY7xIAtIvT0a7+vuF5j
HoWBxgYpFEbOGhbotF9z1bRNc9Ee43FvCHPlP83jvqw1rtZPEr5jSN46GYOLeNJz
3jdMSVTregqp/69k4z9LCxPmnhZjz9Rs+hIhUOBCoiDIx5LOwXqXoUtljXgommWB
y+2+k+RATg9niT6bO8aDDfAC4g4PaZ6wIn9H0r8lgE+h4qGVYXGXvAsiS6yHMXS9
hLh1ca6saOqn0b87B+Z/OZcbyZNaVaUnh85zoG1lUTLakbRG2tu/VojmJIobo9EV
+stax4HtoHSw7vswrF2BXGD948rt1sBmqwnG6zHwC5b2APJfW9iSJ14to+BVGUH4
Qc5ATNluvf/aN3L65vOue9fEc2qg7AR6m4lTsY2lFe3fOW17xT6/NtAKwb6wrwi2
UnhgUPtxUE00+6/aKXmUsOHvGUUQEyerVZpXgde0J9Q6xl3iqU0Zll69aeHuwIsA
EBO9OrILyToBianahvDUKTG6sOp2sScp6Z4tWG/movKuc/zK8ooqcFHLT/eo2obl
jappuAq8QM51xN96cI0/yjW4wVdCl6onik/Kaav8w7akVI778gWd3iufB+d6YVKk
jI2EGxe28yAMNg4uo6ka8wspHWHTmILpHoB+OqlghfZ3voVpQ6dBzgo83yBhsy8h
lggy1WSSUmoaHjsub7qQqckG0L47bH4YfIx9XP7waOMV2HqBOpn/HwI13i4Qmtxg
th1wa2sl05WADbebw2NmLkNp+Oyld3v+FW/MCYP1tdVoEdL+VLZDtox8hmv87i7h
OwMYEp/8unZIIoHDuFms67SeLI+Kg4qslYJ8LFnRvWIZcn4ahew+bg700wonQ2E7
BOOpo2rFQRZXjsXQ7pe3+sCV9nOPEzEfnH1JsaXb89VIDnojVxSwja74OXS5xWcI
zOD+KpiUTkgE3XYpdG0OxwduWg0P75scSEJKsNSoe1Hu6FX2b13Z97dYIUa8paRG
siLdCxCwvDFDR795JGOlHhSDgWKoQps86V1wz33i6FhtpXGje0nMDd0kuoC4i2bh
zSvpFgwE4IylOfk8jChLXQsVVwl+mo10cnNc4tT1+CEwhgIE/vE2Ih0rw2i4/znt
qU/kTJXMGW5agNzqYbUtnxRDjEw/+x6RAa3KEQWFWK0Vgw/bdirugQWmrenvjjZk
+sZQd4y3xW7OxEtg8tE3elimz1pxjUZucVsP0WIApWh6COuKsmHnXrHzccC9ozy6
Bo4co0zCYBQQ7e6tt66exB2G0cA4mK8OkskfAQnABUCkVqtcSUb+zZIQ2p1XvYgN
SQRsOSpWAHzIeffSZwlwON/9sHRIxWbMNaFLZ/dJ9F5A6T379oPDeMf48jyv8sST
b8LuMfPGTfM2D9ytwVs7UNOwOoxO5lIa2pwZtRBmM8qnvOG+xgzhxNgWbCw/UrHc
uYBtqxyusg15b4rdkmiCnA9mdVEEGgjkx2fzCUlmnzoEKInP0hs4o+slmKUWXN/4
GgTCWi+kJDn4uLnVKwOWsz6O6DUn7wv5ZNMzxoOEQBuiFvh8mc7P1Q9gUPR9NLat
m+cOFg4rEjTzno0v0PGAlNJx+7wWCc28q8SA/sU4lyAnZQFffb/+75BSKNnHKPKc
4RRkyHSlAhXe0505NxQE4xyMolcIHUMbcK+5zuXba5dNwR2IS77cuRKe73ReD6v/
8SZKTXFoLAHm3fMq9ynJBw==
`protect END_PROTECTED
