`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gytpZzYMXkWbWmC3d9jbSeJHy/X6JScbLfgMgDRXAM5ASBWtOxgCPmGHt4+1iV9w
tT1r/mpTpKi6bEGn8umU3e7YCBuvDPWiF64c2EZqeI+m+T8xhf11UbA9lWBoY+Af
hAKwSp/klm0vu6Z6rhTEi1n3T/JhwpUHKncTGtrnqBJ/7C9tohwdUkryrB/NeT+e
COTkHnGc1+eouKbmlSON7fgikmjXCy1OIMZTvRg8SfyAcGUFC60Xgx/pHyA1HBkO
X8xT3fGcKBL4mYg7PfoCf7Q+VBhiET7U8movd2AM7ZmXxYTzGISgbm1AwpX8W7w/
/xeIgjO9qeFT7gJQilY/UF0r1sq6LF75wQ1WR7ltSJiCKalLVx2FyKyDusF+hLCQ
1WlKDsPhxrk0TIq1wB7Ekll2V/G5LM8hQVooFNdAy/c0a9lDoKa3ne0JzdQh2Fn2
R5hilvwjZ/VWmgIHIk0ClyxOhpoFtZswc1mcS2wT712hbrEc1KqrDVVhS6mBYHAz
y5oDx9hJqRBTFIvnawz6Ibwvq/lv7uRMuWvBkoLN0Dr6v+8iDcvFuw4Cdx8zPc5e
vQUMBskpSK0KLqNzFEWBmBhG2i2nKn6RVm5ZKAByFx2ERj82oIn7K/0qYmb+49gj
haQ+360HCjF4SQQ2nhegp/mfC290kBfqyf6hGrlbwUXlCK7oIJmfPK4D0vMay8+V
jcir3qTp0zr9iQDZpGk/voEM9qpR73/M/9XFYPKhLZd5rnxWLwiv9Sjm8pwoHNmO
H33kZ/emT4lzuQgpEgfQlOrqcF5DbOBSIvXWPf1OtlgrOtp4QJNk+xb1xhx94f3V
AQOyouz23PL0+ktIY6w/AEduA0PwIk6XqeRCjhGGhz4FRCRR4f/NDe9u1iX7KZmP
+EvwIhAg/p2aSpdBuBWq3uX+YRIvhth63/AogqMVdMMTdsydDMdPoUiUfG1slgjB
wrfevkTRh00G4zcYVEvsExRv2QsFeD3omESuAn2hiHoBc7/osd07IGOL+RfTvpD6
c/Hh+EQy6M17O6xCKouu7EuejAIPEHJu2qsehIDn3UbqfrXKaz4nbNd3RRyWPkwe
5EDVIbpWJEv2cLsxj9VfIzZ/dOh8ZSb2HW34WyACnmILYpGUz1+RJ3rGfyksh84n
Gqw8VnqJk72A+oUu6Wi7ELcUOYoh8q3IPIOLLeA5nQ5qQwCWkC6bYecy7VlCaRXo
wHc79/9T3MVTp5VeeBA27c4u5JrtCmxzZ/hU4xj3AJFGdwqZRohefTAwu2fv3v54
3YaLjg9+4lOcI6zda2v32AzAZIV/9UZe3/kT+atfi5GBoyVzdXpMEqTP3lEPtt7f
Xm3yhhXsKSzf4SIuzHRkg8ZxgCmYNGyJUb30yjTiLjfm7UrIvXZQTWwQ4nmkmYMP
YwncbiGYki6xaCULZJtJAph67q6ElWs0RM6O+SkIjHBoqvlVkOmemJVe+KsbjlrY
C9jQ0KTQyMNNZpJxahg3F7uOQJc7fwoBhEc7cZredohqSm1tmQowrwluUm7gv1E9
uKgqAAmKO3/93VftMw0i7Q5rVW4q+kgOzPModxms36Kaqb+CsIGSbI5x+SXwCc/Z
5vlKxcsYpIuJBYAJJBxsnuiI/bwttQZghEQIa3C2ub9HxiYzWp9qSOWlsqm6jwux
k2a6Uh/e1VwA/P0c9PWj0pXJszFuQUwJdx8/fW+2XzLdKIvk5cZIRWZhwBg1wY/g
BZi2JvlwyCk0iP0eAf8J8rmWtFkJNklbtvmRGaIfN4LzX9KT89Xwyn6ZfSS/KVz8
Am71XWpiqGJKQuQJa8SiCgS6dBgdl48Bs4uoACgepzoBjyx/Vpg3hOS5YVfE5wKJ
rd3YlkvPpGFkj7n9cYiITqrk5lB47IUersGpdofVWtmUnUrVIp5jQ2IM16XmsKMb
HWpd73k17vrjGVM6FAhIymYfBFQ2YUGaRw+RF2dh4UlF68HEkehDuDUl+ZjMLEVk
s7sj+vElpTY4Vc6YVcEzvs7hfNU79Mk4PHG6N7uys5OcizLdQM03zgTXJO06j425
nKfcRwe/rIxwHEXXsmFBh8gLdB02Hs6k+gKimBEcEGPyhJeHCqGhb4UBDHigfjD/
L5HNjeZ4AwWNdMEFO38zWNB+OcoA8sPRcT/84l8En0PqDVRN9u0y29qZwdtef1Ld
prNosFRqM6lPKLV7KkmIp/FtqHsCjgntrImndzc1HJmhzs/tNRPlhBML6GyhPzLg
nYwM9se8F5LHr3f81BIgp7rk/syNQXqBgr71nlmA5kfmh620SblgVchz3JhTttBO
l+p1KfJcq2pVKx5lbwgrKByPwpDtczRaT/odODztxoDPPgPICL+FuD/KJ1SMfEFV
qpAmupGkE9lF6J6bJIeT317xgSf5jnPtkYdogSr1vppjOWUEUsj5p3UxjIV409aY
y9+vnEb4X/l2w8EVq0FgD11QCJ3g5yYkSOPZ9G/ZJnYPJMQbTihh/MrHmYcZw2RB
Z9cbYmKoP5jh6xJl4fF+PGWDb48qDS1ZnDTK6KgMLB3wsA04OLOYLD1kc80oFcmF
c29kd3g2Mvi9+pXYEYzd05HhNduCmFPz/TQ7zEkqKUoS73eVJFk2JuJce9oFC2Su
BFCVTlRzrWcX/k24BALq6podsqnsNOuLkRa3U0GB++GmVLywYecaOzWc7IkVf9tJ
gqtkgfX9JbDy93smTnEXIlXdzA/j2pnJi9ulLzdG6ba4p7DmHXS8St0vJZ3yvAvh
+ORY8LjHOEdtST7iF7eCp9H8t162V3DTAGtu9bEx4bRvN4qA6kBDNLIWW4MYVj9h
OM/45+EGpWvPw6SzhrJqrGctSdaLUFe8XeE7zaSLZwlJCQB8lPHRcdu4gw4uVXct
anAffgTEbSMwrMSuoh/lSUk08XOvvYhYmqLFJ+DRvw7QOBIdAIWze09L9I9E2BDU
5IDpAD5+LQFskDKOEm5StR0IhduZFyVdQ0kx7+YSbiDgms4pnxnQv4ikv1NSLGmj
wteeA8Dn3JAcehU/xLeiSgbHL/ZipXntYgewsKP4ZCTwf5GwVp/azPrsOk6B/LV1
7o3LhmolyT7ZNpiD8/nZU/naGYvhN0We3lGaH8DydKdtrOvEHIQl3WoTezRgdssJ
gMadCo8Uja0+nl59YQdGEC66haPP0a7JivrOEMDOzuzAQRGXW7DCXFOkRzZHlYcP
NzE+fhtoyl1ICRsiLV5C6MmmHXyMXe2lGBndv+HK+7GGyt0oetYyeRxjCJTZ55mG
Eq0bLg11yfHz6fWZSqSyyb2vp0p1w4QK5EbMYXKA/vfloKMnTjYLaLkQEM01neIZ
rjM6EK86/TVfbcL6qAA4mQFx4tbgPsWATYFLxmzyvt8usJOEy4wX7naKuU40lJnQ
GJ2OvXpP7CTld2uHz/2tfKPuZ2S2qan02aEOfftF/Bg8GgR56tcXP+yTvzGpl6xX
VjOsCp1vqJn4tOuNMIGf4hBJmePF7nQCEM4sIrFoA18y3990H4cUOmcjQ7UB3O+2
vHkYfdS6MB25U5hRQEyaLQ==
`protect END_PROTECTED
