`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QAeU4CbnFZhdfin187vyiidjfHO9H4xZ/63IPc/8WcWoyBt8/AuMRnkfQFhMT7ZQ
LcdUZjFWBJhUxQ3Lvgd56R1PMNUwedRf10zMzSNiCwL3HJjszSM/XOhPaGlhIPgl
8shOGRwDH3NzVMNLOQBVKVVXuIIAtZ2Emg1lUNrr25MnrCMsOESODHHGlpoh1B5P
9f+tpsu/UO8LzwFjH2JWtOg6etDLfzp0Z4nKt8dEdunoNIwnY/MIcc6RuDVAp/EL
jFVc42T8gwBu0M090B6g3tBnTIMafbRGBtV+MrP02YVasgTA2XnOMD2cFPokO9mY
JI5L65YvBsij199loyub/MOOj6QA8rqPI5yi3oQ5aH29fHRBFwatLgt2DT3lEE4P
mwBgojuxo+ti4faIZapr0El/0fsaM1Twg3hdv9dI8HZYC6Ui5pNGWGrubkUsDdOx
gVc1IF9ckqVLclToo//XUw+BAaUdW95pdrd7bG6c7qgDJm2HT1hKVhm2NUCgs65Z
52JCLYNTjbYuROSBCPaNo2XeGpciLsolLCGe+yBXSM68ZKXiea/CJTL2zx6dJmoO
vFKRa5J3Bl4gsitJQeRm5SNejT1RmUnUw9iGzKfqZxd73+WJUpqPylk5fkLlHSPW
/XzKNCogrLx/16kHTh3aYQCkfuzhlkvl29FoxziEMupKw2Vwcir79HDhf/HPZqO8
JEkhiMtiMbJYojSHf3uCiSuT6qYeQbACIcm9ITYh6FnbWkY0HrX4jVPxm/nO3ER4
vZUOQsWIH68Hm7z1lhJuURSepIqOLZ3DHN6wzA83fi+FMS/nhV6HeOkxXdP75MOU
Kx8dP/89E8vTYRmBl6ix2uW2WptXasZStG4OAc3QSQEszf45xp8ua0t/EivKn6ok
hwm466xnVZxjKeh2LtMInBnt0QvDhPTpZf+7sQ/9dYQe6w3hNoiTgkZ6PWWHKYmK
9gZAqb6gd/GiltPkiLIv+K2KGFkDFO8wbZM8qbCZVtz0V8uKKxbHky3Wx3NRPScD
xDkWDTLl7nF//6oqe/NEdWYn/e/HWsOZDMpukTvQ8LMC66cRmou4zzR0mj70jlGa
bxTZGnGqmCnbhHQJAk/QboLVy5kXUaWWklRvfOudRuk47LDezl85ir8W/0dgulEs
Vd1iTh3fKSsnmPyu21Uw6x4aMBRoytw/SsqOKkrYQ79OFd3cfHqewJ6QmE5CBw4o
JL8IUYhIP0bvtAdBN4R7DoP/5I3guhGtUFQen/UIVMx0z6cGZKJboNcTo/mRZgSM
0Cqfimfjsk1a1jkfO6jRb8dn7So6u0Rz7Q44mGfNu6qaFu3eUi/wG3P6GDmnFKMJ
Xt6uhUntYN2DHmsGePUxAQoQLMkU4JVGWvYUcuzOBBSVebgFjHfJpL5IbmfcCc9g
01LZkSHSWuaAfYFLZ024cUy6AUzqqxCQu9OBs6HEWFm9e9svCS+YQMvpGfoF+8Ts
oRXwAHn1KBu2Oul4YXyu+KIE/2mc9YY8taaHqpOhmLI8FoMXaatbX3mBDi8aTZbc
50+200uJ3cPi1YpOdTNTG1dfraILEdE2eov27ZBSoMKxKxXjhiAPbosytWQdoLEX
zKoTOhmj9euwfrjDYovp9vOGStru8GWr/8J7ACWv4NmTD7pDrbaRFsvNyU40Cl3S
ovcH2K7pDSUenOGKCIjyM3dhnF0FezTHNi3S0SAWnFpUQbAhY46FWbJe6y28UvMk
F4dMNe9PthhkAIQ3t8MiBTrdvEVIeCSV1DROCZGqU/MIPfpZ3b8QeSqKB1ZcKryK
Lxn3jcRxj6fGXNgt3avUUtQr8Ij3CzDpTbS01zym1zsRl50vsiKCld5Ipzgcj0Pe
u5HY3rrqOU2KeW9NIfZxj16xknqNL3COZKCce2Nkxx0=
`protect END_PROTECTED
