`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MUg71dWbyakFyuYB9SsaDxc7UQbykdQGhbiK76Xq2VbtOkrhCgivJtYa74kmJQgp
ZjvkPkW1dJfumAiNJzg89tMnWV30Uz4rmejuJC6kaaMl/9n1lPAg4VjuICNH/14K
5XMG/IY0dPpkHk5w+O7WvTAneXxfUzLNXtfQIV3QyGsV1INlJ52mUmXihHJbrDYJ
0zWZ4TvxZvBdphO5sGUbKvWLtpn9MEhrI7zBn1OUoOHjnf4x9O6B8GgbtMWkaOhj
bVY1rKUYp+td9bZfIoEDjF2GzJOK4qc5xVVYS/kdFRs3piyha8oTWae2v25oIQwv
4JjE5bVubX0iWUUn/0sw4BzLff8dWIORlF80LWuqpSRpEFz4ZvWlBS73bm6XbL6A
QvTMAvN5k4SrPxX17Yb3TZ1OcFxBrRXRhhe5MBR9kFB9Mt4EZbaetKMhXwmoDvjK
HUnZS/FZ4WGJ3m4FuLbkLB8R2+gJnb/8aJpEEoX+naRdQKi2KhDBbKjNZOt0ajzm
kxy6GRMqMaL9UpqCoqklbw==
`protect END_PROTECTED
