`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EXCGONMOHQ46pw06J3+ZjszsTnw/swfkocyp3vbxf1cEejSqBalcZEjUJs+rrPT
poksEPKQuBvyif6Cs0ZbbIN+mEnrA2v4qkvo6+DQpHnTULNwDIwrnh01Aww+K8AU
qj1u4qL4B0GWQtrTmHjSkm/V4F5AF+ncfSvinFgcj6UBux2TcOLRvD89sGOB/3QI
Ssrx0gFEE1G9Dfs6lKEC+tGNtHtkZRkcnZ0UoyVhbmDXHRcVlvGUnvcJ1JKkEi5S
SMOw+efdRk3m8TApIRgNj2GyOabwMVmD8hEix7oLwsgCPhL+YmkBGBWKt4mk4O3d
hu0l7ib4+BhHUTpzxr+0ySJ7R5HHiWWYX40a7s7aXob0P2KTvzCiXCiqZyPF0TdY
Umd95A+mdFrpCJK2BAZm/AxmsBcf7nPSfReS5EzRWO69vM8ktckBAPIqbE2VMrEo
C37hqxbFRvbixJX9GnCuC77C3CTEsAgGAIRzIX1uYQ+wqf+cUkW5SlvLKw7wu/Xv
TCF4D3zJnkmMxCKpWyXxCVN6dYGxTPF87l4yvRFcil0mFPDuJ/Y2FKFb4pdEImxt
00pZv4gowh7QFB0iFU6XT/PkWhlQEVWAY42at3oLocrfmBIDpGUMTDp3oBIEqZ/v
J5H5up6nLUJ+JCSQ2XZdXlU884ZlUhD0r2mlyVJ6EpkQeReoFj5nTd7ESmadSx0L
9Mz2DfyDQJGrih3Op5L2Las0wojz2YEOup+ZGK85kcDWizmsXWvR+IcHls9vCAYQ
l2YjsTGc3Fq1OZzI+BJL/5bOJFLJQhRd5WNpOQPhGz5JYvMKT7wZt2JYoh9/x/U2
+76FDSk9Uorz0JECQmP9v2K8RH30Jz+v0fMYBiV3BTv6vTyy+dfJ/NeOvyPb+Een
t5KKdr50+iYFifATuLPnWd8HRDzHq3QyCwJQVcvY7UFXAUZuDf0BSB/IBRBSf9Xe
b1B7ut+qFPfkbr0CbaTWzCYoq6Qys8+iXa0pyEFY6Bx2hD80X43oMZPOUzJKf5Gn
y7gVJ3vPNlF44q7DQsTNfH3pWj2BpYnY54VToaqwmI/brcAFxL0R7L3IHjRebKEe
FcRzgH+1gFfMVzGd0AzbBC89DAM5lFyrlzqSzmiSsCPeUqR6kpWUhxCYEVpL37Fw
ULSUmy3gu98flxvVJyDCFDajIYfPTpTOcz0N0LW0A6qqWJf5ScO9KhUyNs2bSTim
T6wIZJjon6nX/XvscpAXPNdml56eJ6hWenzIwUrxbKfi4eN1aVJ+PaH7sEGVBFb1
o8tKM9zEyzbJnx0L9NubzTj84nJnO9rswdHy6mxClawU4aNKAqbzeNxmJNz9SJBF
`protect END_PROTECTED
