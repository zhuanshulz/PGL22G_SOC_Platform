`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YabBv5x9JYmQ9mcbDcC9GKKU44SsmkBcT9FfCCoKZ8A4GRAzx1EjKOSW82WWC6KZ
WPzzNgBotnh0ghjuVrhkpSLWLE5rU4U1JEVlavAE/wSZ7gtdhanA6Ot/p7dt92Ej
jVbv9NsPJWB15PDCO+3+MZyYdxSH8js/mVPaIwfl00wEJM/V/FqmvAL6SrtfF4iS
BzhO6/diX6BNvdHMzSpujyCeIPL6xQFg7ePisBOdmn1okhX0BpJX6guLkiwum0Cm
ToDeP5vigpw1qc8IWHqjWA==
`protect END_PROTECTED
