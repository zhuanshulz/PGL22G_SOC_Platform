`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qb/bFMnCultbuhN7aaLC5qRaDUcsj4yvYl+JoK/RKOPCktqf5Mo/fvKzTp92Z2sJ
ChslkZB34k7WCYH/Gpew+pH0EVNt+IZg57y9wAaomcVUpMKnIz9vhD9ooB9l1LRX
3kCDaAXQW58lpx4mJuJdmqiKPb2og+MHiuGQdExwgnNJQUiycLUkRx6qrARNb59X
01iRIgTVT+y5M8zVRJd/+R0l1r8tkCQZGp2t/jYhrs/ozMFZncFTVTyvbra9tyI0
d3/Gh98LiZBTT1K3hP7YhxAlNU63rezU7VWmYezAB1UGTdwgsU+VEav/WeUD9MAf
bbXhPEV9xLh2fBqVduqvlWUSqc2hoe0quPX2DWq9kXaXosGKcZJtFmikNCJ8QNr5
CeEOZrt2g5vwW2+0HxLmbBJ0HFinNr2nQdDrGuKuspHpWfUYxDLX1GnDgIUELVOQ
se9HyVsjHOrqR1HnkDWHmyZzDcFc7MNtMsum+WhvOsDebblId65t2rQUh6vnZEFz
iGPD2AV7umfvN4kw5BNS2CLDIqfwI/IccHPFoBmuXZOm8LtMqv2irmZlC0gkyZuP
`protect END_PROTECTED
