`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9czoqD9LQlPyTtMeiS2U5W7NrPKk4B7rlCLaFx1XTwe+dx52V8SyHL6KNDa3BMB
0RIQDObi8vRnx1HdApxeECXYM6KQ1Ne1J4c/MioxetF6kcyK+7m197x1DxoshfiX
ts+LbB9TdiAExLtVsHUFX6hnsR6MMR4XDri93tF0y2fM1TAhOda7yW64pSx/Rj2L
8pLeNM61CHGTSpZ1+dhdSz5Pbk6KerOgUFLZD9CVtI2OeU0e3hQ+wqhMrWbb3z0T
asUTkbBJ1TsVb8mQqixITBQ4f9Gg2iaiD2ibzoQzvQ7VL3PkTkLVzGv9u/L5cw7x
44EzQbGefilC6npK+RlZDrLA0o8q4V/eqyPVzvhdoXw/E6H3opkQK2qcY8et9aFz
qFbiddUMBGD1KbPNmla+XtSLyHAwdC0ykl2M2B7/FvWzTSeVEr83QB0foxC+akdb
QYuFpRIYJE1/kE8IMzkBEaMsrfgK/omPOjj7v6tIB1t58WWmSmSdY0miuRBDSlBP
9SRyyKTgWrPpfhYEkNvKB+ppRvw6G6dVIbVLZ7EtaRLf8Xnjz6d8yXmTX+Q2Wdn9
5syZ5zYvQ3eHOyX547xc1N+PBRt8LyVUT2ToqX1VJhOyQV5z2EvH0YJppLlfn/Ds
oOUQZbS/aYoijdI5/sQYob5pung4TtXim04+IfwXPNEg+cPUAe5soNuGCrD0dUfm
YZbBGE5vgy8Clizli+f95Z6qDxJYO7U1pME76uOkzVKwIkSAxSrPDDhqmFRC7q6q
NH3DriQhzdX7+t9RkG7RW1aFRyZV3sl02l1u9sE+SVJpAAc5R4pvnPY1nC/7NLdL
deLLLwBxeGSCEBDvjPCEOPXtJpYoapGwWeU2CK7s64hap/Lr+GYmosr1WlKkBWs0
ID51xJXSnF57Q08i3ITYjEU8CgF5DH2jUd6md5j/UTP7DADoyN575jA806ItWPA7
lgsN40sy+yjzPhh2TzY+fQpyF+N8gdlNd0vKuaa9Yo5W+k/GRqpVz9QJ1cjWmNmi
rg2hTmpKeOAytXHMPqiwzhH1K4CUrv8OQ8qVILm/2BNLAOUvMuK3A1xGYSn4S/mB
GumDniS9NZVUVgwmYEi6bAzyORixqlxJrbNud7uVOF4nwWlL8664yPU9P0MUg0FT
wsyaUqFK2zqSZT4vLvDOp5oAT9zLBzHJKxi7kSZHDZ/6g/ZuWEbOWVO2qRZHg/Xq
kSSwQC3F0cBHt1oXSorw6Y+OVLn0Vs0bJ0TVtKvISlNVs9mPgX6DGE7L0KxkrQ56
HBgFXLlJgKK40kGo1ZEHsK/J+JqxzwUl9NAHvEYVlZ+6tDdCfyNytLeiPBB8KlwL
Y5JMYHSnSPg7o71bKS4UYRHSQudAEZ8eKJ2NEK/oYiZ2TXHu+AHLxQKsExE2s+n0
nNYOyIZ78lD/ymzKb2j0UkW/UWECR3VTKV9oEm4fxXUEC1TZlzfGd7j39tv/Asdl
AGC8hbcVfCXpSoCHUG50QsUBr+3B/jxyDHVlCcnPDuBRz5E7SPD34sdzMz5xjcwx
vK3gy4MGnpjNNwSlvUh3jOrUp9owgygSlT04rdRL/8qGN6384jUVYjELMR+dGB+8
l1g4uywdjw4fb5L5GkYwwhHP/sM5orbHzHqiKLLhSW322r1b9KmhHzUFyhsEDT2x
zSHK2njdmLfNTkwoi01IZ4NllIcZy1l55QD3o4qNWBb8Udqh3P2fWczVs5YBwAG2
mFdT1vVI5kU/+cNN0QgtIr6O+pf/B8/N+tTuiXR8MYvijk8UNQOWnY3T8X+qYLKV
eIsvwZYJx8H/tLTKkvynnIyKpq9J6yA+ehu7aWMJS8Mf6v8CQAJCVlfX+7dJF+Qz
yBZlZ4Oak/Js5dVonSugvjCwHJtdKpnsF3XJVf4xRJMF+MCbIAXJuGWJbgcP51kJ
l2LYLK0HIlvIZJEYy1Ut7Y3QKe3e4krihZI2oqVnvEwKfw5LRFsyuZJoWPDApFSO
gorQgd3On5toHA96NMvNuA==
`protect END_PROTECTED
