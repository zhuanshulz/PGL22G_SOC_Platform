`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFK0HBEjMJM+K/+qJPm8gyRZgaYMqo8qGRRE69RR7YLB9pzFAqgwx1BJ7r90TShf
pdXhvC/198oEe64yWS1zBAr7jMqKYpy0BRb7WPShMJPSa323fHkXZ3/ewnXEE6mT
fgBCWwwpNHfFEiMmpexMMHvRn6ZYqgfRGrJJ1MHAYNHaqdFCbVzWYnDryZLYz39J
lv07n5m3vKsuT0LUVS7ygld8EOWQYxBl8ZyT1zZAc+y8GsD/KCuuK6dmxVOi6OEz
JDV6JqEvBLk1ewGHqjjjyffM8KxW+tkFyxUlMzWjd40BFVkKbWUKcreLFbfcMW58
/9w91vl/nFJ9ThAuSjg/23NkalK0a2WeDPMu15ilLSWcpvPc560g2t+8VU1N4hCa
uCQSHxpRUNdYya5T4dQUE/pk7ptjyLQjpPcJG4s7B5RnlBraFH96o4JqQ4d9rZor
4roebKEoEMMfu3KyRK5F3yRsAMJ7mgsUo96OEo3VYxBHOqaV1SeCiRmxLem6k6qX
BoA5YL6bni/kHwtRcQNEnTZHHybgPr/xwonn3SWjD3tTTompgK8AlpLhRGMw/Rmk
4csY+H9BczNXLpRCjiT7W7LvA0YPkAohRLSw+PDOBAsyglGg4q4vFjHXQi7Ru+zJ
2KqAoua8eRCnJtDQv4ttSGP4U7DcxE62ok+qKlhXQNCgsvvsTMIPT+y4Y45l05uL
wp/McbTLP9lxRd1hd6/D8ob7VM3fh9UAD5Ir1aogLhqPN204wS+BMox/luJUYiJc
RTsZwMGSfbS/ZfQkf+S2RdH2jfHiKu2t6el70JF4WSfpeEAUqpXtypI/dPHTs45J
AshTogSWDTzK0WDug324VF98xVyKS+avNvPrXibT3diu0U0YQ1JVZJlbdAhjoaeL
20RVObPG0CZJ7ScI4V/j28GwfZ4yHTCJmCtG6N8nSLhTmLDgTbVzKeHUu/S3ISBQ
Q3fJJMV72Whjrg4oeQT6s6V+ulWTgotl8QKAQSe4d9PTRUPV9yKac34by3+AveeJ
NggfbovQzYSVT23qeitktV74wTEMHMOudZWrJ50PcsIjNobhmA5Ou1AHKGfcsQY2
NpL4fUMTsC2bY08oMIfE52Mt3hPhzahYC3MbblkW7F5WWXpoR2U/pb1B9aBtlyAz
4lFJBPT3z7KVGdfK0qfDTcUMNRexrhn5w09hkz8LgWkJM+xDQLr4e/AmZfjC82Mh
hDTyH5FfcY7i6TbII4Aq9h/t52h+g5JS+RYZtOqvaqSCuMZMvSpWnbKc0gsed3mx
WID5NHULgXYv9wNuBz47jOzY7zE6XMY0KTnFm7u8lODeE6CzQ5wkd5v3XSd8ewLn
qsnqps74W7TtYLDne4NxhQF0JMwNMeUf4TbOqteL2CfhATUG6y0l9lEDNNlULcl3
r4WgR+vxs/9H4NQCKjIUtui7522pzfX3p9SZvMMqlFj6QvT/OGASvgHbsu5DUho4
Q0nkzHJrgd4ozHdFjMFtmyxnUEXgazlOexsreq0uXEcxa349ZsiCohyKDi3q3wN/
u7Gopz+EICxu5oo6TrsmbIsZRjrXJp7sTO/LFF0HSihF49T3TvcQtKfF/0EbuDrt
NQd18DMrbQoXwkalQ+i+yqKAfOhf7BG2t2fJYLdCTtfTohDGicLrUubnqL4g32Tp
PypdX52ICz/WUjPVJtKMGEEw+j50UfjmF8DcEN9i/r8rIrtCZ2pCv199ANj+7O3w
kqdbX3WISe449dsmPY7GBdMK5RIvDOfLSI1jNYR83wGnJOqKvc3Jo34JZGKgB7EP
D11imzE+CoXIoPgM5UKmLNOrg6Dny49Rxkp4iXoGLPIm4VnTWq3fGmTytXT/ej7w
dKSl5YuWqTMMTyqG+tTeeyLpbwU5FFE9pO2LPioOVMCYPcTY0nKwcNa17ZYovfKZ
bajhtJWcVLO4v48XBmglESIXSfuqppIjztGIPFewFMbMq3eopoYOF6Wk+cBpB2Hn
a+VSlOJl+23RThqSgFpZvo6+UK5aC6rDCnu1TtWkkD6JeTVJ6hV1sSEiWPLwb7Ip
6fM2A0mssGsEIomf/03YYM58yxM4zoTPQuLHfCVRZoEz2ta/8drGdSuRHja5LwNu
H0+OYqQ0dza0fks7kxIshN0gHlBd2lXBFHNj/McWBUjT7IR8RCcxw8k42SBb0IIY
B9zFfL7KoHfcY651FGvfG2+MFJI/8io+Afo0vtRDEccpSByg5mp/zZvRVtbiP0ZP
+2awTtAWLNrXgL8hEWmwXELr1YAiziLZ/HgCO7qEdDyltDCCHVAZ+YxKFZj6xTmz
pw1jOM2PDABjGU4Hsd2fgJzPuJ0k/HexTCItUzGw97Z17EGAgpmat/3apg2dLvDI
DGo+E7HrAYFrtrloocdTQR7ZhI8yhxkZw4+Q++l4qSZJR6YbdZiAU5B8Gzfo395m
wPn+ugpJCmBTAE++L/WqSz6IiWWg/Ghvu522aUVL6o0L2AULV2MAWSuomXh1LCuz
rvk0Subt+C9+Dzyxb/K9TJoxmvX1LGk9O7fKJTZZCXu08hYXYAj2rcMxb66y5Jgu
3m3Sdoud0Vt+C7Jd44gKoj3OjT60n72X9ZPypalvlqU3xuLcdeo1P8GciS32hjJ6
zDBu9mIEUuV3SISS03jtaeTf4R5Yk84IfzskNm4v+29wYipBUlwe3g7YYljv6fN3
ZZMjS+EzyjiIeEFtgMqHmfcWUtpw44yNEdpDVK9yTnF98+wf0isI6RqhU1boF5Pq
eLH1sxShkdj67dC1uBRDJ5WDRhCHr3iPIyKR4JiSBva4IzQlnqaW0CwQ9xTNu2TA
pqzIdgMfIv+3+Y7hRJOthEww4xruBKYbemMtbmX8ErP+KFlgnJdUJbD3asq0Z5I9
98Nni71wUYJ+SkOE1s2R+EVnJDcgFlCtdoHGtknFGEBUthAC/Xm6bex+f4yduyBT
8x/tGK6bvFsRdQSx8UWgLU4nc1NZCPX+jsSoC0tZ2/zbiCwlUIMpdFSIin3BgF7Y
vhxUx97VmEgLPZzl2nbY6z1+H1G0xO9O5AL7nI3eX8xvmoa4ELSRutq+B8ND/BfR
KIqhXK5Fm1UmnuDE/X9uK7NX3jitvD40tGrBPPYMXu8i3YsFrGr6wmJYs0qqZYyE
sb6mJLYYC0M/2jk2EMSmCQaN/VT8eI/VCjsLnDF/rUjFoGUuKUVkjYJOfJVJ73p7
7gevKFL54XzjVIb7LRoEwgpX8s6gGtPapyp5jONXzIIqPp+aFowfphn3JX/FPJ3D
UFUFVzh78YEQzFhcqfnDQVcAci4zQLAqjrjbxpoY3lzcx4gcZUsm7yR0FM/dZNWG
1t45kiMSfSJEBbEPvUg0zJJR6jWTyyokwMM4NN4LqXZHNq/oC47cwLb3hkijEVF0
/NxQh+vGcDE1DwgSerpS3aOa29tvT6YFk3rImSDf4niQSKr8G55SSBrIH4tCapXx
tkSqkmhKERG/nhcR8b0g9jfdB8gYzUTJ76d1xQThponkTQtZeA2FJsiYzHgeIZ3i
ckV6svwrzkLRTyR8x67EO8+1X+KpUQloJVO3JWT9F3wzuGbO+Z/uPS2xhbcFWkBv
urovgXXTOEgtSQpbNdWMQGFf3BAx6fclE/rI7OadCmn5DZiTNVYXjPRSXWE3xDqv
LDmfAza3Dg+iJRkS/hdjxRau+NUjAlHcc7NfR0pFNW7lNuesNiaDtdysB/WhB3o7
XsMyu+AGh2lWnPGEUzJ+HqmqBRc7OzGkI9X2uVLqvFCXNGmhsSWq1qdUDM4Per95
TZSvhFaXkdEk4w+Ni8NuC9mVs8WDCAt5Oy8eDSqZMH5R4O5+5X27nie1lATk6DCb
sNwec4o9Fe01aPh1XSVdiCHfMzxdTmWzuayufwWXIbZYVJ+lZFursYpUL/uVlIcq
z5UjtjmpyhpZPNyIJIv2XT76kkzVm1QPFB8+liD4weTefu8fg0DBJP33dywxhvPy
qu9GGyNw3fVLU+CWo1nOVrpehCpNS8Y7z4+GKR5dxDhyCrCG1avfJ+1sDYrf9CUl
5sCoe9Qb7bE71+FClJmyU8NHIvZu/Ww6Zhiw94KXhTaHXSTSiCMFB+Q2bJSgg1Bm
qZCEHi96f/xJB82xShdxD03Zyb5WUXyU35FXyX8idNHCjLGP6FfUXKDlRQNLJrg/
3xARCoFBIA9xMSYxNaJQzhSC9uLw59b3VnTBqpT6Ox67+0f2PEB58DK2MJhQwQtk
f31uKqUDZ7tZNeYaU17bav6/3Jxneu33SLVrYqytBkc+XoMsGZP/saeRJQ1mQprK
W/N/Ot72qFB3Upy+cL6tl2HCAGxiENzhofCtBMyNJBhIZeJy4vZZwYVDX0GjjTJV
dzzp2G2f8cfoLjIc8hzXrc2V/M/UXJRTp98AlBm8cztfQAAvjBNc+fxPn4ij5R9n
tQ8rWdMb2n/HceKbaig9l1MWjhZBpnUuTz609Ks4eA7sAvIcsJFGtXaorcd/VNBI
UV5hiI+QBWyJsyKdUwDIokYquWq6U4Sx6a7MaUeXccw7IJ/7otlQKEsJRX9JZL5f
HbFFKy8ZVI32O4jkRgROUBrVeYIrwfJ9pxJWAbsyd4GkN1tVsH2VirsYUoywMHSb
8f6Ohuy5rCz2go/axO+d8oKpljr/ARjpIrh1e+OfA0rK9wM2+7I64D20N9eVHZpm
f+xDwvfC8siJKCqWNOA5NnR2l0m3nMu7VkiTypnsR5ZRrNrklWw4NBSacDAxAVIA
8gv4TrDZoVNW7vhfjgZ9is83IFsjUWm2iDf8EPdF6Rts3i1P+OO1lGAaDp8dfbnl
I7fTG+YYIu2UpGi0fLEMPRNNvFT/8C9mu0UDYNd23jJ466dDMKIj7Ok/77ci8EUs
t33BYq9vynIXqBi2mwYGXLuLUz9wIYNB+Hn1dx6ipeK0H9OzfCtMeC8VoER/KqSM
G99yzVSQLnpKiSvxGnU/XZBS7kDzN9In4qZL3eMDgQgEub8ArLQg1iMTU/mSlmCW
Uxk2yATPriWlRUi+mpbrReI8aK/HZAgti9VEDivf/EVVJibNuIHeM0sG4yHrDZPM
e1Iuhnru+Zd5v+e5NjjoMVn6H5TnCMpzb5iXlt2+QhiuNDc2+RSZEQFyypTf9kwd
ANCsvovRlHbYnU4ZfrQ3Z3RRoXWJpItR89cTK6QKzVJd71zNoAp/Dc0YFzwUzhg1
4q475/Tkrzt15OhFI4LMbNsi0OjQUc+YohsoAadP9lDvevmMJ4xDvkobn/SDl1oW
+JAO3syl45l0SMO73FEDV+jtvZKHvoaLGvN7qLM6f4AP6Q/VJ0TzFlGDr18096yl
I7iKF1MqRsD6CWmpDskc83YmwsO9wnLhFQyRoGrfGU+D/Az8hHJbIYPTXStQ1VGl
sA26HFhODyiOineIDj/RXsgwljTGeAuqpsu+0oIne4zCwQKkDU7jwf3FghnxXmlZ
/wwnorBufjNZbR+KfxE1QFtQenNK0UjGZHIiHRadOJq+Gtr6MAeui14VpLx/o2jW
+nksUH9Uh9F23/fda4pbTqHDyztD8qCJyFL8nO9/beoiWf3+QUU7mGt11Ytn/FIW
eIz5CAp3rjyBSGg+dVtSP+jgeQM4Y0CmD/bsU+q+3NCvndAkTmc5DYn5rmSsQbsb
uf27Bz6QhOSwWA9S4Wo21BYZ6POmQkQvrHiO5DnakT5X1G9FusLTCKljSegwYfMJ
aZlQHwhvMod/EJcR8F+GL4zl2UglScBGoKwv54lfZI6E7IFqCk+pdciYKadfnL+d
xx5UcbicM+JkQnZnLEGd9etYXMmzBzIV+1B8jTER3bMOB5rTEUW0vBkHAEZcSola
JPyaFb+h9j05Q8pyzI0V/bp27JYxWmZhBI5aLOGXxYql6s/QdEBPbEOGAHnFOWG3
75riNepgXoS/Vovp+D/1ibcX4igCE2HeREzLPFTwMkAXY3lBqUnxcfS4biMMIoME
ezNarkpfLKRFLZcB+9w/hHgiKXpuGTpwd6DcGokck2X4zqAKQjK1GtilUHQChrzP
I6SLwSKqot0afK4U4fVzxdlb5VR3b4mzsYZLgui6e7gLNUx+llSH3v/UX1RAiWbo
LrkpfptDiUKfGItXbr35KJ4DCvsybi1LAgmOt/uUl/sm7rq01GiDscUADbweKOM2
N447Hs3HimHwKRuEjgiy5nxgZ0V7RubDdjoEr1A7nM8yEh3k6KMRU7TykbpjzpCP
nRLF8izw0DOSaqXF2FEwSrTSDWvioKhnp2uvgYVL9dGRiD8vnOzwSbq2R/ODLo2P
PVh0EQnH5fBRf9eGzvr0QHKNO5ipN5JEn0rvIbk8vA4HzVH0TafwuQEQtVDnRkWI
IY/AOATMuuzwxMYm8w1dY+EZy6LO3mWg5luBedQsFpgWPDOtD+Ol9peMB0/iVvY6
kG8yxc1L9K8j0zQgIN6vnDzXqmF+J69wK63vs4MqYV3Xnrov/+g8t8ViR2tsJfup
EBugsxvpyPvvfivKq0WHnaZ+qsPi8+tKTeoe3dqixHLLULF1qCJllUrGXy1+tVLq
MlrEov2U7UUHl1I0tzTf/4qDl1D2x1AGBjB1SeFzn7cislOHo6bit+kLO+ExNw7d
S49w+l2M65x4M4rMz/D8Ldp6ibegtJQEB/Xj+PBfusvR2UtMO44GAYEq36LyvNm7
0O9UpJ0bDL5gNelrLgYd7oiK+Gh3P7fHDcwCMqM6Xnx/TutXmdJT2FD6Q9I9ghE5
YNEupMqPsgSyM567VUf9SZAD6xJLJmBojRplti+F93LT7YbISxVpWMM2MLDMzLrw
HL7bmtstZk2b9hGBeuLBMiPIZ8YzsbcfExKR6KC+p2xMV/talX8CC3UgfcqAXTBJ
6BGHaW3pJsjz5ia9o7LUm9cWxTjYlnrwTNFLhQaA/TfcryUjeDxxD8XMaj8n02Qd
zEJIFvg1hHflpCPWPcbRkYG/NXvFWKd89q284eoltEqXD4DUJ2yf7FssdtgefYqd
BWTGGnQ9gvrf2WHRXr7qW3qEekVUgBP5c4Uwr5w7cvs9RvmC02VOUy1BPDUWZ+11
lDZ7dME0K83sJT4HE6BaiBL65HUdxSvS3l3YnlaCmY72nDslqtUZkKItova4O822
m3e5SUsZwe8tHp7nWDEDGNfQZAX0sRv+jRI0zcn02FkdOd0G2mYMTjq+cyCYhj9g
TikiBoXlLMWpyIfX++akeJ1iHkRhJX1fK2MmNfo1VVJ9LIgLssNE070PTXqf4VcY
IisfW0wMjcBo2RIhcnADM0f7zgItcjhG8sPDjEUAhX4QjOhX8ixnPnVyAAplwR9e
bEgx1h+bMa3BeB3ujth2a82cgEPswICzRnbRTyM5xR4ulqc1sYenVbp8qhbQahLg
LdOULgcdl0SOLBohk3/4Vx6Rzp8tGXGt1Rm+xJKq4bxaC3TZei0kOOY8+nGSymar
ZAAN7BhMO4Mt7UJLuP7HiI4fldE05+ohmd30vXmGtAzeH1v2bWD2QSUJzUPiulCq
q6OfENWRZwPD8wIcZZ7XqtizEmK0XcuahnAFELrxXRdDhTSZXyE1ogryYTC62MFk
Sv8u4qao1RpjcjMNz3jT6/ugnMO24yoOkzx45z/yDiuaFaj0pWAUDC7Wx5HZxMOj
UJcJTnc+9VSr+ZPY2Qejq7mqobctbB3WzPDOZxawLpt15ey0kOXM6x9DdJLtha7T
iKu3PnCnKiGZaKS3OizRNNDfjMw9Dc0ilaobL7P618HdL5LgBPwF7oAe3l6gLTp5
qevP5NzKpt8nKd4oTwHu2IHxfvWI6GXc8R0qzbC9IshLFKdlzjXDnq5rYFXqow6E
2OZQHU1W+DH4LFJ7/3oSNBSezjdKujiv0uMnas/jsyWIk4wKrym6FC6y5BFy9NfM
SucEgFF8kIHKevOVe8wjgYLCbngDp1a/4pJ4OTZUUuINDcPer0Q2QobVPNsLXpdu
rDrGt5NTyg1wbD08JARdeHIwYyX4/L34OUh8lj1PDlvxPI2I+eIKiFk1XO/bl6wu
Peuk7DbjqQCxkln/NR4aT7VL1A6TNn4Pc2hFReg6IL0Io2TCrHhbdGSiDSXAZyIq
eRGP7e7DIR5ebDsFeMJfTbOAnY3+BFCzdWF6EuU+4UUdqc+X4WYM7ZKE9WzCH1rk
WRJiVEmLSqBUJchFOydrNXpU0fUQmReYNIPIcm7guxMReXoXs83OqIZZ6fYUwsS+
kv0ejaJ2dHEvi/fFYdA+Lb27NclpsogF2Ho9eFwvzo1WrFAUMmZCKjQJ/GYe+9JU
fE3kuI7MS3QogcgkVH5ajdkgvXhkO7IhH84Tdj4g7mZpjHZEARaaqpe8rJM5fL09
so5E5vyrABHv1ryH6qCbZwTrHJIHd9UgcJcurD9qZJP5fa08744ecCDIIH6X2JF7
YVbuiVZJEc3hocovBp92pYbjhPoN0RW3ed+BzmHc/sg0cttV/fYjnBic30wXWWrQ
nLvQttkkVtqgF1MvLuCwx6mGxKweD4aHUQzUQ0qP4iMXYIHY6nYLkqgGvaMmAX0J
vZEmHkDZxuO0FZClXhLL0fr2B2t3qn93NzCDlayY7BGoy/vxn1x/zOX30vx+yK6r
bkJsNEataEHET5s5KO2fOh8a/POqMU8ucpxteW3mQepCPnm8GO5ADe5muxLCQrVI
2fKdjyI7hDyIPg1so+wfsIdkKjNNO331AQgTW8HPrAw4dnQYCUwt9MoKDXTaQ5OV
6B/Ayd/0W2ge/A/Lr5rKVDXs4ZBduM9RbXuU066peK9jpsz15kBalBILKXHt28Gq
CA52iXB/EQCXyxu6VIgK7K6J3mTnY1itdyJkpDXSgqogaHg00bn+h+obYqWG/Zrp
MpjR1u87o5qPnGoX2RdykgOBqBUF2qHS5MuKocfAc4wMbIzYzwl+BJF8bTD5Piki
Qvrq8K0hYgA7rno+IglffGLhDax2Xj6+3tHE6jf6ZLvJz9ApNT5iQwB9uudgRbqJ
2ef8DArebpcfjxEl3iqbRYUWOrmi85kzu7SquHYFRNuZ/M4LMXSSJWlyqSR6hOKl
2zGkMFZDPi8NRHadv62Hvc7/ZI9P+yxUKOzZvKd2sL6/m5A4IPjC+q/9OS6eLKlX
54Q4LOzzwBRgB6cNqOA/suuoqtGknYwc7srgVpeQt4x5MmJVG35ceHOSwa+N6E9i
xi3A3dkKK9UkjKDrt2A3L8kBKQu/eUbNdgJxmI3rvef4+WCGPM7vSAL0BsMGs1+w
fhHEaDarRbEOx2PAWe7EWMVHfCJdH1x9M+hqjpeSxZmXWnoTtt2BjlBuQArtq8jy
qCwXRTXbX1pnhIPu2fjBk7WD1bIH89ztKvQTwVs8SsU17hs3O23FAzNSCqCWa4p/
WqQJEppDUjXJP2nAvR3nrHOfcX26Q0qZGHngSFWA9fOyA2MQ8LA4NHxiL3PAuySx
NNZJ2Nrn5XqvMOTnDrU9aFo95m/SxdqHrboE1Ex5ILpjHYYtshUbedvhQMgn0BcQ
eny2x38Kr3hXMzGEBRkiNyeJOO4kPAFciIGHHzhxV2wgot6jG5VOUAGkaxeNKd1x
AP0DBnhamgdu/cfFn8Hdb+dGGv2CkK/3mageT8m/1kRS+My28boZqEL/wNJnKyD9
+Zs4mQ1paya67k8WtfADbeFo5GcE2iNuKZQv7ZfX2qPFIcEdIOvEFp20Bo4eAouO
x8tn7rbtbG0TeblNCvkEaZA66YMi1MN3LURYHOOVH2tkpEFbIDsmeUB0msx2nhLY
z8mK7Vx6uuM2bMfVuMkndDbUzL0B2w5mXq7jUVtN+cHp1EchbEiAcx2pa9HRIWVx
XwOda/yHG+83SJj7btl8jGAkXQbKcoaowhbkpVa7MgTS3gF90SUpH56AeJmWTcXR
AxDT3kf7soicNhbgNAS8KFvego0iBW8oBP6cKBuw+3Fkug15q6LisPn3c3wPHIDu
vkCDFQgUgA9rVcW7UDObxgXleylSTnAAI3DsFVpFNvF73iiTRm/0sjwIiFrbkjIb
pT6hwATEnOwKYERkWETKFigplABNLejTUJGSL3GtaMfo+5d7ghpZEmzs80oXfkje
Yr/UlAY9QLyQdGmPdgoFwacot8FzA9fqf5p3xSFaVwweN8V+N61YfEXCy6KeyHxo
/GKe1K7HKac0B1qyhW00mT1wVv5XSPkQI3qxGcKl3c7VyQldTetJNtBr3b755XgT
DKejW4+w1KzSCB9nlCsbz5HLFx/3orD87YC9CZw/L8Q4H4H04IGMSq2kirlIoTcK
Ej/ShfFgfPbtiLZ73Iakp8FJIakR6VXCttGIMjL1Nt41uE1aiy5rYqtkKhEUtCrd
FkOJ/KVJ8LZydWVNfXb0pdL2Zqj8VQ3fs4ymQsb6NMtZlRlzZwlWVhtWkbskUL0W
o+gXptizkEih36Vjk8IY+TYSYDRAYHAxRgvHSL9m1u0ahsPD5sK5Dj6y8ke1IRBK
U+5bujVtXDH6ZfcYlWdyIQ2xjdMEobhlmFZtQo++geoRGWi0W9cMP/5+m17S0lS4
+stOC21jOCxt1wWtJeP5+xxZD2Lags5yGyd++GGovIOsbbeoFV9Tq4WQACcnCQhd
F5ckAjOV8vACjrSoxjrxwSCLxvlcOdsODGzJCYhG0zLSEJSoid5Y5OfTLQH3Dbdo
04WLxu4Bbr4AXL40XRxXDIabQ8VdllmCIGXqjtPiQsDmHzkgAi3L7MjNAGpSOyOA
1gGiWMvqlE5gSIghvPGKkKOqXx6y4Ta/1T0+2WjYV/usxW0gFHb97PMW5R76Ziiu
SL4zjdxfBpqM8n4K0WAOVEEyQd/uTQtMsOOLPAPOfk+xfnMtxIvQdndBMYOJCDge
khKFwNn6iFXPiXxQzJ/6cXCg20YVuMFI7T7B7KaB+1yiPCKKRjAMIiNHiieMY5xS
IPp5ENgnjweQIUjNYQ4U85Fil5RDHN9m89HjwT3+w6tWHnv2ojEnI5NHV3HBN2/W
zN6Dth9kx4vqwfVG5nJJvuyu9a38Yq4WIxawJKnkmCEbkTa9KJDULlo9U2P8SYKb
w/Nm1V+k+dG2I3JqaaMS86e45bq3ZXANKw1kcfMnhGDuVWRLeXPPRR/bZTIaThcv
VV7rYVBF+Rf2qtj8KZoUxs9IR0gNNBoEUj2ZNtjM2kOvTQpt5ByjHEwQcLy4a3Kp
C5VL+lWinM/JGdF6b+03EP0DOA5FW91yxtY0GU216rLmIhKAMACRgTCqekE+nNo6
VgtI5NyJ/4vWerojUPJ4tWeECcwrhBW7UlN5Cnqb+4tB7TrNvuXP4MPrR1HPZEhb
sk76XZnJmmXVDsP79HiBB0Ksnd/LDGgifHQnxdtVxWJskNTKAWzntV8XOJOsY+o2
xykIBG/R2SjHDusWu8yrYxGiMCgwr9iPSgSxNvTrxWgjFW2BAt91RLBZFIJq8wOM
NhvcoVScxd/SQAibimfXv7/BiGPb2IDkAg0z+2zv0uClOr/ncugYzhv+EZVPZQUl
xkCIYLE+vDbg3evWM+HI5D0T17wqEEfNhLcihwlZK7yJpPqSbEiD7Ei39EWJlD54
pn9oEX3A2woIQMFgfCd999m5+Kpc3SB+swTyjY3ayj0d2i0R0NhdWxz+Xd2TjUxm
JvcFESNC6E1w66pCdClwTpeisJ/KwOa4UinWmdaoGskLopd3HP56IdViBeRhPq4E
TksaR33SfCAmjsY3FlUKH6AzXgX+QbDcjrOruEAZbp1QFy6joRMyJWZyrx6VnSIk
ihRH38PVv/vHlKuI2TTehXXf15psVnn4FwOScRbePAd7hkEHKzKKD0U/i2mHQdvW
+uswsa8UpavSDoM7OiW+AfLhX1jp0X0ebJ0UxTizc5rpthbtBVA91NfUUc3pZr0n
eYfXRLhDph9bOg+0vxP0hynWwygYbvAuIq2MgMvtJ7PE9tLtpw1ni9lQ64TIie4W
wTKP036erxjhASnOq7tZMicgArgOA4XHh8GAOkDHe4kzWFTW8gSUD61NlB78GWVp
MU3yl5msThkIyv0S9drRWlO5OgXvw334js3qnQC+1UYdoi/pyOoe/Z7l21St06cT
7OmF0wo70ZaHtuorBX2Glj7Mp7TQYRD82XqopDfaMKW/Q5+v1IOfsx2ebSuNBv5K
hCKvKwGLXqb9jMRwqyH/aL0y0jOf5s7PDfM7wdL8CZYW48iI/+/utbmYIKQq1kK7
NCPyNveIS3rOR4HE3nzlQrv/MEjPx16h6lDsSyFIa7wOt7tpNyLCX0yGQpKWE3jX
vQIbrfabSmIJo/h3s69+XebOEzhPutSnTPonnrCLKELWhmPdICALUxNDBWz1O0++
2jo1jvFdUfaDzz1FpiKp+OaKaar7DRLz8HJFQUaOcFcytWxJCiPytIDw17XmDiDy
TjHWPP/eHPDK6TRPxrRYKgXRbSponDEfU47Iszg3x+fDa7YWOHu5CXaaZbLePD5Q
9GRzQP0goBJs9h2W45l++bKfEl81Kr9JMP9HF5ibc6ir/kdH+HFVXjan+G6ZxdU8
Bl5lw63eODC7fz4IOnoD5ixMRXXuHmn1yUogBXbnoTSe0/kmgfcnBwHD8WJrz0/M
YtX53J1RfLi+x0wIW/IkxrVbIsUtjxReetsQZrAQogw6PMQNrYitcXd5XwN3p91B
+Ao9SHCx1EemZcEBIiz5TCxOjA2aJT276Bzl6BBvtkdDhXbAX2jJ0IYfimCk6t61
PSkJThQRw6xdMJIXrt30IdYAcNaOu9kHUqpeT8omVjOpkYdkpa9hwg1TsI5x+Jom
ZYAvkAwsyFV3cl4kbeT/0SAtkHPoJZ5X5PPW8XQP4x8=
`protect END_PROTECTED
