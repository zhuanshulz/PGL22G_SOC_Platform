`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RC5xBKmkN1zSyCX+n6ru6A5AV/D1ESJlme6y67KLy8z+5tXg7zKfacJiagLdhcWg
CaJ9Q0gbqBGr0/Z2qBvVHNMOGvBGmZ3d+VSFnljjS+TNyTFCyHWqQasioIkCLOg2
P6Db07Nx62Jdrqbpq5oyjAfOd5NYMSA2j+FoDRPsGGAHydLVH3Nmd+Gv6mDXxnpZ
N7Kku7SGMbuX/Wt/5o4PMscgFltoTKQGs/peSvYsnwjYcuZrqJfNOLPeoi8N0EWt
5W/nRvehmXkPIeglYmb0vjAuvpb7ZpKjPTEzd3/0UU0pjWdc/ExIujKsivEVrUQy
ypx+PSfiLRQpdDt4VtgY/K6aOKCrEFnL0iyOU5boK2lgdcTlZiwWvddISo9dgKXb
PeR8KYJFti/1pmjrAMykcgo3d+i0Pq89ZDvxCxaq24l9BUnxGNcLXdomVrYjNWEJ
3XBTCSb5uVpd2hqzeE8wfhgvKuqYT+XsGPT4nF5d7JQp/bc4N4IRM2chfHBSmV9c
0l6n/WYwGlKDTdDrHpSc/JQUZHwUCGv6qcK+9gGATzfovXiVkce0bWAA/IXXSzNX
ikD0Qdbj7Du3amklr+ZUnRDBk19afiRP15BMXRd0zMlLw6kEHvHjg040BnicXGb2
onX5b+NGyjfGs7wsaWjr56/UhjgUkh3F+owekzjTmgltaVeAmO7IOHTf/V36ERMf
6FtUUUhHdSTgWsxACg2L5vMZgRByYD5A8SVm1vvxkbhy9Dui+FZ3eRGK5xocKmq9
QmORnyFldmNhCtN7cM6/lw==
`protect END_PROTECTED
