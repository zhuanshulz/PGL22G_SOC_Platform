`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/A+5W6w3k34oymDnXZuuKOItmafpp9ZeuMN+h/9sP1q10u8s82liXDAMCsV9/zCi
/5R16drb5qlSopZupMfVEsPAOgodSt8F4BzognPRBjXi2q8Ufds/sxTne/7HuYuO
/i70Zh4FoI6DOXQAgmGwpt8rvTy23WmNQjiI3Gl69RYJcg0XduA05Lwgr7Fpi5t1
fj2/lnRj1VaooekQPZBYxIyhe7cVHG2Ym2IkVsR0JybY0fVbvHA6+EebrPryuqZ7
MCZohbEX56RjoPcTSTpst1HKxSlzKrpk0caeAKSU+we5LBd6pXFRWj9RrPQAlSbe
3nN3bL+PrEQJbOpPc2Rc4DRfOjYFt+XK1h1I9a8Erp2DoBRrbZ8yFPdDT7NHacAM
sRCr0c1ypx/oI0Eaek2w+ntjAyNcqNiK9+Qg8Lddv5tSZ2yPVsAwMIvNp+ansv0t
QOvInNJSPILP1KNzX95NlSnvYDyjTi6opi64hCShhqPUZhCrUQ2QStBR3ycTVh9W
+p1STqU34ooRWX7bFxWhhI7b0KVYrovU8N0GHznf9fGmzAY5AMQsg8nKDpErWjTX
ipx1pT6kHA/NBsp/IWtsx20JVUoO4A83TnevZpr0jr/HIliEFb0IxEG7UY+Zwham
Tm2ptj8AqpyUwgeIDJ1hBZ9Fy7RM6FHsxCYF4mqRkhQ3DmrH+kpA0tW6Y5SilXvB
PWpsolDF5xCPXZzUofdIFQiTBtRgKrZFqxODp/CoeYK0Uu9806PWV3hjibpIx7Ez
EWY2r7/gxUssmH5l6LamWWi0sKfSm/8oEavuNTE19dkl/r4NKq+C4UALW4p0y8YA
QHzv5BqcE3S7G59qpdGHuzCoXtuGWGN8mMAcm7rvyrpmkmofzJOGMzbiuHnGVNr6
QwdQpVfCiqGUAO9y2cD5a0qj7ALjidOa5Gjm/qKqETuPpMLMUgav5zEaXmkyuUBW
quTxsdV19EWewDxL8S2iZy/tiG1/zmZEEFaJqJBWrbeMI61oh44j+Mx0DhMf5YLP
q0jaEiBUt4MLsxLolehaziYoDZNhJ4b/cCkNuNj2eaINxTL9zURbE65kgV2SH4G0
kQn8611vGgtFtvq7M1miBRd2I/MNstnihmf3yRd2tb+b20sOOjycfYd6QJmJu0u2
RqGyLYiWxZrM0+A0uzNHvmKUK9lK+bIKRLV8ArogSbVZ/gVSusa6/G13Xho0gGxi
6KTBJacYROskXTlixGnQJebRwufc4b4/5/TZhJFN+W8u42np5akbvMa58AoXw7sn
yurtXkHSEW6iZ9is093Ha66S+1opHjIHaLyfNjvNX1O7HiJC1ZQRabRSy0WXZfJC
nMrnXd5uDPJer6AKVcts+++xQaBgciIEAyfEnuIujoiieVa8LdEsuJc4ibfhY85h
UL5R+VpdS8ZQ7aL9TTIsODbciuXLquFwvikkbM9jyOxurrFYPYL19qgCKjxjCSsj
qSybUDyQelnLZkU0bbukgIJAmplvaeYjoaX3vuZ5dD2FhQfonLYgfsZYjNFjX4jb
fAYpMr6sDgIlBDNlncfbJbqDFOWQhS18YEWdQq8mqnR9f0yFnT/C7oaSatRAxbrr
ijRkfdR/TYb5M1TB+Hs2oy6N5p08CffwWdmqWhbpZwYseJlwj8kTzz8ph/3zzz/u
OejOjZHB9+H6BvZfZgpwvOZB17rBF2TwYdcTKQH/11+9YlVYOUSX9a5IRLIJjt5f
EUr645XGWAVwd5RU2KKdv5Iyo4NCA1VYEvtNjY3ja3wO5PpfFjYiCPK9IYseCSMi
s3rPP2fHhNcEevsTLZMfh5wpgRA7Z5CDehTDRSdEpqs0FWV+nNTIDW8G5gX0GhN1
1fbO89Q2Gas3haHMIiDmTvJPMW3gL1S7Ui6b9qax8Wg//pJQfqjVD6kE0p5P1AL2
X5h+ce5pZnxYNPx/+50YEzlAKBkZcOxfzWe8LW2HuJ0GrL33/Jaq/3RNtVlWmrDW
mVcEsXYQXKHoiDmr9lTvKBw9gdMPKI455QcH/yJtueaeeH+jsnA0BMpFhl7SIXwH
9o/YtJKeoFpySeOpak9nDWJ0yo0PSvFWOPWS4DWARtes2qXQtHvt+MCBqFcNIUZ4
iXWWqiiJLzGIiweUs3q8wua/mFJYSNfaWt4vx54tDFBtizARKaCTlJtA3cjGs7Tp
hqf0W0WXWwuIF3namVB6YBkh5/gmTwOxse7FH6Sb0EHb33kQzEN7iRopSIRM9B0a
Jf1ds38ZJ2cv+vH0gQ3lmGcLBjS0SiylpfCDonQ6jqQHfYHSyALnL0r/M3Uk5297
jKG0UJhikcoijgzSE/bCQD4HPXFq2RuUNFYC7jNqLJJ0oPUVXpPjG8GgehDYsJ3p
9HuxQj/biWIt+9daUzfcOBUKY349p5v3jjBOvIcl7uoLkn0R+izo0Y3pQxFK34NO
DjRxhvucjOE2f41c+xWo7XrL3b3L+tUUV74v10T8Fk/h4rLUQsARBzJH8owwp3zb
sKf6UJYOuHQ1afOpffxXFaOJBkU25sson1lj2OfawOo7PyMZrFTVrK/Npn8Ax4xY
60d9tgAx9BaaVvvVOUksPIM8J/aGl6K199MolwgikFA7k/qfx3IzvjweuMwSlc4n
pRvGRuMSI6zu7Sa7p68QnCDqhU7WEe1lj2JCtfFW0WwwunprHeIrYgx5ZNrIVwqY
lXf2Cn7aM/gUVsC+MmC2syPQ6/2GMKX89MqwGLbYJwDHsuInqI2D1X1e2k1SCtD3
wH4ft7ZrlhelixH6aNq4Bc5PPygidK1aomM6TSmNRouySTjFLT1Sr7il9fVcsh5g
W6PY5dk/X2b2h+OuYhBZ4NCRm73fjc13yhkks59ViCaiXIiNRP6sUZ44fKlSqVPl
pimBSwgpKl1vjoMANldRnyE942VpEfxGt5ku4CyYA+WOS++i4RRR0oJgOnS2P5YG
kYk/ENhQZEY9QdXYzc0rVlYroMD5lpjuP7Joc/N8euGX1g1jiCE3QhdLMSik40hQ
T74aJ+SEwmycLnO+30kQBd0y+hxo+wirtRpBA3FU4uch4st5xC94fyTfmkr37erB
R/B91uMuNUb1kLHiJ3I2Y4eUfreod/ogbcmnaHqvZ2xrNMprmvto/PeUDw/IF3QY
VkPJM5A9q5mbqNWOa3AFxVZZgZahkhITGYyQB3ewr4+FN84V2FzjC485nYg53t26
6nGpWJbjUX1SExx4wPuxRGIs6k1YBORgJUaR9uAq86P46PKdj4Vo2bu+KBViOjq9
oxByPp1hwVrEVVE1PFLQvlAfQi7phDawau0GkT/mUcYjxZVicxzn66p44TP2xH+4
8xR/oiWuXMepuSuBSGwUF4VJOxFqyyA3asgUS3qpf0pJlPrUEw6wO9IzRHkM/8Oz
nuYdC9DHpqAKoqlxnepyYlVV+8rPDDYaiE83IU3Bec/at0fe7cogpGMNYEzSS2aV
v+/hqrvFyMs47XVA2ZfttMQuD8DU4yngXENIvWxPQ1r6maDPbGi1xD4S5D+59aKe
BkT9Lz3+00gsFToe9ajY9f+FSbDi+qE0LUxJsHVHfjRHVL8m7D9Lnuc99h4vf14H
DeD42Zsr4wrrxK4PyNcBLLYKxujVdqoaezyNck78aEuGi1ERZ6fX1mdQHKfPEgpv
VFHemTkf5oOZ4jjp7/aOg+Cvb1+peLsDaRkeV/aSHVL31Am6HtRPVWxl3LOZ31aN
2rLUxfh4jyCfl9IXqndXkw2HHY1jgo+3N+4UpnCTR+VorLpbksrInW6hGZ4RBi7o
OfLwKECPHSDdvDbVuUkHZzidr5wyejoyG14FaWaXaDtwvm7tojENhpJEeUrVkGD1
hfZMgkbnFU/VKYrQwd7mV4KXg73Nr3G43o8iOA5Ekxuzqiw75yzjU5goY0aUWQU4
ZPbyZTAbmfVQHawBgK9ZeuVLETx2NX2M715IvWvtCBk3RRlRbiLIYpINgUnF4akE
Cv1d3wD9tzLvMlmUxnyV3uFRyUbTJ4/56rX1q/EPn4InBxfVvypuwbcrWB4UHOx8
4rEuKS9IPGs+PBXe7F5sbCMo58NNhHqRLkIqAVQ2H5LXBrL2DWXn6xb6zorr5L/y
FMy5r+SCXVkcXMtjYQsMJgKPgLmLGaNFrvMx1gnK8O3Sv4nwPMlm1BoJm+Ld3wVn
pTuNfAhSsih/mLud4mluaGVLa1xgUfma+oXdWHnwyF2xnn1XmJll/o5t9gFHxFn1
UiGNqKeZzoaA1nYx4t1IwSdebSeP7RDKKDLt3xOcmAIAEXE8IaLWcU4/5bQUIpBf
ioRBk3oeh+63RsCEqRpKrDrGOF+QoFeEDQ3qcT4ir7wLmBwIeyhJoL4kt01fGQcI
XniG7Pj9YBU8cDwW2iJC9VdDv1ZsTmMCWkIv8faktu03o6V1GHrQHy8D4favREUK
vIeTWG7xskQGOObwkdw6UzXZCGfwzJkyqzBo6/SGS+5hLgzNxyjORQ9KjIKaFl2i
qga91lQvyWEFASZCR7YxljlyHM1D0z2BxEonaouAyk/DfHyBREvjW4bKo9mflmee
fw5mr4j0XbeFuxJCYLIIMtTM9df5qGc4EfIf3vrN3xcN99gPA6o5u5LaHEeGe039
FHTct8cyet7myst4qjaPyl4zJzpKzoBh/b/1aYqnKqaJShL8IPHY5drogkkFAkPa
medL64gHDmzVfS8ck4Cki3tfG+1iYSuK56UD7pTC9UdwGD/IocKW7m9ronxwbXHJ
xU0E4CDJhug5TZZ35+CNWOb8L8foqzycP3Thmij2LNkFp9dBAOEdf/Jpnvk4DTjK
scZmlN9w7ufJbWI+Wf/e+1ywL0GwYG1U1u4RsQ1WBF89+rGoHyHUF28BdELX+s04
KPxVtBobyDBRP0RyBMjBlKjZoX4sDvrxJHwJwZaGUVPxgr2/Ap3LJMcJ5HRnTLio
m0LL96LV1Bup2XhSruOgq00Zabp89FngP8FSQyWsvrDynrhWXYjHLzb2iL4wwNco
xZVgTyg/4kOT1vAWKwn1heW+9p5EYAH/oIApirJeXCHnW2iMPExtDXjoVh9wt99L
iZYJf7Aq8dv9m6iYm9Fg0uc/bEMONDmn/7WyUP4AkkV8R0h3BtWIwp3GyznBHTte
HMXC6zzmp+F4fg0Y/mWllBYlC0SAD9jBEzd8JlvYVFdpfrvFGzJN3NG3jh6F/Mfr
EFB+rjkkl3eQCGmELKpL5vQ+B0us3iS4rY0DdaI+CnXu5agns2SSYdlGYmHYln8n
pmT8tpU4D7ftFb4ns86i+Pl+8DBC4Hlfn466gBk2bHTw6oAHY+t45IMOAYQdHQD1
L/UfG5pwX6TD9T/CFSUjakWrc5vPOvCe4Geu9SYgWeYAvsijbw89SfLIbZLV9gK6
tJNimgpYMq0InQtk32aJYNRb/W9fvxdgE7V1iGY0ZOZoToZqn+RoOZUDqcZPGoLQ
U4iar0olKkn7fyLw1nwuU/mFFSP1D2dTWfHzr0su683zHv97O+WYrPYkhD9asnOL
lsWOiZlGPLBZth3RobAE3FXlXgirM0+rloZ8+110EYr8DiNOgBum6szab9gbNsvF
6KHYoF4GwDpbKoiMIkIZ9w7DHy+S9qUpnBnVxqe4UJ0PLjNqWBCVp5INqyxaiWNm
1lGTnF4Ejr4BZ0fbf6sMxnA0sk7njIx6UuRqDG8YwovUGEe4/WqVAlv5t/t10nx9
ljaZM2srnECm9j1VObJhY+e5MRfK4aXeM/paMeJ+oLqnM67V+K1zCBeoSefvCtuC
OGbIWNjj65mWsFq1AI0pAR8E8EOc2JY4/bhmvDL05chpLAHtR9hBoizfdRpKsOvi
w1aCxdt8oe1Xh65YE4JjYApisWWIhAZqDhy1Rkcr3GZYIlaBk3B6jCnv4O/bF24u
UMXMpZU5GDep3dB9YdPP7EIpz0vqciPmXgUex6mmtueViHMqpVsGpNQQJ4MM0ZZP
KysxtGgswNCCbayGffKErCKkpAiFnRXr1IOOeu2sCpktSBJxKB+dxxCev8zl9zOc
rFjfe0OWazFTTy8uepDGFQ6W3UmqE9z0tqI99pgKl6FQejYRHlUQJZk4Ivx4krfq
BXm4tRgTgvZijXHN0x74CHefDcrarhOO0VbCOFlL/irpq92jqTl4slqtcJF9di3H
wKWFwCIk/nY7JtADY5AadtlWx6LByEYAQbHj/Kx+l6pgQBht7VsVTcQuNqA2juNF
xXcy2G29LAnL12p4qdZRgNYMhlqxYqCft7435Q+tMx2jWzpVyp9zpb5iFT3Ag08a
bMX0o/MtmcgIePSEdj3Rr6MX8/6J0FoZMJBmo765WqvoMkbPH4GY52NsGy9HR6wG
2CMIpNTzkiyws7P9j+pDIIYKxzZ9ZYSuXAH+wdI5V7CjLnvlCwFeb+dbATLRSz2F
hVcW2kLRVnMZGgwH5uujCICbrmLqDfZr1tB/cy9lFRg7zNpTFYhm7Z4EEHbF1aSR
9X/V5+HoR0pcGc036giQmqnaNdOrtPlYfUOtspBFqFJskKWgTZNZQ6llalCAlD3x
wSBGHe9HmKJEFHyWMrHu1eO8nuENVBgJh8s1bKqBcLgT3esC1DYSeeaLWzWAw8Hh
1EfoN5oCQMYFQXYNX+LASbjEHIElvTxQM/8AMtC6wssi7SpbEaF/lHyR8/9YX2Ez
IKCEsFMPBXnBwlfa7ZEVTlvBa3lP+xS8JbwF+OcGPMtSGdLB1Czp1E5gP2rnFr2p
sqVDTIZRllzFKnj5EnMVMpl2Rm9DR/ifo2sAEhHoI5Ko8jDcOyZ5AA5cKhohFQOi
0Vk+lDZ1ImsssKKhxBOAo3qxgSrFHtvfK9h/Dyjrkqv+UoPrtWsrkISkGaJa9qVC
31X4mPCkuacuC9PKGxT3yKcIcmUezWsn18ilEjA1tiEqwGpdIlKzn+oUwikRBo8K
Lo90uSHJ5zHOMy1jmwlQ7/pEDQgoZE5/NLFpEqt8VY6xROK2plN9+e7fzPZr1kso
9hEjygwGkFmeeTvfkNT0Wb3IHKGwa55ss+IjvhWMCgXeoWRkLQyCRIZoiT3k9nne
NrrDjXvmSLlpilHsBPOI6E1Dtk+k9cgdo2WQ9B6dUE9SGFAAfmqnEjGFS+1Kh5ih
a27oYfgg7KtNhJJsenMUQDIQ05y5RHb0F5Sczwilad82lOALMOakF6oxq5xKLOir
vMMBz8sMMghCDmCvjdmZdiKTlwxFXpFdLlc2qcVHG/YIpcnVN0FeQ+YLEvsHj7+t
E69Oswt0/KwU0CLk7ekvw8RmJBTTxVMeBe4vzTZqQzAjvUKqarvjN2OC5cqvrxNu
JNK976j56vGk9LDqjpWYRhbpTnL3md2vjCEuLkZaGCTc52ev+RDHwaYookcYUJwF
d2L06sKE39UR6e5D0G4Rr19bZkrRC1X2RMXlHVcGSaxeQiy6F6cuheqwPsiNlIjP
t2aNaAEuv8SBtrJ4s1nppA9QcoXIyL4FGDMxAjA87WZR2Wvlh3DnR8BTTT0m9W48
gIKo0RXJ19k6AaXJ1RsF50fYY6wv3+6CcPCE162RnUC3YSxoOuLiNIIeJ9p8uiiZ
KG3U4VKzVNcUfjLJOCtIWM6e4jJzWjPYf9bkKhUe/vhpR2DrcXpc1h6f+jN09XdH
nQsw1B9ma2DEfzx6656ApRZcPE1E0R1i/z5Zb1/AwJg5QrGCoHy2u4cU0b+LxBjt
mHoVlYM0TvjkaPBValPfK+HKcTB0zlyqm7CVDP400g7m2KeE5Rvf72nOXO+kxDnF
mArHsiTx4rRsrA9VrHamExzjavZYMlPglUKFTdGZ/1VplNvzMT8c6EfrKSbcWgHi
Kd8WCFmx98Vp1IQ3Ev76lJwtuEF663LUWmRG9THbxU05BKqXNv0lH4DmOmlAhH9z
qMdqwfPAqS981d36Gng926rVGXmmL5zn2tduSkK16mYmVNFwiGGqnTG/GSGCSKtF
pRmP27/rkHvN8CvqyKKfUFjhhhJseXR3SPj5wefzlehqM7vITRK7hjgMNoSQqHeY
g9KCIQNf5/gphm8Tq7oRnVahJJ5+I31b60EYv7yNrejynRK1/dO+uxMqk+EKdnvA
KYiNf0VVnlV5tcW5ylKkcDCyrcbxtrvaojTC0ftt2oMHQ+h30jd5m/5mFq3ghyLG
Hqf7xwu2Ju94oW0LGjMlr9YvuT4I7J9WRo8U5BAIHKZd6ojBDY+OrB+yi2UAy/bL
8w6gtq00wPGuDHtPITW/IFLSo1VxYJMzB89OaDtFrLXh0Yx0mIKY0iiBu+NR6Tyh
Ebf2BgDb/kLM3rV/tMhTNNJKleIfdh5/B/uSgs43jOnDJTvc3eaGt+Vl2L6zTfbz
4u2Izmk6U2ySR7oN0l3wNRlkpyLBZ2LI9h76exgoYWwBYyy7OjvVr8YK72bInmKW
iCVxOZDkGbFZanWxleP9rTXdbhugkiJA9g3O0SZNEUJztkdTVSV8v2cdb2v8W22s
iJcyubsfu+DnTd9YwfLfCcG6isa+16yElOe0UiNaFwy2ecIIhRBxTVmZqFzXh8eX
+0Pp63BoVKMcpIQkPuG3n8GZpJtFOso5nEqmwwX7Vzbn8QEan1jMpi68ww4DHWlq
mwzjX+C9/yNnscICU4qkNdvZnAapml70qFd616SiWkLbql63+vn9I8n5rOzJZUYc
csGkLykjelaCjA27b/lhsbivk5sQJ6RB9EMRcHGzqkdLuojQ7CUETVm6OTwIxUrI
ZaEy7D4wTyZOlqtEtmToyH7bZeVLbJxIsSTDf8HyVrYUyObGVtcYOqO2IeFCI2o6
uppEHGzeojZ6jJIs0n0p5cxK8W6oP7ESzQhkc0c8CC3wcHR0ZXCeZo/JK4B3srvG
TFTleuv/3ITMg9Avj3kA4PRYLBcL7h7c8/yQNJA24ucTkRTO1FP+OXkirDQKzb3W
bQx8AwsA/kQqxFVX3VLMFXINGSYnJvYjazZnhQUGcYB2EeNP0RCW1buu1r8rnmR4
fOnkMnIwoZDwCdcOL9DTA+GhLASXYRSBu9Aa5scwh/7/Cf6XwCgsd2VIeJG1z+yk
aXtj098NaHuDiBxcAJAap6FIAVJKqngmIf9XD5rSzmPT5oZrOzYWh/F5QU65EeI3
4IXhuFofG6oswfWRX9Oq8HS3O2d9/anXcby3ZxM+qofOmd1JXa4wYbNglFXfMnXf
sIU8J4pkqhblwUGKsQOzMumrUQPvTKjd1TtL2bndHB3uGNZCNX21Is9rfcr/Fp1C
EdurpYtH/RHQKGUc++OTyPWvpteJvgv96uhezd/Y4ze8hcTxYKkdAiotTjGPKR66
0Qm+dqsY2u8HUPlHsSFhyEoBgfvRCRoWht0axpuF+xs=
`protect END_PROTECTED
