`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sVSUM/KcIxr6js5YVpxV3mqCzI8hYxygawo2ld1K/EBK5WMNUYbzNrZXe1WtQhpO
e+zpaT9/MVQ1dphZoJND2027kueBxPbjQQO5E7Y7HOvV6ejjfpd2N0wG/PyeppMq
ttU0hu5eThL4snsP9OiOvb0F+K+Z+o0QE0yV8VFjxk3GD+tFQlsUZ9YXmld2N6G7
9vseZo+BLWrdDWxkiXCKHa7ZS30cglpTH3vdk8eXqtg1N7X20cbYQgVGJmAKgtCF
u8BLH4hM6vR749tvk7oqMZSOzPIfifSxRqLOyZ7NcoXbrqpu6HztXDuHElFGK1Eo
zzzSANs+CR/OHgzvhBBZjZz/gAnrUvmXBs4pf3t1f2+naRLXuN5r0k0cQ3x5pVYb
rXa4lAx3uSSgrAxnWldjX43l+DuWxzlJ5Ce4AZHF0G/YpoYUQZ2e0V9C37IqspTw
ZG8bxpRBglmowcP+UPgMvCgJbYfUplRRq6ZMrY6+tp3Qk+pSmqsIqqQjxl02SY7T
IRTNoKiKrBYZL+WgUUj1nhj7GRaSmevyOrS/ppliA54QaPfkbFaOwMk9rIMoCfIW
/nBQqb8sxy2LcQIHDbHTSQonxnNDlMjHULIq32e2HPFdFQV8mBPk830fRMknb0J8
3IYWo9uKoWj4qKTNYJCQP4pRgqE3bYsMPjEVk0GOQ8MXh89B1GnaFUs4BoCMyXoE
0ECDPlqih3AYYfw8fFWHuJjIRuPbIf/Aiipi376GAL3ZmXGDwDMrEk3QfED9G8kp
jwUD6BUOWB2ukfv/mMXW1nPiVK5+0eSOWUhnx9V9VB/bHr4kdQjo+l/Z6nRk18Gk
VGxT83qE6KXwMHm2H8ZNRfypV/VoCFAo06ntJlCRmeI4azqfy+rxNA25labM2jO6
rneDblEQDXm1EjM2EP9itCDCsTT7GX5vU94KfVzemh7yTkInggoHKCI6jVhLznRs
WiuJtoBSEX4XgpBzDbulGDkBDv+AS2gvQv8dl8Hb2oFjlA5sybofjB5Whi/Oo7rF
oxG+KKWrpN31yeRoB7hRusqp7dqnI3B1WrL9ZTDBPCbE1c5peZPcnCfgBZDKypIC
y0UUKhv656jOam5C74B6UQM5wcv1LyAcPV3y16GgShSUD8KNoEMUCabl+61nj+FR
GNgd+I32FR6LDUjG0c0KFlPdj3Ct1r3JRjlPU898ZFMSmKSQ5sjgPVtTNsFGYhxM
1uQVo+HNcLJna7FDzalTY1JA15XcBnXKwTuTJsibN58A8gEefNI9QvRm4wwjTRTg
TZoAtGCrpNw53sUpcjaUIlzTRwkIQHwfspJk8Bzx2h0faxqzVJZMigEC2TnjF5zI
Ezx6dCWUiiz65Lpe07GKUGlBzSIKQpKYYxNEBVa1ZTr0nPJjv3vAGsPIFaRDENMi
lMczpilKnhx7ZK/6Fq0Yq8nvRHKS5gqP8p3q40iKWTL+jd/CFKPZ+B3bCbVA5BpF
O7C6uFvpAPtJWJvURjvxev33wrka+o3qzVA5DD1Z1VV1m8EjLgG9oqKZjyhiLyNA
pnVqY3Ta2+/ZBLrBljw58RZVJmdBr4J+3se4XUISimklk5/xJuDuHDSW+UDxvhIB
xnkcX1cLEZcE/RvUqG1F3qLJVIhvJZMFXQZo6no5VaqcxnBkBKZow01EwB2h4h0B
/bB0+Rf7tFzdXIGuBRSlLLwj91BEDhT6m9SMDG68x+Z8qWEu4jtJn3tbcswDySxF
jzBBaCPuArUPfSCa+EL0hP86x3k4Qur8ZarAj7EjC2NQdBFX//4TMtC1sKb5hnLL
Y+IFhRhy3BxKHkmoFqTsRUhtptWX+wCP41iVKJCo01RpnYH0HkafXrvTcqAkO4Hx
iovxMC7M276/hgwrTUWFNKxSjimhS+G/dLZRrjfjQ+6mCJnj2kzHvM4zsZqTxhNy
cPZnWEhuDNhir1YEwfuT+QcX99UT3TJ1HaRIvJDu5B6wQ+Igc6kKTFW+i/yBPyem
5mCyommA2W54Dh6AUy6Wi7r3iGDHh14qy9fR2opA17tzIJX6dLfuGzkgaQAiP24o
bqkVQoRR7ZgwQL/g+rPxtmrv5yowJDspLMTOprXqAoLrj4F4s+DXlxzm9t5lyqY9
XElUuDRP/096RFK4RdetvrV/p9Wy865Ot71nDU++7iaDTtA/kjhvezVGv55X7K+c
wK7eitByZ/Sb3gn1xLg2YcGj9OuITaZJf67JqOmGtjnpe76XM3MNJ/UMpbtsuUNu
3ZuH1ECHzbGwjljtd1Lqb2Rqjrn957nPYH7Y/++CE+UWQkBnPt1qPV1fdYY5/xjQ
gbZtsFm6XMcKakbINAKg0k05tioeHes/yZFPC47IkB8My97LBt80mRIrMbzHgywX
v8LQ3gGbTiXdxpXlBo2SOQl+889xuPY9TvEZ9Gmlvh9Jd9Z8hmSVw2Zw8kK7Umi2
envDtPakc6/tNePvsyvzr28Imyzuzy1hNUVFNUvOO0xWa0UAZtdfmdnv/nTIxVDi
xdFajrd/7DiNqYGnZ8n/hAcpqfDD85S6o4ahcFP3dJorJgG0WaNEyvKHB/62XQNF
S8KbzBCcOVp4WZuQJqfOvovjTcNp5oaLr4GG8UVpKKY6s1JJRDI8/9Ozqiwhleoj
VZVQoqr/afsd6/uj7cd0QL8UT+43cUokegAKnkf3O0ZV9JIZiwV3u9SJpqjxsYux
QGWW09PznenwPcdoF8wz7UXQIfyrhwryHF5ZrKPrbW5dU9Cp+FgB6k6DqwI9eQaE
I4jNSf6DUGgLVz4TLU3XYLHbwK9YUjAHPhnAPnwTV1LkGx5+Q0RVMonuYOaN9dB6
gkzFt9mCZVUgkhbeAmMl9WIV35Nl1XToUpVP3CdZistUBf7idyT0QmR79SgKaA4X
mMMi8cUGu+gOF6zx0nvVqG3KqYW5Nd4sJrg64k68i6gILQSF6ynMhOmEi8/Eq/oM
3kk/ML+zhxe8Y3S+wZ1KBuFuXG72afm+dRPFMfeJYjF0MlESzMEW1qc7vvyUpunK
Mf7OANdw7yjxbyoUYwrB7GH4nMn51cCD1Nsx/19tdtERI2umSvvmAUvP3Wx/7fkH
hQMEoZo65Zd2j6XtyCO4l1grYTuXe9dBNh5sofULq5flhGtGlOxEf+AHMEx3nRkq
yvltoFY7ciwBoLxqy5aWhfQ1fr004P6C/bk51/RAfEdPFMR3bQ7XfBQKoH7fJqjS
fNef5UhKqYkTsx/nTxl7jUIbj41exO2zpRGn6KMsnVc/NpW45sKBKblEEHhboadK
Obu+69rZg2OXGMZic3bxyEGs1T3eSrsHNhcK4Omid7AeoN3VAZaqf3augvnMfTAh
ynY9qvFAdcv4nkC9Z3E+jorrzku7d0mzQUIHRoXxkdy7rVkFNxChWpOhCJnibRCG
WkheAvf8/mOOcjZv06GAOTA37LgbOxf89v8/EbhurtczPBZJ4vq02Ew+4j2tY7KH
Op7RwnR8PeNX8n0oGTSJ1aWdCwJWgqBew7K1UAlBJuZptUSjtCfAVH0EtA6IYqVy
IzvHdQIkX36Tnk4w9VTBsyF9kN4beRcR5HdPjEldyaIvt0GyQBehHwOPugvDrFkU
uTJ/06Wx16qy4NBMKOdEGUpR4gnksOrchx2w5X00yenB0py2baIdu8GPytMLpSdC
thhgpFdPepBBBBHpJoIEyxAE3iyj/6As1F+AP6fkvQy9KGXAkXzoZ4IXQi10zRly
foda9UxDnutOFRFnJ07PeUJQAz+4/YzuPbMnwNqaY9JRBHD8/HohRhBAhnwAFffT
p36aEHsGiBIwEtq+HYD4LILjEiCp5Zb8dn5hqxahH3GI6IJrQHlK3VsDv+7O4Dvk
QafAmsnDrUMN+233N0cfR3PKE3681sUEP9xjvfRvJJx2twipVrMQ8oJzesQwGVPP
fF17SS+csJwd8CDOExd2NSdB8lGHkM1k/ZHoutBFywYZhjOKfKcEf3jVrhmhcVlK
oBUhX6hwLh0WeQRj7TUiDjyXa7YpJaZOKOWZ4NacFdgZ6w39AlTvGZZCtYd/jJRy
m9cTRgAmX76P9LSFbI2MyOt3z9oYc7YuNdaNVywQk3bNKoM3O9QJDCOrKvuFdSRk
JoFw3/fz7EujaJRRgkQOu1rmICqp6vfu621/zkEJo0oltDPwek/beEUkP2Gg+S0B
hYkQ0eHgf/VpujHvXED65K+dKmLJHjhSw3dLVgDOB8eowzJ2I2fXMf9XD8dI3BZv
mTL9Yke4uX4aDwvwgjPSRwrwk5VcOzR4734C/C4aMNIBwtTdoonlF8ICzAhkzY/A
rbNfVwRQ+fcFLVi7HCoH1Fua5jMZ/Xo91zpY2tppUHqwIKKOSyIHek4YEf+BDtR7
SSOS4SE8T0xyhuzVtGbIA6IiZGPo+sUk6Sb59aIuaIPSRpKMDWSAfqLSFHIkZRo4
4BmdCN4SXvVcCm6A9TWb3jYtBW/BxIoepaNbbS58YZmM1JSAGpQdySwEy5auGUTs
swEtohOCVpIR8X0XLXBEdHaEtiB1MkydlbnPGasiKK/Q3PJbxLDZ7BHWttAPjyAp
kksUmW7gag17RV07o9F0avsweTvS83REOEHE5QrXCLHATlollQ80XBYQHR2K0Kq0
z/OctkzYZ5XLa/jo2en6tD6iStzJydbl3kEB3tqRUZ6EnkQhlCCYng6g6kQBLiBq
kH+4+j0xhGKCNNh0pjqVZPOfzYmApnRAUhSGHYVdPdQPkeuAoGvatNRb2SHb1YSj
GxFMrlkA/R98VCRapdVr7/kf4gvKplPq6oozzTDgs6JPGiUOdYIQTPX20LAwdm7j
RWxF4IHYseMwyHqNw53aSKX7LYzj/+0kSsxAxE2BjkPCofM3VGLD3EE4IuYRKGnR
xtaeZhSIpMHDzOeVRqapmDJAjElyuLQz4NhdnrjwxrLRckfmDfC2uioIJBTPbagf
gi58t7mYgqdwDg2NTprNgAoeTkxfReBY/OZMdwQSAUOYc+VbKeAN71WXIElM+sDi
yCWnp8JscbEqHfDtB5CkPgzEes1G6rto3bx7SqboDdzEH49VkSvP1NFLrMBwN/Pv
f6Q73M/2HNUSgdmq0yFlUx7OjlYHgknyG75BCM0LzMfERyhx/G4zSj7OwNx9vj99
QCYYE9J2mTjuj+Pldn9DSJRuljpDd9eRCZ5zlEoyCo+rnswhqUKOo+Yl50syg5zQ
z0Ri3Wm724WLWAi5ocSf6++sQ3GbISoRNlJNq4DPEKdABTFy2tznfrNsi7BIuvNp
082fMqtEoROk9S39sQSZ12Cnwtflj/j0sfXpJufPmObETUn3w+ARy1LKvRfmCerb
A6SqiP+T0E0GvB7LFLIbDQ3iJwm2KCVDr/0Q1o1E2LLygmobrVMzUm/aVf8dggWA
X2rIvVAchL0aW5a1+icAhySq9GInaRpHvBq5jEH9m7F3dH+ABn+gaZnX/2WsI27/
nGYQj0ELKOMzb/hbTt4wFf+Pcf5qik1wj127+/1Rk9DKCXiStbu/NwfKByhGY/Fk
nbg33F4iCsHlqhiisqiCZTJHOhnDIlAN8L5itA8dHNqc3QLOpyzi3ZfyXc3gzqGx
Bbc7ySnI57c1ciwVjoV5Stl5X0K135+EvjjsaKmQbOAlLNHVPuJxG7MyO7F++oXE
yoLDtU9ImMFRXZBMOkjYq1w+0Sm02LOQdl51nxq+qziezXqTbLku54ibWnZ6THiX
u26EtGO8p4TIZcLzvkasPA==
`protect END_PROTECTED
