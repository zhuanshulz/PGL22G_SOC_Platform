`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5cmeEuM2wXQk7vyRiwD4dQ4uND9SB/c/1rATU2koIqn2xcOmoQkHatzVs40xd0aQ
UZGsqgqIpn8QMZ/k5GcJ3xR6tqPpdDgZM1FKdVSGPdlU48YoRg+BgPVq72IF/o/A
f6B+syawpCL89v/1b9K7WYzNn0d7VZCwyNScPGWn0Pd53k/PNS0IY1p8XbLLRHLv
ZMm8tPKJ7tdfwslDq05gZt/CakMEkhCZyKUAwAdIWgSK31sM93vtF1F2bWGYi4Fp
9UmNChhRFjLYriZe2WW3GNfWnAk19apAZJuOgiTbXjkYOZ/PA1kz7kf5Xe9dJyTs
RPo1C2Jk6BOGoW2j21EG05Rh7DZWGgXfn+3gOLH06kWfyf8R1CylW/FWxcVeryHn
eI5b7aOsZQWt7n/WXABTDtZnth4sJCA6DNa1I9VlucU=
`protect END_PROTECTED
