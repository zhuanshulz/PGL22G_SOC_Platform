`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sw8XEjSGDix+4grLo6fUp0dGwJBY9+ORptKjiiXjrIH0SdyHKauF86byTGAEELtB
Rl4SdZerjAM7FKwm/l+7ck5e2rJKvVsgNJeAEOyTmpSmalmU/7oJk2vBZbklOtOq
SWMqrxm6++NKIA0sdVQgtZgdxH5qi1oaP3axArL0wSM8T69jtI1GbK38eDSwPbXB
7/m4wQmcITvOKsOcOwyaQxy21aaCKRKU5kLuPwF5+CHdjjOFYeSDfhB8zCiZD1Vu
BikhLA6f4CVLHo5RJ47IIFxPF2hrKzlpfBiArlJ4LMSNEXh4kCh0AhQE7UtBiz61
mYOyIcuXUwpQLZAm5RkZxA==
`protect END_PROTECTED
