`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5348baq/9EE7fPCWkq/+zuJfO+RA+xmivcailpz3BctAH/hdPMMxBEBQNxC1Te2
/EcuHC1HRtYK43jEzHDU34rDGLmy+Df1miHdPhZZnV1iDGo05T2pbexuMXO9U1OS
LYJQ9w77GdWq4fiwwuUg6a/vBdkQ6HRw/dWL6+CK9rDz0FEElz1dz1ib85yGXIl8
9M+JcbyBCGwQ1oFyKmmqej/mWNJra0TWWkJKs7ju4mjsu6yD2lrDYKYHdCXjsgRm
vifvzbufv9+7/lDN5FrBzVhwQ6nQKr+aDz3ES6i6R4ftgxAKjJgD1cofHrela5TB
NvktgkAzEPkluStP8HU1wloDerAHd8e4BeUuQYQHnV+tTQeExugtguOM7di2GIf4
ld1PMDZMfV0RLnaC6/VwbvSb8Sn+h4kU3RpOjQEsCl5oK8vuATd0Q1+hBVGSvElz
Ccdf6KVtK7saixXpoFYhuCB6ODoizPU1Ldt2GDpQiwhLG2iBkfYdLAT5l0V624D/
tsWd7DPQix0qV9IV/H39MgRQDfAymMJmIjM273Aj6F5XyaPf1OLQODqTTt/pgp8D
0EKaeSQTWOkFQytB+bFEz1J5JI+zIi6Y0BnlEPawAqgPcJo3usYNZMbYZWPcB0Qg
FsgTa2nhhHNNMRBZusP7Us2D1u38GGYPcmm4Cu277VBYeccLpSnqTkJe/giLysiM
u5J7lKQFW+VwV7oJDSlluiWHBpOrgEvhzapj8AyhONA6MtABi1g0amW/piUyGl/o
l80mxccmjAlRqLVTQiLzx1MyVXUOWTYJ7ujf6oyKIoX71Pav9a0ak509mA4mesec
htA9vsqyvzEe014rjO/Btwo7cFkD/7WFGXb5pPDoYLKHZIGp8s68Pxdv8NCDy8Wd
kbbe0cBQ53/Iu9593G5OnlLCfINQofP366IipcWDehHVf3ArjnPEz6pfEse/XKC0
WztMirHUSse3F1G/vRK7swjHU6gawHpubaQNcILOLgoqaEohqqBWnLey7J9ciC1A
UQ5FrsVyExHbRzXzz16SM5s5WRQyNQmmI6jg+FqXTjr9JRJAxsgCJopLmLq3+HvX
0KJ92UKUn/xrFGJ3FZRNXVupQH03UKnTQbT9/KLJXZZv3sW+//l6p8JmVINKR6lv
KzrwOPXZ1j5MH4wWSSOgZtngdQnBulQDAGHChVDRPmuZAVNsjzhl0rXJlurSDJvb
ZJf9SSc8NlTGpIOyJD9vDoeeeYXijWFyB1XalKYpnUyzg6K4TZ23R4DmE2CuoQxm
1Thh3KJVu8j4pp58Kb6hpw==
`protect END_PROTECTED
