`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNZ3bxCKhrQp1llhr91s5vADJdcuVWlvQ99elb6EIPayrJJ+OARtxQyFCZUH2Awz
rlDD2msVflKWAVNJLnD8HBGzQJYioHC4+qOSvyzfcu+AUuudetcMeL+PTi6iQulO
FBHOlQay21T/FajxCXSojdTQ+sCukly40PutG4YKV6a1if48V+PuwNYnFlQZ2kVs
6EniebMiJO4g00I98wvVf+qJ1lOoOdyjYDlrqjYOl7n+3aIRw3D+HwxGfiSUyxbt
c8GORy7iSacooiAaggJErGoKy/fwbDN3qMDeoCaLIYUCm0xop+hBT+/P0f1NKTn9
GlUYIrn6Vz5JAa9PcY1zy0vtO7hgu9JOLiZSeAt7m5/7CJ1M7DSma76rl08YKLba
2sKtpi8qI4s1yNuqilQh7+ehhTB0XC4yiMvllOKbmnYMkG9kDJOa0p5pCExI1j+J
7+SypQ6izFq0AmRXTOfm/RBbsgv2z/2B9xkDNAe7m7Sh4tRjqB54HwsMYNOu5BgM
e597F+zo4nortbfCrobqf+HTCMw7TEf/e3DYMJK2Gvuom18/JWxFM5s4KFCR5aQY
Q4IM0lc9xUskUH5IGNy+ETn8rKztCLvsO15PI0I+MUO1L69IhWoyvQN5CsTiGQ29
0yHoq7LJHvyZ/MgWyri7BZ+M8ZXgBNevh4t6zgO26+7rXg7kA5WBy25KR0ueCUy5
PV4q2b2qHUNmkZ9npJPo4fwlVQU1VcxdTwGtgBLCGzWT3vkh7Iue6t6nyGYWzBz+
EcSDp0jU1BaeIOsHtbfct3YYJ25CYzD9WrTHHBd2W0FJCYcgbmGfwA10x6CVI1UQ
C4RttD06gkiGorTZBPLb2iUwhpVCFpmREPyf0Wic3Dw4srET/d8ycKB7Np0hLMGZ
TF4MyPG5h7/BcPDZbHorsoNbZagkspGJYivSIb7wFuJmO8TOA8vjMy/nFPnVDUo0
lVqXojOzdxGGIff15KnP9NqKFytBluz7uVZ8aWY0z3MEG18Donce7KFAKlCTpItn
Iwu92kLqob6uMKTJC/qd5kP6Y0r1xqZawphu1OKczehtG3Qivh7AnDJdv0ekpoQe
En4Y/iY6b6ZDcjrioqgN3XMLYkqpw/TXWNkvHGDX+MDKCpetD/f2oTYmpTXm83Oy
jeJX5lrDZonnuPP2Y9JYCX8Jnh5/OlgQ27JG03YNu9px0J7Uh+ZvXLD04liXiCJr
mG5ALCrE2RThAGs9FlfdqyKOx9YNyl6SRSxWHKasAe+mjo6WIN3Fd7vEMN0ZBxMx
flv7HhwTRmT2QpyL0rDbRZ1iSmGT0oyCg0whj9u+pQNyGgu2cMUtgFX2WC8ItydN
BGM1Smex/lhjv2QVa54D8MKNaIAzYTkiJmfXiLDXbeaybJhJamK8bnSnl+0t0Wzo
nBVfdK+5wMHs48lUWySjdytveFrneAtBzEONy9w4E/GhWfeV6FdZp+96VxbstTAJ
o843YZgXOYXSK9LHV7ycShYFg/IqPLqhl/wYVLCSb+wZS+eVNozKJAHXROQdem6e
E2iRK1dHbafqLsgFw0/PAwK/W0BuniXa4NCgiI6EXSAxhtNC5kMJPytPHPHGrcoc
dyhXdshEqeQ0V+oLf+cjMsdKYRfsdNhxJaqe2IrN4se0v4vltFDG+gPWGtwszcnX
fHHS+0vt6uWYstaxb0EBokmndbngiM+D6jtYN4FtcnVcYOjeoarOF0SmBFLqHvB7
QEwwCkFUxJl6+gohu+yGTJuRK9NU6zRLyMVnVObA9AK2Ion7mgT2jLGPQsD4IAOS
wcnnWq417WfVWMH3AFjBksPIs7a7AVzMQJy1I/naeMRDLMLeY90ysrxaHyy9o+//
1hxLbQsROpMJuoagPWjWf3e6eVteBaQ1QUBqfojLfAw7oySZPGw/lspMtg+jTDS8
pBvZPVcLPuIxDb30uNKu9aWjW19b46Umt5Ep/nV3oP02RQJicK8FV/uFkI9x0lIp
SRVyh4EXhcuM5tSxCV8PV7F7dJdcuow56p5A/DiMNlAAAHuU2Xmn2+Ice1OAYuEV
2LYP/Q2Dosm/z6VDjmErtXCg9+rA4z+LaJjq8F9JjrGKR5zYInXj0J0Ljek4iFla
MxxyBwFa6eiiIXefLfwVtpcRqJfvko62qRaT7ekhvQbGtq6M7lMLTSFOlsU9IFmh
mR3HJU5r7slN2/zSRMkVPPeH+gCHCelzarJZe12wicH2TuyWddtGx4f8h4j8/Lfe
Gg0H8Bpe09K64Ru7xNSktS14fIcGS+qScVjHYaHx48iBk2M4aIWZycftslNLoQqN
53V1QlY5u04ssTvaMiMAjRrMBWm/XVegPDJpUsADd15PICzDqbG8iNzzHduhCZn0
HXywNsW8vH+TkOqtr5P0eZRZwXqkuu/Q4eSzVDVcLomhqGnoMgFY7+IMg479rZ0X
NP25H8Fa/yTbptxrrhkRIwo+Lwb3ZR/5yqD1zBqWzQgHJVub1wkzurlRsx0sZJX4
oEZEfNoOtZxL4yaIYLjOJ1e/P+qT9NE6WNgMNHbYclrI2bC5UrGCpal4d75QsYm8
vIdzy0dzbuejojyRf3/+XuFHv90VBbQLP87auWQ9Spa3ymyRPaqYzEvWb+7phS7C
WRkun8sRV+OXtZfzjvNdpDZqNwr5ffsACJoDYByfV/TQNHfc+wKBG6FPTR2SAsJQ
91O8K1yjyyPFmS1Llr6D7uGOiEsf53xvDOJwV/dAyLkd4FuIre/7Jof9vmxaKthW
VGahgCau1QlUSr1xyLYNGA==
`protect END_PROTECTED
