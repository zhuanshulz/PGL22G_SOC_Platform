`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gGELz2Dy0TKslgDamI4XB+oqqVAWFH3sMxQgvq7e4eSTU3odIXtUT3Ifg6szn/jN
smZVTS3piOOlg4oln1+6VwXLYyuayY1ubJ+yhXb8e5i3o2jrZR3e/8/mIs1Jg2EE
HheuvUGdnehSMNoBE1CJ/3NVJuOaxCCpwzzX43Sy4mSxW673iQLWJmofPpK1SShy
iqV6BnlkbXEYmOC1STsXNBhzfdYRk5JKPgmZrevPyTalR4iaqvtJdBacVqpZrhJ4
cBSa6Yd5vDLUq4Nbl3S6g7wCFTPiCrOKspSfrSS0+MX70C9XcOKRzr3be3hzfgWS
CYk8YgYvLj9Amrw/YxaIpmbsvkbteS6aSNTpsODTcV0ofPcoIKnPy/XgQAcl5tEe
MDYJMZzhUQnsTmGGXBriNP3ZQxplFJRrTUsvQG1+w2P1vq8nFZb19losHDXvWR9Y
HBln69uiBVnBXtMJEWNSWbgWPaVcu3cBsdxv7p+D/vriUcGGdvKNFA+xpEc4Tg+k
enaOSulJAKinnzlSFKgp7u8KCDd5LFly3gkIIMexSfUkr1EbesIKpkuHl1QFDPDg
jXIuxpBy7gRoIbQGbrlZdZJT2FUPRAn+nQ6OFjluArcamOwHq2AutTC9RgQF4OTA
6TH63KYhn/movY0hohVBVUJOrsO6v7vvjKGpMxoMAn7qe4S6dSLEWuCNNJ13lJu6
jDuhEfuzIpIqZyoJmPCoalp6FTfYt6w8ZfELv5BTjEm39dUjEz8i7eylhA4HOazf
AyY36KwaySHAJyCCgskzNCzOUYZ9cZhxMX/9huXu96AiL3zzv6oTFiWC33SRnBC9
Q61lqbeq2pI+aF0W1dpClshofD2oapGiDwtmXDVXvXqkxJo9sA0cMWEsiNUKJ4Kl
k81DNPCL2AN85GAkVvgzBYPaAhrLD4SdPRjw2jbC2sCzp65/+kz4gEfm/XARplCM
MMYEMVtJy6RxuRYxQ+plGgVxZaKC13u5TcmzjjJaWQWwKT2CNoBPc2bOypeYiiRF
zy35I5wCEAwQ3bfCEcEv9XgCrvd+TyIxJz68p3oA21LaYkUIwoW4uhozT0qoJJIZ
AxQR/Aj9hLX+/6NTfaPHQFxjb9VCfH763pb2wTsYGxqBXQLpXrxpmANElnk+dhvE
`protect END_PROTECTED
