`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7vmDzHID30g2F9SvdRDiZ/NF2EKdcZV4aiGIDLXmdFIsC8i/GUZ1wIMJh2tAHTcI
9fvmB8sDgvDthV1g9r3/s6Rp6GB+0f+9Vzn1JTnBL/FKpT42FoQ0uYonoVxfOuHv
gaWh4U+HLpFWp/C5bd0qbyw71RNq5Zuvkl5MIr4dh5LGTJ9VklTThP67b2UDznqJ
g7AFAPhPkB+qTgZzizq53KinDGYu49AGwHzMpHVZ0hXT0QhMue4KzB/81d+Zh+7h
YQXsXp3iPQlMwunSDQhodW+mQra4kZ1Jn9os9QNEXz/CPerNHREGi8Es/H7aJggU
HSLZTnCXLEeOOJkqWp+a7wICeSKmD2LCLSUVMIh9NaQghv7axrhhpBhIGXi+kAxf
9CpurKQGvZjLd6BnmzdpcVqkT8f5GseD3roy8kWNci3MdDDXDg9UwnpOjEmmrvk2
TwwAcdNbNaWtLtx0Cng86RfUuynI8IJWINPURQodnTXl4JPRanHJlnZa2dWjiEUc
6VM0PV/2bN3A0svlBS6yRjSDzY4ZVXik+NoSxmts6JNzrUel/SoEmTCZIm4OQbTW
yjve+Ocz9xvK0mLxLmMNjKlQY4taIl4rxGO+v6xvdgCul0ZJrpbkUANszR152r9l
dSn1TCm2e79BWz41jbvtJaXe9ir6tY+sjZd6q/VjAadQMPKOrEQsIoJFao1tHRPf
+aD2pFh+UIyNUcUEuMWHfbJ9x5sfavgYRZRTgmTQ/3M7LN9piw+0Qqrm/KAPR5xF
XZTQE37SZzj1Vjo4Zw+n4JwEJ3zS4RmA/jskM7f9ST42mXbXX2vUouVCFESmkfho
q8mLnbKkxCVVq0sz09DokFjBb262bPyKUfYLyCAGWdo=
`protect END_PROTECTED
