`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uWYoHPfBAEAeJbne1IerENHdVuwe/4zq5CBUKbWf3dWBZL2Kq5wiTNYqz5KJie28
EIiqJ2czWMv0s6TPni8xM7u4sQyDlqYGsxgDOkvQwSmpRJzraFV688LZnXyir+Yw
MoiTwLkfvU4gj23H/+QXkrI4YpDbZdu+6L3Yse6JzoacmkBnd0MPqr3TL0qiaO7o
fIFsM/vgu6N9SW/RqTpppjZdep6ucxOqspZ8TdnJWZtCEvUCTNtnquV9m1djmU1q
RFCkBVjodWSNWr8yjkrntw1qj5+T0kKOX7topKkspJqqo66+axF2+7Ek9jgmbBxx
ydxspS1d00IBb1IpHbyIK8gs2zuZ4kHKaJVQ+f3qgca9ZKnoXTFJb+BeNYZeatoP
KA2wTUbCvbg/C4WC9pzxgjYfsljMVCyZq6dR82Z7op/QRQ1eZ9sQsXoGcFXOkP0h
lLdewPY86yg7opmOJpnrzJfEmWLSlkTbNudTVqhsPvLmYy73kxnm5j1+WVqf17Eb
so87aub28Cm+zq6sedxkvBEyfVuCDesSW2jqcL2WJ0vq0wcD0MCwFgqbUiTp6xAi
yII8beoRe2aIeJujHTNLJuTqHJupH6vGwx0b90mKdkO60co+IKHAbKEC8B5KLf+Z
73DIgJ3rk6AHE0vI38aTkw==
`protect END_PROTECTED
