library verilog;
use verilog.vl_types.all;
entity V_PCIEGEN3 is
    generic(
        PF1_ENABLE      : string  := "TRUE";
        FLT_SHORT_TLP   : string  := "TRUE";
        APP_DEV_NUM     : integer := 0;
        APP_BUS_NUM     : integer := 0;
        DEBUG_INFO_SEL  : integer := 0;
        DYN_DEBUG_SEL_EN: string  := "FALSE";
        GRS_EN          : string  := "FALSE";
        VF_ER_REPORT_EN : string  := "TRUE";
        ATOMIC_DISABLE  : string  := "FALSE";
        VC_DISABLE      : string  := "FALSE";
        SRIOV_DISABLE   : string  := "FALSE";
        BAR_RESIZABLE   : integer := 1365;
        NUM_OF_RBARS    : integer := 27;
        MSI_PVM_DISABLE : integer := 0;
        BAR_MASK_WRITABLE: integer := 0
    );
    port(
        PCLK            : in     vl_logic;
        PCLK_DIV2       : in     vl_logic;
        MEM_CLK         : in     vl_logic;
        USER_CLK        : in     vl_logic;
        BUTTON_RST      : in     vl_logic;
        POWER_UP_RST    : in     vl_logic;
        PERST           : in     vl_logic;
        USER_RST_N      : out    vl_logic;
        TRAINING_RST_N  : out    vl_logic;
        APP_INIT_RST    : in     vl_logic;
        PHY_RST_N       : out    vl_logic;
        DEVICE_TYPE     : in     vl_logic_vector(3 downto 0);
        RX_LANE_FLIP_EN : in     vl_logic;
        TX_LANE_FLIP_EN : in     vl_logic;
        APP_LTSSM_ENABLE: in     vl_logic;
        SMLH_LINK_UP    : out    vl_logic;
        RDLH_LINK_UP    : out    vl_logic;
        APP_REQ_RETRY_EN: in     vl_logic;
        SMLH_LTSSM_STATE: out    vl_logic_vector(5 downto 0);
        CFG_2ND_RESET   : out    vl_logic;
        LINK_REQ_RST    : out    vl_logic;
        APP_PF_REQ_RETRY_EN: in     vl_logic_vector(1 downto 0);
        CFG_VF_BME      : out    vl_logic_vector(5 downto 0);
        APP_VF_REQ_RETRY_EN: in     vl_logic_vector(5 downto 0);
        SMLH_REQ_RST    : out    vl_logic;
        AXIS_MASTER0_TDATA: out    vl_logic_vector(255 downto 0);
        AXIS_MASTER0_TKEEP: out    vl_logic_vector(7 downto 0);
        AXIS_MASTER0_TLAST: out    vl_logic;
        AXIS_MASTER0_TUSER: out    vl_logic_vector(12 downto 0);
        AXIS_MASTER0_TVALID: out    vl_logic;
        AXIS_MASTER0_TREADY: in     vl_logic;
        USER_RCVD_NP_READY: in     vl_logic;
        CORE_AVL_NP_CNT : out    vl_logic_vector(5 downto 0);
        USER_RCVD_P_READY: in     vl_logic;
        CORE_AVL_P_CNT  : out    vl_logic_vector(5 downto 0);
        AXIS_MASTER1_TDATA: out    vl_logic_vector(255 downto 0);
        AXIS_MASTER1_TKEEP: out    vl_logic_vector(7 downto 0);
        AXIS_MASTER1_TUSER: out    vl_logic_vector(33 downto 0);
        AXIS_MASTER1_TVALID: out    vl_logic;
        AXIS_SLAVE0_TDATA: in     vl_logic_vector(255 downto 0);
        AXIS_SLAVE0_TLAST: in     vl_logic;
        AXIS_SLAVE0_TUSER: in     vl_logic_vector(5 downto 0);
        AXIS_SLAVE0_TVALID: in     vl_logic;
        AXIS_SLAVE0_TREADY: out    vl_logic;
        AXIS_SLAVE1_TDATA: in     vl_logic_vector(255 downto 0);
        AXIS_SLAVE1_TLAST: in     vl_logic;
        AXIS_SLAVE1_TUSER: in     vl_logic_vector(5 downto 0);
        AXIS_SLAVE1_TVALID: in     vl_logic;
        AXIS_SLAVE1_TREADY: out    vl_logic;
        AXIS_SLAVE2_TDATA: in     vl_logic_vector(255 downto 0);
        AXIS_SLAVE2_TLAST: in     vl_logic;
        AXIS_SLAVE2_TUSER: in     vl_logic_vector(5 downto 0);
        AXIS_SLAVE2_TVALID: in     vl_logic;
        AXIS_SLAVE2_TREADY: out    vl_logic;
        RADM_CPL_TIMEOUT: out    vl_logic_vector(1 downto 0);
        RADM_TIMEOUT_CPL_ATTR: out    vl_logic_vector(3 downto 0);
        RADM_TIMEOUT_CPL_LEN: out    vl_logic_vector(21 downto 0);
        RADM_TIMEOUT_CPL_TAG: out    vl_logic_vector(15 downto 0);
        RADM_TIMEOUT_CPL_TC: out    vl_logic_vector(5 downto 0);
        RADM_TIMEOUT_FUNC_NUM: out    vl_logic_vector(1 downto 0);
        RADM_TIMEOUT_VFUNC_ACTIVE: out    vl_logic_vector(1 downto 0);
        RADM_TIMEOUT_VFUNC_NUM: out    vl_logic_vector(5 downto 0);
        APP_DBI_RO_WR_DISABLE: in     vl_logic;
        DBI_ADDR        : in     vl_logic_vector(31 downto 0);
        DBI_CS          : in     vl_logic;
        DBI_CS2         : in     vl_logic;
        DBI_DIN         : in     vl_logic_vector(31 downto 0);
        DBI_FUNC_NUM    : in     vl_logic;
        DBI_VFUNC_ACTIVE: in     vl_logic;
        DBI_VFUNC_NUM   : in     vl_logic_vector(2 downto 0);
        DBI_WR          : in     vl_logic_vector(3 downto 0);
        LBC_DBI_ACK     : out    vl_logic;
        LBC_DBI_DOUT    : out    vl_logic_vector(31 downto 0);
        SEDI            : in     vl_logic_vector(1 downto 0);
        SEDI_ACK        : in     vl_logic_vector(1 downto 0);
        SEDO            : out    vl_logic_vector(1 downto 0);
        SEDO_EN         : out    vl_logic_vector(1 downto 0);
        SYS_INT         : in     vl_logic_vector(1 downto 0);
        CFG_INT_DISABLE : out    vl_logic_vector(1 downto 0);
        INT_GRT         : out    vl_logic;
        CFG_MSI_PENDING : in     vl_logic_vector(63 downto 0);
        CFG_VF_MSI_PENDING: in     vl_logic_vector(191 downto 0);
        VEN_MSI_FUNC_NUM: in     vl_logic;
        VEN_MSI_REQ     : in     vl_logic;
        VEN_MSI_TC      : in     vl_logic_vector(2 downto 0);
        VEN_MSI_VECTOR  : in     vl_logic_vector(4 downto 0);
        VEN_MSI_VFUNC_ACTIVE: in     vl_logic;
        VEN_MSI_VFUNC_NUM: in     vl_logic_vector(2 downto 0);
        CFG_MSI_EN      : out    vl_logic_vector(1 downto 0);
        CFG_MSI_MASK_UPDATE: out    vl_logic;
        CFG_MULTI_MSI_EN: out    vl_logic_vector(5 downto 0);
        CFG_VF_MSI_EN   : out    vl_logic_vector(5 downto 0);
        CFG_VF_MULTI_MSI_EN: out    vl_logic_vector(17 downto 0);
        VEN_MSI_GRANT   : out    vl_logic;
        MSIX_ADDR       : in     vl_logic_vector(63 downto 0);
        MSIX_DATA       : in     vl_logic_vector(31 downto 0);
        CFG_MSIX_EN     : out    vl_logic_vector(1 downto 0);
        CFG_MSIX_FUNC_MASK: out    vl_logic_vector(1 downto 0);
        CFG_VF_MSIX_EN  : out    vl_logic_vector(5 downto 0);
        CFG_VF_MSIX_FUNC_MASK: out    vl_logic_vector(5 downto 0);
        CFG_BW_MGT_MSI  : out    vl_logic;
        CFG_LINK_AUTO_BW_MSI: out    vl_logic;
        CFG_PME_MSI     : out    vl_logic_vector(1 downto 0);
        CFG_BW_MGT_INT  : out    vl_logic;
        CFG_LINK_AUTO_BW_INT: out    vl_logic;
        CFG_LINK_EQ_REQ_INT: out    vl_logic;
        CFG_PME_INT     : out    vl_logic_vector(1 downto 0);
        CFG_NF_ERR_RPT_EN: out    vl_logic_vector(1 downto 0);
        CFG_NO_SNOOP_EN : out    vl_logic_vector(1 downto 0);
        CFG_OBFF_EN     : out    vl_logic_vector(1 downto 0);
        CFG_PBUS_DEV_NUM: out    vl_logic_vector(4 downto 0);
        CFG_PBUS_NUM    : out    vl_logic_vector(7 downto 0);
        CFG_MEM_SPACE_EN: out    vl_logic_vector(1 downto 0);
        CFG_EXT_TAG_EN  : out    vl_logic_vector(1 downto 0);
        CFG_F_ERR_RPT_EN: out    vl_logic_vector(1 downto 0);
        CFG_ARI_FWD_EN  : out    vl_logic_vector(1 downto 0);
        CFG_ATOMIC_EGRESS_BLOCK: out    vl_logic_vector(1 downto 0);
        CFG_ATOMIC_REQ_EN: out    vl_logic_vector(1 downto 0);
        CFG_BUS_MASTER_EN: out    vl_logic_vector(1 downto 0);
        CFG_COR_ERR_RPT_EN: out    vl_logic_vector(1 downto 0);
        CFG_CRS_SW_VIS_EN: out    vl_logic_vector(1 downto 0);
        CFG_MAX_PAYLOAD_SIZE: out    vl_logic_vector(5 downto 0);
        CFG_MAX_RD_REQ_SIZE: out    vl_logic_vector(5 downto 0);
        CFG_VF_EN       : out    vl_logic_vector(1 downto 0);
        CFG_TC_ENABLE   : out    vl_logic_vector(7 downto 0);
        CFG_RCB         : out    vl_logic_vector(1 downto 0);
        CFG_REG_SERREN  : out    vl_logic_vector(1 downto 0);
        CFG_RELAX_ORDER_EN: out    vl_logic_vector(1 downto 0);
        RBAR_CTRL_UPDATE: out    vl_logic_vector(1 downto 0);
        APP_CLK_PM_EN   : in     vl_logic;
        APPS_PM_VF_XMT_PME: in     vl_logic_vector(5 downto 0);
        APPS_PM_XMT_PME : in     vl_logic_vector(1 downto 0);
        APPS_PM_XMT_TURNOFF: in     vl_logic;
        APP_UNLOCK_MSG  : in     vl_logic;
        AUX_PM_EN       : out    vl_logic_vector(1 downto 0);
        PM_DSTATE       : out    vl_logic_vector(5 downto 0);
        PM_MASTER_STATE : out    vl_logic_vector(4 downto 0);
        PM_PME_EN       : out    vl_logic_vector(1 downto 0);
        PM_SLAVE_STATE  : out    vl_logic_vector(4 downto 0);
        PM_STATUS       : out    vl_logic_vector(1 downto 0);
        PM_VF_DSTATE    : out    vl_logic_vector(17 downto 0);
        PM_VF_PME_EN    : out    vl_logic_vector(5 downto 0);
        PM_VF_STATUS    : out    vl_logic_vector(5 downto 0);
        PM_XTLH_BLOCK_TLP: out    vl_logic;
        APP_READY_ENTR_L23: in     vl_logic;
        APP_REQ_ENTR_L1 : in     vl_logic;
        APP_REQ_EXIT_L1 : in     vl_logic;
        CFG_PWR_BUDGET_DATA_REG: in     vl_logic_vector(31 downto 0);
        CFG_PWR_BUDGET_FUNC_NUM: in     vl_logic;
        CFG_PWR_BUDGET_VALID: in     vl_logic;
        DPA_SUBSTATE_UPDATE: out    vl_logic_vector(1 downto 0);
        WAKE            : out    vl_logic;
        CFG_PWR_BUDGET_DATA_SEL_REG: out    vl_logic_vector(7 downto 0);
        CFG_PWR_BUDGET_SEL: out    vl_logic_vector(1 downto 0);
        APP_XFER_PENDING: in     vl_logic;
        APP_HDR_LOG     : in     vl_logic_vector(127 downto 0);
        APP_HDR_VALID   : in     vl_logic;
        APP_ERR_ADVISORY: in     vl_logic;
        APP_ERR_BUS     : in     vl_logic_vector(12 downto 0);
        APP_ERR_FUNC_NUM: in     vl_logic;
        APP_ERR_VFUNC_ACTIVE: in     vl_logic;
        APP_ERR_VFUNC_NUM: in     vl_logic_vector(2 downto 0);
        CFG_SEND_COR_ERR: out    vl_logic_vector(1 downto 0);
        CFG_SEND_F_ERR  : out    vl_logic_vector(1 downto 0);
        CFG_SEND_NF_ERR : out    vl_logic_vector(1 downto 0);
        CFG_AER_RC_ERR_INT: out    vl_logic_vector(1 downto 0);
        CFG_AER_RC_ERR_MSI: out    vl_logic_vector(1 downto 0);
        CFG_SYS_ERR_RC  : out    vl_logic_vector(1 downto 0);
        APP_LTR_MSG_FUNC_NUM: in     vl_logic;
        APP_LTR_MSG_LATENCY: in     vl_logic_vector(31 downto 0);
        APP_LTR_MSG_REQ : in     vl_logic;
        APP_LTR_MSG_GRANT: out    vl_logic;
        CFG_LTR_M_EN    : out    vl_logic;
        CFG_DISABLE_LTR_CLR_MSG: out    vl_logic;
        APP_FLR_PF_DONE : in     vl_logic_vector(1 downto 0);
        APP_FLR_VF_DONE : in     vl_logic_vector(5 downto 0);
        CFG_FLR_PF_ACTIVE: out    vl_logic_vector(1 downto 0);
        CFG_FLR_VF_ACTIVE: out    vl_logic_vector(5 downto 0);
        CFG_START_VFI   : out    vl_logic_vector(5 downto 0);
        CFG_NUM_VF      : out    vl_logic_vector(5 downto 0);
        APP_OBFF_CPU_ACTIVE_MSG_REQ: in     vl_logic;
        APP_OBFF_IDLE_MSG_REQ: in     vl_logic;
        APP_OBFF_OBFF_MSG_REQ: in     vl_logic;
        APP_OBFF_MSG_GRANT: out    vl_logic;
        MSG_RCVD        : out    vl_logic;
        MSG_RCVD_DATA   : out    vl_logic_vector(7 downto 0);
        MSG_RCVD_TYPE   : out    vl_logic_vector(4 downto 0);
        APP_RAS_DES_SD_HOLD_LTSSM: in     vl_logic;
        DIAG_CTRL_BUS   : in     vl_logic_vector(2 downto 0);
        DYN_DEBUG_INFO_SEL: in     vl_logic_vector(5 downto 0);
        DEBUG_INFO_MUX  : out    vl_logic_vector(142 downto 0);
        CFG_IDO_CPL_EN  : out    vl_logic_vector(1 downto 0);
        CFG_IDO_REQ_EN  : out    vl_logic_vector(1 downto 0);
        XADM_CPLD_CDTS  : out    vl_logic_vector(11 downto 0);
        XADM_CPLH_CDTS  : out    vl_logic_vector(7 downto 0);
        XADM_NPD_CDTS   : out    vl_logic_vector(11 downto 0);
        XADM_NPH_CDTS   : out    vl_logic_vector(7 downto 0);
        XADM_PD_CDTS    : out    vl_logic_vector(11 downto 0);
        XADM_PH_CDTS    : out    vl_logic_vector(7 downto 0);
        RADM_Q_NOT_EMPTY: out    vl_logic;
        RADM_QOVERFLOW  : out    vl_logic;
        PHY_MAC_DIRFEEDBACK: in     vl_logic_vector(47 downto 0);
        PHY_MAC_FOMFEEDBACK: in     vl_logic_vector(63 downto 0);
        PHY_MAC_LOCALFS : in     vl_logic_vector(47 downto 0);
        PHY_MAC_LOCALLF : in     vl_logic_vector(47 downto 0);
        PHY_MAC_LOCAL_TX_COEF_VALID: in     vl_logic_vector(7 downto 0);
        PHY_MAC_LOCAL_TX_PSET_COEF: in     vl_logic_vector(47 downto 0);
        PHY_MAC_PHYSTATUS: in     vl_logic_vector(7 downto 0);
        PHY_MAC_RXDATA  : in     vl_logic_vector(255 downto 0);
        PHY_MAC_RXDATAK : in     vl_logic_vector(31 downto 0);
        PHY_MAC_RXDATAVALID: in     vl_logic_vector(7 downto 0);
        PHY_MAC_RXELECIDLE: in     vl_logic_vector(7 downto 0);
        PHY_MAC_RXSTARTBLOCK: in     vl_logic_vector(7 downto 0);
        PHY_MAC_RXSTATUS: in     vl_logic_vector(23 downto 0);
        PHY_MAC_RXSYNCHEADER: in     vl_logic_vector(15 downto 0);
        PHY_MAC_RXVALID : in     vl_logic_vector(7 downto 0);
        MAC_PHY_BLOCKALIGNCONTROL: out    vl_logic;
        MAC_PHY_DIRCHANGE: out    vl_logic_vector(7 downto 0);
        MAC_PHY_FS      : out    vl_logic_vector(47 downto 0);
        MAC_PHY_GETLOCAL_PSET_COEF: out    vl_logic_vector(7 downto 0);
        MAC_PHY_INVALID_REQ: out    vl_logic_vector(7 downto 0);
        MAC_PHY_LF      : out    vl_logic_vector(47 downto 0);
        MAC_PHY_LOCAL_PSET_INDEX: out    vl_logic_vector(31 downto 0);
        MAC_PHY_POWERDOWN: out    vl_logic_vector(1 downto 0);
        MAC_PHY_RATE    : out    vl_logic_vector(1 downto 0);
        MAC_PHY_RXEQEVAL: out    vl_logic_vector(7 downto 0);
        MAC_PHY_RXEQINPROGRESS: out    vl_logic_vector(7 downto 0);
        MAC_PHY_RXPOLARITY: out    vl_logic_vector(7 downto 0);
        MAC_PHY_RXPRESETHINT: out    vl_logic_vector(23 downto 0);
        MAC_PHY_TXCOMPLIANCE: out    vl_logic_vector(7 downto 0);
        MAC_PHY_TXDATA  : out    vl_logic_vector(255 downto 0);
        MAC_PHY_TXDATAK : out    vl_logic_vector(31 downto 0);
        MAC_PHY_TXDATAVALID: out    vl_logic_vector(7 downto 0);
        MAC_PHY_TXDEEMPH: out    vl_logic_vector(48 downto 0);
        MAC_PHY_TXDETECTRX_LOOPBACK: out    vl_logic_vector(7 downto 0);
        MAC_PHY_TXELECIDLE_H: out    vl_logic_vector(7 downto 0);
        MAC_PHY_TXELECIDLE_L: out    vl_logic_vector(7 downto 0);
        MAC_PHY_TXMARGIN: out    vl_logic_vector(2 downto 0);
        MAC_PHY_TXSTARTBLOCK: out    vl_logic_vector(7 downto 0);
        MAC_PHY_TXSWING : out    vl_logic;
        MAC_PHY_TXSYNCHEADER: out    vl_logic_vector(15 downto 0);
        PNP_RAM_RD_ADDR : out    vl_logic_vector(9 downto 0);
        PNP_RAM_RD_EN   : out    vl_logic;
        PNP_RAM_WR_ADDR : out    vl_logic_vector(9 downto 0);
        PNP_RAM_WR_DATA : out    vl_logic_vector(134 downto 0);
        PNP_RAM_WR_EN   : out    vl_logic;
        PNP_RAM_RD_DATA : in     vl_logic_vector(134 downto 0);
        RETRYRAM_XDLH_DATA: in     vl_logic_vector(134 downto 0);
        XDLH_RETRYRAM_ADDR: out    vl_logic_vector(9 downto 0);
        XDLH_RETRYRAM_DATA: out    vl_logic_vector(134 downto 0);
        XDLH_RETRYRAM_EN: out    vl_logic;
        XDLH_RETRYRAM_WE: out    vl_logic;
        CFG_PF_TPH_ST_MODE: out    vl_logic_vector(5 downto 0);
        CFG_TPH_REQ_EN  : out    vl_logic_vector(1 downto 0);
        CFG_VF_TPH_REQ_EN: out    vl_logic_vector(5 downto 0);
        CFG_VF_TPH_ST_MODE: out    vl_logic_vector(17 downto 0);
        TPH_RD_DATA_VALID: in     vl_logic;
        TPH_RAM_RD_DATA : in     vl_logic_vector(15 downto 0);
        TPH_RAM_ADDR    : out    vl_logic_vector(4 downto 0);
        TPH_RAM_FUNC_NUM: out    vl_logic_vector(2 downto 0);
        TPH_RAM_FUNC_ACTIVE: out    vl_logic;
        TPH_RAM_WR_BYTE_EN: out    vl_logic_vector(1 downto 0);
        TPH_RAM_WR_DATA : out    vl_logic_vector(15 downto 0);
        TPH_RAM_WR_EN   : out    vl_logic;
        RAM_TEST_EN     : in     vl_logic;
        RAM_TEST_ADDRH  : in     vl_logic;
        RETRY_TEST_DATA_EN: in     vl_logic;
        RAM_TEST_MODE_N : in     vl_logic;
        TEST_MODE_N     : in     vl_logic;
        TEST_RST_N      : in     vl_logic;
        TEST_SE_N       : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PF1_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of FLT_SHORT_TLP : constant is 1;
    attribute mti_svvh_generic_type of APP_DEV_NUM : constant is 2;
    attribute mti_svvh_generic_type of APP_BUS_NUM : constant is 2;
    attribute mti_svvh_generic_type of DEBUG_INFO_SEL : constant is 2;
    attribute mti_svvh_generic_type of DYN_DEBUG_SEL_EN : constant is 1;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of VF_ER_REPORT_EN : constant is 1;
    attribute mti_svvh_generic_type of ATOMIC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of VC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of SRIOV_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of BAR_RESIZABLE : constant is 2;
    attribute mti_svvh_generic_type of NUM_OF_RBARS : constant is 2;
    attribute mti_svvh_generic_type of MSI_PVM_DISABLE : constant is 2;
    attribute mti_svvh_generic_type of BAR_MASK_WRITABLE : constant is 2;
end V_PCIEGEN3;
