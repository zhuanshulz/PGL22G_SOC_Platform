`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dIDQ42l8Ax2u4UCvtblZgkfyV/mRN6GY8h/iRGmexxNk3L7QSLKGFoqMI+fgpOmM
SldxwrAoSOAWv/14Af7p7+DA3xULL41ykjp/6vgtlShf9Ba5C8/bPkWLP9DeOsEd
E7mj4Qre/Fv5rDxtYtu65/gz8Rwvta8BHMEJyXNGQ40ArKz8jO1HzvQ+QTem3rZW
gi0pEfUHT10i7YkFYY/M4BXwbCjEPW8pOBa1ulC7NBb4eY0/V3qRFxBd+XCkpYdt
PhTS2MjfnNpqxJvzllIk7Hi1YepnomCC0eBQXvHQ50KresBIJFC3Iehy/1+q2SZx
DexyRdHkZ81Fa5Qa1t8gIiPr8ePc5G6vAdz19EMGHnwUOSE+sfQTp4CrjjZ7/1wc
ONuHgAde22hqlcPFqX4F+EMZn6XBJi4JRoeirsxtx6FYa4DQmf7dA0aX463FHSKI
s4SaFHRTgbB5VsGvrUbxIBj7xcNt9nW89moR6pvyJ52MToaQinwDpB0wmQkoVNjJ
41G1CxiYhCx8AuRKpENGc8wwftc4Pg9PbiXUtXb1Y+c8qNxQtI2Px3Dq4tDj6U8X
xHVWX1PXVfHNOgb0Hmuz1p4cyCIBuH1v9X7Y4LGvyQM5LX4FB1C4PSxQjLYTQrBz
U4xuT62zN4aYeQ1Sk4vp66bL4zYADEeLqHacc486/KHBmMLZYBXf3IO9hYiudCqs
PMM/9GwSB5K9ueZs2Xr2MptLnmSG23xne5MRnTPROAHas71+It/BBYM4CmpnWpnF
+qB1qYbxlpY8+FrctMcFIpXEenBUo53SJZAcq2zavd2/k8HZ9/aKDQm38I2juSMN
F0d5qxItKkVJffeUAVl6F3mq6UN64nPm4wY8Myr5xxZtxaOdvszcMydPdxLGGavH
DAUPbNp6ymZ27FzhezY+WcXbPVT+xiOhMymkWWdJroaVNG/16fn8dkIoGpG9+Yez
pQPlu59YOrx3Y6Rf2baHwpl6VH/PD4hJELA8AQU8h8zDjgvdue2gY8lLP8AeGOq2
df4p3t7I4HMGv5mnaMxC0bqZwLGlV32TQB4bC5/CSuKtg2bieQgRYAVi0Rc+u8Nd
ZRgG96OQnUjaQ5gGqEfHiaSt5w7tVhzIn8t4C4jfzMGkAQUgBdyWG5ygZaUrWUHx
Siu+y65MPgj9hcAGDGN6FECsKdDI4j6Nnpk0HfBmSTtMlrraNf5ZAQsWNeGwJyc0
tvLTcFGnm4Z5euLcVHnnzUNdmZvw56O8GNn9nQ4pR4aL2t+vzry3lDBwlUKbtk+c
W1B4yuvNwvyUKAVQh6Idhax4T5bp4l8mbYhkP8CtgbE9uWTbJ5DA+B09+cYIs81c
lp1H/+6AMz8htEhQTwv+VlGRnROD5WtmCnmRTV3m+szWlwbFE01YVOgLr2GwGFm6
S/2iw56gw1mT76MzTYDvJWXC0QRm7T6v7gJ9yvk7HZhBRNy3sZv0+3g/AqqSZptp
pylHyWc8PKpxpr6dxBTBPjXb5ByqKTTCwJ33F2hDFCY8StllVVMl6ivPm6fHgEWW
R3XMACz30aUKL3XGtTWFsFZu/Y90uoJ1WdXVN/Jv48zIksdeDOkhYsL75h7RsPqf
8nRgYnFm9+rp2sl2ANhsVsPNAKYr8Q/08B5IXale0CoL8YMN8NwidYy3SIxBRjJM
stZTpoc46MtcpJ4mPgpYYQI+gLJwJ18q21BcKHSTAEFqMwGG9eSL4CgTyPlO8r2B
xM0XoI+erZYpJboorOBQVrX1S05/UWhx3+2puq6jsDFdvqNV6vzlJ0oSmn3EdWtQ
pAcq0q9bTK3C9FhfT4ny68ovKbiJI6duBj2HK8kW2Tggn3z8+GyJ4/40N8cFpGDZ
ZH3vwtENGJNfkJq+Q6zMFwFgPWnkNSRVeiloeNpW006byhC8RuSbmTpQSAE4MqzT
nRLYW0LNTw+Kd5Jm/1AIiO5ppzbkZ07vub8Z2YkLCyNGfx4mF8wiN1Q4sk7x/UPD
hjmLMjalGQfxu6T3uzQLs1zfGKOeCKv4301GlwtUsdlGb3fPftuuwiyJhpS0tUxE
sMhFFdvYOYPoGqxVA7ssazIZr3KiG3lC71g3EswOuj0e6/NFMAuH4ffGjlSTqFC+
vyfsf9gWbdBzkWQqIxdRLBL87CuAXrDuZ3E0LblaGKIfptFhj+bwYkktffAiTZv9
PINgNXMQbCg+uCT7ihmTdwUhQ/vFeRRICAKqhctIclEnWaDnxQGnUuz4D+cSBFbH
/Lr4/eqCYJzCnl67xYS5fFjmjbBbJmh63myosjxTQXFvYMq0GaBae4y6Zi3M7oCM
ZZGJxN4otV0GX6ffwZObGqbznLEBiZ9gX57NmrSjRNiQIyQrSRgGxxX1hVzNrt/K
g8rPPuLlibxMp4GT+44gZS7/cGCAdPg4D1rLnPgLjW7Kx1UcUtULRuVO7kokmaqy
nkUzDyCymNPM+W185GyEwg6kAcfodwezOgsh4/QQH3F+SHb/4xZO/Htx00EOEftC
a/ZfcY3uD9a05DAB0Lqtifw+cmUROTxIaVe7XT9CrdVQnKba3UwGD4ijqFkqhiLu
tpHbqREbXe5zwDJ+5cjQU9HTYHFDtf6cOXlalVcpzh/zzgAJgCvFTKTm2Uknh8KT
x1GhCzK725V3yCZB46ZPkZ0jMRZZrsJlXq5jPGeNmUq4+c0rwW63S2mZi4+Trye2
NHnj7P981NCK+OwZr6SdQvr3La9UnXd5jnsBhWMKBr6yEC3EWOqZQlk5cdEytHYL
tW09VOVMf7NqW8VuEg+8WS3BUBcEnwyPitMq6efPTGhRsdWpn8eL7JO9Zoabzgmg
Zvccq6a8Tbe12PQhC8WK9GcXP9zl51dXaqNbS9Ao25bWmIIRed7L2rE6W6thbs/P
EoBnfzoHRGEwhRT9bYPzAceWNkrxJdIi9qK5laBw3Me8vVSVOUU+hYmcoVWpzjtq
EM4dV/E811b5I4yz3TT9sYPMl9l6xs2KVYLDpl5RfN6pjtzU2XD0QbMWjdOgWe3v
WQgTJmoPK76QfrEgngCi7jrpNCZZVowqGUiXKsrTpvFlS/YO+Bd8lIZCi2tDGwbx
h/mhGa+uiPedLkdom6IsONxtRxc9Xiu3KZaphkVHB8eLHJ4kMpZU0wNryTzYqKcA
E2uQaDalIDAFzYKPbUH6DbLOdeE9uQxyuTitkTK89m7BezleOukvDo70Rf1+T4aF
v0mxJb0/es8uuwRVUESuzXRHmtprR5RgA5+ZTmc+gTM3Kd6ObxNilLi2Rwp0W3dQ
0aQ1HoLkpC+bgFrjPnw/k0uxqdC4YmlX2MBpCyB8L4GjH3FQ6VCyotxCsGdmtDnm
yOxunlSQfAmtRq98Zu2dR/k+FTmaaPEM8RrseSOq9DjzQ8EE8uA+gsHNbUW8ZObN
TIUvBZgsdBSCz+cRPLAfJjiqXAJ94bpvJRmNVLH996osqJR7KICKlIyREsGUpawz
pDkUd8bp0taF696/6y0drCdINhp0FjZ6/LIzeRrBH3zebx9HEg4TJ2f3Qf3tZuii
rBiqBo2pnJTdVfxQEcxBXIaXdSpIlkOIUx7SX4OTmkQ3bjhkdl5F8b9bOE5TkQiR
l/LimqODpusKbrPZ1MmjQ4uQHeuKp180ETjJSSrFGKamt45RmRqPf6DasO5SCoUc
NbZg9kfgw1DpJiMoYd3ep3J+KFurVPhMHf/3EqPPIPIoQGRYcjEQstIRxKsMF2oN
VNuuYqjiO8WzfZ/mHEmLu/Y+dduDHygECY2g1OrNkjPJFqrZ3yKvmObPvPUj5czk
A7IjhSKQknnD0gU4cIVUI37iN9ElyQWl05+djRJjjJhcwYCB7ZMoGmVtn7ZuT5mf
ilHK3mr291e31pHmqat9o1XPuc6DLGJzuBgachEHfi+lH/GDr19RF6VgW8OlnE+b
7C2P06WtC8SmiDGpNu94Ib+4AhP8Kg+EU0H4lZvSyuhyUa0JrX2A9uWTljXrVKHj
65oTcd0vlKJKKjEd8a3Djd1WvV/GVTkfzQLF1zidwI2IvQtt9nCxrKZNd7IOzd2u
I1or9wazKctXP5zZ5walVWYIXOyocJfserO6y5KfcJxl5Set044TZ3VzCgPHpyqn
zZ99xoBKsV91zTk3j8UBySB5k8vc5nXgnacE6/D8YAXOmF4NO2HAbuIQa/VcUKG9
qSPre0s7XYbeGlWx8+U6zJMYFJKrqYWI4dfYkS0tLNJLGfoqCNdQdFtIJlT3aPKN
ltL/3fb9oMF3hg+P+WtjO64hZ5BYmTKPQLj3qYV+PsxxyBfs26Nl1nl6ovIPuXEH
TrwUvwyxCWIwr6wHE1G718yQl/isFz0Ko+I163hvv6U/TbDxblAiz+SGSosisRS+
IezF7ve66lgp6441y/ZPuc9qRZccxHvObIeD/t1YCmf94xVDiTzBhxubAIw/wZxe
3Og56tFqn2VnC/ndzPgp+hWkgG3au1Cd60CT4J5Jx63igSKMwIQwoaN4rjKI0ulH
gHCv36yxSnM2BkbQv/sa8RxoLvPEd5iK1O5h+QW0ObJP8YhXfJZBvO/7qZ1I+NcX
mNqQG8Y5e/nvNhkzOoNPkwm/cXg7N43Swvgpn6Vulkg=
`protect END_PROTECTED
