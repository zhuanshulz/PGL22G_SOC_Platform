`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zyCbJcH7aCecTdhI/TQM4Zs3SyOQ0e8nbT2DtI1NQ0bTU+veUDjdCcjysv6P/qNO
4sfj2NVfspEprl6Cgj2mGMX/GXzdwSjd6nGLgooDNURbGsVI8gIHzojEZX2u37Nr
/r9iWXSY89Xpb2pcj4HNOiPPEz11pk8TBbnr9LnFJ3uzM0/PlpuyFDpn0FWpxo9r
UO0pIc7sQ0QmnONR2C83fdLAKJrf4l0gojX6rdJ7HMVUeTpjGaiuXgrzkYQ+5lHT
dvTzgZnXEsuEQmTX8oCaJXgyjzn2Sx8xge/hJAZWuGAeV9xdputM8Q/XwPARReb6
4mvsR/uv0GkTCv11HfeC1ko7jSkbDwPsW6ByKsrxNB9dPsu5cQknEo0MwdiuF7pl
5oEcjm+uHVU6t7rmy6ggTj3lkakte6zBDGtdVozfupR04xTaXgxD/ar0wCIBpxIL
nIFi/vOBGoT25MCyjdrHHQv6vkMd1HWR1X7ZTpj88jUNmFTtpXOVyusLBqIk/HcU
gLffXHRId+A8tQKse7rJ16RcQPp6OOLAIBWoIwNCvclzhh808k3y9dImDnkEZcVF
C66WVoQsdbl7LL0YzpDQi4bps/gbKpvO/PRMPHuoywr3bzUonqca0TJqg8Lf4fOc
1ldz4iFjj03dVvYo0OUm9s9ZNF2t1Y4swQVQt2tQL/uEtA1YfufGGjzmTboiMboo
aAvFDfstheS7mdr7zgoqxh2UrEi3dXPE3q/e0CpYMaB0W9Zapf3uhRj9hbbrjyEH
aR9J2ZECFYkvSgxHTkcJjpL8qP0KVtjINIRXeeL1rQxPw/HU61G0Icvm+mtMc3Sf
jyNAWxuRtqZ9N9F5NSE4H5cpyt6/Z+DCQWKJ5Yp3AnOQqRDbh6xLXfTLXyoSt1nB
oVw+n2//eAMUIuAue8cS3RVuQhM2Iuybdh2jaNxYaTVqawksUbML3eJuY9Qm8GUZ
VlOZnn8nyGJzNLzxrtj3qBdGY6JoHItfjepP8DEqZL8reMt86pml26ls5g4BqeCG
t4gDW+FrowHHnvRlLjYnivulo7WkkJQxPn1jEJaKTeieAw84z+MBJJf900uA7iYb
dxS1nM0Tk6ezvojAzWZenCKurG0rMkFrspX9j79nL1TpJalPgMV0dnvtOdlRHQgm
pYWwy4Ju2nIxF5/D/lOWpQn3FCr21YTxqUeML89ij7w4X2UVfF1MLgqX2Cw32BCQ
oS77p5+DeFJHmaeBnJ7ASvOQ/+htfx4d+zjrWYlUYn7OmDX+fSYJFGO2juTerthk
uRzWtf/n+JrRLfR2dxY/GK9zLhvF9V3zZpKwtXTwBSJBkwtkMpvhTP6w9nHHtt3o
HHyxZ2myi4f/Rba9mFkxKue8ypUNc+gEcN6sS+9BRNplfKigXYIr3HTcnSmJx4J1
82hNuAZaofgTKFcsNdXxHbiIWs8ZcTYreAjpHS1jXIMwjwke4acqRn/Up2ZjYrmr
GmFYke2W7yKM1EjFZcv9WRKw/iOoF+WOOsU24u4nS6QJpTRATf8T3EdoW5VaB0jU
+HMHNvUQQcNW+M28tFn1Plj9q5soEpdJ6M5bDWoHy3J7kuJsFQIqoCnUQ2Ia94FW
1DYQC0JRupH+UB86c0gvrexRNXeaTq/RnFiU7BbTHDo=
`protect END_PROTECTED
