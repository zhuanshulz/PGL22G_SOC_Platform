`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2vohZfybTtIYnRtUCMkTlhGOf7hi0YD/eFWBpsRJJNoZLAk3dUD2wrdC/Oy8nCKy
1cRAaDDsJSQ/N1csNTEnZacjk1P7SkI+c4NhQ917aIdLreqhNeeUrfxkVMc0vV15
Nn6eX1VztkxXinyrlgrAOL+svDYC/CxJuCUIm6jVm/rd7CbeOI3rLp1tOnjnX/vl
RoPx11sec+KTIeHF9kcWMn6pN1FrRqaA6L0OyJoYfUrSAFGolnoJGZtIladBLPJx
qqUG8gC5S6+bkY0byyNNFD+CSDooPsgdnq5jVEaAGHwNChdAzSM9xkOyIlRQOO06
FQ8gYfxQMUOFMzKqUYZY4OHOE52FekONtsGEI1BUpikRyeL0oZFQ0K5ITt5LHc7v
vYRyySs/6ZHR0oYLkfYc7qSV+tWZUvcpkRD6Sl7LdDsMEB48mQR7W4j01E2qIB5W
BfsfDfPwt5hPkHuF0F8z2qHDryRiE2Jso4R6lbQHafqhwU3/7qV4Pc5Y8TMkK7/B
UuR0Hytt0WZEXl48c02kQy4iZ9sa+3EdB6skLvG/HpApdYAFHjhkMlaL1yKtnYIK
CtM4sRvoHQV2dI5OYLNX+nu/B8mpKNNCp3XUOFhjuMAgSmjoP+iIYcy8ndsum7Wu
9CFKT8uUmTuN7H589N35NftZtPxNNni9eItgYHXmJui34TKET6XPO40ngQIeaiIh
2ZPuRs5mYQxRVktUeA9ZsUGSVZDd29X8iAwB898myzER8sqazIqL0hFc8UITZ6kW
6VLchA5eCXj6O9nzGtJ3/+vENBG98xJ9oXM9OE0UzmuldBWG5WxXaGKS7Q4dObzz
10aC6UXqfbQQ7M/6Adg6Hg1Q52+vizgABKODfO8c+FKzCAdNh1b0pX2t0zELBSQY
MyTu5HaRkwTyyLCrkz2SdPrlHd45M7aBaINVcWGui8pBNdi+313b66vXLfwnSZnM
o+EWvyTaysPKLvGBv0Y8uDYl4sJXnjZ+bs75IEdxkO5LWN94XQu7YcGMRu1DIat8
4VllJdsHujaRurCbFp1qt9FIDJsGrag2kwUjWF9wfJul0fML1qMYCxvvIqKC3Se/
VVczKvf4QCO2ThS/F4T2uvtAxI1srFKeVQVG30QGeH4mUKSfPAT1fZ6sIodGg3Eh
xPOwmSvbiVqEi5SSOEAEaqmH0oH8qaSGg9CYJpmkOUtqA6TuPwNogxHjIuIHdraj
VevLYwKWdOHckmsZP/uIRqeGURt41e8W+ru3SAHqFmGGNqptVGK3J6Sfg161JAWJ
Nlf7BxhHWR5DT0BwQOEJy093BO74voNttCEN7yUvfmWvER9t40S+94rpbe0lYc8l
yuhnWmKV4CbAL1o3wZSjCBwDPRGctkNmoU14PkFhe3aaGTSnk1bj3bLh8HutEYqO
9AmPJMzaRQuknjsxUvSDmKygBwLgFqgNTwtaWUfAQBg072xxulisPK/SmWL/wVne
Cfkj22cdibMy1pPnqkFUIjGHW55DlJQcE+YMavkrHasyGpGq2oWUXgHwCAGadktf
8fgXAOBZ2j4zrYhwwdNDlyjcCbnaUxiPku9zN/jyDYayC5X7pJTbbVPOhFBVXL9V
UjF7f/sX//pV6gATv26J0g1UCja1+VzUf4oFzzVs9zpdTuSTHer1fbuoiphZw96S
L6V4TZe0xjcipmAZxno9dwiRR+Ema7TxUS7qQUW2oWjgcxuLGu2kDFIH34GyhpVl
AC0UI15DhOVV6Ix3cyNuQRYhizT6hWnReOpmtga+Ooho6Jg81PatKNTHVsZ8FkLH
bcAiy2QmQpmuODekDqNHwLlwJKL0RDOFmJdXBsccqx3wFf8YwcN5mVcw6AwGJ9ZJ
rpUhIFZnaqUNqxyR3+ZjtwobYYYO/ECDDqxRr85yGdyMZMDcYvXrzdnxhVdJAd5B
MqRfER98KlW7PW2DIDc+mOqr7X6fjz0reeiFGrESZ4oneOlD3EpKROXkWcTRo1r1
1geqLo+gJnDTFB6s2bfFFp7GEqBoA+8OmOzoWBT0BZMge2fxiQtQ1deegFBAEIAP
vTzNfQs4R2YGM9/1MdA0YS0U8tAQMWgVcno5DcaqQfQbOKdZBzTSDYDhKJFbv/0y
uOWP2NGReextuzGHH0+gkElR2eFELxceXdvLqMe3p99Icw7DRLq/FNniQskML2W2
RM3SxmIxbEaJ2Rs3cchYRoqFSYS/VreL/IRUN+w+Cxq0E4KmvebJQElLz/MPmdNw
iFq7gh4wn5FWvJDOPZgrPc6XEEz81ocIZL9rSVGZ8QHSqIjP+HJdpRUcEkf2x3zS
WBHHy9BEtmiGIm7qccsDlGbjhFBBaZUXoH6iX8cRTLP3Vk/D86WnFrRz0fILBouR
rt4dZZBxNUIWWpMmEbY6qgOxHjWBIBZAohjQ43DOEE4IwSfGVx51QTW1EqDGUI4a
TLLTQ4U1P6ySUA3GYqHxdRMYBQZyL7bVmgDtDkXKozPlzoCP9dFKuK52X6JmCj7m
4YdfRLlwGPHuLNC+MuQzSrBFLUnmrWC5w3wX0kNJeC+HBI12/gFPUd4LqNKS98bo
Pj0fp7xhOfO0RTQvggVyetD/k6aKDvULGNBGQ8kDZPXxz2tp+XyDk1nCzLpDp4KN
oV2eyA61WYt6eN7VGp0DHuuJhIhjZcev7gqYbaTC8IubBRsgiXRdO4jCs+c4qThG
eTNlG3FQBBYdBGnj6NvV5wA9++oavKntWwxZp2Ep+P74f4noV8nbo9fkh9g9P7I+
Ak5HZCKGq1gcLqPc1gJ6K5/dkbmi2PaxJ9T/pCHVMo4MfZH+9YPh3QoGMYVyV+HY
Nb75XoJOBGfmRyRUbkF31JjesGZSfj/qMlCSoGJ1Jak6qB6g/4U9JXk+nkmywPoj
7frhG32LrSfrNjHIKzoriWPJFnmFaSS4yj6SCCxuAmRbdDyjmofubzdB5sb7XKk6
9BsUAjaJh6fe4o/xfssA4ghFipTxYifrUMNaNZVEOt1T7o2qMKuq2pbQLiW4IIvf
8ueX87o8jlLGxN62tqE9CWwHandVl/OBUWRzm02+0blZePc5LzWTwVfzcSiX6hz5
yXzlXn2yr/bfY0CN7FaMZORt5z+L0mA+OMrHU9MRl4y8J970xds6Xf4PL8zrunGP
FQ9OrxS5OzC3cvd6jmEOhepNZLAxes8cJOjN8PFbgwUCcHlUywgxRkqecDmZFQZp
iZcrdMgcMzIQHfunF0elCoC+GU4MlKk46qXXk+b8Bz6FzyM7at9qh/5uKwKo4+uM
ZuZgVkcVqQQYbFJT6ow/3EcXl0dyJH8CDJxNKboePUmTXZfZWYV8DVZte48vMRBZ
MMjN9DF6bMjtGmNDBFqPDxspQsHj2cvd3occvyO8Xm+Kpre0kex1fcLf+QC/0ha7
KG7UY4fgCiDHmphfWkb1F8MawOk7gORPhAeBauvXiTW0JbwxUnoCwqlsDaST1WBi
fdUZT/JL8MGX503DLYnKNW+yMbaGraw/u7IFBGhirbitFXtq8s6D+EMDzPDEHIf2
afwj478m6ZbtyGJFYL2eV6PsOIX5FXBio+n+YsejnvztvBjBD3x0oXlkRw1j7hQn
45QGYxQE03YcMW73a4DaTFJMLktIc/mRvronS3/eB2XxbOW3vkalSRaYeCdvJFHM
4XZCj6iIw8CXR3AheIhoyMjj+rNI0EwZl3gqDxjb71UH6wiRqr1tEvPetYSr2Qab
BhvhYpG1BEgczRD+YlB/UyXWlrBCT+iHXkif6oDQDeN28lr08bVHa+fQB7pf4HAY
9H6hl6o1C5oiCBIOJA+PWnqpWV2b2hlHpkXi+lUASETjY3Z/Puj6tadzyXRYKEUJ
LTDmjqhDOMRoAVZTzY/cSuNJUU1To7lqQW0o+LqAKhLcjFHbj8CFO23A7epXk64u
om7gezjgvAcinh5SomyCeB2Ub+L75NnGf4h/58osZcU5yRs3Jif5Vznzdp7swEYr
GX45T4UBkKQ+YHzgYYJK6prOiG/PmEt3zzDX1uF/uNMYcfQ++ozJXTmyVK1prTBX
KLqBEILJZwYWQewfHx340JIXo2chEfC22kJ3wwZ1VLHl45lRUSKWdyX6gaiBKVVX
syx6jCt1CZ37PxB9IuAr95jGt6JpUNGzLat4RGu6wtwmuHnu9kEYtmsPjouw0rbi
SQYgws0cARhLPt3BD6otXix7WeyacJmRNjsXSYuYD2SbB45zfa2QH1VDLj8kbwUX
iwzvVA3iNn/q0StK5dHuMBMxH79PXuoypNRbrRKGYtNiKCfHkFsRjl2i2MEjD0Jq
ns1IU7LBIY2l4hkXezsBZsLUoPbYR3UGAx59mMCKLVFpLUU2SWYSBJKbk2WqwlEE
WOKVF006iWnXoUe9iR4w85jsghTt2FGksIQyQYp0YzNG+EHu9AMGZXXGD8negFXf
qcBbEHEP7j05D5mXq6bwhCErBlFEFZEopEiiSsjdhB1ykZRsGtkg+My8v/DMNNG+
5A6vl2O1pkxrJbzYvWO+LEtJRgKMNy+KK0rgV/FQ779NJYO8vT9+5xTkhLA1DnhB
DAbfirtbVRPUXjUrlQin8pfJyeY4/Z9JZL/1c1AjHZj6X0uM/ZtL3jrZw4l3NJEI
OpF5RNtEWL7jaCpAF4H55WIX6q+jVKR3H/XvM6jhL3eqsMeXXplfNFaYzpGI77dr
A0gTBKaRyt/s4NJ9Iug/6THHxVnoVsdfzbal3X9M9/0DHJ9h6k9QBQk3Wms4VF46
8rHAr16fNd5OIzXUKvfAOkWGPcnoCYTPEytsUCq/skI0uTpAdZ51DmMkJUsp8IiD
7fRwLBCLiv5C8VRx8SIqDI8uUoYXxBNrcBbxMri/+J2rpqUUHRJC2cptOInE/3AZ
NXuKEQkJ1bL4/D+6uf57QoqeUU7f2r4U5ucD873IFrVgBw7BQd1ueeBVkmWgLKEf
nyVlU53foUeV5MH3L/My1h4c62UDw9SVyz8f8Kte3GTt8bg9hfbR7qUmGlqZ+wHa
DglkSFgNl66vzZwaEYkmWgajjH2NijO6vKN3u7JU3mTf5ExqWctDFcjshVA6Nga8
2wOKmOcBgTfBs3PSWCCkOLZraFwaS96Kn2yJcfNxRDwm4gBTekaeiEaIFd0hFaS7
MevWLB7t256orHueIXja1fMCTilrU4mbL9xoqW//ENgypExm3rb3abag5PaxplZD
MKju5z6wEJnAOtbugWj8cU6ARyNcYMa2b1mCMEPiTlQYF0oomjSlgA5whfTl3Tgp
M1nWMZkDCgtD3jQ2zOo0BWNzHxdIuTBSWXUaEkMD2PWXVmcUs/M/lo0UHrgRAhwi
zDB7+7YSpu90TebvvrEz+pNpeNsJkzmCmSAyi9IBsUEpxswgpymOQ8UUu36A8SeY
vEt0As6OVzpeYeCWK9n0LpMV/deCpJdC4+mWz708AGsPps9c3ppKlA76x3IMFdzf
eJ1EN9yTQDqyDGmOFBpd36grju2UqWrRN0in+GVLTEL808H6mf3FSbbB22+YCIt4
6akSgRNPGDvLN7UavWk2ayaNL6TtzA8Gn7QqkhCCnyVp72/x73Ad+V05EwPjOnQu
B21AvU46aV7tFVepDMxlesb4lEpgDK1dSF/tgP9riz8leIAQNg3KhJepmzAD8XnE
rUJ+GMsWHdwVYFeuZiVO1l94SciU3mLFhfsFJxuzJlXnxQUSnW2zjlR3Q/4IJUhY
ISNWhxgrnfLDzk4P3Hfirk/SDeXZ1zvVS6es1DESbAru1IASNfo+8K7NYFtsXOHN
UsPpZ8z+UDtt/zxsEs5JotXQK+Hcpdo9d5VjbKACdrUdvYBTnP5/EtBi8GWCjuGz
z/8n4k0VrI9ExFOw9UtoGclVJJ3hkEkfrKvFlPRg1rrPl9BoidHwtT863Ka5RnOM
Nqp9fDKZFjcbrp1h9iH93zVZxw9KRCV+aFfErrcqqcrefHo6/t+MPTKGjj90qy44
dH8ODGlHuJalVdZCl/pcaxBlDwN+Zt0gl23+2y3W+iwq33IIUjoOXShBxYJ4rsg4
kDynYgDIfX7k3gnYTgeftS0icTTMJAwvf0uuFT4cMPpSenrBYBoAhLTXG00qVzzr
z89qSf2Arkq6CnHoVNWl00ecXWFZulizvN6dTU9Yo2I+MZYSpuqqE1TEyB/WqyLI
z2kVunzPD5/mh1gqJqTCIQZr8dDXQaSfCnXwlRN2kC9pXOcF/uyEjuh5inFyAM1v
l3bcXZcjcMOXvY+j79LzD1V702zEAI6g5jfgsXyMWe8hP1tm+5tVc7ltphVQEiO8
MAHJ3vViuP/7NwAnTMq8uOODUMELB63Mzy9hHTr6k252wNHXCDCdGIYPlrrF8hPX
pcX471m/ZPZaDTzH+YOJwx8zghbP9k/o+DcJKJmrm/g3sQaXgBtLMkiFMgVQWI5U
GYJcdTwXMj+b0MyN2UsFj8fFdLbKwN47tlNnWFUj5+YE3po2xVpYOTO5Go6fUEK3
7fR8erw5LtBhEsEbn1vjDwkl4VjxYxtswVJbz9Wa0DiS0dJ5MLs/ybWvnnoq0rcC
8UWJPBFN05r/pSEzFEBZ8KU1x4AJ1VznWQISh8Q1CSfkfUyo1c1YTJ3B+thyIR7k
zbPhwc0xwPjmAQvFLhwXQojMW/+nazx68MTmEziuxbBse3bJPeaIvB+gi8zEi4w6
v33+5cGumI/Ri54fL8LrNat2fQuetRoz2TDDVymy2f5ij63ZgTWulv2A86/PCiCW
wxgoC4qKi+WKwBTjYjseYn1ITjQzVZRakOBPFV70hljWJgEWuXjs6Culqcqh15z8
hd7IY/1mgflwzh/LfJFJPGk+8rs3J9kThNV89xMdwhiY8aDQhlZZwzPlfZtSOLWr
laQPw7wAXDYjDKjwgGkCeXU6e/hEQM94QC5idRu4FZbno6L4ilCgMCXNLkY7pdYy
pUHYQB7SyQUe5Vsbm4SEXIdcfkOrVcME+ceZZQ8h+qMYgTKGJQYC2qyi/fbFqQLw
y57V8qh3TlJ601Aw/HjQwFydcyMkD9V2NLgh/nZrsE7S/gBKNPA1sLM/w7x/onNv
x9qtLUQvIGrDCvLsi+vohXY8C18aWVkTYvtV7Oe9on4cu9kgj0Bxs8lcoqavayx+
yJ6w+r6zyN/dwoKzyoqXgNDfqYE/dBYuiyPTVR7Hac3WZv5OUj0OUpRstgLQkOTM
PmLgc3HEObB5dzs2DbzKC/gzBzR9n8DRgEk37saD5qKBA1XCSU95h5/9X9J1bmqm
Y6nyFJNq6l4uHdEtUg2HAmsfC3BXJnBL7a3nz6J+z9WrpjicsBPqJYoo6JWGhlAA
ftpkvErSDmWmi6QktesW/eMjBWDKOO5edZGwVnc+2FBLWbnbre83HQb4CJCrDncE
WK8SvR8KJdwvlDhLuLDHx1pnLFFthYodOS3cVM5PpBOSN7WozvtzAyxACXmCwOg5
oiQr0i5bOUvxvGSjxTsf2q/EitA+bGh+N6HcdyqCUHOIi5csDd3gbssP207ce6F2
4n60qrGwlGZ3TMsA9YxwoFE8QKlDSkkAD59AOgpiNTnjHPpnaW3Se7Oh7+j8I1s6
LPTgEMJEL7fXoT3B2h8YsE1T3+XhNBl1BDfxtLQUfWQR13tHw5SQfX2ZfXVIZuKo
R0AcN7P+xFWe+Y1s1ys3oJaZnTctY2K7wQvMrcYpoCe+ECpDesfbxHC/lBWFi2o9
IOIUnYob5kK1swtLGMqwm6WdQjVhDbgIx7iynmng1FlemWBNhpN74LeFJRCykD/J
Ob5mxaKpdVg6mjZhRHdiFys5mjvnq3HFqr5j+mHpLHRf20/8l8xz1aUu9Sd2syP/
Qk8tMq6TLcnU3PxV701dr0rZMNGofjJ1KTfpcbcKRMPxZsCCfH3mu0k7z8V2Fnhm
gJqfPYh+0nkm0FmUACrt9badgKf9AOrc25WkFrhSI9c=
`protect END_PROTECTED
