`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abYb2LA27W5PMBRkNY1+CJUkq+8lqy3xl6vzmQMaFyYHLkQOU3NsMM8Puf9GaA8W
ve7jxkuVODOIz7vk652aX7y2bIO8/BXwThMWIlV81f096Lu3Cls3FliM/l2G0Ziy
ZubBAhOZOVM5MKprm1Fl6Uika+M4nBOMHXToDWTMeUSUhPvStvrhJTXRkvQ/+aGe
2qyLQJXMvxEVRebfcl7vax2Q3M6eMkj/lxCH1J40t6HY+p7QJuoQvgQebhGf+UNS
+s2K9BKWaGxQz6M37I+NUWYF3ZDeb9SyO9lwjntAWzTv3SxDI8RT4C3koCwIG9qN
l20SJfGr6U82kNjmuGnkUAd0xQl6ZiW2/Jj1vyVAdhz2f3jkdrxDwmaEPLjKF7f9
pqR0+KHhOsItq5bUGQiiCs4Pq7sUChnUf571ZeCGcHGwbDw9/wo/1PicZ5pL9qOU
ubcQvmdLiV+IWRNBUCgISgU1ehtD2dXryMgd21iq4qpIy1xeEkTQ6lECNQXZrnko
j51iw/qT3U8Nk/aS32D/OTz8hMMB41kBXbovQAo+KnppBsWNWG2wRDGeTbRmZBlG
X9zJo/M5nQsPUKvIxMXcrfxC4ljjF9jax+d3ZAxHvJ/Gx8W8eWah6FISPjBxTVb7
C1gQtQYx+Cne4NeJ/KqojvUEQljoal2MpAc+HLcAJRm9zlLUvpjKDduqRhAnUlUp
rih+eLZheUtwvbcKqPHh1fLW/08a/te0IZo4/79D4NQfU/BpqlYuJUaQFhxm/jcO
`protect END_PROTECTED
