`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsOJLzqS+Pf04ZN+a2106G3JexQjrvUH8qX6+rtpSolz20EQBGtN4tt3NGXcQEze
w2tPeZS+wDrx21bVwEOki8thZsM1BOlNbT3VbCFfjcazLs7f7W80X+OVdmcvEsrh
pfvnZWupPiiInbSbH2nDAhPdhHALyopfKjmskytcElhys6zhHhQafDbUT22IHxJ/
q8vbnjhAxZGy0lcohWyBlmBJDooyHRE8AeJAVpQnaglImHC2/r01dVvcM8QY/1Za
9njEgCJA7mh275XPM+1f3w1z5fHDDaj/jwYhSukTVlorfVW5hnldcZAFcKfTEzFi
F/0+6IjaTdZE6mb7Hu0MslCsJsWohNJmfrgYmGdL/sqfP0oraZbVsIShiHQof1Ub
jtt7zBzB7loClO2OMIHYk9tZfK1qFkyVBlUx2YGmvAvs9Sw0kOjFC8vhH78W9UGR
LufnfX3SPmtLLoMp+hOQDLnKP3ymAFqC6VZKLy7LVy7q4ARwBN5HImG530t3HPnd
Ar8x7wNCok+xGjU4+vYlIkGX3P/pjZzS7w+AHhZzRNV1EnBZLWFl3+TypfHbmyul
2ti4DOEoAZQFGWPqIOP4tCHHSjLNfOJAQmR5I1nXcPFsLgId8hOhe3IZw91J5RBI
u4t4l8D1fM32RdbDuNlb4YHlKJQ4gkqUkyNGDzmglwpSR5VzOp4PmMRedLHZldSQ
xRkmHXxLSfvrXw4cOzsizYBTC/b+1GH7ge1ZLSloiYh+ebdDe33Qf972o4WwFQRw
y04yYS+rqH7uG9H4dXDTj5LnwtPr0LFw+bCIsVPmtGmMtiaTHyNy7AWc8doiQbsv
XcNzBFrmG/1sCYvpvmonbe7R5ellwSJ8kgFbdKghfRJFx4p1LZW+4VMDZkpWhyqP
bvdZtD5t+G5kF3P7NxY0mUlHSZIle4HTQhfPOxRkrbrJVlD2pIg/1hZkrWpydkL2
CDlb0KkEihfFVPukDg1GQ4b0gBckhq+3zLH+JZDesuP4BTgwIcqHNR5w/UVZddbU
D0DioI/iAHwHw5Ba4v7dLxVB0TFgoT8m4expNnmbvtCGdUK7WSuS3S7XzjddayTA
ZkWirY0bYPqTYG3uOLm4k1JIy66HkdZt+z5HyibMZIfx6uxlbEEkldYBQp/ScGC8
07jV/osvmICsXcjFXsPoCE6o6hcSP8GUpMmyrg6gjEwh9aU+ktunqclGD6RPtuzd
ZwnCbqwSR6mNuNjDGRHKNrWuLf2aR2ehRNrHNnqIl9gPtcErnDEQgYoOtlUdDZT4
JlcHeWfobaa8SBRm8WDy2erIkGnsjxCuGx242cwZaKlfHRG/iQ6mqw++9F0RlRO2
bHgIRdGdUozasY8hsMe1X+NHxg7F6lZ/F+/la5C+Cb73a7ufVzmU7E0GtTdvz4fn
MCoY7GT8dqSqlHwc1S93wh4mq9PojLqtSIAngw5DsTcNEPCWhCyZFeK9xq+PE3C7
qDfDVSbm36Yk0IKa1NJ2AaTkz0E366NM0EO1WbA9Hq+GPk2plOo4ZjZHKzOGiCOS
zKq3TfwfohRPRy1aFhJ/zUArTaVI7m7O6zdhIEyxvyeWxvmXYaZ5o16rtRHAD+Ha
UG5ZjobAADOo+Uz4fZ/3xZ+hLdzFOpPKaJWYKeDqinRC/vLQUgQiS+r3fJokSHOh
8RStfb4hrlS7S05eGVu6arJ9AveEbVxO6curK0userbnNsLqayTuPecTs+vY58pS
94psFJZgUzpUUdEviWywQY4XgMbah8156bezxaughfoTOHKPosr0tFA8GU8TySil
ngm+hIlli6sqX49exQqm+i2ytDeNhxoSPEeW99Il1IaDGPvFdz/Fk+HMKhvMo+Zn
zMOzqfzXZDtaavoZ8PCpRGrlV8kv95JOpbqPrin5E1n7kqlLkzTpZxUrARGGBBZb
/pSbVDGTPDGWzHYaYFwpLRK/DxTMct57pTpvN6M3Pi7LsG2aOrw2mGp0kr52k4z7
TgcGcBjA6fNLdZJetZp2EzYJerc1KlqDJqQ9hx4bCG0zbIA72sm3tKI8VjdtZW/k
2F2Q/iJlUlamBJxZzAvtsLQa8peQFx9oyfggxhvTzB6EptlT/7P8ovyHAIAtOCz6
XvaX6/F88vY/sg3fJe/FGou9myGMS2rDpVHO73LKw/m6r0MyVM1lPyPXqmKd4kSM
dsyzyYVCSWfbpJnzVjWbQ+l/dZAnYXDGb1pyhtW852bBuS26KxH0BkR7yU0L1IVQ
v7N7VL/HaO8oRuWCTNj9T1Y66yNxBHQejiEv4l837w1hTmDgAScJeL9vZNtVCPbE
DXFticeidZ1yjSGZr+SEmPlnvhyVZAQeI/6U13D/lCaHAonEgERP8IkwrV8ICO90
7yZaAcOg2S2PNXXYxNFNPwv0sHPE5lqYZbhfg99S8Cs2oV5uBZA/GvE3Pm7MqDM5
GuolgXT819DV47XokWahpoXEjjGn+W2qAX0A63bPBazNlvRs2DP+Ox2CbbYok7Rx
7riOVMGX9fUOv+ipFClmI5pQ+PLkURZooNZ/xKA2TTJDyOR6iTba4bxx2yHHWUKU
m0483zaiQ4mSUlHmAxj3wVzQtg3KH3XXiSU7tvAAebS74TYBo88yPwsrGGCz+wpy
acGjIwSu4kNk/ZB/hvJ7/wLLy2KC3uxG0nDrkKdVTPDz6P9aE+85JfQBWmHsS1Y9
CREX9Fg+dRDg397e/T8dzVFqR31xtduyBc1DCcyX3RmOwPsZEi6aavO1MS/ecpy2
zvrfKMaBu4YcMYcp2eWPpbERCq9X3n3v+c/P47cwCfcdGQ45KBSNXioMv/hyBgxc
DI6Rugo0v4rCvvZDH0T/Wxzedw4h41mzqcqYI/j7tjEFlJ8U8hyTK/Ciqh4AAy43
D7OT16VFcshmGAcjoG+uYBc45mObaubG58g6mSJ51IeeDNxYT1iFGHWpW9pyMD42
DXKUUWHGOSvpPNCEW5sLoA9dk3P8mDE6IYe7nFWOqwIbKPVTDgsN6qCkKr4CMvxb
lrjRSVOj9Mzw/gqf3clB+ViMFO2AroSX7gj1T4Ro0g7+aLkIFInQ4Jxhq95tqO3P
P9wYOTToehtF+5Niob4ohkOqtOJlHsigu9k/Aajo4LVrNjLZZIhopSj2IzIKeH1n
k96TQoUgZQDL+Dy1w+jXfAEMadvhcAXtIkgXA4ophNFbAgE6DPM6nzwjMiTyp6Ek
KgJ8J5lzGkeFEA0qEu0lxHRE+ogM8/rAhXG1bixUb1VeYtjeRn9YM1PGyJHyKEmL
f+PabgaK9k1wBi8IZsMdr07wgh0md0PYxB+RgS2SSh9xNRO0O6X9Bgzs0UZa0A0M
ucF42/EYfTxDPMB5huPrSUhum2+UkbNKWbOpPJKMlpfFH77Rku62p6areKycpqkH
qsfwHC68nlCERvoocDETGOUN1yoXmdfOMhNowLgzKvgZqNo8w/tAFpPxoSXjxsaV
nvWR8xBuRAD8ReQwQyBwjGmM9vswEyt7YRrad3d/eIRrYXw58BT+3YvzOmpxoG+n
MKdfgJ2+3aQUglkuUoyMwnuRsGYK9UVxtAPyYBJ8KcT6VOm30cIWBbaTIgjB1C3u
7UXvJFBnBGtLjxwMngmqhn2SpfBqyDEpu/mwx0qT0Xtdyn99hQ+hsDwV3EZPt0az
EHu8QOMu7KJDqa/uK5DGXw==
`protect END_PROTECTED
