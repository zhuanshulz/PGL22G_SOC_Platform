`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh9GtIyzDfp9hj2C0+UQ+xwNaWjkswpy6/XR32Dg8RgzXc9LW1mtpXhuA0Qrw6yl
rz9t5xilSaeVH34wlfAI9nrNsNhfEe6bRlEmL+vZ6WVO2b1c+NDeGNNcDZYjnjkz
R5l7s4/kwuLPSF0T0hx0OgdBEXKVUNZXPAViUM5Dv3JlVliyjxuZOokI5n2nTNU8
sW9RifBa6lj4nAlGrfEK2+Xex/MN3/uR7kDmuMUOeup1VmAmGWI3eNcc3JyxD4JT
4UaFtTLX2YKyVEIRSbw5s7qTJItprV/52CDfqKOl12ztYujW+mVsIdvevk6T6fRi
ZnsgqKbzaFfHXxQSVWTyj8VyRB6uT+QjiK0rE1aXc79WkHXb3JGWCTikkKCjmuVX
wBfpLbXSxy8qfepOOt5HzzQdXUQi/CzSxHzbS2o2dUjNmjroUY5UGKguZczvBFmS
4t5Ly2NVS0sFlr9qmnoxFSBmp4FQE+0jRj4RsIWqbwP47sbmJ2LVq6fzonOFZxg7
+86jTOPJX/IqRy97bm9z4VPZE/m84qM2qx5J3Q1MXY55/jdvrGaaG+eM3K/5em/m
vEI66Sjv+S5xAflVCxaMMVYUj9n6bJE7N0+2B33JAl6B+XkgUc602JD41hGnxKtI
vcmo5wKJXnyPBv/zLe57D/SngDcQ7YZaWno9LxhCMkY0uV10vGPwdT6Y61YzH270
iHOlHSUhUe9RWt6sALItKV14UPxwJfhbt+scmSZGkGN/kDqKRUgVNxq/T95y0+Zr
`protect END_PROTECTED
