`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xzUT3IKGQ0cHG0rx5GKJi6AtwmjuU7XQilKqbmDt3ODv8TwdikkBi5L9yET37bgw
qq4dG+n/8I9fGNeyh/NVtNvc2MOxH+hFE7spUBxyir860Ow+kyCdV3t2oOvymGxF
651WpSGQIr5prIeUbAkEH1zBLQFj5PwWoF6znY5pb7OibrT39GLiftt+EILse7M2
4TnvYuwY6A3YlDkqaGBWYHHmlm6PzXMsK6n4vYiDCDclhaNQBi0brWUH/iqEOC5t
JGcEEh6vjQKqmcrAUGsmnh5b96nSW6w2a/M9ux/R9qG6dQT1aV1YU06beUS7oaIA
lptHQCvJyTs9gvsoZhnFhIj9T+gDBnHG88IgnR1ON0FcJ9oWuVMdj55UWBP8GrEu
97yroWmB05KC00BkRnY7O2iyHcFz8SIOiGiYQsg1Yh55jDnzaqbz6KqbbbA8zlU2
YZVnv9R3vVmsQrIJojd0qoQSI0HKpTxs+Z9jq2JODxvlqFc65ISu1fGrox1h6+kd
uEon/hq1wGrVIsN7dE/ZhlOBuTPgK86Ila1RaNP3NOq5k98xbBklxbXodD9l7WTl
n3g6nZH/uZ0weyLa6Mz/QrmUQWEXF1mTcV9KBrfJ1b5Wx1gosR7dTqnthn3e88L4
Ue0+ufGHKM/k+QyYgJjOWm8XrdRM/Oxq+CPz/ZlwSs+kgaH1auRiiW5pPgljDsZ2
bBhZMicTkwjegvo5+Y6bP8pH/1kK2NybYctY12PKhYc6+2VxYih9NPY9fVj49DyQ
zMvGX7zMpJTKZILceBLwuaViFDoLaE2lMClK2rSoLfPPlYA2jMsrnNhXSMeDXfeo
ypoDvmdArdDZzdW2nwNxJE2DdV5lFBmzG1QeV9o7YmweEPQh9vQrIwJQ1mH6izPs
agSY6NAFqzXjeeAo0AQ+zi2O+K+13qVafKsT9iQ3UPWFNr9ROmT1gIzf4/Ogf6GN
Ev/fBxy6USyrl6nqVSBYkqUSc+Zs064IzmfA372BJrEBQs2BysU1BoypT17hbAwW
6i+hjGeOIlZ+4jVjkSE6uTuGOFnroXpWhsK23ST9qzsXp83/nunFegcwzt+XaSC7
/Bn5Z8kEiYSF9S8EY9036TonXG+7tNzwnqkwRVMFbpyEUDmc+/3LNSv8pt1zyxKY
byPiVyuqldrhPPKizbs3AG9QhsTw3t+CVXKKUkpXGak=
`protect END_PROTECTED
