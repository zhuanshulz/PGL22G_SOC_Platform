`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I4FcEZO9AU7MhzT/NdaU0A8m3oUfmaxv6nUD5yjIk41MpcjAOPclEHzCgzc/gsQv
BIGq3DXIH9k22nVWJfECfiwQhuKdfjIc++L6Gd8WbreEz76Sn63Hw2Lp3JOA3mVG
gIyduSXefmBgb2Jcc1tUh/sprCTg4JIe5c1pXQr4hf7bQRpJx4F0bckhY/M/gKuh
qaA1ih6xfRHt1LxpWH3XGy95C/4J4yFQyA2/bl5qbEtIHsZ2bT6LVllUZZWxjTg+
s3DXAzBczozZV2F0FUx85AeuUoz172ES/EmJKc8ZQwOI+kMjz4RP/5CPzYfp4zZV
82dU0kU2rIEDsMogvYYxDiHr9pcFvC33lTqoEekZImNqV/IxFnF69JJT8O8bLD/L
wTk3m/JkwKS8IYrk0VhEbi5sgh0bXIwBbUjr5Zyhp4tU6x0Z7aKc++CS3kYR6MZc
Dzl8SmJzzQp3uXLZY3z3tt88kIHN9BL5A/OzVf7zq/A6qWbg4aGpGy++CGPekhna
7uMprCIX6U/iH1/jZbk1zpo/d6hnlUVo03NyevCC9B7nhZcyl3mAvvD5bLa25bqs
gJ6nxTOr2QbxW8BD6JlyTthLnXYOvWmzXIRNZDISVe7lYrdQFKfEwLAePmKC8Iwo
2UEXUwPJe3NJn4WVp2xB+R0EO81oi87idscSA1xL03eJJjMaFbnsqgnYBx3nQSIC
B5k5iTmy4jnJlmi2u4fusYp8GzNTOAkPH36EoLgsv9B0jGUpbOajhPDbYHkyJKi0
nQ8OcSMsgg/oSQ9EeE17MsaN4RS+Rt8s2GlyqkJ+JaEBBYe3tzefqiHtejPcDci9
udtceWztqDNfkZYW0k5VrETIacfd5t7qef10s46ECX/T+Ub6/Fpkdnqe6VXnR6Pf
W/RgROaS39d1+1Ff+1+DYc3pENrCQuu+KJrLKurmfeO0UV21Hlo4Kj3UY+5/xwSF
PgZgXPGjOi+kI5jdDrW+jN2mrKsf4xszyVoQIW5lIf64+nbBT6EAwdjSRktPY5oU
PWXQjI6Jl4UY8i2lkIFUkf7bn9iVKRwNC32hT5kjPyfxoOBFiJNIc+ulRxJtTq09
vGt6oohgCcWP/a4/SsxG2vgeSjkDGvLaw4CKRXlk7DhDOBWI5/+xa7N4aCWGCuAC
7ytRAYDl2skyLJzjMmx5Feq0dPtXwsAKOb9ECBXGW0TQNWp/7PrNJmpTeflgKSUo
jh4FjSWkgQaAvTOBOzE4a4VUA30jFH4Zqlz88riRmPWRIKO8gJAGt2DFXytGlkMb
1lNG1As8u7sZ5bR9bffL3Um35JOfgm71In7PNFibpDdUQW5VhQXz9LokOhyRAM6D
4F5DJBq+RlybCnROqlYeJ7etUCuNXjTCx2uCwqWUaEVZ7XRdrS+ceWQ9Of1rWDD8
4KRR8fKKt3+AHoZt7CMY0mI7+UbFQ0U1tWL1UdzNsDHpubfLKlk6tnEq2dqByA+M
1aJHl7/CCJNROx6VjRXG9W6Toiezxo21VQiZ7GhN9INEIG4fgaRld0WIlBdWfgpC
IxCV2ZZa/SkATuFn4XXr49qvzWZo9omS3c0oRDeGQLUkz6FuXWMbVAjIHDBaimYA
qWIqoIXD+U9n8kWgwKe9mIk+dS4pfjgIzx+zWh6A5gyO/oc97OMQqRmvYl+KgwHF
G6GiJUtdWntc0bStNk6uEYDEGp3v4Wg1JSKRQ+uUW4azs9Mun9cszBrR3B4+9O0O
vWQbBHILxmgUFR1G43AiUkQQbxe3GEu+ER0FypHP+CGmwyY4UiXKYv/av8jrEfUL
gwU4NAeVDsZFFdm0uDOqbZwq068Slbn1LMcHG76pvg/pj6As38fUg4+QBMQqZlZl
tnE0HxHo7K1kpKQKrr4/uacTRkljoa1cE2nLKrspjonfxUVWS//rdjaRZn3esVl9
uve3/n8JKTGJX7+5XI1cqZ2ByjwL1Xf5UkF21HDGs07fYysDPxmgQe/wCa2lm/Yu
BvQjxl8ujbhyFPf4IQuTdWr2BJiIj8jIaJ6BNqc70aG4+Ov1AWV5hx3kVL2qGixF
RIAYuBCAre47YtBPHHKNOqBmlihhSOdfyke5FY+IqLgZuTCxzgM0w9HPUtx7RgaV
kR9qgfQKYxumxXVVmIL6d/ecq6vu5LJT+meJJKXhWZfPJCb6ENDD2VIbzPh6Vs4i
XGiOX70NrZBn6NZPqS8sVsDvfcuwbp91aUbR8ikotbJ0xusv8+0qx3+ONf5ct/bS
UK22Ai2KOY+qVIkoBwqLQGG0EtxAvXPT2wg5UDIaVNkT+IFjPVNGpidSBl5WD1Em
AG79Zc3UYXR2OMJaxy0/4J9YKdDtaLV2xIT+8s7OWLM2/wqVZlcWSReKFiLN+Ohg
vtjz5Wpm/PA49ehAbDrpobw2l/bo7dmU1y0e8pElrfUVbcrmulWX7xcmmUMapqiK
LRlcWJFxq06yDt3jcDVffb4bKUx5ExdiR3ehku//XiFcds9033pfsiVehpKnfX97
49USfK3/kICLxOH3V4sTZboauY+zG4jCMjMt6qdul7PxT3I4YApprf5HhbWJSWM/
rbWDbi1F5HCnmeTKooMV4X01nmh4IWEQeI2a6OiChTWffmMM2cu/tqw1zYzLbAH6
a2wZfH9vFiCyGYjeWjhf08um8RJxtgQI0YLX/T4oUdWgKn1+x34Wyn5dTYrbB+5P
8AsfsgblcyXu0WmWQbSl0o2YXiqPdjr+2UZFZZTww56+cLmTcGNHGpCu8Spuo/cb
lXd7BYbFVu8/E9DbpXOqc6mU7OWmrRDYl+a/XcgN+RleeU1/+X6VQS9po8GkwtLO
GclOALgD0oQUVadQjwNhm+ljFK8xqANVWT+ICbspLslXZ+6wClrOqJiDCvqg0/4o
`protect END_PROTECTED
