`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IAEz8qsgTsrPiIjajuUvyexExwJA9lzPsMHejuHQvkAzW4123Q23rZCpqRRw85k/
J7l637Ho6Drb4uCykPKOC6FHIhPUHfJ9/Xh8954z1jwBWeXr4oWvZA4lGRiSxYyJ
ULEHaYnqSwfDDST7Wg17GhDena9QvbiVzy6GYgxOt7A0g2iw7IN8FmgnkNZrQm/d
J6GYKMvSMeBbnRNS4p4Hu+6WN4fQ0gSImerQhogCKVVoV34YtgU5aOaZdNqzNvwF
FcrJ/+g81j9904YLKc3mcaydtPxXI9TkYvcYBWVfon+mqB1IAi478ks3AQ+hmqBl
ogiwuyJLqbxc4tSK5fUHjyyKNJOxjDFWOIWC6NmV3WkZGIN6iylmdm8WBwgZsgVP
2OkaO+xPRXtEV+P0X5ptBBSLVfqI3Iba2AvrJCseNV/9C80dmC4akaq13V4Q+kBz
5cTYbBES0KPxNworDsiXf9KInKpEPcq6YeB4cEaPtzhRJrnp02fml1T7rAZMCV2E
KHavSIBu+DHlJyeyZ+WP/ne8Wxw+F/xJ3huGdpZ8avVPJcGwdYYe12zeIXeQ+GOn
OZ4OvqpekvXHubJ+LchrFlsqnYCHeR7ZEjtRbf3OllWxns0PLPq2cO/o3JK6Cosk
FuKdvFq8R1yRmzXJbYffFDk06lBxy4h/XvYqpComTmofO43i9aQsjgIKipfN+bAA
S6fWElImcDGm9Pd3Tkn4IWsy0p9CigOnuY3RVtULREs9scqXjA1wbEhS4pf6G3MI
Av18nygsVtQSyQyqXwBPNMKdjiXl2AiAbqn0jHKi9B4RYfPvmcCKNZcXLKvimqzl
qdTA8oU4QzRimdFi1nyWScBbeqv2PYTocEwnlzkz7G92tvAaUSEQkPL7+w15H56n
7YL2GOJ32O0pfUVLmtB4mRshA+WAPIM+e7QHmL96lv8fVNOX/RJNToFAVGcdde5R
6uKtKLTFN8klhApxPVuypGC1c9AMbIwnENgiYqv4jtA50fJbiIruSeuSKBaAqtsq
NNpkwoWQBuz2nDh/bR9v2P6JaDYHstfKbSQUH9QcuHr1iYXkoPq6pLatW3Ml1JZM
APjkvEHqBohuyQfhC8U81PMmErv2mR0RbUUzXCxpytZJ0dnZEoC4+/2V8vgxi/kl
Wg4FSKGq7VCqT64o885RP4MUajuc/UADWFsyJhurqyKQrlF3PEyRZ+LxdrCpr+Fb
QIU17mEkgsEP5bxtZrI5qmHXVIFTzpGvhZGngwgGXELV9iQDUV5huyHAzrdbfXRp
kgmb98rcUoxJqpgLyqdMEpQjhOEaAJ1nMyKA+zG1uzw1G3gbxU2vNsZfDKTfDINi
+zyZWj4F+tn/y/2FuR7qh2PpPYeo/SDPXyBstU0RfYI86v/QPgEzSrGANpiJAZut
AR3IKrpYzTibOKrDTl8e4iA2QXwP+usEAaJjG0Ajk5jr6QkLjg4+UHahQnJljgGM
ZoovP2auh232Xlikup5twUUfIRl808jfztjW94J3aeJeV8YBUx8ksxqDP8ehAdtF
Nu2nW4kb7dMsb1Lpfg8cpd2KhATK/Vu0tPrF/Q0lmjzQOq/d66x0BrirPNhzDx6x
VL7chltJARWVF5+sKbMU5B96st2J5DQWjI66oXVuHLvBcsSu3oehTbA8MYBALZXq
bZpofzEjI7+07PMc58ck4apDsVrwUkDEYNz4ekovvM3wQ5cDFhtqEZD2j9AAUEEJ
jKzQ2sSYuHZd23WcAqHZpC1CY4jpXe+pwfNXqliFxKmNL3/LfwHrWDv6VDB0bXIc
+j2y7fcDO4tLYDKKkwdXUePqIBcEgh4DYsd/QTyJcGaTUOeOZDZIwathXVz4Fnca
FeTuVGJY9QudnRWvs3FXboC2C5iASnIqn1rrCnRd8xzRGlRKUvawR6ImovMEc5QW
rAhXa68Do7qkdg+x0r4Fmz7ELNQbn33L710fPIv9R+o=
`protect END_PROTECTED
