`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O3no/bU3A9U/dj2clV2ULs/OZLmyHuPyl6NA2CgAt9gFafO9orqmQ3NqBBWcvMsK
UfVfTuc/j3KxLL7r00+Dmcc6s7maAUMboy+D0t6rbfQbr4RIMVyHMXrBO8vVWESY
axx9f2GZPgEhrQ2HfFT3VEagqIlmv76nOf4lrBng77rumOD6HhTUz75FBJfrtbHF
/Yek7SnpG221oE7AUFpNFY8PCX7ZcFFo5Aq5FgSIPth/ADD1562zs9ju2KehETb0
P9DZLOgdgbnsLLYGamWOXnGMszR6sEkYnuisph/s6REhqrVEvp+gd3ys49sOTznM
5KOwocngYFr4jsjiCb2EIjq/lPZTF8KWWrN2KLPD/7AU0uvGIt2S0f258xCCyy3i
yGEivPFCkBcwWol3XcvWdgfV1ZZebVU1GxJ47902qqBOiHwCxybNdrv/JHd3WbTN
`protect END_PROTECTED
