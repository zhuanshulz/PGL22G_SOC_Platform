`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Z0u9IVsxruu18VdQV5LL/Yasj7BzxjoYTvS90gMpr4Qubps1jn7UdTtyd6qXOFJ
PXdhLzwNjsrnfwJlu+rVT2ihxZzrmkMzwDFWU5t55s8ZcE1gDrqpdPKstl34j1nD
lEtttPMOtDozlVVEfPihVS8+7nNmpFdhCPky2QGb/8vah6A5Nmv+drvU5cQkfdwr
EwgBHpeYGPgPL8I0MpmRM599MBl0TMIEGmSBF9WMTHLJueOxJS82gXU30QoYDbG5
quR2DHbyfd2DIMgoqqzt8VG7eliwtjqEiOYHwh7HRLZlYwSjnNyAhMUbbP+xI7yp
O1eKyQeqf8HW9PDvUIyFD2/RHJn4YWxvuYsHbKCDxZO+4gf7eDvKGFDTo/0SOatK
qArHtiorpTUpyrHX1HZsBRPipKrlFNsvvymInWva+A9v37C+E4K+vhgwHT8YbdN6
15MaHOnLeF5YkamQyLWIzhWH+yLvoN60HeLzhnPqR0+RurtZsAZyXyyWcGApA7RD
LsEao3CSqkJ6bhDUgD5UxrIBHRcjSkl/ef4DI3bhPRcXIFwc4PB7G0RtfgFPTXuQ
/tTCvP+bV3STP5IQ9y0lGe+xBKj75u4RuMVymRUPscINql8vqn4OGqigxGxnSKIG
lG9OKYZV/w6ZTpB8DF0TUR8xodoWOVtlVijrc0qL5a4jNHzOJ39qJA6EDSqaeonP
idIJ2CvvW2qvaKXmiydGi9FWMsm161zZqRd0MyBFswWqe6uRctcQ2iiSXrfLey/F
AXdq23hc2eXl5xKoq/oqbvQH12RKoFPGRMdX5ikb+1nRhEJFqB95VCFN3WmS9P6B
2P2RwxRqEFl2x2eIPt+xpMaH5oKeDk0X25DcUBjHz/RP8ICU+U47qWbyQQqoFKP/
cRk/Y78YJx24ubiZNbm2CT/6NpCgYRR34MGVlnns/B0SsmQ7H616eQgZHfpIjqTj
CIh9AiAeI6LeKXQN4PyPz3M80w8ire1WBQkbQ1lBAtr9viqtAtWfM+xrX9kNQAi7
BfRUuTLBNxXIEkPnwHzlkE6In1BYBEuUYC6c+UGB8SynPRJHX3VFOnkPhGuPppjc
nzeGQgZof2YIutXUCDofvr0vM2cPFAUqN+iqzv+zQWUFxLYM1ttuYAU0A1qbpmpn
yqNd6FvScXVt3K2A9ukgQqsyildP+HZ0sTZgWgPn3r7RSXgL4fR2x66wGmyOQAtE
muJM6SQWfAaPOVPlJpkxtIEWTR18AZrDAZffy0o0Tx+IlDhlvVTp5vQ7gjiRwDMV
AYVDIw4JXSpX+oo1hJwDdi3Vhg1MekVB2TaH7p/119WAHkqKpLYnSsmL2bsKupvI
he4LXPFrf2/aooldDfc4yj8MyicRhE0/rKyZa6eRW7RGvoqXDpXvHZbXL6aYSlyh
OdmY/lLmtnybvIOZjutnAqb3Z/HJipSXAWVxtys1aQqGOc0XN3swbqgVFasvhaBa
O/p8mogxwAOp8GSTcH1e5g==
`protect END_PROTECTED
