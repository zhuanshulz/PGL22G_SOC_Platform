`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4LA91QOBKc3RreyG2qt8J/CQYMhFUN3z98zkCWvsYiDcb/CCqskaEaXsERLcXbjf
tR8CpgjeKMkcIHfetib3xzw1sPVw53/U+Xo004ijlKDj9Cf4ZZoM2VN621bK25na
eP7W/Jl4yVAtsGeCGJVm/yNsqQZX6iY+bOFaNqlSyC0pLd94M0MztrK/sD+YYHkV
AB3i4J+TnZDYTmYOmNqHPgN2qcR76aW2dc5WX7m1eXpZ1ZuZ3MW7aMzsCIaNzQRB
Yb8LIzgZVk+nAGu9cNc07y5j0NQMbXG+o+bXbcdZzQBfRjGitR+g7DOc6+zuphcn
JNIGcS3FZgV4o0ue7hZZEOScGGfpQzDionrt8M17FZgTI8rnm6j64B0G+ZNk0g0D
UHFsWXfDFFJkvf3Ir7MwuYtKksqlmnRQFl9Dxh+BhjAzxK9n7rBqtf+sBVi7OAsW
DpLJiAoitErNGL57ofZB2P99CDTHFDRwGnnsyJH5xdi3njaQz5WfqWgzepD8WZuq
Dy7t7zHU6ZLPLuICPmyQqPu35WuZr/AEyH3d9ni9Bl/CT7nKO50K/3wq9DsrKcKX
mAdYTdju0W4GdDoAi8rYb5THm/TINxQlqR2763JK8gsYEjz07kkIn656HWfsiVtf
mcDTbGZL97NNZjxhAaDF1lL7AWuqv5PO/IQ3NDmokD+ol3YtT/MSqGadCqWEFvB9
4Cm8iIkMMjgjqfrzqI2st9eQuNzYaz6NTmUP4/E8VnJe0d2qWzXVjMn6/DdGz3HK
R8+ecXDbZFS0piYoXpPxE1Kmxkxei7oybPdGgKnPLblqkS5E86Ra5hCs7N/fu3LD
MVcALkWT1uT+Zod60kYmce3MUrH8cFneISd3XT2Y2DQA/dGWYFPn7xqLceJgCZie
jU+KbZSmPoEBvPBlMkmF9jxMgl9DZCi/5rbg5NU7qqSVu5Rck+JvpTIpERxO3ccw
rwZrt/FBGUjTcfdKUoxCQEboDDIJGQrpVaSOIL7yV0++hTDu/rfj85nG0YPBuIud
qynrMJMrrmB417y3mIUA9EfaVFfj7BUmE/HnhoiMCMdlBLi950KgRa4j8TLlwBWg
4Mp85L0THnAfcxg8jrSXEMkmE4Cp8nAuWdB9RX6uXaHHLRCaOfnIeb6t+JW7AMoz
1PMT/6fvu5ROKieIkmzoWwk3XO/FRAYaVdQjyWFPjbm6qchRW/X9vwHatEobpr4L
YsFjfupFePHTRkIoLFiVg9gkrF0qxd1b4FIEP6QSJkOKP+ZU2ajLQMI/HCGOhWEq
wOLB9yk45RzmrTlflYKyOH5x8bGBi8dan9aMP5I4JT8TbF4UzGoDyu63aZeAn1Dp
BX7AVOWmsvUSWYdnz+HQXMhb0Uxtw/4e7RMqtrqlb8b6ZSRio7+K9OiPaBKt9xU3
VcHyLpvLqTIuK9FoStYZ9PZyy6qBcC3+oz5Fpe3TCKJ3ot3zP/N4KyUEgSxAVBgd
z4Fk7Ux17jj9vyInjgluPw==
`protect END_PROTECTED
