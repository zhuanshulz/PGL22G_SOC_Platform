`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JmSCf1bG4uB9lqJO6x17+TRCz1oeiURkcsUP1P7QCojFdMdWFK8bNo4o8Zl35Jk
foQipH9IUbE/jUK77GDZC4iAjIEDvIko7Ksapc2FP+R8tBE9linXjej+p14e5Hk7
PNx6fXp/ibE9027vYlAQhGgL5rjaOPEIfLi6zg4oOPU5BRQb2pt7lsEmQ0cA5zCW
9kYRyi7XSZMnI+SUCmQcJrdNfpkTi94EUYSq4kVFe2aJQ/KSKvOngsS24R4/T+0M
IC+E15CbFlEjERKp0c2KsvMNPMXf23wwQye7O3KB+aX1bnuWmXhoM4MqdldIEQ1B
oh7t0oZNWDD/YwZ3dx4A/dSdzMKFvpTNx02IjCgzmxamyW95i+NlsaiHrxAkxE5y
ZYFyj76Uii4i8tIE8veii+6/PsGWEG29cSJ3wE2262s/CHEs3/dS03LrfaBljU1P
oYnKKs5MfiKWVccxLBN58hv/7m8LNtDoE7cuXLNWiIFIa6YYwgai6XSdVyEBEEsZ
mg2ap2NsF7C2fxP/da1QyHgVmpCZv5Y6zDsLJ0ZY/UvJ/LcmfkFHGuWXqrQqt2rQ
UQt7BIXYheoc/+BfPGRZ/3rlQe97/DvGaddNLvjDMPhhZNr/mNgVVclheq6f4lg7
1YI9Mc0vuFnGHcT7gL7ihWUWurRk0dks4RlMrouOAh5Dr2p8xjtUKGntjYUHGWNJ
ygVG77n+qtpJyjSM6B91DrFgBnruV8QTcMf9rsy4bExajh2kdL79z3/bD1Iy8hbv
kBLFgdRunn2uwvWErkMFjn2anMHm9XRUKARqQCqQ/ryTt4QWWcwrV9GS55DotQT2
6mh1JC9IycO6dTuzIVXgBNkjT426HcoGzH5pL766Mvk5R4D5z75dUHhRvvBEKU/K
CkuDk70opgMP9s+RuqQmkbZbU+WvpIPDnUavFQu1WuYzUyiplWbXZA/o7WbHg6ZX
AEr0BqKcz5jNIE43sDsnEdXbDUKFzHGrVkkkARIR4jyIilDkfc537nSjxBIkFtpI
oOMjdQU7GXQkFbLPT2UmKiBazL6RNINMbkji13Ns3122PkQHTC+HeYKwvbftAnZE
mg+B0r/XpIOm2+kIFRkH3nhmDgwpvdU4XzjlvpAXn+ii+7u6507A5gotl+XJhL8H
dL+ey8J26VYVYg8gtn/t6HYAWU0dgwPCNsWghYF7lJVV5GVolzKgl237nLA28T8Y
BbQDdnquJgQrU7q5uU9qP0E/v7uhKLEkBgICDM7I53xO5OMgPbgB1Hjf6wEviPT6
wL7wIiPA7WrNg3LegSL7ukLtoe2LMGhao8ucBPIRFR4qOi4Ri3r6bAbFpk9rotc4
Nyj3SEeyAR7ajVLNosey8zD//x0DA9o2BdQn2vAGx7EQfyQe5Rt3yya8u9jV7TwM
ZSCvVuFrYJ1mRhWgWRpmWLqMTkjaEXQU86r28gAa4rfO3kEDmukbNYgXJwPo2p/1
eXVj0rjIqrsNAmTOzvbEEVKk+KRCRNMFJlCYwsUFFG/I21pvulgLB4ca0e3i1YZE
JVBZz5Ovoy9fqOoPh6Un3Si0CkGHx9W1S0m5bTcVaov7tA/Ja8i6vH2wB0E7Pviu
WmgHpNcXqzV8+jH9lxAmsRbQ6XVa/XRniG3eUYyhduHiMD4y3ydzxPU8esAta2XY
StzE32xs4L5JbId8JP7OVm7RvY42PtP4aWJEquBDWxCZKeppv2erCQJvx9FEmC6e
h6riL2tb+FaxFCIvYBgF3inl13PYNvCqSpOOPXbXJBHO4lTuWX11HeovqEOLDdC/
QxmhX+T/1IMZQe2zGPoQqmC1LI3vncy0yisD0JzA/mYjkTuA7A5jBeYYGpNuekGe
ImOhZhtfwvmsWuPJfjWPGky0GU/UCKyx0pzrnLN0bVM=
`protect END_PROTECTED
