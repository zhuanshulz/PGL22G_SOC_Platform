`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/c1PIe9pZFZz4ZUM6u5ijG6wKWgxD/MgfE0CuJnQSrCCPEBi+JF9YPBdDu6iSm3
mNMolHwQhMS/tEYsN3bYjPleA7onALrE3a6Y48wlUlEw2hR8MTu8bcgTtZW9KffJ
FdG0+88vCKMoTlxM76z6LeF1OLtNta7M7B6IRc8iP+4g9mjvfcXv0YnK64+6/EGV
A0gwzDIFqqi67palK4WJpN+/Dd20uTQuXkXaG4f8J1EHv89uBq6fz00L+miTAKrU
NUWvnfyMUY/Kzx3JY1a9Cv984hZV6QXZ3R63ukKaj3lmlWRkE4+vyE+7DW70iJGB
6eLIsaLTR0Uc1S6Wu9ptvg==
`protect END_PROTECTED
