`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YY0Xve11dWbOMMFuWGpGmL2wK5tbYxslo8kjqzPFtgScgxBgwkiJT1r2km4rstnW
jsD+jcgSb4mKTJjGw413WclVW26UFx93RE+t8qt8jwBt/sMnJRBvbHiSaJUpWdLI
M7+GfCzzqM4uhhQhnWS8F2dkrRhSmXf7z7OS4AM71Cww2nTYWPgEo1ptNZpFvQVa
ybMlZ94kzngoXgVzky9nxl8bsWuW1dAhp0yYRUOhXtxG0bRKkr2NPmmESPLhZnMD
dwkNwGi/j5RN23ktK/D30oSfAckU/4HwpvksUBVZbU9WgAyZ1DQDC4SmMBToNKCt
IgwRkw2m9xGIBrzNsT4IKzV5MxXjVPQtrqEq0tuNVREsO24pdQyfqzv8oWBFwqjR
RVVli1IEni1IPCy5eis1mmtUbzCqjS1fGWYjxD0NMfLr/3NrDIp510dOecDZppDE
9HjuThz7S62E2Q3Um/c2ygQM2qWmlRfOyclzyMLTJ1qrsuBlmOlIXVhIdFkf9PWa
WK92kuopNTXtYaR5IoDNkhIKi6mjNOr1Eu25WsrKkYH6AvgptLpFN5oefuLg+egd
ZVIfoLlwVaLUKxB6fr6bwlrgRUoCo8XxVc5HSoiMELxmdV9VNdGPod4k15V7JeMx
a41fQk+6LTS+QW6f+zS5SxIx//FKsUIUJfPsyBtF3xrk2GdZNpdFXfD6ZPI/q4JZ
ZYK8HBz3c3J+CBec1Nk8qOlZKGCIoEikOzH145T+oPt7DPa1MoE61a8erdWP4OHm
ymphcrkngyk94BfeopLJAWuRra09YoKVNsoPqp2LkWOFE7m1WF3iDGhVGqS9XEIS
p2JxGqdIn3GDJI8cagJHHxKB5v8ExX9VIX99skYLu0O1yZvuBZpwPzJLCC869oeY
V2bj5WqOo55kCzIa20A2bUImHRibCotkGKGWRlk/Vq8+HdFNLrU8UjpZwdNFri9k
CCebchvTNtBK/zdR7gbG9aeuVI1z7cdVCB0LBhIHIvmUnOS6NcFAkliBhR1J7KGv
uhXIxd5CgeIQZoDPbiMp01p7zZOJGnzijeyZwasIiriM2E/9XXLgrrnPMLYYzkov
hTnuX/RA5ResRXCP+jQolDYoDUxCPSME/v3cJAyBKYlAxXs0aRDoPqFZ7WSzywL2
46RpSgOtB7DCYEAmMLx9oV0i8w85TBrAk0sonV49OwQ5Kqa5xY8w35wRY3CJzsVs
K7seJsa66A0rfUrNWnZazclXZ5vMCPo5wx9Q6/dz0cPrgkPg4/geCesW19kVDgwY
Z2kxOcepKM3+cSiEmmNZxEuQTLKIMMBozJ8Ip1JGCNI+bbTzeWx01BbKTmBe612b
/OK0XF93pB5K82QJxaxx2UJZVt9mFCdQKxpO9z9rat0FH4Ox8p+/lBlwlxHDs2Bt
iGfVHT3shzlsQq0feJFg/5X3Q76h6MX/CtzjDGT1ayaGck6ONlmLCSvOCFbb5qox
CMLDpZK9Mmnptmny5paNYboMs3mA0aHLHki+LFHXUAu6sQpGc7/u+I6jCdPnGa9J
mmKm9EQY4Nu2hOgTmMcNATEwaCFmsquHHig7we2QGldkRRyxgZalRa8d3b28pDyQ
9MjtdKdU33kfayEVi3P98wJ3VomMhpBQqwkkrx/fidhG7nQ75uvEYqVEq/NT5Wpt
FLZgSrUxI00tXNEaJfi220M8N0t/2fQY8N9kzgkiY/s=
`protect END_PROTECTED
