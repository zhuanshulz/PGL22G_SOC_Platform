`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xfvdeHSeGYKCMHB99D+YPX/Xquigyo/SgMLrgpe+efNtJydCJ3FkNoMnDdj1avYL
fL5mJgvDVW2Y8+nOo/o/uc3QD5Jjs3mP503j6ptVZ0RM07GNtmnTlWX1bfPi7M0x
CuTjYtJAznwBAfL5wiVJgyaQa8JeZzT9P1q81GnHYck5ieg81Rxjurv0par8qy7k
Z8JL99LTdnaF9X1Sk07sIvBUBHnqlEaCYsFqFcgcbqcHJzSRaX+RDADo9dL5N/Rf
48Gvz23S4fxFW0HQtXHclGF1oQcdj3GyYp6/QhcOeplUVXbvHkluENVyvpba2UIa
MdSj4cJjuOgN3TysByVqBVfqSp42tSU4dwLJ7osu2HFR8koYiH8qNdGwoODoWq92
Wqhi5G8LmXtoHbCWlikYhsWCsF21lZ6+UBF1hmoju7zv5NcayJwKP0AMWIvUagzX
`protect END_PROTECTED
