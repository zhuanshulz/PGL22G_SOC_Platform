`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7araqI/dr6TFsifijyEGJXAfJyRY1HUDoppXceuk88/gnXCI+B+y1mIvGjM8ruY
4q8vjGe2+ND3LNyjQf8ADxtUzazykrXusDrtMYELNF83x5fXZSICinxH8srZpQrs
3eR/qc88mJuZmHvkeyL8NTPseHWhcPB5lyay0c8UmBv8E87zc2FC8nrKnTA5I4I6
/SbYS/JM1Rl/SJz9hb00+PCJGPKlLGkoXDuXHj/yKXZcvcJOqPKV/hbdooGqCwYj
7hO8jSuZHnh7kbY2lXuEMwxSaSE46NezkOsiQJW9ACfhIAVTKJgnQll8sw0y22vp
VfHru6YLz+ucDY0sE4tTMjjoWnaO1qCyKiGoKfK7/RcMYaFxeSjdiZibdau9//cl
m/AiCmMSwOGaI8Dfj+CkfTd5yv9Id77rfPeTrd4aefRYzzbyp8as1Db/slrbjrtw
uZyY6IamtfysF6oQXv6nWte3StgUrl9nrQWG2IiT/yOhbfQpWP9g8wTyP1jucuwr
7afxV4oGfBYrnA3I4H/5rG30EENmXOTA/j3ea4cm8R1eeB6X/OKf7eyF3fzEkbOg
yNov0ChfjIc9O5C8jJVPgaDLfZT5ktZ4k9DRb3z5RykYAHX3IUoaIG/u9zJX0ROb
QtknBi/3D11utQXUjR1dqYeCpaWcmRnr/0543Bu82+xkJU9kDVqB0vzi5CvVxzMS
kf9MRALBgn2s2nITv3o66diiV/gXjiq8o8ZvF+IkFK/0zkDmBrwaFFtxKZRmYl62
iQjtAOuZ+z74kkp+7nudiyb6AZkjfFOgjzz32VVfLy8KECK/HFyOd/lxk9fJnweo
Z+A5DZ3eT+X1osrE3+tpQE9J3VfluCexExMbQhtRIB7mI994pC/HwghgXtWa6Nli
aLko75U7yxO9StTjq8bTC58mJM9xB7G9+3qm2kzeh/A=
`protect END_PROTECTED
