`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nmcwoRzqmFFDIHa2axu2krkT7/56hrQtHaEL4E/06mR2ZcEAE8E8d023U0pmn9bt
AHsKxyK44BPtt6km4kovmCUEaO2LRCpHWJB1A9hSLZSeekrpwbkwabK9gyzU7+R7
Powyd+FnG+fQrI4GzYuYGzdU8c+UR9uBl4ZtoTgPvD7yV9dMjJonXKI7uSvoRZa1
LZ3lgjYikmJ0Tms+ISZITwAKISvzxxb4qXL5eQoi2uLhMFyTs7l5RHaRxzkTOWbD
ZwHj1rA2qT7KEMlTQfnARHh8LId6aruOtiBxkZ371YjfEZgDPpT9VCJSTt0mnU/t
A5Kv3LbAQ2jUldQD8gkdPykgsyeSm6NC/7VALseKarZKOdkefcxsobLbJzsQaamP
EwP00ibDhyGEn8sLJh+t6gFcw/tmx6UjPu46iQkI3oT/YXhJ7+YXIta03+bu70o2
igeyxEAttm9GtC507B9vMUxvSpkm410mi2BbwhTd6SWNqmoujg8EPxuhxWBfEyRz
zIg+cLf04xu+i9E2bwtBstAd4BBek3AzNtSyHfGqL+x2KvWm4azfHWni6L+YdwF0
BuroSvMiu5zYcCgVM7WfzQOW1gXJJSFmBy89U0xM5iPNUsxq+1OMhuQPsNt12eTV
Bd5Kb92/1UFdkISlAE8F4Ihf53qGVHWM2NcrK40XD04Oko+QnUCWZWIbn0pwNWRM
Pam1OUTFnkJI/ZuYE2K27dND4b6/h9WTuv52h+9JnK0=
`protect END_PROTECTED
