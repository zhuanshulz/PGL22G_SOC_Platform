library verilog;
use verilog.vl_types.all;
entity INT_PREADD_MULTADDACC is
    generic(
        GRS_EN          : string  := "FALSE";
        SYNC_RST        : string  := "FALSE";
        INREG_EN        : string  := "FALSE";
        PREREG_EN       : string  := "FALSE";
        PIPEREG_EN      : string  := "FALSE";
        SIB1_EN         : string  := "FALSE";
        SIC0_EN         : string  := "FALSE";
        SIC1_EN         : string  := "FALSE";
        ADDSUB_OP       : integer := 0;
        ACCUMADDSUB_OP  : integer := 0;
        DYN_OP_ADDSUB   : integer := 1;
        DYN_OP_ACC      : integer := 1;
        ASIZE           : integer := 18;
        BSIZE           : integer := 18;
        PSIZE           : integer := 64;
        PREADD_EN       : integer := 1;
        MASK            : vl_logic_vector;
        DYN_ACC_INIT    : integer := 0;
        ACC_INIT_VALUE  : vl_logic_vector;
        SC_PSE_A0       : vl_logic_vector;
        SC_PSE_A1       : vl_logic_vector;
        SC_PSE_B0       : vl_logic_vector;
        SC_PSE_B1       : vl_logic_vector;
        SC_PSE_C0       : vl_logic_vector;
        SC_PSE_C1       : vl_logic_vector
    );
    port(
        CE              : in     vl_logic;
        RST             : in     vl_logic;
        CLK             : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        A0              : in     vl_logic_vector;
        A1              : in     vl_logic_vector;
        B_SIGNED        : in     vl_logic;
        B0              : in     vl_logic_vector;
        B1              : in     vl_logic_vector;
        C_SIGNED        : in     vl_logic;
        C0              : in     vl_logic_vector;
        C1              : in     vl_logic_vector;
        PREADDSUB       : in     vl_logic_vector(1 downto 0);
        ACCUM_INIT      : in     vl_logic_vector;
        ADDSUB          : in     vl_logic;
        ACCUMADDSUB     : in     vl_logic;
        RELOAD          : in     vl_logic;
        P               : out    vl_logic_vector;
        OVER            : out    vl_logic;
        UNDER           : out    vl_logic;
        R               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of GRS_EN : constant is 1;
    attribute mti_svvh_generic_type of SYNC_RST : constant is 1;
    attribute mti_svvh_generic_type of INREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PREREG_EN : constant is 1;
    attribute mti_svvh_generic_type of PIPEREG_EN : constant is 1;
    attribute mti_svvh_generic_type of SIB1_EN : constant is 1;
    attribute mti_svvh_generic_type of SIC0_EN : constant is 1;
    attribute mti_svvh_generic_type of SIC1_EN : constant is 1;
    attribute mti_svvh_generic_type of ADDSUB_OP : constant is 1;
    attribute mti_svvh_generic_type of ACCUMADDSUB_OP : constant is 1;
    attribute mti_svvh_generic_type of DYN_OP_ADDSUB : constant is 1;
    attribute mti_svvh_generic_type of DYN_OP_ACC : constant is 1;
    attribute mti_svvh_generic_type of ASIZE : constant is 1;
    attribute mti_svvh_generic_type of BSIZE : constant is 1;
    attribute mti_svvh_generic_type of PSIZE : constant is 1;
    attribute mti_svvh_generic_type of PREADD_EN : constant is 2;
    attribute mti_svvh_generic_type of MASK : constant is 4;
    attribute mti_svvh_generic_type of DYN_ACC_INIT : constant is 1;
    attribute mti_svvh_generic_type of ACC_INIT_VALUE : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_A0 : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_A1 : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_B0 : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_B1 : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_C0 : constant is 4;
    attribute mti_svvh_generic_type of SC_PSE_C1 : constant is 4;
end INT_PREADD_MULTADDACC;
