`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M2YC+cDe1aORltAu/cBabSk33V/qExvKqJH12gRmTo50c7U18/1OsUs162B4eVvK
JAXUy/ELI9UJgSdA12b0J0xfaWaYXvW2tJopVXif3d3ujB5n9dMj5GOJm6at8mmt
9wq67pwsK07DIvOrSBMlukmgtEwpX5fVNVz+UoO7lThyAy8tl0vjqd4tNrUZRi0p
Hz5W6rOBY6ap9dyFDOjwI/ajkaiDICDMA1AVieYjnf6yPlSvxpnBMNylV+KGm9V+
w3qVxyL9dA+cUm+kyYE7AFT3iVMZBzXNkbDbDU+v8Cka8nsOQ3L44VfQxSqlvRc0
PmUnu11S/0mgrW/Xds8tVCDJbsFUMREBjWgU/OBRHXbEIvMiKdKO3+gduSouAxQU
hO9e4jXex+fzosbPyHXHhkU/0LjIVjvY6pNFXp3OrkJvLRrQpxpeM+niaUG5SoKC
/B08/5JoS5VhG56fCsweiYrBXeEM2Y94R2+Yx3MUvgvCC4VC9ZVwR31uoOn8uy7i
n6J3mseFwOfytMbAhLgwCpaaDByV5jHog9aVBXpMH9tFeS9+kPAXuvsNHC+yeNNn
JLnMeMrczAe2ZU3803j9h+lLPx3wqkvcLNfi1ljMzGHXphaTBlpx40Oinf/KnG4H
lWdSa+MRFfDWUsAUvVjdLw==
`protect END_PROTECTED
