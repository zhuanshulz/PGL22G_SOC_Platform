`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFzDImk9eZUJ+ya8Nl5kY0ZKel91BGfttu09xvYB3hWqEva7prwpVF9wxGZxau5+
I9y4hVkiuD3QEyz+DUxWmU9MRuiUwFTPVGleC69UC1Ure+dtSgjS3j909fVpTwzX
4KyvyzC9xiEnmcaHGq/9aNxR7Q0OgmCGcOiIU3FWXxBfI6yVa5inDe6v2rPS1voJ
snjCpqsP3lfVNDDWrIzj9+sfn/f3jQPtjgY0G/Xei+VVFOx3LbMYS+2/c4QryyyZ
U0JvVg8EuGosP31uUX3jcqudPUKcuBtgix2JwcWMop7ItjbGn1ZU6nSBu2O1N+Na
fvwq/dAEXmi4pk/2UzWZCJrhdXx6Fd8vDOWx+LcnHPco7F0sxZf59f2rYoDIPH6R
5m5GPUO4ZX5+sAP9ZTAxIH0HeHv+32AkbqYj5NzuMe26BsadgJf3GiuOyEKjKaRU
oo0//X9n3QJxPYGaBsG3qKFw7JCfvZYxDEOAqVFrGlPdUpvdzggQqhAH3P8EeMpA
ay7TqwnODcTslhUGoSee2Pn/z0+YbWnH3tmXVGWCYPl/1tIblhAyVlnW3pEd5u7c
2VlCNfipTUWBMJ5s86j0ckmYPcQ98pfqMYktR1PxXeHsv1jaRP+DLoFmGtsONQ4O
2USee+uPx0fDdM9kN3vkhhf0goQCbd4aeTjJtvZMArw8fnem+apGTa/CXf77raLz
eZ5Dbap7Q1bslPb0a/8EPBBe8LTckaou8MXVLAAHkRNgWNcvwKbvTAlWPXXRIQR/
WtjO5j8lIdX7Ws0hJnNqq67FHnKPjQxVqhdmqLI5THjx8+Dy1aKDh62eqHKP6SVI
9r4rBUJOaf8AJQv6ATW3dbAAO5gXOFNWwTUxXMNzgPSe/oZpKCtjxi7p5TG5AFZU
dw0SHz1lotRyq3lbvjnUiCBTUg0HWV43aqDP7C/Vu8mWzWCXnSf2UFXE98zZrHXP
8tfZlo/UzC8DRAqZbWn45SpAKqMGKBnMuQLbHZkOEBgP5xOar2MEjxGU4e1uOPoI
RU4C3+SvgdDUXxa3/Zbf/IUPR7TmFh24GtxjKlq0yC4DndYENh53bynUyCsDZEXd
0gbLIcUvEibJKTrKb+5Ruy/PRgcVfSHPAmL12nRXdemIitRZn9QSVzPNpq+nEnu3
Pqsh+NYp3Vt0u8Ku3/PAWgP8jfFd2N8uotu699vORdeaFbgOSLVjH5DnTxd9SmqR
2J0CdmCVLwcuXPGBF8r9Q8iT8a34NZKCc0fntwuBa569WtEpiPuKGP5hJcYdgVV7
4LT3jqkuZLcrxX+9h54CEFp4rP/M6VljJ5twSCczTvPeLpT4EktsxEUt6cDc03/l
Yk0zn5gydCXf++iIwkeqiGHjT44UlJzJaInbmXbFqJKFoa7jjjLw4U8jmhfYJfi6
ryp8GZlvXrKoIgOx4/sVF9n6bTuq8oV27M7z5z6UU1D1wN+u9BRKApWxN9Tb1s+K
nzTiek2NRHTpaSUVzUyi7lq+riW+3T+0MhYR8GdayBUFWqu4LUZg//Xt6n81ji73
qWU7X780XO8TM3snPChyH9cX00xoDmHBHC6b4+8ZJa4aShpwKgkm1MjO4NH3PQ/r
dlhU3o/PuGVng5n3sC7OfVMvXmVXLC57q23bjiBT3NUkUKgDr+MyyTapDXohmB0m
4RrLcEjejxtJbig2++QHu9FBHyY1sF4IcwDTAa/tqhX12JYF6sNxeDymd5SP5MLC
1tjH+HaHikyiRVDEdjr9C6ku41VFo81NwZyQFFgOv3YUoH9vC6yufEPtDj2ZeBNt
pzcx5tpUd5k1NiKvDbEk9whJn5WGiyrNSlOko76nOMFa5JRB2YEsLXK+fWR2bywr
yOXB8VIFcgIsHWXfQkRym2D7uKdnrqoWgWLO3umQ3xGQEVlft1L936CbNmTBMyg1
+4/z7jQ+0WKKeFpI/R57fyjCK8O+8A7iPYNso8A90M48OFpRjJh5yQiMIqXGU7HV
ym9KJZEMUj6Mkcax0ys24jswWeVNhHLxAbScL2LTRo9tW/6TYXQAwnERIYUgBM7Z
O8vBLYZfDYjOjLbf1SYex38kneh2cBToJkAiZBfzYl+fM8WFf+peY88MZwMaCvrz
03UY/kxEB5xlfF34ZpxG7WBMQ1npWT1+LWH1/w8OsGhQ60G4XBLJX1jW9KQl1k8Y
19HcCALp8dkt7eXjvA//eqpPB+y4Nkq11jzE0SCSvwIpAjpjKDhAHZ1FenNE/CP9
3DEMVze9N+t3DVDhk6ehBGuriVpvH4X/xSgTBtKd2lkFhU8gktVVOh9g05xNihgY
UPWGOpuDDOmlom8ASjXIOoLwqentd0ZTu1aaLsngyYkcRkDI42dgl80b/GBaqaC9
zusK4ArChAZ7Sh/2pnjopEBPGrfmN+76uuPGzhSlpCd7TfHPfXcvOKbCIHwr4wsD
FCHxEuTn4O2jM1X33om0Et8lpu/Q0HslKT+ZHpCwPADo0KDTK8zEnr8VFOXTCj8F
ZnCCDwNLaqLBcpI0OpADRAhpe3YIlKnWIFgCf+LZKCkRLzR1Iyn3w7f3reFAoxyp
4Xt07eFspVwM8D9S4+v61rcjccFR1hu1/GaXSrQHWkOnjY5xDBk1+xrvStVluN9y
lY09e88rbYroz5q0Xu/v+Wryo6FJA8rmIc0u0lT+qHT9jBj4Z+RmMQ1L7f9iOANy
ETkdhzRlgPzHW4ANjbmsW7wO7ZKyyC8KehA8KXG0IIpH0YN0sKAE39z4kmz9xd3x
x4LhRBSkLPVbey8k8M24iWvi+ZJDsH1B+Z7GPLHb1vYYmNRC49ezXDmTo6/IRHkh
iDREco27BfkwjaVfb1/b54kwCC1koYCPCDbXbS9QOgZVr/WJ4lraY1pr6tjAtVUQ
hmsgTTay8nzKLjhHiXrJRrVu6qk9QdXrnD/7ejaouZqM5LgIEzZID8loLe/q9xFU
dfM80ZNBUKYyzVWf+YmPl2MJ3kTTJvlZieZ6+G7qbmkb6tYxjX9Y1i0ebjBc+G8+
Ba2LUSWFC6D4z673LY9Pt68U7hXPeQigJK8cEf4b/5wI9VL1vRerSNeSd4RhjcCw
AQfFoUhyEOkLWQ0U71hB5urszk68uAUbHxLv65V6iuVHUWi0m/zUFX66osVd/nox
wKb+cNVAjE/HDgXJ9yYifuQHqQylICrUub1uDvwy4KKhvngVZl8/UM4D23UIPrG8
y3f0r/FxIRkigURGYRZbhPPNciMyMHGlRNw4lN9RQRFdG8bQXFKouNdUq+9qPOKu
vmsYs5ZFzCWHRnAtINdfgU6EGi9qt9rRGpRBG+Eeez0g9bxVquY6TcxpRIGKfn5U
T8SQDFY2EjA7Co87NyVlJmW8ji/ibtPE8BZuoGZ/LW7uXnGBP3kHptJHTFFnlnZn
8R4U77YnTDmPbPeG6eShCIaWbtCFqJLRvM0AfYO2x2W23ZvO37nVtAhxUAESvjDQ
gc6aqvV8dDHAVFvVOOI8wdkhMH1XC/iOIUM8a0quMOZTaa/tUvmvqFmiD5WBi2g2
5xe4UuwHcggb2m+cBDQoy1q3iIf31pI4uuzPuFxW83QYw/pn6I0Z34ZXgxVM8rf1
lCAPiyXAJE0cBQMbokWiUEB2EZnH6bDH7iAtWzQsmtf7UUKeir+XDAiRzP/FJtvh
QaXoA5G6DsgWjk7gwBEz4+oUmfXXAq0QxVFda6qp/0DCARkxBvXy1NxockD3Uy4e
mWyQsyEdxCRoP/ROvTEwNB5DMBek0XUX+SRGpPlhLQDCB7CheuEEdep66ApXP1hg
NAa5pYuYo2oHPSXhZeRpdypy50nLRexn+l2YBIm5K+vV0O0lFFvidE8jahkrs6qw
gLSr81snHzyOqi9S+Rj2QskT8SiUr5lUvb3wRJDh4eXFLopKAYHRM8ecuIYCXWBY
+MBxwCJr4nkqUCu+54jXmHIsoT9Z6Mnn76dqJA7ZH8iQve4vwemkkWaNlkuHZfqJ
Gh4i+WFBMFbhkJYdmToeHL7br7N1xVejXhv9eHq1WdnujkKelu2jY0VExRvDa5q7
`protect END_PROTECTED
