`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWD7rc/MctFjVg3+FUCLzhM6H/vYaBzl5c5rIqnFq/XUBU2cPJv3extqVbN7enc2
Q4Qg3pkx8TGbLVtdyqwEG4rZ0nBksFdNaIGswK+a9+ynhwWnLGlvBHA1qwQsOyA4
MFH8fbpE7SpEC9mtK8W5iDR2bm9/Tk86IVEtpfKs3AlcDwfeakBvs74gWM90v84N
r0li89c98nvRZA9sAe5Vj5Jk3FXgCVlHMq6AMWyAZ0pI73UF6b4tSsEBo1MvPo9Z
Aj/XEvkLMKD7+xCm/MgHTrqNQnQRsucM51esGu7LgsH70yKFthvLya5jN3pagrtq
NYTg2K155zPzLJaWeFxq6JKadXjq5uOCznYu9e+VkKI9BOwnDYs9/O7PncFXjtxF
sAysL0rRdN2+AuMhxjxR9BZtwdaAiZ8FzvwSJN5HG4rRN78c5z1s0Z7If2f7Cwmt
v2elXMqQn4S0uNScosvB1NtWlmpI5VJqgJDx3sUMJm+Kh089OuWsNSqGcWEdPJlE
2ogO6Dc+ZQRtAp0YQxplPI/LJxQqfV2ux+wq0IrxYEF85bar37NkplVDlHTt8B77
4B54N25KmAzI015gJthSU9v1IrO1SabQqEhhL3JgD/5P1+sdD2hpOHH2errHWi4y
H012rB4e6bO1LFkzCUQ+rBOMLXd0KAvU0rO8LAWnFnmM3mx42niWhjJM9jGxWoaR
rMo5aB5C7lBK/syOl8vwh3RDxPfoqg5zYHVAMYrpk7c+E61cGppe+HMsGpAqXMdx
pmtU9tU6YY1SAfIBATIBQpNGBZCdjq8oDIXIIhWy6jK44qIuLub+txe9Qpot6sVl
Z91ZSEWiBZmPc4TBQOR+rQGlBqlodVhN+WbYDgGlIxISj9HiyxEt7ZPwn9csHorF
zPrtyC13erOQMXK7a+odiFRavhNrR/9PC9WWLw4MMiaU8ayLnjoT9IoBbsobOdyr
MaVpXX+IfswAHktcKGc1FQ8mCKsPcHMbocjCa2KFC/DcmDiP+D4vIMXXq7ixm98K
LcOZTXDldDB78WBmlaPwM3T2Bds5oRX/2D/88WsGMcOTbrsNvn5IwL+6Yh4FJ+wt
UJs5NZ5t7yuBVhvRhhygudo7Wh8ZVNNNxfyRSXHqD/FUJFYxE904wnf9dEesSvZm
2I/6y/hbp34XM8kZX2faIAjzlq4Tmq0SjXkgv34OhJ4/LbupnCJWy7ZydBnTKu9V
Z2aeC6OlVIJ1osBHGHYTSyVMB7lBNSxiv6pOwP5o5NMQzGgIr8sVukenmyMmywfU
ds6b5iX4mmmzg+ytHjqYRcHQG2Azouh05vleJbcLFVm6E+F20lebgrYkksYEL15S
5TPZZHvD3NKs+LeX2RSTAMUq9HPnj5JLz5K8cKv2Uh0SqGSx99TaMvXlA9iqyALI
QquuHdABw+E51WlxT/kbjsHtrk4RYiLIKh93aGs0pp2wdNdgUgorCEjGItZNJVtu
yPk/nmxLN1gQDt1FvSqwd8dl4prxU6RnJ3iLwjRHzj7OYUj9i3QMJf3BqU7wygeA
VKRAzB9Mf9XcD3Nf9qFn1yUvgFyuF4ofogjn7+99EJ0rhgKJajxe53ymPiJ24UPH
1Nceozsqzf04UNIeHK9KGxROnaYvptMsu6I4Eh301pA5cC1ONa6ZtUGfUJ2u/xPi
W1Gl/VPawauOkxOK7WMQ8BpeCAofMne29qBkj88oL3mfg265LYYQtjl1INRfKCLW
NsCfAOcPvcjjt5kLmHwOe7p3Xv7aoQWQDjOq8PUW686LvKJPRXBzDVqZK/M6BdUn
hnGZXRsRMZHAjgJCNYd277pkKZK8JVOU49ZUSmImeyyOSF3KfJy5/mWbFEQOi3lQ
Vo2e4AM6EzkKVRhO0PmKw2GQbxFHAC9o44nT9hAgYmUOYwZNCP/UuIQyCufzmBSQ
Pod4lvRj8Bd6O4TuZO0AHOxnSvCNMmV9uJlI8XZXyOF0K0TMBZAUb97+ZfCnF28s
eyL+/PHWZwG/o4DDPsXDxGepZah8h7z3iYWQocQtHlerKkZ5fCR2n5k9AuSJM3OD
uDkUaYeHAz43BP7dW41GthrSQ4rTYmu+zRStsnt8VNZhUAlBgGBAERtbJ0zeopSX
2Mo1DoK7Hnh/6zNpCc5/VgEvWIHIxriepLHi1S5ecanUwB586J1MamyVXAhgNfj8
OfseGlq284j1Dhr4Xi1kfdlswSTxbsF1Mp57Q3cKa6GAto3DK7+NuN3VrTPtvcvE
wIWr1AdNtA+Hh9/fiZTqZa4va9USZHJa3m/VUoUOLzd2fZ1ZjGFsTi0mTLKZnyX1
soAID/R0nh2WKgyTc29ipS0+wi3xt3y0uB+eUKm+JirwkeMD0gkNDli4Dj6n+Hkx
L97/t8Y4DmkiLwzDjC9Evk7VfIOxz8XWhxie96UpOBlVcCaV0+ugMcFDSEExV1lA
FTGBOkZVNi3tg2NpCK6VAYvsf2vJNMwETK4Y/NNYp20dTABRxdgdMul8c9SFJlTK
U58aEl/noha1B9HuwcMKsSP/4H9u91HZlvG7montFCTtTsElxuqyaoleysFUIrx6
pXMRjBY8OZVSXjSx4SJM30JZRDUnD+EMz04rB0YPLzLNwQ33dhCvwcXtwXriJ3Y7
TIMs5GRiVL3XdJcdsqrTBowVEGbfPxxWNH1t98QPIzHDR7nxx7QKWI/hTgR+lhSs
YIt9jWZVShu3kyzPEAu6dfdqCiTZU/uGqTl8cD70OXNYIk0B3nqhD2gwob3PN/hg
MwerDLV3mjM2vjFL28iB/KtIrJyW8LdGnyvjjXs23OAeW5FN1XS7vWML45snWu0B
bJH5ovCSdLzz81wIZlaT66/6GVTeeXkAH+6KUKu5igO5IvMxPEt6Tjd8IYduFNW7
iiFVjO/YAQtEmIFRZH/tijhmHHNdkDAdV6VkJikoOileO++janWu2hwjpaJxBZRF
/TIVj6KnFRH9qQrexNesmFC6D56je+/zKil4N6MkRe3pLUg4qJz1rUpsMnOsZ4Lh
hBENnvje9bdYclyJcCp3zK1kTyCOMx/cwj2rBcSnLhZFPNC4sO6qio+CUiv0kM7s
rY4IMNX0fRKx7T0cYvvgDBe5XWOk6Xpg0WNyIiTVwSJb/nNIZSNZjXyOriuEACT6
SxGmVGT1Y0ZvttlDQOmiL/a4PvHIWzrbyoV4Rx8/ZDeFTqQNg323iXPmOZKuqO5S
ohsBzSFqZeIB8D1UzDX8UkG+NXb/5X7xGCUu8FGxhXBtsiaWalj9BqCoY4ZZxOqQ
du1965wfoyqz4+fxW5BvJDetPTphTW5cwrF/UVrCwdhbgtDG4uLYKW74kxYa+2nA
7Yu4e3w3/fiQetAQTnX9ecqDeddnCavDpxOkhGfYpkqnI/5hDOmSDA6KOPFTHnto
CHpsUeKyqQBIcm99tINLwOzZX1lmfqq+/HV9EzTwck/qvkVPlncOUaTjrDvo+Bf2
YVzX4/Dy6mndudHUIF4jTF3+rBa9oJr+a+2oGovsHgo6GfHdOsJfalcq88zW1h9U
4EsTJPdmPY9w9b06yiCTkrZlELlBfxKpw4n4+o1aUWbmGu4zoNj4bzbzmSX2djKb
NS+HTF/0CFSauqwl1NkmicVcEdLAZ5SriqcaLv6Ui5AtprL2B31SgeT09Alp2Jas
6xGvIKT+XP/2/wO471ytRIFJHr8Lx5Gr0+1p8wZt5TZ4ND3k0yqWEOokdzqFg1px
Oo20bOaib1zNnGTucMOXlPH9nUHsL8pEkp9pBZ0cqRnWLz1tHGDskxbe48NSKvof
sgEJmjuQD2KWNwi+Bbi93o/+KTQ+ra7K+sDFys+f3jaW2uheBytDkaGp+jFQpNow
W8pHt+aHfptZb6lsos9YMdgWDtg/7v5QF5fJvB3D0nXixGA0xp6qZl22YqWuqQWz
mBqkS60sxLdKj35pA2fZedaEnBPQPDHJnGh6N8umlzv47r9okJSUQ93kSkFSvTSv
oA/11+5omlfJhmPuBQZ5OVihy//sx0mAixhlw43y+H8SLlLLf1nO83TAIf5JKRLb
4LBNC8nayXrTnYawVPzW4nVkz1iIw/nca92OgTOTkSqNRYGRiTAxo2WlHCqSHmzj
Y88yQFAnbkvmYhT6vXpbeKlGjFGVJj3RC5ajtsQZuDpPaWTmaPYpBCAz5PZXYuj7
0xhN1KHo+aPYdlF1mG+6Rj10lnoqOrCFG7/0dIX2UoOH/z17J2nOiKrbUXPsC5zW
U9HzzjVskLLGezOPrwieBpB4EvWr4EM8nPEoE8nLA6tX4QPYzkCMU2HBZ0afd9aQ
XcVoVqdNfoiv6NVTN+bNjN0gTg9cGmH6bjvs1Di5rSxkX6rjmm3A0J3f4d/gkIQB
AzVoJ5dk9m4bMfn4pF4rvP3mib1r2j0HeSS7jbb6u6lxGfXOJnCMaoJ1mdsngkro
x0GgofHPmfWvssesRNsmU3jEDoKBozW51ZxZVrprdmj31zNDnVIztl5lNXxCPl+o
pTM+7vKAEhFS8qrsC56p6tPayte+kxinbhi6kq2JDFH0eiXtC+lj9GuLvAl1QT3w
UbKNYx/OfAihg53oE8E0/cIuotC7hAWr6tAnmv5ozmmsdmNf2JVSKXu2q7vYEioq
ksqXeHEDwwLwCR1GjD+R0vFkWC9O0hxM3QxG9Gcqq+nLNLfq6eTclsCOawI/i8cJ
xPpJ7utc0TMNdvMFUTsA7RjFyy2Ar5GBZ8WYUkdeseMgV6zgfdDiLYLyE4jcOFjU
c0esEDv0eCQ1r09nZVy3Hkf9ltpBQfN6ilQfblOO8wihFm8i+Y9q57dKcxLZQTSp
SdY0YoaP86O7AQan+EjW/IXEVAS68FGXRTBl/YhwrxRUKAuVATvKHejbhbN9fyiu
0z5dk19BN9L7bMwPeVvsoWVxqnwaLP4zcsaWKOzmT3hQa7j2m/5duqp4+XdCxMJO
OZpnO039RC4dr16xH4KwNzRsvG48FcJ9dBPz3IfUWvOVixiyqXERXoNObZd67NNg
QQ+xTayCbPqOYgozwEiq1+k3tefjIITPZmOGqb1RabMQx0g6YaOSHqti44ua65lg
6blFcxMsoApXahmkQHzn2Bgkib/VkzlYiszNr1dx0/4VGhI9IdIGBkYKcZVtnpuR
zYgBcUa89MEvfin3ECtkXrTbDtGRinYRMegYgG65uESGQGB3DtwFhH143BkGWe8E
nv6eoadqCXxRHxmH+Kj/QGMoDv6OPpWTps8iWkMV44O0gXsOWa2nGeBM5C9PeF73
Cp7aGXVwo70MgE9DKfcvl0n01jbCb5a2OpXSREMx3xsQ/wG4lmOd2mRHBxVjquxm
ddN9uccn+/I3R5j5McAlY5TRkwm5kTEUp/bJAr7yq7xxcNwBwBTgsicSPzy+tIQj
chFx8igObcQNHviz+XrIMSEB9GS8ZH7qvK1zI/3YJBAEQ+BxCIPRxB9GNPh1WShO
5zb32DMgZR+zEfOLErJVsbwDyq8kfOKmU/szqaBuY5+yp67dccuRFvnN9JJUKPZn
5Wb4Ixa2UhKLcV8oAjkC2WX78BxO8pSybGwaJMn4iVIXV6mYNgnH+Ujg+JgHcVFS
/S0h8O363/J6RoeQC7f44mUa7FMLPhqn8wBJtuepXonTipon127/iw0EKx9xcIlv
+0jCsLU5CNYt5Sc3qZwAWryhkhByFc4vsiisPyiQdlYU++5yFPSN80xNJBc6zeeB
5FtuVp3K1pxW6pZVV8xQg7LTZaiO0aNFzpCQ5jmUgjVb5lgeJIdQwwojfcEAJ0Kl
NVi6JNXM+jgCV4F8FFaKxAfCKhGdzX3C4qriOM+6kotPdEHynUWMrjDQNO55zP2o
1tSGui8HF8VqC4wHXVKD+kq/zV+ojl7uUUUMDoj+FVad5thN/KJEsZZlHjRPfUgZ
uR9CDg6rL+Xvoo1PZWelqdCHCRU/NagBF+X/lrJ5qSeVKUX5ffC3OGmqiQtxPb0q
CfUSyWVEOj6RFs0WoDS8pm7SptUWYXSYDDAqfoAxg5qbZPrzGIKflK7QsRslqxnX
xP/aQFSJUQNrh1XzqLiU4fW9Z5VFreygyy6OtWeurnXnduVrZwnFTPiB+89vg3Tf
W8XmIR9FtNFODwxXKIR4vRdEQSEUqp8BcX8jPiOMXvuqHSTXzYo8307gerWQD6my
i3Esxa2KeajybBtZ5CwSwxCCZb/wf1PgMfBWRSrKjFqCc0wZvOgvhR1cyiW5EDw6
ZmjRV8C+XaKg8OxQJ1qmWgwzdIzHu+PhF/yrCSkDPgB33TKxnA4HJtkK0LB+cLIA
vrpRkE0hH2PsHx61RGxP+p7h8rHGZIPQMlYn+Ivbqs+0VgJSeELWw9pSIwQ/TLP+
CQY97sMOZRSLGA7uLKWFRGQkB7/kz1gbsrH26idGvtU4O+8xCXRx7yEN75OiYXRp
fDU3kRb0RIcphQHKgQNWHnD/EM1cm6dsnysS3PBUVnuJ6CU+PdPbIGF04izsAA7t
WgQ6iJhpmSxr67zcDE402Jo6iS04fyE2NBSgyCYISUVcENjnr1Ab0iTuG8WNUePv
o+klsnBQjSZHG4J8z36R6Rh5chQEqzoSrSaIBTrr3sxq5TZB01BwDsFGMG1qhHz1
O+ZpfSLOnC48vtu4gSXSVju8wnE2cZNuPO14UjDAz/FEtlEbv+NeaXpRGXD9coe9
PX18+5hijc+nmH+yWJ9LuAoJujexgVRMJs+xKWouKD1bAsyUO8oZWX4JSwI7sZgf
VDkjbjFL7vMMBzHRlcpG704VKcgbufsDbnkLumFhL7JJVtkSdk64PRtM2h+26Lwc
VrjrL/7W6qS3TBa36+UCfjmpvvIdbbRpnmsa4A8m/SY8SzXMceaUMGQgwsGJDOPm
PZEM6wLES9c0JippEwxDIQAK0haGbu9yzI6Erj1Rz0fD13ITHNFQPY8QCTaGyskQ
E5lxjq7Auw40TFceYq7OZDq3nF5K+mZabSeSigJeACpKP5Xn6oYJuNZX2sFtdwUa
/MfqVXmHVDe3/epP2m6CcHa9EP1pWayUTPKhwG/gIMU+QQq0ZsdlB26ICY5Fkw8X
xByL+HNDn2G6DDX64EwN38ADh6ywYYvJxoW+cJ6Hb0DakZasQV0fyBlFIbfRIf2H
B84nhaNSMrR8gF97MaKDr9i49izJHEsce/maMM2rjEdzHcBkDxR0BAZ+t6tUqaP3
G/IRqTsSx249ywJlliVHscOu/8qucYoF+usyxwz7qwV0sY6W8L3GAh0RTggqFYqF
43Jz2K9E334dldloy5BnN3p+EDbmf71ahO+cSTuHYkH+kFIQ2r/IPAJ9vl2MzZ2Z
D3zQMC1HwAiXxnvPZkLtVQdRfi3QzOEQl/NZ40Q85Db35HMZAaEWCe/5xMLLaYy0
iYHEHFeEyEQSEwbNAWAC1SpRytFuhTLuBt4q3gStwkfkoFTtSdBqDihFKGYG2cS5
wNGi9he004n8vSWnYo2I/D+LYDAimRapfhWYn/Ol+G3vnCEAR/46dyKSzsVBSKtj
ZMX3i25is2nAm0rGDGLsu3qR3GoPJLDR7IhmMlKz0lnZ9uTEVXf9ukELLn7FwQiO
HL6cYgOcM3JjBgzGwuQHAg2cyQvCiZaxppwFcHTzShVg7ahLCWc4CBTyXHeUKKNY
kZuhlcmk6MSCvKdZPaxXSPz/8e5HQ3iWRjVaWAmOf1cvQzKmoNVRrn5/OfGgWhUl
wI0KdCB0eSXbT9tJ3NMdal1TuHX2WXXgnUWkdzTFv3VrNps3CZUuUIM6UxFh1LGa
PPTQ84XbI14kBnqMEhhxpEKS9VNt3oAcx0ytnwD99PIAsfIHOwKiTTMk+C5NOfZv
OKCdEW5hYfBlQndJPJZ+8/kKZ9L9wg/xEGC2UeBce+obX4SrQ/08pDjQrvhEQQ4R
t2Dtfe1dm0qvuA0gxbs5d1GrVRYJTHgaHwEo/lXI0q9dUFvv15Q9QrKlPd5x9Ov1
7qImogz8+6y9EKl6lx2W1AUlRvghe69+d/b1Iw7XsdqPreuAW45xzWulw9rG11+y
1d0lusX3C1zUTrGZeIKV2tSBL04MR3KGNKSO2IiRy7SQnEYz679MxR9+zpt3dBs/
PzUoi5b8DnX0XfMYlxZ7FCoFKIyV+VEQQal33814pjMHok52MwqIp1fd94ae6wm6
xz9dY0ao2tHXiJNdJlFW+zIPM6ahgtGW/7vOqS1mo8zbxfuta69khpGeFj8bRtWO
tqSqG1nxhQGR16o8nran5HvzyaOhWwqmP9hWha7mgwyKbn9HG9sewBf7rnjWyXnS
6ZlDWsjeqIJGqZR7MWcLPXgzyr33jXtimav3qWVEwAqAR3DpOjZN9w0168APs4G2
aEW/48VvTPyL7DL3smXfASudVUZFvW2EWnPgJyzYVCx6GVf5xUeBTyU5X5wpID0d
KfNaDlOSicrzZleN7RnXzMtsiyx5pNjrnKGkHUVhYRdXeknPsAWUUryJgJWSTLQ2
xMB4Mpwkw4kWlXrz8fDgTvgnvBOjdQY9xcdQ8BC9M8GDZWp3Rikmqt1/k+2O0nT2
4zvzep2b0fTqirI9LDAcTUzfpg8W+BP44c/oT9/6HV3E0oCYY87SmUaqkiV4xyhh
MD4RJzMaIGFQIlKZ4zafE5gOkhUFOAGdt4NE8tprV0Y52TpqYzeTZzWMemTZp+cK
u4XalU7xxrAnuxZFxLh1z4hQAT2e+5ED1i21kL9+LbFzAVhm+GxGddbW3E0tT27+
hTNRk430cfKeQ0G1G4ZGCkmxMDq6quyV5uOeiLbzQysuxWFaAqqgrdRYqL1U1oH/
3gfTDJkrD6C0O3wUfOJDdxjYmo6h4RZ/NWhmx18BEEn6jdachXWRLLZ1owKLl+j+
F7uySmdZkl1hBeke6RF0JGjS+KG/xL1wvm7TmEfLJEp2rrUM/JMXWN+fzY6gvn5M
d9l5Zv5jJFF3xWqh1/E3Ahqdvh0lubbU0WpBL2CTG+Tgf2tGHLEdx8Xzo1ISdnRq
I+t+QqtPjv/CcjQLAFnjSOTeRjvrhuBKYmxF1LQp+Od28v37bvSLzwhdeqS55QZR
To2V44GkbMYm1v2TcbNr3yLTF/b7PImyrKKOEL/zBUsvrOjhKdNRZTGOEl04xkUV
YTrOFEijvvAOu+ZX0HT7z/NIKHDhBQE9EW2hj1AvVMWSwwTp9WtSwmFLjigJlb8z
rCYd9h1sV3RvA/sVVI8Ujl0rOvb/j7iTC2qGfkcmm1+K3eGQ8Ci9tsneR2Y5xNYV
TBUNf3qXNNtZpNZKI38a4FPoNJKa/+pbCTujZ6VBskEHnwwXTDRQis5uil15gbOS
fpTjLS8LlId5mDXCS7me8TEAX1nqoB/0lo1uL+iMilV2bF4EMUGhDseIv0Xlta66
iSfkBLXr0+hcnn8OrQpN5x81EWx7w0GyXO3+2aPf4y7EqlkDsUL95VRzamRGPB9o
z8lN0F4Vz7yD0IkCPl10n447UUdedLDpixe3vfs8mKRAwWeGi4a5iY04OqSU3wc3
QpBs1UllrvvP92kBfLUj/fJpq6KhgJJB52BmhOawoYhNcAxQUfHq9jJtz+YogrUO
fE1O9sylu9qOlULXIowThlCmfaQGBZ0AlbIfET4LyJxrwQ+WHooFsCZTwnHNibKK
52FbQuM/Jy5AGm7rOy0MI4UIFMRRJZuT+qZjTp4myoi79SoAO8V61pxa4uJTT/9f
yn0wekLqaslk+L6acgn2GQcJiDsiOyEigc10pty75RUs63pQjxHcY6Zlb5LrkjmY
khAtQsvpqInqL1bU053gitNe4EBz3SWYyH4jUNXXhOT0ApvxEn/gELEeT3Om4KWR
elNFY/K2tz1aBjL/amrgoY/8XgHVKCdTUcsTMLY5Rde1rfe6c/d+jLmTdULORMfS
s9rpC3aTKD6Ol4tv7fDm19zGK5c5cJEkuvXfsFvp5z+I6jBV1ksPycL1Y/h76qvQ
m1Nx3IqbbijRvf8SiDDleKqko7vvJVyuPeW2a39dn0lBYPf7fsRQtJ3Zgr9F7/wM
jmgnQRQPVl4VH33RmhJl/wlZVa4ViNwwgzz7qyRpkPUNt43m8fNW/pcDTO9cZ1Xb
wqMY5fedJChJbiRIHdTVFH3rtC3uGqev5yRNMJD6kLRGjrTbjARfpo1tka7TM6no
L+gCjoZYTcMkW1ewZKxKLJ2QakFV9qn0S0ft6uJqqrX8cStSXPLBTtr6wm64FoHB
HSlmYbFcSjioGMnvi/YuQ0DL4c0CYYOa+SR+LHpNoGibflmRcMWjQj390+v7wox9
onvp7Ia9+D5JHzg6t30bM+X2PMH9ntgpv7OYmHQ5BIrpvurF0gwrKfbuHyJRCBm0
`protect END_PROTECTED
