`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4/8fVJazQIk0K6YazpQcu7Yi/iLMkhJ78G4h5dboeKfoodH3pb5l2o5KdTnYVMAu
WMCHUbhfYmDSUKhcyzO+ytHuLTzAP5BeREHaB/5xNOGxuLkZg98ZkE+t/g727RgN
lyhbaCOGYVOL/eMolAJMOby8NVS3+cy8sZSQ2YOitunkpAv94BRgVcNRINphDULT
5lhkA8Bcrs4uh7qYvKGzRz2GMloyTJdtTwI18hLKmBdoxNXInZtJ9LgpRPEnzy+b
MlOuCAEayIrNEJBZbZfF1j8dFRjOnPL5v4lInGQOXQoT5HbDYiZEy9P71818XBsZ
HmrZ1+9EYPuGy3AVMvOejgRsqi9tWK7D/OzHc8e3KqqcuhjeGNq+Gg6MdjIeVPuc
MlukZrLnjBq/zlCmXihAdt7SJvBSIaOTohnLjXdlCzrkWMI8yT1EOb0HlqiIibIC
wtFFCZjYdMsvwSC6JuBhiFQs+2bl2prkh4nAB1kb6tbexBxp9dZTdrUBY37BF/rb
uYyVyV7c+FnygejQf/szTuEI4RbjPM4F47O86SUkFb0+AuRY5eDdn5iJcmc3c5xc
p+XEX3T9ecK3xegEopTx5TR6v2E1a+pjQFeECzqyCMOiH8UwpDF0pHSlh1hDtpvw
I6I5nhW/GOPVWO3o0UbAs7Z7bZKWgbYcFtsZHakXiXKmgInBI0nz+YEvk8i8M70A
aE7aGRiB+lwSjIQDMfObSrLomfSLGGMv6XDty54w68jDAF2NvaQ/mKxMEwHL0R/y
EGzQyq1jhOroDUabOeJ8ka5QT9gQO6mLHbiz8AtDNXtgawMfiS4QHSKhdpd5GwOE
XlXPo1Yry1FxNNFTlHFEVd5sB0hWiAD3L3l8txlQB7p7Kp3Rt+j2gZ7b1TCUdELA
h4ErkiVNhooPWMFd8zCHtfWWtlisQevt06u0uDCbwKJnh8dbzbaT/4Qa2tCRfxcB
EgFiNuyDEELfwObvpM6wfZKGrwPicE/w3gCDR11PnDzeR3N82HC9+07Pcu6YAVXP
Xcp5Pd8SPC8+wXsVBHHkp3jAoVj9NyTAv2pIWRhxJB8CvvBmBXJo07NZ/FmjsEem
V9iB+MgsJp9bBtcTGiAOxBLMhwZr4AmIePAIGiQj/buPS3QZ8hQR42fid1LX4N3/
M+jtsmmyT/tCH9/apMhs2kNUro+O6CEfiKpuzjjmPFcuEd7hMUjIT5q8K8t2MzW5
LJddqv7Cab87x2cwefa6cLvQrF73gsed1JJeToa/K66+rivY5w1ZAgDuVJV4p7CC
2MrjPbrqJeWzyQSnXoc5LPgreiS9MIRcefXos/bmYHCzTYLWt0AeA5FPqb+7wLWl
l0LuoEVhDcRBa1QwPbaYhmVBlmis31wO1lCrAW1PHyoLDQK9MhLNUtiI52z+EJ+X
TVejwcbcg3SVIoza6bY6HnnFpXEjLGcqHDeEZg7iSkxh1M1dHt4ElGlh8Ps/DzcH
vAZ3IbOnWt5JZpgSMs/fXtubYaYeeZUWupAJ5VCGQl/SCyW18MExIgudQMevLuIT
348UeknycI/I1u34BezB2ZkI+AE2D2IxA7OHzlWIG9XU+mltTH83RS/xgSvICIWf
zhh6kuw3aDlAjvpAq76GldXklQrRuN+cwHBtl+I0ycMUOH/jjidPcJ7WaxosNf3B
0+xLJ8liWUqVzZFtVGf4qxskOD29rudLdbdydOyCTKGxbqLAyZBZo5zuDalLMfzz
7PvKEkT8YoEeYkmiQXLY/LYcK7Xz5Fid2eOMI2Xegt1GavvQgwcg553+2RZi/REa
fkIPSirOldGTaPvBEPgN364//fV2BBr3EHAhF+ahE+UpzRk2l+hKlEsGfrDB4/vw
isNwsJUGZApiPKzqsKJm1IIfFav8hs4mcrjjaZyfXpCGH9xQeOZXPe7Oc6268EI1
YzFPv1tSnQfwp6y3T8dHDPiLdZnJOqz7HQRSRc8s9Gux4fLCugaZ5M5KYGUG6TBT
do3wI+GbvJND5C826UwzY2jcWDNg5B4KkmQN3mVL7MTd9GZjIGtQ1FrPEtCsq8Sq
wMHeD3HS6/5/bbAXqe8OoKtJqNxuX3OY8j27knzhHqNzrCvAcvIaqsnLdozbW5dV
B6IcXaysIyhz58nsx3mQRCMQ9XEuNjo8OvP5PtmrwkVlu71581eyQzjgjlN1hXnA
tb/8+SgvHPSa0PYv0YQ0xAotGEc92KqVipEvVzpL5PDsnpv7shfyb8oGDFpKKM3F
7fPzxHuj1uL6L/rVDcwboIOvqFx3pIxBi94clENxUmH31lAOWxPnjYh0DJ5m02gr
N+7v0epaKjHcxQe/1karEbnX9GUTEm4fNMgC6/LaAMJJxvVFAMYBFk4p28JsDKni
OzEly8BlGHFrf8I5uB58LmdLb8wX1qLSrGIc+QauFcq4A4pMbR7sVal0nF91v69s
k34uwwiin7PmXlDKxYm+11/f1P0+3s0WGXP8jFdAbIfRJfkWeXkcMcvpFXjmLKga
`protect END_PROTECTED
