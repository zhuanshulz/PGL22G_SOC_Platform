`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
40MYWzqj0lh0uRwRDJNgmjZVXolhyVlWJ1/K3xvGOOiqNd4mUP3VMsttvp49ltBl
MpM5Jofm1g3h28j+7M+60VYutFzf6Aidc+uWaJCXon1s9PKtA4fq6cFzJZ+nVQG3
rR98P4ztGhoT729KRgxTA09jfB+vKskDjeZV2x/qJNJkKZpqtnqp47qdettC/RST
iMNRIWTryF+ZZWm2YkhP8jdtMMD0Guiddk8AR1d235a+FQrEz3r1jhS3mTBwjP33
c29ytag1dGpTxeFtxiiOnsTZ9NbnM7EKAbA8rDFMS1v9Sf1wBx1iCzeTlSemGp1Q
fN/F4aOMztbWvELvXnjFEbp0u4CdcQPYOOD3tTgSMCyJZJdNSkQoU/HG3o+CgY+a
ZQS436yICCIRqKnTCA2pwHjRlbJrWtOyhv9a5d6IkjNDKcxtYF5kLWS93O8UverS
ToMzFLyxDy6UthSD+NIFqDpfA3WKxdrC5n2tKpu3bHMgE08yAJ1qtz4Y1lkgLCxL
cPdwlCyVgHPPB3YNP+R/PuKUznCJNmzpl6ZCBEQoN+kqxdGhvOvPl9PciVwndAN9
xE/zG6c6h1mKj3hoEniaE1xY1ATeZRB9jHPn74r9rVJSPzYO50+im9GFM6liJGSV
N967I2/oe+ZUm+53V4RaP2W/Ru7JRO8gNrzn5jS0em9O4eRbNlxLfQ7BEFCyIIE6
7YSMyfxBke3Io/5ysgJKEZN4zOfBHSPqcfFEYqoeHA/IrBGIgw+CSbV+FikrOQBW
+0NCOsb8dm9ef62fKi34vi5p8prz3ynZyHzHud4hsI0gOewwuirQn1BIqr4eEfnc
lvxOM66gRGHrXCMjnQf56E2AKbYcKgtXLaXS3L8T4hzPU9lxsT1xlgXOKS6WiS7q
MBAdAHq1d9fNCB+hE63gEXXkVUx/EiFD+s/0U6cOwhAXRtSHzubueAEkIIFKASV8
59WuktoAcmCXQrbKdxaKBciVKldiHL8+qO67j8NCBwSqgpR6qsjKBX+lyto+6gIy
sPOcwEHvVTl2hDk2Po/QSID5PnRjRukUQvM+FFAyYGjjbIuegp4bgJBK25rZtLlh
7ITzygsp+zFwKNuin21H/L1XthA7gLajO+ogX71EaddFtN3c8urS3t+C7jPZ77DZ
p6ckmOTYllceummFNE7kRGCO+NF5D8I/LYA71z99sDsxWituWJSHfmKLxEtUml5Q
nZTlueuIiL91b1srwNGDgaQWx7htS1h5E00zCmlaYf23NgUXLZs7DPJs7as5S+7N
Kyxm+f9onN8kKV7pB+Izi03iL+5UFMxumdcVBfCv9EyLrkz7UmaXInfbP+EIyZ4t
H1PTHY+mECzu+/8GMrWKNNGa5w+IQE0oNMVoDOA6snX4EVvO/LWMugoLU6ho6WvG
GDbinhjjTQhL3sOs+EwYGjHlaYia/0BjJ64D+Sjtm4b1aZO2VlzZ6TtLBRInLd8d
U+ImXYSH1T4kqS+oWmc30gjorpK0GyIzL27/Po00SUFYF3fcdYrNCxTHkDLsHeiX
FE5m8nF/LfcJ11rQlJRtunZjpaAelNwdOOmffC+AqF+z+E6isCYEET5goOlNOPCb
/SBVYwMlSqOi20jDaRvDSXkM9+9kxATkfTDmDLbqCX0OFU8wukMINDIUxBCRt79h
8NbJGZxLCuL9z1GktQlyc064RKPovuQAtG3n/etW9y+8f4XwzzxxRNI0M0syNVsQ
el9lonR1lXYo9t4nws5BQD/6pDG9b01LhOfCe9sWft+O//k43zZIh7YB1nBa6J1O
EZ130vckwJ/8IgJSKUUq96PK+py3FMROalMf0l3Fsl2bpbnemuF08XPNl7XrJi2N
v53gpJlY/tT5vCQYqveqnYwfynOrLGN8bCAxP4EREKVFJBUtrE9l1LsvESCj/a+X
N+BWmNf5XFGPXhd/Epl5Ydj8iWHM2i0ViSOG6nMF+F6eg7IER+Ng0KWxm7Uub7LS
RmvPT8bcnEG8U5bz84dvXXS9O4Qo+s7B5KEeXo6m1xtQP1vf6bnS6GTBhDrMOxtR
LvQggSDVHyCtFnU9w/i89OHsZCLhMjtSKNzCd4Z6G1s6DNkq0TBnHK0J5Y0pwKsR
o7vVopzp8lWyeMcKwZjvrVEQP3WyPwu+BTyYg2I4BgnHPiSd8av4H4iAFVCbsaOs
NmJju+MSHDU9YmT/3Ttd0NvafxScyM7Ybxz2yz3oRDtmkkJgJOx69mBvk3DPcAtS
yB+C7D7gYbgReMmAxbOAuFWce/JWfKcHQx6cEY8N0/kTkVzIbKMtpirvmoCZxnxf
d/NmmaNkI3lyCeesPTGfvxyKyYJPTF0OPK+n+fMeB4rnO6W8eQZc9Wy5vtCTQtO6
DrTraZiALBES1/8w7KG8pVieI7a6DosFx41YszZ3FCWpyVy2jRdo8eTk64bjM3Ca
11YZeSSlnXsLzq0hZ6ZwjgHu0Lg+Hn7OkvTdIjBUzezZC1kZrXWKSvS8K27plENJ
iHLTxKGP+r2x0EmNHRDth1NWIRDU8TJzTnxi+nqC9mf0RGW2UyFJSR/Goo/4jsRt
Q5Og1R07QAm0mjnIHF1IAotNuVCLkrRBQ794U5dEAsBvwQFCN8nL3MrYy0ZcjVeu
9T8MKlrvx99eGBx8CqH0bN1pUwNCSi0nOKjKUUbrhYX6TsgDc0o5bYjsQvJJyWyV
bRAkqljBOXO+ZuJ1jU7zGx7HMLRiiLtcyR7R6ikh2xPHa0iNo/N0GzGTLRNo/DnQ
UDAV8HGJP8KcZy0YOGTYr8JI6c4fWv/6eBtVv78mAWI63H9n4Wr8LFIhgdRxmBYm
9o97Pn61ipTCquamwpkabuX+jR+5SZmypNaB0rMo3aEPijU0fHvTucGYcRWP5pVF
rWt4/S1tUS6PtW4X0Y4wcDsk0nNXTVsWWir9a8V8mQgvBE7GY4S1p+n7Iy6eu1Ux
MROzGC0geQwINodN7GlZzL6iOE8lor55qH1xZ5URaW2k8fdvK51DgRvuqRXRL7lQ
rnaaYA1HM2iPfdCVwMjqCgEEJSc0Kp5f9jo9dFNGqMcopFhN5feG0XU1I+WKoao9
CRjMBiGkXoV51e0aY0oAnKbMe+aYyH9D/sxu3bEEgBNIOS1jwBNMat6EPtrUdpJ2
oOlAB7oqs7GQCIXYpLyaaG4qfKxEML3RIerLn7da4sn6rubTvXF1M2G1Bd9IGbI7
FQ1dD+HmGUp7Hx55qhdc6E+q5elSaZAtpB95aM8RhRO9yMd3CElmiIf71UZMjW6a
PSQR+fgUF8Yruicp3Y9nu8A/VHl3IBhGkDp12Euqt7DNwoTJRkq5aHosCeTEiJjh
yOJTCLxGfBYNcyHfwDJJx0DM00u4fKLuDsp4KwUUJi/ReAsODr6bxP9ev20JZoDW
UA+ov8k4h1cAwgSPUomBQ5NeUp5NgoR8oUWMoBW1wmrrmLgIT9rZPp6o5Yhq4tdp
hhhRwqVMMMeqJSB6s9gRCKihbB+sttoF/U2h14bkqGPjq3kB9fuJYlDlt52MuHh4
vNhSjnjq+xQrZBNFSZQSUENVfrB/Py1CCgGFQTnrAKpumpP/b7pH4l+CfZ69nAad
AyQeIbkc5gULqDc9HtdLk4hYJSZwN58xcXO2KalvyEdIDkyT3ng5/v0dshURRTRI
cBnCYQdvOC8c4BAeEomPOBnL74fF5Joy4fLvmRvjRDKlJrbKyw7SsFgIBh9Vo+VI
8fQ2Wne7/cQ7P6z0uVH86wpLCQACFqKp04n5A/GJ7o5T7V8Gk9oYEGwm2I4dj2cu
Tq9XXAthZii48KC6cJQ5hjqwilcPTVGeol5qGhkdPkli5iPGj1iwOvZNI8FqSp4A
qjXmydPswm0SFq+pAI2U//7c8ZQOuyh5hvdJHdh43uzuJqubL2kH62MrmCmOr0fV
rTwJDxuCS7J1F85Acbj8FSMPH57NfwyLKDJBvOW1/fwz/yW+n9lwP6KHqilBbaiB
cuaYfIqnLkDKeXoVEKA9m4znHBzfGhStWmVxybaOe5KZ0+a7hhRdFvp6KZrLc4zf
z/TwuRFvE2gA3HVJ/5ulOkAAAqpNZogLqg42hdH2BC1UAb7HDZAjwaWorbRjGs+l
cO9AeiaGRJcEQkSL3SC1bhLHkqq+2B8cg9NXgaQANqoZUefSxswlqroWg0aDvtIY
ekjoHCJrigHT2NbcZoqjFb4hF3xq5rvfiam2k7Qc2PQagjEBgzuBQ+ZOTdKSciEx
EIMR292mc4shPmHeSRbepYPBXVzYYuKwOvCWLm3DABfsUaaOcNgvF1JcTYFJFPaa
mFuYQXL3i5qHCS1duBK8N93g8i44nVRDiCiXq6BhPkKfKBfTz3OEy3ErgJ2VZDsW
c3EWr0Q0GlsE8yKz4ZRp9vqJpBovl8MKVF9c+lPs6mHQgRgP9AJi7EvghQVukf2W
qw3ONeHbB4KmX6mzC9H2InVSBwds7gpAToUiBhUoFok6oTs/KyvXuxIsr8hbnYsu
YAoNzysZ+CVcscBsYwEdvLULN+lEOWWkFsLz+A8RNC5jXlGJUvlqt274EYiHnaUB
JNMqGXY4p5Ba/8a5wX6eFE7jn480gMdYTeqZVrOZhYrDkT1aZa62xpY4HxYYEsUp
/z4nALq5bJpebo3ygVgRvtdLWLMbr+KenH5Ef28sLmwyD9zNFbfwoTbVlkx6VZq2
6RuUYvhLTJlFh2iAsvL0zZJ1manHHiA18qGfCgCwMqhCtvhwhVKJDEb0CpDPU4rU
PGwB3h60oWvh1PwaYrG/DA1niDUr2rc9f/Oble4TMfdTWpqEyURMCJ3dd4DWqkdf
PgLokpEvplk7Ju0pEc/E9Unv9GxdYRKw8fsK1z4F0twzODQBd1rNJbdSOuz1AXyZ
xy6Mf5z5O20SH9tSW5zNPGlDJHhblFuzVJtqm9uOnqRNcCshbTN5XIvPN8zGLk+P
WcE1uNyk97uan7XAV1RfWFjB4TXdlzUJC1oRSyMqDNTfMRZR6LCjW3sUb+WzuqOl
RqqwNjaafxpnwgE6fnYL3W9btqWXbVXGXe7q26FfmwqDPfBeG7Lr+oWPD5f84icA
r0pHSz169apnwfxUPL9+JuveWaaKr8LhOiwRBUKvPEh7VECz2pVl7aVFHNUv5lNn
nApna9hkMC+dIzvVOFn2oyco6WFxYI7/mq/uhCx/roIUhKFr8qgI9aivoDsTYOC8
xGeQH9+lRQYZXSu/dPmaOhILsrWj7q2c2M+Aann5fJTuyUrR+QsqUiEfS83nJJxW
lWTion/1DtpCTlcXOFG6jG79kixEZLGwfLXTK4a8upCNjvT67QV4+24kVJ1SNOHL
/UE53fD3hA6Ce3ZVI/d3BLrWISfHTtWQokEVCRR9VnNP8RvvGfADf3o4HffxNYg+
WJ4osG5tjxD7od8WV78ZsYPwHCYG7CVZxFayvRuZg5U/0AJoXDl9lDLhIaSgGJuG
XPsuFYNVuqGGebAbxWW0OigsKn7oBhpu91PAkb53TjgOMjB6R5HFLNBIhZTf4iI2
jopzcvXdqBXcl2xHEior9XdHbRhwNwnYVaDlYzd00KIelDw18Yd5Iq247RbEGHjz
45z89FxdXwZd8Tj+LgMLglnzuV0ftznKr2DezkcfrwlqKHAn+epa7L5Dr3wM1Mi3
0zkRkcfHhEIoBpfFxiWs0UWRRvwDmLLcjpdfBrB8lk3mRymYiIVJ7DaFQdYlJwQS
DDTj9MYpoZyDM3/fIZEHmQDGG3XWshUGf4PpdP6FW6kpj2rEm9L1amtzsm+BnvXw
U/7H3I3VpeoXoKaFNM2g8hb+6mPMq7XdAaIaY+xf8I7L7lPmJGcxemdKCgZHCXYW
QPylZ6Vj7fjLxa0dmWtg4la3bUSyaK0lbcjhkeFkqGBbyiIlfbMwfAp7bOM9hwPT
hKwzJpuVCyCFRWP+8byUOkf3bLYB0wz9+xj6/2892Yv0Abh2ttZVVEeR//hFsgJ/
VvXrJefIuT9vOSijtxNlKyF/LYgVhH6oooCsSBJ/6WXbrjaK87+PPm0O3KAHnB38
Jr9zYwmhdLhga30zxLiIE4PO0Mmx8kHqRqjz0sP5MTT/uR528FMw6qTS1UScE0Wx
k/KchHhFg5RL3880PhuwK1ym69EGLubfiAwYyKRIS+TEWi6HEmdSbJgk6vwKWeLc
VYPwCfQXB2a/vdYb0kx6XMbhST1FtpEyvctMD3jwV0ZmzGY65vM6tgemZPvgkY6n
vww1JAZADPZ/wKfL2tyRyXgkI641SlRathmByWvRsBc81uQuiTS37Z8a7d2ZL9ff
YHDH7MxUJVBHG4Lv271PPT3UIkSzsn0R6KZOy7yjIbLW4dSI8GQWImAPD8LqQg5I
He6lFGOqUboW/WmQQZqoY1O1TRL3M9PHFILq7WTu0RJ9rh1YnWZVG2jVkg704Vto
21kvf8SjB9uU9tE/MgURyiFUTyskX0MNxojslzCzFYA3amdmbad7WySZF40BTQtG
Yk15xUFeUFINBUgEHRgDdQ==
`protect END_PROTECTED
