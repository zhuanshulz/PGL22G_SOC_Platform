`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqikGaaOwO/B+XDonPP1Qbwd3jbsmE38TIUP7rmorObcSClNEtEOu1IGFKKiC+3c
+1H781pljAidca9aBlBBuorvdO1hu/JlwQyno2tUd5F0G4K2a+EzssMkn9UJOUQX
Bn3G2m5OB3LhmPpjpGrPNqtQpKMPrpVNTwuslqkHjcGDB6tufGe8tttwlHk438b/
GVhGGyfPeKPwD8qnzZrXg42p9S7O2bMQxfjRfFK0PaiO2SM+Q6FBzrv85a6xipDq
pZEg1rS7K6ltScL/kcOsnA==
`protect END_PROTECTED
