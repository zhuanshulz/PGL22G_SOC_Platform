`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pr89jdlKNVH0Xfw80/wopWMa1mbMAo+UE+dJ5F4dJ7ZWSwMrmCi5GkQ+rF+/OZom
MwtAMnmYfbBZpVLpnIpyio2KiniKyri9vSy3yUxykB3ob3M1jgqyXTlaULG5VT0p
Na3YR4Eho72C4jl+lxBY5v2HLtdett6XhkY2OQdZv+ncYUqyqIyxwRWYrm2P6gCa
YeaaE+tZ9QBglaGskX6TnGDD+TB4hF3+tHN0pielSUhSy7WPxF4UB44CsD9xcOPw
ZQhS3YNVzN/v8KT9R779thRzqSu5ChiGRH951ijNDUbL0BGS+g/KEA70Pfw2JnTb
uoMohzbIqeYiUNPY/FMC3gagj3mPoMOmtn8cZRz3o3HMcdF7ysMiqj342zzyMjva
i7Xilhvx7YTDk4T5FlY5fdyWTIDvlZPEc7YGd7WP3XjhRUz/OQKsxl3DphgFJRFN
91y4VGxop0i0o8b53UqaKdvWvEvWxHRCQGpNyp6/JUXbW84BlCMpBA1VajQ/6mKi
7Les14iBrfGpv8adsWY+wb9z8GMtMC8Oep1Ec8adE4EZOPPcAeCjsINhBR/pnQuS
7XkV+FuYoLDCe86x2ZLnUY+FnK3KhFqTYB5R+hC4TwQygdHqWIhkckzDAIMb1iEb
gkZ/XTopIOaLMNfbFMde8JMqVgCBUNhTv/PjF3Pb1/VpC04s2joso4tDhgbXkLaX
hzvklYGzd8Z6WYer2Y1JZdoXIlXBkKw3H4Xyfclc5pAHahTGI5ZYSTas4zVhVJAj
tEt++tMYZhjmQGzyHWBcBI8zN4MpkouzInZ2IYTfYcOZbd0PEG+eF01nccD8pST2
O5bfd4y4yydzxuZpUX4Ul8ekwV0UAR1Y6OBKB0gUg7oMGw5UgF3GcyxJsm49AatT
0CeNDdtG+cj4erJaStIBd2SEwR+FwD0dflYTk6r8soYdkMmkSHw69gkw+RrKSv0K
ywd7UzbvUWl1FtU50j9VtpRQvqvAVtWU42V90ES0+tR7zS4W0CcA+kpxX94r9NVP
GGXPMq8kz5C1JJ+fvF0JK2hqyiuHAsRJF6dWOJay3YkZXWIUYGbp1akLjYGDZ/sH
vaN3TargRmug3HPw1MaMbYdrNwEVcjhuUxnfexWh5YGUJmEQCxQk6nRkmoxk9WhV
ugDKklHmld0IE6x2LCnHa8CeZVXm725DdiPD3y0X06PtER8OTBBYqrNsPdv6CW00
n+IMti8oFdtbABcfrEpEvkF/RDoxs8+o+Hm/mcfptiMYOSGGWK2kiPI4rBFmR0lv
6lOoZfKlgDNNdsBWlTYEOPWYEo7KZwgOgH0xKSOuXPybN3kgahW6vOloeUVA+W1/
XYSwAF6i5ogQFncR/iN9x6ha1zL+8YQEaVIXk6DS4rgbZjD8n4Bu7Wk820WtjVmO
0JpLSqGSrfGzU99la/5HcZbQQuqxp9c2sfbpZxHsdtuKlwJrdAQQLYXHu5LV2e5u
3TFX9mWzOhKqnQTGaVatBt1AbARMXjrammWTmCkAtMkUYJzHf8+aGAxd8CcMRpzj
GTgjEkBoOyt72cpDshb94XEHWQcFaqCAsGj+0YFi+ikXlDiREim7gpPhTO6B9CpX
s09IfELzAxxpgWeFxQLIgWX06OjhgmpFJjDXjDNq7TBLkUyF8NxMOlFptZqfebiT
1GR3qF/EQ8CKdil0FveW1DVLnmTsxoFl+552FM6wAoUoIG2gRUiHi5pWE2zp8lIh
/NSpjdMxn2YrG0ZnICPgrtbmQxNyAXdy5xgIAn1ACKxceEkw4Hi/0nLv8es6/mL4
TG7DpedW9xQeMSbUQ1UoK43sLKsEA8zluc31X8MZ4hvyQiuZE+DdIICxfCXo8685
hySYIGqcl7swSu/IuUbpBCV1T7bSFVAjsPl835VZmz60ZjC0UO/+/K+jZ9A3g/dE
knsjrcUbGOmn1LSyR5uZh7i9hMs9Vi9GmJcP60jmEA4ZnPPaJPXMwWDE1mN3A1Os
4sx/OT8j8c06ex7h8rglTkvWl+S2rqXt3XMC7Mb0fg5QoAKHXMdxhXoJ2bygz9iZ
cPB2MI/yAJPIdEMoTOfWROQ3PCMKAZyBtJcEl9WLOPZiEy2/GGUAfH9bXEYP2Mbf
hYmPoL+1dk8p4oBS0UDByEbC5+zMx0uj2+mtNF0bMWuti+CedC2WHeRHWoWuiO0C
WR9sD4DmYxQ1dUti2VipWx9o6xvX4RWvp0TijPB6E2HcJXFOIW1IQlsJK+o+j4gO
WQvYDaI8SrNweRvj/dZrqZZlOWL51vrD17mzyzN7u0b3FbrTdqnBVnkUj/qLuuFT
`protect END_PROTECTED
