`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JT5eEvGWtoOj0Yo3/CTNt118dcojY0rrmwBEAL48hTVWAjpASUkJoYoDLSUHK2q9
jL4pQGwL44YWs3bEw3sCNJpRretHOiQgi9t1J27yWSGZBGqypJIGd0IXo7O5Xze/
V4LOUpX119wegQ8IIDChV0V7yTw0t8fPY0apd21pVG1RzqWQ5IEnq+r2XE6ee41t
yhkXuuoobjVbkgKnRIf/kOxjSQP5FQpzUaO/XzuKDKE3OoQKsbJ4fgLGOj6XhOZ7
BUpHfjAbwzKHlRstV38oNm273BZgHexxn6NhxBWquc0GPvJJKdYBNmZyoxIA3Gl1
6873cK7VQXdySrWXcJzQubdxD/LoNqNAuHMhFFnzWXEzkL79lW11p/JLlKGw5kCp
Vi05a9op8CMYLj2hROTyRoaHbiDci+C1sesLyzabJ2VtC837spUzeAjuTQk8K7qF
7QbHLMIE3FU6Oc+W/GPHciAl+lx4wAbv1FXKin0H9IjxNVbq2zTAZgYnqYtyQmMZ
pfkTTukKbNEZn9mMCSVWr34wUlZwfep0orz8NANd+y0G5lzbgLemDl6r+uU081+Q
JSJsnR02h0hc8ZWxudssScPSiRLvXtMt6FXNxX7swrd721WPVISgXf5QUbb6Oejs
3NdBIDMjM+bBPpkSPMkRDdkUhYZdosLY2h/2Ce/zJZwe08LluLMYi2jubmzDV/f1
tvvFPou/PIfl0RPthQIFajt5rfve2EeT1XEW/yx3s4zFKIDMKKopxhgKDiBjYUGL
14OId6edPMKuolR8DbgzflUUSGg1OXtSpAMhbfLcFyUxLZAZp3oYHMeLuVoTJqIK
ZNY1eMGA0F02/on93C2wtFdDEVKZjFZX9EYnIbQRi8Yodrym9PQvxQgiJd9HYd/0
N9XNZwkLVUDA4koocRAILrn1NtXsAzbstNzoWI7E4V1p98pP+kbClfa7UX2nE1uQ
9RSGSO79do8VgwseGNt0rBW4xt3D4Uv0i7ScIcFKAdnLUyKeeGqPOLwle6qiwR5i
yg/g5R3egnAwI/yBldBUDMzFTglKqg/EPcikaLSPai7/qlKewwBZBTP54hD+bbxw
`protect END_PROTECTED
