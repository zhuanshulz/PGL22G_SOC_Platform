`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YWCV5xgx8OIfnEFvI6IJnRdliNq9tPC6htE1JmHGF5B+m84d6kN1rcM8HmQNruZg
iIk+3RWebViyEx+8+SIVI47Il6OekruY/nQta8N+GI0BbRgsVgky6ujoVzEAx+SS
FRk8pfCxrrcZsT5xsnEMV8KXXJGPJCxu4LSJNgHl1Hp9t4vPpY6AiEVH1jAUUFxC
dieeLeRhRSYQ9K59y/Y+9KMg1RJfhAmgpOq2wZNqYW457d8VQdJVfAbbT3YyzIbj
MZOdt7eSLCEjlkUE1ZMzKlw5ekPDbKEhdortpX4/+ekRogZ68TmPJECHWm4V1All
as2n8TGBEjtq77MxREm0e5jwzkXljvrQ7wr11rD2MV67OHF1Y6UE2CHXOrQ7FBxL
qlzklTDGQxE3uZRLfSg8gjpHcjCHCx4xf6dt/Do1XQEgfjVQGCdgkX7JzhQjUHJm
dp5pmkd4X4LDtcMEbhosEPa8O3pzQmCcfQux5sv0beIcHMoD/dKQaujQ95/Qfs8k
mTSffkufQLgZp82/c9MVFwNY8zNdVFurSqI+j5zCYVtWEd1H5T1nvjsW5g0bykAO
X00Is1DL2R9kHU1G2A7gmiOh1iGIF4NthYHTiZ1QFzxOQ8gzagP2aPHs6u39t8Uc
hCwQwScxabzWwiMWp5yuLjwee294PIiuv99X43EL+AkbqtyLvGh2M0NNOKXYMcZd
AiwwDKqJurB0LQO/SpUyGRxKASOmp1DqTnrndHGOz8N21mqeHx0IrKD15V7aPLSZ
jZC6V2eAXKGx29nDIbKdydJRZNMRigRiS4kSmaFUwP8lno55fNQxUlxCmGEp14o0
c2mPN44coTOJwRulJfjYjF5DabgZrC301hfEYZW38LEtjldbQeWfnAyEYp6nO9AW
7K+qmxCLuqvhvBhdMOt1WyWstkcxQvbmEhTvIHGTCCWvXHuhOPRQUUqJYmBvA/kD
ZHqkPk2unJ9Ofc/reNjEa5YzbQQi2aBmmKOGYte5ISwssd0ZVACazHJnNZ2Dcn7M
zC1QBNY3f858HWgi19+ohN7kEeafu3uTQjZdvtHuYW3D36n1fwIkRwFsTxsx0z4y
euNiBpNCBVrdQkcHSE0q/h6n9d9mcMq91jyk7j7mEfbxRgFZw0WtDHRMI7v56VA3
KUwr2It3xaFuX2NFa59XB9SKkeCt4Cg7gX1cXjczNzJhB8LhxcA3kshwbcNIIdHM
kx5WI6bz+APD5mZGxS06gPX9YCJW1ZG0qedn3giA8A9z2cIlhA06nfcBR6TOaZgo
f4RNIwDj4FKCTkrIGb/ZXZKxBCUrDDyJ/1yYFa1K1JDFmbCJb84NLh12sng02YB3
kkJ9X7/cMWCi+p8JeDCLlN4Jf4BpOukyr2WFtNUpPXxZc9xYP8TxqSghmaeIKzTZ
fYbYvhEH1knuhmnmyDzEJ0qD0GeRDm0NV7ypRFuts8YDSUaGpvRE4BBdawvDPNQW
zJH12AFJnN6SxQ3nBsHOkMpUwUTynYZiuqw5fWUWTCzetiYcKGKFB3ub5qlYkMXY
X3w5eMICkqwfodYqSYRe3DT2ArtCdEu6tMzW8FQUR0CTHL2lEj/IHPoP8cBaaZYo
560BQdGafaubooD8N9xuuK2Zic58YXgpuEzyUV6Kn29z8EqnnlJd87mtMggG/d9k
h12g8kVtcKwsJ8ey1FVHSdYgXyJIiwGC4JL0+e+F+ux6BMYeAYtxWJjBWJR9o86S
797YKHzSwnbJxJQJS7KwxkvlswqgNAMvcJ0+S9TGG8jqRggAM/dhV7vuqT9KGTAy
dY5kXcwSwqVoptfj8XxA4ElRoYVltGfQu7u/wVRJu3fAnqE51EFa8++Xd75XQKzv
IujF6aFt6wAN6lZllBsHC8V0lpPhOinnEmN9Eofy3+OzrPzDgfAFfRe7lKT0QnbO
lCbkf1MjXtVZMLcwlHy9X5KlguskA1jeQ0qG4eJAseWVZ8dxUdcA2SeS9V0HWKyJ
rzTw6Kk3hL6u35T66bkFmDKdMKboyEcoscynnlywbBzYP3xoyxVbsIhiO5ZFTxQl
z83AUoPq78Unot6igB3WORmF5gVUUTfPE7Z2elXwae+OYfZu2d/5Mo7GZURhFwvU
ZxZZa9Q10245YV++CvUBKe49u78KBT5cRtvg/qZHvFtuRiXdj0hGKthgWLsN8GUd
3bLEc9t4E9v+VVukshNYlq0VAof0jpLX0cpdi84B8zX8oS2DmDwVLC8Heg3b73xd
j8MOglzMtOVIPK9ysFJHfKi4goWhW7q1mswmvrDO99xEP7i1qjqKz01Ye4ZKm2Uh
`protect END_PROTECTED
