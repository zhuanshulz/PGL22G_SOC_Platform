`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6oN1YtYkL0muu7qcmtGrg3lJlck+ngeUp/+EE50wmPkqmUhvgp9MnmuDqKFiI4Y
sVT0jfyOEnF+ufXlDjnI4OETaxvkXteb92Q79HlUDRtH3qfasOIYfHSMwq8KWryL
095JyzpuheRXiZ6Ft4qD3kfpXSlvzcue0vN/vRSJLsxJQUJ7PmnU4XExndtBeb7v
Y4ttdQZmRwfgzsA/+avFfLVuQubOO8w4zYCDoUY/MyVSWoyNrc8jzTBM9IuywPTL
v7//4WKUsrkfmWK661Cw9gB+i0+8JndsLAb9CSxqIaghR1RGIdGQj7ieA8nvqtHJ
ETSiXNiElCTqViXDyDlklVMAyGHxXzQxlyVwF6TdEi/sOx8WgSeZT31kmleh78XD
SM0GCdGZXVdr95q7B0U3pKNeSE0F3Ny0yG/UGg/KdxyyUSspCTsqGOBRb6/xYaFu
tH8/FYtVeMi69wJCRmkTM3kEsdfQhdTNszEX+2YhE/Dwx2dNNxCBYHvohiGos9r1
NYuH29A7fJMmJ7VJ9Hejf6lit6NFGNSCbi5i4wbPCeLqTdGEBywBKHZ6Hg/ZCnHc
mte0KIbtcqiyxZOHfjb9uZideTbqdtwbDmw5WqJkkEURjHe/xio4FRcQopKnZvz3
YMJgWMpzXb9E0pXfdB/I2SdrK+zAF7bDBtF5/epbzEEvyrwwovCAbu6mprb144DK
iAfAklLVgIPi2gNLfTBR9FttCcGEhns+5XAo5dF4mx9p2n4TLh7dAylNpBwcusvN
7gDnDkDaUAzs/Auf/O8uOa44dmSVihpQ7hCxvkmUJAnsc3YLQ1kBxAZZFV5EmB1D
0CoKxch/+WOnEz5DslEJXxTmhazS1jU3PmOk/oiShjm2k7rOYs51EJlr1wcVDW1l
8XZfoCfO/Ttq+j8yRxWgzJkt7xwwG+QOu+28MItUW/cm2DlpRL6V6fwfyVBi1pN9
FaN/LlpUzV4bZ2p7BNuuYjSZm9jrKqJB0Xh+a+yxotaNEte0qKSK3jirGNBLRNUg
gTSYTlhFTxdncsS/bux8gYH13FlkVlrbYCmFgyZCEqjaXzL2zyKWYfIeR8LJF41/
pFX2PXX+3dCXsZ6ZcguiC5KOfcrms09ZAd+6IA2hqlpZ42Kq/wCh6BwyljbjwiJn
O/5bmdVBehwtnww+PBpfvoLM0Qp/iMjPVoFNki7xyYpgeCCIcUf+hTIJcpSNrJ3E
roMXhhCNsIA6g993ZRuUiowRAQ+Rk2SLS7ySoNU4GrlX2CWKLmRRKNnK9CfhD5Xk
KUfAXc9yjyO5mI1tNIzyhQ7qjYv24FjRnlAOpubCN//zSS4/4nvJpAi7fHflMUv8
c/DrrJj/dBYnsqAFsK+i3L5UHVaqbqJ7qaMRbDv/Zz97HjyqLEu/jeIunQHjywiy
l4/lZRY73881kG41p81XneTA13rf942XJXN8NYcc5mhRKO27hTfN/fizw/H+rbZK
usOs7/k3JP8I/0fqGK2RFnByhAr5qipKGZ4WMywTGGxT95RDXgyInKW4VIadxiLE
PQLRCAx5anucLSs1ZPdIagk6Q7IRdhpbywbcuOIoUkyeIED/8CCEHksQGBeZUCKi
1lOU6zckAq+N9NsE9xBqM/J0uRsokimqGL1/nw+vWzn1Anw6IGantedCSr9KCGup
keIcVXYpDfaAH+M1g4SJL1l6y65ZhqWq9Ps0VmNM1e9C0+4FQRZinGdK0w2oOk+B
+h/ccFdpgzFDCKDgGhdx23WwBv5THO1nAKdkp0Vz1bKbTbB6wHwdjvransDSxcAF
LCPGPiVnNInCxPU1utu6QmKq9WYYBoFPb+iSGx3oA3u4Bo7zvzjad+s1dc73V7mi
5g/5mEzUamuPupgLMqQCs49C+Ruh9Q9c8vUEeCuDznGbOTLg9FiT45J599y2NDdc
tbsI1Kc3wSvzSMsoUnbiazlKexeXMEv42Q4v8YxQ6fGURrv29XGfoJ1sppRwJOXj
9a7uJ7mVZrsVMjLI6nD5htk1B/WGMpEIT2NcWjfONrR/clPPK2kejjkkoEcKb3lA
fFRPTqG/Ac/+wDKUsNrVbLjkGXoQOg5vu9XZ0N1ezqi3CJBVyZyVJiwAndEAOrfb
Mps0ipDwRcg37StXUAQg0/iXonufHaapZqEAcxY8BdnfV8epbRJ38ZM3g5nIflgC
LoVlT5/fIoSWSDrx26JG1asXoH2c62UHWnsODXa2Yl9p1mBXXStDEUKIt/TRpX52
YmLKiC1zo9gUUIfv3bOQ/Q==
`protect END_PROTECTED
