`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BUk6t+dHqnaaIuvvhgRtjcurNKX+v8nKspmHJn8LfSRIoylRwgkHAJO02vq90QCn
klWWn9d7s/U1WmM7Ifg0KvSd937TiGO1DnhXJ+LfBWCsDbpsbbFie481bvVf5R4K
VM4OYa62Z7VRyN0uPWWPylSE+S5CRlkl29wlMe64geXPaE9rY9AnvAstt2tK7+Xa
EnSpyIVLqlN0CJtE1NiVOxBFDf1XhPGMUx13EQmReK+MGf4olF4Bu1AKPv4bw0FF
4xidKGsUfhkj6gmvrOyYY64Q76S0nE7cNL9oMDYOwDBhlKii/61XtYFUXx0Ba8Vb
qwzJZA9tGjQUEBWeVViiROEgjyu6wnKqUtCzBwxA6l5ouymceEnj/NJwcOkaz700
R0y75eFBo/4CjkrM1cZe4i7g3n3gGbUbio42630auvoHkXBWg8Q0brKxxqWcaNKn
0MJ7BtWUI7I2m3ropiFQXlwf7WYJKWWBp/ghOmGcOPsNvUCq/iORyscfkE/3/2ti
jcVQJoQRjK+B0VBt4VqC1o/tOTVZ3ZykYb4RzpS9YfKG1H9jQJ9JI9IUl+o4GM4o
5Jh8IzQMc6UzrMIParrwTQIOYgewf+b6egEugzYjqBN2V7iEHlkH/v7pHyyYvq1+
FegLt8CBn4++IqhHDuNY5KNGoVAEd408TbXItQNcrct8SWESPlNEjr0QSbdvxHx6
i4FjNb1rBtUVR97Ljewywj8KyB0Hk1Qtzf+lJu5W2BDY9jhKq3w46PjPOI8PHwF7
YOy2mHGe8sK2xQl/ql81b8zU67LIPxx7WKAkAFlJZYQ+p9LgC3HGz5indP6yR5SZ
qCyAsebbuXVuxQVD2cj3ZQaWBhMgQWcfmrrsrAGAbMbBI/I6FiCjg7jzs9OwxfgS
Ku0PS+zYo7Gyh0mh2cYDwj2F8Wod/zvjNbNmcrvqlTMszjNn/jkfl1bz2SrkusQW
kXxf31mx2Yx/S+88MQ29zLw2swA7SSwHL/Rrg8fHuAg=
`protect END_PROTECTED
