`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0SZT161ebnR3NTcf4pxNbRcCqua6EHGanPe/jj1K4Lg4diDqRiuKSTnv/Ovrsg8o
V/WLdETxGeaupBcjXMgZvc8BQdB97BoG5m/6g8ka7lz0fFxgsX0QxQocai9SWJBI
TY/NxM9G+fs3VBxzNGleEs2LpF2pAzSe0FBoAvDxLSX6yQO0RNAGIxP6Sp/lggxP
K2hiP+Ry0GifhGb9U5lG1Es+Flj55X+BBgWHgdb45900KjlBniZxA6cAkk2ixxyj
U9zH6fU3nHy6l4P+HAXZ+wRTf4c8NL9ONCdLxQpyBKodz4Z8edMl8wZDQXoeRJY9
QOGSipIBssnp0InojRQgLJ5NfoGdoGIYZUNGdO3FMS42ae9YMBp3xvoBsG1CAzqH
zF63QgS8Ojoa7jFYA2yJrPgXUmQSYnk47hUvZZ3GsgNI1U9Erpy3B2Ff9hH6fG7R
xLQwdFSVAP7zAvVV/lJe2fH8kQvc5EH4Y/aIq2yaX7+ZPVcPA/NQv4WmPrDc04U8
vYvS+Tac7xdovSFSAD0Th+MCy8cMHJMVbYvFcY2lXMP99b5BfokS8AhkZ/YDf6YP
z/S8rtVISRxD80GZKqkTW4yqQzW1gzOSzJRAclaBorv9ls2Bx/ly/2fmhSa8aqF/
qS0rwl6evnRQZ7ic7CPVYDYWhMp9PdyUo9i5eK6qk9Ego9GUCu6AvFzrV054KQJV
`protect END_PROTECTED
