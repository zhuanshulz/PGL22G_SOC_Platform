`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flJan6xyi31je6vugBMyjbB0Bj0HOOn4YgB9ZhqoBuK8R1w8CJ+rvio912GttkHU
vWTWLf65lrI0wTnhyRrdRA1pnbc9PtsdR21uSjzyTR5d+Ad3Xh+X5akWw7NkMT49
O1A+bafj9B3I017Azhnhvp0Nh+OSlXOqSo35t4aK6ju4DiRdslLE0NAolAWaRMNr
rbj3lW5rz75LcVSJILkjA5QIYrCpOsVkZFHSvv5dOQmBsj0fP9XERFaA9E6KbRLf
oT8ZfoI2ZI1V7Tdvd7sKuQh/W9SpoP0/XEOIwi1O+oQLZ+QKjdogroD6OsoybJLS
uzu23JAdYFq87oKvcrripF3QXkm4tsBSwCnwF1CKTGM=
`protect END_PROTECTED
