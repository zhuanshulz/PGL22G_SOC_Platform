`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m/5OJyFxaZRRVhCjl7JXR/YNS/tGxK1SC/OVeQRPWoLAnX3K46IqZMLLqy94RY1b
jO9g4NKppVfFhe64YEGpYQPkBO3zjhZ0fs1rTN+LZjuWae/dVeMHeqs5DFn1yuLG
iGmuaj/iSffHaxygHBQybVN8YlVs0OiJSnn1GDODvc77CRzmp9FOxB0eaTA/yWXF
vICOEjiinfUbXx0FFwRJhO7gIF+3WfLKJjQqbQRt5OsMKTUHxDUEQboRO3Gsh4oc
Sy57LZ9fa8Ds6nq3McSHvvw8MUehjXe2F9XvEvr3mNj9LDbijM+dmNodv+o8oZq1
mHFJ8ceUUuQAzgVC3vOoHaXnjw9tO7KHbll2A0IV19a3clE9XJm2fOd14nGxlNAk
NKmSjgJwOkN2oCdj6Hqg2Cgwqw0ZwX7wZoJT4i+Ffe5FBigD9yEzDD0+/e8VCSBf
lX1Y+8OrE7Rt90NjutuGsALci4CO7R18SDqXREFa2GHOtx7Km+qFvBfJR5R2Vhmd
nIXh3cPBP9IAuHbQedRNKtwFUHmdLtbl7zCzBtR6aJnsdZfJH3dwekuWf35F8E+e
UEPJWb43i7Hq8BBn+UKui0CVVqG8tySq6evls3pU/aoxy9VQJC+nkWe7LdKpQmXS
GMIHyvlJg+uMQXU05l89z980R8mlCOJHGzP+8iT1sZSou9B87uMTJNmw5Oa49xmY
qKSU+wefta2n/c1bBMrXNlWG8fN4buNnTA2uJFb8SJFuCo5sUEvMxGKjN0hXD2Wj
uqP09yBeexjsZ/dHgT4cG5WijTL12zU3wuGktlvxiNIGJ8ShC0LfoX2d7ej2ulom
cE+mBlgg8wk4apWfQhZlhYxbRVZ4wKupBRhsCDYyE2Pt8RbNIbCsr8waBa4gD0il
9BRAHlv38TWSgAy1w+YIDgMuxFbXYqb1+PyYlHES2JK57u02enwI9OrzuYfpGQ0O
5KslSHuq8YzqE+Cehfcvns8ScnLT0szkOrzUWa6Rjo9IpWj62c7hnmrNKNuTHTfG
V/L80dn+6QsV+81HI8+gZvOgWBfL2xCIDoLCHYTS3Xwc0aiX/NI5YEdj0+e/nFDY
eYSuXwMluNVy7bb9ph3Hq8cL8/EN5rWvvd7O0ZOFNmRjFerMJLrI0Z8tF3szlqR5
rs2QJWRPRsVh12TNUegJMrm5+Uk9T2BPglPwkFQljVgIDDgcgVJBfUrvwXXbYvV/
1+w0oCdjmauYUYlufoP2c7/YqkQMnLFfv5v3XAJvXhdOp8WQNhCbo+iQiaIJUVof
XdsIXscS/9GdCe+N7CNBYIwjQNk0P2jbYLmul5J80Sw0lUhzux5KRg2R95/zjVwc
71ZwIBB8NtEEw08q8RcoeZtkcaylZYIPFIGp5xO83T3S9Nu3V4ZkwKtWf9o49YHC
Ndsxb9uhs/OIQ0UqBnwNRDyWXI3aFpXEOoUXv9x9lk135tS7gbuXR9u2A9J/dXqL
8Gi/syCo8mmI3DVSqkHXXh1VBdiHSbuaeFCotLPJwovgTWO8ecjynZ5OoJuNCJwU
rg/XS7Ia5QjeL8QNThm3ty/wxD01ojS8WvjyazwYUYT+rn3JnVAXHsdohjROSbeX
RPPxRCgkbmRO6osITKrhBByzcq39z7f76T8OssWVHv1j8Bv8PuMO/lC1tuj8I1WK
qyfQ8dVFYwvMyLFllQk4sxnvvymMiUWx83NBWkplBrDGqK+EJJjVVS0R7lf7l4Ab
w1n/dHMu5MT97jgQy4AbGThR1jo+0oxvkL5U4zEK8d3Axmt5aQElTbDvr02KwNbO
Mki4z37Q3D+XVCYIgJP7obOmfcfZvwO5eiEqSgAbKq7Iu4v0YK9TJvgB59hWv9P1
1LYcviZE612rknAEI35gQPYb2nAoqd4zla/u2DLTMAiDD8Zt0Kaf67za2OnNhaN9
dgGpHNV6g51MP0PTPjQJTqdbbhqnb7bON3/QVeVh7GhWOTGxOAS4C9+/aKUykdIQ
PBYA2tnKtcBXwjchPEWgTS4SLQ2aZCBpQCK+rXeAPQtNZAQlRxeO1fL8qb5gCh89
7fDxhQ2Rh1bNJKoUz2CvorxnFaTHHa4pPcKM79s+EJ4TyQx8sd/YXcZa927QDJlJ
D5ZW4PssdAMMSvwhPzOjw5NmMklhFsrbmG+VAqs/9t4WSoGuFu7+phfgvJlyBocG
5UThxGyy8f5JTlmeRTUE9eVdFRiIbExW0apkns0GB1k88YZ3EjmQjVXSgD0n0hI5
9PUmCPTVc0DyikmyX+7MlG6YzbrE8+j65vrskrpAfO/tKTf7fTVhp0HOd5R011F4
mzig1dS+CmPmNa0//gTQHrZTYtjBwo/lCWRtaM/UbWRt3hR9+ViEZeWroeenEc0O
PAb+dAVNBunizCfyU4F/QKiW7XTDlTgcUrZv4FmWNhQ0VYnEN6ZRFrJXIr0IoVZI
6TIoCimdDZ8QZevniBqDM9Zi3M6Rxr0Qc6ysjl8Wj3mM6Tdi5mtJHIX7lQiBR/nX
hiP45r1rPVtskqfcTLjM91nSlNz1AZq+oYD0PgGLSnh/jIKMHJcUwKpqz/TYDMtM
BN3qPlHfax2zXKCJ9uJ7IAPADYFnm+ODBli+7psN5WVQih6CyvYigQf7lt0j27zN
fzIGECtUahn8Jy/R9T2VrQckMrMlw3Oo184yDVZ/Go8qzsCuTm75QdZNxNHJrZ1n
Fm7JdxnS5NuhLhOeJ1mMVyFUJnllMuryHkANXWgmYZ27NgPzbbKuqLav67cRCW45
WgbKk8X1ZO6NcOyoOBBW6Rj73CpNY2IGfMJ/rcWd6ZnAKbHbYz7VBt5M//U8DgSX
fWq82vlo9edhtFHaz9bAFH5yuSvOs+bbPmbliOSuJtjyOQDlUmSAl6saPkdyDjIy
`protect END_PROTECTED
