`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
izR7l0ibw0gveVg1DiIL69BiLRaKAq+/zDsesJG4WQknhWAUi5zANyRTg1s9ivVd
maFG3K9RP7Soe/vfDUIqopx118umsVB+dzWDDoSaWJXSV2wRe7yp8ubfZwmh1FLX
WihKuNv2YPODyDbhGM5YBJ/xXF352GA9mZE8UD2VFWN0ROFxvyMghZ8RQF+/byvd
gEWgjRzUKRecXd09iCA4VMiMAWqrdN5ZrU3n08JqgkkoeBeOQl25zayg2cJkOLXv
jnODBYGr2SfFNY75aRfo/FVHks/gZhWj7zapOpPUvOiYM1ULwMnivzngk5w4rsdP
RwHtkxs4s+zb16tRHl9K/56R7hZCNztOUlyprPzANDrOz1nmf5UW3W14BDcz3sGg
u0wPF86xZ1heO8KmX8UMqEZasoem9F6erENW2eZfA1n/x1XtH88sHyHASyAbyWLL
oUU3CQeATTnAHgi7sNMgXF4iaD9OwSjJ7Wh4SAGc1h0OxhPP36UH5D5+n0iKSRce
3QNSD4FAFyCvJ/FrggrAvXg1TixzyeqsLyPrWBeqEJ0=
`protect END_PROTECTED
