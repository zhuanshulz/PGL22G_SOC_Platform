`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CihmEb/GvBZnB4gSqzLNpPcFkf6o6GiUdFttq+DIvep7t5uhb74ZPmFNok3Ba02c
Ce8Sgo2ZgedhgP8NNO8vLuiopwbzOi4pqF1w0/YsOP7IDUoCEe9OQ9sDS/HQl0Zf
lJiVdH26NwoyRkHAHTQ0PFXQSefVSQcpHpTn4/w5ctKdF8F+6TXLXb0uXlHKUdCT
06M4dHRclGAGAmZlDCIMcOmhd5py0LPUygsmAuqOt4zFOsTxVFO/vxzfoN6Z4iPO
gTFF1zbbP+cfYpUNCCJnlO66TxEruFGmkvDGg/9ZvDz7cWe3sa3YUaZmw4TDjmBZ
fdMtV6baxs6kUwUeHVe4L40V0fm0g8KOjTwiWlbWbiNjDuyH0hty3i78JafVPYqf
8L1ohN9IuKfG6SNavxjqSu6u0OpFDFpplwijUnimJYyELY8+0/jEUmO9x75s89F2
`protect END_PROTECTED
