`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+7bp/VMSWPlS6h0ICDXIc6a9XCaidXIx2cIKad40RH1J/6CpqPyac3JHeIFmTVJE
1itmxrIJpw27qfxfwxSvuPKMjRq6P2I28IXj78CAkRKYcN5PnshDcie2mwbUJ0nB
bbFhmMwBj/CWyU+zqMrXE9TEKzOcLmsI8kf8SsKI8XVkojUKt6hwJXnMrrM18KlG
ae7gMn+UFuAMm0tjShvh159E5o5O8IhTvbbU/66ALJyWsJ4NLoo2+E+fe53ZSEr2
Dd3lz+l3JfnVcS1HcJzjdM7q9LtqR2XA2t3qba318wZ7Tjss4nlWiRn+6zCD23ID
kXMtAKuiygKUjsf1cECDuoH1x3WGAP/KlUDlYdIlWjw6d1bwLR3DJ0ShqfyGoq27
FCok3RRVgyMp80kX6MBtjuEqm94L5CRQJ9Kju/ADszmxU79f3kEv4EAdPSjhFoLi
0Cu3X4P2cREZZqJYl63G6ykG4wgOgD6HpAixsvsqroCYjrE7aR5sWgSWlIOa/4vd
HSYnWwCcXG/PP11D6XWfwkU7A35WQrISNT4sWP1czc1HY4WqVxuk0DkYsxNO4mzB
E2z8QjvGwO5wLxsDwuW3QgOGu1vQMD4UNMQr0kISUOfMoUnVoFFWnriSmnONF2+q
vBxRHX6PkNDwQEic9jRq8pHe1Pgvs4hCA7lLje6JHFoUctQttBudXvl/38314ghj
cjI6yYCrjrHlieoown15byjM18CGuo2SzkrICiS6ybQ8dBRzuhsoOyHuZX2JGEai
5EOv2cir2Crpil/mt0oesPc+p15A18XoEy8Mwx+XOdxbMlvUG1kUPV2b1nO2O6dW
wPS6PeTIw0eQY8r3RrOW39fFfCcUKZA6cbOahncDr+ZSu2p7O1P9ZcNQg7OCKMjK
ycLQjW+i7pu+i1U3kUnKAyy8eIHPvf2p4cJw3lSA7xSW6A0oMLgBhni0FqzmhxLI
TGItPuwQukq3WyknZjHdVg==
`protect END_PROTECTED
