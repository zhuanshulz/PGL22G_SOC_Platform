`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TfPHwwEpYGlI3w7cgySPmoOUwWimusL1ZSlyymtPCssCh67UvIBcnm2B5eC6fHsE
R08LcLgcjS/nF+EGpUq79HNkKosJ+dT2w2wIJ/pGp3Nlt6eJ9zAN5L6x87FbUUqi
h5uawxXCQiNs1t6l61GOL8ecRfQ5k6EDKZu+sWbV+sE0R8ndQDUgkAOz+ExFjrEW
r0QrKOjBt8wuSn0vdjNN5judjw/Kr+UuavDMbaCz8/scs/eE7NbgEuH7z0UrHbRq
BdMiFBKjUn6ulZ5ZbEWFnA==
`protect END_PROTECTED
