`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y3rdyimoPf+0qnw4D60+8ouMeYpNj7iwfifA4+cEW877JqWkj8UgfqQFJf76tv8n
s31cxpqFqWLSksfIjnmp8mYP9OnAKA10/vM35pvQ7I0581lWNzEM9fj24JlaS9uG
a6LrfFo1KgugwbXg7SRdKIijPEnP7E7QH1W1TzSsiafGmhxPyYmExlugEYGZ8WSE
7vJtxeCO6Fiu+N3eso3q/eZfGgCUlylM6Pc6uDkwYg6WAplr9JssKFFi5eeUTiIJ
lNaU/eUt3lDm6AKX002xHg==
`protect END_PROTECTED
