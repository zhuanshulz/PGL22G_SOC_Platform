`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FMhpJU+p996Aof6ipivk6h4j7dL0mvzrEKpcAiO5hfY5C6j+/Cv2B+x/HrjscRPf
pZ69HMOCUnBLbtMJ34QKTcmTTyXGU9uEjOaUwm6j5rEi2ZGkQSZc6kPEbA05qo5S
vhcFzDLyOJDm80wYGWHvIPWMCQhoEPXFUTQltWBrZlDElL0Wo70s/PMA4cjh0lY1
J/c65G6sRgijpO9b2tYjCjzY/QDFw8WND4mNyuyJV4OB4OAAFer7HLtNJY9VQbXS
15YqAc+j38SMX2J9QsjD8s+Tbm1Q4gWMELlOq8CvGYRl0d6spj4wpRiGOkQWj5T/
o2yMQMksOF6LBEnl2LKU4KvgaUBXn9aTf3th2YIRhYwrshftI3B+u1IafJ4obeYu
9m5P3NKccY4FwhkzzfB9NntFlJBeVQsSgcY9u4qz9Fb7bpU1nORxRsJrNzOe3at5
d4k4CMA3HzpydsD/GO6Z4q6Xa3Kr/vf2ZYbe5TcU9KlffCUOKAzMaC5dwnVRhUfR
nITCklZuw976/LXi2MdYDQ==
`protect END_PROTECTED
