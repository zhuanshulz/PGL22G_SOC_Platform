`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JrUD5LELOf+QGUBk3A2esyXkTTEyssejgc7IBZleq5f25b5JhRr32dsyX2pnPpqc
aiVUFkotYujlwTYRetkP18idog65WqQeRCJIPus9gjREaYWTCPrBsoKPs5KPG5dA
mWLKPsL9Tkpk1AFuSQ8pmnJgcXaMNVY1VGpEv459hqJtDGiEAG4OAmpzMMpEcIxu
Jh9/gujNi/+S7W4YLKm7o4HXwxGFOdGjjDoXk5CNwP2dP0KfVTi8xQYuYzSnJh5F
Hk6ACdlsW8ESX2SaJQOVUCva4fww5dCw0WJvc3xFYwKZSBCQARzMgWTZCHFOu3m4
RtqDq3mzBMjDrdOUvm4sEfJ3zNT4dkxs+E1Yl17nIb9dol9kJSOkfqPPYanN4DND
Cenu1PAIqo0vuq0U4pEasZPyycJiqJGuW//SKrcjfiqqShYkKFc0PG0FPOryQD5K
qpl3AlQyFCj/sW0/kbxNoe0qs+CvJAWbyVe0vt6yypzKnGZ9HsaFNb+hoOSWdhDa
EkmaTtV1Qe5xYmdJ6xNafOzXzWDzuqIH+yxUK+cq8RQpegvnSQ3B8FnAWoNw3zzc
HI3ad5VJICPuI4gNGzvDM22UltWBG1vsGN+xmAh4tWe/iLwEvdCMItWwkRVi44e4
q54WO3ZvE8t2OQmBT1yDCkcy/HGZMfr7iA3h3XVUlDPoNtSRaEuHnG7Dzsf7h5JQ
`protect END_PROTECTED
