`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMXKoHSrchgokWJY6PwsykWXJ6+cG490UmIOCcw6vTlaLUQntG/E/4hcfssNk9ki
JxXAk4flyuSP0p8gk21bHqc40ZcNPKQoXtUXGLzMl+ZL/ssvcIuCALDOQ+p/Goan
DM1z2LHkHAQOnx5rKUyESjr5DSH4PMq7tjGV+D2QEVVCaKjXGphBZA4yZQFZJuK7
bpzEqnAvcfGUx8Pu5m4yLInof+G2UH0+PVMSrsHfGepuEuvxq3soRwyQl1lc2gPH
qj4I3p6TJKmnTSTq/6lXRkgCSPhsPCW3GimLPX1idns2nG5wSA5Akf18s6/IhrQJ
IEq9AlHuQBebARQJGx9ss9/GX1YDpbUhraO6/f7v+GkwQCjZj8n7PDMR1hcVKRNT
2ZxZcaw+zYz0BVbAAOo9BpSTdDba47q+86H+Iuz+CeXNd4yzoSh0tWGMhyVpjdrY
P1BPlI0VsP0AXCMmxBvZNpsUicJesTQMXdjsgTGUv9/uNdLjteK6zF7pszirkAg9
Uk8S5JPK4vpJdjIrPd25o8eHaZ7kSvF4Y2l0BnrMnxpwo5x0SIqZYInYcnt/g14q
2PySVXE8Pg9x2l+kCybzO7u0g/N7FlvSZ/VV+DnZI7By+77AMciOc3bJrQxaDYsQ
aFJy/aTXQZaoDt+HOZbUFzWQH36ZsHIN8lqxeSoRfIoFEE3W+blPhdj63fzib7U9
u+3vzoGS/WU75vRt97MNHg==
`protect END_PROTECTED
