`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LXtyYnR7dzu6NITmEvcc5j4eOAlPM/CEmsEEjDM0QfFMBeMJs6El8NQu/KkCIuJl
bwqqlsTphWZNde4lfKI9/1amglWITPPxc2XWdr0y5rv0Hdh38wgP5NoBICt+iBeZ
5PnIk4CgTaJqRvOlJIMwu43woSc7fHUdTxZjgFVsSwYfX4PgK5DYykIAI4yyFRcf
4yCRToi09xRhQU5tRs3GIl1uoLxAJa2oYXm1dAuzqUFeBWrINnXQemd1dCbD+FuP
jIZBKtZUwb+mn6nsn8I957mpeWI5ujZVtmmMARKdjd8S6h9iLbOzLSN86RHnzE5o
kvQV32KpO1UFLheGw2X0/AZdK3PTiRypOoO4FEjgTNCvLDZTqgA3YuMPB84YVPvr
rHwrJtwKmswfKjWMuqm2DznWtDWGIouxa4aaDGJgYwgioc9R7Zz4POsIfcIEtsBY
bkYfiu1crmnjjawBoaGC8S/SIEW2yijKUnPIGfxsde5jMuLwCVyLrYR8dH+c/a8E
H9ctqJFM9gmiJGRGH8zSBfMe0op+mE0VdxmfxxGh009d4NlJPvsKu3lwD44xerLd
KZ798VJjrZYfZyLa1zripFZ3zKq3IA+JGID15Qgx3EzRXqffKa2CIW5wlnUM1F2h
aN/ySoOkAJm4LOnc3o4CB/DdH4toMninIbxL5KMehG/T4cXggwEmU4P61CBPGO1q
fcOPhp3Diood3G4CDGeiQhYQ+fncHlA0DBYlmtGu6x536ae3uagQM9hlMBJ0Q9jI
gl0VAuu6lXV9bOQ90C/csfU8zvNSZqcwyj7L9AR9VnMKVzA+7tv60/sriduZ8F/5
0qnkI/FDxIFQiJG6uXcGUtyh3YbHd7jp/SUufZUSrnR8OuKMDDTpss0M16f4IzT/
cHSDHbO4HMc/F8yVBTAaz10u6nn7nj7BXaVCVWiIeB8+uVgfAGLHGJjDApgUrwYF
EX803ihIgdYv9pA4k3uT69aqZBcoRck/3r6dLjRrBjVuEudQoBghlsjgY5rGpAXo
j4MiAsxzl3h0PC1NSEAMq8BDSiL9ShOGdd1z/AHFXUkrAf4WpJGvazz5u9JNj1ar
PhP89WGpodOY639xDdQ3bXbR4NzWAUpCcLL0cUUZ92882fMbtKWZNxVmB/p/YGPL
YJj10CyQjvPRlYAf7NL5urESKd1t9dRixgwUjdf2i6lzg0rUFIA8oYW48UlyrEdw
zFyTx+PblIz16JVSlMB0vw==
`protect END_PROTECTED
